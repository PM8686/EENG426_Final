magic
tech sky130l
timestamp 1731220651
<< m1 >>
rect 2048 2447 2052 2475
rect 504 2359 508 2387
rect 576 2359 580 2387
rect 648 2359 652 2387
rect 928 2359 932 2387
rect 1488 2363 1492 2391
rect 1536 2363 1540 2391
rect 1592 2363 1596 2391
rect 1648 2363 1652 2391
rect 1768 2363 1772 2391
rect 1832 2363 1836 2391
rect 1904 2363 1908 2391
rect 2080 2363 2084 2391
rect 2392 2339 2396 2391
rect 760 2211 764 2239
rect 920 2211 924 2239
rect 1368 2223 1372 2251
rect 1440 2223 1444 2251
rect 1664 2223 1668 2251
rect 1736 2223 1740 2251
rect 1872 2223 1876 2251
rect 1944 2223 1948 2251
rect 2024 2223 2028 2251
rect 2112 2223 2116 2251
rect 2208 2223 2212 2251
rect 264 2099 268 2187
rect 552 2159 556 2191
rect 256 2067 260 2095
rect 376 2067 380 2095
rect 584 2067 588 2155
rect 768 2067 772 2095
rect 824 2067 828 2095
rect 872 2067 876 2095
rect 920 2067 924 2095
rect 968 2067 972 2095
rect 1024 2067 1028 2095
rect 1472 2079 1476 2107
rect 1528 2079 1532 2107
rect 1600 2079 1604 2107
rect 1680 2079 1684 2107
rect 1768 2079 1772 2107
rect 2032 2079 2036 2107
rect 2136 2079 2140 2107
rect 2208 2079 2212 2107
rect 664 2011 668 2039
rect 248 1927 252 1955
rect 304 1927 308 1955
rect 376 1927 380 1955
rect 1952 1943 1956 1971
rect 2128 1943 2132 1971
rect 2176 1943 2180 1971
rect 552 1783 556 1811
rect 600 1783 604 1811
rect 656 1783 660 1811
rect 792 1783 796 1811
rect 1008 1783 1012 1811
rect 1432 1795 1436 1823
rect 1480 1795 1484 1823
rect 1536 1795 1540 1823
rect 1592 1795 1596 1823
rect 1704 1795 1708 1883
rect 1928 1795 1932 1823
rect 480 1643 484 1671
rect 528 1643 532 1671
rect 624 1643 628 1671
rect 872 1643 876 1671
rect 1536 1643 1540 1671
rect 1592 1643 1596 1671
rect 1656 1643 1660 1671
rect 1840 1643 1844 1671
rect 1896 1643 1900 1727
rect 2008 1643 2012 1671
rect 2064 1643 2068 1671
rect 168 1587 172 1603
rect 1664 1595 1668 1639
rect 232 1499 236 1527
rect 296 1499 300 1527
rect 376 1499 380 1527
rect 472 1499 476 1527
rect 568 1499 572 1527
rect 768 1499 772 1527
rect 856 1499 860 1527
rect 1792 1503 1796 1531
rect 1904 1503 1908 1531
rect 1136 1443 1140 1471
rect 1856 1439 1860 1459
rect 656 1355 660 1383
rect 720 1355 724 1383
rect 784 1355 788 1383
rect 1376 1347 1380 1375
rect 1584 1347 1588 1375
rect 1672 1347 1676 1375
rect 1936 1347 1940 1375
rect 2024 1347 2028 1375
rect 2184 1347 2188 1375
rect 2344 1347 2348 1427
rect 296 1211 300 1239
rect 360 1211 364 1239
rect 776 1211 780 1239
rect 1824 1203 1828 1231
rect 1872 1203 1876 1231
rect 1936 1203 1940 1231
rect 2072 1203 2076 1231
rect 2328 1203 2332 1231
rect 168 1067 172 1095
rect 248 1067 252 1095
rect 336 1067 340 1095
rect 808 1067 812 1095
rect 872 1067 876 1095
rect 936 1067 940 1095
rect 992 1067 996 1095
rect 1120 1067 1124 1095
rect 1568 1055 1572 1083
rect 1632 1055 1636 1083
rect 1696 1055 1700 1083
rect 1824 1055 1828 1083
rect 1888 1055 1892 1083
rect 2056 1055 2060 1083
rect 2112 1055 2116 1083
rect 2288 1055 2292 1083
rect 664 1011 668 1039
rect 1968 991 1972 1019
rect 328 915 332 943
rect 376 915 380 943
rect 432 915 436 943
rect 840 915 844 943
rect 920 915 924 943
rect 992 915 996 943
rect 1120 915 1124 943
rect 1496 899 1500 987
rect 1576 899 1580 927
rect 1672 899 1676 927
rect 1768 899 1772 927
rect 2056 899 2060 927
rect 296 851 300 883
rect 576 771 580 799
rect 720 771 724 799
rect 784 771 788 799
rect 960 771 964 799
rect 1016 771 1020 799
rect 2184 783 2188 867
rect 1512 751 1516 779
rect 1656 751 1660 779
rect 1808 751 1812 779
rect 1856 751 1860 779
rect 1920 751 1924 779
rect 1984 751 1988 779
rect 2224 751 2228 779
rect 168 719 172 735
rect 264 627 268 655
rect 376 627 380 655
rect 800 627 804 655
rect 936 627 940 655
rect 1000 627 1004 655
rect 1120 627 1124 655
rect 1672 615 1676 643
rect 1720 615 1724 643
rect 1776 615 1780 643
rect 1832 615 1836 643
rect 1984 615 1988 643
rect 2216 555 2220 611
rect 2392 587 2396 643
rect 184 487 188 515
rect 384 487 388 515
rect 448 487 452 515
rect 512 487 516 515
rect 728 487 732 515
rect 1032 487 1036 515
rect 1520 471 1524 499
rect 1568 471 1572 499
rect 1624 471 1628 499
rect 1680 471 1684 499
rect 2056 471 2060 499
rect 368 347 372 375
rect 432 347 436 375
rect 952 347 956 375
rect 1008 347 1012 375
rect 1640 335 1644 363
rect 1952 335 1956 363
rect 1544 275 1548 291
rect 344 195 348 223
rect 424 195 428 223
rect 496 195 500 223
rect 560 195 564 223
rect 624 195 628 223
rect 768 195 772 223
rect 816 195 820 223
rect 864 195 868 223
rect 912 195 916 223
rect 960 195 964 223
rect 1008 195 1012 223
rect 1440 187 1444 215
rect 1488 187 1492 215
rect 1544 187 1548 215
rect 1600 187 1604 215
rect 1664 187 1668 215
rect 1808 187 1812 215
rect 1888 187 1892 215
rect 1976 187 1980 215
rect 2064 187 2068 215
<< m2c >>
rect 256 2479 260 2483
rect 296 2479 300 2483
rect 336 2479 340 2483
rect 376 2479 380 2483
rect 424 2479 428 2483
rect 480 2479 484 2483
rect 536 2479 540 2483
rect 600 2479 604 2483
rect 664 2479 668 2483
rect 728 2479 732 2483
rect 792 2479 796 2483
rect 848 2479 852 2483
rect 904 2479 908 2483
rect 952 2479 956 2483
rect 1000 2479 1004 2483
rect 1048 2479 1052 2483
rect 1096 2479 1100 2483
rect 1136 2479 1140 2483
rect 1176 2479 1180 2483
rect 1216 2479 1220 2483
rect 1328 2475 1332 2479
rect 1368 2475 1372 2479
rect 1408 2475 1412 2479
rect 1464 2475 1468 2479
rect 1536 2475 1540 2479
rect 1608 2475 1612 2479
rect 1688 2475 1692 2479
rect 1760 2475 1764 2479
rect 1832 2475 1836 2479
rect 1912 2475 1916 2479
rect 1992 2475 1996 2479
rect 2048 2475 2052 2479
rect 2088 2475 2092 2479
rect 2192 2475 2196 2479
rect 2296 2475 2300 2479
rect 256 2447 260 2451
rect 296 2447 300 2451
rect 336 2447 340 2451
rect 376 2447 380 2451
rect 424 2447 428 2451
rect 480 2447 484 2451
rect 536 2447 540 2451
rect 600 2447 604 2451
rect 664 2447 668 2451
rect 728 2447 732 2451
rect 792 2447 796 2451
rect 848 2447 852 2451
rect 904 2447 908 2451
rect 952 2447 956 2451
rect 1000 2447 1004 2451
rect 1048 2447 1052 2451
rect 1096 2447 1100 2451
rect 1136 2447 1140 2451
rect 1176 2447 1180 2451
rect 1216 2447 1220 2451
rect 1328 2443 1332 2447
rect 1368 2443 1372 2447
rect 1408 2443 1412 2447
rect 1464 2443 1468 2447
rect 1536 2443 1540 2447
rect 1608 2443 1612 2447
rect 1688 2443 1692 2447
rect 1760 2443 1764 2447
rect 1832 2443 1836 2447
rect 1912 2443 1916 2447
rect 1992 2443 1996 2447
rect 2048 2443 2052 2447
rect 2088 2443 2092 2447
rect 2192 2443 2196 2447
rect 2296 2443 2300 2447
rect 2384 2443 2388 2447
rect 1400 2391 1404 2395
rect 1440 2391 1444 2395
rect 1480 2391 1484 2395
rect 1488 2391 1492 2395
rect 1528 2391 1532 2395
rect 1536 2391 1540 2395
rect 1584 2391 1588 2395
rect 1592 2391 1596 2395
rect 1640 2391 1644 2395
rect 1648 2391 1652 2395
rect 1704 2391 1708 2395
rect 1760 2391 1764 2395
rect 1768 2391 1772 2395
rect 1824 2391 1828 2395
rect 1832 2391 1836 2395
rect 1896 2391 1900 2395
rect 1904 2391 1908 2395
rect 1976 2391 1980 2395
rect 2072 2391 2076 2395
rect 2080 2391 2084 2395
rect 2176 2391 2180 2395
rect 2288 2391 2292 2395
rect 2384 2391 2388 2395
rect 2392 2391 2396 2395
rect 224 2387 228 2391
rect 288 2387 292 2391
rect 352 2387 356 2391
rect 424 2387 428 2391
rect 496 2387 500 2391
rect 504 2387 508 2391
rect 568 2387 572 2391
rect 576 2387 580 2391
rect 640 2387 644 2391
rect 648 2387 652 2391
rect 712 2387 716 2391
rect 776 2387 780 2391
rect 848 2387 852 2391
rect 920 2387 924 2391
rect 928 2387 932 2391
rect 992 2387 996 2391
rect 1400 2359 1404 2363
rect 1440 2359 1444 2363
rect 1480 2359 1484 2363
rect 1488 2359 1492 2363
rect 1528 2359 1532 2363
rect 1536 2359 1540 2363
rect 1584 2359 1588 2363
rect 1592 2359 1596 2363
rect 1640 2359 1644 2363
rect 1648 2359 1652 2363
rect 1704 2359 1708 2363
rect 1760 2359 1764 2363
rect 1768 2359 1772 2363
rect 1824 2359 1828 2363
rect 1832 2359 1836 2363
rect 1896 2359 1900 2363
rect 1904 2359 1908 2363
rect 1976 2359 1980 2363
rect 2072 2359 2076 2363
rect 2080 2359 2084 2363
rect 2176 2359 2180 2363
rect 2288 2359 2292 2363
rect 2384 2359 2388 2363
rect 224 2355 228 2359
rect 288 2355 292 2359
rect 352 2355 356 2359
rect 424 2355 428 2359
rect 496 2355 500 2359
rect 504 2355 508 2359
rect 568 2355 572 2359
rect 576 2355 580 2359
rect 640 2355 644 2359
rect 648 2355 652 2359
rect 712 2355 716 2359
rect 776 2355 780 2359
rect 848 2355 852 2359
rect 920 2355 924 2359
rect 928 2355 932 2359
rect 992 2355 996 2359
rect 1352 2335 1356 2339
rect 1408 2335 1412 2339
rect 1464 2335 1468 2339
rect 1528 2335 1532 2339
rect 1600 2335 1604 2339
rect 1672 2335 1676 2339
rect 1744 2335 1748 2339
rect 1824 2335 1828 2339
rect 1904 2335 1908 2339
rect 1992 2335 1996 2339
rect 2088 2335 2092 2339
rect 2192 2335 2196 2339
rect 2296 2335 2300 2339
rect 2384 2335 2388 2339
rect 2392 2335 2396 2339
rect 296 2331 300 2335
rect 352 2331 356 2335
rect 424 2331 428 2335
rect 496 2331 500 2335
rect 576 2331 580 2335
rect 656 2331 660 2335
rect 736 2331 740 2335
rect 808 2331 812 2335
rect 880 2331 884 2335
rect 944 2331 948 2335
rect 1016 2331 1020 2335
rect 1088 2331 1092 2335
rect 1352 2303 1356 2307
rect 1408 2303 1412 2307
rect 1464 2303 1468 2307
rect 1528 2303 1532 2307
rect 1600 2303 1604 2307
rect 1672 2303 1676 2307
rect 1744 2303 1748 2307
rect 1824 2303 1828 2307
rect 1904 2303 1908 2307
rect 1992 2303 1996 2307
rect 2088 2303 2092 2307
rect 2192 2303 2196 2307
rect 2296 2303 2300 2307
rect 2384 2303 2388 2307
rect 296 2299 300 2303
rect 352 2299 356 2303
rect 424 2299 428 2303
rect 496 2299 500 2303
rect 576 2299 580 2303
rect 656 2299 660 2303
rect 736 2299 740 2303
rect 808 2299 812 2303
rect 880 2299 884 2303
rect 944 2299 948 2303
rect 1016 2299 1020 2303
rect 1088 2299 1092 2303
rect 1360 2251 1364 2255
rect 1368 2251 1372 2255
rect 1432 2251 1436 2255
rect 1440 2251 1444 2255
rect 1512 2251 1516 2255
rect 1584 2251 1588 2255
rect 1656 2251 1660 2255
rect 1664 2251 1668 2255
rect 1728 2251 1732 2255
rect 1736 2251 1740 2255
rect 1800 2251 1804 2255
rect 1864 2251 1868 2255
rect 1872 2251 1876 2255
rect 1936 2251 1940 2255
rect 1944 2251 1948 2255
rect 2016 2251 2020 2255
rect 2024 2251 2028 2255
rect 2104 2251 2108 2255
rect 2112 2251 2116 2255
rect 2200 2251 2204 2255
rect 2208 2251 2212 2255
rect 2304 2251 2308 2255
rect 2384 2251 2388 2255
rect 168 2239 172 2243
rect 208 2239 212 2243
rect 248 2239 252 2243
rect 304 2239 308 2243
rect 360 2239 364 2243
rect 432 2239 436 2243
rect 504 2239 508 2243
rect 584 2239 588 2243
rect 672 2239 676 2243
rect 752 2239 756 2243
rect 760 2239 764 2243
rect 832 2239 836 2243
rect 912 2239 916 2243
rect 920 2239 924 2243
rect 992 2239 996 2243
rect 1072 2239 1076 2243
rect 1152 2239 1156 2243
rect 1360 2219 1364 2223
rect 1368 2219 1372 2223
rect 1432 2219 1436 2223
rect 1440 2219 1444 2223
rect 1512 2219 1516 2223
rect 1584 2219 1588 2223
rect 1656 2219 1660 2223
rect 1664 2219 1668 2223
rect 1728 2219 1732 2223
rect 1736 2219 1740 2223
rect 1800 2219 1804 2223
rect 1864 2219 1868 2223
rect 1872 2219 1876 2223
rect 1936 2219 1940 2223
rect 1944 2219 1948 2223
rect 2016 2219 2020 2223
rect 2024 2219 2028 2223
rect 2104 2219 2108 2223
rect 2112 2219 2116 2223
rect 2200 2219 2204 2223
rect 2208 2219 2212 2223
rect 2304 2219 2308 2223
rect 2384 2219 2388 2223
rect 168 2207 172 2211
rect 208 2207 212 2211
rect 248 2207 252 2211
rect 304 2207 308 2211
rect 360 2207 364 2211
rect 432 2207 436 2211
rect 504 2207 508 2211
rect 584 2207 588 2211
rect 672 2207 676 2211
rect 752 2207 756 2211
rect 760 2207 764 2211
rect 832 2207 836 2211
rect 912 2207 916 2211
rect 920 2207 924 2211
rect 992 2209 996 2213
rect 1072 2207 1076 2211
rect 1152 2207 1156 2211
rect 552 2191 556 2195
rect 1400 2191 1404 2195
rect 1464 2191 1468 2195
rect 1536 2191 1540 2195
rect 1616 2191 1620 2195
rect 1696 2191 1700 2195
rect 1776 2191 1780 2195
rect 1856 2191 1860 2195
rect 1928 2191 1932 2195
rect 1992 2191 1996 2195
rect 2056 2191 2060 2195
rect 2120 2191 2124 2195
rect 2192 2191 2196 2195
rect 2264 2191 2268 2195
rect 2336 2191 2340 2195
rect 2384 2191 2388 2195
rect 160 2187 164 2191
rect 232 2187 236 2191
rect 264 2187 268 2191
rect 304 2187 308 2191
rect 384 2187 388 2191
rect 464 2187 468 2191
rect 544 2187 548 2191
rect 160 2155 164 2159
rect 232 2155 236 2159
rect 624 2187 628 2191
rect 704 2187 708 2191
rect 784 2187 788 2191
rect 856 2187 860 2191
rect 928 2187 932 2191
rect 1000 2187 1004 2191
rect 1072 2187 1076 2191
rect 1144 2187 1148 2191
rect 1400 2159 1404 2163
rect 1464 2159 1468 2163
rect 1536 2159 1540 2163
rect 1616 2159 1620 2163
rect 1696 2159 1700 2163
rect 1776 2159 1780 2163
rect 1856 2159 1860 2163
rect 1928 2159 1932 2163
rect 1992 2159 1996 2163
rect 2056 2159 2060 2163
rect 2120 2159 2124 2163
rect 2192 2159 2196 2163
rect 2264 2159 2268 2163
rect 2336 2159 2340 2163
rect 2384 2159 2388 2163
rect 304 2155 308 2159
rect 384 2155 388 2159
rect 464 2155 468 2159
rect 544 2155 548 2159
rect 552 2155 556 2159
rect 584 2155 588 2159
rect 624 2155 628 2159
rect 704 2155 708 2159
rect 784 2155 788 2159
rect 856 2155 860 2159
rect 928 2155 932 2159
rect 1000 2155 1004 2159
rect 1072 2155 1076 2159
rect 1144 2155 1148 2159
rect 160 2095 164 2099
rect 216 2095 220 2099
rect 256 2095 260 2099
rect 264 2095 268 2099
rect 296 2095 300 2099
rect 368 2095 372 2099
rect 376 2095 380 2099
rect 440 2095 444 2099
rect 504 2095 508 2099
rect 568 2095 572 2099
rect 160 2063 164 2067
rect 216 2063 220 2067
rect 256 2063 260 2067
rect 296 2063 300 2067
rect 368 2063 372 2067
rect 376 2063 380 2067
rect 440 2065 444 2069
rect 1424 2107 1428 2111
rect 1464 2107 1468 2111
rect 1472 2107 1476 2111
rect 1520 2107 1524 2111
rect 1528 2107 1532 2111
rect 1592 2107 1596 2111
rect 1600 2107 1604 2111
rect 1672 2107 1676 2111
rect 1680 2107 1684 2111
rect 1760 2107 1764 2111
rect 1768 2107 1772 2111
rect 1848 2107 1852 2111
rect 1936 2107 1940 2111
rect 2024 2107 2028 2111
rect 2032 2107 2036 2111
rect 2112 2107 2116 2111
rect 2136 2107 2140 2111
rect 2200 2107 2204 2111
rect 2208 2107 2212 2111
rect 2296 2107 2300 2111
rect 2384 2107 2388 2111
rect 632 2095 636 2099
rect 696 2095 700 2099
rect 760 2095 764 2099
rect 768 2095 772 2099
rect 816 2095 820 2099
rect 824 2095 828 2099
rect 864 2095 868 2099
rect 872 2095 876 2099
rect 912 2095 916 2099
rect 920 2095 924 2099
rect 960 2095 964 2099
rect 968 2095 972 2099
rect 1016 2095 1020 2099
rect 1024 2095 1028 2099
rect 1072 2095 1076 2099
rect 1424 2075 1428 2079
rect 1464 2075 1468 2079
rect 1472 2075 1476 2079
rect 1520 2075 1524 2079
rect 1528 2075 1532 2079
rect 1592 2075 1596 2079
rect 1600 2075 1604 2079
rect 1672 2075 1676 2079
rect 1680 2075 1684 2079
rect 1760 2075 1764 2079
rect 1768 2075 1772 2079
rect 1848 2075 1852 2079
rect 1936 2075 1940 2079
rect 2024 2075 2028 2079
rect 2032 2075 2036 2079
rect 2112 2075 2116 2079
rect 2136 2075 2140 2079
rect 2200 2075 2204 2079
rect 2208 2075 2212 2079
rect 2296 2075 2300 2079
rect 2384 2075 2388 2079
rect 504 2063 508 2067
rect 568 2063 572 2067
rect 584 2063 588 2067
rect 632 2063 636 2067
rect 696 2063 700 2067
rect 760 2063 764 2067
rect 768 2063 772 2067
rect 816 2063 820 2067
rect 824 2063 828 2067
rect 864 2063 868 2067
rect 872 2063 876 2067
rect 912 2063 916 2067
rect 920 2063 924 2067
rect 960 2063 964 2067
rect 968 2063 972 2067
rect 1016 2063 1020 2067
rect 1024 2063 1028 2067
rect 1072 2063 1076 2067
rect 2064 2055 2068 2059
rect 2104 2055 2108 2059
rect 2144 2055 2148 2059
rect 2184 2055 2188 2059
rect 2224 2055 2228 2059
rect 2264 2055 2268 2059
rect 2304 2055 2308 2059
rect 2344 2055 2348 2059
rect 2384 2055 2388 2059
rect 160 2039 164 2043
rect 200 2039 204 2043
rect 240 2039 244 2043
rect 304 2039 308 2043
rect 376 2039 380 2043
rect 448 2039 452 2043
rect 512 2039 516 2043
rect 576 2039 580 2043
rect 640 2039 644 2043
rect 664 2039 668 2043
rect 704 2039 708 2043
rect 768 2039 772 2043
rect 840 2039 844 2043
rect 2064 2023 2068 2027
rect 2104 2023 2108 2027
rect 2144 2023 2148 2027
rect 2184 2023 2188 2027
rect 2224 2023 2228 2027
rect 2264 2023 2268 2027
rect 2304 2023 2308 2027
rect 2344 2023 2348 2027
rect 2384 2023 2388 2027
rect 160 2007 164 2011
rect 200 2007 204 2011
rect 240 2007 244 2011
rect 304 2007 308 2011
rect 376 2007 380 2011
rect 448 2007 452 2011
rect 512 2007 516 2011
rect 576 2007 580 2011
rect 640 2007 644 2011
rect 664 2007 668 2011
rect 704 2007 708 2011
rect 768 2007 772 2011
rect 840 2007 844 2011
rect 1424 1971 1428 1975
rect 1464 1971 1468 1975
rect 1504 1971 1508 1975
rect 1544 1971 1548 1975
rect 1584 1971 1588 1975
rect 1624 1971 1628 1975
rect 1664 1971 1668 1975
rect 1704 1971 1708 1975
rect 1744 1971 1748 1975
rect 1792 1971 1796 1975
rect 1848 1971 1852 1975
rect 1896 1971 1900 1975
rect 1944 1971 1948 1975
rect 1952 1971 1956 1975
rect 1992 1971 1996 1975
rect 2040 1971 2044 1975
rect 2080 1971 2084 1975
rect 2120 1971 2124 1975
rect 2128 1971 2132 1975
rect 2168 1971 2172 1975
rect 2176 1971 2180 1975
rect 2216 1971 2220 1975
rect 2264 1971 2268 1975
rect 2304 1971 2308 1975
rect 2344 1971 2348 1975
rect 2384 1971 2388 1975
rect 160 1955 164 1959
rect 200 1955 204 1959
rect 240 1955 244 1959
rect 248 1955 252 1959
rect 296 1955 300 1959
rect 304 1955 308 1959
rect 368 1955 372 1959
rect 376 1955 380 1959
rect 440 1955 444 1959
rect 520 1955 524 1959
rect 600 1955 604 1959
rect 672 1955 676 1959
rect 744 1955 748 1959
rect 816 1955 820 1959
rect 888 1955 892 1959
rect 960 1955 964 1959
rect 1032 1955 1036 1959
rect 1424 1939 1428 1943
rect 1464 1939 1468 1943
rect 1504 1939 1508 1943
rect 1544 1939 1548 1943
rect 1584 1939 1588 1943
rect 1624 1939 1628 1943
rect 1664 1939 1668 1943
rect 1704 1939 1708 1943
rect 1744 1939 1748 1943
rect 1792 1939 1796 1943
rect 1848 1939 1852 1943
rect 1896 1939 1900 1943
rect 1944 1939 1948 1943
rect 1952 1939 1956 1943
rect 1992 1939 1996 1943
rect 2040 1939 2044 1943
rect 2080 1939 2084 1943
rect 2120 1939 2124 1943
rect 2128 1939 2132 1943
rect 2168 1939 2172 1943
rect 2176 1939 2180 1943
rect 2216 1939 2220 1943
rect 2264 1939 2268 1943
rect 2304 1939 2308 1943
rect 2344 1939 2348 1943
rect 2384 1939 2388 1943
rect 160 1923 164 1927
rect 200 1923 204 1927
rect 240 1923 244 1927
rect 248 1923 252 1927
rect 296 1923 300 1927
rect 304 1923 308 1927
rect 368 1923 372 1927
rect 376 1923 380 1927
rect 440 1923 444 1927
rect 520 1923 524 1927
rect 600 1923 604 1927
rect 672 1923 676 1927
rect 744 1923 748 1927
rect 816 1923 820 1927
rect 888 1923 892 1927
rect 960 1923 964 1927
rect 1032 1923 1036 1927
rect 1368 1915 1372 1919
rect 1408 1915 1412 1919
rect 1448 1915 1452 1919
rect 1488 1915 1492 1919
rect 1536 1915 1540 1919
rect 1592 1915 1596 1919
rect 1656 1915 1660 1919
rect 1736 1915 1740 1919
rect 1832 1915 1836 1919
rect 1944 1915 1948 1919
rect 2056 1915 2060 1919
rect 2176 1915 2180 1919
rect 272 1899 276 1903
rect 312 1899 316 1903
rect 352 1899 356 1903
rect 392 1899 396 1903
rect 440 1899 444 1903
rect 496 1899 500 1903
rect 560 1899 564 1903
rect 624 1899 628 1903
rect 688 1899 692 1903
rect 752 1899 756 1903
rect 816 1899 820 1903
rect 880 1899 884 1903
rect 944 1899 948 1903
rect 1008 1901 1012 1905
rect 1080 1899 1084 1903
rect 1152 1899 1156 1903
rect 1368 1883 1372 1887
rect 1408 1883 1412 1887
rect 1448 1883 1452 1887
rect 1488 1883 1492 1887
rect 1536 1883 1540 1887
rect 1592 1883 1596 1887
rect 1656 1883 1660 1887
rect 1704 1883 1708 1887
rect 1736 1883 1740 1887
rect 1832 1883 1836 1887
rect 1944 1883 1948 1887
rect 2056 1883 2060 1887
rect 2176 1883 2180 1887
rect 272 1869 276 1873
rect 312 1867 316 1871
rect 352 1867 356 1871
rect 392 1867 396 1871
rect 440 1867 444 1871
rect 496 1867 500 1871
rect 560 1867 564 1871
rect 624 1867 628 1871
rect 688 1867 692 1871
rect 752 1867 756 1871
rect 816 1867 820 1871
rect 880 1867 884 1871
rect 944 1867 948 1871
rect 1008 1867 1012 1871
rect 1080 1867 1084 1871
rect 1152 1867 1156 1871
rect 1384 1823 1388 1827
rect 1424 1823 1428 1827
rect 1432 1823 1436 1827
rect 1472 1823 1476 1827
rect 1480 1823 1484 1827
rect 1528 1823 1532 1827
rect 1536 1823 1540 1827
rect 1584 1823 1588 1827
rect 1592 1823 1596 1827
rect 1640 1823 1644 1827
rect 1696 1823 1700 1827
rect 424 1811 428 1815
rect 464 1811 468 1815
rect 504 1811 508 1815
rect 544 1811 548 1815
rect 552 1811 556 1815
rect 592 1811 596 1815
rect 600 1811 604 1815
rect 648 1811 652 1815
rect 656 1811 660 1815
rect 712 1811 716 1815
rect 784 1811 788 1815
rect 792 1811 796 1815
rect 856 1811 860 1815
rect 928 1811 932 1815
rect 1000 1811 1004 1815
rect 1008 1811 1012 1815
rect 1072 1811 1076 1815
rect 1152 1811 1156 1815
rect 1216 1811 1220 1815
rect 424 1779 428 1783
rect 464 1779 468 1783
rect 504 1779 508 1783
rect 544 1779 548 1783
rect 552 1779 556 1783
rect 592 1779 596 1783
rect 600 1779 604 1783
rect 648 1779 652 1783
rect 656 1779 660 1783
rect 712 1779 716 1783
rect 784 1779 788 1783
rect 792 1779 796 1783
rect 856 1781 860 1785
rect 1752 1823 1756 1827
rect 1808 1823 1812 1827
rect 1864 1823 1868 1827
rect 1920 1823 1924 1827
rect 1928 1823 1932 1827
rect 1976 1823 1980 1827
rect 1384 1791 1388 1795
rect 1424 1791 1428 1795
rect 1432 1791 1436 1795
rect 1472 1791 1476 1795
rect 1480 1791 1484 1795
rect 1528 1791 1532 1795
rect 1536 1791 1540 1795
rect 1584 1791 1588 1795
rect 1592 1791 1596 1795
rect 1640 1791 1644 1795
rect 1696 1791 1700 1795
rect 1704 1791 1708 1795
rect 1752 1791 1756 1795
rect 1808 1791 1812 1795
rect 1864 1791 1868 1795
rect 1920 1791 1924 1795
rect 1928 1791 1932 1795
rect 1976 1791 1980 1795
rect 928 1779 932 1783
rect 1000 1779 1004 1783
rect 1008 1779 1012 1783
rect 1072 1779 1076 1783
rect 1152 1779 1156 1783
rect 1216 1779 1220 1783
rect 432 1759 436 1763
rect 472 1759 476 1763
rect 512 1759 516 1763
rect 552 1759 556 1763
rect 592 1759 596 1763
rect 632 1759 636 1763
rect 672 1759 676 1763
rect 720 1759 724 1763
rect 776 1759 780 1763
rect 832 1759 836 1763
rect 896 1759 900 1763
rect 960 1759 964 1763
rect 1024 1759 1028 1763
rect 1096 1759 1100 1763
rect 1168 1759 1172 1763
rect 1216 1759 1220 1763
rect 1328 1759 1332 1763
rect 1368 1759 1372 1763
rect 1416 1759 1420 1763
rect 1480 1759 1484 1763
rect 1544 1759 1548 1763
rect 1608 1759 1612 1763
rect 1672 1759 1676 1763
rect 1728 1759 1732 1763
rect 1784 1759 1788 1763
rect 1832 1759 1836 1763
rect 1888 1759 1892 1763
rect 1944 1759 1948 1763
rect 2000 1759 2004 1763
rect 432 1727 436 1731
rect 472 1727 476 1731
rect 512 1727 516 1731
rect 552 1727 556 1731
rect 592 1727 596 1731
rect 632 1727 636 1731
rect 672 1727 676 1731
rect 720 1727 724 1731
rect 776 1727 780 1731
rect 832 1727 836 1731
rect 896 1727 900 1731
rect 960 1727 964 1731
rect 1024 1727 1028 1731
rect 1096 1727 1100 1731
rect 1168 1727 1172 1731
rect 1216 1727 1220 1731
rect 1328 1727 1332 1731
rect 1368 1727 1372 1731
rect 1416 1727 1420 1731
rect 1480 1727 1484 1731
rect 1544 1727 1548 1731
rect 1608 1727 1612 1731
rect 1672 1727 1676 1731
rect 1728 1727 1732 1731
rect 1784 1727 1788 1731
rect 1832 1727 1836 1731
rect 1888 1727 1892 1731
rect 1896 1727 1900 1731
rect 1944 1727 1948 1731
rect 2000 1727 2004 1731
rect 304 1671 308 1675
rect 344 1671 348 1675
rect 384 1671 388 1675
rect 424 1671 428 1675
rect 472 1671 476 1675
rect 480 1671 484 1675
rect 520 1671 524 1675
rect 528 1671 532 1675
rect 568 1671 572 1675
rect 616 1671 620 1675
rect 624 1671 628 1675
rect 664 1671 668 1675
rect 712 1671 716 1675
rect 760 1671 764 1675
rect 808 1671 812 1675
rect 864 1671 868 1675
rect 872 1671 876 1675
rect 920 1671 924 1675
rect 1328 1671 1332 1675
rect 1368 1671 1372 1675
rect 1408 1671 1412 1675
rect 1448 1671 1452 1675
rect 1488 1671 1492 1675
rect 1528 1671 1532 1675
rect 1536 1671 1540 1675
rect 1584 1671 1588 1675
rect 1592 1671 1596 1675
rect 1648 1671 1652 1675
rect 1656 1671 1660 1675
rect 1712 1671 1716 1675
rect 1776 1671 1780 1675
rect 1832 1671 1836 1675
rect 1840 1671 1844 1675
rect 1888 1671 1892 1675
rect 1944 1671 1948 1675
rect 2000 1671 2004 1675
rect 2008 1671 2012 1675
rect 2056 1671 2060 1675
rect 2064 1671 2068 1675
rect 2112 1671 2116 1675
rect 304 1639 308 1643
rect 344 1639 348 1643
rect 384 1639 388 1643
rect 424 1639 428 1643
rect 472 1639 476 1643
rect 480 1639 484 1643
rect 520 1639 524 1643
rect 528 1639 532 1643
rect 568 1639 572 1643
rect 616 1639 620 1643
rect 624 1639 628 1643
rect 664 1639 668 1643
rect 712 1639 716 1643
rect 760 1639 764 1643
rect 808 1639 812 1643
rect 864 1639 868 1643
rect 872 1639 876 1643
rect 920 1639 924 1643
rect 1328 1639 1332 1643
rect 1368 1639 1372 1643
rect 1408 1639 1412 1643
rect 1448 1639 1452 1643
rect 1488 1639 1492 1643
rect 1528 1639 1532 1643
rect 1536 1639 1540 1643
rect 1584 1639 1588 1643
rect 1592 1639 1596 1643
rect 1648 1639 1652 1643
rect 1656 1639 1660 1643
rect 1664 1639 1668 1643
rect 1712 1639 1716 1643
rect 1776 1639 1780 1643
rect 1832 1639 1836 1643
rect 1840 1639 1844 1643
rect 1888 1639 1892 1643
rect 1896 1639 1900 1643
rect 1944 1639 1948 1643
rect 2000 1639 2004 1643
rect 2008 1639 2012 1643
rect 2056 1639 2060 1643
rect 2064 1639 2068 1643
rect 2112 1639 2116 1643
rect 160 1615 164 1619
rect 200 1615 204 1619
rect 240 1615 244 1619
rect 280 1615 284 1619
rect 336 1615 340 1619
rect 416 1615 420 1619
rect 496 1615 500 1619
rect 584 1615 588 1619
rect 664 1615 668 1619
rect 744 1615 748 1619
rect 816 1615 820 1619
rect 880 1615 884 1619
rect 944 1615 948 1619
rect 1008 1615 1012 1619
rect 1072 1615 1076 1619
rect 1328 1615 1332 1619
rect 1368 1615 1372 1619
rect 1408 1617 1412 1621
rect 1448 1615 1452 1619
rect 1488 1615 1492 1619
rect 1528 1615 1532 1619
rect 1584 1615 1588 1619
rect 1656 1615 1660 1619
rect 168 1603 172 1607
rect 1728 1615 1732 1619
rect 1808 1615 1812 1619
rect 1880 1615 1884 1619
rect 1952 1615 1956 1619
rect 2024 1615 2028 1619
rect 2088 1615 2092 1619
rect 2152 1615 2156 1619
rect 2216 1615 2220 1619
rect 2280 1615 2284 1619
rect 2344 1615 2348 1619
rect 2384 1615 2388 1619
rect 1664 1591 1668 1595
rect 160 1583 164 1587
rect 168 1583 172 1587
rect 200 1583 204 1587
rect 240 1583 244 1587
rect 280 1583 284 1587
rect 336 1583 340 1587
rect 416 1583 420 1587
rect 496 1583 500 1587
rect 584 1583 588 1587
rect 664 1583 668 1587
rect 744 1583 748 1587
rect 816 1583 820 1587
rect 880 1583 884 1587
rect 944 1583 948 1587
rect 1008 1583 1012 1587
rect 1072 1583 1076 1587
rect 1328 1583 1332 1587
rect 1368 1583 1372 1587
rect 1408 1583 1412 1587
rect 1448 1583 1452 1587
rect 1488 1583 1492 1587
rect 1528 1583 1532 1587
rect 1584 1583 1588 1587
rect 1656 1583 1660 1587
rect 1728 1583 1732 1587
rect 1808 1583 1812 1587
rect 1880 1583 1884 1587
rect 1952 1583 1956 1587
rect 2024 1583 2028 1587
rect 2088 1583 2092 1587
rect 2152 1583 2156 1587
rect 2216 1583 2220 1587
rect 2280 1583 2284 1587
rect 2344 1583 2348 1587
rect 2384 1583 2388 1587
rect 1496 1531 1500 1535
rect 1648 1531 1652 1535
rect 1784 1531 1788 1535
rect 1792 1531 1796 1535
rect 1896 1531 1900 1535
rect 1904 1531 1908 1535
rect 1992 1531 1996 1535
rect 2080 1531 2084 1535
rect 2152 1531 2156 1535
rect 2216 1531 2220 1535
rect 2280 1531 2284 1535
rect 2344 1531 2348 1535
rect 2384 1531 2388 1535
rect 176 1527 180 1531
rect 224 1527 228 1531
rect 232 1527 236 1531
rect 288 1527 292 1531
rect 296 1527 300 1531
rect 368 1527 372 1531
rect 376 1527 380 1531
rect 464 1527 468 1531
rect 472 1527 476 1531
rect 560 1527 564 1531
rect 568 1527 572 1531
rect 664 1527 668 1531
rect 760 1527 764 1531
rect 768 1527 772 1531
rect 848 1527 852 1531
rect 856 1527 860 1531
rect 928 1527 932 1531
rect 1000 1527 1004 1531
rect 1072 1527 1076 1531
rect 1144 1527 1148 1531
rect 1216 1527 1220 1531
rect 1496 1499 1500 1503
rect 1648 1499 1652 1503
rect 1784 1499 1788 1503
rect 1792 1499 1796 1503
rect 1896 1499 1900 1503
rect 1904 1499 1908 1503
rect 1992 1499 1996 1503
rect 2080 1499 2084 1503
rect 2152 1499 2156 1503
rect 2216 1499 2220 1503
rect 2280 1499 2284 1503
rect 2344 1499 2348 1503
rect 2384 1499 2388 1503
rect 176 1495 180 1499
rect 224 1495 228 1499
rect 232 1495 236 1499
rect 288 1495 292 1499
rect 296 1495 300 1499
rect 368 1495 372 1499
rect 376 1495 380 1499
rect 464 1495 468 1499
rect 472 1495 476 1499
rect 560 1495 564 1499
rect 568 1495 572 1499
rect 664 1495 668 1499
rect 760 1495 764 1499
rect 768 1495 772 1499
rect 848 1495 852 1499
rect 856 1495 860 1499
rect 928 1495 932 1499
rect 1000 1495 1004 1499
rect 1072 1495 1076 1499
rect 1144 1495 1148 1499
rect 1216 1495 1220 1499
rect 344 1471 348 1475
rect 384 1471 388 1475
rect 424 1471 428 1475
rect 472 1471 476 1475
rect 528 1471 532 1475
rect 584 1471 588 1475
rect 640 1471 644 1475
rect 696 1471 700 1475
rect 760 1471 764 1475
rect 824 1471 828 1475
rect 880 1471 884 1475
rect 936 1471 940 1475
rect 992 1471 996 1475
rect 1048 1471 1052 1475
rect 1112 1471 1116 1475
rect 1136 1471 1140 1475
rect 1176 1471 1180 1475
rect 1216 1471 1220 1475
rect 1328 1459 1332 1463
rect 1400 1459 1404 1463
rect 1504 1459 1508 1463
rect 1608 1459 1612 1463
rect 1712 1459 1716 1463
rect 1808 1459 1812 1463
rect 1856 1459 1860 1463
rect 1896 1459 1900 1463
rect 1976 1459 1980 1463
rect 2056 1459 2060 1463
rect 2128 1459 2132 1463
rect 2192 1459 2196 1463
rect 2264 1459 2268 1463
rect 2336 1459 2340 1463
rect 2384 1459 2388 1463
rect 344 1439 348 1443
rect 384 1439 388 1443
rect 424 1439 428 1443
rect 472 1439 476 1443
rect 528 1439 532 1443
rect 584 1439 588 1443
rect 640 1439 644 1443
rect 696 1439 700 1443
rect 760 1439 764 1443
rect 824 1439 828 1443
rect 880 1439 884 1443
rect 936 1439 940 1443
rect 992 1439 996 1443
rect 1048 1439 1052 1443
rect 1112 1439 1116 1443
rect 1136 1439 1140 1443
rect 1176 1439 1180 1443
rect 1216 1439 1220 1443
rect 1856 1435 1860 1439
rect 1328 1427 1332 1431
rect 1400 1427 1404 1431
rect 1504 1427 1508 1431
rect 1608 1427 1612 1431
rect 1712 1427 1716 1431
rect 1808 1427 1812 1431
rect 1896 1429 1900 1433
rect 1976 1427 1980 1431
rect 2056 1427 2060 1431
rect 2128 1427 2132 1431
rect 2192 1427 2196 1431
rect 2264 1427 2268 1431
rect 2336 1427 2340 1431
rect 2344 1427 2348 1431
rect 2384 1427 2388 1431
rect 288 1383 292 1387
rect 328 1383 332 1387
rect 368 1383 372 1387
rect 416 1383 420 1387
rect 472 1383 476 1387
rect 528 1383 532 1387
rect 584 1383 588 1387
rect 648 1383 652 1387
rect 656 1383 660 1387
rect 712 1383 716 1387
rect 720 1383 724 1387
rect 776 1383 780 1387
rect 784 1383 788 1387
rect 840 1383 844 1387
rect 904 1383 908 1387
rect 976 1383 980 1387
rect 1048 1383 1052 1387
rect 1328 1375 1332 1379
rect 1368 1375 1372 1379
rect 1376 1375 1380 1379
rect 1424 1375 1428 1379
rect 1496 1375 1500 1379
rect 1576 1375 1580 1379
rect 1584 1375 1588 1379
rect 1664 1375 1668 1379
rect 1672 1375 1676 1379
rect 1752 1375 1756 1379
rect 1840 1375 1844 1379
rect 1928 1375 1932 1379
rect 1936 1375 1940 1379
rect 2016 1375 2020 1379
rect 2024 1375 2028 1379
rect 2096 1375 2100 1379
rect 2176 1375 2180 1379
rect 2184 1375 2188 1379
rect 2248 1375 2252 1379
rect 2328 1375 2332 1379
rect 288 1351 292 1355
rect 328 1351 332 1355
rect 368 1351 372 1355
rect 416 1351 420 1355
rect 472 1351 476 1355
rect 528 1351 532 1355
rect 584 1351 588 1355
rect 648 1351 652 1355
rect 656 1351 660 1355
rect 712 1351 716 1355
rect 720 1351 724 1355
rect 776 1351 780 1355
rect 784 1351 788 1355
rect 840 1351 844 1355
rect 904 1351 908 1355
rect 976 1351 980 1355
rect 1048 1351 1052 1355
rect 2384 1375 2388 1379
rect 1328 1343 1332 1347
rect 1368 1343 1372 1347
rect 1376 1343 1380 1347
rect 1424 1343 1428 1347
rect 1496 1343 1500 1347
rect 1576 1343 1580 1347
rect 1584 1343 1588 1347
rect 1664 1343 1668 1347
rect 1672 1343 1676 1347
rect 1752 1343 1756 1347
rect 1840 1343 1844 1347
rect 1928 1343 1932 1347
rect 1936 1343 1940 1347
rect 2016 1343 2020 1347
rect 2024 1343 2028 1347
rect 2096 1343 2100 1347
rect 2176 1343 2180 1347
rect 2184 1343 2188 1347
rect 2248 1343 2252 1347
rect 2328 1343 2332 1347
rect 2344 1343 2348 1347
rect 2384 1343 2388 1347
rect 160 1327 164 1331
rect 200 1327 204 1331
rect 240 1327 244 1331
rect 280 1327 284 1331
rect 352 1327 356 1331
rect 432 1327 436 1331
rect 520 1327 524 1331
rect 608 1327 612 1331
rect 696 1327 700 1331
rect 784 1327 788 1331
rect 864 1327 868 1331
rect 944 1327 948 1331
rect 1032 1327 1036 1331
rect 1120 1327 1124 1331
rect 1472 1319 1476 1323
rect 1512 1319 1516 1323
rect 1552 1321 1556 1325
rect 1592 1319 1596 1323
rect 1640 1319 1644 1323
rect 1696 1319 1700 1323
rect 1744 1319 1748 1323
rect 1800 1319 1804 1323
rect 1856 1319 1860 1323
rect 1928 1319 1932 1323
rect 2008 1319 2012 1323
rect 2096 1319 2100 1323
rect 2192 1319 2196 1323
rect 2296 1319 2300 1323
rect 2384 1319 2388 1323
rect 160 1295 164 1299
rect 200 1295 204 1299
rect 240 1295 244 1299
rect 280 1295 284 1299
rect 352 1295 356 1299
rect 432 1295 436 1299
rect 520 1295 524 1299
rect 608 1295 612 1299
rect 696 1295 700 1299
rect 784 1295 788 1299
rect 864 1295 868 1299
rect 944 1295 948 1299
rect 1032 1295 1036 1299
rect 1120 1295 1124 1299
rect 1472 1287 1476 1291
rect 1512 1287 1516 1291
rect 1552 1287 1556 1291
rect 1592 1287 1596 1291
rect 1640 1287 1644 1291
rect 1696 1287 1700 1291
rect 1744 1287 1748 1291
rect 1800 1287 1804 1291
rect 1856 1287 1860 1291
rect 1928 1287 1932 1291
rect 2008 1287 2012 1291
rect 2096 1287 2100 1291
rect 2192 1287 2196 1291
rect 2296 1287 2300 1291
rect 2384 1287 2388 1291
rect 160 1239 164 1243
rect 200 1239 204 1243
rect 272 1239 276 1243
rect 296 1239 300 1243
rect 352 1239 356 1243
rect 360 1239 364 1243
rect 440 1239 444 1243
rect 528 1239 532 1243
rect 616 1239 620 1243
rect 696 1239 700 1243
rect 768 1239 772 1243
rect 776 1239 780 1243
rect 840 1239 844 1243
rect 904 1239 908 1243
rect 968 1239 972 1243
rect 1032 1239 1036 1243
rect 1096 1239 1100 1243
rect 1536 1231 1540 1235
rect 1576 1231 1580 1235
rect 1616 1231 1620 1235
rect 1656 1231 1660 1235
rect 1696 1231 1700 1235
rect 1736 1231 1740 1235
rect 1776 1231 1780 1235
rect 1816 1231 1820 1235
rect 1824 1231 1828 1235
rect 1864 1231 1868 1235
rect 1872 1231 1876 1235
rect 1928 1231 1932 1235
rect 1936 1231 1940 1235
rect 1992 1231 1996 1235
rect 2064 1231 2068 1235
rect 2072 1231 2076 1235
rect 2144 1231 2148 1235
rect 2232 1231 2236 1235
rect 2320 1231 2324 1235
rect 2328 1231 2332 1235
rect 2384 1231 2388 1235
rect 160 1207 164 1211
rect 200 1207 204 1211
rect 272 1207 276 1211
rect 296 1207 300 1211
rect 352 1207 356 1211
rect 360 1207 364 1211
rect 440 1207 444 1211
rect 528 1207 532 1211
rect 616 1207 620 1211
rect 696 1207 700 1211
rect 768 1207 772 1211
rect 776 1207 780 1211
rect 840 1207 844 1211
rect 904 1207 908 1211
rect 968 1207 972 1211
rect 1032 1207 1036 1211
rect 1096 1207 1100 1211
rect 1536 1199 1540 1203
rect 1576 1199 1580 1203
rect 1616 1199 1620 1203
rect 1656 1199 1660 1203
rect 1696 1199 1700 1203
rect 1736 1199 1740 1203
rect 1776 1199 1780 1203
rect 1816 1199 1820 1203
rect 1824 1199 1828 1203
rect 1864 1199 1868 1203
rect 1872 1199 1876 1203
rect 1928 1199 1932 1203
rect 1936 1199 1940 1203
rect 1992 1199 1996 1203
rect 2064 1199 2068 1203
rect 2072 1199 2076 1203
rect 2144 1199 2148 1203
rect 2232 1199 2236 1203
rect 2320 1199 2324 1203
rect 2328 1199 2332 1203
rect 2384 1199 2388 1203
rect 160 1179 164 1183
rect 200 1179 204 1183
rect 256 1179 260 1183
rect 328 1179 332 1183
rect 408 1179 412 1183
rect 496 1179 500 1183
rect 584 1179 588 1183
rect 664 1179 668 1183
rect 744 1179 748 1183
rect 824 1179 828 1183
rect 896 1179 900 1183
rect 960 1179 964 1183
rect 1016 1179 1020 1183
rect 1072 1179 1076 1183
rect 1128 1179 1132 1183
rect 1176 1179 1180 1183
rect 1216 1179 1220 1183
rect 1584 1175 1588 1179
rect 1624 1175 1628 1179
rect 1664 1175 1668 1179
rect 1704 1175 1708 1179
rect 1744 1175 1748 1179
rect 1784 1175 1788 1179
rect 1824 1175 1828 1179
rect 1880 1175 1884 1179
rect 1952 1175 1956 1179
rect 2048 1175 2052 1179
rect 2160 1175 2164 1179
rect 2280 1175 2284 1179
rect 2384 1175 2388 1179
rect 160 1147 164 1151
rect 200 1147 204 1151
rect 256 1147 260 1151
rect 328 1147 332 1151
rect 408 1147 412 1151
rect 496 1147 500 1151
rect 584 1147 588 1151
rect 664 1147 668 1151
rect 744 1147 748 1151
rect 824 1147 828 1151
rect 896 1147 900 1151
rect 960 1147 964 1151
rect 1016 1147 1020 1151
rect 1072 1147 1076 1151
rect 1128 1147 1132 1151
rect 1176 1147 1180 1151
rect 1216 1147 1220 1151
rect 1584 1143 1588 1147
rect 1624 1143 1628 1147
rect 1664 1143 1668 1147
rect 1704 1143 1708 1147
rect 1744 1143 1748 1147
rect 1784 1143 1788 1147
rect 1824 1143 1828 1147
rect 1880 1143 1884 1147
rect 1952 1143 1956 1147
rect 2048 1143 2052 1147
rect 2160 1143 2164 1147
rect 2280 1143 2284 1147
rect 2384 1143 2388 1147
rect 160 1095 164 1099
rect 168 1095 172 1099
rect 240 1095 244 1099
rect 248 1095 252 1099
rect 328 1095 332 1099
rect 336 1095 340 1099
rect 416 1095 420 1099
rect 504 1095 508 1099
rect 584 1095 588 1099
rect 664 1095 668 1099
rect 736 1095 740 1099
rect 800 1095 804 1099
rect 808 1095 812 1099
rect 864 1095 868 1099
rect 872 1095 876 1099
rect 928 1095 932 1099
rect 936 1095 940 1099
rect 984 1095 988 1099
rect 992 1095 996 1099
rect 1048 1095 1052 1099
rect 1112 1095 1116 1099
rect 1120 1095 1124 1099
rect 1176 1095 1180 1099
rect 1216 1095 1220 1099
rect 1560 1083 1564 1087
rect 1568 1083 1572 1087
rect 1624 1083 1628 1087
rect 1632 1083 1636 1087
rect 1688 1083 1692 1087
rect 1696 1083 1700 1087
rect 1752 1083 1756 1087
rect 1816 1083 1820 1087
rect 1824 1083 1828 1087
rect 1880 1083 1884 1087
rect 1888 1083 1892 1087
rect 1936 1083 1940 1087
rect 1992 1083 1996 1087
rect 2048 1083 2052 1087
rect 2056 1083 2060 1087
rect 2104 1083 2108 1087
rect 2112 1083 2116 1087
rect 2160 1083 2164 1087
rect 2216 1083 2220 1087
rect 2280 1083 2284 1087
rect 2288 1083 2292 1087
rect 2344 1083 2348 1087
rect 2384 1083 2388 1087
rect 160 1063 164 1067
rect 168 1063 172 1067
rect 240 1063 244 1067
rect 248 1063 252 1067
rect 328 1063 332 1067
rect 336 1063 340 1067
rect 416 1063 420 1067
rect 504 1063 508 1067
rect 584 1063 588 1067
rect 664 1063 668 1067
rect 736 1063 740 1067
rect 800 1063 804 1067
rect 808 1063 812 1067
rect 864 1063 868 1067
rect 872 1063 876 1067
rect 928 1063 932 1067
rect 936 1063 940 1067
rect 984 1063 988 1067
rect 992 1063 996 1067
rect 1048 1063 1052 1067
rect 1112 1063 1116 1067
rect 1120 1063 1124 1067
rect 1176 1063 1180 1067
rect 1216 1063 1220 1067
rect 1560 1051 1564 1055
rect 1568 1051 1572 1055
rect 1624 1051 1628 1055
rect 1632 1051 1636 1055
rect 1688 1051 1692 1055
rect 1696 1051 1700 1055
rect 1752 1051 1756 1055
rect 1816 1051 1820 1055
rect 1824 1051 1828 1055
rect 1880 1051 1884 1055
rect 1888 1051 1892 1055
rect 1936 1051 1940 1055
rect 1992 1051 1996 1055
rect 2048 1051 2052 1055
rect 2056 1051 2060 1055
rect 2104 1051 2108 1055
rect 2112 1051 2116 1055
rect 2160 1051 2164 1055
rect 2216 1051 2220 1055
rect 2280 1051 2284 1055
rect 2288 1051 2292 1055
rect 2344 1051 2348 1055
rect 2384 1051 2388 1055
rect 224 1039 228 1043
rect 264 1039 268 1043
rect 312 1039 316 1043
rect 368 1039 372 1043
rect 416 1039 420 1043
rect 464 1039 468 1043
rect 512 1039 516 1043
rect 560 1041 564 1045
rect 608 1039 612 1043
rect 656 1039 660 1043
rect 664 1039 668 1043
rect 704 1039 708 1043
rect 752 1039 756 1043
rect 808 1039 812 1043
rect 864 1039 868 1043
rect 920 1039 924 1043
rect 984 1039 988 1043
rect 1048 1039 1052 1043
rect 1112 1039 1116 1043
rect 1176 1039 1180 1043
rect 1216 1039 1220 1043
rect 1528 1019 1532 1023
rect 1648 1019 1652 1023
rect 1760 1019 1764 1023
rect 1856 1019 1860 1023
rect 1944 1019 1948 1023
rect 1968 1019 1972 1023
rect 2024 1021 2028 1025
rect 2096 1019 2100 1023
rect 2168 1019 2172 1023
rect 2232 1019 2236 1023
rect 2304 1019 2308 1023
rect 224 1007 228 1011
rect 264 1007 268 1011
rect 312 1007 316 1011
rect 368 1007 372 1011
rect 416 1007 420 1011
rect 464 1007 468 1011
rect 512 1007 516 1011
rect 560 1007 564 1011
rect 608 1007 612 1011
rect 656 1007 660 1011
rect 664 1007 668 1011
rect 704 1007 708 1011
rect 752 1007 756 1011
rect 808 1007 812 1011
rect 864 1007 868 1011
rect 920 1007 924 1011
rect 984 1007 988 1011
rect 1048 1007 1052 1011
rect 1112 1007 1116 1011
rect 1176 1007 1180 1011
rect 1216 1007 1220 1011
rect 1496 987 1500 991
rect 1528 987 1532 991
rect 1648 987 1652 991
rect 1760 987 1764 991
rect 1856 987 1860 991
rect 1944 987 1948 991
rect 1968 987 1972 991
rect 2024 987 2028 991
rect 2096 987 2100 991
rect 2168 987 2172 991
rect 2232 987 2236 991
rect 2304 987 2308 991
rect 320 943 324 947
rect 328 943 332 947
rect 368 943 372 947
rect 376 943 380 947
rect 424 943 428 947
rect 432 943 436 947
rect 496 943 500 947
rect 576 943 580 947
rect 664 943 668 947
rect 752 943 756 947
rect 832 943 836 947
rect 840 943 844 947
rect 912 943 916 947
rect 920 943 924 947
rect 984 943 988 947
rect 992 943 996 947
rect 1048 943 1052 947
rect 1112 943 1116 947
rect 1120 943 1124 947
rect 1176 943 1180 947
rect 1216 943 1220 947
rect 1344 927 1348 931
rect 1384 927 1388 931
rect 1424 927 1428 931
rect 1488 927 1492 931
rect 320 911 324 915
rect 328 911 332 915
rect 368 911 372 915
rect 376 911 380 915
rect 424 911 428 915
rect 432 911 436 915
rect 496 911 500 915
rect 576 911 580 915
rect 664 911 668 915
rect 752 911 756 915
rect 832 911 836 915
rect 840 911 844 915
rect 912 911 916 915
rect 920 911 924 915
rect 984 911 988 915
rect 992 911 996 915
rect 1048 911 1052 915
rect 1112 911 1116 915
rect 1120 911 1124 915
rect 1176 911 1180 915
rect 1216 911 1220 915
rect 1568 927 1572 931
rect 1576 927 1580 931
rect 1664 927 1668 931
rect 1672 927 1676 931
rect 1760 927 1764 931
rect 1768 927 1772 931
rect 1864 927 1868 931
rect 1960 927 1964 931
rect 2048 927 2052 931
rect 2056 927 2060 931
rect 2128 927 2132 931
rect 2200 927 2204 931
rect 2264 927 2268 931
rect 2336 927 2340 931
rect 2384 927 2388 931
rect 1344 895 1348 899
rect 1384 895 1388 899
rect 1424 895 1428 899
rect 1488 895 1492 899
rect 1496 895 1500 899
rect 1568 895 1572 899
rect 1576 895 1580 899
rect 1664 895 1668 899
rect 1672 895 1676 899
rect 1760 895 1764 899
rect 1768 895 1772 899
rect 1864 895 1868 899
rect 1960 895 1964 899
rect 2048 895 2052 899
rect 2056 895 2060 899
rect 2128 895 2132 899
rect 2200 895 2204 899
rect 2264 895 2268 899
rect 2336 895 2340 899
rect 2384 895 2388 899
rect 280 883 284 887
rect 296 883 300 887
rect 336 883 340 887
rect 400 883 404 887
rect 480 883 484 887
rect 560 883 564 887
rect 648 883 652 887
rect 736 883 740 887
rect 816 883 820 887
rect 888 883 892 887
rect 960 883 964 887
rect 1024 883 1028 887
rect 1080 883 1084 887
rect 1144 883 1148 887
rect 1208 883 1212 887
rect 280 851 284 855
rect 1360 867 1364 871
rect 1400 867 1404 871
rect 1440 867 1444 871
rect 1496 867 1500 871
rect 1560 867 1564 871
rect 1632 867 1636 871
rect 1704 867 1708 871
rect 1776 867 1780 871
rect 1848 867 1852 871
rect 1920 867 1924 871
rect 1984 867 1988 871
rect 2048 867 2052 871
rect 2112 867 2116 871
rect 2168 867 2172 871
rect 2184 867 2188 871
rect 2224 867 2228 871
rect 2280 867 2284 871
rect 2344 867 2348 871
rect 2384 867 2388 871
rect 336 851 340 855
rect 400 851 404 855
rect 480 851 484 855
rect 560 851 564 855
rect 648 851 652 855
rect 736 851 740 855
rect 816 851 820 855
rect 888 851 892 855
rect 960 851 964 855
rect 1024 851 1028 855
rect 1080 851 1084 855
rect 1144 851 1148 855
rect 1208 851 1212 855
rect 296 847 300 851
rect 1360 835 1364 839
rect 1400 835 1404 839
rect 1440 835 1444 839
rect 1496 835 1500 839
rect 1560 835 1564 839
rect 1632 835 1636 839
rect 1704 835 1708 839
rect 1776 835 1780 839
rect 1848 835 1852 839
rect 1920 837 1924 841
rect 1984 835 1988 839
rect 2048 835 2052 839
rect 2112 835 2116 839
rect 2168 835 2172 839
rect 216 799 220 803
rect 272 799 276 803
rect 336 799 340 803
rect 408 799 412 803
rect 488 799 492 803
rect 568 799 572 803
rect 576 799 580 803
rect 640 799 644 803
rect 712 799 716 803
rect 720 799 724 803
rect 776 799 780 803
rect 784 799 788 803
rect 840 799 844 803
rect 896 799 900 803
rect 952 799 956 803
rect 960 799 964 803
rect 1008 799 1012 803
rect 1016 799 1020 803
rect 1072 799 1076 803
rect 2224 835 2228 839
rect 2280 835 2284 839
rect 2344 835 2348 839
rect 2384 835 2388 839
rect 1328 779 1332 783
rect 1368 779 1372 783
rect 1432 779 1436 783
rect 1504 779 1508 783
rect 1512 779 1516 783
rect 1576 779 1580 783
rect 1648 779 1652 783
rect 1656 779 1660 783
rect 1720 779 1724 783
rect 1784 779 1788 783
rect 1808 779 1812 783
rect 1848 779 1852 783
rect 1856 779 1860 783
rect 1912 779 1916 783
rect 1920 779 1924 783
rect 1976 779 1980 783
rect 1984 779 1988 783
rect 2048 779 2052 783
rect 2128 779 2132 783
rect 2184 779 2188 783
rect 2216 779 2220 783
rect 2224 779 2228 783
rect 2304 779 2308 783
rect 2384 779 2388 783
rect 216 767 220 771
rect 272 767 276 771
rect 336 767 340 771
rect 408 767 412 771
rect 488 767 492 771
rect 568 767 572 771
rect 576 767 580 771
rect 640 767 644 771
rect 712 767 716 771
rect 720 767 724 771
rect 776 767 780 771
rect 784 767 788 771
rect 840 767 844 771
rect 896 767 900 771
rect 952 767 956 771
rect 960 767 964 771
rect 1008 767 1012 771
rect 1016 767 1020 771
rect 1072 767 1076 771
rect 160 747 164 751
rect 200 747 204 751
rect 240 747 244 751
rect 304 747 308 751
rect 376 747 380 751
rect 448 747 452 751
rect 520 747 524 751
rect 584 747 588 751
rect 648 747 652 751
rect 720 747 724 751
rect 808 747 812 751
rect 904 747 908 751
rect 1008 747 1012 751
rect 1120 747 1124 751
rect 1216 747 1220 751
rect 1328 747 1332 751
rect 1368 747 1372 751
rect 1432 747 1436 751
rect 1504 747 1508 751
rect 1512 747 1516 751
rect 1576 747 1580 751
rect 1648 747 1652 751
rect 1656 747 1660 751
rect 1720 747 1724 751
rect 1784 747 1788 751
rect 1808 747 1812 751
rect 1848 747 1852 751
rect 1856 747 1860 751
rect 1912 747 1916 751
rect 1920 747 1924 751
rect 1976 747 1980 751
rect 1984 747 1988 751
rect 2048 747 2052 751
rect 2128 747 2132 751
rect 2216 747 2220 751
rect 2224 747 2228 751
rect 2304 747 2308 751
rect 2384 747 2388 751
rect 168 735 172 739
rect 1328 727 1332 731
rect 1392 727 1396 731
rect 1480 727 1484 731
rect 1560 727 1564 731
rect 1640 727 1644 731
rect 1720 727 1724 731
rect 1800 727 1804 731
rect 1880 727 1884 731
rect 1968 727 1972 731
rect 2056 727 2060 731
rect 2144 727 2148 731
rect 2232 727 2236 731
rect 2320 727 2324 731
rect 2384 727 2388 731
rect 160 715 164 719
rect 168 715 172 719
rect 200 715 204 719
rect 240 715 244 719
rect 304 715 308 719
rect 376 715 380 719
rect 448 715 452 719
rect 520 715 524 719
rect 584 715 588 719
rect 648 715 652 719
rect 720 715 724 719
rect 808 715 812 719
rect 904 715 908 719
rect 1008 715 1012 719
rect 1120 715 1124 719
rect 1216 715 1220 719
rect 1328 695 1332 699
rect 1392 695 1396 699
rect 1480 695 1484 699
rect 1560 695 1564 699
rect 1640 695 1644 699
rect 1720 695 1724 699
rect 1800 695 1804 699
rect 1880 695 1884 699
rect 1968 695 1972 699
rect 2056 695 2060 699
rect 2144 695 2148 699
rect 2232 695 2236 699
rect 2320 695 2324 699
rect 2384 695 2388 699
rect 160 655 164 659
rect 200 655 204 659
rect 256 655 260 659
rect 264 655 268 659
rect 312 655 316 659
rect 368 655 372 659
rect 376 655 380 659
rect 424 655 428 659
rect 480 655 484 659
rect 528 655 532 659
rect 584 655 588 659
rect 648 655 652 659
rect 720 655 724 659
rect 792 655 796 659
rect 800 655 804 659
rect 864 655 868 659
rect 928 655 932 659
rect 936 655 940 659
rect 992 655 996 659
rect 1000 655 1004 659
rect 1048 655 1052 659
rect 1112 655 1116 659
rect 1120 655 1124 659
rect 1176 655 1180 659
rect 1216 655 1220 659
rect 1616 643 1620 647
rect 1664 643 1668 647
rect 1672 643 1676 647
rect 1712 643 1716 647
rect 1720 643 1724 647
rect 1768 643 1772 647
rect 1776 643 1780 647
rect 1824 643 1828 647
rect 1832 643 1836 647
rect 1896 643 1900 647
rect 1976 643 1980 647
rect 1984 643 1988 647
rect 2072 643 2076 647
rect 2176 643 2180 647
rect 2288 643 2292 647
rect 2384 643 2388 647
rect 2392 643 2396 647
rect 160 623 164 627
rect 200 623 204 627
rect 256 623 260 627
rect 264 623 268 627
rect 312 623 316 627
rect 368 623 372 627
rect 376 623 380 627
rect 424 623 428 627
rect 480 623 484 627
rect 528 623 532 627
rect 584 623 588 627
rect 648 623 652 627
rect 720 623 724 627
rect 792 623 796 627
rect 800 623 804 627
rect 864 623 868 627
rect 928 623 932 627
rect 936 623 940 627
rect 992 623 996 627
rect 1000 623 1004 627
rect 1048 623 1052 627
rect 1112 623 1116 627
rect 1120 623 1124 627
rect 1176 623 1180 627
rect 1216 623 1220 627
rect 1616 611 1620 615
rect 1664 611 1668 615
rect 1672 611 1676 615
rect 1712 611 1716 615
rect 1720 611 1724 615
rect 1768 611 1772 615
rect 1776 611 1780 615
rect 1824 611 1828 615
rect 1832 611 1836 615
rect 1896 611 1900 615
rect 1976 611 1980 615
rect 1984 611 1988 615
rect 2072 611 2076 615
rect 2176 611 2180 615
rect 2216 611 2220 615
rect 2288 611 2292 615
rect 2384 611 2388 615
rect 160 603 164 607
rect 208 603 212 607
rect 280 603 284 607
rect 352 603 356 607
rect 424 603 428 607
rect 504 603 508 607
rect 584 603 588 607
rect 664 603 668 607
rect 744 603 748 607
rect 824 603 828 607
rect 904 603 908 607
rect 976 603 980 607
rect 1040 603 1044 607
rect 1104 603 1108 607
rect 1168 603 1172 607
rect 1216 603 1220 607
rect 1584 583 1588 587
rect 1624 583 1628 587
rect 1664 583 1668 587
rect 1704 583 1708 587
rect 1744 583 1748 587
rect 1784 583 1788 587
rect 1832 583 1836 587
rect 1880 583 1884 587
rect 1936 583 1940 587
rect 1992 583 1996 587
rect 2056 583 2060 587
rect 2120 583 2124 587
rect 2192 583 2196 587
rect 160 571 164 575
rect 208 571 212 575
rect 280 571 284 575
rect 352 571 356 575
rect 424 571 428 575
rect 504 571 508 575
rect 584 571 588 575
rect 664 571 668 575
rect 744 571 748 575
rect 824 571 828 575
rect 904 571 908 575
rect 976 571 980 575
rect 1040 571 1044 575
rect 1104 571 1108 575
rect 1168 571 1172 575
rect 1216 571 1220 575
rect 2264 583 2268 587
rect 2336 583 2340 587
rect 2384 583 2388 587
rect 2392 583 2396 587
rect 1584 551 1588 555
rect 1624 551 1628 555
rect 1664 551 1668 555
rect 1704 551 1708 555
rect 1744 551 1748 555
rect 1784 551 1788 555
rect 1832 551 1836 555
rect 1880 551 1884 555
rect 1936 551 1940 555
rect 1992 551 1996 555
rect 2056 551 2060 555
rect 2120 551 2124 555
rect 2192 551 2196 555
rect 2216 551 2220 555
rect 2264 551 2268 555
rect 2336 551 2340 555
rect 2384 551 2388 555
rect 176 515 180 519
rect 184 515 188 519
rect 248 515 252 519
rect 312 515 316 519
rect 376 515 380 519
rect 384 515 388 519
rect 440 515 444 519
rect 448 515 452 519
rect 504 515 508 519
rect 512 515 516 519
rect 576 515 580 519
rect 648 515 652 519
rect 720 515 724 519
rect 728 515 732 519
rect 792 515 796 519
rect 864 515 868 519
rect 944 515 948 519
rect 1024 515 1028 519
rect 1032 515 1036 519
rect 1104 515 1108 519
rect 1432 499 1436 503
rect 1472 499 1476 503
rect 1512 499 1516 503
rect 1520 499 1524 503
rect 1560 499 1564 503
rect 1568 499 1572 503
rect 1616 499 1620 503
rect 1624 499 1628 503
rect 1672 499 1676 503
rect 1680 499 1684 503
rect 1736 499 1740 503
rect 1808 499 1812 503
rect 1888 499 1892 503
rect 1968 499 1972 503
rect 2048 499 2052 503
rect 2056 499 2060 503
rect 2128 499 2132 503
rect 2216 499 2220 503
rect 2312 499 2316 503
rect 2384 499 2388 503
rect 176 483 180 487
rect 184 483 188 487
rect 248 483 252 487
rect 312 483 316 487
rect 376 483 380 487
rect 384 483 388 487
rect 440 483 444 487
rect 448 483 452 487
rect 504 483 508 487
rect 512 483 516 487
rect 576 483 580 487
rect 648 483 652 487
rect 720 483 724 487
rect 728 483 732 487
rect 792 483 796 487
rect 864 483 868 487
rect 944 483 948 487
rect 1024 483 1028 487
rect 1032 483 1036 487
rect 1104 483 1108 487
rect 264 465 268 469
rect 1432 467 1436 471
rect 1472 467 1476 471
rect 1512 467 1516 471
rect 1520 467 1524 471
rect 1560 467 1564 471
rect 1568 467 1572 471
rect 1616 467 1620 471
rect 1624 467 1628 471
rect 1672 467 1676 471
rect 1680 467 1684 471
rect 1736 467 1740 471
rect 1808 467 1812 471
rect 1888 467 1892 471
rect 1968 467 1972 471
rect 2048 467 2052 471
rect 2056 467 2060 471
rect 2128 467 2132 471
rect 2216 467 2220 471
rect 2312 467 2316 471
rect 2384 467 2388 471
rect 304 463 308 467
rect 352 463 356 467
rect 408 463 412 467
rect 464 463 468 467
rect 528 463 532 467
rect 592 463 596 467
rect 656 463 660 467
rect 720 463 724 467
rect 784 463 788 467
rect 848 463 852 467
rect 912 463 916 467
rect 976 463 980 467
rect 1040 463 1044 467
rect 1328 447 1332 451
rect 1368 447 1372 451
rect 1408 447 1412 451
rect 1472 447 1476 451
rect 1560 447 1564 451
rect 1656 447 1660 451
rect 1760 447 1764 451
rect 1856 447 1860 451
rect 1944 447 1948 451
rect 2024 449 2028 453
rect 2096 447 2100 451
rect 2160 447 2164 451
rect 2224 447 2228 451
rect 2280 447 2284 451
rect 2344 447 2348 451
rect 2384 447 2388 451
rect 264 431 268 435
rect 304 431 308 435
rect 352 431 356 435
rect 408 431 412 435
rect 464 431 468 435
rect 528 431 532 435
rect 592 431 596 435
rect 656 431 660 435
rect 720 431 724 435
rect 784 431 788 435
rect 848 431 852 435
rect 912 431 916 435
rect 976 431 980 435
rect 1040 431 1044 435
rect 1328 415 1332 419
rect 1368 415 1372 419
rect 1408 415 1412 419
rect 1472 415 1476 419
rect 1560 415 1564 419
rect 1656 415 1660 419
rect 1760 415 1764 419
rect 1856 415 1860 419
rect 1944 415 1948 419
rect 2024 415 2028 419
rect 2096 415 2100 419
rect 2160 415 2164 419
rect 2224 415 2228 419
rect 2280 415 2284 419
rect 2344 415 2348 419
rect 2384 415 2388 419
rect 168 375 172 379
rect 208 375 212 379
rect 248 375 252 379
rect 296 375 300 379
rect 360 375 364 379
rect 368 375 372 379
rect 424 375 428 379
rect 432 375 436 379
rect 496 375 500 379
rect 568 375 572 379
rect 640 375 644 379
rect 712 375 716 379
rect 776 375 780 379
rect 832 375 836 379
rect 888 375 892 379
rect 944 375 948 379
rect 952 375 956 379
rect 1000 375 1004 379
rect 1008 375 1012 379
rect 1056 375 1060 379
rect 168 343 172 347
rect 208 343 212 347
rect 248 343 252 347
rect 296 343 300 347
rect 360 343 364 347
rect 368 343 372 347
rect 424 343 428 347
rect 432 343 436 347
rect 496 343 500 347
rect 568 345 572 349
rect 1384 363 1388 367
rect 1424 363 1428 367
rect 1464 363 1468 367
rect 1512 363 1516 367
rect 1568 363 1572 367
rect 1632 363 1636 367
rect 1640 363 1644 367
rect 1704 363 1708 367
rect 1784 363 1788 367
rect 1864 363 1868 367
rect 1944 363 1948 367
rect 1952 363 1956 367
rect 2024 363 2028 367
rect 2104 363 2108 367
rect 2184 363 2188 367
rect 2272 363 2276 367
rect 2360 363 2364 367
rect 640 343 644 347
rect 712 343 716 347
rect 776 343 780 347
rect 832 343 836 347
rect 888 343 892 347
rect 944 343 948 347
rect 952 343 956 347
rect 1000 343 1004 347
rect 1008 343 1012 347
rect 1056 343 1060 347
rect 1384 331 1388 335
rect 1424 331 1428 335
rect 1464 331 1468 335
rect 1512 331 1516 335
rect 1568 331 1572 335
rect 1632 331 1636 335
rect 1640 331 1644 335
rect 1704 331 1708 335
rect 1784 331 1788 335
rect 1864 331 1868 335
rect 1944 331 1948 335
rect 1952 331 1956 335
rect 2024 331 2028 335
rect 2104 331 2108 335
rect 2184 331 2188 335
rect 2272 331 2276 335
rect 2360 331 2364 335
rect 160 315 164 319
rect 200 315 204 319
rect 240 315 244 319
rect 280 315 284 319
rect 320 315 324 319
rect 360 315 364 319
rect 416 315 420 319
rect 472 315 476 319
rect 520 315 524 319
rect 568 315 572 319
rect 616 315 620 319
rect 664 315 668 319
rect 712 315 716 319
rect 760 315 764 319
rect 808 315 812 319
rect 864 315 868 319
rect 1536 303 1540 307
rect 1576 303 1580 307
rect 1616 303 1620 307
rect 1656 303 1660 307
rect 1696 303 1700 307
rect 1736 303 1740 307
rect 1776 303 1780 307
rect 1816 303 1820 307
rect 1864 303 1868 307
rect 1928 303 1932 307
rect 1992 303 1996 307
rect 2064 303 2068 307
rect 2144 303 2148 307
rect 2224 303 2228 307
rect 2304 303 2308 307
rect 2384 303 2388 307
rect 1544 291 1548 295
rect 160 283 164 287
rect 200 283 204 287
rect 240 283 244 287
rect 280 283 284 287
rect 320 283 324 287
rect 360 283 364 287
rect 416 283 420 287
rect 472 283 476 287
rect 520 283 524 287
rect 568 283 572 287
rect 616 283 620 287
rect 664 283 668 287
rect 712 283 716 287
rect 760 283 764 287
rect 808 283 812 287
rect 864 283 868 287
rect 1536 271 1540 275
rect 1544 271 1548 275
rect 1576 271 1580 275
rect 1616 271 1620 275
rect 1656 271 1660 275
rect 1696 271 1700 275
rect 1736 271 1740 275
rect 1776 271 1780 275
rect 1816 271 1820 275
rect 1864 271 1868 275
rect 1928 271 1932 275
rect 1992 271 1996 275
rect 2064 271 2068 275
rect 2144 271 2148 275
rect 2224 271 2228 275
rect 2304 271 2308 275
rect 2384 271 2388 275
rect 160 223 164 227
rect 248 223 252 227
rect 336 223 340 227
rect 344 223 348 227
rect 416 223 420 227
rect 424 223 428 227
rect 488 223 492 227
rect 496 223 500 227
rect 552 223 556 227
rect 560 223 564 227
rect 616 223 620 227
rect 624 223 628 227
rect 672 223 676 227
rect 720 223 724 227
rect 760 223 764 227
rect 768 223 772 227
rect 808 223 812 227
rect 816 223 820 227
rect 856 223 860 227
rect 864 223 868 227
rect 904 223 908 227
rect 912 223 916 227
rect 952 223 956 227
rect 960 223 964 227
rect 1000 223 1004 227
rect 1008 223 1012 227
rect 1048 223 1052 227
rect 1392 215 1396 219
rect 1432 215 1436 219
rect 1440 215 1444 219
rect 1480 215 1484 219
rect 1488 215 1492 219
rect 1536 215 1540 219
rect 1544 215 1548 219
rect 1592 215 1596 219
rect 1600 215 1604 219
rect 1656 215 1660 219
rect 1664 215 1668 219
rect 1728 215 1732 219
rect 1800 215 1804 219
rect 1808 215 1812 219
rect 1880 215 1884 219
rect 1888 215 1892 219
rect 1968 215 1972 219
rect 1976 215 1980 219
rect 2056 215 2060 219
rect 2064 215 2068 219
rect 2144 215 2148 219
rect 2232 215 2236 219
rect 2320 215 2324 219
rect 2384 215 2388 219
rect 160 191 164 195
rect 248 191 252 195
rect 336 191 340 195
rect 344 191 348 195
rect 416 191 420 195
rect 424 191 428 195
rect 488 191 492 195
rect 496 191 500 195
rect 552 191 556 195
rect 560 191 564 195
rect 616 191 620 195
rect 624 191 628 195
rect 672 191 676 195
rect 720 191 724 195
rect 760 191 764 195
rect 768 191 772 195
rect 808 191 812 195
rect 816 191 820 195
rect 856 191 860 195
rect 864 191 868 195
rect 904 191 908 195
rect 912 191 916 195
rect 952 191 956 195
rect 960 191 964 195
rect 1000 191 1004 195
rect 1008 191 1012 195
rect 1048 191 1052 195
rect 1392 183 1396 187
rect 1432 183 1436 187
rect 1440 183 1444 187
rect 1480 183 1484 187
rect 1488 183 1492 187
rect 1536 183 1540 187
rect 1544 183 1548 187
rect 1592 183 1596 187
rect 1600 183 1604 187
rect 1656 183 1660 187
rect 1664 183 1668 187
rect 1728 183 1732 187
rect 1800 183 1804 187
rect 1808 183 1812 187
rect 1880 183 1884 187
rect 1888 183 1892 187
rect 1968 183 1972 187
rect 1976 183 1980 187
rect 2056 183 2060 187
rect 2064 183 2068 187
rect 2144 183 2148 187
rect 2232 183 2236 187
rect 2320 183 2324 187
rect 2384 183 2388 187
rect 1328 155 1332 159
rect 1368 155 1372 159
rect 1408 155 1412 159
rect 1448 155 1452 159
rect 1488 155 1492 159
rect 1544 155 1548 159
rect 1608 155 1612 159
rect 1672 155 1676 159
rect 1736 155 1740 159
rect 1800 155 1804 159
rect 1856 155 1860 159
rect 1912 155 1916 159
rect 1960 155 1964 159
rect 2000 155 2004 159
rect 2040 155 2044 159
rect 2080 155 2084 159
rect 2120 155 2124 159
rect 2168 155 2172 159
rect 2216 155 2220 159
rect 2264 155 2268 159
rect 2304 155 2308 159
rect 2344 155 2348 159
rect 2384 155 2388 159
rect 176 139 180 143
rect 216 139 220 143
rect 256 139 260 143
rect 296 139 300 143
rect 336 139 340 143
rect 376 139 380 143
rect 416 139 420 143
rect 456 139 460 143
rect 496 139 500 143
rect 536 139 540 143
rect 576 139 580 143
rect 616 139 620 143
rect 656 139 660 143
rect 696 139 700 143
rect 736 139 740 143
rect 776 139 780 143
rect 816 139 820 143
rect 856 139 860 143
rect 896 139 900 143
rect 936 139 940 143
rect 976 139 980 143
rect 1016 139 1020 143
rect 1056 139 1060 143
rect 1096 139 1100 143
rect 1136 139 1140 143
rect 1176 139 1180 143
rect 1216 139 1220 143
rect 1328 123 1332 127
rect 1368 123 1372 127
rect 1408 123 1412 127
rect 1448 123 1452 127
rect 1488 123 1492 127
rect 1544 123 1548 127
rect 1608 123 1612 127
rect 1672 123 1676 127
rect 1736 123 1740 127
rect 1800 123 1804 127
rect 1856 123 1860 127
rect 1912 123 1916 127
rect 1960 123 1964 127
rect 2000 123 2004 127
rect 2040 123 2044 127
rect 2080 123 2084 127
rect 2120 123 2124 127
rect 2168 123 2172 127
rect 2216 123 2220 127
rect 2264 123 2268 127
rect 2304 123 2308 127
rect 2344 123 2348 127
rect 2384 123 2388 127
rect 216 107 220 111
rect 256 107 260 111
rect 296 107 300 111
rect 336 107 340 111
rect 376 107 380 111
rect 416 107 420 111
rect 456 107 460 111
rect 496 107 500 111
rect 536 107 540 111
rect 576 107 580 111
rect 616 107 620 111
rect 656 107 660 111
rect 696 107 700 111
rect 736 107 740 111
rect 776 107 780 111
rect 816 107 820 111
rect 856 107 860 111
rect 896 107 900 111
rect 936 107 940 111
rect 976 107 980 111
rect 1016 107 1020 111
rect 1056 107 1060 111
rect 1096 107 1100 111
rect 1136 107 1140 111
rect 1176 107 1180 111
rect 1216 107 1220 111
<< m2 >>
rect 326 2487 332 2488
rect 326 2486 327 2487
rect 304 2484 327 2486
rect 255 2483 264 2484
rect 230 2479 236 2480
rect 230 2475 231 2479
rect 235 2475 236 2479
rect 255 2479 256 2483
rect 263 2479 264 2483
rect 295 2483 301 2484
rect 255 2478 264 2479
rect 270 2479 276 2480
rect 230 2474 236 2475
rect 270 2475 271 2479
rect 275 2475 276 2479
rect 295 2479 296 2483
rect 300 2482 301 2483
rect 304 2482 306 2484
rect 326 2483 327 2484
rect 331 2483 332 2487
rect 358 2487 364 2488
rect 358 2486 359 2487
rect 344 2484 359 2486
rect 326 2482 332 2483
rect 335 2483 341 2484
rect 300 2480 306 2482
rect 300 2479 301 2480
rect 295 2478 301 2479
rect 310 2479 316 2480
rect 270 2474 276 2475
rect 310 2475 311 2479
rect 315 2475 316 2479
rect 335 2479 336 2483
rect 340 2482 341 2483
rect 344 2482 346 2484
rect 358 2483 359 2484
rect 363 2483 364 2487
rect 782 2487 788 2488
rect 782 2486 783 2487
rect 760 2484 783 2486
rect 358 2482 364 2483
rect 375 2483 381 2484
rect 340 2480 346 2482
rect 340 2479 341 2480
rect 335 2478 341 2479
rect 350 2479 356 2480
rect 310 2474 316 2475
rect 350 2475 351 2479
rect 355 2475 356 2479
rect 375 2479 376 2483
rect 380 2482 381 2483
rect 390 2483 396 2484
rect 390 2482 391 2483
rect 380 2480 391 2482
rect 380 2479 381 2480
rect 375 2478 381 2479
rect 390 2479 391 2480
rect 395 2479 396 2483
rect 423 2483 429 2484
rect 390 2478 396 2479
rect 398 2479 404 2480
rect 350 2474 356 2475
rect 398 2475 399 2479
rect 403 2475 404 2479
rect 423 2479 424 2483
rect 428 2482 429 2483
rect 446 2483 452 2484
rect 446 2482 447 2483
rect 428 2480 447 2482
rect 428 2479 429 2480
rect 423 2478 429 2479
rect 446 2479 447 2480
rect 451 2479 452 2483
rect 479 2483 485 2484
rect 446 2478 452 2479
rect 454 2479 460 2480
rect 398 2474 404 2475
rect 454 2475 455 2479
rect 459 2475 460 2479
rect 479 2479 480 2483
rect 484 2482 485 2483
rect 502 2483 508 2484
rect 502 2482 503 2483
rect 484 2480 503 2482
rect 484 2479 485 2480
rect 479 2478 485 2479
rect 502 2479 503 2480
rect 507 2479 508 2483
rect 535 2483 541 2484
rect 502 2478 508 2479
rect 510 2479 516 2480
rect 454 2474 460 2475
rect 510 2475 511 2479
rect 515 2475 516 2479
rect 535 2479 536 2483
rect 540 2482 541 2483
rect 566 2483 572 2484
rect 566 2482 567 2483
rect 540 2480 567 2482
rect 540 2479 541 2480
rect 535 2478 541 2479
rect 566 2479 567 2480
rect 571 2479 572 2483
rect 599 2483 605 2484
rect 566 2478 572 2479
rect 574 2479 580 2480
rect 510 2474 516 2475
rect 574 2475 575 2479
rect 579 2475 580 2479
rect 599 2479 600 2483
rect 604 2482 605 2483
rect 630 2483 636 2484
rect 630 2482 631 2483
rect 604 2480 631 2482
rect 604 2479 605 2480
rect 599 2478 605 2479
rect 630 2479 631 2480
rect 635 2479 636 2483
rect 650 2483 656 2484
rect 630 2478 636 2479
rect 638 2479 644 2480
rect 574 2474 580 2475
rect 638 2475 639 2479
rect 643 2475 644 2479
rect 650 2479 651 2483
rect 655 2482 656 2483
rect 663 2483 669 2484
rect 663 2482 664 2483
rect 655 2480 664 2482
rect 655 2479 656 2480
rect 650 2478 656 2479
rect 663 2479 664 2480
rect 668 2479 669 2483
rect 727 2483 733 2484
rect 663 2478 669 2479
rect 702 2479 708 2480
rect 638 2474 644 2475
rect 702 2475 703 2479
rect 707 2475 708 2479
rect 727 2479 728 2483
rect 732 2482 733 2483
rect 760 2482 762 2484
rect 782 2483 783 2484
rect 787 2483 788 2487
rect 1126 2487 1132 2488
rect 1126 2486 1127 2487
rect 1104 2484 1127 2486
rect 782 2482 788 2483
rect 791 2483 797 2484
rect 732 2480 762 2482
rect 732 2479 733 2480
rect 727 2478 733 2479
rect 766 2479 772 2480
rect 702 2474 708 2475
rect 766 2475 767 2479
rect 771 2475 772 2479
rect 791 2479 792 2483
rect 796 2482 797 2483
rect 814 2483 820 2484
rect 814 2482 815 2483
rect 796 2480 815 2482
rect 796 2479 797 2480
rect 791 2478 797 2479
rect 814 2479 815 2480
rect 819 2479 820 2483
rect 847 2483 853 2484
rect 814 2478 820 2479
rect 822 2479 828 2480
rect 766 2474 772 2475
rect 822 2475 823 2479
rect 827 2475 828 2479
rect 847 2479 848 2483
rect 852 2482 853 2483
rect 870 2483 876 2484
rect 870 2482 871 2483
rect 852 2480 871 2482
rect 852 2479 853 2480
rect 847 2478 853 2479
rect 870 2479 871 2480
rect 875 2479 876 2483
rect 903 2483 909 2484
rect 870 2478 876 2479
rect 878 2479 884 2480
rect 822 2474 828 2475
rect 878 2475 879 2479
rect 883 2475 884 2479
rect 903 2479 904 2483
rect 908 2482 909 2483
rect 918 2483 924 2484
rect 918 2482 919 2483
rect 908 2480 919 2482
rect 908 2479 909 2480
rect 903 2478 909 2479
rect 918 2479 919 2480
rect 923 2479 924 2483
rect 951 2483 957 2484
rect 918 2478 924 2479
rect 926 2479 932 2480
rect 878 2474 884 2475
rect 926 2475 927 2479
rect 931 2475 932 2479
rect 951 2479 952 2483
rect 956 2482 957 2483
rect 966 2483 972 2484
rect 966 2482 967 2483
rect 956 2480 967 2482
rect 956 2479 957 2480
rect 951 2478 957 2479
rect 966 2479 967 2480
rect 971 2479 972 2483
rect 999 2483 1005 2484
rect 966 2478 972 2479
rect 974 2479 980 2480
rect 926 2474 932 2475
rect 974 2475 975 2479
rect 979 2475 980 2479
rect 999 2479 1000 2483
rect 1004 2482 1005 2483
rect 1014 2483 1020 2484
rect 1014 2482 1015 2483
rect 1004 2480 1015 2482
rect 1004 2479 1005 2480
rect 999 2478 1005 2479
rect 1014 2479 1015 2480
rect 1019 2479 1020 2483
rect 1047 2483 1053 2484
rect 1014 2478 1020 2479
rect 1022 2479 1028 2480
rect 974 2474 980 2475
rect 1022 2475 1023 2479
rect 1027 2475 1028 2479
rect 1047 2479 1048 2483
rect 1052 2482 1053 2483
rect 1062 2483 1068 2484
rect 1062 2482 1063 2483
rect 1052 2480 1063 2482
rect 1052 2479 1053 2480
rect 1047 2478 1053 2479
rect 1062 2479 1063 2480
rect 1067 2479 1068 2483
rect 1095 2483 1101 2484
rect 1062 2478 1068 2479
rect 1070 2479 1076 2480
rect 1022 2474 1028 2475
rect 1070 2475 1071 2479
rect 1075 2475 1076 2479
rect 1095 2479 1096 2483
rect 1100 2482 1101 2483
rect 1104 2482 1106 2484
rect 1126 2483 1127 2484
rect 1131 2483 1132 2487
rect 1166 2487 1172 2488
rect 1166 2486 1167 2487
rect 1144 2484 1167 2486
rect 1126 2482 1132 2483
rect 1135 2483 1141 2484
rect 1100 2480 1106 2482
rect 1100 2479 1101 2480
rect 1095 2478 1101 2479
rect 1110 2479 1116 2480
rect 1070 2474 1076 2475
rect 1110 2475 1111 2479
rect 1115 2475 1116 2479
rect 1135 2479 1136 2483
rect 1140 2482 1141 2483
rect 1144 2482 1146 2484
rect 1166 2483 1167 2484
rect 1171 2483 1172 2487
rect 1202 2487 1208 2488
rect 1202 2486 1203 2487
rect 1184 2484 1203 2486
rect 1166 2482 1172 2483
rect 1175 2483 1181 2484
rect 1140 2480 1146 2482
rect 1140 2479 1141 2480
rect 1135 2478 1141 2479
rect 1150 2479 1156 2480
rect 1110 2474 1116 2475
rect 1150 2475 1151 2479
rect 1155 2475 1156 2479
rect 1175 2479 1176 2483
rect 1180 2482 1181 2483
rect 1184 2482 1186 2484
rect 1202 2483 1203 2484
rect 1207 2483 1208 2487
rect 1202 2482 1208 2483
rect 1215 2483 1221 2484
rect 1180 2480 1186 2482
rect 1180 2479 1181 2480
rect 1175 2478 1181 2479
rect 1190 2479 1196 2480
rect 1150 2474 1156 2475
rect 1190 2475 1191 2479
rect 1195 2475 1196 2479
rect 1215 2479 1216 2483
rect 1220 2482 1221 2483
rect 1318 2483 1324 2484
rect 1318 2482 1319 2483
rect 1220 2480 1319 2482
rect 1220 2479 1221 2480
rect 1215 2478 1221 2479
rect 1318 2479 1319 2480
rect 1323 2479 1324 2483
rect 1358 2483 1364 2484
rect 1358 2482 1359 2483
rect 1336 2480 1359 2482
rect 1318 2478 1324 2479
rect 1327 2479 1333 2480
rect 1190 2474 1196 2475
rect 1302 2475 1308 2476
rect 1302 2471 1303 2475
rect 1307 2471 1308 2475
rect 1327 2475 1328 2479
rect 1332 2478 1333 2479
rect 1336 2478 1338 2480
rect 1358 2479 1359 2480
rect 1363 2479 1364 2483
rect 1398 2483 1404 2484
rect 1398 2482 1399 2483
rect 1376 2480 1399 2482
rect 1358 2478 1364 2479
rect 1367 2479 1373 2480
rect 1332 2476 1338 2478
rect 1332 2475 1333 2476
rect 1327 2474 1333 2475
rect 1342 2475 1348 2476
rect 1302 2470 1308 2471
rect 1342 2471 1343 2475
rect 1347 2471 1348 2475
rect 1367 2475 1368 2479
rect 1372 2478 1373 2479
rect 1376 2478 1378 2480
rect 1398 2479 1399 2480
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1407 2479 1413 2480
rect 1372 2476 1378 2478
rect 1372 2475 1373 2476
rect 1367 2474 1373 2475
rect 1382 2475 1388 2476
rect 1342 2470 1348 2471
rect 1382 2471 1383 2475
rect 1387 2471 1388 2475
rect 1407 2475 1408 2479
rect 1412 2478 1413 2479
rect 1430 2479 1436 2480
rect 1430 2478 1431 2479
rect 1412 2476 1431 2478
rect 1412 2475 1413 2476
rect 1407 2474 1413 2475
rect 1430 2475 1431 2476
rect 1435 2475 1436 2479
rect 1463 2479 1469 2480
rect 1430 2474 1436 2475
rect 1438 2475 1444 2476
rect 1382 2470 1388 2471
rect 1438 2471 1439 2475
rect 1443 2471 1444 2475
rect 1463 2475 1464 2479
rect 1468 2478 1469 2479
rect 1502 2479 1508 2480
rect 1502 2478 1503 2479
rect 1468 2476 1503 2478
rect 1468 2475 1469 2476
rect 1463 2474 1469 2475
rect 1502 2475 1503 2476
rect 1507 2475 1508 2479
rect 1535 2479 1541 2480
rect 1502 2474 1508 2475
rect 1510 2475 1516 2476
rect 1438 2470 1444 2471
rect 1510 2471 1511 2475
rect 1515 2471 1516 2475
rect 1535 2475 1536 2479
rect 1540 2478 1541 2479
rect 1574 2479 1580 2480
rect 1574 2478 1575 2479
rect 1540 2476 1575 2478
rect 1540 2475 1541 2476
rect 1535 2474 1541 2475
rect 1574 2475 1575 2476
rect 1579 2475 1580 2479
rect 1607 2479 1613 2480
rect 1574 2474 1580 2475
rect 1582 2475 1588 2476
rect 1510 2470 1516 2471
rect 1582 2471 1583 2475
rect 1587 2471 1588 2475
rect 1607 2475 1608 2479
rect 1612 2478 1613 2479
rect 1654 2479 1660 2480
rect 1654 2478 1655 2479
rect 1612 2476 1655 2478
rect 1612 2475 1613 2476
rect 1607 2474 1613 2475
rect 1654 2475 1655 2476
rect 1659 2475 1660 2479
rect 1686 2479 1693 2480
rect 1654 2474 1660 2475
rect 1662 2475 1668 2476
rect 1582 2470 1588 2471
rect 1662 2471 1663 2475
rect 1667 2471 1668 2475
rect 1686 2475 1687 2479
rect 1692 2475 1693 2479
rect 1759 2479 1765 2480
rect 1686 2474 1693 2475
rect 1734 2475 1740 2476
rect 1662 2470 1668 2471
rect 1734 2471 1735 2475
rect 1739 2471 1740 2475
rect 1759 2475 1760 2479
rect 1764 2478 1765 2479
rect 1798 2479 1804 2480
rect 1798 2478 1799 2479
rect 1764 2476 1799 2478
rect 1764 2475 1765 2476
rect 1759 2474 1765 2475
rect 1798 2475 1799 2476
rect 1803 2475 1804 2479
rect 1831 2479 1837 2480
rect 1798 2474 1804 2475
rect 1806 2475 1812 2476
rect 1734 2470 1740 2471
rect 1806 2471 1807 2475
rect 1811 2471 1812 2475
rect 1831 2475 1832 2479
rect 1836 2478 1837 2479
rect 1878 2479 1884 2480
rect 1878 2478 1879 2479
rect 1836 2476 1879 2478
rect 1836 2475 1837 2476
rect 1831 2474 1837 2475
rect 1878 2475 1879 2476
rect 1883 2475 1884 2479
rect 1911 2479 1917 2480
rect 1878 2474 1884 2475
rect 1886 2475 1892 2476
rect 1806 2470 1812 2471
rect 1886 2471 1887 2475
rect 1891 2471 1892 2475
rect 1911 2475 1912 2479
rect 1916 2478 1917 2479
rect 1958 2479 1964 2480
rect 1958 2478 1959 2479
rect 1916 2476 1959 2478
rect 1916 2475 1917 2476
rect 1911 2474 1917 2475
rect 1958 2475 1959 2476
rect 1963 2475 1964 2479
rect 1991 2479 1997 2480
rect 1958 2474 1964 2475
rect 1966 2475 1972 2476
rect 1886 2470 1892 2471
rect 1966 2471 1967 2475
rect 1971 2471 1972 2475
rect 1991 2475 1992 2479
rect 1996 2478 1997 2479
rect 2047 2479 2053 2480
rect 2047 2478 2048 2479
rect 1996 2476 2048 2478
rect 1996 2475 1997 2476
rect 1991 2474 1997 2475
rect 2047 2475 2048 2476
rect 2052 2475 2053 2479
rect 2087 2479 2093 2480
rect 2047 2474 2053 2475
rect 2062 2475 2068 2476
rect 1966 2470 1972 2471
rect 2062 2471 2063 2475
rect 2067 2471 2068 2475
rect 2087 2475 2088 2479
rect 2092 2478 2093 2479
rect 2158 2479 2164 2480
rect 2158 2478 2159 2479
rect 2092 2476 2159 2478
rect 2092 2475 2093 2476
rect 2087 2474 2093 2475
rect 2158 2475 2159 2476
rect 2163 2475 2164 2479
rect 2191 2479 2197 2480
rect 2158 2474 2164 2475
rect 2166 2475 2172 2476
rect 2062 2470 2068 2471
rect 2166 2471 2167 2475
rect 2171 2471 2172 2475
rect 2191 2475 2192 2479
rect 2196 2478 2197 2479
rect 2262 2479 2268 2480
rect 2262 2478 2263 2479
rect 2196 2476 2263 2478
rect 2196 2475 2197 2476
rect 2191 2474 2197 2475
rect 2262 2475 2263 2476
rect 2267 2475 2268 2479
rect 2286 2479 2292 2480
rect 2262 2474 2268 2475
rect 2270 2475 2276 2476
rect 2166 2470 2172 2471
rect 2270 2471 2271 2475
rect 2275 2471 2276 2475
rect 2286 2475 2287 2479
rect 2291 2478 2292 2479
rect 2295 2479 2301 2480
rect 2295 2478 2296 2479
rect 2291 2476 2296 2478
rect 2291 2475 2292 2476
rect 2286 2474 2292 2475
rect 2295 2475 2296 2476
rect 2300 2475 2301 2479
rect 2295 2474 2301 2475
rect 2358 2475 2364 2476
rect 2270 2470 2276 2471
rect 2358 2471 2359 2475
rect 2363 2471 2364 2475
rect 2358 2470 2364 2471
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 1238 2456 1244 2457
rect 1238 2452 1239 2456
rect 1243 2452 1244 2456
rect 110 2451 116 2452
rect 242 2451 248 2452
rect 242 2447 243 2451
rect 247 2450 248 2451
rect 255 2451 261 2452
rect 255 2450 256 2451
rect 247 2448 256 2450
rect 247 2447 248 2448
rect 242 2446 248 2447
rect 255 2447 256 2448
rect 260 2447 261 2451
rect 255 2446 261 2447
rect 266 2451 272 2452
rect 266 2447 267 2451
rect 271 2450 272 2451
rect 295 2451 301 2452
rect 295 2450 296 2451
rect 271 2448 296 2450
rect 271 2447 272 2448
rect 266 2446 272 2447
rect 295 2447 296 2448
rect 300 2447 301 2451
rect 295 2446 301 2447
rect 326 2451 332 2452
rect 326 2447 327 2451
rect 331 2450 332 2451
rect 335 2451 341 2452
rect 335 2450 336 2451
rect 331 2448 336 2450
rect 331 2447 332 2448
rect 326 2446 332 2447
rect 335 2447 336 2448
rect 340 2447 341 2451
rect 335 2446 341 2447
rect 358 2451 364 2452
rect 358 2447 359 2451
rect 363 2450 364 2451
rect 375 2451 381 2452
rect 375 2450 376 2451
rect 363 2448 376 2450
rect 363 2447 364 2448
rect 358 2446 364 2447
rect 375 2447 376 2448
rect 380 2447 381 2451
rect 375 2446 381 2447
rect 390 2451 396 2452
rect 390 2447 391 2451
rect 395 2450 396 2451
rect 423 2451 429 2452
rect 423 2450 424 2451
rect 395 2448 424 2450
rect 395 2447 396 2448
rect 390 2446 396 2447
rect 423 2447 424 2448
rect 428 2447 429 2451
rect 423 2446 429 2447
rect 446 2451 452 2452
rect 446 2447 447 2451
rect 451 2450 452 2451
rect 479 2451 485 2452
rect 479 2450 480 2451
rect 451 2448 480 2450
rect 451 2447 452 2448
rect 446 2446 452 2447
rect 479 2447 480 2448
rect 484 2447 485 2451
rect 479 2446 485 2447
rect 502 2451 508 2452
rect 502 2447 503 2451
rect 507 2450 508 2451
rect 535 2451 541 2452
rect 535 2450 536 2451
rect 507 2448 536 2450
rect 507 2447 508 2448
rect 502 2446 508 2447
rect 535 2447 536 2448
rect 540 2447 541 2451
rect 535 2446 541 2447
rect 566 2451 572 2452
rect 566 2447 567 2451
rect 571 2450 572 2451
rect 599 2451 605 2452
rect 599 2450 600 2451
rect 571 2448 600 2450
rect 571 2447 572 2448
rect 566 2446 572 2447
rect 599 2447 600 2448
rect 604 2447 605 2451
rect 599 2446 605 2447
rect 630 2451 636 2452
rect 630 2447 631 2451
rect 635 2450 636 2451
rect 663 2451 669 2452
rect 663 2450 664 2451
rect 635 2448 664 2450
rect 635 2447 636 2448
rect 630 2446 636 2447
rect 663 2447 664 2448
rect 668 2447 669 2451
rect 663 2446 669 2447
rect 727 2451 733 2452
rect 727 2447 728 2451
rect 732 2450 733 2451
rect 774 2451 780 2452
rect 774 2450 775 2451
rect 732 2448 775 2450
rect 732 2447 733 2448
rect 727 2446 733 2447
rect 774 2447 775 2448
rect 779 2447 780 2451
rect 774 2446 780 2447
rect 782 2451 788 2452
rect 782 2447 783 2451
rect 787 2450 788 2451
rect 791 2451 797 2452
rect 791 2450 792 2451
rect 787 2448 792 2450
rect 787 2447 788 2448
rect 782 2446 788 2447
rect 791 2447 792 2448
rect 796 2447 797 2451
rect 791 2446 797 2447
rect 814 2451 820 2452
rect 814 2447 815 2451
rect 819 2450 820 2451
rect 847 2451 853 2452
rect 847 2450 848 2451
rect 819 2448 848 2450
rect 819 2447 820 2448
rect 814 2446 820 2447
rect 847 2447 848 2448
rect 852 2447 853 2451
rect 847 2446 853 2447
rect 870 2451 876 2452
rect 870 2447 871 2451
rect 875 2450 876 2451
rect 903 2451 909 2452
rect 903 2450 904 2451
rect 875 2448 904 2450
rect 875 2447 876 2448
rect 870 2446 876 2447
rect 903 2447 904 2448
rect 908 2447 909 2451
rect 903 2446 909 2447
rect 918 2451 924 2452
rect 918 2447 919 2451
rect 923 2450 924 2451
rect 951 2451 957 2452
rect 951 2450 952 2451
rect 923 2448 952 2450
rect 923 2447 924 2448
rect 918 2446 924 2447
rect 951 2447 952 2448
rect 956 2447 957 2451
rect 951 2446 957 2447
rect 966 2451 972 2452
rect 966 2447 967 2451
rect 971 2450 972 2451
rect 999 2451 1005 2452
rect 999 2450 1000 2451
rect 971 2448 1000 2450
rect 971 2447 972 2448
rect 966 2446 972 2447
rect 999 2447 1000 2448
rect 1004 2447 1005 2451
rect 999 2446 1005 2447
rect 1014 2451 1020 2452
rect 1014 2447 1015 2451
rect 1019 2450 1020 2451
rect 1047 2451 1053 2452
rect 1047 2450 1048 2451
rect 1019 2448 1048 2450
rect 1019 2447 1020 2448
rect 1014 2446 1020 2447
rect 1047 2447 1048 2448
rect 1052 2447 1053 2451
rect 1047 2446 1053 2447
rect 1062 2451 1068 2452
rect 1062 2447 1063 2451
rect 1067 2450 1068 2451
rect 1095 2451 1101 2452
rect 1095 2450 1096 2451
rect 1067 2448 1096 2450
rect 1067 2447 1068 2448
rect 1062 2446 1068 2447
rect 1095 2447 1096 2448
rect 1100 2447 1101 2451
rect 1095 2446 1101 2447
rect 1126 2451 1132 2452
rect 1126 2447 1127 2451
rect 1131 2450 1132 2451
rect 1135 2451 1141 2452
rect 1135 2450 1136 2451
rect 1131 2448 1136 2450
rect 1131 2447 1132 2448
rect 1126 2446 1132 2447
rect 1135 2447 1136 2448
rect 1140 2447 1141 2451
rect 1135 2446 1141 2447
rect 1166 2451 1172 2452
rect 1166 2447 1167 2451
rect 1171 2450 1172 2451
rect 1175 2451 1181 2452
rect 1175 2450 1176 2451
rect 1171 2448 1176 2450
rect 1171 2447 1172 2448
rect 1166 2446 1172 2447
rect 1175 2447 1176 2448
rect 1180 2447 1181 2451
rect 1175 2446 1181 2447
rect 1202 2451 1208 2452
rect 1202 2447 1203 2451
rect 1207 2450 1208 2451
rect 1215 2451 1221 2452
rect 1238 2451 1244 2452
rect 1278 2452 1284 2453
rect 1215 2450 1216 2451
rect 1207 2448 1216 2450
rect 1207 2447 1208 2448
rect 1202 2446 1208 2447
rect 1215 2447 1216 2448
rect 1220 2447 1221 2451
rect 1278 2448 1279 2452
rect 1283 2448 1284 2452
rect 2406 2452 2412 2453
rect 2406 2448 2407 2452
rect 2411 2448 2412 2452
rect 1278 2447 1284 2448
rect 1318 2447 1324 2448
rect 1215 2446 1221 2447
rect 1318 2443 1319 2447
rect 1323 2446 1324 2447
rect 1327 2447 1333 2448
rect 1327 2446 1328 2447
rect 1323 2444 1328 2446
rect 1323 2443 1324 2444
rect 1318 2442 1324 2443
rect 1327 2443 1328 2444
rect 1332 2443 1333 2447
rect 1327 2442 1333 2443
rect 1358 2447 1364 2448
rect 1358 2443 1359 2447
rect 1363 2446 1364 2447
rect 1367 2447 1373 2448
rect 1367 2446 1368 2447
rect 1363 2444 1368 2446
rect 1363 2443 1364 2444
rect 1358 2442 1364 2443
rect 1367 2443 1368 2444
rect 1372 2443 1373 2447
rect 1367 2442 1373 2443
rect 1398 2447 1404 2448
rect 1398 2443 1399 2447
rect 1403 2446 1404 2447
rect 1407 2447 1413 2448
rect 1407 2446 1408 2447
rect 1403 2444 1408 2446
rect 1403 2443 1404 2444
rect 1398 2442 1404 2443
rect 1407 2443 1408 2444
rect 1412 2443 1413 2447
rect 1407 2442 1413 2443
rect 1430 2447 1436 2448
rect 1430 2443 1431 2447
rect 1435 2446 1436 2447
rect 1463 2447 1469 2448
rect 1463 2446 1464 2447
rect 1435 2444 1464 2446
rect 1435 2443 1436 2444
rect 1430 2442 1436 2443
rect 1463 2443 1464 2444
rect 1468 2443 1469 2447
rect 1463 2442 1469 2443
rect 1502 2447 1508 2448
rect 1502 2443 1503 2447
rect 1507 2446 1508 2447
rect 1535 2447 1541 2448
rect 1535 2446 1536 2447
rect 1507 2444 1536 2446
rect 1507 2443 1508 2444
rect 1502 2442 1508 2443
rect 1535 2443 1536 2444
rect 1540 2443 1541 2447
rect 1535 2442 1541 2443
rect 1574 2447 1580 2448
rect 1574 2443 1575 2447
rect 1579 2446 1580 2447
rect 1607 2447 1613 2448
rect 1607 2446 1608 2447
rect 1579 2444 1608 2446
rect 1579 2443 1580 2444
rect 1574 2442 1580 2443
rect 1607 2443 1608 2444
rect 1612 2443 1613 2447
rect 1607 2442 1613 2443
rect 1654 2447 1660 2448
rect 1654 2443 1655 2447
rect 1659 2446 1660 2447
rect 1687 2447 1693 2448
rect 1687 2446 1688 2447
rect 1659 2444 1688 2446
rect 1659 2443 1660 2444
rect 1654 2442 1660 2443
rect 1687 2443 1688 2444
rect 1692 2443 1693 2447
rect 1687 2442 1693 2443
rect 1759 2447 1765 2448
rect 1759 2443 1760 2447
rect 1764 2446 1765 2447
rect 1798 2447 1804 2448
rect 1764 2444 1795 2446
rect 1764 2443 1765 2444
rect 1759 2442 1765 2443
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 1238 2439 1244 2440
rect 1238 2435 1239 2439
rect 1243 2435 1244 2439
rect 1793 2438 1795 2444
rect 1798 2443 1799 2447
rect 1803 2446 1804 2447
rect 1831 2447 1837 2448
rect 1831 2446 1832 2447
rect 1803 2444 1832 2446
rect 1803 2443 1804 2444
rect 1798 2442 1804 2443
rect 1831 2443 1832 2444
rect 1836 2443 1837 2447
rect 1831 2442 1837 2443
rect 1878 2447 1884 2448
rect 1878 2443 1879 2447
rect 1883 2446 1884 2447
rect 1911 2447 1917 2448
rect 1911 2446 1912 2447
rect 1883 2444 1912 2446
rect 1883 2443 1884 2444
rect 1878 2442 1884 2443
rect 1911 2443 1912 2444
rect 1916 2443 1917 2447
rect 1911 2442 1917 2443
rect 1958 2447 1964 2448
rect 1958 2443 1959 2447
rect 1963 2446 1964 2447
rect 1991 2447 1997 2448
rect 1991 2446 1992 2447
rect 1963 2444 1992 2446
rect 1963 2443 1964 2444
rect 1958 2442 1964 2443
rect 1991 2443 1992 2444
rect 1996 2443 1997 2447
rect 1991 2442 1997 2443
rect 2047 2447 2053 2448
rect 2047 2443 2048 2447
rect 2052 2446 2053 2447
rect 2087 2447 2093 2448
rect 2087 2446 2088 2447
rect 2052 2444 2088 2446
rect 2052 2443 2053 2444
rect 2047 2442 2053 2443
rect 2087 2443 2088 2444
rect 2092 2443 2093 2447
rect 2087 2442 2093 2443
rect 2158 2447 2164 2448
rect 2158 2443 2159 2447
rect 2163 2446 2164 2447
rect 2191 2447 2197 2448
rect 2191 2446 2192 2447
rect 2163 2444 2192 2446
rect 2163 2443 2164 2444
rect 2158 2442 2164 2443
rect 2191 2443 2192 2444
rect 2196 2443 2197 2447
rect 2191 2442 2197 2443
rect 2262 2447 2268 2448
rect 2262 2443 2263 2447
rect 2267 2446 2268 2447
rect 2295 2447 2301 2448
rect 2295 2446 2296 2447
rect 2267 2444 2296 2446
rect 2267 2443 2268 2444
rect 2262 2442 2268 2443
rect 2295 2443 2296 2444
rect 2300 2443 2301 2447
rect 2295 2442 2301 2443
rect 2382 2447 2389 2448
rect 2406 2447 2412 2448
rect 2382 2443 2383 2447
rect 2388 2443 2389 2447
rect 2382 2442 2389 2443
rect 1974 2439 1980 2440
rect 1974 2438 1975 2439
rect 1793 2436 1975 2438
rect 1238 2434 1244 2435
rect 1278 2435 1284 2436
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 270 2432 276 2433
rect 270 2428 271 2432
rect 275 2428 276 2432
rect 270 2427 276 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 350 2432 356 2433
rect 350 2428 351 2432
rect 355 2428 356 2432
rect 350 2427 356 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 454 2432 460 2433
rect 454 2428 455 2432
rect 459 2428 460 2432
rect 454 2427 460 2428
rect 510 2432 516 2433
rect 510 2428 511 2432
rect 515 2428 516 2432
rect 510 2427 516 2428
rect 574 2432 580 2433
rect 574 2428 575 2432
rect 579 2428 580 2432
rect 574 2427 580 2428
rect 638 2432 644 2433
rect 638 2428 639 2432
rect 643 2428 644 2432
rect 638 2427 644 2428
rect 702 2432 708 2433
rect 702 2428 703 2432
rect 707 2428 708 2432
rect 702 2427 708 2428
rect 766 2432 772 2433
rect 766 2428 767 2432
rect 771 2428 772 2432
rect 766 2427 772 2428
rect 822 2432 828 2433
rect 822 2428 823 2432
rect 827 2428 828 2432
rect 822 2427 828 2428
rect 878 2432 884 2433
rect 878 2428 879 2432
rect 883 2428 884 2432
rect 878 2427 884 2428
rect 926 2432 932 2433
rect 926 2428 927 2432
rect 931 2428 932 2432
rect 926 2427 932 2428
rect 974 2432 980 2433
rect 974 2428 975 2432
rect 979 2428 980 2432
rect 974 2427 980 2428
rect 1022 2432 1028 2433
rect 1022 2428 1023 2432
rect 1027 2428 1028 2432
rect 1022 2427 1028 2428
rect 1070 2432 1076 2433
rect 1070 2428 1071 2432
rect 1075 2428 1076 2432
rect 1070 2427 1076 2428
rect 1110 2432 1116 2433
rect 1110 2428 1111 2432
rect 1115 2428 1116 2432
rect 1110 2427 1116 2428
rect 1150 2432 1156 2433
rect 1150 2428 1151 2432
rect 1155 2428 1156 2432
rect 1150 2427 1156 2428
rect 1190 2432 1196 2433
rect 1190 2428 1191 2432
rect 1195 2428 1196 2432
rect 1278 2431 1279 2435
rect 1283 2431 1284 2435
rect 1974 2435 1975 2436
rect 1979 2435 1980 2439
rect 1974 2434 1980 2435
rect 2406 2435 2412 2436
rect 1278 2430 1284 2431
rect 2406 2431 2407 2435
rect 2411 2431 2412 2435
rect 2406 2430 2412 2431
rect 1190 2427 1196 2428
rect 1302 2428 1308 2429
rect 1302 2424 1303 2428
rect 1307 2424 1308 2428
rect 1302 2423 1308 2424
rect 1342 2428 1348 2429
rect 1342 2424 1343 2428
rect 1347 2424 1348 2428
rect 1342 2423 1348 2424
rect 1382 2428 1388 2429
rect 1382 2424 1383 2428
rect 1387 2424 1388 2428
rect 1382 2423 1388 2424
rect 1438 2428 1444 2429
rect 1438 2424 1439 2428
rect 1443 2424 1444 2428
rect 1438 2423 1444 2424
rect 1510 2428 1516 2429
rect 1510 2424 1511 2428
rect 1515 2424 1516 2428
rect 1510 2423 1516 2424
rect 1582 2428 1588 2429
rect 1582 2424 1583 2428
rect 1587 2424 1588 2428
rect 1582 2423 1588 2424
rect 1662 2428 1668 2429
rect 1662 2424 1663 2428
rect 1667 2424 1668 2428
rect 1662 2423 1668 2424
rect 1734 2428 1740 2429
rect 1734 2424 1735 2428
rect 1739 2424 1740 2428
rect 1734 2423 1740 2424
rect 1806 2428 1812 2429
rect 1806 2424 1807 2428
rect 1811 2424 1812 2428
rect 1806 2423 1812 2424
rect 1886 2428 1892 2429
rect 1886 2424 1887 2428
rect 1891 2424 1892 2428
rect 1886 2423 1892 2424
rect 1966 2428 1972 2429
rect 1966 2424 1967 2428
rect 1971 2424 1972 2428
rect 1966 2423 1972 2424
rect 2062 2428 2068 2429
rect 2062 2424 2063 2428
rect 2067 2424 2068 2428
rect 2062 2423 2068 2424
rect 2166 2428 2172 2429
rect 2166 2424 2167 2428
rect 2171 2424 2172 2428
rect 2166 2423 2172 2424
rect 2270 2428 2276 2429
rect 2270 2424 2271 2428
rect 2275 2424 2276 2428
rect 2270 2423 2276 2424
rect 2358 2428 2364 2429
rect 2358 2424 2359 2428
rect 2363 2424 2364 2428
rect 2358 2423 2364 2424
rect 1374 2416 1380 2417
rect 198 2412 204 2413
rect 198 2408 199 2412
rect 203 2408 204 2412
rect 198 2407 204 2408
rect 262 2412 268 2413
rect 262 2408 263 2412
rect 267 2408 268 2412
rect 262 2407 268 2408
rect 326 2412 332 2413
rect 326 2408 327 2412
rect 331 2408 332 2412
rect 326 2407 332 2408
rect 398 2412 404 2413
rect 398 2408 399 2412
rect 403 2408 404 2412
rect 398 2407 404 2408
rect 470 2412 476 2413
rect 470 2408 471 2412
rect 475 2408 476 2412
rect 470 2407 476 2408
rect 542 2412 548 2413
rect 542 2408 543 2412
rect 547 2408 548 2412
rect 542 2407 548 2408
rect 614 2412 620 2413
rect 614 2408 615 2412
rect 619 2408 620 2412
rect 614 2407 620 2408
rect 686 2412 692 2413
rect 686 2408 687 2412
rect 691 2408 692 2412
rect 686 2407 692 2408
rect 750 2412 756 2413
rect 750 2408 751 2412
rect 755 2408 756 2412
rect 750 2407 756 2408
rect 822 2412 828 2413
rect 822 2408 823 2412
rect 827 2408 828 2412
rect 822 2407 828 2408
rect 894 2412 900 2413
rect 894 2408 895 2412
rect 899 2408 900 2412
rect 894 2407 900 2408
rect 966 2412 972 2413
rect 966 2408 967 2412
rect 971 2408 972 2412
rect 1374 2412 1375 2416
rect 1379 2412 1380 2416
rect 1374 2411 1380 2412
rect 1414 2416 1420 2417
rect 1414 2412 1415 2416
rect 1419 2412 1420 2416
rect 1414 2411 1420 2412
rect 1454 2416 1460 2417
rect 1454 2412 1455 2416
rect 1459 2412 1460 2416
rect 1454 2411 1460 2412
rect 1502 2416 1508 2417
rect 1502 2412 1503 2416
rect 1507 2412 1508 2416
rect 1502 2411 1508 2412
rect 1558 2416 1564 2417
rect 1558 2412 1559 2416
rect 1563 2412 1564 2416
rect 1558 2411 1564 2412
rect 1614 2416 1620 2417
rect 1614 2412 1615 2416
rect 1619 2412 1620 2416
rect 1614 2411 1620 2412
rect 1678 2416 1684 2417
rect 1678 2412 1679 2416
rect 1683 2412 1684 2416
rect 1678 2411 1684 2412
rect 1734 2416 1740 2417
rect 1734 2412 1735 2416
rect 1739 2412 1740 2416
rect 1734 2411 1740 2412
rect 1798 2416 1804 2417
rect 1798 2412 1799 2416
rect 1803 2412 1804 2416
rect 1798 2411 1804 2412
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 1950 2416 1956 2417
rect 1950 2412 1951 2416
rect 1955 2412 1956 2416
rect 1950 2411 1956 2412
rect 2046 2416 2052 2417
rect 2046 2412 2047 2416
rect 2051 2412 2052 2416
rect 2046 2411 2052 2412
rect 2150 2416 2156 2417
rect 2150 2412 2151 2416
rect 2155 2412 2156 2416
rect 2150 2411 2156 2412
rect 2262 2416 2268 2417
rect 2262 2412 2263 2416
rect 2267 2412 2268 2416
rect 2262 2411 2268 2412
rect 2358 2416 2364 2417
rect 2358 2412 2359 2416
rect 2363 2412 2364 2416
rect 2358 2411 2364 2412
rect 966 2407 972 2408
rect 1278 2409 1284 2410
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 110 2400 116 2401
rect 1238 2405 1244 2406
rect 1238 2401 1239 2405
rect 1243 2401 1244 2405
rect 1278 2405 1279 2409
rect 1283 2405 1284 2409
rect 1278 2404 1284 2405
rect 2406 2409 2412 2410
rect 2406 2405 2407 2409
rect 2411 2405 2412 2409
rect 2406 2404 2412 2405
rect 1686 2403 1692 2404
rect 1686 2402 1687 2403
rect 1238 2400 1244 2401
rect 1416 2400 1687 2402
rect 650 2399 656 2400
rect 650 2398 651 2399
rect 497 2396 651 2398
rect 497 2392 499 2396
rect 650 2395 651 2396
rect 655 2395 656 2399
rect 650 2394 656 2395
rect 1399 2395 1405 2396
rect 1278 2392 1284 2393
rect 223 2391 229 2392
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 223 2387 224 2391
rect 228 2390 229 2391
rect 278 2391 284 2392
rect 278 2390 279 2391
rect 228 2388 279 2390
rect 228 2387 229 2388
rect 223 2386 229 2387
rect 278 2387 279 2388
rect 283 2387 284 2391
rect 278 2386 284 2387
rect 287 2391 293 2392
rect 287 2387 288 2391
rect 292 2390 293 2391
rect 342 2391 348 2392
rect 342 2390 343 2391
rect 292 2388 343 2390
rect 292 2387 293 2388
rect 287 2386 293 2387
rect 342 2387 343 2388
rect 347 2387 348 2391
rect 342 2386 348 2387
rect 351 2391 357 2392
rect 351 2387 352 2391
rect 356 2390 357 2391
rect 414 2391 420 2392
rect 414 2390 415 2391
rect 356 2388 415 2390
rect 356 2387 357 2388
rect 351 2386 357 2387
rect 414 2387 415 2388
rect 419 2387 420 2391
rect 414 2386 420 2387
rect 422 2391 429 2392
rect 422 2387 423 2391
rect 428 2387 429 2391
rect 422 2386 429 2387
rect 495 2391 501 2392
rect 495 2387 496 2391
rect 500 2387 501 2391
rect 495 2386 501 2387
rect 503 2391 509 2392
rect 503 2387 504 2391
rect 508 2390 509 2391
rect 567 2391 573 2392
rect 567 2390 568 2391
rect 508 2388 568 2390
rect 508 2387 509 2388
rect 503 2386 509 2387
rect 567 2387 568 2388
rect 572 2387 573 2391
rect 567 2386 573 2387
rect 575 2391 581 2392
rect 575 2387 576 2391
rect 580 2390 581 2391
rect 639 2391 645 2392
rect 639 2390 640 2391
rect 580 2388 640 2390
rect 580 2387 581 2388
rect 575 2386 581 2387
rect 639 2387 640 2388
rect 644 2387 645 2391
rect 639 2386 645 2387
rect 647 2391 653 2392
rect 647 2387 648 2391
rect 652 2390 653 2391
rect 711 2391 717 2392
rect 711 2390 712 2391
rect 652 2388 712 2390
rect 652 2387 653 2388
rect 647 2386 653 2387
rect 711 2387 712 2388
rect 716 2387 717 2391
rect 711 2386 717 2387
rect 775 2391 781 2392
rect 775 2387 776 2391
rect 780 2390 781 2391
rect 838 2391 844 2392
rect 838 2390 839 2391
rect 780 2388 839 2390
rect 780 2387 781 2388
rect 775 2386 781 2387
rect 838 2387 839 2388
rect 843 2387 844 2391
rect 838 2386 844 2387
rect 847 2391 853 2392
rect 847 2387 848 2391
rect 852 2390 853 2391
rect 906 2391 912 2392
rect 852 2388 902 2390
rect 852 2387 853 2388
rect 847 2386 853 2387
rect 110 2383 116 2384
rect 900 2382 902 2388
rect 906 2387 907 2391
rect 911 2390 912 2391
rect 919 2391 925 2392
rect 919 2390 920 2391
rect 911 2388 920 2390
rect 911 2387 912 2388
rect 906 2386 912 2387
rect 919 2387 920 2388
rect 924 2387 925 2391
rect 919 2386 925 2387
rect 927 2391 933 2392
rect 927 2387 928 2391
rect 932 2390 933 2391
rect 991 2391 997 2392
rect 991 2390 992 2391
rect 932 2388 992 2390
rect 932 2387 933 2388
rect 927 2386 933 2387
rect 991 2387 992 2388
rect 996 2387 997 2391
rect 991 2386 997 2387
rect 1238 2388 1244 2389
rect 1238 2384 1239 2388
rect 1243 2384 1244 2388
rect 1278 2388 1279 2392
rect 1283 2388 1284 2392
rect 1399 2391 1400 2395
rect 1404 2394 1405 2395
rect 1416 2394 1418 2400
rect 1686 2399 1687 2400
rect 1691 2399 1692 2403
rect 1686 2398 1692 2399
rect 1404 2392 1418 2394
rect 1422 2395 1428 2396
rect 1404 2391 1405 2392
rect 1399 2390 1405 2391
rect 1422 2391 1423 2395
rect 1427 2394 1428 2395
rect 1439 2395 1445 2396
rect 1439 2394 1440 2395
rect 1427 2392 1440 2394
rect 1427 2391 1428 2392
rect 1422 2390 1428 2391
rect 1439 2391 1440 2392
rect 1444 2391 1445 2395
rect 1439 2390 1445 2391
rect 1462 2395 1468 2396
rect 1462 2391 1463 2395
rect 1467 2394 1468 2395
rect 1479 2395 1485 2396
rect 1479 2394 1480 2395
rect 1467 2392 1480 2394
rect 1467 2391 1468 2392
rect 1462 2390 1468 2391
rect 1479 2391 1480 2392
rect 1484 2391 1485 2395
rect 1479 2390 1485 2391
rect 1487 2395 1493 2396
rect 1487 2391 1488 2395
rect 1492 2394 1493 2395
rect 1527 2395 1533 2396
rect 1527 2394 1528 2395
rect 1492 2392 1528 2394
rect 1492 2391 1493 2392
rect 1487 2390 1493 2391
rect 1527 2391 1528 2392
rect 1532 2391 1533 2395
rect 1527 2390 1533 2391
rect 1535 2395 1541 2396
rect 1535 2391 1536 2395
rect 1540 2394 1541 2395
rect 1583 2395 1589 2396
rect 1583 2394 1584 2395
rect 1540 2392 1584 2394
rect 1540 2391 1541 2392
rect 1535 2390 1541 2391
rect 1583 2391 1584 2392
rect 1588 2391 1589 2395
rect 1583 2390 1589 2391
rect 1591 2395 1597 2396
rect 1591 2391 1592 2395
rect 1596 2394 1597 2395
rect 1639 2395 1645 2396
rect 1639 2394 1640 2395
rect 1596 2392 1640 2394
rect 1596 2391 1597 2392
rect 1591 2390 1597 2391
rect 1639 2391 1640 2392
rect 1644 2391 1645 2395
rect 1639 2390 1645 2391
rect 1647 2395 1653 2396
rect 1647 2391 1648 2395
rect 1652 2394 1653 2395
rect 1703 2395 1709 2396
rect 1703 2394 1704 2395
rect 1652 2392 1704 2394
rect 1652 2391 1653 2392
rect 1647 2390 1653 2391
rect 1703 2391 1704 2392
rect 1708 2391 1709 2395
rect 1703 2390 1709 2391
rect 1759 2395 1765 2396
rect 1759 2391 1760 2395
rect 1764 2391 1765 2395
rect 1759 2390 1765 2391
rect 1767 2395 1773 2396
rect 1767 2391 1768 2395
rect 1772 2394 1773 2395
rect 1823 2395 1829 2396
rect 1823 2394 1824 2395
rect 1772 2392 1824 2394
rect 1772 2391 1773 2392
rect 1767 2390 1773 2391
rect 1823 2391 1824 2392
rect 1828 2391 1829 2395
rect 1823 2390 1829 2391
rect 1831 2395 1837 2396
rect 1831 2391 1832 2395
rect 1836 2394 1837 2395
rect 1895 2395 1901 2396
rect 1895 2394 1896 2395
rect 1836 2392 1896 2394
rect 1836 2391 1837 2392
rect 1831 2390 1837 2391
rect 1895 2391 1896 2392
rect 1900 2391 1901 2395
rect 1895 2390 1901 2391
rect 1903 2395 1909 2396
rect 1903 2391 1904 2395
rect 1908 2394 1909 2395
rect 1975 2395 1981 2396
rect 1975 2394 1976 2395
rect 1908 2392 1976 2394
rect 1908 2391 1909 2392
rect 1903 2390 1909 2391
rect 1975 2391 1976 2392
rect 1980 2391 1981 2395
rect 1975 2390 1981 2391
rect 2071 2395 2077 2396
rect 2071 2391 2072 2395
rect 2076 2391 2077 2395
rect 2071 2390 2077 2391
rect 2079 2395 2085 2396
rect 2079 2391 2080 2395
rect 2084 2394 2085 2395
rect 2175 2395 2181 2396
rect 2175 2394 2176 2395
rect 2084 2392 2176 2394
rect 2084 2391 2085 2392
rect 2079 2390 2085 2391
rect 2175 2391 2176 2392
rect 2180 2391 2181 2395
rect 2175 2390 2181 2391
rect 2286 2395 2293 2396
rect 2286 2391 2287 2395
rect 2292 2391 2293 2395
rect 2286 2390 2293 2391
rect 2383 2395 2389 2396
rect 2383 2391 2384 2395
rect 2388 2394 2389 2395
rect 2391 2395 2397 2396
rect 2391 2394 2392 2395
rect 2388 2392 2392 2394
rect 2388 2391 2389 2392
rect 2383 2390 2389 2391
rect 2391 2391 2392 2392
rect 2396 2391 2397 2395
rect 2391 2390 2397 2391
rect 2406 2392 2412 2393
rect 1278 2387 1284 2388
rect 1760 2386 1762 2390
rect 1902 2387 1908 2388
rect 1902 2386 1903 2387
rect 1760 2384 1903 2386
rect 990 2383 996 2384
rect 1238 2383 1244 2384
rect 1902 2383 1903 2384
rect 1907 2383 1908 2387
rect 2072 2386 2074 2390
rect 2406 2388 2407 2392
rect 2411 2388 2412 2392
rect 2286 2387 2292 2388
rect 2406 2387 2412 2388
rect 2286 2386 2287 2387
rect 2072 2384 2287 2386
rect 990 2382 991 2383
rect 900 2380 991 2382
rect 990 2379 991 2380
rect 995 2379 996 2383
rect 1902 2382 1908 2383
rect 2286 2383 2287 2384
rect 2291 2383 2292 2387
rect 2286 2382 2292 2383
rect 990 2378 996 2379
rect 1374 2369 1380 2370
rect 198 2365 204 2366
rect 198 2361 199 2365
rect 203 2361 204 2365
rect 198 2360 204 2361
rect 262 2365 268 2366
rect 262 2361 263 2365
rect 267 2361 268 2365
rect 262 2360 268 2361
rect 326 2365 332 2366
rect 326 2361 327 2365
rect 331 2361 332 2365
rect 326 2360 332 2361
rect 398 2365 404 2366
rect 398 2361 399 2365
rect 403 2361 404 2365
rect 398 2360 404 2361
rect 470 2365 476 2366
rect 470 2361 471 2365
rect 475 2361 476 2365
rect 470 2360 476 2361
rect 542 2365 548 2366
rect 542 2361 543 2365
rect 547 2361 548 2365
rect 542 2360 548 2361
rect 614 2365 620 2366
rect 614 2361 615 2365
rect 619 2361 620 2365
rect 614 2360 620 2361
rect 686 2365 692 2366
rect 686 2361 687 2365
rect 691 2361 692 2365
rect 686 2360 692 2361
rect 750 2365 756 2366
rect 750 2361 751 2365
rect 755 2361 756 2365
rect 750 2360 756 2361
rect 822 2365 828 2366
rect 822 2361 823 2365
rect 827 2361 828 2365
rect 822 2360 828 2361
rect 894 2365 900 2366
rect 894 2361 895 2365
rect 899 2361 900 2365
rect 894 2360 900 2361
rect 966 2365 972 2366
rect 966 2361 967 2365
rect 971 2361 972 2365
rect 1374 2365 1375 2369
rect 1379 2365 1380 2369
rect 1374 2364 1380 2365
rect 1414 2369 1420 2370
rect 1414 2365 1415 2369
rect 1419 2365 1420 2369
rect 1414 2364 1420 2365
rect 1454 2369 1460 2370
rect 1454 2365 1455 2369
rect 1459 2365 1460 2369
rect 1454 2364 1460 2365
rect 1502 2369 1508 2370
rect 1502 2365 1503 2369
rect 1507 2365 1508 2369
rect 1502 2364 1508 2365
rect 1558 2369 1564 2370
rect 1558 2365 1559 2369
rect 1563 2365 1564 2369
rect 1558 2364 1564 2365
rect 1614 2369 1620 2370
rect 1614 2365 1615 2369
rect 1619 2365 1620 2369
rect 1614 2364 1620 2365
rect 1678 2369 1684 2370
rect 1678 2365 1679 2369
rect 1683 2365 1684 2369
rect 1678 2364 1684 2365
rect 1734 2369 1740 2370
rect 1734 2365 1735 2369
rect 1739 2365 1740 2369
rect 1734 2364 1740 2365
rect 1798 2369 1804 2370
rect 1798 2365 1799 2369
rect 1803 2365 1804 2369
rect 1798 2364 1804 2365
rect 1870 2369 1876 2370
rect 1870 2365 1871 2369
rect 1875 2365 1876 2369
rect 1870 2364 1876 2365
rect 1950 2369 1956 2370
rect 1950 2365 1951 2369
rect 1955 2365 1956 2369
rect 1950 2364 1956 2365
rect 2046 2369 2052 2370
rect 2046 2365 2047 2369
rect 2051 2365 2052 2369
rect 2046 2364 2052 2365
rect 2150 2369 2156 2370
rect 2150 2365 2151 2369
rect 2155 2365 2156 2369
rect 2150 2364 2156 2365
rect 2262 2369 2268 2370
rect 2262 2365 2263 2369
rect 2267 2365 2268 2369
rect 2262 2364 2268 2365
rect 2358 2369 2364 2370
rect 2358 2365 2359 2369
rect 2363 2365 2364 2369
rect 2358 2364 2364 2365
rect 966 2360 972 2361
rect 1399 2363 1405 2364
rect 223 2359 229 2360
rect 223 2355 224 2359
rect 228 2358 229 2359
rect 242 2359 248 2360
rect 242 2358 243 2359
rect 228 2356 243 2358
rect 228 2355 229 2356
rect 223 2354 229 2355
rect 242 2355 243 2356
rect 247 2355 248 2359
rect 242 2354 248 2355
rect 278 2359 284 2360
rect 278 2355 279 2359
rect 283 2358 284 2359
rect 287 2359 293 2360
rect 287 2358 288 2359
rect 283 2356 288 2358
rect 283 2355 284 2356
rect 278 2354 284 2355
rect 287 2355 288 2356
rect 292 2355 293 2359
rect 287 2354 293 2355
rect 342 2359 348 2360
rect 342 2355 343 2359
rect 347 2358 348 2359
rect 351 2359 357 2360
rect 351 2358 352 2359
rect 347 2356 352 2358
rect 347 2355 348 2356
rect 342 2354 348 2355
rect 351 2355 352 2356
rect 356 2355 357 2359
rect 351 2354 357 2355
rect 414 2359 420 2360
rect 414 2355 415 2359
rect 419 2358 420 2359
rect 423 2359 429 2360
rect 423 2358 424 2359
rect 419 2356 424 2358
rect 419 2355 420 2356
rect 414 2354 420 2355
rect 423 2355 424 2356
rect 428 2355 429 2359
rect 423 2354 429 2355
rect 495 2359 501 2360
rect 495 2355 496 2359
rect 500 2358 501 2359
rect 503 2359 509 2360
rect 503 2358 504 2359
rect 500 2356 504 2358
rect 500 2355 501 2356
rect 495 2354 501 2355
rect 503 2355 504 2356
rect 508 2355 509 2359
rect 503 2354 509 2355
rect 567 2359 573 2360
rect 567 2355 568 2359
rect 572 2358 573 2359
rect 575 2359 581 2360
rect 575 2358 576 2359
rect 572 2356 576 2358
rect 572 2355 573 2356
rect 567 2354 573 2355
rect 575 2355 576 2356
rect 580 2355 581 2359
rect 575 2354 581 2355
rect 639 2359 645 2360
rect 639 2355 640 2359
rect 644 2358 645 2359
rect 647 2359 653 2360
rect 647 2358 648 2359
rect 644 2356 648 2358
rect 644 2355 645 2356
rect 639 2354 645 2355
rect 647 2355 648 2356
rect 652 2355 653 2359
rect 647 2354 653 2355
rect 711 2359 717 2360
rect 711 2355 712 2359
rect 716 2358 717 2359
rect 734 2359 740 2360
rect 734 2358 735 2359
rect 716 2356 735 2358
rect 716 2355 717 2356
rect 711 2354 717 2355
rect 734 2355 735 2356
rect 739 2355 740 2359
rect 734 2354 740 2355
rect 774 2359 781 2360
rect 774 2355 775 2359
rect 780 2355 781 2359
rect 774 2354 781 2355
rect 838 2359 844 2360
rect 838 2355 839 2359
rect 843 2358 844 2359
rect 847 2359 853 2360
rect 847 2358 848 2359
rect 843 2356 848 2358
rect 843 2355 844 2356
rect 838 2354 844 2355
rect 847 2355 848 2356
rect 852 2355 853 2359
rect 847 2354 853 2355
rect 919 2359 925 2360
rect 919 2355 920 2359
rect 924 2358 925 2359
rect 927 2359 933 2360
rect 927 2358 928 2359
rect 924 2356 928 2358
rect 924 2355 925 2356
rect 919 2354 925 2355
rect 927 2355 928 2356
rect 932 2355 933 2359
rect 927 2354 933 2355
rect 990 2359 997 2360
rect 990 2355 991 2359
rect 996 2355 997 2359
rect 1399 2359 1400 2363
rect 1404 2362 1405 2363
rect 1422 2363 1428 2364
rect 1422 2362 1423 2363
rect 1404 2360 1423 2362
rect 1404 2359 1405 2360
rect 1399 2358 1405 2359
rect 1422 2359 1423 2360
rect 1427 2359 1428 2363
rect 1422 2358 1428 2359
rect 1439 2363 1445 2364
rect 1439 2359 1440 2363
rect 1444 2362 1445 2363
rect 1462 2363 1468 2364
rect 1462 2362 1463 2363
rect 1444 2360 1463 2362
rect 1444 2359 1445 2360
rect 1439 2358 1445 2359
rect 1462 2359 1463 2360
rect 1467 2359 1468 2363
rect 1462 2358 1468 2359
rect 1479 2363 1485 2364
rect 1479 2359 1480 2363
rect 1484 2362 1485 2363
rect 1487 2363 1493 2364
rect 1487 2362 1488 2363
rect 1484 2360 1488 2362
rect 1484 2359 1485 2360
rect 1479 2358 1485 2359
rect 1487 2359 1488 2360
rect 1492 2359 1493 2363
rect 1487 2358 1493 2359
rect 1527 2363 1533 2364
rect 1527 2359 1528 2363
rect 1532 2362 1533 2363
rect 1535 2363 1541 2364
rect 1535 2362 1536 2363
rect 1532 2360 1536 2362
rect 1532 2359 1533 2360
rect 1527 2358 1533 2359
rect 1535 2359 1536 2360
rect 1540 2359 1541 2363
rect 1535 2358 1541 2359
rect 1583 2363 1589 2364
rect 1583 2359 1584 2363
rect 1588 2362 1589 2363
rect 1591 2363 1597 2364
rect 1591 2362 1592 2363
rect 1588 2360 1592 2362
rect 1588 2359 1589 2360
rect 1583 2358 1589 2359
rect 1591 2359 1592 2360
rect 1596 2359 1597 2363
rect 1591 2358 1597 2359
rect 1639 2363 1645 2364
rect 1639 2359 1640 2363
rect 1644 2362 1645 2363
rect 1647 2363 1653 2364
rect 1647 2362 1648 2363
rect 1644 2360 1648 2362
rect 1644 2359 1645 2360
rect 1639 2358 1645 2359
rect 1647 2359 1648 2360
rect 1652 2359 1653 2363
rect 1647 2358 1653 2359
rect 1658 2363 1664 2364
rect 1658 2359 1659 2363
rect 1663 2362 1664 2363
rect 1703 2363 1709 2364
rect 1703 2362 1704 2363
rect 1663 2360 1704 2362
rect 1663 2359 1664 2360
rect 1658 2358 1664 2359
rect 1703 2359 1704 2360
rect 1708 2359 1709 2363
rect 1703 2358 1709 2359
rect 1759 2363 1765 2364
rect 1759 2359 1760 2363
rect 1764 2362 1765 2363
rect 1767 2363 1773 2364
rect 1767 2362 1768 2363
rect 1764 2360 1768 2362
rect 1764 2359 1765 2360
rect 1759 2358 1765 2359
rect 1767 2359 1768 2360
rect 1772 2359 1773 2363
rect 1767 2358 1773 2359
rect 1823 2363 1829 2364
rect 1823 2359 1824 2363
rect 1828 2362 1829 2363
rect 1831 2363 1837 2364
rect 1831 2362 1832 2363
rect 1828 2360 1832 2362
rect 1828 2359 1829 2360
rect 1823 2358 1829 2359
rect 1831 2359 1832 2360
rect 1836 2359 1837 2363
rect 1831 2358 1837 2359
rect 1895 2363 1901 2364
rect 1895 2359 1896 2363
rect 1900 2362 1901 2363
rect 1903 2363 1909 2364
rect 1903 2362 1904 2363
rect 1900 2360 1904 2362
rect 1900 2359 1901 2360
rect 1895 2358 1901 2359
rect 1903 2359 1904 2360
rect 1908 2359 1909 2363
rect 1903 2358 1909 2359
rect 1974 2363 1981 2364
rect 1974 2359 1975 2363
rect 1980 2359 1981 2363
rect 1974 2358 1981 2359
rect 2071 2363 2077 2364
rect 2071 2359 2072 2363
rect 2076 2362 2077 2363
rect 2079 2363 2085 2364
rect 2079 2362 2080 2363
rect 2076 2360 2080 2362
rect 2076 2359 2077 2360
rect 2071 2358 2077 2359
rect 2079 2359 2080 2360
rect 2084 2359 2085 2363
rect 2079 2358 2085 2359
rect 2175 2363 2181 2364
rect 2175 2359 2176 2363
rect 2180 2362 2181 2363
rect 2186 2363 2192 2364
rect 2186 2362 2187 2363
rect 2180 2360 2187 2362
rect 2180 2359 2181 2360
rect 2175 2358 2181 2359
rect 2186 2359 2187 2360
rect 2191 2359 2192 2363
rect 2186 2358 2192 2359
rect 2286 2363 2293 2364
rect 2286 2359 2287 2363
rect 2292 2359 2293 2363
rect 2286 2358 2293 2359
rect 2382 2363 2389 2364
rect 2382 2359 2383 2363
rect 2388 2359 2389 2363
rect 2382 2358 2389 2359
rect 990 2354 997 2355
rect 1351 2339 1360 2340
rect 295 2335 301 2336
rect 270 2331 276 2332
rect 270 2327 271 2331
rect 275 2327 276 2331
rect 295 2331 296 2335
rect 300 2334 301 2335
rect 318 2335 324 2336
rect 318 2334 319 2335
rect 300 2332 319 2334
rect 300 2331 301 2332
rect 295 2330 301 2331
rect 318 2331 319 2332
rect 323 2331 324 2335
rect 351 2335 357 2336
rect 318 2330 324 2331
rect 326 2331 332 2332
rect 270 2326 276 2327
rect 326 2327 327 2331
rect 331 2327 332 2331
rect 351 2331 352 2335
rect 356 2334 357 2335
rect 390 2335 396 2336
rect 390 2334 391 2335
rect 356 2332 391 2334
rect 356 2331 357 2332
rect 351 2330 357 2331
rect 390 2331 391 2332
rect 395 2331 396 2335
rect 422 2335 429 2336
rect 390 2330 396 2331
rect 398 2331 404 2332
rect 326 2326 332 2327
rect 398 2327 399 2331
rect 403 2327 404 2331
rect 422 2331 423 2335
rect 428 2331 429 2335
rect 482 2335 488 2336
rect 422 2330 429 2331
rect 470 2331 476 2332
rect 398 2326 404 2327
rect 470 2327 471 2331
rect 475 2327 476 2331
rect 482 2331 483 2335
rect 487 2334 488 2335
rect 495 2335 501 2336
rect 495 2334 496 2335
rect 487 2332 496 2334
rect 487 2331 488 2332
rect 482 2330 488 2331
rect 495 2331 496 2332
rect 500 2331 501 2335
rect 562 2335 568 2336
rect 495 2330 501 2331
rect 550 2331 556 2332
rect 470 2326 476 2327
rect 550 2327 551 2331
rect 555 2327 556 2331
rect 562 2331 563 2335
rect 567 2334 568 2335
rect 575 2335 581 2336
rect 575 2334 576 2335
rect 567 2332 576 2334
rect 567 2331 568 2332
rect 562 2330 568 2331
rect 575 2331 576 2332
rect 580 2331 581 2335
rect 655 2335 661 2336
rect 575 2330 581 2331
rect 630 2331 636 2332
rect 550 2326 556 2327
rect 630 2327 631 2331
rect 635 2327 636 2331
rect 655 2331 656 2335
rect 660 2334 661 2335
rect 670 2335 676 2336
rect 670 2334 671 2335
rect 660 2332 671 2334
rect 660 2331 661 2332
rect 655 2330 661 2331
rect 670 2331 671 2332
rect 675 2331 676 2335
rect 722 2335 728 2336
rect 670 2330 676 2331
rect 710 2331 716 2332
rect 630 2326 636 2327
rect 710 2327 711 2331
rect 715 2327 716 2331
rect 722 2331 723 2335
rect 727 2334 728 2335
rect 735 2335 741 2336
rect 735 2334 736 2335
rect 727 2332 736 2334
rect 727 2331 728 2332
rect 722 2330 728 2331
rect 735 2331 736 2332
rect 740 2331 741 2335
rect 807 2335 813 2336
rect 735 2330 741 2331
rect 782 2331 788 2332
rect 710 2326 716 2327
rect 782 2327 783 2331
rect 787 2327 788 2331
rect 807 2331 808 2335
rect 812 2334 813 2335
rect 846 2335 852 2336
rect 846 2334 847 2335
rect 812 2332 847 2334
rect 812 2331 813 2332
rect 807 2330 813 2331
rect 846 2331 847 2332
rect 851 2331 852 2335
rect 879 2335 885 2336
rect 846 2330 852 2331
rect 854 2331 860 2332
rect 782 2326 788 2327
rect 854 2327 855 2331
rect 859 2327 860 2331
rect 879 2331 880 2335
rect 884 2334 885 2335
rect 906 2335 912 2336
rect 906 2334 907 2335
rect 884 2332 907 2334
rect 884 2331 885 2332
rect 879 2330 885 2331
rect 906 2331 907 2332
rect 911 2331 912 2335
rect 930 2335 936 2336
rect 906 2330 912 2331
rect 918 2331 924 2332
rect 854 2326 860 2327
rect 918 2327 919 2331
rect 923 2327 924 2331
rect 930 2331 931 2335
rect 935 2334 936 2335
rect 943 2335 949 2336
rect 943 2334 944 2335
rect 935 2332 944 2334
rect 935 2331 936 2332
rect 930 2330 936 2331
rect 943 2331 944 2332
rect 948 2331 949 2335
rect 1015 2335 1021 2336
rect 943 2330 949 2331
rect 990 2331 996 2332
rect 918 2326 924 2327
rect 990 2327 991 2331
rect 995 2327 996 2331
rect 1015 2331 1016 2335
rect 1020 2334 1021 2335
rect 1054 2335 1060 2336
rect 1054 2334 1055 2335
rect 1020 2332 1055 2334
rect 1020 2331 1021 2332
rect 1015 2330 1021 2331
rect 1054 2331 1055 2332
rect 1059 2331 1060 2335
rect 1074 2335 1080 2336
rect 1054 2330 1060 2331
rect 1062 2331 1068 2332
rect 990 2326 996 2327
rect 1062 2327 1063 2331
rect 1067 2327 1068 2331
rect 1074 2331 1075 2335
rect 1079 2334 1080 2335
rect 1087 2335 1093 2336
rect 1087 2334 1088 2335
rect 1079 2332 1088 2334
rect 1079 2331 1080 2332
rect 1074 2330 1080 2331
rect 1087 2331 1088 2332
rect 1092 2331 1093 2335
rect 1087 2330 1093 2331
rect 1326 2335 1332 2336
rect 1326 2331 1327 2335
rect 1331 2331 1332 2335
rect 1351 2335 1352 2339
rect 1359 2335 1360 2339
rect 1394 2339 1400 2340
rect 1351 2334 1360 2335
rect 1382 2335 1388 2336
rect 1326 2330 1332 2331
rect 1382 2331 1383 2335
rect 1387 2331 1388 2335
rect 1394 2335 1395 2339
rect 1399 2338 1400 2339
rect 1407 2339 1413 2340
rect 1407 2338 1408 2339
rect 1399 2336 1408 2338
rect 1399 2335 1400 2336
rect 1394 2334 1400 2335
rect 1407 2335 1408 2336
rect 1412 2335 1413 2339
rect 1450 2339 1456 2340
rect 1407 2334 1413 2335
rect 1438 2335 1444 2336
rect 1382 2330 1388 2331
rect 1438 2331 1439 2335
rect 1443 2331 1444 2335
rect 1450 2335 1451 2339
rect 1455 2338 1456 2339
rect 1463 2339 1469 2340
rect 1463 2338 1464 2339
rect 1455 2336 1464 2338
rect 1455 2335 1456 2336
rect 1450 2334 1456 2335
rect 1463 2335 1464 2336
rect 1468 2335 1469 2339
rect 1514 2339 1520 2340
rect 1463 2334 1469 2335
rect 1502 2335 1508 2336
rect 1438 2330 1444 2331
rect 1502 2331 1503 2335
rect 1507 2331 1508 2335
rect 1514 2335 1515 2339
rect 1519 2338 1520 2339
rect 1527 2339 1533 2340
rect 1527 2338 1528 2339
rect 1519 2336 1528 2338
rect 1519 2335 1520 2336
rect 1514 2334 1520 2335
rect 1527 2335 1528 2336
rect 1532 2335 1533 2339
rect 1586 2339 1592 2340
rect 1527 2334 1533 2335
rect 1574 2335 1580 2336
rect 1502 2330 1508 2331
rect 1574 2331 1575 2335
rect 1579 2331 1580 2335
rect 1586 2335 1587 2339
rect 1591 2338 1592 2339
rect 1599 2339 1605 2340
rect 1599 2338 1600 2339
rect 1591 2336 1600 2338
rect 1591 2335 1592 2336
rect 1586 2334 1592 2335
rect 1599 2335 1600 2336
rect 1604 2335 1605 2339
rect 1671 2339 1677 2340
rect 1599 2334 1605 2335
rect 1646 2335 1652 2336
rect 1574 2330 1580 2331
rect 1646 2331 1647 2335
rect 1651 2331 1652 2335
rect 1671 2335 1672 2339
rect 1676 2338 1677 2339
rect 1710 2339 1716 2340
rect 1710 2338 1711 2339
rect 1676 2336 1711 2338
rect 1676 2335 1677 2336
rect 1671 2334 1677 2335
rect 1710 2335 1711 2336
rect 1715 2335 1716 2339
rect 1743 2339 1749 2340
rect 1710 2334 1716 2335
rect 1718 2335 1724 2336
rect 1646 2330 1652 2331
rect 1718 2331 1719 2335
rect 1723 2331 1724 2335
rect 1743 2335 1744 2339
rect 1748 2338 1749 2339
rect 1790 2339 1796 2340
rect 1790 2338 1791 2339
rect 1748 2336 1791 2338
rect 1748 2335 1749 2336
rect 1743 2334 1749 2335
rect 1790 2335 1791 2336
rect 1795 2335 1796 2339
rect 1823 2339 1829 2340
rect 1790 2334 1796 2335
rect 1798 2335 1804 2336
rect 1718 2330 1724 2331
rect 1798 2331 1799 2335
rect 1803 2331 1804 2335
rect 1823 2335 1824 2339
rect 1828 2338 1829 2339
rect 1870 2339 1876 2340
rect 1870 2338 1871 2339
rect 1828 2336 1871 2338
rect 1828 2335 1829 2336
rect 1823 2334 1829 2335
rect 1870 2335 1871 2336
rect 1875 2335 1876 2339
rect 1902 2339 1909 2340
rect 1870 2334 1876 2335
rect 1878 2335 1884 2336
rect 1798 2330 1804 2331
rect 1878 2331 1879 2335
rect 1883 2331 1884 2335
rect 1902 2335 1903 2339
rect 1908 2335 1909 2339
rect 1978 2339 1984 2340
rect 1902 2334 1909 2335
rect 1966 2335 1972 2336
rect 1878 2330 1884 2331
rect 1966 2331 1967 2335
rect 1971 2331 1972 2335
rect 1978 2335 1979 2339
rect 1983 2338 1984 2339
rect 1991 2339 1997 2340
rect 1991 2338 1992 2339
rect 1983 2336 1992 2338
rect 1983 2335 1984 2336
rect 1978 2334 1984 2335
rect 1991 2335 1992 2336
rect 1996 2335 1997 2339
rect 2074 2339 2080 2340
rect 1991 2334 1997 2335
rect 2062 2335 2068 2336
rect 1966 2330 1972 2331
rect 2062 2331 2063 2335
rect 2067 2331 2068 2335
rect 2074 2335 2075 2339
rect 2079 2338 2080 2339
rect 2087 2339 2093 2340
rect 2087 2338 2088 2339
rect 2079 2336 2088 2338
rect 2079 2335 2080 2336
rect 2074 2334 2080 2335
rect 2087 2335 2088 2336
rect 2092 2335 2093 2339
rect 2178 2339 2184 2340
rect 2087 2334 2093 2335
rect 2166 2335 2172 2336
rect 2062 2330 2068 2331
rect 2166 2331 2167 2335
rect 2171 2331 2172 2335
rect 2178 2335 2179 2339
rect 2183 2338 2184 2339
rect 2191 2339 2197 2340
rect 2191 2338 2192 2339
rect 2183 2336 2192 2338
rect 2183 2335 2184 2336
rect 2178 2334 2184 2335
rect 2191 2335 2192 2336
rect 2196 2335 2197 2339
rect 2295 2339 2301 2340
rect 2191 2334 2197 2335
rect 2270 2335 2276 2336
rect 2166 2330 2172 2331
rect 2270 2331 2271 2335
rect 2275 2331 2276 2335
rect 2295 2335 2296 2339
rect 2300 2338 2301 2339
rect 2350 2339 2356 2340
rect 2350 2338 2351 2339
rect 2300 2336 2351 2338
rect 2300 2335 2301 2336
rect 2295 2334 2301 2335
rect 2350 2335 2351 2336
rect 2355 2335 2356 2339
rect 2383 2339 2389 2340
rect 2350 2334 2356 2335
rect 2358 2335 2364 2336
rect 2270 2330 2276 2331
rect 2358 2331 2359 2335
rect 2363 2331 2364 2335
rect 2383 2335 2384 2339
rect 2388 2338 2389 2339
rect 2391 2339 2397 2340
rect 2391 2338 2392 2339
rect 2388 2336 2392 2338
rect 2388 2335 2389 2336
rect 2383 2334 2389 2335
rect 2391 2335 2392 2336
rect 2396 2335 2397 2339
rect 2391 2334 2397 2335
rect 2358 2330 2364 2331
rect 1062 2326 1068 2327
rect 1278 2312 1284 2313
rect 482 2311 488 2312
rect 482 2310 483 2311
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 308 2308 483 2310
rect 110 2303 116 2304
rect 295 2303 301 2304
rect 295 2299 296 2303
rect 300 2302 301 2303
rect 308 2302 310 2308
rect 482 2307 483 2308
rect 487 2307 488 2311
rect 930 2311 936 2312
rect 930 2310 931 2311
rect 482 2306 488 2307
rect 840 2308 931 2310
rect 300 2300 310 2302
rect 318 2303 324 2304
rect 300 2299 301 2300
rect 295 2298 301 2299
rect 318 2299 319 2303
rect 323 2302 324 2303
rect 351 2303 357 2304
rect 351 2302 352 2303
rect 323 2300 352 2302
rect 323 2299 324 2300
rect 318 2298 324 2299
rect 351 2299 352 2300
rect 356 2299 357 2303
rect 351 2298 357 2299
rect 390 2303 396 2304
rect 390 2299 391 2303
rect 395 2302 396 2303
rect 423 2303 429 2304
rect 423 2302 424 2303
rect 395 2300 424 2302
rect 395 2299 396 2300
rect 390 2298 396 2299
rect 423 2299 424 2300
rect 428 2299 429 2303
rect 423 2298 429 2299
rect 495 2303 501 2304
rect 495 2299 496 2303
rect 500 2302 501 2303
rect 562 2303 568 2304
rect 562 2302 563 2303
rect 500 2300 563 2302
rect 500 2299 501 2300
rect 495 2298 501 2299
rect 562 2299 563 2300
rect 567 2299 568 2303
rect 562 2298 568 2299
rect 575 2303 584 2304
rect 575 2299 576 2303
rect 583 2299 584 2303
rect 575 2298 584 2299
rect 655 2303 661 2304
rect 655 2299 656 2303
rect 660 2302 661 2303
rect 722 2303 728 2304
rect 722 2302 723 2303
rect 660 2300 723 2302
rect 660 2299 661 2300
rect 655 2298 661 2299
rect 722 2299 723 2300
rect 727 2299 728 2303
rect 722 2298 728 2299
rect 734 2303 741 2304
rect 734 2299 735 2303
rect 740 2299 741 2303
rect 734 2298 741 2299
rect 807 2303 813 2304
rect 807 2299 808 2303
rect 812 2302 813 2303
rect 840 2302 842 2308
rect 930 2307 931 2308
rect 935 2307 936 2311
rect 1074 2311 1080 2312
rect 1074 2310 1075 2311
rect 930 2306 936 2307
rect 1001 2308 1075 2310
rect 812 2300 842 2302
rect 846 2303 852 2304
rect 812 2299 813 2300
rect 807 2298 813 2299
rect 846 2299 847 2303
rect 851 2302 852 2303
rect 879 2303 885 2304
rect 879 2302 880 2303
rect 851 2300 880 2302
rect 851 2299 852 2300
rect 846 2298 852 2299
rect 879 2299 880 2300
rect 884 2299 885 2303
rect 879 2298 885 2299
rect 943 2303 949 2304
rect 943 2299 944 2303
rect 948 2302 949 2303
rect 1001 2302 1003 2308
rect 1074 2307 1075 2308
rect 1079 2307 1080 2311
rect 1074 2306 1080 2307
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1278 2308 1279 2312
rect 1283 2308 1284 2312
rect 2406 2312 2412 2313
rect 2406 2308 2407 2312
rect 2411 2308 2412 2312
rect 1278 2307 1284 2308
rect 1351 2307 1357 2308
rect 948 2300 1003 2302
rect 1006 2303 1012 2304
rect 948 2299 949 2300
rect 943 2298 949 2299
rect 1006 2299 1007 2303
rect 1011 2302 1012 2303
rect 1015 2303 1021 2304
rect 1015 2302 1016 2303
rect 1011 2300 1016 2302
rect 1011 2299 1012 2300
rect 1006 2298 1012 2299
rect 1015 2299 1016 2300
rect 1020 2299 1021 2303
rect 1015 2298 1021 2299
rect 1054 2303 1060 2304
rect 1054 2299 1055 2303
rect 1059 2302 1060 2303
rect 1087 2303 1093 2304
rect 1238 2303 1244 2304
rect 1351 2303 1352 2307
rect 1356 2306 1357 2307
rect 1394 2307 1400 2308
rect 1394 2306 1395 2307
rect 1356 2304 1395 2306
rect 1356 2303 1357 2304
rect 1087 2302 1088 2303
rect 1059 2300 1088 2302
rect 1059 2299 1060 2300
rect 1054 2298 1060 2299
rect 1087 2299 1088 2300
rect 1092 2299 1093 2303
rect 1351 2302 1357 2303
rect 1394 2303 1395 2304
rect 1399 2303 1400 2307
rect 1394 2302 1400 2303
rect 1407 2307 1413 2308
rect 1407 2303 1408 2307
rect 1412 2306 1413 2307
rect 1450 2307 1456 2308
rect 1450 2306 1451 2307
rect 1412 2304 1451 2306
rect 1412 2303 1413 2304
rect 1407 2302 1413 2303
rect 1450 2303 1451 2304
rect 1455 2303 1456 2307
rect 1450 2302 1456 2303
rect 1463 2307 1469 2308
rect 1463 2303 1464 2307
rect 1468 2306 1469 2307
rect 1514 2307 1520 2308
rect 1514 2306 1515 2307
rect 1468 2304 1515 2306
rect 1468 2303 1469 2304
rect 1463 2302 1469 2303
rect 1514 2303 1515 2304
rect 1519 2303 1520 2307
rect 1514 2302 1520 2303
rect 1527 2307 1533 2308
rect 1527 2303 1528 2307
rect 1532 2306 1533 2307
rect 1586 2307 1592 2308
rect 1586 2306 1587 2307
rect 1532 2304 1587 2306
rect 1532 2303 1533 2304
rect 1527 2302 1533 2303
rect 1586 2303 1587 2304
rect 1591 2303 1592 2307
rect 1586 2302 1592 2303
rect 1599 2307 1605 2308
rect 1599 2303 1600 2307
rect 1604 2306 1605 2307
rect 1658 2307 1664 2308
rect 1658 2306 1659 2307
rect 1604 2304 1659 2306
rect 1604 2303 1605 2304
rect 1599 2302 1605 2303
rect 1658 2303 1659 2304
rect 1663 2303 1664 2307
rect 1658 2302 1664 2303
rect 1671 2307 1677 2308
rect 1671 2303 1672 2307
rect 1676 2306 1677 2307
rect 1710 2307 1716 2308
rect 1676 2304 1707 2306
rect 1676 2303 1677 2304
rect 1671 2302 1677 2303
rect 1087 2298 1093 2299
rect 1705 2298 1707 2304
rect 1710 2303 1711 2307
rect 1715 2306 1716 2307
rect 1743 2307 1749 2308
rect 1743 2306 1744 2307
rect 1715 2304 1744 2306
rect 1715 2303 1716 2304
rect 1710 2302 1716 2303
rect 1743 2303 1744 2304
rect 1748 2303 1749 2307
rect 1743 2302 1749 2303
rect 1790 2307 1796 2308
rect 1790 2303 1791 2307
rect 1795 2306 1796 2307
rect 1823 2307 1829 2308
rect 1823 2306 1824 2307
rect 1795 2304 1824 2306
rect 1795 2303 1796 2304
rect 1790 2302 1796 2303
rect 1823 2303 1824 2304
rect 1828 2303 1829 2307
rect 1823 2302 1829 2303
rect 1870 2307 1876 2308
rect 1870 2303 1871 2307
rect 1875 2306 1876 2307
rect 1903 2307 1909 2308
rect 1903 2306 1904 2307
rect 1875 2304 1904 2306
rect 1875 2303 1876 2304
rect 1870 2302 1876 2303
rect 1903 2303 1904 2304
rect 1908 2303 1909 2307
rect 1903 2302 1909 2303
rect 1991 2307 1997 2308
rect 1991 2303 1992 2307
rect 1996 2306 1997 2307
rect 2074 2307 2080 2308
rect 2074 2306 2075 2307
rect 1996 2304 2075 2306
rect 1996 2303 1997 2304
rect 1991 2302 1997 2303
rect 2074 2303 2075 2304
rect 2079 2303 2080 2307
rect 2074 2302 2080 2303
rect 2087 2307 2093 2308
rect 2087 2303 2088 2307
rect 2092 2306 2093 2307
rect 2178 2307 2184 2308
rect 2178 2306 2179 2307
rect 2092 2304 2179 2306
rect 2092 2303 2093 2304
rect 2087 2302 2093 2303
rect 2178 2303 2179 2304
rect 2183 2303 2184 2307
rect 2178 2302 2184 2303
rect 2186 2307 2197 2308
rect 2186 2303 2187 2307
rect 2191 2303 2192 2307
rect 2196 2303 2197 2307
rect 2186 2302 2197 2303
rect 2295 2307 2301 2308
rect 2295 2303 2296 2307
rect 2300 2306 2301 2307
rect 2342 2307 2348 2308
rect 2342 2306 2343 2307
rect 2300 2304 2343 2306
rect 2300 2303 2301 2304
rect 2295 2302 2301 2303
rect 2342 2303 2343 2304
rect 2347 2303 2348 2307
rect 2342 2302 2348 2303
rect 2350 2307 2356 2308
rect 2350 2303 2351 2307
rect 2355 2306 2356 2307
rect 2383 2307 2389 2308
rect 2406 2307 2412 2308
rect 2383 2306 2384 2307
rect 2355 2304 2384 2306
rect 2355 2303 2356 2304
rect 2350 2302 2356 2303
rect 2383 2303 2384 2304
rect 2388 2303 2389 2307
rect 2383 2302 2389 2303
rect 1790 2299 1796 2300
rect 1790 2298 1791 2299
rect 1705 2296 1791 2298
rect 1278 2295 1284 2296
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 1238 2291 1244 2292
rect 1238 2287 1239 2291
rect 1243 2287 1244 2291
rect 1278 2291 1279 2295
rect 1283 2291 1284 2295
rect 1790 2295 1791 2296
rect 1795 2295 1796 2299
rect 1790 2294 1796 2295
rect 2406 2295 2412 2296
rect 1278 2290 1284 2291
rect 2406 2291 2407 2295
rect 2411 2291 2412 2295
rect 2406 2290 2412 2291
rect 1238 2286 1244 2287
rect 1326 2288 1332 2289
rect 270 2284 276 2285
rect 270 2280 271 2284
rect 275 2280 276 2284
rect 270 2279 276 2280
rect 326 2284 332 2285
rect 326 2280 327 2284
rect 331 2280 332 2284
rect 326 2279 332 2280
rect 398 2284 404 2285
rect 398 2280 399 2284
rect 403 2280 404 2284
rect 398 2279 404 2280
rect 470 2284 476 2285
rect 470 2280 471 2284
rect 475 2280 476 2284
rect 470 2279 476 2280
rect 550 2284 556 2285
rect 550 2280 551 2284
rect 555 2280 556 2284
rect 550 2279 556 2280
rect 630 2284 636 2285
rect 630 2280 631 2284
rect 635 2280 636 2284
rect 630 2279 636 2280
rect 710 2284 716 2285
rect 710 2280 711 2284
rect 715 2280 716 2284
rect 710 2279 716 2280
rect 782 2284 788 2285
rect 782 2280 783 2284
rect 787 2280 788 2284
rect 782 2279 788 2280
rect 854 2284 860 2285
rect 854 2280 855 2284
rect 859 2280 860 2284
rect 854 2279 860 2280
rect 918 2284 924 2285
rect 918 2280 919 2284
rect 923 2280 924 2284
rect 918 2279 924 2280
rect 990 2284 996 2285
rect 990 2280 991 2284
rect 995 2280 996 2284
rect 990 2279 996 2280
rect 1062 2284 1068 2285
rect 1062 2280 1063 2284
rect 1067 2280 1068 2284
rect 1326 2284 1327 2288
rect 1331 2284 1332 2288
rect 1326 2283 1332 2284
rect 1382 2288 1388 2289
rect 1382 2284 1383 2288
rect 1387 2284 1388 2288
rect 1382 2283 1388 2284
rect 1438 2288 1444 2289
rect 1438 2284 1439 2288
rect 1443 2284 1444 2288
rect 1438 2283 1444 2284
rect 1502 2288 1508 2289
rect 1502 2284 1503 2288
rect 1507 2284 1508 2288
rect 1502 2283 1508 2284
rect 1574 2288 1580 2289
rect 1574 2284 1575 2288
rect 1579 2284 1580 2288
rect 1574 2283 1580 2284
rect 1646 2288 1652 2289
rect 1646 2284 1647 2288
rect 1651 2284 1652 2288
rect 1646 2283 1652 2284
rect 1718 2288 1724 2289
rect 1718 2284 1719 2288
rect 1723 2284 1724 2288
rect 1718 2283 1724 2284
rect 1798 2288 1804 2289
rect 1798 2284 1799 2288
rect 1803 2284 1804 2288
rect 1798 2283 1804 2284
rect 1878 2288 1884 2289
rect 1878 2284 1879 2288
rect 1883 2284 1884 2288
rect 1878 2283 1884 2284
rect 1966 2288 1972 2289
rect 1966 2284 1967 2288
rect 1971 2284 1972 2288
rect 1966 2283 1972 2284
rect 2062 2288 2068 2289
rect 2062 2284 2063 2288
rect 2067 2284 2068 2288
rect 2062 2283 2068 2284
rect 2166 2288 2172 2289
rect 2166 2284 2167 2288
rect 2171 2284 2172 2288
rect 2166 2283 2172 2284
rect 2270 2288 2276 2289
rect 2270 2284 2271 2288
rect 2275 2284 2276 2288
rect 2270 2283 2276 2284
rect 2358 2288 2364 2289
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 1062 2279 1068 2280
rect 1334 2276 1340 2277
rect 1334 2272 1335 2276
rect 1339 2272 1340 2276
rect 1334 2271 1340 2272
rect 1406 2276 1412 2277
rect 1406 2272 1407 2276
rect 1411 2272 1412 2276
rect 1406 2271 1412 2272
rect 1486 2276 1492 2277
rect 1486 2272 1487 2276
rect 1491 2272 1492 2276
rect 1486 2271 1492 2272
rect 1558 2276 1564 2277
rect 1558 2272 1559 2276
rect 1563 2272 1564 2276
rect 1558 2271 1564 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1702 2276 1708 2277
rect 1702 2272 1703 2276
rect 1707 2272 1708 2276
rect 1702 2271 1708 2272
rect 1774 2276 1780 2277
rect 1774 2272 1775 2276
rect 1779 2272 1780 2276
rect 1774 2271 1780 2272
rect 1838 2276 1844 2277
rect 1838 2272 1839 2276
rect 1843 2272 1844 2276
rect 1838 2271 1844 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1990 2276 1996 2277
rect 1990 2272 1991 2276
rect 1995 2272 1996 2276
rect 1990 2271 1996 2272
rect 2078 2276 2084 2277
rect 2078 2272 2079 2276
rect 2083 2272 2084 2276
rect 2078 2271 2084 2272
rect 2174 2276 2180 2277
rect 2174 2272 2175 2276
rect 2179 2272 2180 2276
rect 2174 2271 2180 2272
rect 2278 2276 2284 2277
rect 2278 2272 2279 2276
rect 2283 2272 2284 2276
rect 2278 2271 2284 2272
rect 2358 2276 2364 2277
rect 2358 2272 2359 2276
rect 2363 2272 2364 2276
rect 2358 2271 2364 2272
rect 1278 2269 1284 2270
rect 1278 2265 1279 2269
rect 1283 2265 1284 2269
rect 142 2264 148 2265
rect 142 2260 143 2264
rect 147 2260 148 2264
rect 142 2259 148 2260
rect 182 2264 188 2265
rect 182 2260 183 2264
rect 187 2260 188 2264
rect 182 2259 188 2260
rect 222 2264 228 2265
rect 222 2260 223 2264
rect 227 2260 228 2264
rect 222 2259 228 2260
rect 278 2264 284 2265
rect 278 2260 279 2264
rect 283 2260 284 2264
rect 278 2259 284 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 406 2264 412 2265
rect 406 2260 407 2264
rect 411 2260 412 2264
rect 406 2259 412 2260
rect 478 2264 484 2265
rect 478 2260 479 2264
rect 483 2260 484 2264
rect 478 2259 484 2260
rect 558 2264 564 2265
rect 558 2260 559 2264
rect 563 2260 564 2264
rect 558 2259 564 2260
rect 646 2264 652 2265
rect 646 2260 647 2264
rect 651 2260 652 2264
rect 646 2259 652 2260
rect 726 2264 732 2265
rect 726 2260 727 2264
rect 731 2260 732 2264
rect 726 2259 732 2260
rect 806 2264 812 2265
rect 806 2260 807 2264
rect 811 2260 812 2264
rect 806 2259 812 2260
rect 886 2264 892 2265
rect 886 2260 887 2264
rect 891 2260 892 2264
rect 886 2259 892 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 1046 2264 1052 2265
rect 1046 2260 1047 2264
rect 1051 2260 1052 2264
rect 1046 2259 1052 2260
rect 1126 2264 1132 2265
rect 1278 2264 1284 2265
rect 2406 2269 2412 2270
rect 2406 2265 2407 2269
rect 2411 2265 2412 2269
rect 2406 2264 2412 2265
rect 1126 2260 1127 2264
rect 1131 2260 1132 2264
rect 1978 2263 1984 2264
rect 1978 2262 1979 2263
rect 1126 2259 1132 2260
rect 1864 2260 1979 2262
rect 110 2257 116 2258
rect 110 2253 111 2257
rect 115 2253 116 2257
rect 110 2252 116 2253
rect 1238 2257 1244 2258
rect 1238 2253 1239 2257
rect 1243 2253 1244 2257
rect 1864 2256 1866 2260
rect 1978 2259 1979 2260
rect 1983 2259 1984 2263
rect 1978 2258 1984 2259
rect 1354 2255 1365 2256
rect 1238 2252 1244 2253
rect 1278 2252 1284 2253
rect 1278 2248 1279 2252
rect 1283 2248 1284 2252
rect 1354 2251 1355 2255
rect 1359 2251 1360 2255
rect 1364 2251 1365 2255
rect 1354 2250 1365 2251
rect 1367 2255 1373 2256
rect 1367 2251 1368 2255
rect 1372 2254 1373 2255
rect 1431 2255 1437 2256
rect 1431 2254 1432 2255
rect 1372 2252 1432 2254
rect 1372 2251 1373 2252
rect 1367 2250 1373 2251
rect 1431 2251 1432 2252
rect 1436 2251 1437 2255
rect 1431 2250 1437 2251
rect 1439 2255 1445 2256
rect 1439 2251 1440 2255
rect 1444 2254 1445 2255
rect 1511 2255 1517 2256
rect 1511 2254 1512 2255
rect 1444 2252 1512 2254
rect 1444 2251 1445 2252
rect 1439 2250 1445 2251
rect 1511 2251 1512 2252
rect 1516 2251 1517 2255
rect 1511 2250 1517 2251
rect 1583 2255 1589 2256
rect 1583 2251 1584 2255
rect 1588 2254 1589 2255
rect 1614 2255 1620 2256
rect 1614 2254 1615 2255
rect 1588 2252 1615 2254
rect 1588 2251 1589 2252
rect 1583 2250 1589 2251
rect 1614 2251 1615 2252
rect 1619 2251 1620 2255
rect 1614 2250 1620 2251
rect 1622 2255 1628 2256
rect 1622 2251 1623 2255
rect 1627 2254 1628 2255
rect 1655 2255 1661 2256
rect 1655 2254 1656 2255
rect 1627 2252 1656 2254
rect 1627 2251 1628 2252
rect 1622 2250 1628 2251
rect 1655 2251 1656 2252
rect 1660 2251 1661 2255
rect 1655 2250 1661 2251
rect 1663 2255 1669 2256
rect 1663 2251 1664 2255
rect 1668 2254 1669 2255
rect 1727 2255 1733 2256
rect 1727 2254 1728 2255
rect 1668 2252 1728 2254
rect 1668 2251 1669 2252
rect 1663 2250 1669 2251
rect 1727 2251 1728 2252
rect 1732 2251 1733 2255
rect 1727 2250 1733 2251
rect 1735 2255 1741 2256
rect 1735 2251 1736 2255
rect 1740 2254 1741 2255
rect 1799 2255 1805 2256
rect 1799 2254 1800 2255
rect 1740 2252 1800 2254
rect 1740 2251 1741 2252
rect 1735 2250 1741 2251
rect 1799 2251 1800 2252
rect 1804 2251 1805 2255
rect 1799 2250 1805 2251
rect 1863 2255 1869 2256
rect 1863 2251 1864 2255
rect 1868 2251 1869 2255
rect 1863 2250 1869 2251
rect 1871 2255 1877 2256
rect 1871 2251 1872 2255
rect 1876 2254 1877 2255
rect 1935 2255 1941 2256
rect 1935 2254 1936 2255
rect 1876 2252 1936 2254
rect 1876 2251 1877 2252
rect 1871 2250 1877 2251
rect 1935 2251 1936 2252
rect 1940 2251 1941 2255
rect 1935 2250 1941 2251
rect 1943 2255 1949 2256
rect 1943 2251 1944 2255
rect 1948 2254 1949 2255
rect 2015 2255 2021 2256
rect 2015 2254 2016 2255
rect 1948 2252 2016 2254
rect 1948 2251 1949 2252
rect 1943 2250 1949 2251
rect 2015 2251 2016 2252
rect 2020 2251 2021 2255
rect 2015 2250 2021 2251
rect 2023 2255 2029 2256
rect 2023 2251 2024 2255
rect 2028 2254 2029 2255
rect 2103 2255 2109 2256
rect 2103 2254 2104 2255
rect 2028 2252 2104 2254
rect 2028 2251 2029 2252
rect 2023 2250 2029 2251
rect 2103 2251 2104 2252
rect 2108 2251 2109 2255
rect 2103 2250 2109 2251
rect 2111 2255 2117 2256
rect 2111 2251 2112 2255
rect 2116 2254 2117 2255
rect 2199 2255 2205 2256
rect 2199 2254 2200 2255
rect 2116 2252 2200 2254
rect 2116 2251 2117 2252
rect 2111 2250 2117 2251
rect 2199 2251 2200 2252
rect 2204 2251 2205 2255
rect 2199 2250 2205 2251
rect 2207 2255 2213 2256
rect 2207 2251 2208 2255
rect 2212 2254 2213 2255
rect 2303 2255 2309 2256
rect 2303 2254 2304 2255
rect 2212 2252 2304 2254
rect 2212 2251 2213 2252
rect 2207 2250 2213 2251
rect 2303 2251 2304 2252
rect 2308 2251 2309 2255
rect 2303 2250 2309 2251
rect 2382 2255 2389 2256
rect 2382 2251 2383 2255
rect 2388 2251 2389 2255
rect 2382 2250 2389 2251
rect 2406 2252 2412 2253
rect 1278 2247 1284 2248
rect 2406 2248 2407 2252
rect 2411 2248 2412 2252
rect 2406 2247 2412 2248
rect 167 2243 173 2244
rect 110 2240 116 2241
rect 110 2236 111 2240
rect 115 2236 116 2240
rect 167 2239 168 2243
rect 172 2242 173 2243
rect 198 2243 204 2244
rect 198 2242 199 2243
rect 172 2240 199 2242
rect 172 2239 173 2240
rect 167 2238 173 2239
rect 198 2239 199 2240
rect 203 2239 204 2243
rect 198 2238 204 2239
rect 207 2243 213 2244
rect 207 2239 208 2243
rect 212 2242 213 2243
rect 238 2243 244 2244
rect 238 2242 239 2243
rect 212 2240 239 2242
rect 212 2239 213 2240
rect 207 2238 213 2239
rect 238 2239 239 2240
rect 243 2239 244 2243
rect 238 2238 244 2239
rect 247 2243 253 2244
rect 247 2239 248 2243
rect 252 2242 253 2243
rect 294 2243 300 2244
rect 294 2242 295 2243
rect 252 2240 295 2242
rect 252 2239 253 2240
rect 247 2238 253 2239
rect 294 2239 295 2240
rect 299 2239 300 2243
rect 294 2238 300 2239
rect 303 2243 309 2244
rect 303 2239 304 2243
rect 308 2242 309 2243
rect 350 2243 356 2244
rect 350 2242 351 2243
rect 308 2240 351 2242
rect 308 2239 309 2240
rect 303 2238 309 2239
rect 350 2239 351 2240
rect 355 2239 356 2243
rect 350 2238 356 2239
rect 359 2243 365 2244
rect 359 2239 360 2243
rect 364 2242 365 2243
rect 378 2243 384 2244
rect 378 2242 379 2243
rect 364 2240 379 2242
rect 364 2239 365 2240
rect 359 2238 365 2239
rect 378 2239 379 2240
rect 383 2239 384 2243
rect 378 2238 384 2239
rect 386 2243 392 2244
rect 386 2239 387 2243
rect 391 2242 392 2243
rect 431 2243 437 2244
rect 431 2242 432 2243
rect 391 2240 432 2242
rect 391 2239 392 2240
rect 386 2238 392 2239
rect 431 2239 432 2240
rect 436 2239 437 2243
rect 431 2238 437 2239
rect 503 2243 509 2244
rect 503 2239 504 2243
rect 508 2242 509 2243
rect 542 2243 548 2244
rect 542 2242 543 2243
rect 508 2240 543 2242
rect 508 2239 509 2240
rect 503 2238 509 2239
rect 542 2239 543 2240
rect 547 2239 548 2243
rect 542 2238 548 2239
rect 550 2243 556 2244
rect 550 2239 551 2243
rect 555 2242 556 2243
rect 583 2243 589 2244
rect 583 2242 584 2243
rect 555 2240 584 2242
rect 555 2239 556 2240
rect 550 2238 556 2239
rect 583 2239 584 2240
rect 588 2239 589 2243
rect 583 2238 589 2239
rect 670 2243 677 2244
rect 670 2239 671 2243
rect 676 2239 677 2243
rect 670 2238 677 2239
rect 686 2243 692 2244
rect 686 2239 687 2243
rect 691 2242 692 2243
rect 751 2243 757 2244
rect 751 2242 752 2243
rect 691 2240 752 2242
rect 691 2239 692 2240
rect 686 2238 692 2239
rect 751 2239 752 2240
rect 756 2239 757 2243
rect 751 2238 757 2239
rect 759 2243 765 2244
rect 759 2239 760 2243
rect 764 2242 765 2243
rect 831 2243 837 2244
rect 831 2242 832 2243
rect 764 2240 832 2242
rect 764 2239 765 2240
rect 759 2238 765 2239
rect 831 2239 832 2240
rect 836 2239 837 2243
rect 831 2238 837 2239
rect 911 2243 917 2244
rect 911 2239 912 2243
rect 916 2239 917 2243
rect 911 2238 917 2239
rect 919 2243 925 2244
rect 919 2239 920 2243
rect 924 2242 925 2243
rect 991 2243 997 2244
rect 991 2242 992 2243
rect 924 2240 992 2242
rect 924 2239 925 2240
rect 919 2238 925 2239
rect 991 2239 992 2240
rect 996 2239 997 2243
rect 991 2238 997 2239
rect 1071 2243 1077 2244
rect 1071 2239 1072 2243
rect 1076 2242 1077 2243
rect 1134 2243 1140 2244
rect 1134 2242 1135 2243
rect 1076 2240 1135 2242
rect 1076 2239 1077 2240
rect 1071 2238 1077 2239
rect 1134 2239 1135 2240
rect 1139 2239 1140 2243
rect 1134 2238 1140 2239
rect 1142 2243 1148 2244
rect 1142 2239 1143 2243
rect 1147 2242 1148 2243
rect 1151 2243 1157 2244
rect 1151 2242 1152 2243
rect 1147 2240 1152 2242
rect 1147 2239 1148 2240
rect 1142 2238 1148 2239
rect 1151 2239 1152 2240
rect 1156 2239 1157 2243
rect 1151 2238 1157 2239
rect 1238 2240 1244 2241
rect 110 2235 116 2236
rect 912 2234 914 2238
rect 1238 2236 1239 2240
rect 1243 2236 1244 2240
rect 1070 2235 1076 2236
rect 1238 2235 1244 2236
rect 1070 2234 1071 2235
rect 912 2232 1071 2234
rect 1070 2231 1071 2232
rect 1075 2231 1076 2235
rect 1070 2230 1076 2231
rect 1334 2229 1340 2230
rect 1334 2225 1335 2229
rect 1339 2225 1340 2229
rect 1334 2224 1340 2225
rect 1406 2229 1412 2230
rect 1406 2225 1407 2229
rect 1411 2225 1412 2229
rect 1406 2224 1412 2225
rect 1486 2229 1492 2230
rect 1486 2225 1487 2229
rect 1491 2225 1492 2229
rect 1486 2224 1492 2225
rect 1558 2229 1564 2230
rect 1558 2225 1559 2229
rect 1563 2225 1564 2229
rect 1558 2224 1564 2225
rect 1630 2229 1636 2230
rect 1630 2225 1631 2229
rect 1635 2225 1636 2229
rect 1630 2224 1636 2225
rect 1702 2229 1708 2230
rect 1702 2225 1703 2229
rect 1707 2225 1708 2229
rect 1702 2224 1708 2225
rect 1774 2229 1780 2230
rect 1774 2225 1775 2229
rect 1779 2225 1780 2229
rect 1774 2224 1780 2225
rect 1838 2229 1844 2230
rect 1838 2225 1839 2229
rect 1843 2225 1844 2229
rect 1838 2224 1844 2225
rect 1910 2229 1916 2230
rect 1910 2225 1911 2229
rect 1915 2225 1916 2229
rect 1910 2224 1916 2225
rect 1990 2229 1996 2230
rect 1990 2225 1991 2229
rect 1995 2225 1996 2229
rect 1990 2224 1996 2225
rect 2078 2229 2084 2230
rect 2078 2225 2079 2229
rect 2083 2225 2084 2229
rect 2078 2224 2084 2225
rect 2174 2229 2180 2230
rect 2174 2225 2175 2229
rect 2179 2225 2180 2229
rect 2174 2224 2180 2225
rect 2278 2229 2284 2230
rect 2278 2225 2279 2229
rect 2283 2225 2284 2229
rect 2278 2224 2284 2225
rect 2358 2229 2364 2230
rect 2358 2225 2359 2229
rect 2363 2225 2364 2229
rect 2358 2224 2364 2225
rect 1359 2223 1365 2224
rect 1359 2219 1360 2223
rect 1364 2222 1365 2223
rect 1367 2223 1373 2224
rect 1367 2222 1368 2223
rect 1364 2220 1368 2222
rect 1364 2219 1365 2220
rect 1359 2218 1365 2219
rect 1367 2219 1368 2220
rect 1372 2219 1373 2223
rect 1367 2218 1373 2219
rect 1431 2223 1437 2224
rect 1431 2219 1432 2223
rect 1436 2222 1437 2223
rect 1439 2223 1445 2224
rect 1439 2222 1440 2223
rect 1436 2220 1440 2222
rect 1436 2219 1437 2220
rect 1431 2218 1437 2219
rect 1439 2219 1440 2220
rect 1444 2219 1445 2223
rect 1439 2218 1445 2219
rect 1511 2223 1517 2224
rect 1511 2219 1512 2223
rect 1516 2222 1517 2223
rect 1534 2223 1540 2224
rect 1534 2222 1535 2223
rect 1516 2220 1535 2222
rect 1516 2219 1517 2220
rect 1511 2218 1517 2219
rect 1534 2219 1535 2220
rect 1539 2219 1540 2223
rect 1534 2218 1540 2219
rect 1583 2223 1589 2224
rect 1583 2219 1584 2223
rect 1588 2222 1589 2223
rect 1622 2223 1628 2224
rect 1622 2222 1623 2223
rect 1588 2220 1623 2222
rect 1588 2219 1589 2220
rect 1583 2218 1589 2219
rect 1622 2219 1623 2220
rect 1627 2219 1628 2223
rect 1622 2218 1628 2219
rect 1655 2223 1661 2224
rect 1655 2219 1656 2223
rect 1660 2222 1661 2223
rect 1663 2223 1669 2224
rect 1663 2222 1664 2223
rect 1660 2220 1664 2222
rect 1660 2219 1661 2220
rect 1655 2218 1661 2219
rect 1663 2219 1664 2220
rect 1668 2219 1669 2223
rect 1663 2218 1669 2219
rect 1727 2223 1733 2224
rect 1727 2219 1728 2223
rect 1732 2222 1733 2223
rect 1735 2223 1741 2224
rect 1735 2222 1736 2223
rect 1732 2220 1736 2222
rect 1732 2219 1733 2220
rect 1727 2218 1733 2219
rect 1735 2219 1736 2220
rect 1740 2219 1741 2223
rect 1735 2218 1741 2219
rect 1790 2223 1796 2224
rect 1790 2219 1791 2223
rect 1795 2222 1796 2223
rect 1799 2223 1805 2224
rect 1799 2222 1800 2223
rect 1795 2220 1800 2222
rect 1795 2219 1796 2220
rect 1790 2218 1796 2219
rect 1799 2219 1800 2220
rect 1804 2219 1805 2223
rect 1799 2218 1805 2219
rect 1863 2223 1869 2224
rect 1863 2219 1864 2223
rect 1868 2222 1869 2223
rect 1871 2223 1877 2224
rect 1871 2222 1872 2223
rect 1868 2220 1872 2222
rect 1868 2219 1869 2220
rect 1863 2218 1869 2219
rect 1871 2219 1872 2220
rect 1876 2219 1877 2223
rect 1871 2218 1877 2219
rect 1935 2223 1941 2224
rect 1935 2219 1936 2223
rect 1940 2222 1941 2223
rect 1943 2223 1949 2224
rect 1943 2222 1944 2223
rect 1940 2220 1944 2222
rect 1940 2219 1941 2220
rect 1935 2218 1941 2219
rect 1943 2219 1944 2220
rect 1948 2219 1949 2223
rect 1943 2218 1949 2219
rect 2015 2223 2021 2224
rect 2015 2219 2016 2223
rect 2020 2222 2021 2223
rect 2023 2223 2029 2224
rect 2023 2222 2024 2223
rect 2020 2220 2024 2222
rect 2020 2219 2021 2220
rect 2015 2218 2021 2219
rect 2023 2219 2024 2220
rect 2028 2219 2029 2223
rect 2023 2218 2029 2219
rect 2103 2223 2109 2224
rect 2103 2219 2104 2223
rect 2108 2222 2109 2223
rect 2111 2223 2117 2224
rect 2111 2222 2112 2223
rect 2108 2220 2112 2222
rect 2108 2219 2109 2220
rect 2103 2218 2109 2219
rect 2111 2219 2112 2220
rect 2116 2219 2117 2223
rect 2111 2218 2117 2219
rect 2199 2223 2205 2224
rect 2199 2219 2200 2223
rect 2204 2222 2205 2223
rect 2207 2223 2213 2224
rect 2207 2222 2208 2223
rect 2204 2220 2208 2222
rect 2204 2219 2205 2220
rect 2199 2218 2205 2219
rect 2207 2219 2208 2220
rect 2212 2219 2213 2223
rect 2207 2218 2213 2219
rect 2303 2223 2309 2224
rect 2303 2219 2304 2223
rect 2308 2219 2309 2223
rect 2303 2218 2309 2219
rect 2342 2223 2348 2224
rect 2342 2219 2343 2223
rect 2347 2222 2348 2223
rect 2383 2223 2389 2224
rect 2383 2222 2384 2223
rect 2347 2220 2384 2222
rect 2347 2219 2348 2220
rect 2342 2218 2348 2219
rect 2383 2219 2384 2220
rect 2388 2219 2389 2223
rect 2383 2218 2389 2219
rect 142 2217 148 2218
rect 142 2213 143 2217
rect 147 2213 148 2217
rect 142 2212 148 2213
rect 182 2217 188 2218
rect 182 2213 183 2217
rect 187 2213 188 2217
rect 182 2212 188 2213
rect 222 2217 228 2218
rect 222 2213 223 2217
rect 227 2213 228 2217
rect 222 2212 228 2213
rect 278 2217 284 2218
rect 278 2213 279 2217
rect 283 2213 284 2217
rect 278 2212 284 2213
rect 334 2217 340 2218
rect 334 2213 335 2217
rect 339 2213 340 2217
rect 334 2212 340 2213
rect 406 2217 412 2218
rect 406 2213 407 2217
rect 411 2213 412 2217
rect 406 2212 412 2213
rect 478 2217 484 2218
rect 478 2213 479 2217
rect 483 2213 484 2217
rect 478 2212 484 2213
rect 558 2217 564 2218
rect 558 2213 559 2217
rect 563 2213 564 2217
rect 558 2212 564 2213
rect 646 2217 652 2218
rect 646 2213 647 2217
rect 651 2213 652 2217
rect 646 2212 652 2213
rect 726 2217 732 2218
rect 726 2213 727 2217
rect 731 2213 732 2217
rect 726 2212 732 2213
rect 806 2217 812 2218
rect 806 2213 807 2217
rect 811 2213 812 2217
rect 806 2212 812 2213
rect 886 2217 892 2218
rect 886 2213 887 2217
rect 891 2213 892 2217
rect 886 2212 892 2213
rect 966 2217 972 2218
rect 966 2213 967 2217
rect 971 2213 972 2217
rect 1046 2217 1052 2218
rect 1006 2215 1012 2216
rect 1006 2214 1007 2215
rect 966 2212 972 2213
rect 991 2213 1007 2214
rect 162 2211 173 2212
rect 162 2207 163 2211
rect 167 2207 168 2211
rect 172 2207 173 2211
rect 162 2206 173 2207
rect 198 2211 204 2212
rect 198 2207 199 2211
rect 203 2210 204 2211
rect 207 2211 213 2212
rect 207 2210 208 2211
rect 203 2208 208 2210
rect 203 2207 204 2208
rect 198 2206 204 2207
rect 207 2207 208 2208
rect 212 2207 213 2211
rect 207 2206 213 2207
rect 238 2211 244 2212
rect 238 2207 239 2211
rect 243 2210 244 2211
rect 247 2211 253 2212
rect 247 2210 248 2211
rect 243 2208 248 2210
rect 243 2207 244 2208
rect 238 2206 244 2207
rect 247 2207 248 2208
rect 252 2207 253 2211
rect 247 2206 253 2207
rect 294 2211 300 2212
rect 294 2207 295 2211
rect 299 2210 300 2211
rect 303 2211 309 2212
rect 303 2210 304 2211
rect 299 2208 304 2210
rect 299 2207 300 2208
rect 294 2206 300 2207
rect 303 2207 304 2208
rect 308 2207 309 2211
rect 303 2206 309 2207
rect 350 2211 356 2212
rect 350 2207 351 2211
rect 355 2210 356 2211
rect 359 2211 365 2212
rect 359 2210 360 2211
rect 355 2208 360 2210
rect 355 2207 356 2208
rect 350 2206 356 2207
rect 359 2207 360 2208
rect 364 2207 365 2211
rect 359 2206 365 2207
rect 378 2211 384 2212
rect 378 2207 379 2211
rect 383 2210 384 2211
rect 431 2211 437 2212
rect 431 2210 432 2211
rect 383 2208 432 2210
rect 383 2207 384 2208
rect 378 2206 384 2207
rect 431 2207 432 2208
rect 436 2207 437 2211
rect 431 2206 437 2207
rect 503 2211 509 2212
rect 503 2207 504 2211
rect 508 2210 509 2211
rect 550 2211 556 2212
rect 550 2210 551 2211
rect 508 2208 551 2210
rect 508 2207 509 2208
rect 503 2206 509 2207
rect 550 2207 551 2208
rect 555 2207 556 2211
rect 550 2206 556 2207
rect 578 2211 589 2212
rect 578 2207 579 2211
rect 583 2207 584 2211
rect 588 2207 589 2211
rect 578 2206 589 2207
rect 671 2211 677 2212
rect 671 2207 672 2211
rect 676 2210 677 2211
rect 686 2211 692 2212
rect 686 2210 687 2211
rect 676 2208 687 2210
rect 676 2207 677 2208
rect 671 2206 677 2207
rect 686 2207 687 2208
rect 691 2207 692 2211
rect 686 2206 692 2207
rect 751 2211 757 2212
rect 751 2207 752 2211
rect 756 2210 757 2211
rect 759 2211 765 2212
rect 759 2210 760 2211
rect 756 2208 760 2210
rect 756 2207 757 2208
rect 751 2206 757 2207
rect 759 2207 760 2208
rect 764 2207 765 2211
rect 759 2206 765 2207
rect 831 2211 837 2212
rect 831 2207 832 2211
rect 836 2210 837 2211
rect 854 2211 860 2212
rect 854 2210 855 2211
rect 836 2208 855 2210
rect 836 2207 837 2208
rect 831 2206 837 2207
rect 854 2207 855 2208
rect 859 2207 860 2211
rect 854 2206 860 2207
rect 911 2211 917 2212
rect 911 2207 912 2211
rect 916 2210 917 2211
rect 919 2211 925 2212
rect 919 2210 920 2211
rect 916 2208 920 2210
rect 916 2207 917 2208
rect 911 2206 917 2207
rect 919 2207 920 2208
rect 924 2207 925 2211
rect 991 2209 992 2213
rect 996 2212 1007 2213
rect 996 2209 997 2212
rect 1006 2211 1007 2212
rect 1011 2211 1012 2215
rect 1046 2213 1047 2217
rect 1051 2213 1052 2217
rect 1046 2212 1052 2213
rect 1126 2217 1132 2218
rect 1126 2213 1127 2217
rect 1131 2213 1132 2217
rect 1126 2212 1132 2213
rect 1858 2215 1864 2216
rect 1006 2210 1012 2211
rect 1070 2211 1077 2212
rect 991 2208 997 2209
rect 919 2206 925 2207
rect 1070 2207 1071 2211
rect 1076 2207 1077 2211
rect 1070 2206 1077 2207
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2210 1140 2211
rect 1151 2211 1157 2212
rect 1151 2210 1152 2211
rect 1139 2208 1152 2210
rect 1139 2207 1140 2208
rect 1134 2206 1140 2207
rect 1151 2207 1152 2208
rect 1156 2207 1157 2211
rect 1858 2211 1859 2215
rect 1863 2214 1864 2215
rect 2305 2214 2307 2218
rect 1863 2212 2307 2214
rect 1863 2211 1864 2212
rect 1858 2210 1864 2211
rect 1151 2206 1157 2207
rect 551 2195 557 2196
rect 159 2191 165 2192
rect 134 2187 140 2188
rect 134 2183 135 2187
rect 139 2183 140 2187
rect 159 2187 160 2191
rect 164 2190 165 2191
rect 198 2191 204 2192
rect 198 2190 199 2191
rect 164 2188 199 2190
rect 164 2187 165 2188
rect 159 2186 165 2187
rect 198 2187 199 2188
rect 203 2187 204 2191
rect 231 2191 237 2192
rect 198 2186 204 2187
rect 206 2187 212 2188
rect 134 2182 140 2183
rect 206 2183 207 2187
rect 211 2183 212 2187
rect 231 2187 232 2191
rect 236 2190 237 2191
rect 263 2191 269 2192
rect 263 2190 264 2191
rect 236 2188 264 2190
rect 236 2187 237 2188
rect 231 2186 237 2187
rect 263 2187 264 2188
rect 268 2187 269 2191
rect 303 2191 309 2192
rect 263 2186 269 2187
rect 278 2187 284 2188
rect 206 2182 212 2183
rect 278 2183 279 2187
rect 283 2183 284 2187
rect 303 2187 304 2191
rect 308 2190 309 2191
rect 350 2191 356 2192
rect 350 2190 351 2191
rect 308 2188 351 2190
rect 308 2187 309 2188
rect 303 2186 309 2187
rect 350 2187 351 2188
rect 355 2187 356 2191
rect 383 2191 392 2192
rect 350 2186 356 2187
rect 358 2187 364 2188
rect 278 2182 284 2183
rect 358 2183 359 2187
rect 363 2183 364 2187
rect 383 2187 384 2191
rect 391 2187 392 2191
rect 450 2191 456 2192
rect 383 2186 392 2187
rect 438 2187 444 2188
rect 358 2182 364 2183
rect 438 2183 439 2187
rect 443 2183 444 2187
rect 450 2187 451 2191
rect 455 2190 456 2191
rect 463 2191 469 2192
rect 463 2190 464 2191
rect 455 2188 464 2190
rect 455 2187 456 2188
rect 450 2186 456 2187
rect 463 2187 464 2188
rect 468 2187 469 2191
rect 542 2191 549 2192
rect 463 2186 469 2187
rect 518 2187 524 2188
rect 438 2182 444 2183
rect 518 2183 519 2187
rect 523 2183 524 2187
rect 542 2187 543 2191
rect 548 2187 549 2191
rect 551 2191 552 2195
rect 556 2194 557 2195
rect 1399 2195 1405 2196
rect 556 2192 610 2194
rect 556 2191 557 2192
rect 551 2190 557 2191
rect 608 2190 610 2192
rect 623 2191 629 2192
rect 623 2190 624 2191
rect 608 2188 624 2190
rect 542 2186 549 2187
rect 598 2187 604 2188
rect 518 2182 524 2183
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 623 2187 624 2188
rect 628 2187 629 2191
rect 703 2191 709 2192
rect 623 2186 629 2187
rect 678 2187 684 2188
rect 598 2182 604 2183
rect 678 2183 679 2187
rect 683 2183 684 2187
rect 703 2187 704 2191
rect 708 2190 709 2191
rect 746 2191 752 2192
rect 746 2190 747 2191
rect 708 2188 747 2190
rect 708 2187 709 2188
rect 703 2186 709 2187
rect 746 2187 747 2188
rect 751 2187 752 2191
rect 770 2191 776 2192
rect 746 2186 752 2187
rect 758 2187 764 2188
rect 678 2182 684 2183
rect 758 2183 759 2187
rect 763 2183 764 2187
rect 770 2187 771 2191
rect 775 2190 776 2191
rect 783 2191 789 2192
rect 783 2190 784 2191
rect 775 2188 784 2190
rect 775 2187 776 2188
rect 770 2186 776 2187
rect 783 2187 784 2188
rect 788 2187 789 2191
rect 842 2191 848 2192
rect 783 2186 789 2187
rect 830 2187 836 2188
rect 758 2182 764 2183
rect 830 2183 831 2187
rect 835 2183 836 2187
rect 842 2187 843 2191
rect 847 2190 848 2191
rect 855 2191 861 2192
rect 855 2190 856 2191
rect 847 2188 856 2190
rect 847 2187 848 2188
rect 842 2186 848 2187
rect 855 2187 856 2188
rect 860 2187 861 2191
rect 927 2191 933 2192
rect 855 2186 861 2187
rect 902 2187 908 2188
rect 830 2182 836 2183
rect 902 2183 903 2187
rect 907 2183 908 2187
rect 927 2187 928 2191
rect 932 2190 933 2191
rect 966 2191 972 2192
rect 966 2190 967 2191
rect 932 2188 967 2190
rect 932 2187 933 2188
rect 927 2186 933 2187
rect 966 2187 967 2188
rect 971 2187 972 2191
rect 999 2191 1005 2192
rect 966 2186 972 2187
rect 974 2187 980 2188
rect 902 2182 908 2183
rect 974 2183 975 2187
rect 979 2183 980 2187
rect 999 2187 1000 2191
rect 1004 2190 1005 2191
rect 1038 2191 1044 2192
rect 1038 2190 1039 2191
rect 1004 2188 1039 2190
rect 1004 2187 1005 2188
rect 999 2186 1005 2187
rect 1038 2187 1039 2188
rect 1043 2187 1044 2191
rect 1071 2191 1077 2192
rect 1038 2186 1044 2187
rect 1046 2187 1052 2188
rect 974 2182 980 2183
rect 1046 2183 1047 2187
rect 1051 2183 1052 2187
rect 1071 2187 1072 2191
rect 1076 2190 1077 2191
rect 1110 2191 1116 2192
rect 1110 2190 1111 2191
rect 1076 2188 1111 2190
rect 1076 2187 1077 2188
rect 1071 2186 1077 2187
rect 1110 2187 1111 2188
rect 1115 2187 1116 2191
rect 1142 2191 1149 2192
rect 1110 2186 1116 2187
rect 1118 2187 1124 2188
rect 1046 2182 1052 2183
rect 1118 2183 1119 2187
rect 1123 2183 1124 2187
rect 1142 2187 1143 2191
rect 1148 2187 1149 2191
rect 1142 2186 1149 2187
rect 1374 2191 1380 2192
rect 1374 2187 1375 2191
rect 1379 2187 1380 2191
rect 1399 2191 1400 2195
rect 1404 2194 1405 2195
rect 1422 2195 1428 2196
rect 1422 2194 1423 2195
rect 1404 2192 1423 2194
rect 1404 2191 1405 2192
rect 1399 2190 1405 2191
rect 1422 2191 1423 2192
rect 1427 2191 1428 2195
rect 1450 2195 1456 2196
rect 1422 2190 1428 2191
rect 1438 2191 1444 2192
rect 1374 2186 1380 2187
rect 1438 2187 1439 2191
rect 1443 2187 1444 2191
rect 1450 2191 1451 2195
rect 1455 2194 1456 2195
rect 1463 2195 1469 2196
rect 1463 2194 1464 2195
rect 1455 2192 1464 2194
rect 1455 2191 1456 2192
rect 1450 2190 1456 2191
rect 1463 2191 1464 2192
rect 1468 2191 1469 2195
rect 1522 2195 1528 2196
rect 1463 2190 1469 2191
rect 1510 2191 1516 2192
rect 1438 2186 1444 2187
rect 1510 2187 1511 2191
rect 1515 2187 1516 2191
rect 1522 2191 1523 2195
rect 1527 2194 1528 2195
rect 1535 2195 1541 2196
rect 1535 2194 1536 2195
rect 1527 2192 1536 2194
rect 1527 2191 1528 2192
rect 1522 2190 1528 2191
rect 1535 2191 1536 2192
rect 1540 2191 1541 2195
rect 1614 2195 1621 2196
rect 1535 2190 1541 2191
rect 1590 2191 1596 2192
rect 1510 2186 1516 2187
rect 1590 2187 1591 2191
rect 1595 2187 1596 2191
rect 1614 2191 1615 2195
rect 1620 2191 1621 2195
rect 1682 2195 1688 2196
rect 1614 2190 1621 2191
rect 1670 2191 1676 2192
rect 1590 2186 1596 2187
rect 1670 2187 1671 2191
rect 1675 2187 1676 2191
rect 1682 2191 1683 2195
rect 1687 2194 1688 2195
rect 1695 2195 1701 2196
rect 1695 2194 1696 2195
rect 1687 2192 1696 2194
rect 1687 2191 1688 2192
rect 1682 2190 1688 2191
rect 1695 2191 1696 2192
rect 1700 2191 1701 2195
rect 1762 2195 1768 2196
rect 1695 2190 1701 2191
rect 1750 2191 1756 2192
rect 1670 2186 1676 2187
rect 1750 2187 1751 2191
rect 1755 2187 1756 2191
rect 1762 2191 1763 2195
rect 1767 2194 1768 2195
rect 1775 2195 1781 2196
rect 1775 2194 1776 2195
rect 1767 2192 1776 2194
rect 1767 2191 1768 2192
rect 1762 2190 1768 2191
rect 1775 2191 1776 2192
rect 1780 2191 1781 2195
rect 1855 2195 1861 2196
rect 1775 2190 1781 2191
rect 1830 2191 1836 2192
rect 1750 2186 1756 2187
rect 1830 2187 1831 2191
rect 1835 2187 1836 2191
rect 1855 2191 1856 2195
rect 1860 2194 1861 2195
rect 1894 2195 1900 2196
rect 1894 2194 1895 2195
rect 1860 2192 1895 2194
rect 1860 2191 1861 2192
rect 1855 2190 1861 2191
rect 1894 2191 1895 2192
rect 1899 2191 1900 2195
rect 1927 2195 1933 2196
rect 1894 2190 1900 2191
rect 1902 2191 1908 2192
rect 1830 2186 1836 2187
rect 1902 2187 1903 2191
rect 1907 2187 1908 2191
rect 1927 2191 1928 2195
rect 1932 2194 1933 2195
rect 1958 2195 1964 2196
rect 1958 2194 1959 2195
rect 1932 2192 1959 2194
rect 1932 2191 1933 2192
rect 1927 2190 1933 2191
rect 1958 2191 1959 2192
rect 1963 2191 1964 2195
rect 1991 2195 1997 2196
rect 1958 2190 1964 2191
rect 1966 2191 1972 2192
rect 1902 2186 1908 2187
rect 1966 2187 1967 2191
rect 1971 2187 1972 2191
rect 1991 2191 1992 2195
rect 1996 2194 1997 2195
rect 2022 2195 2028 2196
rect 2022 2194 2023 2195
rect 1996 2192 2023 2194
rect 1996 2191 1997 2192
rect 1991 2190 1997 2191
rect 2022 2191 2023 2192
rect 2027 2191 2028 2195
rect 2055 2195 2061 2196
rect 2022 2190 2028 2191
rect 2030 2191 2036 2192
rect 1966 2186 1972 2187
rect 2030 2187 2031 2191
rect 2035 2187 2036 2191
rect 2055 2191 2056 2195
rect 2060 2194 2061 2195
rect 2086 2195 2092 2196
rect 2086 2194 2087 2195
rect 2060 2192 2087 2194
rect 2060 2191 2061 2192
rect 2055 2190 2061 2191
rect 2086 2191 2087 2192
rect 2091 2191 2092 2195
rect 2119 2195 2125 2196
rect 2086 2190 2092 2191
rect 2094 2191 2100 2192
rect 2030 2186 2036 2187
rect 2094 2187 2095 2191
rect 2099 2187 2100 2191
rect 2119 2191 2120 2195
rect 2124 2194 2125 2195
rect 2158 2195 2164 2196
rect 2158 2194 2159 2195
rect 2124 2192 2159 2194
rect 2124 2191 2125 2192
rect 2119 2190 2125 2191
rect 2158 2191 2159 2192
rect 2163 2191 2164 2195
rect 2191 2195 2197 2196
rect 2158 2190 2164 2191
rect 2166 2191 2172 2192
rect 2094 2186 2100 2187
rect 2166 2187 2167 2191
rect 2171 2187 2172 2191
rect 2191 2191 2192 2195
rect 2196 2194 2197 2195
rect 2230 2195 2236 2196
rect 2230 2194 2231 2195
rect 2196 2192 2231 2194
rect 2196 2191 2197 2192
rect 2191 2190 2197 2191
rect 2230 2191 2231 2192
rect 2235 2191 2236 2195
rect 2250 2195 2256 2196
rect 2230 2190 2236 2191
rect 2238 2191 2244 2192
rect 2166 2186 2172 2187
rect 2238 2187 2239 2191
rect 2243 2187 2244 2191
rect 2250 2191 2251 2195
rect 2255 2194 2256 2195
rect 2263 2195 2269 2196
rect 2263 2194 2264 2195
rect 2255 2192 2264 2194
rect 2255 2191 2256 2192
rect 2250 2190 2256 2191
rect 2263 2191 2264 2192
rect 2268 2191 2269 2195
rect 2335 2195 2341 2196
rect 2263 2190 2269 2191
rect 2310 2191 2316 2192
rect 2238 2186 2244 2187
rect 2310 2187 2311 2191
rect 2315 2187 2316 2191
rect 2335 2191 2336 2195
rect 2340 2194 2341 2195
rect 2350 2195 2356 2196
rect 2350 2194 2351 2195
rect 2340 2192 2351 2194
rect 2340 2191 2341 2192
rect 2335 2190 2341 2191
rect 2350 2191 2351 2192
rect 2355 2191 2356 2195
rect 2382 2195 2389 2196
rect 2350 2190 2356 2191
rect 2358 2191 2364 2192
rect 2310 2186 2316 2187
rect 2358 2187 2359 2191
rect 2363 2187 2364 2191
rect 2382 2191 2383 2195
rect 2388 2191 2389 2195
rect 2382 2190 2389 2191
rect 2358 2186 2364 2187
rect 1118 2182 1124 2183
rect 1278 2168 1284 2169
rect 450 2167 456 2168
rect 450 2166 451 2167
rect 110 2164 116 2165
rect 110 2160 111 2164
rect 115 2160 116 2164
rect 344 2164 451 2166
rect 110 2159 116 2160
rect 159 2159 168 2160
rect 159 2155 160 2159
rect 167 2155 168 2159
rect 159 2154 168 2155
rect 198 2159 204 2160
rect 198 2155 199 2159
rect 203 2158 204 2159
rect 231 2159 237 2160
rect 231 2158 232 2159
rect 203 2156 232 2158
rect 203 2155 204 2156
rect 198 2154 204 2155
rect 231 2155 232 2156
rect 236 2155 237 2159
rect 231 2154 237 2155
rect 303 2159 309 2160
rect 303 2155 304 2159
rect 308 2158 309 2159
rect 344 2158 346 2164
rect 450 2163 451 2164
rect 455 2163 456 2167
rect 450 2162 456 2163
rect 1238 2164 1244 2165
rect 1238 2160 1239 2164
rect 1243 2160 1244 2164
rect 1278 2164 1279 2168
rect 1283 2164 1284 2168
rect 2406 2168 2412 2169
rect 2406 2164 2407 2168
rect 2411 2164 2412 2168
rect 1278 2163 1284 2164
rect 1399 2163 1405 2164
rect 308 2156 346 2158
rect 350 2159 356 2160
rect 308 2155 309 2156
rect 303 2154 309 2155
rect 350 2155 351 2159
rect 355 2158 356 2159
rect 383 2159 389 2160
rect 383 2158 384 2159
rect 355 2156 384 2158
rect 355 2155 356 2156
rect 350 2154 356 2155
rect 383 2155 384 2156
rect 388 2155 389 2159
rect 383 2154 389 2155
rect 450 2159 456 2160
rect 450 2155 451 2159
rect 455 2158 456 2159
rect 463 2159 469 2160
rect 463 2158 464 2159
rect 455 2156 464 2158
rect 455 2155 456 2156
rect 450 2154 456 2155
rect 463 2155 464 2156
rect 468 2155 469 2159
rect 463 2154 469 2155
rect 543 2159 549 2160
rect 543 2155 544 2159
rect 548 2158 549 2159
rect 551 2159 557 2160
rect 551 2158 552 2159
rect 548 2156 552 2158
rect 548 2155 549 2156
rect 543 2154 549 2155
rect 551 2155 552 2156
rect 556 2155 557 2159
rect 551 2154 557 2155
rect 583 2159 589 2160
rect 583 2155 584 2159
rect 588 2158 589 2159
rect 623 2159 629 2160
rect 623 2158 624 2159
rect 588 2156 624 2158
rect 588 2155 589 2156
rect 583 2154 589 2155
rect 623 2155 624 2156
rect 628 2155 629 2159
rect 623 2154 629 2155
rect 703 2159 709 2160
rect 703 2155 704 2159
rect 708 2158 709 2159
rect 770 2159 776 2160
rect 770 2158 771 2159
rect 708 2156 771 2158
rect 708 2155 709 2156
rect 703 2154 709 2155
rect 770 2155 771 2156
rect 775 2155 776 2159
rect 770 2154 776 2155
rect 783 2159 789 2160
rect 783 2155 784 2159
rect 788 2158 789 2159
rect 842 2159 848 2160
rect 842 2158 843 2159
rect 788 2156 843 2158
rect 788 2155 789 2156
rect 783 2154 789 2155
rect 842 2155 843 2156
rect 847 2155 848 2159
rect 842 2154 848 2155
rect 854 2159 861 2160
rect 854 2155 855 2159
rect 860 2155 861 2159
rect 854 2154 861 2155
rect 927 2159 933 2160
rect 927 2155 928 2159
rect 932 2158 933 2159
rect 966 2159 972 2160
rect 932 2156 962 2158
rect 932 2155 933 2156
rect 927 2154 933 2155
rect 960 2150 962 2156
rect 966 2155 967 2159
rect 971 2158 972 2159
rect 999 2159 1005 2160
rect 999 2158 1000 2159
rect 971 2156 1000 2158
rect 971 2155 972 2156
rect 966 2154 972 2155
rect 999 2155 1000 2156
rect 1004 2155 1005 2159
rect 999 2154 1005 2155
rect 1038 2159 1044 2160
rect 1038 2155 1039 2159
rect 1043 2158 1044 2159
rect 1071 2159 1077 2160
rect 1071 2158 1072 2159
rect 1043 2156 1072 2158
rect 1043 2155 1044 2156
rect 1038 2154 1044 2155
rect 1071 2155 1072 2156
rect 1076 2155 1077 2159
rect 1071 2154 1077 2155
rect 1110 2159 1116 2160
rect 1110 2155 1111 2159
rect 1115 2158 1116 2159
rect 1143 2159 1149 2160
rect 1238 2159 1244 2160
rect 1399 2159 1400 2163
rect 1404 2162 1405 2163
rect 1450 2163 1456 2164
rect 1450 2162 1451 2163
rect 1404 2160 1451 2162
rect 1404 2159 1405 2160
rect 1143 2158 1144 2159
rect 1115 2156 1144 2158
rect 1115 2155 1116 2156
rect 1110 2154 1116 2155
rect 1143 2155 1144 2156
rect 1148 2155 1149 2159
rect 1399 2158 1405 2159
rect 1450 2159 1451 2160
rect 1455 2159 1456 2163
rect 1450 2158 1456 2159
rect 1463 2163 1469 2164
rect 1463 2159 1464 2163
rect 1468 2162 1469 2163
rect 1522 2163 1528 2164
rect 1522 2162 1523 2163
rect 1468 2160 1523 2162
rect 1468 2159 1469 2160
rect 1463 2158 1469 2159
rect 1522 2159 1523 2160
rect 1527 2159 1528 2163
rect 1522 2158 1528 2159
rect 1534 2163 1541 2164
rect 1534 2159 1535 2163
rect 1540 2159 1541 2163
rect 1534 2158 1541 2159
rect 1615 2163 1621 2164
rect 1615 2159 1616 2163
rect 1620 2162 1621 2163
rect 1682 2163 1688 2164
rect 1682 2162 1683 2163
rect 1620 2160 1683 2162
rect 1620 2159 1621 2160
rect 1615 2158 1621 2159
rect 1682 2159 1683 2160
rect 1687 2159 1688 2163
rect 1682 2158 1688 2159
rect 1695 2163 1701 2164
rect 1695 2159 1696 2163
rect 1700 2162 1701 2163
rect 1762 2163 1768 2164
rect 1762 2162 1763 2163
rect 1700 2160 1763 2162
rect 1700 2159 1701 2160
rect 1695 2158 1701 2159
rect 1762 2159 1763 2160
rect 1767 2159 1768 2163
rect 1762 2158 1768 2159
rect 1775 2163 1781 2164
rect 1775 2159 1776 2163
rect 1780 2162 1781 2163
rect 1846 2163 1852 2164
rect 1846 2162 1847 2163
rect 1780 2160 1847 2162
rect 1780 2159 1781 2160
rect 1775 2158 1781 2159
rect 1846 2159 1847 2160
rect 1851 2159 1852 2163
rect 1846 2158 1852 2159
rect 1855 2163 1864 2164
rect 1855 2159 1856 2163
rect 1863 2159 1864 2163
rect 1855 2158 1864 2159
rect 1894 2163 1900 2164
rect 1894 2159 1895 2163
rect 1899 2162 1900 2163
rect 1927 2163 1933 2164
rect 1927 2162 1928 2163
rect 1899 2160 1928 2162
rect 1899 2159 1900 2160
rect 1894 2158 1900 2159
rect 1927 2159 1928 2160
rect 1932 2159 1933 2163
rect 1927 2158 1933 2159
rect 1958 2163 1964 2164
rect 1958 2159 1959 2163
rect 1963 2162 1964 2163
rect 1991 2163 1997 2164
rect 1991 2162 1992 2163
rect 1963 2160 1992 2162
rect 1963 2159 1964 2160
rect 1958 2158 1964 2159
rect 1991 2159 1992 2160
rect 1996 2159 1997 2163
rect 1991 2158 1997 2159
rect 2022 2163 2028 2164
rect 2022 2159 2023 2163
rect 2027 2162 2028 2163
rect 2055 2163 2061 2164
rect 2055 2162 2056 2163
rect 2027 2160 2056 2162
rect 2027 2159 2028 2160
rect 2022 2158 2028 2159
rect 2055 2159 2056 2160
rect 2060 2159 2061 2163
rect 2055 2158 2061 2159
rect 2086 2163 2092 2164
rect 2086 2159 2087 2163
rect 2091 2162 2092 2163
rect 2119 2163 2125 2164
rect 2119 2162 2120 2163
rect 2091 2160 2120 2162
rect 2091 2159 2092 2160
rect 2086 2158 2092 2159
rect 2119 2159 2120 2160
rect 2124 2159 2125 2163
rect 2119 2158 2125 2159
rect 2158 2163 2164 2164
rect 2158 2159 2159 2163
rect 2163 2162 2164 2163
rect 2191 2163 2197 2164
rect 2191 2162 2192 2163
rect 2163 2160 2192 2162
rect 2163 2159 2164 2160
rect 2158 2158 2164 2159
rect 2191 2159 2192 2160
rect 2196 2159 2197 2163
rect 2191 2158 2197 2159
rect 2230 2163 2236 2164
rect 2230 2159 2231 2163
rect 2235 2162 2236 2163
rect 2263 2163 2269 2164
rect 2263 2162 2264 2163
rect 2235 2160 2264 2162
rect 2235 2159 2236 2160
rect 2230 2158 2236 2159
rect 2263 2159 2264 2160
rect 2268 2159 2269 2163
rect 2263 2158 2269 2159
rect 2335 2163 2344 2164
rect 2335 2159 2336 2163
rect 2343 2159 2344 2163
rect 2335 2158 2344 2159
rect 2350 2163 2356 2164
rect 2350 2159 2351 2163
rect 2355 2162 2356 2163
rect 2383 2163 2389 2164
rect 2406 2163 2412 2164
rect 2383 2162 2384 2163
rect 2355 2160 2384 2162
rect 2355 2159 2356 2160
rect 2350 2158 2356 2159
rect 2383 2159 2384 2160
rect 2388 2159 2389 2163
rect 2383 2158 2389 2159
rect 1143 2154 1149 2155
rect 1070 2151 1076 2152
rect 1070 2150 1071 2151
rect 960 2148 1071 2150
rect 110 2147 116 2148
rect 110 2143 111 2147
rect 115 2143 116 2147
rect 1070 2147 1071 2148
rect 1075 2147 1076 2151
rect 1278 2151 1284 2152
rect 1070 2146 1076 2147
rect 1238 2147 1244 2148
rect 110 2142 116 2143
rect 1238 2143 1239 2147
rect 1243 2143 1244 2147
rect 1278 2147 1279 2151
rect 1283 2147 1284 2151
rect 1278 2146 1284 2147
rect 2406 2151 2412 2152
rect 2406 2147 2407 2151
rect 2411 2147 2412 2151
rect 2406 2146 2412 2147
rect 1238 2142 1244 2143
rect 1374 2144 1380 2145
rect 134 2140 140 2141
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 206 2140 212 2141
rect 206 2136 207 2140
rect 211 2136 212 2140
rect 206 2135 212 2136
rect 278 2140 284 2141
rect 278 2136 279 2140
rect 283 2136 284 2140
rect 278 2135 284 2136
rect 358 2140 364 2141
rect 358 2136 359 2140
rect 363 2136 364 2140
rect 358 2135 364 2136
rect 438 2140 444 2141
rect 438 2136 439 2140
rect 443 2136 444 2140
rect 438 2135 444 2136
rect 518 2140 524 2141
rect 518 2136 519 2140
rect 523 2136 524 2140
rect 518 2135 524 2136
rect 598 2140 604 2141
rect 598 2136 599 2140
rect 603 2136 604 2140
rect 598 2135 604 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 758 2140 764 2141
rect 758 2136 759 2140
rect 763 2136 764 2140
rect 758 2135 764 2136
rect 830 2140 836 2141
rect 830 2136 831 2140
rect 835 2136 836 2140
rect 830 2135 836 2136
rect 902 2140 908 2141
rect 902 2136 903 2140
rect 907 2136 908 2140
rect 902 2135 908 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1046 2140 1052 2141
rect 1046 2136 1047 2140
rect 1051 2136 1052 2140
rect 1046 2135 1052 2136
rect 1118 2140 1124 2141
rect 1118 2136 1119 2140
rect 1123 2136 1124 2140
rect 1374 2140 1375 2144
rect 1379 2140 1380 2144
rect 1374 2139 1380 2140
rect 1438 2144 1444 2145
rect 1438 2140 1439 2144
rect 1443 2140 1444 2144
rect 1438 2139 1444 2140
rect 1510 2144 1516 2145
rect 1510 2140 1511 2144
rect 1515 2140 1516 2144
rect 1510 2139 1516 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1670 2144 1676 2145
rect 1670 2140 1671 2144
rect 1675 2140 1676 2144
rect 1670 2139 1676 2140
rect 1750 2144 1756 2145
rect 1750 2140 1751 2144
rect 1755 2140 1756 2144
rect 1750 2139 1756 2140
rect 1830 2144 1836 2145
rect 1830 2140 1831 2144
rect 1835 2140 1836 2144
rect 1830 2139 1836 2140
rect 1902 2144 1908 2145
rect 1902 2140 1903 2144
rect 1907 2140 1908 2144
rect 1902 2139 1908 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2030 2144 2036 2145
rect 2030 2140 2031 2144
rect 2035 2140 2036 2144
rect 2030 2139 2036 2140
rect 2094 2144 2100 2145
rect 2094 2140 2095 2144
rect 2099 2140 2100 2144
rect 2094 2139 2100 2140
rect 2166 2144 2172 2145
rect 2166 2140 2167 2144
rect 2171 2140 2172 2144
rect 2166 2139 2172 2140
rect 2238 2144 2244 2145
rect 2238 2140 2239 2144
rect 2243 2140 2244 2144
rect 2238 2139 2244 2140
rect 2310 2144 2316 2145
rect 2310 2140 2311 2144
rect 2315 2140 2316 2144
rect 2310 2139 2316 2140
rect 2358 2144 2364 2145
rect 2358 2140 2359 2144
rect 2363 2140 2364 2144
rect 2358 2139 2364 2140
rect 1118 2135 1124 2136
rect 1398 2132 1404 2133
rect 1398 2128 1399 2132
rect 1403 2128 1404 2132
rect 1398 2127 1404 2128
rect 1438 2132 1444 2133
rect 1438 2128 1439 2132
rect 1443 2128 1444 2132
rect 1438 2127 1444 2128
rect 1494 2132 1500 2133
rect 1494 2128 1495 2132
rect 1499 2128 1500 2132
rect 1494 2127 1500 2128
rect 1566 2132 1572 2133
rect 1566 2128 1567 2132
rect 1571 2128 1572 2132
rect 1566 2127 1572 2128
rect 1646 2132 1652 2133
rect 1646 2128 1647 2132
rect 1651 2128 1652 2132
rect 1646 2127 1652 2128
rect 1734 2132 1740 2133
rect 1734 2128 1735 2132
rect 1739 2128 1740 2132
rect 1734 2127 1740 2128
rect 1822 2132 1828 2133
rect 1822 2128 1823 2132
rect 1827 2128 1828 2132
rect 1822 2127 1828 2128
rect 1910 2132 1916 2133
rect 1910 2128 1911 2132
rect 1915 2128 1916 2132
rect 1910 2127 1916 2128
rect 1998 2132 2004 2133
rect 1998 2128 1999 2132
rect 2003 2128 2004 2132
rect 1998 2127 2004 2128
rect 2086 2132 2092 2133
rect 2086 2128 2087 2132
rect 2091 2128 2092 2132
rect 2086 2127 2092 2128
rect 2174 2132 2180 2133
rect 2174 2128 2175 2132
rect 2179 2128 2180 2132
rect 2174 2127 2180 2128
rect 2270 2132 2276 2133
rect 2270 2128 2271 2132
rect 2275 2128 2276 2132
rect 2270 2127 2276 2128
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 1278 2125 1284 2126
rect 1278 2121 1279 2125
rect 1283 2121 1284 2125
rect 134 2120 140 2121
rect 134 2116 135 2120
rect 139 2116 140 2120
rect 134 2115 140 2116
rect 190 2120 196 2121
rect 190 2116 191 2120
rect 195 2116 196 2120
rect 190 2115 196 2116
rect 270 2120 276 2121
rect 270 2116 271 2120
rect 275 2116 276 2120
rect 270 2115 276 2116
rect 342 2120 348 2121
rect 342 2116 343 2120
rect 347 2116 348 2120
rect 342 2115 348 2116
rect 414 2120 420 2121
rect 414 2116 415 2120
rect 419 2116 420 2120
rect 414 2115 420 2116
rect 478 2120 484 2121
rect 478 2116 479 2120
rect 483 2116 484 2120
rect 478 2115 484 2116
rect 542 2120 548 2121
rect 542 2116 543 2120
rect 547 2116 548 2120
rect 542 2115 548 2116
rect 606 2120 612 2121
rect 606 2116 607 2120
rect 611 2116 612 2120
rect 606 2115 612 2116
rect 670 2120 676 2121
rect 670 2116 671 2120
rect 675 2116 676 2120
rect 670 2115 676 2116
rect 734 2120 740 2121
rect 734 2116 735 2120
rect 739 2116 740 2120
rect 734 2115 740 2116
rect 790 2120 796 2121
rect 790 2116 791 2120
rect 795 2116 796 2120
rect 790 2115 796 2116
rect 838 2120 844 2121
rect 838 2116 839 2120
rect 843 2116 844 2120
rect 838 2115 844 2116
rect 886 2120 892 2121
rect 886 2116 887 2120
rect 891 2116 892 2120
rect 886 2115 892 2116
rect 934 2120 940 2121
rect 934 2116 935 2120
rect 939 2116 940 2120
rect 934 2115 940 2116
rect 990 2120 996 2121
rect 990 2116 991 2120
rect 995 2116 996 2120
rect 990 2115 996 2116
rect 1046 2120 1052 2121
rect 1278 2120 1284 2121
rect 2406 2125 2412 2126
rect 2406 2121 2407 2125
rect 2411 2121 2412 2125
rect 2406 2120 2412 2121
rect 1046 2116 1047 2120
rect 1051 2116 1052 2120
rect 1046 2115 1052 2116
rect 110 2113 116 2114
rect 110 2109 111 2113
rect 115 2109 116 2113
rect 110 2108 116 2109
rect 1238 2113 1244 2114
rect 1238 2109 1239 2113
rect 1243 2109 1244 2113
rect 1422 2111 1429 2112
rect 1238 2108 1244 2109
rect 1278 2108 1284 2109
rect 1278 2104 1279 2108
rect 1283 2104 1284 2108
rect 1422 2107 1423 2111
rect 1428 2107 1429 2111
rect 1422 2106 1429 2107
rect 1446 2111 1452 2112
rect 1446 2107 1447 2111
rect 1451 2110 1452 2111
rect 1463 2111 1469 2112
rect 1463 2110 1464 2111
rect 1451 2108 1464 2110
rect 1451 2107 1452 2108
rect 1446 2106 1452 2107
rect 1463 2107 1464 2108
rect 1468 2107 1469 2111
rect 1463 2106 1469 2107
rect 1471 2111 1477 2112
rect 1471 2107 1472 2111
rect 1476 2110 1477 2111
rect 1519 2111 1525 2112
rect 1519 2110 1520 2111
rect 1476 2108 1520 2110
rect 1476 2107 1477 2108
rect 1471 2106 1477 2107
rect 1519 2107 1520 2108
rect 1524 2107 1525 2111
rect 1519 2106 1525 2107
rect 1527 2111 1533 2112
rect 1527 2107 1528 2111
rect 1532 2110 1533 2111
rect 1591 2111 1597 2112
rect 1591 2110 1592 2111
rect 1532 2108 1592 2110
rect 1532 2107 1533 2108
rect 1527 2106 1533 2107
rect 1591 2107 1592 2108
rect 1596 2107 1597 2111
rect 1591 2106 1597 2107
rect 1599 2111 1605 2112
rect 1599 2107 1600 2111
rect 1604 2110 1605 2111
rect 1671 2111 1677 2112
rect 1671 2110 1672 2111
rect 1604 2108 1672 2110
rect 1604 2107 1605 2108
rect 1599 2106 1605 2107
rect 1671 2107 1672 2108
rect 1676 2107 1677 2111
rect 1671 2106 1677 2107
rect 1679 2111 1685 2112
rect 1679 2107 1680 2111
rect 1684 2110 1685 2111
rect 1759 2111 1765 2112
rect 1759 2110 1760 2111
rect 1684 2108 1760 2110
rect 1684 2107 1685 2108
rect 1679 2106 1685 2107
rect 1759 2107 1760 2108
rect 1764 2107 1765 2111
rect 1759 2106 1765 2107
rect 1767 2111 1773 2112
rect 1767 2107 1768 2111
rect 1772 2110 1773 2111
rect 1847 2111 1853 2112
rect 1847 2110 1848 2111
rect 1772 2108 1848 2110
rect 1772 2107 1773 2108
rect 1767 2106 1773 2107
rect 1847 2107 1848 2108
rect 1852 2107 1853 2111
rect 1847 2106 1853 2107
rect 1935 2111 1944 2112
rect 1935 2107 1936 2111
rect 1943 2107 1944 2111
rect 1935 2106 1944 2107
rect 1946 2111 1952 2112
rect 1946 2107 1947 2111
rect 1951 2110 1952 2111
rect 2023 2111 2029 2112
rect 2023 2110 2024 2111
rect 1951 2108 2024 2110
rect 1951 2107 1952 2108
rect 1946 2106 1952 2107
rect 2023 2107 2024 2108
rect 2028 2107 2029 2111
rect 2023 2106 2029 2107
rect 2031 2111 2037 2112
rect 2031 2107 2032 2111
rect 2036 2110 2037 2111
rect 2111 2111 2117 2112
rect 2111 2110 2112 2111
rect 2036 2108 2112 2110
rect 2036 2107 2037 2108
rect 2031 2106 2037 2107
rect 2111 2107 2112 2108
rect 2116 2107 2117 2111
rect 2111 2106 2117 2107
rect 2135 2111 2141 2112
rect 2135 2107 2136 2111
rect 2140 2110 2141 2111
rect 2199 2111 2205 2112
rect 2199 2110 2200 2111
rect 2140 2108 2200 2110
rect 2140 2107 2141 2108
rect 2135 2106 2141 2107
rect 2199 2107 2200 2108
rect 2204 2107 2205 2111
rect 2199 2106 2205 2107
rect 2207 2111 2213 2112
rect 2207 2107 2208 2111
rect 2212 2110 2213 2111
rect 2295 2111 2301 2112
rect 2295 2110 2296 2111
rect 2212 2108 2296 2110
rect 2212 2107 2213 2108
rect 2207 2106 2213 2107
rect 2295 2107 2296 2108
rect 2300 2107 2301 2111
rect 2295 2106 2301 2107
rect 2346 2111 2352 2112
rect 2346 2107 2347 2111
rect 2351 2110 2352 2111
rect 2383 2111 2389 2112
rect 2383 2110 2384 2111
rect 2351 2108 2384 2110
rect 2351 2107 2352 2108
rect 2346 2106 2352 2107
rect 2383 2107 2384 2108
rect 2388 2107 2389 2111
rect 2383 2106 2389 2107
rect 2406 2108 2412 2109
rect 1278 2103 1284 2104
rect 2406 2104 2407 2108
rect 2411 2104 2412 2108
rect 2406 2103 2412 2104
rect 159 2099 165 2100
rect 110 2096 116 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 159 2095 160 2099
rect 164 2098 165 2099
rect 206 2099 212 2100
rect 206 2098 207 2099
rect 164 2096 207 2098
rect 164 2095 165 2096
rect 159 2094 165 2095
rect 206 2095 207 2096
rect 211 2095 212 2099
rect 206 2094 212 2095
rect 215 2099 221 2100
rect 215 2095 216 2099
rect 220 2098 221 2099
rect 255 2099 261 2100
rect 255 2098 256 2099
rect 220 2096 256 2098
rect 220 2095 221 2096
rect 215 2094 221 2095
rect 255 2095 256 2096
rect 260 2095 261 2099
rect 255 2094 261 2095
rect 263 2099 269 2100
rect 263 2095 264 2099
rect 268 2098 269 2099
rect 295 2099 301 2100
rect 295 2098 296 2099
rect 268 2096 296 2098
rect 268 2095 269 2096
rect 263 2094 269 2095
rect 295 2095 296 2096
rect 300 2095 301 2099
rect 295 2094 301 2095
rect 367 2099 373 2100
rect 367 2095 368 2099
rect 372 2095 373 2099
rect 367 2094 373 2095
rect 375 2099 381 2100
rect 375 2095 376 2099
rect 380 2098 381 2099
rect 439 2099 445 2100
rect 439 2098 440 2099
rect 380 2096 440 2098
rect 380 2095 381 2096
rect 375 2094 381 2095
rect 439 2095 440 2096
rect 444 2095 445 2099
rect 439 2094 445 2095
rect 503 2099 512 2100
rect 503 2095 504 2099
rect 511 2095 512 2099
rect 503 2094 512 2095
rect 567 2099 573 2100
rect 567 2095 568 2099
rect 572 2098 573 2099
rect 622 2099 628 2100
rect 622 2098 623 2099
rect 572 2096 623 2098
rect 572 2095 573 2096
rect 567 2094 573 2095
rect 622 2095 623 2096
rect 627 2095 628 2099
rect 622 2094 628 2095
rect 631 2099 637 2100
rect 631 2095 632 2099
rect 636 2098 637 2099
rect 686 2099 692 2100
rect 686 2098 687 2099
rect 636 2096 687 2098
rect 636 2095 637 2096
rect 631 2094 637 2095
rect 686 2095 687 2096
rect 691 2095 692 2099
rect 686 2094 692 2095
rect 695 2099 704 2100
rect 695 2095 696 2099
rect 703 2095 704 2099
rect 695 2094 704 2095
rect 746 2099 752 2100
rect 746 2095 747 2099
rect 751 2098 752 2099
rect 759 2099 765 2100
rect 759 2098 760 2099
rect 751 2096 760 2098
rect 751 2095 752 2096
rect 746 2094 752 2095
rect 759 2095 760 2096
rect 764 2095 765 2099
rect 759 2094 765 2095
rect 767 2099 773 2100
rect 767 2095 768 2099
rect 772 2098 773 2099
rect 815 2099 821 2100
rect 815 2098 816 2099
rect 772 2096 816 2098
rect 772 2095 773 2096
rect 767 2094 773 2095
rect 815 2095 816 2096
rect 820 2095 821 2099
rect 815 2094 821 2095
rect 823 2099 829 2100
rect 823 2095 824 2099
rect 828 2098 829 2099
rect 863 2099 869 2100
rect 863 2098 864 2099
rect 828 2096 864 2098
rect 828 2095 829 2096
rect 823 2094 829 2095
rect 863 2095 864 2096
rect 868 2095 869 2099
rect 863 2094 869 2095
rect 871 2099 877 2100
rect 871 2095 872 2099
rect 876 2098 877 2099
rect 911 2099 917 2100
rect 911 2098 912 2099
rect 876 2096 912 2098
rect 876 2095 877 2096
rect 871 2094 877 2095
rect 911 2095 912 2096
rect 916 2095 917 2099
rect 911 2094 917 2095
rect 919 2099 925 2100
rect 919 2095 920 2099
rect 924 2098 925 2099
rect 959 2099 965 2100
rect 959 2098 960 2099
rect 924 2096 960 2098
rect 924 2095 925 2096
rect 919 2094 925 2095
rect 959 2095 960 2096
rect 964 2095 965 2099
rect 959 2094 965 2095
rect 967 2099 973 2100
rect 967 2095 968 2099
rect 972 2098 973 2099
rect 1015 2099 1021 2100
rect 1015 2098 1016 2099
rect 972 2096 1016 2098
rect 972 2095 973 2096
rect 967 2094 973 2095
rect 1015 2095 1016 2096
rect 1020 2095 1021 2099
rect 1015 2094 1021 2095
rect 1023 2099 1029 2100
rect 1023 2095 1024 2099
rect 1028 2098 1029 2099
rect 1071 2099 1077 2100
rect 1071 2098 1072 2099
rect 1028 2096 1072 2098
rect 1028 2095 1029 2096
rect 1023 2094 1029 2095
rect 1071 2095 1072 2096
rect 1076 2095 1077 2099
rect 1071 2094 1077 2095
rect 1238 2096 1244 2097
rect 110 2091 116 2092
rect 369 2090 371 2094
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 498 2091 504 2092
rect 1238 2091 1244 2092
rect 498 2090 499 2091
rect 369 2088 499 2090
rect 498 2087 499 2088
rect 503 2087 504 2091
rect 498 2086 504 2087
rect 1398 2085 1404 2086
rect 1398 2081 1399 2085
rect 1403 2081 1404 2085
rect 1398 2080 1404 2081
rect 1438 2085 1444 2086
rect 1438 2081 1439 2085
rect 1443 2081 1444 2085
rect 1438 2080 1444 2081
rect 1494 2085 1500 2086
rect 1494 2081 1495 2085
rect 1499 2081 1500 2085
rect 1494 2080 1500 2081
rect 1566 2085 1572 2086
rect 1566 2081 1567 2085
rect 1571 2081 1572 2085
rect 1566 2080 1572 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1734 2085 1740 2086
rect 1734 2081 1735 2085
rect 1739 2081 1740 2085
rect 1734 2080 1740 2081
rect 1822 2085 1828 2086
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1822 2080 1828 2081
rect 1910 2085 1916 2086
rect 1910 2081 1911 2085
rect 1915 2081 1916 2085
rect 1910 2080 1916 2081
rect 1998 2085 2004 2086
rect 1998 2081 1999 2085
rect 2003 2081 2004 2085
rect 1998 2080 2004 2081
rect 2086 2085 2092 2086
rect 2086 2081 2087 2085
rect 2091 2081 2092 2085
rect 2086 2080 2092 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 1423 2079 1429 2080
rect 1423 2075 1424 2079
rect 1428 2078 1429 2079
rect 1446 2079 1452 2080
rect 1446 2078 1447 2079
rect 1428 2076 1447 2078
rect 1428 2075 1429 2076
rect 1423 2074 1429 2075
rect 1446 2075 1447 2076
rect 1451 2075 1452 2079
rect 1446 2074 1452 2075
rect 1463 2079 1469 2080
rect 1463 2075 1464 2079
rect 1468 2078 1469 2079
rect 1471 2079 1477 2080
rect 1471 2078 1472 2079
rect 1468 2076 1472 2078
rect 1468 2075 1469 2076
rect 1463 2074 1469 2075
rect 1471 2075 1472 2076
rect 1476 2075 1477 2079
rect 1471 2074 1477 2075
rect 1519 2079 1525 2080
rect 1519 2075 1520 2079
rect 1524 2078 1525 2079
rect 1527 2079 1533 2080
rect 1527 2078 1528 2079
rect 1524 2076 1528 2078
rect 1524 2075 1525 2076
rect 1519 2074 1525 2075
rect 1527 2075 1528 2076
rect 1532 2075 1533 2079
rect 1527 2074 1533 2075
rect 1591 2079 1597 2080
rect 1591 2075 1592 2079
rect 1596 2078 1597 2079
rect 1599 2079 1605 2080
rect 1599 2078 1600 2079
rect 1596 2076 1600 2078
rect 1596 2075 1597 2076
rect 1591 2074 1597 2075
rect 1599 2075 1600 2076
rect 1604 2075 1605 2079
rect 1599 2074 1605 2075
rect 1671 2079 1677 2080
rect 1671 2075 1672 2079
rect 1676 2078 1677 2079
rect 1679 2079 1685 2080
rect 1679 2078 1680 2079
rect 1676 2076 1680 2078
rect 1676 2075 1677 2076
rect 1671 2074 1677 2075
rect 1679 2075 1680 2076
rect 1684 2075 1685 2079
rect 1679 2074 1685 2075
rect 1759 2079 1765 2080
rect 1759 2075 1760 2079
rect 1764 2078 1765 2079
rect 1767 2079 1773 2080
rect 1767 2078 1768 2079
rect 1764 2076 1768 2078
rect 1764 2075 1765 2076
rect 1759 2074 1765 2075
rect 1767 2075 1768 2076
rect 1772 2075 1773 2079
rect 1767 2074 1773 2075
rect 1846 2079 1853 2080
rect 1846 2075 1847 2079
rect 1852 2075 1853 2079
rect 1846 2074 1853 2075
rect 1935 2079 1941 2080
rect 1935 2075 1936 2079
rect 1940 2078 1941 2079
rect 1946 2079 1952 2080
rect 1946 2078 1947 2079
rect 1940 2076 1947 2078
rect 1940 2075 1941 2076
rect 1935 2074 1941 2075
rect 1946 2075 1947 2076
rect 1951 2075 1952 2079
rect 1946 2074 1952 2075
rect 2023 2079 2029 2080
rect 2023 2075 2024 2079
rect 2028 2078 2029 2079
rect 2031 2079 2037 2080
rect 2031 2078 2032 2079
rect 2028 2076 2032 2078
rect 2028 2075 2029 2076
rect 2023 2074 2029 2075
rect 2031 2075 2032 2076
rect 2036 2075 2037 2079
rect 2031 2074 2037 2075
rect 2111 2079 2117 2080
rect 2111 2075 2112 2079
rect 2116 2078 2117 2079
rect 2135 2079 2141 2080
rect 2135 2078 2136 2079
rect 2116 2076 2136 2078
rect 2116 2075 2117 2076
rect 2111 2074 2117 2075
rect 2135 2075 2136 2076
rect 2140 2075 2141 2079
rect 2135 2074 2141 2075
rect 2199 2079 2205 2080
rect 2199 2075 2200 2079
rect 2204 2078 2205 2079
rect 2207 2079 2213 2080
rect 2207 2078 2208 2079
rect 2204 2076 2208 2078
rect 2204 2075 2205 2076
rect 2199 2074 2205 2075
rect 2207 2075 2208 2076
rect 2212 2075 2213 2079
rect 2295 2079 2301 2080
rect 2295 2078 2296 2079
rect 2207 2074 2213 2075
rect 2216 2076 2296 2078
rect 134 2073 140 2074
rect 134 2069 135 2073
rect 139 2069 140 2073
rect 134 2068 140 2069
rect 190 2073 196 2074
rect 190 2069 191 2073
rect 195 2069 196 2073
rect 190 2068 196 2069
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 342 2073 348 2074
rect 342 2069 343 2073
rect 347 2069 348 2073
rect 342 2068 348 2069
rect 414 2073 420 2074
rect 414 2069 415 2073
rect 419 2069 420 2073
rect 478 2073 484 2074
rect 450 2071 456 2072
rect 450 2070 451 2071
rect 414 2068 420 2069
rect 439 2069 451 2070
rect 158 2067 165 2068
rect 158 2063 159 2067
rect 164 2063 165 2067
rect 158 2062 165 2063
rect 206 2067 212 2068
rect 206 2063 207 2067
rect 211 2066 212 2067
rect 215 2067 221 2068
rect 215 2066 216 2067
rect 211 2064 216 2066
rect 211 2063 212 2064
rect 206 2062 212 2063
rect 215 2063 216 2064
rect 220 2063 221 2067
rect 215 2062 221 2063
rect 255 2067 261 2068
rect 255 2063 256 2067
rect 260 2066 261 2067
rect 295 2067 301 2068
rect 295 2066 296 2067
rect 260 2064 296 2066
rect 260 2063 261 2064
rect 255 2062 261 2063
rect 295 2063 296 2064
rect 300 2063 301 2067
rect 295 2062 301 2063
rect 367 2067 373 2068
rect 367 2063 368 2067
rect 372 2066 373 2067
rect 375 2067 381 2068
rect 375 2066 376 2067
rect 372 2064 376 2066
rect 372 2063 373 2064
rect 367 2062 373 2063
rect 375 2063 376 2064
rect 380 2063 381 2067
rect 439 2065 440 2069
rect 444 2068 451 2069
rect 444 2065 445 2068
rect 450 2067 451 2068
rect 455 2067 456 2071
rect 478 2069 479 2073
rect 483 2069 484 2073
rect 478 2068 484 2069
rect 542 2073 548 2074
rect 542 2069 543 2073
rect 547 2069 548 2073
rect 542 2068 548 2069
rect 606 2073 612 2074
rect 606 2069 607 2073
rect 611 2069 612 2073
rect 606 2068 612 2069
rect 670 2073 676 2074
rect 670 2069 671 2073
rect 675 2069 676 2073
rect 670 2068 676 2069
rect 734 2073 740 2074
rect 734 2069 735 2073
rect 739 2069 740 2073
rect 734 2068 740 2069
rect 790 2073 796 2074
rect 790 2069 791 2073
rect 795 2069 796 2073
rect 790 2068 796 2069
rect 838 2073 844 2074
rect 838 2069 839 2073
rect 843 2069 844 2073
rect 838 2068 844 2069
rect 886 2073 892 2074
rect 886 2069 887 2073
rect 891 2069 892 2073
rect 886 2068 892 2069
rect 934 2073 940 2074
rect 934 2069 935 2073
rect 939 2069 940 2073
rect 934 2068 940 2069
rect 990 2073 996 2074
rect 990 2069 991 2073
rect 995 2069 996 2073
rect 990 2068 996 2069
rect 1046 2073 1052 2074
rect 1046 2069 1047 2073
rect 1051 2069 1052 2073
rect 1046 2068 1052 2069
rect 2106 2071 2112 2072
rect 450 2066 456 2067
rect 498 2067 509 2068
rect 439 2064 445 2065
rect 375 2062 381 2063
rect 498 2063 499 2067
rect 503 2063 504 2067
rect 508 2063 509 2067
rect 498 2062 509 2063
rect 567 2067 573 2068
rect 567 2063 568 2067
rect 572 2066 573 2067
rect 583 2067 589 2068
rect 583 2066 584 2067
rect 572 2064 584 2066
rect 572 2063 573 2064
rect 567 2062 573 2063
rect 583 2063 584 2064
rect 588 2063 589 2067
rect 583 2062 589 2063
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2066 628 2067
rect 631 2067 637 2068
rect 631 2066 632 2067
rect 627 2064 632 2066
rect 627 2063 628 2064
rect 622 2062 628 2063
rect 631 2063 632 2064
rect 636 2063 637 2067
rect 631 2062 637 2063
rect 686 2067 692 2068
rect 686 2063 687 2067
rect 691 2066 692 2067
rect 695 2067 701 2068
rect 695 2066 696 2067
rect 691 2064 696 2066
rect 691 2063 692 2064
rect 686 2062 692 2063
rect 695 2063 696 2064
rect 700 2063 701 2067
rect 695 2062 701 2063
rect 759 2067 765 2068
rect 759 2063 760 2067
rect 764 2066 765 2067
rect 767 2067 773 2068
rect 767 2066 768 2067
rect 764 2064 768 2066
rect 764 2063 765 2064
rect 759 2062 765 2063
rect 767 2063 768 2064
rect 772 2063 773 2067
rect 767 2062 773 2063
rect 815 2067 821 2068
rect 815 2063 816 2067
rect 820 2066 821 2067
rect 823 2067 829 2068
rect 823 2066 824 2067
rect 820 2064 824 2066
rect 820 2063 821 2064
rect 815 2062 821 2063
rect 823 2063 824 2064
rect 828 2063 829 2067
rect 823 2062 829 2063
rect 863 2067 869 2068
rect 863 2063 864 2067
rect 868 2066 869 2067
rect 871 2067 877 2068
rect 871 2066 872 2067
rect 868 2064 872 2066
rect 868 2063 869 2064
rect 863 2062 869 2063
rect 871 2063 872 2064
rect 876 2063 877 2067
rect 871 2062 877 2063
rect 911 2067 917 2068
rect 911 2063 912 2067
rect 916 2066 917 2067
rect 919 2067 925 2068
rect 919 2066 920 2067
rect 916 2064 920 2066
rect 916 2063 917 2064
rect 911 2062 917 2063
rect 919 2063 920 2064
rect 924 2063 925 2067
rect 919 2062 925 2063
rect 959 2067 965 2068
rect 959 2063 960 2067
rect 964 2066 965 2067
rect 967 2067 973 2068
rect 967 2066 968 2067
rect 964 2064 968 2066
rect 964 2063 965 2064
rect 959 2062 965 2063
rect 967 2063 968 2064
rect 972 2063 973 2067
rect 967 2062 973 2063
rect 1015 2067 1021 2068
rect 1015 2063 1016 2067
rect 1020 2066 1021 2067
rect 1023 2067 1029 2068
rect 1023 2066 1024 2067
rect 1020 2064 1024 2066
rect 1020 2063 1021 2064
rect 1015 2062 1021 2063
rect 1023 2063 1024 2064
rect 1028 2063 1029 2067
rect 1023 2062 1029 2063
rect 1070 2067 1077 2068
rect 1070 2063 1071 2067
rect 1076 2063 1077 2067
rect 2106 2067 2107 2071
rect 2111 2070 2112 2071
rect 2216 2070 2218 2076
rect 2295 2075 2296 2076
rect 2300 2075 2301 2079
rect 2295 2074 2301 2075
rect 2338 2079 2344 2080
rect 2338 2075 2339 2079
rect 2343 2078 2344 2079
rect 2383 2079 2389 2080
rect 2383 2078 2384 2079
rect 2343 2076 2384 2078
rect 2343 2075 2344 2076
rect 2338 2074 2344 2075
rect 2383 2075 2384 2076
rect 2388 2075 2389 2079
rect 2383 2074 2389 2075
rect 2111 2068 2218 2070
rect 2111 2067 2112 2068
rect 2106 2066 2112 2067
rect 1070 2062 1077 2063
rect 1942 2063 1948 2064
rect 1942 2059 1943 2063
rect 1947 2062 1948 2063
rect 2206 2063 2212 2064
rect 2206 2062 2207 2063
rect 1947 2060 2050 2062
rect 2192 2060 2207 2062
rect 1947 2059 1948 2060
rect 1942 2058 1948 2059
rect 2048 2058 2050 2060
rect 2063 2059 2069 2060
rect 2063 2058 2064 2059
rect 2048 2056 2064 2058
rect 2038 2055 2044 2056
rect 2038 2051 2039 2055
rect 2043 2051 2044 2055
rect 2063 2055 2064 2056
rect 2068 2055 2069 2059
rect 2090 2059 2096 2060
rect 2063 2054 2069 2055
rect 2078 2055 2084 2056
rect 2038 2050 2044 2051
rect 2078 2051 2079 2055
rect 2083 2051 2084 2055
rect 2090 2055 2091 2059
rect 2095 2058 2096 2059
rect 2103 2059 2109 2060
rect 2103 2058 2104 2059
rect 2095 2056 2104 2058
rect 2095 2055 2096 2056
rect 2090 2054 2096 2055
rect 2103 2055 2104 2056
rect 2108 2055 2109 2059
rect 2143 2059 2152 2060
rect 2103 2054 2109 2055
rect 2118 2055 2124 2056
rect 2078 2050 2084 2051
rect 2118 2051 2119 2055
rect 2123 2051 2124 2055
rect 2143 2055 2144 2059
rect 2151 2055 2152 2059
rect 2183 2059 2189 2060
rect 2143 2054 2152 2055
rect 2158 2055 2164 2056
rect 2118 2050 2124 2051
rect 2158 2051 2159 2055
rect 2163 2051 2164 2055
rect 2183 2055 2184 2059
rect 2188 2058 2189 2059
rect 2192 2058 2194 2060
rect 2206 2059 2207 2060
rect 2211 2059 2212 2063
rect 2254 2063 2260 2064
rect 2254 2062 2255 2063
rect 2232 2060 2255 2062
rect 2206 2058 2212 2059
rect 2223 2059 2229 2060
rect 2188 2056 2194 2058
rect 2188 2055 2189 2056
rect 2183 2054 2189 2055
rect 2198 2055 2204 2056
rect 2158 2050 2164 2051
rect 2198 2051 2199 2055
rect 2203 2051 2204 2055
rect 2223 2055 2224 2059
rect 2228 2058 2229 2059
rect 2232 2058 2234 2060
rect 2254 2059 2255 2060
rect 2259 2059 2260 2063
rect 2254 2058 2260 2059
rect 2263 2059 2272 2060
rect 2228 2056 2234 2058
rect 2228 2055 2229 2056
rect 2223 2054 2229 2055
rect 2238 2055 2244 2056
rect 2198 2050 2204 2051
rect 2238 2051 2239 2055
rect 2243 2051 2244 2055
rect 2263 2055 2264 2059
rect 2271 2055 2272 2059
rect 2294 2059 2300 2060
rect 2263 2054 2272 2055
rect 2278 2055 2284 2056
rect 2238 2050 2244 2051
rect 2278 2051 2279 2055
rect 2283 2051 2284 2055
rect 2294 2055 2295 2059
rect 2299 2058 2300 2059
rect 2303 2059 2309 2060
rect 2303 2058 2304 2059
rect 2299 2056 2304 2058
rect 2299 2055 2300 2056
rect 2294 2054 2300 2055
rect 2303 2055 2304 2056
rect 2308 2055 2309 2059
rect 2343 2059 2352 2060
rect 2303 2054 2309 2055
rect 2318 2055 2324 2056
rect 2278 2050 2284 2051
rect 2318 2051 2319 2055
rect 2323 2051 2324 2055
rect 2343 2055 2344 2059
rect 2351 2055 2352 2059
rect 2370 2059 2376 2060
rect 2343 2054 2352 2055
rect 2358 2055 2364 2056
rect 2318 2050 2324 2051
rect 2358 2051 2359 2055
rect 2363 2051 2364 2055
rect 2370 2055 2371 2059
rect 2375 2058 2376 2059
rect 2383 2059 2389 2060
rect 2383 2058 2384 2059
rect 2375 2056 2384 2058
rect 2375 2055 2376 2056
rect 2370 2054 2376 2055
rect 2383 2055 2384 2056
rect 2388 2055 2389 2059
rect 2383 2054 2389 2055
rect 2358 2050 2364 2051
rect 182 2047 188 2048
rect 182 2046 183 2047
rect 161 2044 183 2046
rect 159 2043 165 2044
rect 134 2039 140 2040
rect 134 2035 135 2039
rect 139 2035 140 2039
rect 159 2039 160 2043
rect 164 2039 165 2043
rect 182 2043 183 2044
rect 187 2043 188 2047
rect 182 2042 188 2043
rect 199 2043 208 2044
rect 159 2038 165 2039
rect 174 2039 180 2040
rect 134 2034 140 2035
rect 174 2035 175 2039
rect 179 2035 180 2039
rect 199 2039 200 2043
rect 207 2039 208 2043
rect 239 2043 245 2044
rect 199 2038 208 2039
rect 214 2039 220 2040
rect 174 2034 180 2035
rect 214 2035 215 2039
rect 219 2035 220 2039
rect 239 2039 240 2043
rect 244 2042 245 2043
rect 270 2043 276 2044
rect 270 2042 271 2043
rect 244 2040 271 2042
rect 244 2039 245 2040
rect 239 2038 245 2039
rect 270 2039 271 2040
rect 275 2039 276 2043
rect 303 2043 309 2044
rect 270 2038 276 2039
rect 278 2039 284 2040
rect 214 2034 220 2035
rect 278 2035 279 2039
rect 283 2035 284 2039
rect 303 2039 304 2043
rect 308 2042 309 2043
rect 342 2043 348 2044
rect 342 2042 343 2043
rect 308 2040 343 2042
rect 308 2039 309 2040
rect 303 2038 309 2039
rect 342 2039 343 2040
rect 347 2039 348 2043
rect 375 2043 381 2044
rect 342 2038 348 2039
rect 350 2039 356 2040
rect 278 2034 284 2035
rect 350 2035 351 2039
rect 355 2035 356 2039
rect 375 2039 376 2043
rect 380 2042 381 2043
rect 414 2043 420 2044
rect 414 2042 415 2043
rect 380 2040 415 2042
rect 380 2039 381 2040
rect 375 2038 381 2039
rect 414 2039 415 2040
rect 419 2039 420 2043
rect 434 2043 440 2044
rect 414 2038 420 2039
rect 422 2039 428 2040
rect 350 2034 356 2035
rect 422 2035 423 2039
rect 427 2035 428 2039
rect 434 2039 435 2043
rect 439 2042 440 2043
rect 447 2043 453 2044
rect 447 2042 448 2043
rect 439 2040 448 2042
rect 439 2039 440 2040
rect 434 2038 440 2039
rect 447 2039 448 2040
rect 452 2039 453 2043
rect 506 2043 517 2044
rect 447 2038 453 2039
rect 486 2039 492 2040
rect 422 2034 428 2035
rect 486 2035 487 2039
rect 491 2035 492 2039
rect 506 2039 507 2043
rect 511 2039 512 2043
rect 516 2039 517 2043
rect 562 2043 568 2044
rect 506 2038 517 2039
rect 550 2039 556 2040
rect 486 2034 492 2035
rect 550 2035 551 2039
rect 555 2035 556 2039
rect 562 2039 563 2043
rect 567 2042 568 2043
rect 575 2043 581 2044
rect 575 2042 576 2043
rect 567 2040 576 2042
rect 567 2039 568 2040
rect 562 2038 568 2039
rect 575 2039 576 2040
rect 580 2039 581 2043
rect 639 2043 645 2044
rect 575 2038 581 2039
rect 614 2039 620 2040
rect 550 2034 556 2035
rect 614 2035 615 2039
rect 619 2035 620 2039
rect 639 2039 640 2043
rect 644 2042 645 2043
rect 663 2043 669 2044
rect 663 2042 664 2043
rect 644 2040 664 2042
rect 644 2039 645 2040
rect 639 2038 645 2039
rect 663 2039 664 2040
rect 668 2039 669 2043
rect 698 2043 709 2044
rect 663 2038 669 2039
rect 678 2039 684 2040
rect 614 2034 620 2035
rect 678 2035 679 2039
rect 683 2035 684 2039
rect 698 2039 699 2043
rect 703 2039 704 2043
rect 708 2039 709 2043
rect 754 2043 760 2044
rect 698 2038 709 2039
rect 742 2039 748 2040
rect 678 2034 684 2035
rect 742 2035 743 2039
rect 747 2035 748 2039
rect 754 2039 755 2043
rect 759 2042 760 2043
rect 767 2043 773 2044
rect 767 2042 768 2043
rect 759 2040 768 2042
rect 759 2039 760 2040
rect 754 2038 760 2039
rect 767 2039 768 2040
rect 772 2039 773 2043
rect 826 2043 832 2044
rect 767 2038 773 2039
rect 814 2039 820 2040
rect 742 2034 748 2035
rect 814 2035 815 2039
rect 819 2035 820 2039
rect 826 2039 827 2043
rect 831 2042 832 2043
rect 839 2043 845 2044
rect 839 2042 840 2043
rect 831 2040 840 2042
rect 831 2039 832 2040
rect 826 2038 832 2039
rect 839 2039 840 2040
rect 844 2039 845 2043
rect 839 2038 845 2039
rect 814 2034 820 2035
rect 2146 2035 2152 2036
rect 1278 2032 1284 2033
rect 1278 2028 1279 2032
rect 1283 2028 1284 2032
rect 2146 2031 2147 2035
rect 2151 2034 2152 2035
rect 2266 2035 2272 2036
rect 2151 2032 2186 2034
rect 2151 2031 2152 2032
rect 2146 2030 2152 2031
rect 2184 2028 2186 2032
rect 2266 2031 2267 2035
rect 2271 2034 2272 2035
rect 2271 2032 2307 2034
rect 2271 2031 2272 2032
rect 2266 2030 2272 2031
rect 2305 2028 2307 2032
rect 2406 2032 2412 2033
rect 2406 2028 2407 2032
rect 2411 2028 2412 2032
rect 1278 2027 1284 2028
rect 2063 2027 2069 2028
rect 2063 2023 2064 2027
rect 2068 2026 2069 2027
rect 2090 2027 2096 2028
rect 2090 2026 2091 2027
rect 2068 2024 2091 2026
rect 2068 2023 2069 2024
rect 2063 2022 2069 2023
rect 2090 2023 2091 2024
rect 2095 2023 2096 2027
rect 2090 2022 2096 2023
rect 2103 2027 2112 2028
rect 2103 2023 2104 2027
rect 2111 2023 2112 2027
rect 2103 2022 2112 2023
rect 2143 2027 2149 2028
rect 2143 2023 2144 2027
rect 2148 2026 2149 2027
rect 2183 2027 2189 2028
rect 2148 2024 2179 2026
rect 2148 2023 2149 2024
rect 2143 2022 2149 2023
rect 754 2019 760 2020
rect 754 2018 755 2019
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 577 2016 755 2018
rect 577 2012 579 2016
rect 754 2015 755 2016
rect 759 2015 760 2019
rect 2177 2018 2179 2024
rect 2183 2023 2184 2027
rect 2188 2023 2189 2027
rect 2183 2022 2189 2023
rect 2206 2027 2212 2028
rect 2206 2023 2207 2027
rect 2211 2026 2212 2027
rect 2223 2027 2229 2028
rect 2223 2026 2224 2027
rect 2211 2024 2224 2026
rect 2211 2023 2212 2024
rect 2206 2022 2212 2023
rect 2223 2023 2224 2024
rect 2228 2023 2229 2027
rect 2223 2022 2229 2023
rect 2254 2027 2260 2028
rect 2254 2023 2255 2027
rect 2259 2026 2260 2027
rect 2263 2027 2269 2028
rect 2263 2026 2264 2027
rect 2259 2024 2264 2026
rect 2259 2023 2260 2024
rect 2254 2022 2260 2023
rect 2263 2023 2264 2024
rect 2268 2023 2269 2027
rect 2263 2022 2269 2023
rect 2303 2027 2309 2028
rect 2303 2023 2304 2027
rect 2308 2023 2309 2027
rect 2303 2022 2309 2023
rect 2343 2027 2349 2028
rect 2343 2023 2344 2027
rect 2348 2026 2349 2027
rect 2370 2027 2376 2028
rect 2370 2026 2371 2027
rect 2348 2024 2371 2026
rect 2348 2023 2349 2024
rect 2343 2022 2349 2023
rect 2370 2023 2371 2024
rect 2375 2023 2376 2027
rect 2370 2022 2376 2023
rect 2382 2027 2389 2028
rect 2406 2027 2412 2028
rect 2382 2023 2383 2027
rect 2388 2023 2389 2027
rect 2382 2022 2389 2023
rect 2214 2019 2220 2020
rect 2214 2018 2215 2019
rect 754 2014 760 2015
rect 1238 2016 1244 2017
rect 2177 2016 2215 2018
rect 1238 2012 1239 2016
rect 1243 2012 1244 2016
rect 110 2011 116 2012
rect 158 2011 165 2012
rect 158 2007 159 2011
rect 164 2007 165 2011
rect 158 2006 165 2007
rect 182 2011 188 2012
rect 182 2007 183 2011
rect 187 2010 188 2011
rect 199 2011 205 2012
rect 199 2010 200 2011
rect 187 2008 200 2010
rect 187 2007 188 2008
rect 182 2006 188 2007
rect 199 2007 200 2008
rect 204 2007 205 2011
rect 199 2006 205 2007
rect 210 2011 216 2012
rect 210 2007 211 2011
rect 215 2010 216 2011
rect 239 2011 245 2012
rect 239 2010 240 2011
rect 215 2008 240 2010
rect 215 2007 216 2008
rect 210 2006 216 2007
rect 239 2007 240 2008
rect 244 2007 245 2011
rect 239 2006 245 2007
rect 270 2011 276 2012
rect 270 2007 271 2011
rect 275 2010 276 2011
rect 303 2011 309 2012
rect 303 2010 304 2011
rect 275 2008 304 2010
rect 275 2007 276 2008
rect 270 2006 276 2007
rect 303 2007 304 2008
rect 308 2007 309 2011
rect 303 2006 309 2007
rect 342 2011 348 2012
rect 342 2007 343 2011
rect 347 2010 348 2011
rect 375 2011 381 2012
rect 375 2010 376 2011
rect 347 2008 376 2010
rect 347 2007 348 2008
rect 342 2006 348 2007
rect 375 2007 376 2008
rect 380 2007 381 2011
rect 375 2006 381 2007
rect 414 2011 420 2012
rect 414 2007 415 2011
rect 419 2010 420 2011
rect 447 2011 453 2012
rect 447 2010 448 2011
rect 419 2008 448 2010
rect 419 2007 420 2008
rect 414 2006 420 2007
rect 447 2007 448 2008
rect 452 2007 453 2011
rect 447 2006 453 2007
rect 511 2011 517 2012
rect 511 2007 512 2011
rect 516 2010 517 2011
rect 562 2011 568 2012
rect 562 2010 563 2011
rect 516 2008 563 2010
rect 516 2007 517 2008
rect 511 2006 517 2007
rect 562 2007 563 2008
rect 567 2007 568 2011
rect 562 2006 568 2007
rect 575 2011 581 2012
rect 575 2007 576 2011
rect 580 2007 581 2011
rect 575 2006 581 2007
rect 602 2011 608 2012
rect 602 2007 603 2011
rect 607 2010 608 2011
rect 639 2011 645 2012
rect 639 2010 640 2011
rect 607 2008 640 2010
rect 607 2007 608 2008
rect 602 2006 608 2007
rect 639 2007 640 2008
rect 644 2007 645 2011
rect 639 2006 645 2007
rect 663 2011 669 2012
rect 663 2007 664 2011
rect 668 2010 669 2011
rect 703 2011 709 2012
rect 703 2010 704 2011
rect 668 2008 704 2010
rect 668 2007 669 2008
rect 663 2006 669 2007
rect 703 2007 704 2008
rect 708 2007 709 2011
rect 703 2006 709 2007
rect 767 2011 773 2012
rect 767 2007 768 2011
rect 772 2010 773 2011
rect 822 2011 828 2012
rect 822 2010 823 2011
rect 772 2008 823 2010
rect 772 2007 773 2008
rect 767 2006 773 2007
rect 822 2007 823 2008
rect 827 2007 828 2011
rect 822 2006 828 2007
rect 830 2011 836 2012
rect 830 2007 831 2011
rect 835 2010 836 2011
rect 839 2011 845 2012
rect 1238 2011 1244 2012
rect 1278 2015 1284 2016
rect 1278 2011 1279 2015
rect 1283 2011 1284 2015
rect 2214 2015 2215 2016
rect 2219 2015 2220 2019
rect 2214 2014 2220 2015
rect 2406 2015 2412 2016
rect 839 2010 840 2011
rect 835 2008 840 2010
rect 835 2007 836 2008
rect 830 2006 836 2007
rect 839 2007 840 2008
rect 844 2007 845 2011
rect 1278 2010 1284 2011
rect 2406 2011 2407 2015
rect 2411 2011 2412 2015
rect 2406 2010 2412 2011
rect 839 2006 845 2007
rect 2038 2008 2044 2009
rect 2038 2004 2039 2008
rect 2043 2004 2044 2008
rect 2038 2003 2044 2004
rect 2078 2008 2084 2009
rect 2078 2004 2079 2008
rect 2083 2004 2084 2008
rect 2078 2003 2084 2004
rect 2118 2008 2124 2009
rect 2118 2004 2119 2008
rect 2123 2004 2124 2008
rect 2118 2003 2124 2004
rect 2158 2008 2164 2009
rect 2158 2004 2159 2008
rect 2163 2004 2164 2008
rect 2158 2003 2164 2004
rect 2198 2008 2204 2009
rect 2198 2004 2199 2008
rect 2203 2004 2204 2008
rect 2198 2003 2204 2004
rect 2238 2008 2244 2009
rect 2238 2004 2239 2008
rect 2243 2004 2244 2008
rect 2238 2003 2244 2004
rect 2278 2008 2284 2009
rect 2278 2004 2279 2008
rect 2283 2004 2284 2008
rect 2278 2003 2284 2004
rect 2318 2008 2324 2009
rect 2318 2004 2319 2008
rect 2323 2004 2324 2008
rect 2318 2003 2324 2004
rect 2358 2008 2364 2009
rect 2358 2004 2359 2008
rect 2363 2004 2364 2008
rect 2358 2003 2364 2004
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 1238 1999 1244 2000
rect 1238 1995 1239 1999
rect 1243 1995 1244 1999
rect 1238 1994 1244 1995
rect 1398 1996 1404 1997
rect 134 1992 140 1993
rect 134 1988 135 1992
rect 139 1988 140 1992
rect 134 1987 140 1988
rect 174 1992 180 1993
rect 174 1988 175 1992
rect 179 1988 180 1992
rect 174 1987 180 1988
rect 214 1992 220 1993
rect 214 1988 215 1992
rect 219 1988 220 1992
rect 214 1987 220 1988
rect 278 1992 284 1993
rect 278 1988 279 1992
rect 283 1988 284 1992
rect 278 1987 284 1988
rect 350 1992 356 1993
rect 350 1988 351 1992
rect 355 1988 356 1992
rect 350 1987 356 1988
rect 422 1992 428 1993
rect 422 1988 423 1992
rect 427 1988 428 1992
rect 422 1987 428 1988
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 550 1992 556 1993
rect 550 1988 551 1992
rect 555 1988 556 1992
rect 550 1987 556 1988
rect 614 1992 620 1993
rect 614 1988 615 1992
rect 619 1988 620 1992
rect 614 1987 620 1988
rect 678 1992 684 1993
rect 678 1988 679 1992
rect 683 1988 684 1992
rect 678 1987 684 1988
rect 742 1992 748 1993
rect 742 1988 743 1992
rect 747 1988 748 1992
rect 742 1987 748 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 1398 1992 1399 1996
rect 1403 1992 1404 1996
rect 1398 1991 1404 1992
rect 1438 1996 1444 1997
rect 1438 1992 1439 1996
rect 1443 1992 1444 1996
rect 1438 1991 1444 1992
rect 1478 1996 1484 1997
rect 1478 1992 1479 1996
rect 1483 1992 1484 1996
rect 1478 1991 1484 1992
rect 1518 1996 1524 1997
rect 1518 1992 1519 1996
rect 1523 1992 1524 1996
rect 1518 1991 1524 1992
rect 1558 1996 1564 1997
rect 1558 1992 1559 1996
rect 1563 1992 1564 1996
rect 1558 1991 1564 1992
rect 1598 1996 1604 1997
rect 1598 1992 1599 1996
rect 1603 1992 1604 1996
rect 1598 1991 1604 1992
rect 1638 1996 1644 1997
rect 1638 1992 1639 1996
rect 1643 1992 1644 1996
rect 1638 1991 1644 1992
rect 1678 1996 1684 1997
rect 1678 1992 1679 1996
rect 1683 1992 1684 1996
rect 1678 1991 1684 1992
rect 1718 1996 1724 1997
rect 1718 1992 1719 1996
rect 1723 1992 1724 1996
rect 1718 1991 1724 1992
rect 1766 1996 1772 1997
rect 1766 1992 1767 1996
rect 1771 1992 1772 1996
rect 1766 1991 1772 1992
rect 1822 1996 1828 1997
rect 1822 1992 1823 1996
rect 1827 1992 1828 1996
rect 1822 1991 1828 1992
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 1918 1996 1924 1997
rect 1918 1992 1919 1996
rect 1923 1992 1924 1996
rect 1918 1991 1924 1992
rect 1966 1996 1972 1997
rect 1966 1992 1967 1996
rect 1971 1992 1972 1996
rect 1966 1991 1972 1992
rect 2014 1996 2020 1997
rect 2014 1992 2015 1996
rect 2019 1992 2020 1996
rect 2014 1991 2020 1992
rect 2054 1996 2060 1997
rect 2054 1992 2055 1996
rect 2059 1992 2060 1996
rect 2054 1991 2060 1992
rect 2094 1996 2100 1997
rect 2094 1992 2095 1996
rect 2099 1992 2100 1996
rect 2094 1991 2100 1992
rect 2142 1996 2148 1997
rect 2142 1992 2143 1996
rect 2147 1992 2148 1996
rect 2142 1991 2148 1992
rect 2190 1996 2196 1997
rect 2190 1992 2191 1996
rect 2195 1992 2196 1996
rect 2190 1991 2196 1992
rect 2238 1996 2244 1997
rect 2238 1992 2239 1996
rect 2243 1992 2244 1996
rect 2238 1991 2244 1992
rect 2278 1996 2284 1997
rect 2278 1992 2279 1996
rect 2283 1992 2284 1996
rect 2278 1991 2284 1992
rect 2318 1996 2324 1997
rect 2318 1992 2319 1996
rect 2323 1992 2324 1996
rect 2318 1991 2324 1992
rect 2358 1996 2364 1997
rect 2358 1992 2359 1996
rect 2363 1992 2364 1996
rect 2358 1991 2364 1992
rect 814 1987 820 1988
rect 1278 1989 1284 1990
rect 1278 1985 1279 1989
rect 1283 1985 1284 1989
rect 1278 1984 1284 1985
rect 2406 1989 2412 1990
rect 2406 1985 2407 1989
rect 2411 1985 2412 1989
rect 2406 1984 2412 1985
rect 134 1980 140 1981
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 174 1980 180 1981
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 214 1980 220 1981
rect 214 1976 215 1980
rect 219 1976 220 1980
rect 214 1975 220 1976
rect 270 1980 276 1981
rect 270 1976 271 1980
rect 275 1976 276 1980
rect 270 1975 276 1976
rect 342 1980 348 1981
rect 342 1976 343 1980
rect 347 1976 348 1980
rect 342 1975 348 1976
rect 414 1980 420 1981
rect 414 1976 415 1980
rect 419 1976 420 1980
rect 414 1975 420 1976
rect 494 1980 500 1981
rect 494 1976 495 1980
rect 499 1976 500 1980
rect 494 1975 500 1976
rect 574 1980 580 1981
rect 574 1976 575 1980
rect 579 1976 580 1980
rect 574 1975 580 1976
rect 646 1980 652 1981
rect 646 1976 647 1980
rect 651 1976 652 1980
rect 646 1975 652 1976
rect 718 1980 724 1981
rect 718 1976 719 1980
rect 723 1976 724 1980
rect 718 1975 724 1976
rect 790 1980 796 1981
rect 790 1976 791 1980
rect 795 1976 796 1980
rect 790 1975 796 1976
rect 862 1980 868 1981
rect 862 1976 863 1980
rect 867 1976 868 1980
rect 862 1975 868 1976
rect 934 1980 940 1981
rect 934 1976 935 1980
rect 939 1976 940 1980
rect 934 1975 940 1976
rect 1006 1980 1012 1981
rect 1006 1976 1007 1980
rect 1011 1976 1012 1980
rect 1006 1975 1012 1976
rect 1423 1975 1429 1976
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 110 1968 116 1969
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1278 1972 1284 1973
rect 1278 1968 1279 1972
rect 1283 1968 1284 1972
rect 1423 1971 1424 1975
rect 1428 1974 1429 1975
rect 1446 1975 1452 1976
rect 1428 1972 1442 1974
rect 1428 1971 1429 1972
rect 1423 1970 1429 1971
rect 434 1967 440 1968
rect 1278 1967 1284 1968
rect 434 1966 435 1967
rect 161 1964 435 1966
rect 161 1960 163 1964
rect 434 1963 435 1964
rect 439 1963 440 1967
rect 1440 1966 1442 1972
rect 1446 1971 1447 1975
rect 1451 1974 1452 1975
rect 1463 1975 1469 1976
rect 1463 1974 1464 1975
rect 1451 1972 1464 1974
rect 1451 1971 1452 1972
rect 1446 1970 1452 1971
rect 1463 1971 1464 1972
rect 1468 1971 1469 1975
rect 1463 1970 1469 1971
rect 1486 1975 1492 1976
rect 1486 1971 1487 1975
rect 1491 1974 1492 1975
rect 1503 1975 1509 1976
rect 1503 1974 1504 1975
rect 1491 1972 1504 1974
rect 1491 1971 1492 1972
rect 1486 1970 1492 1971
rect 1503 1971 1504 1972
rect 1508 1971 1509 1975
rect 1503 1970 1509 1971
rect 1543 1975 1549 1976
rect 1543 1971 1544 1975
rect 1548 1974 1549 1975
rect 1574 1975 1580 1976
rect 1574 1974 1575 1975
rect 1548 1972 1575 1974
rect 1548 1971 1549 1972
rect 1543 1970 1549 1971
rect 1574 1971 1575 1972
rect 1579 1971 1580 1975
rect 1574 1970 1580 1971
rect 1583 1975 1589 1976
rect 1583 1971 1584 1975
rect 1588 1974 1589 1975
rect 1614 1975 1620 1976
rect 1614 1974 1615 1975
rect 1588 1972 1615 1974
rect 1588 1971 1589 1972
rect 1583 1970 1589 1971
rect 1614 1971 1615 1972
rect 1619 1971 1620 1975
rect 1614 1970 1620 1971
rect 1623 1975 1629 1976
rect 1623 1971 1624 1975
rect 1628 1974 1629 1975
rect 1654 1975 1660 1976
rect 1654 1974 1655 1975
rect 1628 1972 1655 1974
rect 1628 1971 1629 1972
rect 1623 1970 1629 1971
rect 1654 1971 1655 1972
rect 1659 1971 1660 1975
rect 1654 1970 1660 1971
rect 1663 1975 1669 1976
rect 1663 1971 1664 1975
rect 1668 1974 1669 1975
rect 1694 1975 1700 1976
rect 1694 1974 1695 1975
rect 1668 1972 1695 1974
rect 1668 1971 1669 1972
rect 1663 1970 1669 1971
rect 1694 1971 1695 1972
rect 1699 1971 1700 1975
rect 1694 1970 1700 1971
rect 1703 1975 1709 1976
rect 1703 1971 1704 1975
rect 1708 1974 1709 1975
rect 1734 1975 1740 1976
rect 1734 1974 1735 1975
rect 1708 1972 1735 1974
rect 1708 1971 1709 1972
rect 1703 1970 1709 1971
rect 1734 1971 1735 1972
rect 1739 1971 1740 1975
rect 1734 1970 1740 1971
rect 1743 1975 1749 1976
rect 1743 1971 1744 1975
rect 1748 1974 1749 1975
rect 1782 1975 1788 1976
rect 1782 1974 1783 1975
rect 1748 1972 1783 1974
rect 1748 1971 1749 1972
rect 1743 1970 1749 1971
rect 1782 1971 1783 1972
rect 1787 1971 1788 1975
rect 1782 1970 1788 1971
rect 1791 1975 1797 1976
rect 1791 1971 1792 1975
rect 1796 1974 1797 1975
rect 1838 1975 1844 1976
rect 1838 1974 1839 1975
rect 1796 1972 1839 1974
rect 1796 1971 1797 1972
rect 1791 1970 1797 1971
rect 1838 1971 1839 1972
rect 1843 1971 1844 1975
rect 1838 1970 1844 1971
rect 1847 1975 1853 1976
rect 1847 1971 1848 1975
rect 1852 1974 1853 1975
rect 1878 1975 1884 1976
rect 1878 1974 1879 1975
rect 1852 1972 1879 1974
rect 1852 1971 1853 1972
rect 1847 1970 1853 1971
rect 1878 1971 1879 1972
rect 1883 1971 1884 1975
rect 1878 1970 1884 1971
rect 1895 1975 1901 1976
rect 1895 1971 1896 1975
rect 1900 1974 1901 1975
rect 1942 1975 1949 1976
rect 1900 1972 1938 1974
rect 1900 1971 1901 1972
rect 1895 1970 1901 1971
rect 1542 1967 1548 1968
rect 1542 1966 1543 1967
rect 1440 1964 1543 1966
rect 434 1962 440 1963
rect 1542 1963 1543 1964
rect 1547 1963 1548 1967
rect 1936 1966 1938 1972
rect 1942 1971 1943 1975
rect 1948 1971 1949 1975
rect 1942 1970 1949 1971
rect 1951 1975 1957 1976
rect 1951 1971 1952 1975
rect 1956 1974 1957 1975
rect 1991 1975 1997 1976
rect 1991 1974 1992 1975
rect 1956 1972 1992 1974
rect 1956 1971 1957 1972
rect 1951 1970 1957 1971
rect 1991 1971 1992 1972
rect 1996 1971 1997 1975
rect 1991 1970 1997 1971
rect 2022 1975 2028 1976
rect 2022 1971 2023 1975
rect 2027 1974 2028 1975
rect 2039 1975 2045 1976
rect 2039 1974 2040 1975
rect 2027 1972 2040 1974
rect 2027 1971 2028 1972
rect 2022 1970 2028 1971
rect 2039 1971 2040 1972
rect 2044 1971 2045 1975
rect 2039 1970 2045 1971
rect 2079 1975 2088 1976
rect 2079 1971 2080 1975
rect 2087 1971 2088 1975
rect 2079 1970 2088 1971
rect 2102 1975 2108 1976
rect 2102 1971 2103 1975
rect 2107 1974 2108 1975
rect 2119 1975 2125 1976
rect 2119 1974 2120 1975
rect 2107 1972 2120 1974
rect 2107 1971 2108 1972
rect 2102 1970 2108 1971
rect 2119 1971 2120 1972
rect 2124 1971 2125 1975
rect 2119 1970 2125 1971
rect 2127 1975 2133 1976
rect 2127 1971 2128 1975
rect 2132 1974 2133 1975
rect 2167 1975 2173 1976
rect 2167 1974 2168 1975
rect 2132 1972 2168 1974
rect 2132 1971 2133 1972
rect 2127 1970 2133 1971
rect 2167 1971 2168 1972
rect 2172 1971 2173 1975
rect 2167 1970 2173 1971
rect 2175 1975 2181 1976
rect 2175 1971 2176 1975
rect 2180 1974 2181 1975
rect 2215 1975 2221 1976
rect 2215 1974 2216 1975
rect 2180 1972 2216 1974
rect 2180 1971 2181 1972
rect 2175 1970 2181 1971
rect 2215 1971 2216 1972
rect 2220 1971 2221 1975
rect 2215 1970 2221 1971
rect 2263 1975 2269 1976
rect 2263 1971 2264 1975
rect 2268 1974 2269 1975
rect 2294 1975 2300 1976
rect 2294 1974 2295 1975
rect 2268 1972 2295 1974
rect 2268 1971 2269 1972
rect 2263 1970 2269 1971
rect 2294 1971 2295 1972
rect 2299 1971 2300 1975
rect 2294 1970 2300 1971
rect 2303 1975 2309 1976
rect 2303 1971 2304 1975
rect 2308 1971 2309 1975
rect 2303 1970 2309 1971
rect 2326 1975 2332 1976
rect 2326 1971 2327 1975
rect 2331 1974 2332 1975
rect 2343 1975 2349 1976
rect 2343 1974 2344 1975
rect 2331 1972 2344 1974
rect 2331 1971 2332 1972
rect 2326 1970 2332 1971
rect 2343 1971 2344 1972
rect 2348 1971 2349 1975
rect 2343 1970 2349 1971
rect 2366 1975 2372 1976
rect 2366 1971 2367 1975
rect 2371 1974 2372 1975
rect 2383 1975 2389 1976
rect 2383 1974 2384 1975
rect 2371 1972 2384 1974
rect 2371 1971 2372 1972
rect 2366 1970 2372 1971
rect 2383 1971 2384 1972
rect 2388 1971 2389 1975
rect 2383 1970 2389 1971
rect 2406 1972 2412 1973
rect 2046 1967 2052 1968
rect 2046 1966 2047 1967
rect 1936 1964 2047 1966
rect 1542 1962 1548 1963
rect 2046 1963 2047 1964
rect 2051 1963 2052 1967
rect 2046 1962 2052 1963
rect 2286 1967 2292 1968
rect 2286 1963 2287 1967
rect 2291 1966 2292 1967
rect 2304 1966 2306 1970
rect 2406 1968 2407 1972
rect 2411 1968 2412 1972
rect 2406 1967 2412 1968
rect 2291 1964 2306 1966
rect 2291 1963 2292 1964
rect 2286 1962 2292 1963
rect 159 1959 165 1960
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 159 1955 160 1959
rect 164 1955 165 1959
rect 159 1954 165 1955
rect 182 1959 188 1960
rect 182 1955 183 1959
rect 187 1958 188 1959
rect 199 1959 205 1960
rect 199 1958 200 1959
rect 187 1956 200 1958
rect 187 1955 188 1956
rect 182 1954 188 1955
rect 199 1955 200 1956
rect 204 1955 205 1959
rect 199 1954 205 1955
rect 222 1959 228 1960
rect 222 1955 223 1959
rect 227 1958 228 1959
rect 239 1959 245 1960
rect 239 1958 240 1959
rect 227 1956 240 1958
rect 227 1955 228 1956
rect 222 1954 228 1955
rect 239 1955 240 1956
rect 244 1955 245 1959
rect 239 1954 245 1955
rect 247 1959 253 1960
rect 247 1955 248 1959
rect 252 1958 253 1959
rect 295 1959 301 1960
rect 295 1958 296 1959
rect 252 1956 296 1958
rect 252 1955 253 1956
rect 247 1954 253 1955
rect 295 1955 296 1956
rect 300 1955 301 1959
rect 295 1954 301 1955
rect 303 1959 309 1960
rect 303 1955 304 1959
rect 308 1958 309 1959
rect 367 1959 373 1960
rect 367 1958 368 1959
rect 308 1956 368 1958
rect 308 1955 309 1956
rect 303 1954 309 1955
rect 367 1955 368 1956
rect 372 1955 373 1959
rect 367 1954 373 1955
rect 375 1959 381 1960
rect 375 1955 376 1959
rect 380 1958 381 1959
rect 439 1959 445 1960
rect 439 1958 440 1959
rect 380 1956 440 1958
rect 380 1955 381 1956
rect 375 1954 381 1955
rect 439 1955 440 1956
rect 444 1955 445 1959
rect 519 1959 525 1960
rect 519 1958 520 1959
rect 439 1954 445 1955
rect 472 1956 520 1958
rect 110 1951 116 1952
rect 438 1951 444 1952
rect 438 1947 439 1951
rect 443 1950 444 1951
rect 472 1950 474 1956
rect 519 1955 520 1956
rect 524 1955 525 1959
rect 519 1954 525 1955
rect 599 1959 605 1960
rect 599 1955 600 1959
rect 604 1958 605 1959
rect 662 1959 668 1960
rect 662 1958 663 1959
rect 604 1956 663 1958
rect 604 1955 605 1956
rect 599 1954 605 1955
rect 662 1955 663 1956
rect 667 1955 668 1959
rect 662 1954 668 1955
rect 671 1959 677 1960
rect 671 1955 672 1959
rect 676 1958 677 1959
rect 682 1959 688 1960
rect 682 1958 683 1959
rect 676 1956 683 1958
rect 676 1955 677 1956
rect 671 1954 677 1955
rect 682 1955 683 1956
rect 687 1955 688 1959
rect 682 1954 688 1955
rect 690 1959 696 1960
rect 690 1955 691 1959
rect 695 1958 696 1959
rect 743 1959 749 1960
rect 743 1958 744 1959
rect 695 1956 744 1958
rect 695 1955 696 1956
rect 690 1954 696 1955
rect 743 1955 744 1956
rect 748 1955 749 1959
rect 743 1954 749 1955
rect 815 1959 821 1960
rect 815 1955 816 1959
rect 820 1958 821 1959
rect 878 1959 884 1960
rect 878 1958 879 1959
rect 820 1956 879 1958
rect 820 1955 821 1956
rect 815 1954 821 1955
rect 878 1955 879 1956
rect 883 1955 884 1959
rect 878 1954 884 1955
rect 887 1959 893 1960
rect 887 1955 888 1959
rect 892 1958 893 1959
rect 950 1959 956 1960
rect 950 1958 951 1959
rect 892 1956 951 1958
rect 892 1955 893 1956
rect 887 1954 893 1955
rect 950 1955 951 1956
rect 955 1955 956 1959
rect 950 1954 956 1955
rect 959 1959 965 1960
rect 959 1955 960 1959
rect 964 1958 965 1959
rect 1014 1959 1020 1960
rect 1014 1958 1015 1959
rect 964 1956 1015 1958
rect 964 1955 965 1956
rect 959 1954 965 1955
rect 1014 1955 1015 1956
rect 1019 1955 1020 1959
rect 1014 1954 1020 1955
rect 1022 1959 1028 1960
rect 1022 1955 1023 1959
rect 1027 1958 1028 1959
rect 1031 1959 1037 1960
rect 1031 1958 1032 1959
rect 1027 1956 1032 1958
rect 1027 1955 1028 1956
rect 1022 1954 1028 1955
rect 1031 1955 1032 1956
rect 1036 1955 1037 1959
rect 1031 1954 1037 1955
rect 1238 1956 1244 1957
rect 1238 1952 1239 1956
rect 1243 1952 1244 1956
rect 1238 1951 1244 1952
rect 443 1948 474 1950
rect 1398 1949 1404 1950
rect 443 1947 444 1948
rect 438 1946 444 1947
rect 1398 1945 1399 1949
rect 1403 1945 1404 1949
rect 1398 1944 1404 1945
rect 1438 1949 1444 1950
rect 1438 1945 1439 1949
rect 1443 1945 1444 1949
rect 1438 1944 1444 1945
rect 1478 1949 1484 1950
rect 1478 1945 1479 1949
rect 1483 1945 1484 1949
rect 1478 1944 1484 1945
rect 1518 1949 1524 1950
rect 1518 1945 1519 1949
rect 1523 1945 1524 1949
rect 1518 1944 1524 1945
rect 1558 1949 1564 1950
rect 1558 1945 1559 1949
rect 1563 1945 1564 1949
rect 1558 1944 1564 1945
rect 1598 1949 1604 1950
rect 1598 1945 1599 1949
rect 1603 1945 1604 1949
rect 1598 1944 1604 1945
rect 1638 1949 1644 1950
rect 1638 1945 1639 1949
rect 1643 1945 1644 1949
rect 1638 1944 1644 1945
rect 1678 1949 1684 1950
rect 1678 1945 1679 1949
rect 1683 1945 1684 1949
rect 1678 1944 1684 1945
rect 1718 1949 1724 1950
rect 1718 1945 1719 1949
rect 1723 1945 1724 1949
rect 1718 1944 1724 1945
rect 1766 1949 1772 1950
rect 1766 1945 1767 1949
rect 1771 1945 1772 1949
rect 1766 1944 1772 1945
rect 1822 1949 1828 1950
rect 1822 1945 1823 1949
rect 1827 1945 1828 1949
rect 1822 1944 1828 1945
rect 1870 1949 1876 1950
rect 1870 1945 1871 1949
rect 1875 1945 1876 1949
rect 1870 1944 1876 1945
rect 1918 1949 1924 1950
rect 1918 1945 1919 1949
rect 1923 1945 1924 1949
rect 1918 1944 1924 1945
rect 1966 1949 1972 1950
rect 1966 1945 1967 1949
rect 1971 1945 1972 1949
rect 1966 1944 1972 1945
rect 2014 1949 2020 1950
rect 2014 1945 2015 1949
rect 2019 1945 2020 1949
rect 2014 1944 2020 1945
rect 2054 1949 2060 1950
rect 2054 1945 2055 1949
rect 2059 1945 2060 1949
rect 2054 1944 2060 1945
rect 2094 1949 2100 1950
rect 2094 1945 2095 1949
rect 2099 1945 2100 1949
rect 2094 1944 2100 1945
rect 2142 1949 2148 1950
rect 2142 1945 2143 1949
rect 2147 1945 2148 1949
rect 2142 1944 2148 1945
rect 2190 1949 2196 1950
rect 2190 1945 2191 1949
rect 2195 1945 2196 1949
rect 2190 1944 2196 1945
rect 2238 1949 2244 1950
rect 2238 1945 2239 1949
rect 2243 1945 2244 1949
rect 2238 1944 2244 1945
rect 2278 1949 2284 1950
rect 2278 1945 2279 1949
rect 2283 1945 2284 1949
rect 2278 1944 2284 1945
rect 2318 1949 2324 1950
rect 2318 1945 2319 1949
rect 2323 1945 2324 1949
rect 2318 1944 2324 1945
rect 2358 1949 2364 1950
rect 2358 1945 2359 1949
rect 2363 1945 2364 1949
rect 2358 1944 2364 1945
rect 1423 1943 1429 1944
rect 1423 1939 1424 1943
rect 1428 1942 1429 1943
rect 1446 1943 1452 1944
rect 1446 1942 1447 1943
rect 1428 1940 1447 1942
rect 1428 1939 1429 1940
rect 1423 1938 1429 1939
rect 1446 1939 1447 1940
rect 1451 1939 1452 1943
rect 1446 1938 1452 1939
rect 1463 1943 1469 1944
rect 1463 1939 1464 1943
rect 1468 1942 1469 1943
rect 1486 1943 1492 1944
rect 1486 1942 1487 1943
rect 1468 1940 1487 1942
rect 1468 1939 1469 1940
rect 1463 1938 1469 1939
rect 1486 1939 1487 1940
rect 1491 1939 1492 1943
rect 1486 1938 1492 1939
rect 1503 1943 1509 1944
rect 1503 1939 1504 1943
rect 1508 1942 1509 1943
rect 1534 1943 1540 1944
rect 1534 1942 1535 1943
rect 1508 1940 1535 1942
rect 1508 1939 1509 1940
rect 1503 1938 1509 1939
rect 1534 1939 1535 1940
rect 1539 1939 1540 1943
rect 1534 1938 1540 1939
rect 1542 1943 1549 1944
rect 1542 1939 1543 1943
rect 1548 1939 1549 1943
rect 1542 1938 1549 1939
rect 1574 1943 1580 1944
rect 1574 1939 1575 1943
rect 1579 1942 1580 1943
rect 1583 1943 1589 1944
rect 1583 1942 1584 1943
rect 1579 1940 1584 1942
rect 1579 1939 1580 1940
rect 1574 1938 1580 1939
rect 1583 1939 1584 1940
rect 1588 1939 1589 1943
rect 1583 1938 1589 1939
rect 1614 1943 1620 1944
rect 1614 1939 1615 1943
rect 1619 1942 1620 1943
rect 1623 1943 1629 1944
rect 1623 1942 1624 1943
rect 1619 1940 1624 1942
rect 1619 1939 1620 1940
rect 1614 1938 1620 1939
rect 1623 1939 1624 1940
rect 1628 1939 1629 1943
rect 1623 1938 1629 1939
rect 1654 1943 1660 1944
rect 1654 1939 1655 1943
rect 1659 1942 1660 1943
rect 1663 1943 1669 1944
rect 1663 1942 1664 1943
rect 1659 1940 1664 1942
rect 1659 1939 1660 1940
rect 1654 1938 1660 1939
rect 1663 1939 1664 1940
rect 1668 1939 1669 1943
rect 1663 1938 1669 1939
rect 1694 1943 1700 1944
rect 1694 1939 1695 1943
rect 1699 1942 1700 1943
rect 1703 1943 1709 1944
rect 1703 1942 1704 1943
rect 1699 1940 1704 1942
rect 1699 1939 1700 1940
rect 1694 1938 1700 1939
rect 1703 1939 1704 1940
rect 1708 1939 1709 1943
rect 1703 1938 1709 1939
rect 1734 1943 1740 1944
rect 1734 1939 1735 1943
rect 1739 1942 1740 1943
rect 1743 1943 1749 1944
rect 1743 1942 1744 1943
rect 1739 1940 1744 1942
rect 1739 1939 1740 1940
rect 1734 1938 1740 1939
rect 1743 1939 1744 1940
rect 1748 1939 1749 1943
rect 1743 1938 1749 1939
rect 1782 1943 1788 1944
rect 1782 1939 1783 1943
rect 1787 1942 1788 1943
rect 1791 1943 1797 1944
rect 1791 1942 1792 1943
rect 1787 1940 1792 1942
rect 1787 1939 1788 1940
rect 1782 1938 1788 1939
rect 1791 1939 1792 1940
rect 1796 1939 1797 1943
rect 1791 1938 1797 1939
rect 1838 1943 1844 1944
rect 1838 1939 1839 1943
rect 1843 1942 1844 1943
rect 1847 1943 1853 1944
rect 1847 1942 1848 1943
rect 1843 1940 1848 1942
rect 1843 1939 1844 1940
rect 1838 1938 1844 1939
rect 1847 1939 1848 1940
rect 1852 1939 1853 1943
rect 1847 1938 1853 1939
rect 1878 1943 1884 1944
rect 1878 1939 1879 1943
rect 1883 1942 1884 1943
rect 1895 1943 1901 1944
rect 1895 1942 1896 1943
rect 1883 1940 1896 1942
rect 1883 1939 1884 1940
rect 1878 1938 1884 1939
rect 1895 1939 1896 1940
rect 1900 1939 1901 1943
rect 1895 1938 1901 1939
rect 1943 1943 1949 1944
rect 1943 1939 1944 1943
rect 1948 1942 1949 1943
rect 1951 1943 1957 1944
rect 1951 1942 1952 1943
rect 1948 1940 1952 1942
rect 1948 1939 1949 1940
rect 1943 1938 1949 1939
rect 1951 1939 1952 1940
rect 1956 1939 1957 1943
rect 1951 1938 1957 1939
rect 1991 1943 1997 1944
rect 1991 1939 1992 1943
rect 1996 1942 1997 1943
rect 2022 1943 2028 1944
rect 2022 1942 2023 1943
rect 1996 1940 2023 1942
rect 1996 1939 1997 1940
rect 1991 1938 1997 1939
rect 2022 1939 2023 1940
rect 2027 1939 2028 1943
rect 2022 1938 2028 1939
rect 2039 1943 2045 1944
rect 2039 1939 2040 1943
rect 2044 1942 2045 1943
rect 2070 1943 2076 1944
rect 2070 1942 2071 1943
rect 2044 1940 2071 1942
rect 2044 1939 2045 1940
rect 2039 1938 2045 1939
rect 2070 1939 2071 1940
rect 2075 1939 2076 1943
rect 2070 1938 2076 1939
rect 2079 1943 2085 1944
rect 2079 1939 2080 1943
rect 2084 1942 2085 1943
rect 2102 1943 2108 1944
rect 2102 1942 2103 1943
rect 2084 1940 2103 1942
rect 2084 1939 2085 1940
rect 2079 1938 2085 1939
rect 2102 1939 2103 1940
rect 2107 1939 2108 1943
rect 2102 1938 2108 1939
rect 2119 1943 2125 1944
rect 2119 1939 2120 1943
rect 2124 1942 2125 1943
rect 2127 1943 2133 1944
rect 2127 1942 2128 1943
rect 2124 1940 2128 1942
rect 2124 1939 2125 1940
rect 2119 1938 2125 1939
rect 2127 1939 2128 1940
rect 2132 1939 2133 1943
rect 2127 1938 2133 1939
rect 2167 1943 2173 1944
rect 2167 1939 2168 1943
rect 2172 1942 2173 1943
rect 2175 1943 2181 1944
rect 2175 1942 2176 1943
rect 2172 1940 2176 1942
rect 2172 1939 2173 1940
rect 2167 1938 2173 1939
rect 2175 1939 2176 1940
rect 2180 1939 2181 1943
rect 2175 1938 2181 1939
rect 2214 1943 2221 1944
rect 2214 1939 2215 1943
rect 2220 1939 2221 1943
rect 2214 1938 2221 1939
rect 2263 1943 2269 1944
rect 2263 1939 2264 1943
rect 2268 1942 2269 1943
rect 2286 1943 2292 1944
rect 2286 1942 2287 1943
rect 2268 1940 2287 1942
rect 2268 1939 2269 1940
rect 2263 1938 2269 1939
rect 2286 1939 2287 1940
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 2303 1943 2309 1944
rect 2303 1939 2304 1943
rect 2308 1942 2309 1943
rect 2326 1943 2332 1944
rect 2326 1942 2327 1943
rect 2308 1940 2327 1942
rect 2308 1939 2309 1940
rect 2303 1938 2309 1939
rect 2326 1939 2327 1940
rect 2331 1939 2332 1943
rect 2326 1938 2332 1939
rect 2343 1943 2349 1944
rect 2343 1939 2344 1943
rect 2348 1942 2349 1943
rect 2366 1943 2372 1944
rect 2366 1942 2367 1943
rect 2348 1940 2367 1942
rect 2348 1939 2349 1940
rect 2343 1938 2349 1939
rect 2366 1939 2367 1940
rect 2371 1939 2372 1943
rect 2366 1938 2372 1939
rect 2382 1943 2389 1944
rect 2382 1939 2383 1943
rect 2388 1939 2389 1943
rect 2382 1938 2389 1939
rect 134 1933 140 1934
rect 134 1929 135 1933
rect 139 1929 140 1933
rect 134 1928 140 1929
rect 174 1933 180 1934
rect 174 1929 175 1933
rect 179 1929 180 1933
rect 174 1928 180 1929
rect 214 1933 220 1934
rect 214 1929 215 1933
rect 219 1929 220 1933
rect 214 1928 220 1929
rect 270 1933 276 1934
rect 270 1929 271 1933
rect 275 1929 276 1933
rect 270 1928 276 1929
rect 342 1933 348 1934
rect 342 1929 343 1933
rect 347 1929 348 1933
rect 342 1928 348 1929
rect 414 1933 420 1934
rect 414 1929 415 1933
rect 419 1929 420 1933
rect 414 1928 420 1929
rect 494 1933 500 1934
rect 494 1929 495 1933
rect 499 1929 500 1933
rect 494 1928 500 1929
rect 574 1933 580 1934
rect 574 1929 575 1933
rect 579 1929 580 1933
rect 574 1928 580 1929
rect 646 1933 652 1934
rect 646 1929 647 1933
rect 651 1929 652 1933
rect 646 1928 652 1929
rect 718 1933 724 1934
rect 718 1929 719 1933
rect 723 1929 724 1933
rect 718 1928 724 1929
rect 790 1933 796 1934
rect 790 1929 791 1933
rect 795 1929 796 1933
rect 790 1928 796 1929
rect 862 1933 868 1934
rect 862 1929 863 1933
rect 867 1929 868 1933
rect 862 1928 868 1929
rect 934 1933 940 1934
rect 934 1929 935 1933
rect 939 1929 940 1933
rect 934 1928 940 1929
rect 1006 1933 1012 1934
rect 1006 1929 1007 1933
rect 1011 1929 1012 1933
rect 1006 1928 1012 1929
rect 159 1927 165 1928
rect 159 1923 160 1927
rect 164 1926 165 1927
rect 182 1927 188 1928
rect 182 1926 183 1927
rect 164 1924 183 1926
rect 164 1923 165 1924
rect 159 1922 165 1923
rect 182 1923 183 1924
rect 187 1923 188 1927
rect 182 1922 188 1923
rect 199 1927 205 1928
rect 199 1923 200 1927
rect 204 1926 205 1927
rect 222 1927 228 1928
rect 222 1926 223 1927
rect 204 1924 223 1926
rect 204 1923 205 1924
rect 199 1922 205 1923
rect 222 1923 223 1924
rect 227 1923 228 1927
rect 222 1922 228 1923
rect 239 1927 245 1928
rect 239 1923 240 1927
rect 244 1926 245 1927
rect 247 1927 253 1928
rect 247 1926 248 1927
rect 244 1924 248 1926
rect 244 1923 245 1924
rect 239 1922 245 1923
rect 247 1923 248 1924
rect 252 1923 253 1927
rect 247 1922 253 1923
rect 295 1927 301 1928
rect 295 1923 296 1927
rect 300 1926 301 1927
rect 303 1927 309 1928
rect 303 1926 304 1927
rect 300 1924 304 1926
rect 300 1923 301 1924
rect 295 1922 301 1923
rect 303 1923 304 1924
rect 308 1923 309 1927
rect 303 1922 309 1923
rect 367 1927 373 1928
rect 367 1923 368 1927
rect 372 1926 373 1927
rect 375 1927 381 1928
rect 375 1926 376 1927
rect 372 1924 376 1926
rect 372 1923 373 1924
rect 367 1922 373 1923
rect 375 1923 376 1924
rect 380 1923 381 1927
rect 375 1922 381 1923
rect 438 1927 445 1928
rect 438 1923 439 1927
rect 444 1923 445 1927
rect 519 1927 525 1928
rect 519 1926 520 1927
rect 438 1922 445 1923
rect 448 1924 520 1926
rect 294 1919 300 1920
rect 294 1915 295 1919
rect 299 1918 300 1919
rect 448 1918 450 1924
rect 519 1923 520 1924
rect 524 1923 525 1927
rect 519 1922 525 1923
rect 599 1927 608 1928
rect 599 1923 600 1927
rect 607 1923 608 1927
rect 599 1922 608 1923
rect 662 1927 668 1928
rect 662 1923 663 1927
rect 667 1926 668 1927
rect 671 1927 677 1928
rect 671 1926 672 1927
rect 667 1924 672 1926
rect 667 1923 668 1924
rect 662 1922 668 1923
rect 671 1923 672 1924
rect 676 1923 677 1927
rect 671 1922 677 1923
rect 682 1927 688 1928
rect 682 1923 683 1927
rect 687 1926 688 1927
rect 743 1927 749 1928
rect 743 1926 744 1927
rect 687 1924 744 1926
rect 687 1923 688 1924
rect 682 1922 688 1923
rect 743 1923 744 1924
rect 748 1923 749 1927
rect 743 1922 749 1923
rect 815 1927 821 1928
rect 815 1923 816 1927
rect 820 1926 821 1927
rect 830 1927 836 1928
rect 830 1926 831 1927
rect 820 1924 831 1926
rect 820 1923 821 1924
rect 815 1922 821 1923
rect 830 1923 831 1924
rect 835 1923 836 1927
rect 830 1922 836 1923
rect 878 1927 884 1928
rect 878 1923 879 1927
rect 883 1926 884 1927
rect 887 1927 893 1928
rect 887 1926 888 1927
rect 883 1924 888 1926
rect 883 1923 884 1924
rect 878 1922 884 1923
rect 887 1923 888 1924
rect 892 1923 893 1927
rect 887 1922 893 1923
rect 950 1927 956 1928
rect 950 1923 951 1927
rect 955 1926 956 1927
rect 959 1927 965 1928
rect 959 1926 960 1927
rect 955 1924 960 1926
rect 955 1923 956 1924
rect 950 1922 956 1923
rect 959 1923 960 1924
rect 964 1923 965 1927
rect 959 1922 965 1923
rect 1014 1927 1020 1928
rect 1014 1923 1015 1927
rect 1019 1926 1020 1927
rect 1031 1927 1037 1928
rect 1031 1926 1032 1927
rect 1019 1924 1032 1926
rect 1019 1923 1020 1924
rect 1014 1922 1020 1923
rect 1031 1923 1032 1924
rect 1036 1923 1037 1927
rect 1031 1922 1037 1923
rect 2082 1923 2088 1924
rect 299 1916 450 1918
rect 1367 1919 1376 1920
rect 299 1915 300 1916
rect 294 1914 300 1915
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1367 1915 1368 1919
rect 1375 1915 1376 1919
rect 1394 1919 1400 1920
rect 1367 1914 1376 1915
rect 1382 1915 1388 1916
rect 1342 1910 1348 1911
rect 1382 1911 1383 1915
rect 1387 1911 1388 1915
rect 1394 1915 1395 1919
rect 1399 1918 1400 1919
rect 1407 1919 1413 1920
rect 1407 1918 1408 1919
rect 1399 1916 1408 1918
rect 1399 1915 1400 1916
rect 1394 1914 1400 1915
rect 1407 1915 1408 1916
rect 1412 1915 1413 1919
rect 1434 1919 1440 1920
rect 1407 1914 1413 1915
rect 1422 1915 1428 1916
rect 1382 1910 1388 1911
rect 1422 1911 1423 1915
rect 1427 1911 1428 1915
rect 1434 1915 1435 1919
rect 1439 1918 1440 1919
rect 1447 1919 1453 1920
rect 1447 1918 1448 1919
rect 1439 1916 1448 1918
rect 1439 1915 1440 1916
rect 1434 1914 1440 1915
rect 1447 1915 1448 1916
rect 1452 1915 1453 1919
rect 1474 1919 1480 1920
rect 1447 1914 1453 1915
rect 1462 1915 1468 1916
rect 1422 1910 1428 1911
rect 1462 1911 1463 1915
rect 1467 1911 1468 1915
rect 1474 1915 1475 1919
rect 1479 1918 1480 1919
rect 1487 1919 1493 1920
rect 1487 1918 1488 1919
rect 1479 1916 1488 1918
rect 1479 1915 1480 1916
rect 1474 1914 1480 1915
rect 1487 1915 1488 1916
rect 1492 1915 1493 1919
rect 1535 1919 1541 1920
rect 1487 1914 1493 1915
rect 1510 1915 1516 1916
rect 1462 1910 1468 1911
rect 1510 1911 1511 1915
rect 1515 1911 1516 1915
rect 1535 1915 1536 1919
rect 1540 1918 1541 1919
rect 1558 1919 1564 1920
rect 1558 1918 1559 1919
rect 1540 1916 1559 1918
rect 1540 1915 1541 1916
rect 1535 1914 1541 1915
rect 1558 1915 1559 1916
rect 1563 1915 1564 1919
rect 1591 1919 1597 1920
rect 1558 1914 1564 1915
rect 1566 1915 1572 1916
rect 1510 1910 1516 1911
rect 1566 1911 1567 1915
rect 1571 1911 1572 1915
rect 1591 1915 1592 1919
rect 1596 1918 1597 1919
rect 1622 1919 1628 1920
rect 1622 1918 1623 1919
rect 1596 1916 1623 1918
rect 1596 1915 1597 1916
rect 1591 1914 1597 1915
rect 1622 1915 1623 1916
rect 1627 1915 1628 1919
rect 1642 1919 1648 1920
rect 1622 1914 1628 1915
rect 1630 1915 1636 1916
rect 1566 1910 1572 1911
rect 1630 1911 1631 1915
rect 1635 1911 1636 1915
rect 1642 1915 1643 1919
rect 1647 1918 1648 1919
rect 1655 1919 1661 1920
rect 1655 1918 1656 1919
rect 1647 1916 1656 1918
rect 1647 1915 1648 1916
rect 1642 1914 1648 1915
rect 1655 1915 1656 1916
rect 1660 1915 1661 1919
rect 1735 1919 1741 1920
rect 1655 1914 1661 1915
rect 1710 1915 1716 1916
rect 1630 1910 1636 1911
rect 1710 1911 1711 1915
rect 1715 1911 1716 1915
rect 1735 1915 1736 1919
rect 1740 1918 1741 1919
rect 1798 1919 1804 1920
rect 1798 1918 1799 1919
rect 1740 1916 1799 1918
rect 1740 1915 1741 1916
rect 1735 1914 1741 1915
rect 1798 1915 1799 1916
rect 1803 1915 1804 1919
rect 1831 1919 1837 1920
rect 1798 1914 1804 1915
rect 1806 1915 1812 1916
rect 1710 1910 1716 1911
rect 1806 1911 1807 1915
rect 1811 1911 1812 1915
rect 1831 1915 1832 1919
rect 1836 1918 1837 1919
rect 1910 1919 1916 1920
rect 1910 1918 1911 1919
rect 1836 1916 1911 1918
rect 1836 1915 1837 1916
rect 1831 1914 1837 1915
rect 1910 1915 1911 1916
rect 1915 1915 1916 1919
rect 1943 1919 1949 1920
rect 1910 1914 1916 1915
rect 1918 1915 1924 1916
rect 1806 1910 1812 1911
rect 1918 1911 1919 1915
rect 1923 1911 1924 1915
rect 1943 1915 1944 1919
rect 1948 1918 1949 1919
rect 2022 1919 2028 1920
rect 2022 1918 2023 1919
rect 1948 1916 2023 1918
rect 1948 1915 1949 1916
rect 1943 1914 1949 1915
rect 2022 1915 2023 1916
rect 2027 1915 2028 1919
rect 2046 1919 2052 1920
rect 2022 1914 2028 1915
rect 2030 1915 2036 1916
rect 1918 1910 1924 1911
rect 2030 1911 2031 1915
rect 2035 1911 2036 1915
rect 2046 1915 2047 1919
rect 2051 1918 2052 1919
rect 2055 1919 2061 1920
rect 2055 1918 2056 1919
rect 2051 1916 2056 1918
rect 2051 1915 2052 1916
rect 2046 1914 2052 1915
rect 2055 1915 2056 1916
rect 2060 1915 2061 1919
rect 2082 1919 2083 1923
rect 2087 1922 2088 1923
rect 2087 1920 2162 1922
rect 2087 1919 2088 1920
rect 2082 1918 2088 1919
rect 2160 1918 2162 1920
rect 2175 1919 2181 1920
rect 2175 1918 2176 1919
rect 2160 1916 2176 1918
rect 2055 1914 2061 1915
rect 2150 1915 2156 1916
rect 2030 1910 2036 1911
rect 2150 1911 2151 1915
rect 2155 1911 2156 1915
rect 2175 1915 2176 1916
rect 2180 1915 2181 1919
rect 2175 1914 2181 1915
rect 2150 1910 2156 1911
rect 302 1907 308 1908
rect 302 1906 303 1907
rect 280 1904 303 1906
rect 271 1903 277 1904
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1895 252 1899
rect 271 1899 272 1903
rect 276 1902 277 1903
rect 280 1902 282 1904
rect 302 1903 303 1904
rect 307 1903 308 1907
rect 1022 1907 1028 1908
rect 1022 1906 1023 1907
rect 1007 1905 1023 1906
rect 302 1902 308 1903
rect 311 1903 320 1904
rect 276 1900 282 1902
rect 276 1899 277 1900
rect 271 1898 277 1899
rect 286 1899 292 1900
rect 246 1894 252 1895
rect 286 1895 287 1899
rect 291 1895 292 1899
rect 311 1899 312 1903
rect 319 1899 320 1903
rect 351 1903 360 1904
rect 311 1898 320 1899
rect 326 1899 332 1900
rect 286 1894 292 1895
rect 326 1895 327 1899
rect 331 1895 332 1899
rect 351 1899 352 1903
rect 359 1899 360 1903
rect 391 1903 397 1904
rect 351 1898 360 1899
rect 366 1899 372 1900
rect 326 1894 332 1895
rect 366 1895 367 1899
rect 371 1895 372 1899
rect 391 1899 392 1903
rect 396 1902 397 1903
rect 406 1903 412 1904
rect 406 1902 407 1903
rect 396 1900 407 1902
rect 396 1899 397 1900
rect 391 1898 397 1899
rect 406 1899 407 1900
rect 411 1899 412 1903
rect 439 1903 445 1904
rect 406 1898 412 1899
rect 414 1899 420 1900
rect 366 1894 372 1895
rect 414 1895 415 1899
rect 419 1895 420 1899
rect 439 1899 440 1903
rect 444 1902 445 1903
rect 462 1903 468 1904
rect 462 1902 463 1903
rect 444 1900 463 1902
rect 444 1899 445 1900
rect 439 1898 445 1899
rect 462 1899 463 1900
rect 467 1899 468 1903
rect 495 1903 501 1904
rect 462 1898 468 1899
rect 470 1899 476 1900
rect 414 1894 420 1895
rect 470 1895 471 1899
rect 475 1895 476 1899
rect 495 1899 496 1903
rect 500 1902 501 1903
rect 526 1903 532 1904
rect 526 1902 527 1903
rect 500 1900 527 1902
rect 500 1899 501 1900
rect 495 1898 501 1899
rect 526 1899 527 1900
rect 531 1899 532 1903
rect 559 1903 565 1904
rect 526 1898 532 1899
rect 534 1899 540 1900
rect 470 1894 476 1895
rect 534 1895 535 1899
rect 539 1895 540 1899
rect 559 1899 560 1903
rect 564 1902 565 1903
rect 590 1903 596 1904
rect 590 1902 591 1903
rect 564 1900 591 1902
rect 564 1899 565 1900
rect 559 1898 565 1899
rect 590 1899 591 1900
rect 595 1899 596 1903
rect 610 1903 616 1904
rect 590 1898 596 1899
rect 598 1899 604 1900
rect 534 1894 540 1895
rect 598 1895 599 1899
rect 603 1895 604 1899
rect 610 1899 611 1903
rect 615 1902 616 1903
rect 623 1903 629 1904
rect 623 1902 624 1903
rect 615 1900 624 1902
rect 615 1899 616 1900
rect 610 1898 616 1899
rect 623 1899 624 1900
rect 628 1899 629 1903
rect 687 1903 696 1904
rect 623 1898 629 1899
rect 662 1899 668 1900
rect 598 1894 604 1895
rect 662 1895 663 1899
rect 667 1895 668 1899
rect 687 1899 688 1903
rect 695 1899 696 1903
rect 738 1903 744 1904
rect 687 1898 696 1899
rect 726 1899 732 1900
rect 662 1894 668 1895
rect 726 1895 727 1899
rect 731 1895 732 1899
rect 738 1899 739 1903
rect 743 1902 744 1903
rect 751 1903 757 1904
rect 751 1902 752 1903
rect 743 1900 752 1902
rect 743 1899 744 1900
rect 738 1898 744 1899
rect 751 1899 752 1900
rect 756 1899 757 1903
rect 802 1903 808 1904
rect 751 1898 757 1899
rect 790 1899 796 1900
rect 726 1894 732 1895
rect 790 1895 791 1899
rect 795 1895 796 1899
rect 802 1899 803 1903
rect 807 1902 808 1903
rect 815 1903 821 1904
rect 815 1902 816 1903
rect 807 1900 816 1902
rect 807 1899 808 1900
rect 802 1898 808 1899
rect 815 1899 816 1900
rect 820 1899 821 1903
rect 866 1903 872 1904
rect 815 1898 821 1899
rect 854 1899 860 1900
rect 790 1894 796 1895
rect 854 1895 855 1899
rect 859 1895 860 1899
rect 866 1899 867 1903
rect 871 1902 872 1903
rect 879 1903 885 1904
rect 879 1902 880 1903
rect 871 1900 880 1902
rect 871 1899 872 1900
rect 866 1898 872 1899
rect 879 1899 880 1900
rect 884 1899 885 1903
rect 943 1903 949 1904
rect 879 1898 885 1899
rect 918 1899 924 1900
rect 854 1894 860 1895
rect 918 1895 919 1899
rect 923 1895 924 1899
rect 943 1899 944 1903
rect 948 1902 949 1903
rect 974 1903 980 1904
rect 974 1902 975 1903
rect 948 1900 975 1902
rect 948 1899 949 1900
rect 943 1898 949 1899
rect 974 1899 975 1900
rect 979 1899 980 1903
rect 1007 1901 1008 1905
rect 1012 1904 1023 1905
rect 1012 1901 1013 1904
rect 1022 1903 1023 1904
rect 1027 1903 1028 1907
rect 1022 1902 1028 1903
rect 1079 1903 1085 1904
rect 1007 1900 1013 1901
rect 974 1898 980 1899
rect 982 1899 988 1900
rect 918 1894 924 1895
rect 982 1895 983 1899
rect 987 1895 988 1899
rect 982 1894 988 1895
rect 1054 1899 1060 1900
rect 1054 1895 1055 1899
rect 1059 1895 1060 1899
rect 1079 1899 1080 1903
rect 1084 1902 1085 1903
rect 1118 1903 1124 1904
rect 1118 1902 1119 1903
rect 1084 1900 1119 1902
rect 1084 1899 1085 1900
rect 1079 1898 1085 1899
rect 1118 1899 1119 1900
rect 1123 1899 1124 1903
rect 1138 1903 1144 1904
rect 1118 1898 1124 1899
rect 1126 1899 1132 1900
rect 1054 1894 1060 1895
rect 1126 1895 1127 1899
rect 1131 1895 1132 1899
rect 1138 1899 1139 1903
rect 1143 1902 1144 1903
rect 1151 1903 1157 1904
rect 1151 1902 1152 1903
rect 1143 1900 1152 1902
rect 1143 1899 1144 1900
rect 1138 1898 1144 1899
rect 1151 1899 1152 1900
rect 1156 1899 1157 1903
rect 1151 1898 1157 1899
rect 1126 1894 1132 1895
rect 1642 1895 1648 1896
rect 1642 1894 1643 1895
rect 1278 1892 1284 1893
rect 1278 1888 1279 1892
rect 1283 1888 1284 1892
rect 1528 1892 1643 1894
rect 1278 1887 1284 1888
rect 1367 1887 1373 1888
rect 1367 1883 1368 1887
rect 1372 1886 1373 1887
rect 1394 1887 1400 1888
rect 1394 1886 1395 1887
rect 1372 1884 1395 1886
rect 1372 1883 1373 1884
rect 1367 1882 1373 1883
rect 1394 1883 1395 1884
rect 1399 1883 1400 1887
rect 1394 1882 1400 1883
rect 1407 1887 1413 1888
rect 1407 1883 1408 1887
rect 1412 1886 1413 1887
rect 1434 1887 1440 1888
rect 1434 1886 1435 1887
rect 1412 1884 1435 1886
rect 1412 1883 1413 1884
rect 1407 1882 1413 1883
rect 1434 1883 1435 1884
rect 1439 1883 1440 1887
rect 1434 1882 1440 1883
rect 1447 1887 1453 1888
rect 1447 1883 1448 1887
rect 1452 1886 1453 1887
rect 1474 1887 1480 1888
rect 1474 1886 1475 1887
rect 1452 1884 1475 1886
rect 1452 1883 1453 1884
rect 1447 1882 1453 1883
rect 1474 1883 1475 1884
rect 1479 1883 1480 1887
rect 1474 1882 1480 1883
rect 1487 1887 1493 1888
rect 1487 1883 1488 1887
rect 1492 1886 1493 1887
rect 1528 1886 1530 1892
rect 1642 1891 1643 1892
rect 1647 1891 1648 1895
rect 1642 1890 1648 1891
rect 2406 1892 2412 1893
rect 2406 1888 2407 1892
rect 2411 1888 2412 1892
rect 1492 1884 1530 1886
rect 1534 1887 1541 1888
rect 1492 1883 1493 1884
rect 1487 1882 1493 1883
rect 1534 1883 1535 1887
rect 1540 1883 1541 1887
rect 1534 1882 1541 1883
rect 1558 1887 1564 1888
rect 1558 1883 1559 1887
rect 1563 1886 1564 1887
rect 1591 1887 1597 1888
rect 1591 1886 1592 1887
rect 1563 1884 1592 1886
rect 1563 1883 1564 1884
rect 1558 1882 1564 1883
rect 1591 1883 1592 1884
rect 1596 1883 1597 1887
rect 1591 1882 1597 1883
rect 1622 1887 1628 1888
rect 1622 1883 1623 1887
rect 1627 1886 1628 1887
rect 1655 1887 1661 1888
rect 1655 1886 1656 1887
rect 1627 1884 1656 1886
rect 1627 1883 1628 1884
rect 1622 1882 1628 1883
rect 1655 1883 1656 1884
rect 1660 1883 1661 1887
rect 1655 1882 1661 1883
rect 1703 1887 1709 1888
rect 1703 1883 1704 1887
rect 1708 1886 1709 1887
rect 1735 1887 1741 1888
rect 1735 1886 1736 1887
rect 1708 1884 1736 1886
rect 1708 1883 1709 1884
rect 1703 1882 1709 1883
rect 1735 1883 1736 1884
rect 1740 1883 1741 1887
rect 1735 1882 1741 1883
rect 1798 1887 1804 1888
rect 1798 1883 1799 1887
rect 1803 1886 1804 1887
rect 1831 1887 1837 1888
rect 1831 1886 1832 1887
rect 1803 1884 1832 1886
rect 1803 1883 1804 1884
rect 1798 1882 1804 1883
rect 1831 1883 1832 1884
rect 1836 1883 1837 1887
rect 1831 1882 1837 1883
rect 1910 1887 1916 1888
rect 1910 1883 1911 1887
rect 1915 1886 1916 1887
rect 1943 1887 1949 1888
rect 1943 1886 1944 1887
rect 1915 1884 1944 1886
rect 1915 1883 1916 1884
rect 1910 1882 1916 1883
rect 1943 1883 1944 1884
rect 1948 1883 1949 1887
rect 1943 1882 1949 1883
rect 2022 1887 2028 1888
rect 2022 1883 2023 1887
rect 2027 1886 2028 1887
rect 2055 1887 2061 1888
rect 2055 1886 2056 1887
rect 2027 1884 2056 1886
rect 2027 1883 2028 1884
rect 2022 1882 2028 1883
rect 2055 1883 2056 1884
rect 2060 1883 2061 1887
rect 2055 1882 2061 1883
rect 2070 1887 2076 1888
rect 2070 1883 2071 1887
rect 2075 1886 2076 1887
rect 2175 1887 2181 1888
rect 2406 1887 2412 1888
rect 2175 1886 2176 1887
rect 2075 1884 2176 1886
rect 2075 1883 2076 1884
rect 2070 1882 2076 1883
rect 2175 1883 2176 1884
rect 2180 1883 2181 1887
rect 2175 1882 2181 1883
rect 314 1879 320 1880
rect 110 1876 116 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 294 1875 300 1876
rect 294 1874 295 1875
rect 110 1871 116 1872
rect 271 1873 295 1874
rect 271 1869 272 1873
rect 276 1872 295 1873
rect 276 1869 277 1872
rect 294 1871 295 1872
rect 299 1871 300 1875
rect 314 1875 315 1879
rect 319 1878 320 1879
rect 1138 1879 1144 1880
rect 1138 1878 1139 1879
rect 319 1875 321 1878
rect 314 1874 321 1875
rect 294 1870 300 1871
rect 302 1871 308 1872
rect 271 1868 277 1869
rect 302 1867 303 1871
rect 307 1870 308 1871
rect 311 1871 317 1872
rect 311 1870 312 1871
rect 307 1868 312 1870
rect 307 1867 308 1868
rect 302 1866 308 1867
rect 311 1867 312 1868
rect 316 1867 317 1871
rect 319 1870 321 1874
rect 968 1876 1139 1878
rect 351 1871 357 1872
rect 351 1870 352 1871
rect 319 1868 352 1870
rect 311 1866 317 1867
rect 351 1867 352 1868
rect 356 1867 357 1871
rect 351 1866 357 1867
rect 362 1871 368 1872
rect 362 1867 363 1871
rect 367 1870 368 1871
rect 391 1871 397 1872
rect 391 1870 392 1871
rect 367 1868 392 1870
rect 367 1867 368 1868
rect 362 1866 368 1867
rect 391 1867 392 1868
rect 396 1867 397 1871
rect 391 1866 397 1867
rect 406 1871 412 1872
rect 406 1867 407 1871
rect 411 1870 412 1871
rect 439 1871 445 1872
rect 439 1870 440 1871
rect 411 1868 440 1870
rect 411 1867 412 1868
rect 406 1866 412 1867
rect 439 1867 440 1868
rect 444 1867 445 1871
rect 439 1866 445 1867
rect 462 1871 468 1872
rect 462 1867 463 1871
rect 467 1870 468 1871
rect 495 1871 501 1872
rect 495 1870 496 1871
rect 467 1868 496 1870
rect 467 1867 468 1868
rect 462 1866 468 1867
rect 495 1867 496 1868
rect 500 1867 501 1871
rect 495 1866 501 1867
rect 526 1871 532 1872
rect 526 1867 527 1871
rect 531 1870 532 1871
rect 559 1871 565 1872
rect 559 1870 560 1871
rect 531 1868 560 1870
rect 531 1867 532 1868
rect 526 1866 532 1867
rect 559 1867 560 1868
rect 564 1867 565 1871
rect 559 1866 565 1867
rect 590 1871 596 1872
rect 590 1867 591 1871
rect 595 1870 596 1871
rect 623 1871 629 1872
rect 623 1870 624 1871
rect 595 1868 624 1870
rect 595 1867 596 1868
rect 590 1866 596 1867
rect 623 1867 624 1868
rect 628 1867 629 1871
rect 623 1866 629 1867
rect 687 1871 693 1872
rect 687 1867 688 1871
rect 692 1870 693 1871
rect 738 1871 744 1872
rect 738 1870 739 1871
rect 692 1868 739 1870
rect 692 1867 693 1868
rect 687 1866 693 1867
rect 738 1867 739 1868
rect 743 1867 744 1871
rect 738 1866 744 1867
rect 751 1871 757 1872
rect 751 1867 752 1871
rect 756 1870 757 1871
rect 802 1871 808 1872
rect 802 1870 803 1871
rect 756 1868 803 1870
rect 756 1867 757 1868
rect 751 1866 757 1867
rect 802 1867 803 1868
rect 807 1867 808 1871
rect 802 1866 808 1867
rect 815 1871 821 1872
rect 815 1867 816 1871
rect 820 1870 821 1871
rect 862 1871 868 1872
rect 862 1870 863 1871
rect 820 1868 863 1870
rect 820 1867 821 1868
rect 815 1866 821 1867
rect 862 1867 863 1868
rect 867 1867 868 1871
rect 862 1866 868 1867
rect 870 1871 876 1872
rect 870 1867 871 1871
rect 875 1870 876 1871
rect 879 1871 885 1872
rect 879 1870 880 1871
rect 875 1868 880 1870
rect 875 1867 876 1868
rect 870 1866 876 1867
rect 879 1867 880 1868
rect 884 1867 885 1871
rect 879 1866 885 1867
rect 943 1871 949 1872
rect 943 1867 944 1871
rect 948 1870 949 1871
rect 968 1870 970 1876
rect 1138 1875 1139 1876
rect 1143 1875 1144 1879
rect 1138 1874 1144 1875
rect 1238 1876 1244 1877
rect 1238 1872 1239 1876
rect 1243 1872 1244 1876
rect 948 1868 970 1870
rect 974 1871 980 1872
rect 948 1867 949 1868
rect 943 1866 949 1867
rect 974 1867 975 1871
rect 979 1870 980 1871
rect 1007 1871 1013 1872
rect 1007 1870 1008 1871
rect 979 1868 1008 1870
rect 979 1867 980 1868
rect 974 1866 980 1867
rect 1007 1867 1008 1868
rect 1012 1867 1013 1871
rect 1007 1866 1013 1867
rect 1070 1871 1076 1872
rect 1070 1867 1071 1871
rect 1075 1870 1076 1871
rect 1079 1871 1085 1872
rect 1079 1870 1080 1871
rect 1075 1868 1080 1870
rect 1075 1867 1076 1868
rect 1070 1866 1076 1867
rect 1079 1867 1080 1868
rect 1084 1867 1085 1871
rect 1079 1866 1085 1867
rect 1118 1871 1124 1872
rect 1118 1867 1119 1871
rect 1123 1870 1124 1871
rect 1151 1871 1157 1872
rect 1238 1871 1244 1872
rect 1278 1875 1284 1876
rect 1278 1871 1279 1875
rect 1283 1871 1284 1875
rect 1151 1870 1152 1871
rect 1123 1868 1152 1870
rect 1123 1867 1124 1868
rect 1118 1866 1124 1867
rect 1151 1867 1152 1868
rect 1156 1867 1157 1871
rect 1278 1870 1284 1871
rect 2406 1875 2412 1876
rect 2406 1871 2407 1875
rect 2411 1871 2412 1875
rect 2406 1870 2412 1871
rect 1151 1866 1157 1867
rect 1342 1868 1348 1869
rect 1342 1864 1343 1868
rect 1347 1864 1348 1868
rect 1342 1863 1348 1864
rect 1382 1868 1388 1869
rect 1382 1864 1383 1868
rect 1387 1864 1388 1868
rect 1382 1863 1388 1864
rect 1422 1868 1428 1869
rect 1422 1864 1423 1868
rect 1427 1864 1428 1868
rect 1422 1863 1428 1864
rect 1462 1868 1468 1869
rect 1462 1864 1463 1868
rect 1467 1864 1468 1868
rect 1462 1863 1468 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1566 1868 1572 1869
rect 1566 1864 1567 1868
rect 1571 1864 1572 1868
rect 1566 1863 1572 1864
rect 1630 1868 1636 1869
rect 1630 1864 1631 1868
rect 1635 1864 1636 1868
rect 1630 1863 1636 1864
rect 1710 1868 1716 1869
rect 1710 1864 1711 1868
rect 1715 1864 1716 1868
rect 1710 1863 1716 1864
rect 1806 1868 1812 1869
rect 1806 1864 1807 1868
rect 1811 1864 1812 1868
rect 1806 1863 1812 1864
rect 1918 1868 1924 1869
rect 1918 1864 1919 1868
rect 1923 1864 1924 1868
rect 1918 1863 1924 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2150 1868 2156 1869
rect 2150 1864 2151 1868
rect 2155 1864 2156 1868
rect 2150 1863 2156 1864
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 110 1854 116 1855
rect 1238 1859 1244 1860
rect 1238 1855 1239 1859
rect 1243 1855 1244 1859
rect 1238 1854 1244 1855
rect 246 1852 252 1853
rect 246 1848 247 1852
rect 251 1848 252 1852
rect 246 1847 252 1848
rect 286 1852 292 1853
rect 286 1848 287 1852
rect 291 1848 292 1852
rect 286 1847 292 1848
rect 326 1852 332 1853
rect 326 1848 327 1852
rect 331 1848 332 1852
rect 326 1847 332 1848
rect 366 1852 372 1853
rect 366 1848 367 1852
rect 371 1848 372 1852
rect 366 1847 372 1848
rect 414 1852 420 1853
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 470 1852 476 1853
rect 470 1848 471 1852
rect 475 1848 476 1852
rect 470 1847 476 1848
rect 534 1852 540 1853
rect 534 1848 535 1852
rect 539 1848 540 1852
rect 534 1847 540 1848
rect 598 1852 604 1853
rect 598 1848 599 1852
rect 603 1848 604 1852
rect 598 1847 604 1848
rect 662 1852 668 1853
rect 662 1848 663 1852
rect 667 1848 668 1852
rect 662 1847 668 1848
rect 726 1852 732 1853
rect 726 1848 727 1852
rect 731 1848 732 1852
rect 726 1847 732 1848
rect 790 1852 796 1853
rect 790 1848 791 1852
rect 795 1848 796 1852
rect 790 1847 796 1848
rect 854 1852 860 1853
rect 854 1848 855 1852
rect 859 1848 860 1852
rect 854 1847 860 1848
rect 918 1852 924 1853
rect 918 1848 919 1852
rect 923 1848 924 1852
rect 918 1847 924 1848
rect 982 1852 988 1853
rect 982 1848 983 1852
rect 987 1848 988 1852
rect 982 1847 988 1848
rect 1054 1852 1060 1853
rect 1054 1848 1055 1852
rect 1059 1848 1060 1852
rect 1054 1847 1060 1848
rect 1126 1852 1132 1853
rect 1126 1848 1127 1852
rect 1131 1848 1132 1852
rect 1126 1847 1132 1848
rect 1358 1848 1364 1849
rect 1358 1844 1359 1848
rect 1363 1844 1364 1848
rect 1358 1843 1364 1844
rect 1398 1848 1404 1849
rect 1398 1844 1399 1848
rect 1403 1844 1404 1848
rect 1398 1843 1404 1844
rect 1446 1848 1452 1849
rect 1446 1844 1447 1848
rect 1451 1844 1452 1848
rect 1446 1843 1452 1844
rect 1502 1848 1508 1849
rect 1502 1844 1503 1848
rect 1507 1844 1508 1848
rect 1502 1843 1508 1844
rect 1558 1848 1564 1849
rect 1558 1844 1559 1848
rect 1563 1844 1564 1848
rect 1558 1843 1564 1844
rect 1614 1848 1620 1849
rect 1614 1844 1615 1848
rect 1619 1844 1620 1848
rect 1614 1843 1620 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1726 1848 1732 1849
rect 1726 1844 1727 1848
rect 1731 1844 1732 1848
rect 1726 1843 1732 1844
rect 1782 1848 1788 1849
rect 1782 1844 1783 1848
rect 1787 1844 1788 1848
rect 1782 1843 1788 1844
rect 1838 1848 1844 1849
rect 1838 1844 1839 1848
rect 1843 1844 1844 1848
rect 1838 1843 1844 1844
rect 1894 1848 1900 1849
rect 1894 1844 1895 1848
rect 1899 1844 1900 1848
rect 1894 1843 1900 1844
rect 1950 1848 1956 1849
rect 1950 1844 1951 1848
rect 1955 1844 1956 1848
rect 1950 1843 1956 1844
rect 1278 1841 1284 1842
rect 1278 1837 1279 1841
rect 1283 1837 1284 1841
rect 398 1836 404 1837
rect 398 1832 399 1836
rect 403 1832 404 1836
rect 398 1831 404 1832
rect 438 1836 444 1837
rect 438 1832 439 1836
rect 443 1832 444 1836
rect 438 1831 444 1832
rect 478 1836 484 1837
rect 478 1832 479 1836
rect 483 1832 484 1836
rect 478 1831 484 1832
rect 518 1836 524 1837
rect 518 1832 519 1836
rect 523 1832 524 1836
rect 518 1831 524 1832
rect 566 1836 572 1837
rect 566 1832 567 1836
rect 571 1832 572 1836
rect 566 1831 572 1832
rect 622 1836 628 1837
rect 622 1832 623 1836
rect 627 1832 628 1836
rect 622 1831 628 1832
rect 686 1836 692 1837
rect 686 1832 687 1836
rect 691 1832 692 1836
rect 686 1831 692 1832
rect 758 1836 764 1837
rect 758 1832 759 1836
rect 763 1832 764 1836
rect 758 1831 764 1832
rect 830 1836 836 1837
rect 830 1832 831 1836
rect 835 1832 836 1836
rect 830 1831 836 1832
rect 902 1836 908 1837
rect 902 1832 903 1836
rect 907 1832 908 1836
rect 902 1831 908 1832
rect 974 1836 980 1837
rect 974 1832 975 1836
rect 979 1832 980 1836
rect 974 1831 980 1832
rect 1046 1836 1052 1837
rect 1046 1832 1047 1836
rect 1051 1832 1052 1836
rect 1046 1831 1052 1832
rect 1126 1836 1132 1837
rect 1126 1832 1127 1836
rect 1131 1832 1132 1836
rect 1126 1831 1132 1832
rect 1190 1836 1196 1837
rect 1278 1836 1284 1837
rect 2406 1841 2412 1842
rect 2406 1837 2407 1841
rect 2411 1837 2412 1841
rect 2406 1836 2412 1837
rect 1190 1832 1191 1836
rect 1195 1832 1196 1836
rect 1190 1831 1196 1832
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 1238 1829 1244 1830
rect 1238 1825 1239 1829
rect 1243 1825 1244 1829
rect 1370 1827 1376 1828
rect 1238 1824 1244 1825
rect 1278 1824 1284 1825
rect 610 1823 616 1824
rect 610 1822 611 1823
rect 440 1820 611 1822
rect 423 1815 429 1816
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 423 1811 424 1815
rect 428 1814 429 1815
rect 440 1814 442 1820
rect 610 1819 611 1820
rect 615 1819 616 1823
rect 1278 1820 1279 1824
rect 1283 1820 1284 1824
rect 1370 1823 1371 1827
rect 1375 1826 1376 1827
rect 1383 1827 1389 1828
rect 1383 1826 1384 1827
rect 1375 1824 1384 1826
rect 1375 1823 1376 1824
rect 1370 1822 1376 1823
rect 1383 1823 1384 1824
rect 1388 1823 1389 1827
rect 1383 1822 1389 1823
rect 1406 1827 1412 1828
rect 1406 1823 1407 1827
rect 1411 1826 1412 1827
rect 1423 1827 1429 1828
rect 1423 1826 1424 1827
rect 1411 1824 1424 1826
rect 1411 1823 1412 1824
rect 1406 1822 1412 1823
rect 1423 1823 1424 1824
rect 1428 1823 1429 1827
rect 1423 1822 1429 1823
rect 1431 1827 1437 1828
rect 1431 1823 1432 1827
rect 1436 1826 1437 1827
rect 1471 1827 1477 1828
rect 1471 1826 1472 1827
rect 1436 1824 1472 1826
rect 1436 1823 1437 1824
rect 1431 1822 1437 1823
rect 1471 1823 1472 1824
rect 1476 1823 1477 1827
rect 1471 1822 1477 1823
rect 1479 1827 1485 1828
rect 1479 1823 1480 1827
rect 1484 1826 1485 1827
rect 1527 1827 1533 1828
rect 1527 1826 1528 1827
rect 1484 1824 1528 1826
rect 1484 1823 1485 1824
rect 1479 1822 1485 1823
rect 1527 1823 1528 1824
rect 1532 1823 1533 1827
rect 1527 1822 1533 1823
rect 1535 1827 1541 1828
rect 1535 1823 1536 1827
rect 1540 1826 1541 1827
rect 1583 1827 1589 1828
rect 1583 1826 1584 1827
rect 1540 1824 1584 1826
rect 1540 1823 1541 1824
rect 1535 1822 1541 1823
rect 1583 1823 1584 1824
rect 1588 1823 1589 1827
rect 1583 1822 1589 1823
rect 1591 1827 1597 1828
rect 1591 1823 1592 1827
rect 1596 1826 1597 1827
rect 1639 1827 1645 1828
rect 1639 1826 1640 1827
rect 1596 1824 1640 1826
rect 1596 1823 1597 1824
rect 1591 1822 1597 1823
rect 1639 1823 1640 1824
rect 1644 1823 1645 1827
rect 1639 1822 1645 1823
rect 1695 1827 1701 1828
rect 1695 1823 1696 1827
rect 1700 1826 1701 1827
rect 1742 1827 1748 1828
rect 1742 1826 1743 1827
rect 1700 1824 1743 1826
rect 1700 1823 1701 1824
rect 1695 1822 1701 1823
rect 1742 1823 1743 1824
rect 1747 1823 1748 1827
rect 1742 1822 1748 1823
rect 1751 1827 1757 1828
rect 1751 1823 1752 1827
rect 1756 1826 1757 1827
rect 1798 1827 1804 1828
rect 1798 1826 1799 1827
rect 1756 1824 1799 1826
rect 1756 1823 1757 1824
rect 1751 1822 1757 1823
rect 1798 1823 1799 1824
rect 1803 1823 1804 1827
rect 1798 1822 1804 1823
rect 1807 1827 1813 1828
rect 1807 1823 1808 1827
rect 1812 1826 1813 1827
rect 1854 1827 1860 1828
rect 1854 1826 1855 1827
rect 1812 1824 1855 1826
rect 1812 1823 1813 1824
rect 1807 1822 1813 1823
rect 1854 1823 1855 1824
rect 1859 1823 1860 1827
rect 1854 1822 1860 1823
rect 1863 1827 1869 1828
rect 1863 1823 1864 1827
rect 1868 1826 1869 1827
rect 1902 1827 1908 1828
rect 1868 1824 1898 1826
rect 1868 1823 1869 1824
rect 1863 1822 1869 1823
rect 1278 1819 1284 1820
rect 610 1818 616 1819
rect 1896 1818 1898 1824
rect 1902 1823 1903 1827
rect 1907 1826 1908 1827
rect 1919 1827 1925 1828
rect 1919 1826 1920 1827
rect 1907 1824 1920 1826
rect 1907 1823 1908 1824
rect 1902 1822 1908 1823
rect 1919 1823 1920 1824
rect 1924 1823 1925 1827
rect 1919 1822 1925 1823
rect 1927 1827 1933 1828
rect 1927 1823 1928 1827
rect 1932 1826 1933 1827
rect 1975 1827 1981 1828
rect 1975 1826 1976 1827
rect 1932 1824 1976 1826
rect 1932 1823 1933 1824
rect 1927 1822 1933 1823
rect 1975 1823 1976 1824
rect 1980 1823 1981 1827
rect 1975 1822 1981 1823
rect 2406 1824 2412 1825
rect 2406 1820 2407 1824
rect 2411 1820 2412 1824
rect 1974 1819 1980 1820
rect 2406 1819 2412 1820
rect 1974 1818 1975 1819
rect 1896 1816 1975 1818
rect 428 1812 442 1814
rect 446 1815 452 1816
rect 428 1811 429 1812
rect 423 1810 429 1811
rect 446 1811 447 1815
rect 451 1814 452 1815
rect 463 1815 469 1816
rect 463 1814 464 1815
rect 451 1812 464 1814
rect 451 1811 452 1812
rect 446 1810 452 1811
rect 463 1811 464 1812
rect 468 1811 469 1815
rect 463 1810 469 1811
rect 486 1815 492 1816
rect 486 1811 487 1815
rect 491 1814 492 1815
rect 503 1815 509 1816
rect 503 1814 504 1815
rect 491 1812 504 1814
rect 491 1811 492 1812
rect 486 1810 492 1811
rect 503 1811 504 1812
rect 508 1811 509 1815
rect 503 1810 509 1811
rect 526 1815 532 1816
rect 526 1811 527 1815
rect 531 1814 532 1815
rect 543 1815 549 1816
rect 543 1814 544 1815
rect 531 1812 544 1814
rect 531 1811 532 1812
rect 526 1810 532 1811
rect 543 1811 544 1812
rect 548 1811 549 1815
rect 543 1810 549 1811
rect 551 1815 557 1816
rect 551 1811 552 1815
rect 556 1814 557 1815
rect 591 1815 597 1816
rect 591 1814 592 1815
rect 556 1812 592 1814
rect 556 1811 557 1812
rect 551 1810 557 1811
rect 591 1811 592 1812
rect 596 1811 597 1815
rect 591 1810 597 1811
rect 599 1815 605 1816
rect 599 1811 600 1815
rect 604 1814 605 1815
rect 647 1815 653 1816
rect 647 1814 648 1815
rect 604 1812 648 1814
rect 604 1811 605 1812
rect 599 1810 605 1811
rect 647 1811 648 1812
rect 652 1811 653 1815
rect 647 1810 653 1811
rect 655 1815 661 1816
rect 655 1811 656 1815
rect 660 1814 661 1815
rect 711 1815 717 1816
rect 711 1814 712 1815
rect 660 1812 712 1814
rect 660 1811 661 1812
rect 655 1810 661 1811
rect 711 1811 712 1812
rect 716 1811 717 1815
rect 711 1810 717 1811
rect 783 1815 789 1816
rect 783 1811 784 1815
rect 788 1811 789 1815
rect 783 1810 789 1811
rect 791 1815 797 1816
rect 791 1811 792 1815
rect 796 1814 797 1815
rect 855 1815 861 1816
rect 855 1814 856 1815
rect 796 1812 856 1814
rect 796 1811 797 1812
rect 791 1810 797 1811
rect 855 1811 856 1812
rect 860 1811 861 1815
rect 855 1810 861 1811
rect 927 1815 933 1816
rect 927 1811 928 1815
rect 932 1814 933 1815
rect 958 1815 964 1816
rect 958 1814 959 1815
rect 932 1812 959 1814
rect 932 1811 933 1812
rect 927 1810 933 1811
rect 958 1811 959 1812
rect 963 1811 964 1815
rect 958 1810 964 1811
rect 999 1815 1005 1816
rect 999 1811 1000 1815
rect 1004 1811 1005 1815
rect 999 1810 1005 1811
rect 1007 1815 1013 1816
rect 1007 1811 1008 1815
rect 1012 1814 1013 1815
rect 1071 1815 1077 1816
rect 1071 1814 1072 1815
rect 1012 1812 1072 1814
rect 1012 1811 1013 1812
rect 1007 1810 1013 1811
rect 1071 1811 1072 1812
rect 1076 1811 1077 1815
rect 1071 1810 1077 1811
rect 1151 1815 1157 1816
rect 1151 1811 1152 1815
rect 1156 1814 1157 1815
rect 1206 1815 1212 1816
rect 1206 1814 1207 1815
rect 1156 1812 1207 1814
rect 1156 1811 1157 1812
rect 1151 1810 1157 1811
rect 1206 1811 1207 1812
rect 1211 1811 1212 1815
rect 1206 1810 1212 1811
rect 1215 1815 1221 1816
rect 1215 1811 1216 1815
rect 1220 1811 1221 1815
rect 1974 1815 1975 1816
rect 1979 1815 1980 1819
rect 1974 1814 1980 1815
rect 1215 1810 1221 1811
rect 1238 1812 1244 1813
rect 110 1807 116 1808
rect 784 1806 786 1810
rect 926 1807 932 1808
rect 926 1806 927 1807
rect 784 1804 927 1806
rect 926 1803 927 1804
rect 931 1803 932 1807
rect 1000 1806 1002 1810
rect 1150 1807 1156 1808
rect 1150 1806 1151 1807
rect 1000 1804 1151 1806
rect 926 1802 932 1803
rect 1150 1803 1151 1804
rect 1155 1803 1156 1807
rect 1150 1802 1156 1803
rect 1170 1807 1176 1808
rect 1170 1803 1171 1807
rect 1175 1806 1176 1807
rect 1217 1806 1219 1810
rect 1238 1808 1239 1812
rect 1243 1808 1244 1812
rect 1238 1807 1244 1808
rect 1175 1804 1219 1806
rect 1175 1803 1176 1804
rect 1170 1802 1176 1803
rect 1358 1801 1364 1802
rect 1358 1797 1359 1801
rect 1363 1797 1364 1801
rect 1358 1796 1364 1797
rect 1398 1801 1404 1802
rect 1398 1797 1399 1801
rect 1403 1797 1404 1801
rect 1398 1796 1404 1797
rect 1446 1801 1452 1802
rect 1446 1797 1447 1801
rect 1451 1797 1452 1801
rect 1446 1796 1452 1797
rect 1502 1801 1508 1802
rect 1502 1797 1503 1801
rect 1507 1797 1508 1801
rect 1502 1796 1508 1797
rect 1558 1801 1564 1802
rect 1558 1797 1559 1801
rect 1563 1797 1564 1801
rect 1558 1796 1564 1797
rect 1614 1801 1620 1802
rect 1614 1797 1615 1801
rect 1619 1797 1620 1801
rect 1614 1796 1620 1797
rect 1670 1801 1676 1802
rect 1670 1797 1671 1801
rect 1675 1797 1676 1801
rect 1670 1796 1676 1797
rect 1726 1801 1732 1802
rect 1726 1797 1727 1801
rect 1731 1797 1732 1801
rect 1726 1796 1732 1797
rect 1782 1801 1788 1802
rect 1782 1797 1783 1801
rect 1787 1797 1788 1801
rect 1782 1796 1788 1797
rect 1838 1801 1844 1802
rect 1838 1797 1839 1801
rect 1843 1797 1844 1801
rect 1838 1796 1844 1797
rect 1894 1801 1900 1802
rect 1894 1797 1895 1801
rect 1899 1797 1900 1801
rect 1894 1796 1900 1797
rect 1950 1801 1956 1802
rect 1950 1797 1951 1801
rect 1955 1797 1956 1801
rect 1950 1796 1956 1797
rect 1383 1795 1389 1796
rect 1383 1791 1384 1795
rect 1388 1794 1389 1795
rect 1406 1795 1412 1796
rect 1406 1794 1407 1795
rect 1388 1792 1407 1794
rect 1388 1791 1389 1792
rect 1383 1790 1389 1791
rect 1406 1791 1407 1792
rect 1411 1791 1412 1795
rect 1406 1790 1412 1791
rect 1423 1795 1429 1796
rect 1423 1791 1424 1795
rect 1428 1794 1429 1795
rect 1431 1795 1437 1796
rect 1431 1794 1432 1795
rect 1428 1792 1432 1794
rect 1428 1791 1429 1792
rect 1423 1790 1429 1791
rect 1431 1791 1432 1792
rect 1436 1791 1437 1795
rect 1431 1790 1437 1791
rect 1471 1795 1477 1796
rect 1471 1791 1472 1795
rect 1476 1794 1477 1795
rect 1479 1795 1485 1796
rect 1479 1794 1480 1795
rect 1476 1792 1480 1794
rect 1476 1791 1477 1792
rect 1471 1790 1477 1791
rect 1479 1791 1480 1792
rect 1484 1791 1485 1795
rect 1479 1790 1485 1791
rect 1527 1795 1533 1796
rect 1527 1791 1528 1795
rect 1532 1794 1533 1795
rect 1535 1795 1541 1796
rect 1535 1794 1536 1795
rect 1532 1792 1536 1794
rect 1532 1791 1533 1792
rect 1527 1790 1533 1791
rect 1535 1791 1536 1792
rect 1540 1791 1541 1795
rect 1535 1790 1541 1791
rect 1583 1795 1589 1796
rect 1583 1791 1584 1795
rect 1588 1794 1589 1795
rect 1591 1795 1597 1796
rect 1591 1794 1592 1795
rect 1588 1792 1592 1794
rect 1588 1791 1589 1792
rect 1583 1790 1589 1791
rect 1591 1791 1592 1792
rect 1596 1791 1597 1795
rect 1591 1790 1597 1791
rect 1602 1795 1608 1796
rect 1602 1791 1603 1795
rect 1607 1794 1608 1795
rect 1639 1795 1645 1796
rect 1639 1794 1640 1795
rect 1607 1792 1640 1794
rect 1607 1791 1608 1792
rect 1602 1790 1608 1791
rect 1639 1791 1640 1792
rect 1644 1791 1645 1795
rect 1639 1790 1645 1791
rect 1695 1795 1701 1796
rect 1695 1791 1696 1795
rect 1700 1794 1701 1795
rect 1703 1795 1709 1796
rect 1703 1794 1704 1795
rect 1700 1792 1704 1794
rect 1700 1791 1701 1792
rect 1695 1790 1701 1791
rect 1703 1791 1704 1792
rect 1708 1791 1709 1795
rect 1703 1790 1709 1791
rect 1742 1795 1748 1796
rect 1742 1791 1743 1795
rect 1747 1794 1748 1795
rect 1751 1795 1757 1796
rect 1751 1794 1752 1795
rect 1747 1792 1752 1794
rect 1747 1791 1748 1792
rect 1742 1790 1748 1791
rect 1751 1791 1752 1792
rect 1756 1791 1757 1795
rect 1751 1790 1757 1791
rect 1798 1795 1804 1796
rect 1798 1791 1799 1795
rect 1803 1794 1804 1795
rect 1807 1795 1813 1796
rect 1807 1794 1808 1795
rect 1803 1792 1808 1794
rect 1803 1791 1804 1792
rect 1798 1790 1804 1791
rect 1807 1791 1808 1792
rect 1812 1791 1813 1795
rect 1807 1790 1813 1791
rect 1854 1795 1860 1796
rect 1854 1791 1855 1795
rect 1859 1794 1860 1795
rect 1863 1795 1869 1796
rect 1863 1794 1864 1795
rect 1859 1792 1864 1794
rect 1859 1791 1860 1792
rect 1854 1790 1860 1791
rect 1863 1791 1864 1792
rect 1868 1791 1869 1795
rect 1863 1790 1869 1791
rect 1919 1795 1925 1796
rect 1919 1791 1920 1795
rect 1924 1794 1925 1795
rect 1927 1795 1933 1796
rect 1927 1794 1928 1795
rect 1924 1792 1928 1794
rect 1924 1791 1925 1792
rect 1919 1790 1925 1791
rect 1927 1791 1928 1792
rect 1932 1791 1933 1795
rect 1927 1790 1933 1791
rect 1974 1795 1981 1796
rect 1974 1791 1975 1795
rect 1980 1791 1981 1795
rect 1974 1790 1981 1791
rect 398 1789 404 1790
rect 398 1785 399 1789
rect 403 1785 404 1789
rect 398 1784 404 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 478 1789 484 1790
rect 478 1785 479 1789
rect 483 1785 484 1789
rect 478 1784 484 1785
rect 518 1789 524 1790
rect 518 1785 519 1789
rect 523 1785 524 1789
rect 518 1784 524 1785
rect 566 1789 572 1790
rect 566 1785 567 1789
rect 571 1785 572 1789
rect 566 1784 572 1785
rect 622 1789 628 1790
rect 622 1785 623 1789
rect 627 1785 628 1789
rect 622 1784 628 1785
rect 686 1789 692 1790
rect 686 1785 687 1789
rect 691 1785 692 1789
rect 686 1784 692 1785
rect 758 1789 764 1790
rect 758 1785 759 1789
rect 763 1785 764 1789
rect 758 1784 764 1785
rect 830 1789 836 1790
rect 830 1785 831 1789
rect 835 1785 836 1789
rect 902 1789 908 1790
rect 870 1787 876 1788
rect 870 1786 871 1787
rect 830 1784 836 1785
rect 855 1785 871 1786
rect 423 1783 429 1784
rect 423 1779 424 1783
rect 428 1782 429 1783
rect 446 1783 452 1784
rect 446 1782 447 1783
rect 428 1780 447 1782
rect 428 1779 429 1780
rect 423 1778 429 1779
rect 446 1779 447 1780
rect 451 1779 452 1783
rect 446 1778 452 1779
rect 463 1783 469 1784
rect 463 1779 464 1783
rect 468 1782 469 1783
rect 486 1783 492 1784
rect 486 1782 487 1783
rect 468 1780 487 1782
rect 468 1779 469 1780
rect 463 1778 469 1779
rect 486 1779 487 1780
rect 491 1779 492 1783
rect 486 1778 492 1779
rect 503 1783 509 1784
rect 503 1779 504 1783
rect 508 1782 509 1783
rect 526 1783 532 1784
rect 526 1782 527 1783
rect 508 1780 527 1782
rect 508 1779 509 1780
rect 503 1778 509 1779
rect 526 1779 527 1780
rect 531 1779 532 1783
rect 526 1778 532 1779
rect 543 1783 549 1784
rect 543 1779 544 1783
rect 548 1782 549 1783
rect 551 1783 557 1784
rect 551 1782 552 1783
rect 548 1780 552 1782
rect 548 1779 549 1780
rect 543 1778 549 1779
rect 551 1779 552 1780
rect 556 1779 557 1783
rect 551 1778 557 1779
rect 591 1783 597 1784
rect 591 1779 592 1783
rect 596 1782 597 1783
rect 599 1783 605 1784
rect 599 1782 600 1783
rect 596 1780 600 1782
rect 596 1779 597 1780
rect 591 1778 597 1779
rect 599 1779 600 1780
rect 604 1779 605 1783
rect 599 1778 605 1779
rect 647 1783 653 1784
rect 647 1779 648 1783
rect 652 1782 653 1783
rect 655 1783 661 1784
rect 655 1782 656 1783
rect 652 1780 656 1782
rect 652 1779 653 1780
rect 647 1778 653 1779
rect 655 1779 656 1780
rect 660 1779 661 1783
rect 655 1778 661 1779
rect 674 1783 680 1784
rect 674 1779 675 1783
rect 679 1782 680 1783
rect 711 1783 717 1784
rect 711 1782 712 1783
rect 679 1780 712 1782
rect 679 1779 680 1780
rect 674 1778 680 1779
rect 711 1779 712 1780
rect 716 1779 717 1783
rect 711 1778 717 1779
rect 783 1783 789 1784
rect 783 1779 784 1783
rect 788 1782 789 1783
rect 791 1783 797 1784
rect 791 1782 792 1783
rect 788 1780 792 1782
rect 788 1779 789 1780
rect 783 1778 789 1779
rect 791 1779 792 1780
rect 796 1779 797 1783
rect 855 1781 856 1785
rect 860 1784 871 1785
rect 860 1781 861 1784
rect 870 1783 871 1784
rect 875 1783 876 1787
rect 902 1785 903 1789
rect 907 1785 908 1789
rect 902 1784 908 1785
rect 974 1789 980 1790
rect 974 1785 975 1789
rect 979 1785 980 1789
rect 974 1784 980 1785
rect 1046 1789 1052 1790
rect 1046 1785 1047 1789
rect 1051 1785 1052 1789
rect 1046 1784 1052 1785
rect 1126 1789 1132 1790
rect 1126 1785 1127 1789
rect 1131 1785 1132 1789
rect 1126 1784 1132 1785
rect 1190 1789 1196 1790
rect 1190 1785 1191 1789
rect 1195 1785 1196 1789
rect 1190 1784 1196 1785
rect 870 1782 876 1783
rect 926 1783 933 1784
rect 855 1780 861 1781
rect 791 1778 797 1779
rect 926 1779 927 1783
rect 932 1779 933 1783
rect 926 1778 933 1779
rect 999 1783 1005 1784
rect 999 1779 1000 1783
rect 1004 1782 1005 1783
rect 1007 1783 1013 1784
rect 1007 1782 1008 1783
rect 1004 1780 1008 1782
rect 1004 1779 1005 1780
rect 999 1778 1005 1779
rect 1007 1779 1008 1780
rect 1012 1779 1013 1783
rect 1007 1778 1013 1779
rect 1070 1783 1077 1784
rect 1070 1779 1071 1783
rect 1076 1779 1077 1783
rect 1070 1778 1077 1779
rect 1150 1783 1157 1784
rect 1150 1779 1151 1783
rect 1156 1779 1157 1783
rect 1150 1778 1157 1779
rect 1206 1783 1212 1784
rect 1206 1779 1207 1783
rect 1211 1782 1212 1783
rect 1215 1783 1221 1784
rect 1215 1782 1216 1783
rect 1211 1780 1216 1782
rect 1211 1779 1212 1780
rect 1206 1778 1212 1779
rect 1215 1779 1216 1780
rect 1220 1779 1221 1783
rect 1215 1778 1221 1779
rect 431 1763 440 1764
rect 406 1759 412 1760
rect 406 1755 407 1759
rect 411 1755 412 1759
rect 431 1759 432 1763
rect 439 1759 440 1763
rect 458 1763 464 1764
rect 431 1758 440 1759
rect 446 1759 452 1760
rect 406 1754 412 1755
rect 446 1755 447 1759
rect 451 1755 452 1759
rect 458 1759 459 1763
rect 463 1762 464 1763
rect 471 1763 477 1764
rect 471 1762 472 1763
rect 463 1760 472 1762
rect 463 1759 464 1760
rect 458 1758 464 1759
rect 471 1759 472 1760
rect 476 1759 477 1763
rect 498 1763 504 1764
rect 471 1758 477 1759
rect 486 1759 492 1760
rect 446 1754 452 1755
rect 486 1755 487 1759
rect 491 1755 492 1759
rect 498 1759 499 1763
rect 503 1762 504 1763
rect 511 1763 517 1764
rect 511 1762 512 1763
rect 503 1760 512 1762
rect 503 1759 504 1760
rect 498 1758 504 1759
rect 511 1759 512 1760
rect 516 1759 517 1763
rect 538 1763 544 1764
rect 511 1758 517 1759
rect 526 1759 532 1760
rect 486 1754 492 1755
rect 526 1755 527 1759
rect 531 1755 532 1759
rect 538 1759 539 1763
rect 543 1762 544 1763
rect 551 1763 557 1764
rect 551 1762 552 1763
rect 543 1760 552 1762
rect 543 1759 544 1760
rect 538 1758 544 1759
rect 551 1759 552 1760
rect 556 1759 557 1763
rect 578 1763 584 1764
rect 551 1758 557 1759
rect 566 1759 572 1760
rect 526 1754 532 1755
rect 566 1755 567 1759
rect 571 1755 572 1759
rect 578 1759 579 1763
rect 583 1762 584 1763
rect 591 1763 597 1764
rect 591 1762 592 1763
rect 583 1760 592 1762
rect 583 1759 584 1760
rect 578 1758 584 1759
rect 591 1759 592 1760
rect 596 1759 597 1763
rect 618 1763 624 1764
rect 591 1758 597 1759
rect 606 1759 612 1760
rect 566 1754 572 1755
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 618 1759 619 1763
rect 623 1762 624 1763
rect 631 1763 637 1764
rect 631 1762 632 1763
rect 623 1760 632 1762
rect 623 1759 624 1760
rect 618 1758 624 1759
rect 631 1759 632 1760
rect 636 1759 637 1763
rect 658 1763 664 1764
rect 631 1758 637 1759
rect 646 1759 652 1760
rect 606 1754 612 1755
rect 646 1755 647 1759
rect 651 1755 652 1759
rect 658 1759 659 1763
rect 663 1762 664 1763
rect 671 1763 677 1764
rect 671 1762 672 1763
rect 663 1760 672 1762
rect 663 1759 664 1760
rect 658 1758 664 1759
rect 671 1759 672 1760
rect 676 1759 677 1763
rect 719 1763 725 1764
rect 671 1758 677 1759
rect 694 1759 700 1760
rect 646 1754 652 1755
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 719 1759 720 1763
rect 724 1762 725 1763
rect 742 1763 748 1764
rect 742 1762 743 1763
rect 724 1760 743 1762
rect 724 1759 725 1760
rect 719 1758 725 1759
rect 742 1759 743 1760
rect 747 1759 748 1763
rect 775 1763 781 1764
rect 742 1758 748 1759
rect 750 1759 756 1760
rect 694 1754 700 1755
rect 750 1755 751 1759
rect 755 1755 756 1759
rect 775 1759 776 1763
rect 780 1762 781 1763
rect 798 1763 804 1764
rect 798 1762 799 1763
rect 780 1760 799 1762
rect 780 1759 781 1760
rect 775 1758 781 1759
rect 798 1759 799 1760
rect 803 1759 804 1763
rect 831 1763 837 1764
rect 798 1758 804 1759
rect 806 1759 812 1760
rect 750 1754 756 1755
rect 806 1755 807 1759
rect 811 1755 812 1759
rect 831 1759 832 1763
rect 836 1762 837 1763
rect 862 1763 868 1764
rect 862 1762 863 1763
rect 836 1760 863 1762
rect 836 1759 837 1760
rect 831 1758 837 1759
rect 862 1759 863 1760
rect 867 1759 868 1763
rect 895 1763 901 1764
rect 862 1758 868 1759
rect 870 1759 876 1760
rect 806 1754 812 1755
rect 870 1755 871 1759
rect 875 1755 876 1759
rect 895 1759 896 1763
rect 900 1762 901 1763
rect 926 1763 932 1764
rect 926 1762 927 1763
rect 900 1760 927 1762
rect 900 1759 901 1760
rect 895 1758 901 1759
rect 926 1759 927 1760
rect 931 1759 932 1763
rect 958 1763 965 1764
rect 926 1758 932 1759
rect 934 1759 940 1760
rect 870 1754 876 1755
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 958 1759 959 1763
rect 964 1759 965 1763
rect 1023 1763 1029 1764
rect 958 1758 965 1759
rect 998 1759 1004 1760
rect 934 1754 940 1755
rect 998 1755 999 1759
rect 1003 1755 1004 1759
rect 1023 1759 1024 1763
rect 1028 1762 1029 1763
rect 1095 1763 1101 1764
rect 1028 1760 1066 1762
rect 1028 1759 1029 1760
rect 1023 1758 1029 1759
rect 998 1754 1004 1755
rect 1064 1750 1066 1760
rect 1070 1759 1076 1760
rect 1070 1755 1071 1759
rect 1075 1755 1076 1759
rect 1095 1759 1096 1763
rect 1100 1762 1101 1763
rect 1126 1763 1132 1764
rect 1126 1762 1127 1763
rect 1100 1760 1127 1762
rect 1100 1759 1101 1760
rect 1095 1758 1101 1759
rect 1126 1759 1127 1760
rect 1131 1759 1132 1763
rect 1167 1763 1176 1764
rect 1126 1758 1132 1759
rect 1142 1759 1148 1760
rect 1070 1754 1076 1755
rect 1142 1755 1143 1759
rect 1147 1755 1148 1759
rect 1167 1759 1168 1763
rect 1175 1759 1176 1763
rect 1202 1763 1208 1764
rect 1167 1758 1176 1759
rect 1190 1759 1196 1760
rect 1142 1754 1148 1755
rect 1190 1755 1191 1759
rect 1195 1755 1196 1759
rect 1202 1759 1203 1763
rect 1207 1762 1208 1763
rect 1215 1763 1221 1764
rect 1215 1762 1216 1763
rect 1207 1760 1216 1762
rect 1207 1759 1208 1760
rect 1202 1758 1208 1759
rect 1215 1759 1216 1760
rect 1220 1759 1221 1763
rect 1314 1763 1320 1764
rect 1215 1758 1221 1759
rect 1302 1759 1308 1760
rect 1190 1754 1196 1755
rect 1302 1755 1303 1759
rect 1307 1755 1308 1759
rect 1314 1759 1315 1763
rect 1319 1762 1320 1763
rect 1327 1763 1333 1764
rect 1327 1762 1328 1763
rect 1319 1760 1328 1762
rect 1319 1759 1320 1760
rect 1314 1758 1320 1759
rect 1327 1759 1328 1760
rect 1332 1759 1333 1763
rect 1354 1763 1360 1764
rect 1327 1758 1333 1759
rect 1342 1759 1348 1760
rect 1302 1754 1308 1755
rect 1342 1755 1343 1759
rect 1347 1755 1348 1759
rect 1354 1759 1355 1763
rect 1359 1762 1360 1763
rect 1367 1763 1373 1764
rect 1367 1762 1368 1763
rect 1359 1760 1368 1762
rect 1359 1759 1360 1760
rect 1354 1758 1360 1759
rect 1367 1759 1368 1760
rect 1372 1759 1373 1763
rect 1415 1763 1421 1764
rect 1367 1758 1373 1759
rect 1390 1759 1396 1760
rect 1342 1754 1348 1755
rect 1390 1755 1391 1759
rect 1395 1755 1396 1759
rect 1415 1759 1416 1763
rect 1420 1762 1421 1763
rect 1446 1763 1452 1764
rect 1446 1762 1447 1763
rect 1420 1760 1447 1762
rect 1420 1759 1421 1760
rect 1415 1758 1421 1759
rect 1446 1759 1447 1760
rect 1451 1759 1452 1763
rect 1479 1763 1485 1764
rect 1446 1758 1452 1759
rect 1454 1759 1460 1760
rect 1390 1754 1396 1755
rect 1454 1755 1455 1759
rect 1459 1755 1460 1759
rect 1479 1759 1480 1763
rect 1484 1762 1485 1763
rect 1510 1763 1516 1764
rect 1510 1762 1511 1763
rect 1484 1760 1511 1762
rect 1484 1759 1485 1760
rect 1479 1758 1485 1759
rect 1510 1759 1511 1760
rect 1515 1759 1516 1763
rect 1543 1763 1549 1764
rect 1510 1758 1516 1759
rect 1518 1759 1524 1760
rect 1454 1754 1460 1755
rect 1518 1755 1519 1759
rect 1523 1755 1524 1759
rect 1543 1759 1544 1763
rect 1548 1762 1549 1763
rect 1574 1763 1580 1764
rect 1574 1762 1575 1763
rect 1548 1760 1575 1762
rect 1548 1759 1549 1760
rect 1543 1758 1549 1759
rect 1574 1759 1575 1760
rect 1579 1759 1580 1763
rect 1594 1763 1600 1764
rect 1574 1758 1580 1759
rect 1582 1759 1588 1760
rect 1518 1754 1524 1755
rect 1582 1755 1583 1759
rect 1587 1755 1588 1759
rect 1594 1759 1595 1763
rect 1599 1762 1600 1763
rect 1607 1763 1613 1764
rect 1607 1762 1608 1763
rect 1599 1760 1608 1762
rect 1599 1759 1600 1760
rect 1594 1758 1600 1759
rect 1607 1759 1608 1760
rect 1612 1759 1613 1763
rect 1671 1763 1677 1764
rect 1607 1758 1613 1759
rect 1646 1759 1652 1760
rect 1582 1754 1588 1755
rect 1646 1755 1647 1759
rect 1651 1755 1652 1759
rect 1671 1759 1672 1763
rect 1676 1762 1677 1763
rect 1694 1763 1700 1764
rect 1694 1762 1695 1763
rect 1676 1760 1695 1762
rect 1676 1759 1677 1760
rect 1671 1758 1677 1759
rect 1694 1759 1695 1760
rect 1699 1759 1700 1763
rect 1727 1763 1733 1764
rect 1694 1758 1700 1759
rect 1702 1759 1708 1760
rect 1646 1754 1652 1755
rect 1702 1755 1703 1759
rect 1707 1755 1708 1759
rect 1727 1759 1728 1763
rect 1732 1762 1733 1763
rect 1750 1763 1756 1764
rect 1750 1762 1751 1763
rect 1732 1760 1751 1762
rect 1732 1759 1733 1760
rect 1727 1758 1733 1759
rect 1750 1759 1751 1760
rect 1755 1759 1756 1763
rect 1783 1763 1789 1764
rect 1750 1758 1756 1759
rect 1758 1759 1764 1760
rect 1702 1754 1708 1755
rect 1758 1755 1759 1759
rect 1763 1755 1764 1759
rect 1783 1759 1784 1763
rect 1788 1762 1789 1763
rect 1798 1763 1804 1764
rect 1798 1762 1799 1763
rect 1788 1760 1799 1762
rect 1788 1759 1789 1760
rect 1783 1758 1789 1759
rect 1798 1759 1799 1760
rect 1803 1759 1804 1763
rect 1831 1763 1837 1764
rect 1831 1762 1832 1763
rect 1816 1760 1832 1762
rect 1798 1758 1804 1759
rect 1806 1759 1812 1760
rect 1758 1754 1764 1755
rect 1806 1755 1807 1759
rect 1811 1755 1812 1759
rect 1806 1754 1812 1755
rect 1094 1751 1100 1752
rect 1094 1750 1095 1751
rect 1064 1748 1095 1750
rect 1094 1747 1095 1748
rect 1099 1747 1100 1751
rect 1094 1746 1100 1747
rect 1674 1751 1680 1752
rect 1674 1747 1675 1751
rect 1679 1750 1680 1751
rect 1816 1750 1818 1760
rect 1831 1759 1832 1760
rect 1836 1759 1837 1763
rect 1887 1763 1893 1764
rect 1831 1758 1837 1759
rect 1862 1759 1868 1760
rect 1862 1755 1863 1759
rect 1867 1755 1868 1759
rect 1887 1759 1888 1763
rect 1892 1762 1893 1763
rect 1902 1763 1908 1764
rect 1902 1762 1903 1763
rect 1892 1760 1903 1762
rect 1892 1759 1893 1760
rect 1887 1758 1893 1759
rect 1902 1759 1903 1760
rect 1907 1759 1908 1763
rect 1943 1763 1949 1764
rect 1902 1758 1908 1759
rect 1918 1759 1924 1760
rect 1862 1754 1868 1755
rect 1918 1755 1919 1759
rect 1923 1755 1924 1759
rect 1943 1759 1944 1763
rect 1948 1762 1949 1763
rect 1966 1763 1972 1764
rect 1966 1762 1967 1763
rect 1948 1760 1967 1762
rect 1948 1759 1949 1760
rect 1943 1758 1949 1759
rect 1966 1759 1967 1760
rect 1971 1759 1972 1763
rect 1999 1763 2005 1764
rect 1966 1758 1972 1759
rect 1974 1759 1980 1760
rect 1918 1754 1924 1755
rect 1974 1755 1975 1759
rect 1979 1755 1980 1759
rect 1974 1754 1980 1755
rect 1999 1759 2000 1763
rect 2004 1759 2005 1763
rect 1999 1758 2005 1759
rect 1679 1748 1818 1750
rect 1830 1751 1836 1752
rect 1679 1747 1680 1748
rect 1674 1746 1680 1747
rect 1830 1747 1831 1751
rect 1835 1750 1836 1751
rect 1999 1750 2001 1758
rect 1835 1748 2001 1750
rect 1835 1747 1836 1748
rect 1830 1746 1836 1747
rect 1202 1739 1208 1740
rect 1202 1738 1203 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 1088 1736 1203 1738
rect 110 1731 116 1732
rect 431 1731 437 1732
rect 431 1727 432 1731
rect 436 1730 437 1731
rect 458 1731 464 1732
rect 458 1730 459 1731
rect 436 1728 459 1730
rect 436 1727 437 1728
rect 431 1726 437 1727
rect 458 1727 459 1728
rect 463 1727 464 1731
rect 458 1726 464 1727
rect 471 1731 477 1732
rect 471 1727 472 1731
rect 476 1730 477 1731
rect 498 1731 504 1732
rect 498 1730 499 1731
rect 476 1728 499 1730
rect 476 1727 477 1728
rect 471 1726 477 1727
rect 498 1727 499 1728
rect 503 1727 504 1731
rect 498 1726 504 1727
rect 511 1731 517 1732
rect 511 1727 512 1731
rect 516 1730 517 1731
rect 538 1731 544 1732
rect 538 1730 539 1731
rect 516 1728 539 1730
rect 516 1727 517 1728
rect 511 1726 517 1727
rect 538 1727 539 1728
rect 543 1727 544 1731
rect 538 1726 544 1727
rect 551 1731 557 1732
rect 551 1727 552 1731
rect 556 1730 557 1731
rect 578 1731 584 1732
rect 578 1730 579 1731
rect 556 1728 579 1730
rect 556 1727 557 1728
rect 551 1726 557 1727
rect 578 1727 579 1728
rect 583 1727 584 1731
rect 578 1726 584 1727
rect 591 1731 597 1732
rect 591 1727 592 1731
rect 596 1730 597 1731
rect 618 1731 624 1732
rect 618 1730 619 1731
rect 596 1728 619 1730
rect 596 1727 597 1728
rect 591 1726 597 1727
rect 618 1727 619 1728
rect 623 1727 624 1731
rect 618 1726 624 1727
rect 631 1731 637 1732
rect 631 1727 632 1731
rect 636 1730 637 1731
rect 658 1731 664 1732
rect 658 1730 659 1731
rect 636 1728 659 1730
rect 636 1727 637 1728
rect 631 1726 637 1727
rect 658 1727 659 1728
rect 663 1727 664 1731
rect 658 1726 664 1727
rect 671 1731 680 1732
rect 671 1727 672 1731
rect 679 1727 680 1731
rect 671 1726 680 1727
rect 702 1731 708 1732
rect 702 1727 703 1731
rect 707 1730 708 1731
rect 719 1731 725 1732
rect 719 1730 720 1731
rect 707 1728 720 1730
rect 707 1727 708 1728
rect 702 1726 708 1727
rect 719 1727 720 1728
rect 724 1727 725 1731
rect 719 1726 725 1727
rect 742 1731 748 1732
rect 742 1727 743 1731
rect 747 1730 748 1731
rect 775 1731 781 1732
rect 775 1730 776 1731
rect 747 1728 776 1730
rect 747 1727 748 1728
rect 742 1726 748 1727
rect 775 1727 776 1728
rect 780 1727 781 1731
rect 775 1726 781 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1730 804 1731
rect 831 1731 837 1732
rect 831 1730 832 1731
rect 803 1728 832 1730
rect 803 1727 804 1728
rect 798 1726 804 1727
rect 831 1727 832 1728
rect 836 1727 837 1731
rect 831 1726 837 1727
rect 862 1731 868 1732
rect 862 1727 863 1731
rect 867 1730 868 1731
rect 895 1731 901 1732
rect 895 1730 896 1731
rect 867 1728 896 1730
rect 867 1727 868 1728
rect 862 1726 868 1727
rect 895 1727 896 1728
rect 900 1727 901 1731
rect 895 1726 901 1727
rect 926 1731 932 1732
rect 926 1727 927 1731
rect 931 1730 932 1731
rect 959 1731 965 1732
rect 959 1730 960 1731
rect 931 1728 960 1730
rect 931 1727 932 1728
rect 926 1726 932 1727
rect 959 1727 960 1728
rect 964 1727 965 1731
rect 959 1726 965 1727
rect 1023 1731 1029 1732
rect 1023 1727 1024 1731
rect 1028 1730 1029 1731
rect 1088 1730 1090 1736
rect 1202 1735 1203 1736
rect 1207 1735 1208 1739
rect 1602 1739 1608 1740
rect 1602 1738 1603 1739
rect 1202 1734 1208 1735
rect 1238 1736 1244 1737
rect 1238 1732 1239 1736
rect 1243 1732 1244 1736
rect 1028 1728 1090 1730
rect 1094 1731 1101 1732
rect 1028 1727 1029 1728
rect 1023 1726 1029 1727
rect 1094 1727 1095 1731
rect 1100 1727 1101 1731
rect 1094 1726 1101 1727
rect 1126 1731 1132 1732
rect 1126 1727 1127 1731
rect 1131 1730 1132 1731
rect 1167 1731 1173 1732
rect 1167 1730 1168 1731
rect 1131 1728 1168 1730
rect 1131 1727 1132 1728
rect 1126 1726 1132 1727
rect 1167 1727 1168 1728
rect 1172 1727 1173 1731
rect 1167 1726 1173 1727
rect 1215 1731 1221 1732
rect 1238 1731 1244 1732
rect 1278 1736 1284 1737
rect 1278 1732 1279 1736
rect 1283 1732 1284 1736
rect 1440 1736 1603 1738
rect 1278 1731 1284 1732
rect 1327 1731 1333 1732
rect 1215 1727 1216 1731
rect 1220 1727 1221 1731
rect 1215 1726 1221 1727
rect 1314 1727 1320 1728
rect 1314 1726 1315 1727
rect 1217 1724 1315 1726
rect 1314 1723 1315 1724
rect 1319 1723 1320 1727
rect 1327 1727 1328 1731
rect 1332 1730 1333 1731
rect 1354 1731 1360 1732
rect 1354 1730 1355 1731
rect 1332 1728 1355 1730
rect 1332 1727 1333 1728
rect 1327 1726 1333 1727
rect 1354 1727 1355 1728
rect 1359 1727 1360 1731
rect 1354 1726 1360 1727
rect 1366 1731 1373 1732
rect 1366 1727 1367 1731
rect 1372 1727 1373 1731
rect 1366 1726 1373 1727
rect 1415 1731 1421 1732
rect 1415 1727 1416 1731
rect 1420 1730 1421 1731
rect 1440 1730 1442 1736
rect 1602 1735 1603 1736
rect 1607 1735 1608 1739
rect 1602 1734 1608 1735
rect 1798 1739 1804 1740
rect 1798 1735 1799 1739
rect 1803 1738 1804 1739
rect 1803 1736 1842 1738
rect 1803 1735 1804 1736
rect 1798 1734 1804 1735
rect 1420 1728 1442 1730
rect 1446 1731 1452 1732
rect 1420 1727 1421 1728
rect 1415 1726 1421 1727
rect 1446 1727 1447 1731
rect 1451 1730 1452 1731
rect 1479 1731 1485 1732
rect 1479 1730 1480 1731
rect 1451 1728 1480 1730
rect 1451 1727 1452 1728
rect 1446 1726 1452 1727
rect 1479 1727 1480 1728
rect 1484 1727 1485 1731
rect 1479 1726 1485 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1730 1516 1731
rect 1543 1731 1549 1732
rect 1543 1730 1544 1731
rect 1515 1728 1544 1730
rect 1515 1727 1516 1728
rect 1510 1726 1516 1727
rect 1543 1727 1544 1728
rect 1548 1727 1549 1731
rect 1543 1726 1549 1727
rect 1574 1731 1580 1732
rect 1574 1727 1575 1731
rect 1579 1730 1580 1731
rect 1607 1731 1613 1732
rect 1607 1730 1608 1731
rect 1579 1728 1608 1730
rect 1579 1727 1580 1728
rect 1574 1726 1580 1727
rect 1607 1727 1608 1728
rect 1612 1727 1613 1731
rect 1607 1726 1613 1727
rect 1671 1731 1680 1732
rect 1671 1727 1672 1731
rect 1679 1727 1680 1731
rect 1671 1726 1680 1727
rect 1694 1731 1700 1732
rect 1694 1727 1695 1731
rect 1699 1730 1700 1731
rect 1727 1731 1733 1732
rect 1727 1730 1728 1731
rect 1699 1728 1728 1730
rect 1699 1727 1700 1728
rect 1694 1726 1700 1727
rect 1727 1727 1728 1728
rect 1732 1727 1733 1731
rect 1727 1726 1733 1727
rect 1750 1731 1756 1732
rect 1750 1727 1751 1731
rect 1755 1730 1756 1731
rect 1783 1731 1789 1732
rect 1783 1730 1784 1731
rect 1755 1728 1784 1730
rect 1755 1727 1756 1728
rect 1750 1726 1756 1727
rect 1783 1727 1784 1728
rect 1788 1727 1789 1731
rect 1783 1726 1789 1727
rect 1830 1731 1837 1732
rect 1830 1727 1831 1731
rect 1836 1727 1837 1731
rect 1840 1730 1842 1736
rect 2406 1736 2412 1737
rect 2406 1732 2407 1736
rect 2411 1732 2412 1736
rect 1887 1731 1893 1732
rect 1887 1730 1888 1731
rect 1840 1728 1888 1730
rect 1830 1726 1837 1727
rect 1887 1727 1888 1728
rect 1892 1727 1893 1731
rect 1887 1726 1893 1727
rect 1895 1731 1901 1732
rect 1895 1727 1896 1731
rect 1900 1730 1901 1731
rect 1943 1731 1949 1732
rect 1943 1730 1944 1731
rect 1900 1728 1944 1730
rect 1900 1727 1901 1728
rect 1895 1726 1901 1727
rect 1943 1727 1944 1728
rect 1948 1727 1949 1731
rect 1943 1726 1949 1727
rect 1966 1731 1972 1732
rect 1966 1727 1967 1731
rect 1971 1730 1972 1731
rect 1999 1731 2005 1732
rect 2406 1731 2412 1732
rect 1999 1730 2000 1731
rect 1971 1728 2000 1730
rect 1971 1727 1972 1728
rect 1966 1726 1972 1727
rect 1999 1727 2000 1728
rect 2004 1727 2005 1731
rect 1999 1726 2005 1727
rect 1314 1722 1320 1723
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 110 1714 116 1715
rect 1238 1719 1244 1720
rect 1238 1715 1239 1719
rect 1243 1715 1244 1719
rect 1238 1714 1244 1715
rect 1278 1719 1284 1720
rect 1278 1715 1279 1719
rect 1283 1715 1284 1719
rect 1278 1714 1284 1715
rect 2406 1719 2412 1720
rect 2406 1715 2407 1719
rect 2411 1715 2412 1719
rect 2406 1714 2412 1715
rect 406 1712 412 1713
rect 406 1708 407 1712
rect 411 1708 412 1712
rect 406 1707 412 1708
rect 446 1712 452 1713
rect 446 1708 447 1712
rect 451 1708 452 1712
rect 446 1707 452 1708
rect 486 1712 492 1713
rect 486 1708 487 1712
rect 491 1708 492 1712
rect 486 1707 492 1708
rect 526 1712 532 1713
rect 526 1708 527 1712
rect 531 1708 532 1712
rect 526 1707 532 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 606 1712 612 1713
rect 606 1708 607 1712
rect 611 1708 612 1712
rect 606 1707 612 1708
rect 646 1712 652 1713
rect 646 1708 647 1712
rect 651 1708 652 1712
rect 646 1707 652 1708
rect 694 1712 700 1713
rect 694 1708 695 1712
rect 699 1708 700 1712
rect 694 1707 700 1708
rect 750 1712 756 1713
rect 750 1708 751 1712
rect 755 1708 756 1712
rect 750 1707 756 1708
rect 806 1712 812 1713
rect 806 1708 807 1712
rect 811 1708 812 1712
rect 806 1707 812 1708
rect 870 1712 876 1713
rect 870 1708 871 1712
rect 875 1708 876 1712
rect 870 1707 876 1708
rect 934 1712 940 1713
rect 934 1708 935 1712
rect 939 1708 940 1712
rect 934 1707 940 1708
rect 998 1712 1004 1713
rect 998 1708 999 1712
rect 1003 1708 1004 1712
rect 998 1707 1004 1708
rect 1070 1712 1076 1713
rect 1070 1708 1071 1712
rect 1075 1708 1076 1712
rect 1070 1707 1076 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1190 1712 1196 1713
rect 1190 1708 1191 1712
rect 1195 1708 1196 1712
rect 1190 1707 1196 1708
rect 1302 1712 1308 1713
rect 1302 1708 1303 1712
rect 1307 1708 1308 1712
rect 1302 1707 1308 1708
rect 1342 1712 1348 1713
rect 1342 1708 1343 1712
rect 1347 1708 1348 1712
rect 1342 1707 1348 1708
rect 1390 1712 1396 1713
rect 1390 1708 1391 1712
rect 1395 1708 1396 1712
rect 1390 1707 1396 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1518 1712 1524 1713
rect 1518 1708 1519 1712
rect 1523 1708 1524 1712
rect 1518 1707 1524 1708
rect 1582 1712 1588 1713
rect 1582 1708 1583 1712
rect 1587 1708 1588 1712
rect 1582 1707 1588 1708
rect 1646 1712 1652 1713
rect 1646 1708 1647 1712
rect 1651 1708 1652 1712
rect 1646 1707 1652 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 1702 1707 1708 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1806 1712 1812 1713
rect 1806 1708 1807 1712
rect 1811 1708 1812 1712
rect 1806 1707 1812 1708
rect 1862 1712 1868 1713
rect 1862 1708 1863 1712
rect 1867 1708 1868 1712
rect 1862 1707 1868 1708
rect 1918 1712 1924 1713
rect 1918 1708 1919 1712
rect 1923 1708 1924 1712
rect 1918 1707 1924 1708
rect 1974 1712 1980 1713
rect 1974 1708 1975 1712
rect 1979 1708 1980 1712
rect 1974 1707 1980 1708
rect 278 1696 284 1697
rect 278 1692 279 1696
rect 283 1692 284 1696
rect 278 1691 284 1692
rect 318 1696 324 1697
rect 318 1692 319 1696
rect 323 1692 324 1696
rect 318 1691 324 1692
rect 358 1696 364 1697
rect 358 1692 359 1696
rect 363 1692 364 1696
rect 358 1691 364 1692
rect 398 1696 404 1697
rect 398 1692 399 1696
rect 403 1692 404 1696
rect 398 1691 404 1692
rect 446 1696 452 1697
rect 446 1692 447 1696
rect 451 1692 452 1696
rect 446 1691 452 1692
rect 494 1696 500 1697
rect 494 1692 495 1696
rect 499 1692 500 1696
rect 494 1691 500 1692
rect 542 1696 548 1697
rect 542 1692 543 1696
rect 547 1692 548 1696
rect 542 1691 548 1692
rect 590 1696 596 1697
rect 590 1692 591 1696
rect 595 1692 596 1696
rect 590 1691 596 1692
rect 638 1696 644 1697
rect 638 1692 639 1696
rect 643 1692 644 1696
rect 638 1691 644 1692
rect 686 1696 692 1697
rect 686 1692 687 1696
rect 691 1692 692 1696
rect 686 1691 692 1692
rect 734 1696 740 1697
rect 734 1692 735 1696
rect 739 1692 740 1696
rect 734 1691 740 1692
rect 782 1696 788 1697
rect 782 1692 783 1696
rect 787 1692 788 1696
rect 782 1691 788 1692
rect 838 1696 844 1697
rect 838 1692 839 1696
rect 843 1692 844 1696
rect 838 1691 844 1692
rect 894 1696 900 1697
rect 894 1692 895 1696
rect 899 1692 900 1696
rect 894 1691 900 1692
rect 1302 1696 1308 1697
rect 1302 1692 1303 1696
rect 1307 1692 1308 1696
rect 1302 1691 1308 1692
rect 1342 1696 1348 1697
rect 1342 1692 1343 1696
rect 1347 1692 1348 1696
rect 1342 1691 1348 1692
rect 1382 1696 1388 1697
rect 1382 1692 1383 1696
rect 1387 1692 1388 1696
rect 1382 1691 1388 1692
rect 1422 1696 1428 1697
rect 1422 1692 1423 1696
rect 1427 1692 1428 1696
rect 1422 1691 1428 1692
rect 1462 1696 1468 1697
rect 1462 1692 1463 1696
rect 1467 1692 1468 1696
rect 1462 1691 1468 1692
rect 1502 1696 1508 1697
rect 1502 1692 1503 1696
rect 1507 1692 1508 1696
rect 1502 1691 1508 1692
rect 1558 1696 1564 1697
rect 1558 1692 1559 1696
rect 1563 1692 1564 1696
rect 1558 1691 1564 1692
rect 1622 1696 1628 1697
rect 1622 1692 1623 1696
rect 1627 1692 1628 1696
rect 1622 1691 1628 1692
rect 1686 1696 1692 1697
rect 1686 1692 1687 1696
rect 1691 1692 1692 1696
rect 1686 1691 1692 1692
rect 1750 1696 1756 1697
rect 1750 1692 1751 1696
rect 1755 1692 1756 1696
rect 1750 1691 1756 1692
rect 1806 1696 1812 1697
rect 1806 1692 1807 1696
rect 1811 1692 1812 1696
rect 1806 1691 1812 1692
rect 1862 1696 1868 1697
rect 1862 1692 1863 1696
rect 1867 1692 1868 1696
rect 1862 1691 1868 1692
rect 1918 1696 1924 1697
rect 1918 1692 1919 1696
rect 1923 1692 1924 1696
rect 1918 1691 1924 1692
rect 1974 1696 1980 1697
rect 1974 1692 1975 1696
rect 1979 1692 1980 1696
rect 1974 1691 1980 1692
rect 2030 1696 2036 1697
rect 2030 1692 2031 1696
rect 2035 1692 2036 1696
rect 2030 1691 2036 1692
rect 2086 1696 2092 1697
rect 2086 1692 2087 1696
rect 2091 1692 2092 1696
rect 2086 1691 2092 1692
rect 110 1689 116 1690
rect 110 1685 111 1689
rect 115 1685 116 1689
rect 110 1684 116 1685
rect 1238 1689 1244 1690
rect 1238 1685 1239 1689
rect 1243 1685 1244 1689
rect 1238 1684 1244 1685
rect 1278 1689 1284 1690
rect 1278 1685 1279 1689
rect 1283 1685 1284 1689
rect 1278 1684 1284 1685
rect 2406 1689 2412 1690
rect 2406 1685 2407 1689
rect 2411 1685 2412 1689
rect 2406 1684 2412 1685
rect 566 1683 572 1684
rect 566 1682 567 1683
rect 428 1680 567 1682
rect 428 1676 430 1680
rect 566 1679 567 1680
rect 571 1679 572 1683
rect 1594 1683 1600 1684
rect 1594 1682 1595 1683
rect 566 1678 572 1679
rect 1528 1680 1595 1682
rect 1528 1676 1530 1680
rect 1594 1679 1595 1680
rect 1599 1679 1600 1683
rect 2110 1683 2116 1684
rect 2110 1682 2111 1683
rect 1594 1678 1600 1679
rect 1948 1680 2111 1682
rect 1948 1676 1950 1680
rect 2110 1679 2111 1680
rect 2115 1679 2116 1683
rect 2110 1678 2116 1679
rect 303 1675 309 1676
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 303 1671 304 1675
rect 308 1674 309 1675
rect 330 1675 336 1676
rect 308 1672 321 1674
rect 308 1671 309 1672
rect 303 1670 309 1671
rect 110 1667 116 1668
rect 319 1666 321 1672
rect 330 1671 331 1675
rect 335 1674 336 1675
rect 343 1675 349 1676
rect 343 1674 344 1675
rect 335 1672 344 1674
rect 335 1671 336 1672
rect 330 1670 336 1671
rect 343 1671 344 1672
rect 348 1671 349 1675
rect 343 1670 349 1671
rect 366 1675 372 1676
rect 366 1671 367 1675
rect 371 1674 372 1675
rect 383 1675 389 1676
rect 383 1674 384 1675
rect 371 1672 384 1674
rect 371 1671 372 1672
rect 366 1670 372 1671
rect 383 1671 384 1672
rect 388 1671 389 1675
rect 383 1670 389 1671
rect 423 1675 430 1676
rect 423 1671 424 1675
rect 428 1672 430 1675
rect 434 1675 440 1676
rect 428 1671 429 1672
rect 423 1670 429 1671
rect 434 1671 435 1675
rect 439 1674 440 1675
rect 471 1675 477 1676
rect 471 1674 472 1675
rect 439 1672 472 1674
rect 439 1671 440 1672
rect 434 1670 440 1671
rect 471 1671 472 1672
rect 476 1671 477 1675
rect 471 1670 477 1671
rect 479 1675 485 1676
rect 479 1671 480 1675
rect 484 1674 485 1675
rect 519 1675 525 1676
rect 519 1674 520 1675
rect 484 1672 520 1674
rect 484 1671 485 1672
rect 479 1670 485 1671
rect 519 1671 520 1672
rect 524 1671 525 1675
rect 519 1670 525 1671
rect 527 1675 533 1676
rect 527 1671 528 1675
rect 532 1674 533 1675
rect 567 1675 573 1676
rect 567 1674 568 1675
rect 532 1672 568 1674
rect 532 1671 533 1672
rect 527 1670 533 1671
rect 567 1671 568 1672
rect 572 1671 573 1675
rect 567 1670 573 1671
rect 615 1675 621 1676
rect 615 1671 616 1675
rect 620 1671 621 1675
rect 615 1670 621 1671
rect 623 1675 629 1676
rect 623 1671 624 1675
rect 628 1674 629 1675
rect 663 1675 669 1676
rect 663 1674 664 1675
rect 628 1672 664 1674
rect 628 1671 629 1672
rect 623 1670 629 1671
rect 663 1671 664 1672
rect 668 1671 669 1675
rect 663 1670 669 1671
rect 711 1675 717 1676
rect 711 1671 712 1675
rect 716 1674 717 1675
rect 750 1675 756 1676
rect 750 1674 751 1675
rect 716 1672 751 1674
rect 716 1671 717 1672
rect 711 1670 717 1671
rect 750 1671 751 1672
rect 755 1671 756 1675
rect 750 1670 756 1671
rect 759 1675 765 1676
rect 759 1671 760 1675
rect 764 1674 765 1675
rect 798 1675 804 1676
rect 798 1674 799 1675
rect 764 1672 799 1674
rect 764 1671 765 1672
rect 759 1670 765 1671
rect 798 1671 799 1672
rect 803 1671 804 1675
rect 798 1670 804 1671
rect 807 1675 813 1676
rect 807 1671 808 1675
rect 812 1674 813 1675
rect 818 1675 824 1676
rect 812 1671 814 1674
rect 807 1670 814 1671
rect 818 1671 819 1675
rect 823 1674 824 1675
rect 863 1675 869 1676
rect 863 1674 864 1675
rect 823 1672 864 1674
rect 823 1671 824 1672
rect 818 1670 824 1671
rect 863 1671 864 1672
rect 868 1671 869 1675
rect 863 1670 869 1671
rect 871 1675 877 1676
rect 871 1671 872 1675
rect 876 1674 877 1675
rect 919 1675 925 1676
rect 919 1674 920 1675
rect 876 1672 920 1674
rect 876 1671 877 1672
rect 871 1670 877 1671
rect 919 1671 920 1672
rect 924 1671 925 1675
rect 1327 1675 1333 1676
rect 919 1670 925 1671
rect 1238 1672 1244 1673
rect 422 1667 428 1668
rect 422 1666 423 1667
rect 319 1664 423 1666
rect 422 1663 423 1664
rect 427 1663 428 1667
rect 616 1666 618 1670
rect 710 1667 716 1668
rect 710 1666 711 1667
rect 616 1664 711 1666
rect 422 1662 428 1663
rect 710 1663 711 1664
rect 715 1663 716 1667
rect 812 1666 814 1670
rect 1238 1668 1239 1672
rect 1243 1668 1244 1672
rect 918 1667 924 1668
rect 1238 1667 1244 1668
rect 1278 1672 1284 1673
rect 1278 1668 1279 1672
rect 1283 1668 1284 1672
rect 1327 1671 1328 1675
rect 1332 1674 1333 1675
rect 1350 1675 1356 1676
rect 1332 1672 1346 1674
rect 1332 1671 1333 1672
rect 1327 1670 1333 1671
rect 1278 1667 1284 1668
rect 918 1666 919 1667
rect 812 1664 919 1666
rect 710 1662 716 1663
rect 918 1663 919 1664
rect 923 1663 924 1667
rect 1344 1666 1346 1672
rect 1350 1671 1351 1675
rect 1355 1674 1356 1675
rect 1367 1675 1373 1676
rect 1367 1674 1368 1675
rect 1355 1672 1368 1674
rect 1355 1671 1356 1672
rect 1350 1670 1356 1671
rect 1367 1671 1368 1672
rect 1372 1671 1373 1675
rect 1367 1670 1373 1671
rect 1407 1675 1413 1676
rect 1407 1671 1408 1675
rect 1412 1674 1413 1675
rect 1430 1675 1436 1676
rect 1412 1672 1426 1674
rect 1412 1671 1413 1672
rect 1407 1670 1413 1671
rect 1406 1667 1412 1668
rect 1406 1666 1407 1667
rect 1344 1664 1407 1666
rect 918 1662 924 1663
rect 1406 1663 1407 1664
rect 1411 1663 1412 1667
rect 1424 1666 1426 1672
rect 1430 1671 1431 1675
rect 1435 1674 1436 1675
rect 1447 1675 1453 1676
rect 1447 1674 1448 1675
rect 1435 1672 1448 1674
rect 1435 1671 1436 1672
rect 1430 1670 1436 1671
rect 1447 1671 1448 1672
rect 1452 1671 1453 1675
rect 1447 1670 1453 1671
rect 1470 1675 1476 1676
rect 1470 1671 1471 1675
rect 1475 1674 1476 1675
rect 1487 1675 1493 1676
rect 1487 1674 1488 1675
rect 1475 1672 1488 1674
rect 1475 1671 1476 1672
rect 1470 1670 1476 1671
rect 1487 1671 1488 1672
rect 1492 1671 1493 1675
rect 1487 1670 1493 1671
rect 1527 1675 1533 1676
rect 1527 1671 1528 1675
rect 1532 1671 1533 1675
rect 1527 1670 1533 1671
rect 1535 1675 1541 1676
rect 1535 1671 1536 1675
rect 1540 1674 1541 1675
rect 1583 1675 1589 1676
rect 1583 1674 1584 1675
rect 1540 1672 1584 1674
rect 1540 1671 1541 1672
rect 1535 1670 1541 1671
rect 1583 1671 1584 1672
rect 1588 1671 1589 1675
rect 1583 1670 1589 1671
rect 1591 1675 1597 1676
rect 1591 1671 1592 1675
rect 1596 1674 1597 1675
rect 1647 1675 1653 1676
rect 1647 1674 1648 1675
rect 1596 1672 1648 1674
rect 1596 1671 1597 1672
rect 1591 1670 1597 1671
rect 1647 1671 1648 1672
rect 1652 1671 1653 1675
rect 1647 1670 1653 1671
rect 1655 1675 1661 1676
rect 1655 1671 1656 1675
rect 1660 1674 1661 1675
rect 1711 1675 1717 1676
rect 1711 1674 1712 1675
rect 1660 1672 1712 1674
rect 1660 1671 1661 1672
rect 1655 1670 1661 1671
rect 1711 1671 1712 1672
rect 1716 1671 1717 1675
rect 1711 1670 1717 1671
rect 1775 1675 1781 1676
rect 1775 1671 1776 1675
rect 1780 1674 1781 1675
rect 1786 1675 1792 1676
rect 1780 1671 1782 1674
rect 1775 1670 1782 1671
rect 1786 1671 1787 1675
rect 1791 1674 1792 1675
rect 1831 1675 1837 1676
rect 1831 1674 1832 1675
rect 1791 1672 1832 1674
rect 1791 1671 1792 1672
rect 1786 1670 1792 1671
rect 1831 1671 1832 1672
rect 1836 1671 1837 1675
rect 1831 1670 1837 1671
rect 1839 1675 1845 1676
rect 1839 1671 1840 1675
rect 1844 1674 1845 1675
rect 1887 1675 1893 1676
rect 1887 1674 1888 1675
rect 1844 1672 1888 1674
rect 1844 1671 1845 1672
rect 1839 1670 1845 1671
rect 1887 1671 1888 1672
rect 1892 1671 1893 1675
rect 1887 1670 1893 1671
rect 1943 1675 1950 1676
rect 1943 1671 1944 1675
rect 1948 1672 1950 1675
rect 1954 1675 1960 1676
rect 1948 1671 1949 1672
rect 1943 1670 1949 1671
rect 1954 1671 1955 1675
rect 1959 1674 1960 1675
rect 1999 1675 2005 1676
rect 1999 1674 2000 1675
rect 1959 1672 2000 1674
rect 1959 1671 1960 1672
rect 1954 1670 1960 1671
rect 1999 1671 2000 1672
rect 2004 1671 2005 1675
rect 1999 1670 2005 1671
rect 2007 1675 2013 1676
rect 2007 1671 2008 1675
rect 2012 1674 2013 1675
rect 2055 1675 2061 1676
rect 2055 1674 2056 1675
rect 2012 1672 2056 1674
rect 2012 1671 2013 1672
rect 2007 1670 2013 1671
rect 2055 1671 2056 1672
rect 2060 1671 2061 1675
rect 2055 1670 2061 1671
rect 2063 1675 2069 1676
rect 2063 1671 2064 1675
rect 2068 1674 2069 1675
rect 2111 1675 2117 1676
rect 2111 1674 2112 1675
rect 2068 1672 2112 1674
rect 2068 1671 2069 1672
rect 2063 1670 2069 1671
rect 2111 1671 2112 1672
rect 2116 1671 2117 1675
rect 2111 1670 2117 1671
rect 2406 1672 2412 1673
rect 1486 1667 1492 1668
rect 1486 1666 1487 1667
rect 1424 1664 1487 1666
rect 1406 1662 1412 1663
rect 1486 1663 1487 1664
rect 1491 1663 1492 1667
rect 1780 1666 1782 1670
rect 2406 1668 2407 1672
rect 2411 1668 2412 1672
rect 1942 1667 1948 1668
rect 2406 1667 2412 1668
rect 1942 1666 1943 1667
rect 1780 1664 1943 1666
rect 1486 1662 1492 1663
rect 1942 1663 1943 1664
rect 1947 1663 1948 1667
rect 1942 1662 1948 1663
rect 278 1649 284 1650
rect 278 1645 279 1649
rect 283 1645 284 1649
rect 278 1644 284 1645
rect 318 1649 324 1650
rect 318 1645 319 1649
rect 323 1645 324 1649
rect 318 1644 324 1645
rect 358 1649 364 1650
rect 358 1645 359 1649
rect 363 1645 364 1649
rect 358 1644 364 1645
rect 398 1649 404 1650
rect 398 1645 399 1649
rect 403 1645 404 1649
rect 398 1644 404 1645
rect 446 1649 452 1650
rect 446 1645 447 1649
rect 451 1645 452 1649
rect 446 1644 452 1645
rect 494 1649 500 1650
rect 494 1645 495 1649
rect 499 1645 500 1649
rect 494 1644 500 1645
rect 542 1649 548 1650
rect 542 1645 543 1649
rect 547 1645 548 1649
rect 542 1644 548 1645
rect 590 1649 596 1650
rect 590 1645 591 1649
rect 595 1645 596 1649
rect 590 1644 596 1645
rect 638 1649 644 1650
rect 638 1645 639 1649
rect 643 1645 644 1649
rect 638 1644 644 1645
rect 686 1649 692 1650
rect 686 1645 687 1649
rect 691 1645 692 1649
rect 686 1644 692 1645
rect 734 1649 740 1650
rect 734 1645 735 1649
rect 739 1645 740 1649
rect 734 1644 740 1645
rect 782 1649 788 1650
rect 782 1645 783 1649
rect 787 1645 788 1649
rect 782 1644 788 1645
rect 838 1649 844 1650
rect 838 1645 839 1649
rect 843 1645 844 1649
rect 838 1644 844 1645
rect 894 1649 900 1650
rect 894 1645 895 1649
rect 899 1645 900 1649
rect 894 1644 900 1645
rect 1302 1649 1308 1650
rect 1302 1645 1303 1649
rect 1307 1645 1308 1649
rect 1302 1644 1308 1645
rect 1342 1649 1348 1650
rect 1342 1645 1343 1649
rect 1347 1645 1348 1649
rect 1342 1644 1348 1645
rect 1382 1649 1388 1650
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1422 1649 1428 1650
rect 1422 1645 1423 1649
rect 1427 1645 1428 1649
rect 1422 1644 1428 1645
rect 1462 1649 1468 1650
rect 1462 1645 1463 1649
rect 1467 1645 1468 1649
rect 1462 1644 1468 1645
rect 1502 1649 1508 1650
rect 1502 1645 1503 1649
rect 1507 1645 1508 1649
rect 1502 1644 1508 1645
rect 1558 1649 1564 1650
rect 1558 1645 1559 1649
rect 1563 1645 1564 1649
rect 1558 1644 1564 1645
rect 1622 1649 1628 1650
rect 1622 1645 1623 1649
rect 1627 1645 1628 1649
rect 1622 1644 1628 1645
rect 1686 1649 1692 1650
rect 1686 1645 1687 1649
rect 1691 1645 1692 1649
rect 1686 1644 1692 1645
rect 1750 1649 1756 1650
rect 1750 1645 1751 1649
rect 1755 1645 1756 1649
rect 1750 1644 1756 1645
rect 1806 1649 1812 1650
rect 1806 1645 1807 1649
rect 1811 1645 1812 1649
rect 1806 1644 1812 1645
rect 1862 1649 1868 1650
rect 1862 1645 1863 1649
rect 1867 1645 1868 1649
rect 1862 1644 1868 1645
rect 1918 1649 1924 1650
rect 1918 1645 1919 1649
rect 1923 1645 1924 1649
rect 1918 1644 1924 1645
rect 1974 1649 1980 1650
rect 1974 1645 1975 1649
rect 1979 1645 1980 1649
rect 1974 1644 1980 1645
rect 2030 1649 2036 1650
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2030 1644 2036 1645
rect 2086 1649 2092 1650
rect 2086 1645 2087 1649
rect 2091 1645 2092 1649
rect 2086 1644 2092 1645
rect 303 1643 309 1644
rect 303 1639 304 1643
rect 308 1642 309 1643
rect 330 1643 336 1644
rect 330 1642 331 1643
rect 308 1640 331 1642
rect 308 1639 309 1640
rect 303 1638 309 1639
rect 330 1639 331 1640
rect 335 1639 336 1643
rect 330 1638 336 1639
rect 343 1643 349 1644
rect 343 1639 344 1643
rect 348 1642 349 1643
rect 366 1643 372 1644
rect 366 1642 367 1643
rect 348 1640 367 1642
rect 348 1639 349 1640
rect 343 1638 349 1639
rect 366 1639 367 1640
rect 371 1639 372 1643
rect 366 1638 372 1639
rect 383 1643 389 1644
rect 383 1639 384 1643
rect 388 1642 389 1643
rect 406 1643 412 1644
rect 406 1642 407 1643
rect 388 1640 407 1642
rect 388 1639 389 1640
rect 383 1638 389 1639
rect 406 1639 407 1640
rect 411 1639 412 1643
rect 406 1638 412 1639
rect 422 1643 429 1644
rect 422 1639 423 1643
rect 428 1639 429 1643
rect 422 1638 429 1639
rect 471 1643 477 1644
rect 471 1639 472 1643
rect 476 1642 477 1643
rect 479 1643 485 1644
rect 479 1642 480 1643
rect 476 1640 480 1642
rect 476 1639 477 1640
rect 471 1638 477 1639
rect 479 1639 480 1640
rect 484 1639 485 1643
rect 479 1638 485 1639
rect 519 1643 525 1644
rect 519 1639 520 1643
rect 524 1642 525 1643
rect 527 1643 533 1644
rect 527 1642 528 1643
rect 524 1640 528 1642
rect 524 1639 525 1640
rect 519 1638 525 1639
rect 527 1639 528 1640
rect 532 1639 533 1643
rect 527 1638 533 1639
rect 566 1643 573 1644
rect 566 1639 567 1643
rect 572 1639 573 1643
rect 566 1638 573 1639
rect 615 1643 621 1644
rect 615 1639 616 1643
rect 620 1642 621 1643
rect 623 1643 629 1644
rect 623 1642 624 1643
rect 620 1640 624 1642
rect 620 1639 621 1640
rect 615 1638 621 1639
rect 623 1639 624 1640
rect 628 1639 629 1643
rect 623 1638 629 1639
rect 663 1643 669 1644
rect 663 1639 664 1643
rect 668 1642 669 1643
rect 702 1643 708 1644
rect 702 1642 703 1643
rect 668 1640 703 1642
rect 668 1639 669 1640
rect 663 1638 669 1639
rect 702 1639 703 1640
rect 707 1639 708 1643
rect 702 1638 708 1639
rect 710 1643 717 1644
rect 710 1639 711 1643
rect 716 1639 717 1643
rect 710 1638 717 1639
rect 750 1643 756 1644
rect 750 1639 751 1643
rect 755 1642 756 1643
rect 759 1643 765 1644
rect 759 1642 760 1643
rect 755 1640 760 1642
rect 755 1639 756 1640
rect 750 1638 756 1639
rect 759 1639 760 1640
rect 764 1639 765 1643
rect 759 1638 765 1639
rect 798 1643 804 1644
rect 798 1639 799 1643
rect 803 1642 804 1643
rect 807 1643 813 1644
rect 807 1642 808 1643
rect 803 1640 808 1642
rect 803 1639 804 1640
rect 798 1638 804 1639
rect 807 1639 808 1640
rect 812 1639 813 1643
rect 807 1638 813 1639
rect 863 1643 869 1644
rect 863 1639 864 1643
rect 868 1642 869 1643
rect 871 1643 877 1644
rect 871 1642 872 1643
rect 868 1640 872 1642
rect 868 1639 869 1640
rect 863 1638 869 1639
rect 871 1639 872 1640
rect 876 1639 877 1643
rect 871 1638 877 1639
rect 918 1643 925 1644
rect 918 1639 919 1643
rect 924 1639 925 1643
rect 918 1638 925 1639
rect 1327 1643 1333 1644
rect 1327 1639 1328 1643
rect 1332 1642 1333 1643
rect 1350 1643 1356 1644
rect 1350 1642 1351 1643
rect 1332 1640 1351 1642
rect 1332 1639 1333 1640
rect 1327 1638 1333 1639
rect 1350 1639 1351 1640
rect 1355 1639 1356 1643
rect 1350 1638 1356 1639
rect 1366 1643 1373 1644
rect 1366 1639 1367 1643
rect 1372 1639 1373 1643
rect 1366 1638 1373 1639
rect 1406 1643 1413 1644
rect 1406 1639 1407 1643
rect 1412 1639 1413 1643
rect 1406 1638 1413 1639
rect 1447 1643 1453 1644
rect 1447 1639 1448 1643
rect 1452 1642 1453 1643
rect 1470 1643 1476 1644
rect 1470 1642 1471 1643
rect 1452 1640 1471 1642
rect 1452 1639 1453 1640
rect 1447 1638 1453 1639
rect 1470 1639 1471 1640
rect 1475 1639 1476 1643
rect 1470 1638 1476 1639
rect 1486 1643 1493 1644
rect 1486 1639 1487 1643
rect 1492 1639 1493 1643
rect 1486 1638 1493 1639
rect 1527 1643 1533 1644
rect 1527 1639 1528 1643
rect 1532 1642 1533 1643
rect 1535 1643 1541 1644
rect 1535 1642 1536 1643
rect 1532 1640 1536 1642
rect 1532 1639 1533 1640
rect 1527 1638 1533 1639
rect 1535 1639 1536 1640
rect 1540 1639 1541 1643
rect 1535 1638 1541 1639
rect 1583 1643 1589 1644
rect 1583 1639 1584 1643
rect 1588 1642 1589 1643
rect 1591 1643 1597 1644
rect 1591 1642 1592 1643
rect 1588 1640 1592 1642
rect 1588 1639 1589 1640
rect 1583 1638 1589 1639
rect 1591 1639 1592 1640
rect 1596 1639 1597 1643
rect 1591 1638 1597 1639
rect 1647 1643 1653 1644
rect 1647 1639 1648 1643
rect 1652 1642 1653 1643
rect 1655 1643 1661 1644
rect 1655 1642 1656 1643
rect 1652 1640 1656 1642
rect 1652 1639 1653 1640
rect 1647 1638 1653 1639
rect 1655 1639 1656 1640
rect 1660 1639 1661 1643
rect 1655 1638 1661 1639
rect 1663 1643 1669 1644
rect 1663 1639 1664 1643
rect 1668 1642 1669 1643
rect 1711 1643 1717 1644
rect 1711 1642 1712 1643
rect 1668 1640 1712 1642
rect 1668 1639 1669 1640
rect 1663 1638 1669 1639
rect 1711 1639 1712 1640
rect 1716 1639 1717 1643
rect 1711 1638 1717 1639
rect 1775 1643 1781 1644
rect 1775 1639 1776 1643
rect 1780 1642 1781 1643
rect 1786 1643 1792 1644
rect 1786 1642 1787 1643
rect 1780 1640 1787 1642
rect 1780 1639 1781 1640
rect 1775 1638 1781 1639
rect 1786 1639 1787 1640
rect 1791 1639 1792 1643
rect 1786 1638 1792 1639
rect 1831 1643 1837 1644
rect 1831 1639 1832 1643
rect 1836 1642 1837 1643
rect 1839 1643 1845 1644
rect 1839 1642 1840 1643
rect 1836 1640 1840 1642
rect 1836 1639 1837 1640
rect 1831 1638 1837 1639
rect 1839 1639 1840 1640
rect 1844 1639 1845 1643
rect 1839 1638 1845 1639
rect 1887 1643 1893 1644
rect 1887 1639 1888 1643
rect 1892 1642 1893 1643
rect 1895 1643 1901 1644
rect 1895 1642 1896 1643
rect 1892 1640 1896 1642
rect 1892 1639 1893 1640
rect 1887 1638 1893 1639
rect 1895 1639 1896 1640
rect 1900 1639 1901 1643
rect 1895 1638 1901 1639
rect 1942 1643 1949 1644
rect 1942 1639 1943 1643
rect 1948 1639 1949 1643
rect 1942 1638 1949 1639
rect 1999 1643 2005 1644
rect 1999 1639 2000 1643
rect 2004 1642 2005 1643
rect 2007 1643 2013 1644
rect 2007 1642 2008 1643
rect 2004 1640 2008 1642
rect 2004 1639 2005 1640
rect 1999 1638 2005 1639
rect 2007 1639 2008 1640
rect 2012 1639 2013 1643
rect 2007 1638 2013 1639
rect 2055 1643 2061 1644
rect 2055 1639 2056 1643
rect 2060 1642 2061 1643
rect 2063 1643 2069 1644
rect 2063 1642 2064 1643
rect 2060 1640 2064 1642
rect 2060 1639 2061 1640
rect 2055 1638 2061 1639
rect 2063 1639 2064 1640
rect 2068 1639 2069 1643
rect 2063 1638 2069 1639
rect 2110 1643 2117 1644
rect 2110 1639 2111 1643
rect 2116 1639 2117 1643
rect 2110 1638 2117 1639
rect 1358 1623 1364 1624
rect 1358 1622 1359 1623
rect 1336 1620 1359 1622
rect 159 1619 168 1620
rect 134 1615 140 1616
rect 134 1611 135 1615
rect 139 1611 140 1615
rect 159 1615 160 1619
rect 167 1615 168 1619
rect 186 1619 192 1620
rect 159 1614 168 1615
rect 174 1615 180 1616
rect 134 1610 140 1611
rect 174 1611 175 1615
rect 179 1611 180 1615
rect 186 1615 187 1619
rect 191 1618 192 1619
rect 199 1619 205 1620
rect 199 1618 200 1619
rect 191 1616 200 1618
rect 191 1615 192 1616
rect 186 1614 192 1615
rect 199 1615 200 1616
rect 204 1615 205 1619
rect 239 1619 245 1620
rect 199 1614 205 1615
rect 214 1615 220 1616
rect 174 1610 180 1611
rect 214 1611 215 1615
rect 219 1611 220 1615
rect 239 1615 240 1619
rect 244 1615 245 1619
rect 266 1619 272 1620
rect 239 1614 245 1615
rect 254 1615 260 1616
rect 214 1610 220 1611
rect 167 1607 173 1608
rect 167 1603 168 1607
rect 172 1606 173 1607
rect 241 1606 243 1614
rect 254 1611 255 1615
rect 259 1611 260 1615
rect 266 1615 267 1619
rect 271 1618 272 1619
rect 279 1619 285 1620
rect 279 1618 280 1619
rect 271 1616 280 1618
rect 271 1615 272 1616
rect 266 1614 272 1615
rect 279 1615 280 1616
rect 284 1615 285 1619
rect 326 1619 332 1620
rect 279 1614 285 1615
rect 310 1615 316 1616
rect 254 1610 260 1611
rect 310 1611 311 1615
rect 315 1611 316 1615
rect 326 1615 327 1619
rect 331 1618 332 1619
rect 335 1619 341 1620
rect 335 1618 336 1619
rect 331 1616 336 1618
rect 331 1615 332 1616
rect 326 1614 332 1615
rect 335 1615 336 1616
rect 340 1615 341 1619
rect 415 1619 421 1620
rect 335 1614 341 1615
rect 390 1615 396 1616
rect 310 1610 316 1611
rect 390 1611 391 1615
rect 395 1611 396 1615
rect 415 1615 416 1619
rect 420 1618 421 1619
rect 462 1619 468 1620
rect 462 1618 463 1619
rect 420 1616 463 1618
rect 420 1615 421 1616
rect 415 1614 421 1615
rect 462 1615 463 1616
rect 467 1615 468 1619
rect 495 1619 501 1620
rect 462 1614 468 1615
rect 470 1615 476 1616
rect 390 1610 396 1611
rect 470 1611 471 1615
rect 475 1611 476 1615
rect 495 1615 496 1619
rect 500 1618 501 1619
rect 550 1619 556 1620
rect 550 1618 551 1619
rect 500 1616 551 1618
rect 500 1615 501 1616
rect 495 1614 501 1615
rect 550 1615 551 1616
rect 555 1615 556 1619
rect 570 1619 576 1620
rect 550 1614 556 1615
rect 558 1615 564 1616
rect 470 1610 476 1611
rect 558 1611 559 1615
rect 563 1611 564 1615
rect 570 1615 571 1619
rect 575 1618 576 1619
rect 583 1619 589 1620
rect 583 1618 584 1619
rect 575 1616 584 1618
rect 575 1615 576 1616
rect 570 1614 576 1615
rect 583 1615 584 1616
rect 588 1615 589 1619
rect 663 1619 669 1620
rect 583 1614 589 1615
rect 638 1615 644 1616
rect 558 1610 564 1611
rect 638 1611 639 1615
rect 643 1611 644 1615
rect 663 1615 664 1619
rect 668 1618 669 1619
rect 710 1619 716 1620
rect 710 1618 711 1619
rect 668 1616 711 1618
rect 668 1615 669 1616
rect 663 1614 669 1615
rect 710 1615 711 1616
rect 715 1615 716 1619
rect 743 1619 749 1620
rect 710 1614 716 1615
rect 718 1615 724 1616
rect 638 1610 644 1611
rect 718 1611 719 1615
rect 723 1611 724 1615
rect 743 1615 744 1619
rect 748 1618 749 1619
rect 782 1619 788 1620
rect 782 1618 783 1619
rect 748 1616 783 1618
rect 748 1615 749 1616
rect 743 1614 749 1615
rect 782 1615 783 1616
rect 787 1615 788 1619
rect 815 1619 824 1620
rect 782 1614 788 1615
rect 790 1615 796 1616
rect 718 1610 724 1611
rect 790 1611 791 1615
rect 795 1611 796 1615
rect 815 1615 816 1619
rect 823 1615 824 1619
rect 866 1619 872 1620
rect 815 1614 824 1615
rect 854 1615 860 1616
rect 790 1610 796 1611
rect 854 1611 855 1615
rect 859 1611 860 1615
rect 866 1615 867 1619
rect 871 1618 872 1619
rect 879 1619 885 1620
rect 879 1618 880 1619
rect 871 1616 880 1618
rect 871 1615 872 1616
rect 866 1614 872 1615
rect 879 1615 880 1616
rect 884 1615 885 1619
rect 943 1619 949 1620
rect 879 1614 885 1615
rect 918 1615 924 1616
rect 854 1610 860 1611
rect 918 1611 919 1615
rect 923 1611 924 1615
rect 943 1615 944 1619
rect 948 1618 949 1619
rect 974 1619 980 1620
rect 974 1618 975 1619
rect 948 1616 975 1618
rect 948 1615 949 1616
rect 943 1614 949 1615
rect 974 1615 975 1616
rect 979 1615 980 1619
rect 1007 1619 1013 1620
rect 974 1614 980 1615
rect 982 1615 988 1616
rect 918 1610 924 1611
rect 982 1611 983 1615
rect 987 1611 988 1615
rect 1007 1615 1008 1619
rect 1012 1618 1013 1619
rect 1038 1619 1044 1620
rect 1038 1618 1039 1619
rect 1012 1616 1039 1618
rect 1012 1615 1013 1616
rect 1007 1614 1013 1615
rect 1038 1615 1039 1616
rect 1043 1615 1044 1619
rect 1058 1619 1064 1620
rect 1038 1614 1044 1615
rect 1046 1615 1052 1616
rect 982 1610 988 1611
rect 1046 1611 1047 1615
rect 1051 1611 1052 1615
rect 1058 1615 1059 1619
rect 1063 1618 1064 1619
rect 1071 1619 1077 1620
rect 1071 1618 1072 1619
rect 1063 1616 1072 1618
rect 1063 1615 1064 1616
rect 1058 1614 1064 1615
rect 1071 1615 1072 1616
rect 1076 1615 1077 1619
rect 1327 1619 1333 1620
rect 1071 1614 1077 1615
rect 1302 1615 1308 1616
rect 1046 1610 1052 1611
rect 1302 1611 1303 1615
rect 1307 1611 1308 1615
rect 1327 1615 1328 1619
rect 1332 1618 1333 1619
rect 1336 1618 1338 1620
rect 1358 1619 1359 1620
rect 1363 1619 1364 1623
rect 1398 1623 1404 1624
rect 1398 1622 1399 1623
rect 1376 1620 1399 1622
rect 1358 1618 1364 1619
rect 1367 1619 1373 1620
rect 1332 1616 1338 1618
rect 1332 1615 1333 1616
rect 1327 1614 1333 1615
rect 1342 1615 1348 1616
rect 1302 1610 1308 1611
rect 1342 1611 1343 1615
rect 1347 1611 1348 1615
rect 1367 1615 1368 1619
rect 1372 1618 1373 1619
rect 1376 1618 1378 1620
rect 1398 1619 1399 1620
rect 1403 1619 1404 1623
rect 1430 1623 1436 1624
rect 1430 1622 1431 1623
rect 1398 1618 1404 1619
rect 1407 1621 1431 1622
rect 1372 1616 1378 1618
rect 1407 1617 1408 1621
rect 1412 1620 1431 1621
rect 1412 1617 1413 1620
rect 1430 1619 1431 1620
rect 1435 1619 1436 1623
rect 1430 1618 1436 1619
rect 1438 1619 1444 1620
rect 1407 1616 1413 1617
rect 1372 1615 1373 1616
rect 1367 1614 1373 1615
rect 1382 1615 1388 1616
rect 1342 1610 1348 1611
rect 1382 1611 1383 1615
rect 1387 1611 1388 1615
rect 1382 1610 1388 1611
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 1438 1615 1439 1619
rect 1443 1618 1444 1619
rect 1447 1619 1453 1620
rect 1447 1618 1448 1619
rect 1443 1616 1448 1618
rect 1443 1615 1444 1616
rect 1438 1614 1444 1615
rect 1447 1615 1448 1616
rect 1452 1615 1453 1619
rect 1474 1619 1480 1620
rect 1447 1614 1453 1615
rect 1462 1615 1468 1616
rect 1422 1610 1428 1611
rect 1462 1611 1463 1615
rect 1467 1611 1468 1615
rect 1474 1615 1475 1619
rect 1479 1618 1480 1619
rect 1487 1619 1493 1620
rect 1487 1618 1488 1619
rect 1479 1616 1488 1618
rect 1479 1615 1480 1616
rect 1474 1614 1480 1615
rect 1487 1615 1488 1616
rect 1492 1615 1493 1619
rect 1514 1619 1520 1620
rect 1487 1614 1493 1615
rect 1502 1615 1508 1616
rect 1462 1610 1468 1611
rect 1502 1611 1503 1615
rect 1507 1611 1508 1615
rect 1514 1615 1515 1619
rect 1519 1618 1520 1619
rect 1527 1619 1533 1620
rect 1527 1618 1528 1619
rect 1519 1616 1528 1618
rect 1519 1615 1520 1616
rect 1514 1614 1520 1615
rect 1527 1615 1528 1616
rect 1532 1615 1533 1619
rect 1583 1619 1589 1620
rect 1527 1614 1533 1615
rect 1558 1615 1564 1616
rect 1502 1610 1508 1611
rect 1558 1611 1559 1615
rect 1563 1611 1564 1615
rect 1583 1615 1584 1619
rect 1588 1618 1589 1619
rect 1622 1619 1628 1620
rect 1622 1618 1623 1619
rect 1588 1616 1623 1618
rect 1588 1615 1589 1616
rect 1583 1614 1589 1615
rect 1622 1615 1623 1616
rect 1627 1615 1628 1619
rect 1655 1619 1661 1620
rect 1622 1614 1628 1615
rect 1630 1615 1636 1616
rect 1558 1610 1564 1611
rect 1630 1611 1631 1615
rect 1635 1611 1636 1615
rect 1655 1615 1656 1619
rect 1660 1618 1661 1619
rect 1694 1619 1700 1620
rect 1694 1618 1695 1619
rect 1660 1616 1695 1618
rect 1660 1615 1661 1616
rect 1655 1614 1661 1615
rect 1694 1615 1695 1616
rect 1699 1615 1700 1619
rect 1727 1619 1733 1620
rect 1694 1614 1700 1615
rect 1702 1615 1708 1616
rect 1630 1610 1636 1611
rect 1702 1611 1703 1615
rect 1707 1611 1708 1615
rect 1727 1615 1728 1619
rect 1732 1618 1733 1619
rect 1774 1619 1780 1620
rect 1774 1618 1775 1619
rect 1732 1616 1775 1618
rect 1732 1615 1733 1616
rect 1727 1614 1733 1615
rect 1774 1615 1775 1616
rect 1779 1615 1780 1619
rect 1794 1619 1800 1620
rect 1774 1614 1780 1615
rect 1782 1615 1788 1616
rect 1702 1610 1708 1611
rect 1782 1611 1783 1615
rect 1787 1611 1788 1615
rect 1794 1615 1795 1619
rect 1799 1618 1800 1619
rect 1807 1619 1813 1620
rect 1807 1618 1808 1619
rect 1799 1616 1808 1618
rect 1799 1615 1800 1616
rect 1794 1614 1800 1615
rect 1807 1615 1808 1616
rect 1812 1615 1813 1619
rect 1879 1619 1885 1620
rect 1807 1614 1813 1615
rect 1854 1615 1860 1616
rect 1782 1610 1788 1611
rect 1854 1611 1855 1615
rect 1859 1611 1860 1615
rect 1879 1615 1880 1619
rect 1884 1618 1885 1619
rect 1918 1619 1924 1620
rect 1918 1618 1919 1619
rect 1884 1616 1919 1618
rect 1884 1615 1885 1616
rect 1879 1614 1885 1615
rect 1918 1615 1919 1616
rect 1923 1615 1924 1619
rect 1951 1619 1960 1620
rect 1918 1614 1924 1615
rect 1926 1615 1932 1616
rect 1854 1610 1860 1611
rect 1926 1611 1927 1615
rect 1931 1611 1932 1615
rect 1951 1615 1952 1619
rect 1959 1615 1960 1619
rect 2010 1619 2016 1620
rect 1951 1614 1960 1615
rect 1998 1615 2004 1616
rect 1926 1610 1932 1611
rect 1998 1611 1999 1615
rect 2003 1611 2004 1615
rect 2010 1615 2011 1619
rect 2015 1618 2016 1619
rect 2023 1619 2029 1620
rect 2023 1618 2024 1619
rect 2015 1616 2024 1618
rect 2015 1615 2016 1616
rect 2010 1614 2016 1615
rect 2023 1615 2024 1616
rect 2028 1615 2029 1619
rect 2087 1619 2093 1620
rect 2023 1614 2029 1615
rect 2062 1615 2068 1616
rect 1998 1610 2004 1611
rect 2062 1611 2063 1615
rect 2067 1611 2068 1615
rect 2087 1615 2088 1619
rect 2092 1618 2093 1619
rect 2118 1619 2124 1620
rect 2118 1618 2119 1619
rect 2092 1616 2119 1618
rect 2092 1615 2093 1616
rect 2087 1614 2093 1615
rect 2118 1615 2119 1616
rect 2123 1615 2124 1619
rect 2151 1619 2157 1620
rect 2118 1614 2124 1615
rect 2126 1615 2132 1616
rect 2062 1610 2068 1611
rect 2126 1611 2127 1615
rect 2131 1611 2132 1615
rect 2151 1615 2152 1619
rect 2156 1618 2157 1619
rect 2182 1619 2188 1620
rect 2182 1618 2183 1619
rect 2156 1616 2183 1618
rect 2156 1615 2157 1616
rect 2151 1614 2157 1615
rect 2182 1615 2183 1616
rect 2187 1615 2188 1619
rect 2202 1619 2208 1620
rect 2182 1614 2188 1615
rect 2190 1615 2196 1616
rect 2126 1610 2132 1611
rect 2190 1611 2191 1615
rect 2195 1611 2196 1615
rect 2202 1615 2203 1619
rect 2207 1618 2208 1619
rect 2215 1619 2221 1620
rect 2215 1618 2216 1619
rect 2207 1616 2216 1618
rect 2207 1615 2208 1616
rect 2202 1614 2208 1615
rect 2215 1615 2216 1616
rect 2220 1615 2221 1619
rect 2278 1619 2285 1620
rect 2215 1614 2221 1615
rect 2254 1615 2260 1616
rect 2190 1610 2196 1611
rect 2254 1611 2255 1615
rect 2259 1611 2260 1615
rect 2278 1615 2279 1619
rect 2284 1615 2285 1619
rect 2330 1619 2336 1620
rect 2278 1614 2285 1615
rect 2318 1615 2324 1616
rect 2254 1610 2260 1611
rect 2318 1611 2319 1615
rect 2323 1611 2324 1615
rect 2330 1615 2331 1619
rect 2335 1618 2336 1619
rect 2343 1619 2349 1620
rect 2343 1618 2344 1619
rect 2335 1616 2344 1618
rect 2335 1615 2336 1616
rect 2330 1614 2336 1615
rect 2343 1615 2344 1616
rect 2348 1615 2349 1619
rect 2370 1619 2376 1620
rect 2343 1614 2349 1615
rect 2358 1615 2364 1616
rect 2318 1610 2324 1611
rect 2358 1611 2359 1615
rect 2363 1611 2364 1615
rect 2370 1615 2371 1619
rect 2375 1618 2376 1619
rect 2383 1619 2389 1620
rect 2383 1618 2384 1619
rect 2375 1616 2384 1618
rect 2375 1615 2376 1616
rect 2370 1614 2376 1615
rect 2383 1615 2384 1616
rect 2388 1615 2389 1619
rect 2383 1614 2389 1615
rect 2358 1610 2364 1611
rect 172 1604 243 1606
rect 172 1603 173 1604
rect 167 1602 173 1603
rect 162 1595 168 1596
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 162 1591 163 1595
rect 167 1594 168 1595
rect 570 1595 576 1596
rect 570 1594 571 1595
rect 167 1592 203 1594
rect 167 1591 168 1592
rect 162 1590 168 1591
rect 201 1588 203 1592
rect 400 1592 571 1594
rect 110 1587 116 1588
rect 159 1587 165 1588
rect 159 1583 160 1587
rect 164 1586 165 1587
rect 167 1587 173 1588
rect 167 1586 168 1587
rect 164 1584 168 1586
rect 164 1583 165 1584
rect 159 1582 165 1583
rect 167 1583 168 1584
rect 172 1583 173 1587
rect 167 1582 173 1583
rect 199 1587 205 1588
rect 199 1583 200 1587
rect 204 1583 205 1587
rect 199 1582 205 1583
rect 239 1587 245 1588
rect 239 1583 240 1587
rect 244 1586 245 1587
rect 266 1587 272 1588
rect 266 1586 267 1587
rect 244 1584 267 1586
rect 244 1583 245 1584
rect 239 1582 245 1583
rect 266 1583 267 1584
rect 271 1583 272 1587
rect 266 1582 272 1583
rect 279 1587 285 1588
rect 279 1583 280 1587
rect 284 1586 285 1587
rect 326 1587 332 1588
rect 326 1586 327 1587
rect 284 1584 327 1586
rect 284 1583 285 1584
rect 279 1582 285 1583
rect 326 1583 327 1584
rect 331 1583 332 1587
rect 326 1582 332 1583
rect 335 1587 341 1588
rect 335 1583 336 1587
rect 340 1586 341 1587
rect 400 1586 402 1592
rect 570 1591 571 1592
rect 575 1591 576 1595
rect 866 1595 872 1596
rect 866 1594 867 1595
rect 570 1590 576 1591
rect 665 1592 867 1594
rect 665 1588 667 1592
rect 866 1591 867 1592
rect 871 1591 872 1595
rect 1058 1595 1064 1596
rect 1058 1594 1059 1595
rect 866 1590 872 1591
rect 924 1592 1059 1594
rect 340 1584 402 1586
rect 406 1587 412 1588
rect 340 1583 341 1584
rect 335 1582 341 1583
rect 406 1583 407 1587
rect 411 1586 412 1587
rect 415 1587 421 1588
rect 415 1586 416 1587
rect 411 1584 416 1586
rect 411 1583 412 1584
rect 406 1582 412 1583
rect 415 1583 416 1584
rect 420 1583 421 1587
rect 415 1582 421 1583
rect 462 1587 468 1588
rect 462 1583 463 1587
rect 467 1586 468 1587
rect 495 1587 501 1588
rect 495 1586 496 1587
rect 467 1584 496 1586
rect 467 1583 468 1584
rect 462 1582 468 1583
rect 495 1583 496 1584
rect 500 1583 501 1587
rect 495 1582 501 1583
rect 550 1587 556 1588
rect 550 1583 551 1587
rect 555 1586 556 1587
rect 583 1587 589 1588
rect 583 1586 584 1587
rect 555 1584 584 1586
rect 555 1583 556 1584
rect 550 1582 556 1583
rect 583 1583 584 1584
rect 588 1583 589 1587
rect 583 1582 589 1583
rect 663 1587 669 1588
rect 663 1583 664 1587
rect 668 1583 669 1587
rect 663 1582 669 1583
rect 710 1587 716 1588
rect 710 1583 711 1587
rect 715 1586 716 1587
rect 743 1587 749 1588
rect 743 1586 744 1587
rect 715 1584 744 1586
rect 715 1583 716 1584
rect 710 1582 716 1583
rect 743 1583 744 1584
rect 748 1583 749 1587
rect 743 1582 749 1583
rect 782 1587 788 1588
rect 782 1583 783 1587
rect 787 1586 788 1587
rect 815 1587 821 1588
rect 815 1586 816 1587
rect 787 1584 816 1586
rect 787 1583 788 1584
rect 782 1582 788 1583
rect 815 1583 816 1584
rect 820 1583 821 1587
rect 815 1582 821 1583
rect 879 1587 885 1588
rect 879 1583 880 1587
rect 884 1586 885 1587
rect 924 1586 926 1592
rect 1058 1591 1059 1592
rect 1063 1591 1064 1595
rect 1438 1595 1444 1596
rect 1438 1594 1439 1595
rect 1058 1590 1064 1591
rect 1238 1592 1244 1593
rect 1238 1588 1239 1592
rect 1243 1588 1244 1592
rect 884 1584 926 1586
rect 930 1587 936 1588
rect 884 1583 885 1584
rect 879 1582 885 1583
rect 930 1583 931 1587
rect 935 1586 936 1587
rect 943 1587 949 1588
rect 943 1586 944 1587
rect 935 1584 944 1586
rect 935 1583 936 1584
rect 930 1582 936 1583
rect 943 1583 944 1584
rect 948 1583 949 1587
rect 943 1582 949 1583
rect 974 1587 980 1588
rect 974 1583 975 1587
rect 979 1586 980 1587
rect 1007 1587 1013 1588
rect 1007 1586 1008 1587
rect 979 1584 1008 1586
rect 979 1583 980 1584
rect 974 1582 980 1583
rect 1007 1583 1008 1584
rect 1012 1583 1013 1587
rect 1007 1582 1013 1583
rect 1038 1587 1044 1588
rect 1038 1583 1039 1587
rect 1043 1586 1044 1587
rect 1071 1587 1077 1588
rect 1238 1587 1244 1588
rect 1278 1592 1284 1593
rect 1278 1588 1279 1592
rect 1283 1588 1284 1592
rect 1352 1592 1439 1594
rect 1278 1587 1284 1588
rect 1327 1587 1333 1588
rect 1071 1586 1072 1587
rect 1043 1584 1072 1586
rect 1043 1583 1044 1584
rect 1038 1582 1044 1583
rect 1071 1583 1072 1584
rect 1076 1583 1077 1587
rect 1071 1582 1077 1583
rect 1327 1583 1328 1587
rect 1332 1586 1333 1587
rect 1352 1586 1354 1592
rect 1438 1591 1439 1592
rect 1443 1591 1444 1595
rect 1514 1595 1520 1596
rect 1514 1594 1515 1595
rect 1438 1590 1444 1591
rect 1504 1592 1515 1594
rect 1332 1584 1354 1586
rect 1358 1587 1364 1588
rect 1332 1583 1333 1584
rect 1327 1582 1333 1583
rect 1358 1583 1359 1587
rect 1363 1586 1364 1587
rect 1367 1587 1373 1588
rect 1367 1586 1368 1587
rect 1363 1584 1368 1586
rect 1363 1583 1364 1584
rect 1358 1582 1364 1583
rect 1367 1583 1368 1584
rect 1372 1583 1373 1587
rect 1367 1582 1373 1583
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1586 1404 1587
rect 1407 1587 1413 1588
rect 1407 1586 1408 1587
rect 1403 1584 1408 1586
rect 1403 1583 1404 1584
rect 1398 1582 1404 1583
rect 1407 1583 1408 1584
rect 1412 1583 1413 1587
rect 1407 1582 1413 1583
rect 1447 1587 1453 1588
rect 1447 1583 1448 1587
rect 1452 1586 1453 1587
rect 1474 1587 1480 1588
rect 1474 1586 1475 1587
rect 1452 1584 1475 1586
rect 1452 1583 1453 1584
rect 1447 1582 1453 1583
rect 1474 1583 1475 1584
rect 1479 1583 1480 1587
rect 1474 1582 1480 1583
rect 1487 1587 1493 1588
rect 1487 1583 1488 1587
rect 1492 1586 1493 1587
rect 1504 1586 1506 1592
rect 1514 1591 1515 1592
rect 1519 1591 1520 1595
rect 1663 1595 1669 1596
rect 1663 1594 1664 1595
rect 1514 1590 1520 1591
rect 1585 1592 1664 1594
rect 1585 1588 1587 1592
rect 1663 1591 1664 1592
rect 1668 1591 1669 1595
rect 2010 1595 2016 1596
rect 2010 1594 2011 1595
rect 1663 1590 1669 1591
rect 1881 1592 2011 1594
rect 1881 1588 1883 1592
rect 2010 1591 2011 1592
rect 2015 1591 2016 1595
rect 2202 1595 2208 1596
rect 2202 1594 2203 1595
rect 2010 1590 2016 1591
rect 2036 1592 2203 1594
rect 1492 1584 1506 1586
rect 1510 1587 1516 1588
rect 1492 1583 1493 1584
rect 1487 1582 1493 1583
rect 1510 1583 1511 1587
rect 1515 1586 1516 1587
rect 1527 1587 1533 1588
rect 1527 1586 1528 1587
rect 1515 1584 1528 1586
rect 1515 1583 1516 1584
rect 1510 1582 1516 1583
rect 1527 1583 1528 1584
rect 1532 1583 1533 1587
rect 1527 1582 1533 1583
rect 1583 1587 1589 1588
rect 1583 1583 1584 1587
rect 1588 1583 1589 1587
rect 1583 1582 1589 1583
rect 1622 1587 1628 1588
rect 1622 1583 1623 1587
rect 1627 1586 1628 1587
rect 1655 1587 1661 1588
rect 1655 1586 1656 1587
rect 1627 1584 1656 1586
rect 1627 1583 1628 1584
rect 1622 1582 1628 1583
rect 1655 1583 1656 1584
rect 1660 1583 1661 1587
rect 1655 1582 1661 1583
rect 1694 1587 1700 1588
rect 1694 1583 1695 1587
rect 1699 1586 1700 1587
rect 1727 1587 1733 1588
rect 1727 1586 1728 1587
rect 1699 1584 1728 1586
rect 1699 1583 1700 1584
rect 1694 1582 1700 1583
rect 1727 1583 1728 1584
rect 1732 1583 1733 1587
rect 1727 1582 1733 1583
rect 1774 1587 1780 1588
rect 1774 1583 1775 1587
rect 1779 1586 1780 1587
rect 1807 1587 1813 1588
rect 1807 1586 1808 1587
rect 1779 1584 1808 1586
rect 1779 1583 1780 1584
rect 1774 1582 1780 1583
rect 1807 1583 1808 1584
rect 1812 1583 1813 1587
rect 1807 1582 1813 1583
rect 1879 1587 1885 1588
rect 1879 1583 1880 1587
rect 1884 1583 1885 1587
rect 1879 1582 1885 1583
rect 1918 1587 1924 1588
rect 1918 1583 1919 1587
rect 1923 1586 1924 1587
rect 1951 1587 1957 1588
rect 1951 1586 1952 1587
rect 1923 1584 1952 1586
rect 1923 1583 1924 1584
rect 1918 1582 1924 1583
rect 1951 1583 1952 1584
rect 1956 1583 1957 1587
rect 1951 1582 1957 1583
rect 2023 1587 2029 1588
rect 2023 1583 2024 1587
rect 2028 1586 2029 1587
rect 2036 1586 2038 1592
rect 2202 1591 2203 1592
rect 2207 1591 2208 1595
rect 2202 1590 2208 1591
rect 2406 1592 2412 1593
rect 2406 1588 2407 1592
rect 2411 1588 2412 1592
rect 2028 1584 2038 1586
rect 2042 1587 2048 1588
rect 2028 1583 2029 1584
rect 2023 1582 2029 1583
rect 2042 1583 2043 1587
rect 2047 1586 2048 1587
rect 2087 1587 2093 1588
rect 2087 1586 2088 1587
rect 2047 1584 2088 1586
rect 2047 1583 2048 1584
rect 2042 1582 2048 1583
rect 2087 1583 2088 1584
rect 2092 1583 2093 1587
rect 2087 1582 2093 1583
rect 2118 1587 2124 1588
rect 2118 1583 2119 1587
rect 2123 1586 2124 1587
rect 2151 1587 2157 1588
rect 2151 1586 2152 1587
rect 2123 1584 2152 1586
rect 2123 1583 2124 1584
rect 2118 1582 2124 1583
rect 2151 1583 2152 1584
rect 2156 1583 2157 1587
rect 2151 1582 2157 1583
rect 2182 1587 2188 1588
rect 2182 1583 2183 1587
rect 2187 1586 2188 1587
rect 2215 1587 2221 1588
rect 2215 1586 2216 1587
rect 2187 1584 2216 1586
rect 2187 1583 2188 1584
rect 2182 1582 2188 1583
rect 2215 1583 2216 1584
rect 2220 1583 2221 1587
rect 2215 1582 2221 1583
rect 2279 1587 2285 1588
rect 2279 1583 2280 1587
rect 2284 1586 2285 1587
rect 2330 1587 2336 1588
rect 2330 1586 2331 1587
rect 2284 1584 2331 1586
rect 2284 1583 2285 1584
rect 2279 1582 2285 1583
rect 2330 1583 2331 1584
rect 2335 1583 2336 1587
rect 2330 1582 2336 1583
rect 2343 1587 2349 1588
rect 2343 1583 2344 1587
rect 2348 1586 2349 1587
rect 2370 1587 2376 1588
rect 2370 1586 2371 1587
rect 2348 1584 2371 1586
rect 2348 1583 2349 1584
rect 2343 1582 2349 1583
rect 2370 1583 2371 1584
rect 2375 1583 2376 1587
rect 2370 1582 2376 1583
rect 2383 1587 2389 1588
rect 2406 1587 2412 1588
rect 2383 1583 2384 1587
rect 2388 1583 2389 1587
rect 2383 1582 2389 1583
rect 2346 1579 2352 1580
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 110 1570 116 1571
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1278 1575 1284 1576
rect 1278 1571 1279 1575
rect 1283 1571 1284 1575
rect 2346 1575 2347 1579
rect 2351 1578 2352 1579
rect 2385 1578 2387 1582
rect 2351 1576 2387 1578
rect 2351 1575 2352 1576
rect 2346 1574 2352 1575
rect 2406 1575 2412 1576
rect 1278 1570 1284 1571
rect 2406 1571 2407 1575
rect 2411 1571 2412 1575
rect 2406 1570 2412 1571
rect 134 1568 140 1569
rect 134 1564 135 1568
rect 139 1564 140 1568
rect 134 1563 140 1564
rect 174 1568 180 1569
rect 174 1564 175 1568
rect 179 1564 180 1568
rect 174 1563 180 1564
rect 214 1568 220 1569
rect 214 1564 215 1568
rect 219 1564 220 1568
rect 214 1563 220 1564
rect 254 1568 260 1569
rect 254 1564 255 1568
rect 259 1564 260 1568
rect 254 1563 260 1564
rect 310 1568 316 1569
rect 310 1564 311 1568
rect 315 1564 316 1568
rect 310 1563 316 1564
rect 390 1568 396 1569
rect 390 1564 391 1568
rect 395 1564 396 1568
rect 390 1563 396 1564
rect 470 1568 476 1569
rect 470 1564 471 1568
rect 475 1564 476 1568
rect 470 1563 476 1564
rect 558 1568 564 1569
rect 558 1564 559 1568
rect 563 1564 564 1568
rect 558 1563 564 1564
rect 638 1568 644 1569
rect 638 1564 639 1568
rect 643 1564 644 1568
rect 638 1563 644 1564
rect 718 1568 724 1569
rect 718 1564 719 1568
rect 723 1564 724 1568
rect 718 1563 724 1564
rect 790 1568 796 1569
rect 790 1564 791 1568
rect 795 1564 796 1568
rect 790 1563 796 1564
rect 854 1568 860 1569
rect 854 1564 855 1568
rect 859 1564 860 1568
rect 854 1563 860 1564
rect 918 1568 924 1569
rect 918 1564 919 1568
rect 923 1564 924 1568
rect 918 1563 924 1564
rect 982 1568 988 1569
rect 982 1564 983 1568
rect 987 1564 988 1568
rect 982 1563 988 1564
rect 1046 1568 1052 1569
rect 1046 1564 1047 1568
rect 1051 1564 1052 1568
rect 1046 1563 1052 1564
rect 1302 1568 1308 1569
rect 1302 1564 1303 1568
rect 1307 1564 1308 1568
rect 1302 1563 1308 1564
rect 1342 1568 1348 1569
rect 1342 1564 1343 1568
rect 1347 1564 1348 1568
rect 1342 1563 1348 1564
rect 1382 1568 1388 1569
rect 1382 1564 1383 1568
rect 1387 1564 1388 1568
rect 1382 1563 1388 1564
rect 1422 1568 1428 1569
rect 1422 1564 1423 1568
rect 1427 1564 1428 1568
rect 1422 1563 1428 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1502 1568 1508 1569
rect 1502 1564 1503 1568
rect 1507 1564 1508 1568
rect 1502 1563 1508 1564
rect 1558 1568 1564 1569
rect 1558 1564 1559 1568
rect 1563 1564 1564 1568
rect 1558 1563 1564 1564
rect 1630 1568 1636 1569
rect 1630 1564 1631 1568
rect 1635 1564 1636 1568
rect 1630 1563 1636 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1782 1568 1788 1569
rect 1782 1564 1783 1568
rect 1787 1564 1788 1568
rect 1782 1563 1788 1564
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1926 1568 1932 1569
rect 1926 1564 1927 1568
rect 1931 1564 1932 1568
rect 1926 1563 1932 1564
rect 1998 1568 2004 1569
rect 1998 1564 1999 1568
rect 2003 1564 2004 1568
rect 1998 1563 2004 1564
rect 2062 1568 2068 1569
rect 2062 1564 2063 1568
rect 2067 1564 2068 1568
rect 2062 1563 2068 1564
rect 2126 1568 2132 1569
rect 2126 1564 2127 1568
rect 2131 1564 2132 1568
rect 2126 1563 2132 1564
rect 2190 1568 2196 1569
rect 2190 1564 2191 1568
rect 2195 1564 2196 1568
rect 2190 1563 2196 1564
rect 2254 1568 2260 1569
rect 2254 1564 2255 1568
rect 2259 1564 2260 1568
rect 2254 1563 2260 1564
rect 2318 1568 2324 1569
rect 2318 1564 2319 1568
rect 2323 1564 2324 1568
rect 2318 1563 2324 1564
rect 2358 1568 2364 1569
rect 2358 1564 2359 1568
rect 2363 1564 2364 1568
rect 2358 1563 2364 1564
rect 1470 1556 1476 1557
rect 150 1552 156 1553
rect 150 1548 151 1552
rect 155 1548 156 1552
rect 150 1547 156 1548
rect 198 1552 204 1553
rect 198 1548 199 1552
rect 203 1548 204 1552
rect 198 1547 204 1548
rect 262 1552 268 1553
rect 262 1548 263 1552
rect 267 1548 268 1552
rect 262 1547 268 1548
rect 342 1552 348 1553
rect 342 1548 343 1552
rect 347 1548 348 1552
rect 342 1547 348 1548
rect 438 1552 444 1553
rect 438 1548 439 1552
rect 443 1548 444 1552
rect 438 1547 444 1548
rect 534 1552 540 1553
rect 534 1548 535 1552
rect 539 1548 540 1552
rect 534 1547 540 1548
rect 638 1552 644 1553
rect 638 1548 639 1552
rect 643 1548 644 1552
rect 638 1547 644 1548
rect 734 1552 740 1553
rect 734 1548 735 1552
rect 739 1548 740 1552
rect 734 1547 740 1548
rect 822 1552 828 1553
rect 822 1548 823 1552
rect 827 1548 828 1552
rect 822 1547 828 1548
rect 902 1552 908 1553
rect 902 1548 903 1552
rect 907 1548 908 1552
rect 902 1547 908 1548
rect 974 1552 980 1553
rect 974 1548 975 1552
rect 979 1548 980 1552
rect 974 1547 980 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1118 1552 1124 1553
rect 1118 1548 1119 1552
rect 1123 1548 1124 1552
rect 1118 1547 1124 1548
rect 1190 1552 1196 1553
rect 1190 1548 1191 1552
rect 1195 1548 1196 1552
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1758 1556 1764 1557
rect 1758 1552 1759 1556
rect 1763 1552 1764 1556
rect 1758 1551 1764 1552
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 1966 1556 1972 1557
rect 1966 1552 1967 1556
rect 1971 1552 1972 1556
rect 1966 1551 1972 1552
rect 2054 1556 2060 1557
rect 2054 1552 2055 1556
rect 2059 1552 2060 1556
rect 2054 1551 2060 1552
rect 2126 1556 2132 1557
rect 2126 1552 2127 1556
rect 2131 1552 2132 1556
rect 2126 1551 2132 1552
rect 2190 1556 2196 1557
rect 2190 1552 2191 1556
rect 2195 1552 2196 1556
rect 2190 1551 2196 1552
rect 2254 1556 2260 1557
rect 2254 1552 2255 1556
rect 2259 1552 2260 1556
rect 2254 1551 2260 1552
rect 2318 1556 2324 1557
rect 2318 1552 2319 1556
rect 2323 1552 2324 1556
rect 2318 1551 2324 1552
rect 2358 1556 2364 1557
rect 2358 1552 2359 1556
rect 2363 1552 2364 1556
rect 2358 1551 2364 1552
rect 1190 1547 1196 1548
rect 1278 1549 1284 1550
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 110 1540 116 1541
rect 1238 1545 1244 1546
rect 1238 1541 1239 1545
rect 1243 1541 1244 1545
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1278 1544 1284 1545
rect 2406 1549 2412 1550
rect 2406 1545 2407 1549
rect 2411 1545 2412 1549
rect 2406 1544 2412 1545
rect 1794 1543 1800 1544
rect 1794 1542 1795 1543
rect 1238 1540 1244 1541
rect 1732 1540 1795 1542
rect 1495 1535 1501 1536
rect 1278 1532 1284 1533
rect 175 1531 181 1532
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 175 1527 176 1531
rect 180 1530 181 1531
rect 186 1531 192 1532
rect 186 1530 187 1531
rect 180 1528 187 1530
rect 180 1527 181 1528
rect 175 1526 181 1527
rect 186 1527 187 1528
rect 191 1527 192 1531
rect 186 1526 192 1527
rect 206 1531 212 1532
rect 206 1527 207 1531
rect 211 1530 212 1531
rect 223 1531 229 1532
rect 223 1530 224 1531
rect 211 1528 224 1530
rect 211 1527 212 1528
rect 206 1526 212 1527
rect 223 1527 224 1528
rect 228 1527 229 1531
rect 223 1526 229 1527
rect 231 1531 237 1532
rect 231 1527 232 1531
rect 236 1530 237 1531
rect 287 1531 293 1532
rect 287 1530 288 1531
rect 236 1528 288 1530
rect 236 1527 237 1528
rect 231 1526 237 1527
rect 287 1527 288 1528
rect 292 1527 293 1531
rect 287 1526 293 1527
rect 295 1531 301 1532
rect 295 1527 296 1531
rect 300 1530 301 1531
rect 367 1531 373 1532
rect 367 1530 368 1531
rect 300 1528 368 1530
rect 300 1527 301 1528
rect 295 1526 301 1527
rect 367 1527 368 1528
rect 372 1527 373 1531
rect 367 1526 373 1527
rect 375 1531 381 1532
rect 375 1527 376 1531
rect 380 1530 381 1531
rect 463 1531 469 1532
rect 463 1530 464 1531
rect 380 1528 464 1530
rect 380 1527 381 1528
rect 375 1526 381 1527
rect 463 1527 464 1528
rect 468 1527 469 1531
rect 463 1526 469 1527
rect 471 1531 477 1532
rect 471 1527 472 1531
rect 476 1530 477 1531
rect 559 1531 565 1532
rect 559 1530 560 1531
rect 476 1528 560 1530
rect 476 1527 477 1528
rect 471 1526 477 1527
rect 559 1527 560 1528
rect 564 1527 565 1531
rect 559 1526 565 1527
rect 567 1531 573 1532
rect 567 1527 568 1531
rect 572 1530 573 1531
rect 663 1531 669 1532
rect 663 1530 664 1531
rect 572 1528 664 1530
rect 572 1527 573 1528
rect 567 1526 573 1527
rect 663 1527 664 1528
rect 668 1527 669 1531
rect 663 1526 669 1527
rect 759 1531 765 1532
rect 759 1527 760 1531
rect 764 1527 765 1531
rect 759 1526 765 1527
rect 767 1531 773 1532
rect 767 1527 768 1531
rect 772 1530 773 1531
rect 847 1531 853 1532
rect 847 1530 848 1531
rect 772 1528 848 1530
rect 772 1527 773 1528
rect 767 1526 773 1527
rect 847 1527 848 1528
rect 852 1527 853 1531
rect 847 1526 853 1527
rect 855 1531 861 1532
rect 855 1527 856 1531
rect 860 1530 861 1531
rect 927 1531 933 1532
rect 927 1530 928 1531
rect 860 1528 928 1530
rect 860 1527 861 1528
rect 855 1526 861 1527
rect 927 1527 928 1528
rect 932 1527 933 1531
rect 927 1526 933 1527
rect 999 1531 1005 1532
rect 999 1527 1000 1531
rect 1004 1530 1005 1531
rect 1062 1531 1068 1532
rect 1062 1530 1063 1531
rect 1004 1528 1063 1530
rect 1004 1527 1005 1528
rect 999 1526 1005 1527
rect 1062 1527 1063 1528
rect 1067 1527 1068 1531
rect 1062 1526 1068 1527
rect 1071 1531 1077 1532
rect 1071 1527 1072 1531
rect 1076 1530 1077 1531
rect 1134 1531 1140 1532
rect 1134 1530 1135 1531
rect 1076 1528 1135 1530
rect 1076 1527 1077 1528
rect 1071 1526 1077 1527
rect 1134 1527 1135 1528
rect 1139 1527 1140 1531
rect 1134 1526 1140 1527
rect 1143 1531 1149 1532
rect 1143 1527 1144 1531
rect 1148 1530 1149 1531
rect 1206 1531 1212 1532
rect 1206 1530 1207 1531
rect 1148 1528 1207 1530
rect 1148 1527 1149 1528
rect 1143 1526 1149 1527
rect 1206 1527 1207 1528
rect 1211 1527 1212 1531
rect 1206 1526 1212 1527
rect 1215 1531 1221 1532
rect 1215 1527 1216 1531
rect 1220 1527 1221 1531
rect 1215 1526 1221 1527
rect 1238 1528 1244 1529
rect 110 1523 116 1524
rect 760 1522 762 1526
rect 998 1523 1004 1524
rect 998 1522 999 1523
rect 760 1520 999 1522
rect 998 1519 999 1520
rect 1003 1519 1004 1523
rect 998 1518 1004 1519
rect 1178 1523 1184 1524
rect 1178 1519 1179 1523
rect 1183 1522 1184 1523
rect 1217 1522 1219 1526
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1278 1528 1279 1532
rect 1283 1528 1284 1532
rect 1495 1531 1496 1535
rect 1500 1534 1501 1535
rect 1638 1535 1644 1536
rect 1638 1534 1639 1535
rect 1500 1532 1639 1534
rect 1500 1531 1501 1532
rect 1495 1530 1501 1531
rect 1638 1531 1639 1532
rect 1643 1531 1644 1535
rect 1638 1530 1644 1531
rect 1647 1535 1653 1536
rect 1647 1531 1648 1535
rect 1652 1534 1653 1535
rect 1732 1534 1734 1540
rect 1794 1539 1795 1540
rect 1799 1539 1800 1543
rect 1794 1538 1800 1539
rect 1652 1532 1734 1534
rect 1783 1535 1789 1536
rect 1652 1531 1653 1532
rect 1647 1530 1653 1531
rect 1783 1531 1784 1535
rect 1788 1531 1789 1535
rect 1783 1530 1789 1531
rect 1791 1535 1797 1536
rect 1791 1531 1792 1535
rect 1796 1534 1797 1535
rect 1895 1535 1901 1536
rect 1895 1534 1896 1535
rect 1796 1532 1896 1534
rect 1796 1531 1797 1532
rect 1791 1530 1797 1531
rect 1895 1531 1896 1532
rect 1900 1531 1901 1535
rect 1895 1530 1901 1531
rect 1903 1535 1909 1536
rect 1903 1531 1904 1535
rect 1908 1534 1909 1535
rect 1991 1535 1997 1536
rect 1991 1534 1992 1535
rect 1908 1532 1992 1534
rect 1908 1531 1909 1532
rect 1903 1530 1909 1531
rect 1991 1531 1992 1532
rect 1996 1531 1997 1535
rect 1991 1530 1997 1531
rect 2079 1535 2085 1536
rect 2079 1531 2080 1535
rect 2084 1534 2085 1535
rect 2142 1535 2148 1536
rect 2142 1534 2143 1535
rect 2084 1532 2143 1534
rect 2084 1531 2085 1532
rect 2079 1530 2085 1531
rect 2142 1531 2143 1532
rect 2147 1531 2148 1535
rect 2142 1530 2148 1531
rect 2151 1535 2157 1536
rect 2151 1531 2152 1535
rect 2156 1534 2157 1535
rect 2206 1535 2212 1536
rect 2206 1534 2207 1535
rect 2156 1532 2207 1534
rect 2156 1531 2157 1532
rect 2151 1530 2157 1531
rect 2206 1531 2207 1532
rect 2211 1531 2212 1535
rect 2206 1530 2212 1531
rect 2215 1535 2221 1536
rect 2215 1531 2216 1535
rect 2220 1534 2221 1535
rect 2270 1535 2276 1536
rect 2270 1534 2271 1535
rect 2220 1532 2271 1534
rect 2220 1531 2221 1532
rect 2215 1530 2221 1531
rect 2270 1531 2271 1532
rect 2275 1531 2276 1535
rect 2270 1530 2276 1531
rect 2278 1535 2285 1536
rect 2278 1531 2279 1535
rect 2284 1531 2285 1535
rect 2278 1530 2285 1531
rect 2343 1535 2349 1536
rect 2343 1531 2344 1535
rect 2348 1534 2349 1535
rect 2374 1535 2380 1536
rect 2374 1534 2375 1535
rect 2348 1532 2375 1534
rect 2348 1531 2349 1532
rect 2343 1530 2349 1531
rect 2374 1531 2375 1532
rect 2379 1531 2380 1535
rect 2374 1530 2380 1531
rect 2382 1535 2389 1536
rect 2382 1531 2383 1535
rect 2388 1531 2389 1535
rect 2382 1530 2389 1531
rect 2406 1532 2412 1533
rect 1278 1527 1284 1528
rect 1785 1526 1787 1530
rect 2406 1528 2407 1532
rect 2411 1528 2412 1532
rect 2078 1527 2084 1528
rect 2406 1527 2412 1528
rect 2078 1526 2079 1527
rect 1785 1524 2079 1526
rect 1238 1523 1244 1524
rect 2078 1523 2079 1524
rect 2083 1523 2084 1527
rect 2078 1522 2084 1523
rect 1183 1520 1219 1522
rect 1183 1519 1184 1520
rect 1178 1518 1184 1519
rect 1470 1509 1476 1510
rect 150 1505 156 1506
rect 150 1501 151 1505
rect 155 1501 156 1505
rect 150 1500 156 1501
rect 198 1505 204 1506
rect 198 1501 199 1505
rect 203 1501 204 1505
rect 198 1500 204 1501
rect 262 1505 268 1506
rect 262 1501 263 1505
rect 267 1501 268 1505
rect 262 1500 268 1501
rect 342 1505 348 1506
rect 342 1501 343 1505
rect 347 1501 348 1505
rect 342 1500 348 1501
rect 438 1505 444 1506
rect 438 1501 439 1505
rect 443 1501 444 1505
rect 438 1500 444 1501
rect 534 1505 540 1506
rect 534 1501 535 1505
rect 539 1501 540 1505
rect 534 1500 540 1501
rect 638 1505 644 1506
rect 638 1501 639 1505
rect 643 1501 644 1505
rect 638 1500 644 1501
rect 734 1505 740 1506
rect 734 1501 735 1505
rect 739 1501 740 1505
rect 734 1500 740 1501
rect 822 1505 828 1506
rect 822 1501 823 1505
rect 827 1501 828 1505
rect 822 1500 828 1501
rect 902 1505 908 1506
rect 902 1501 903 1505
rect 907 1501 908 1505
rect 902 1500 908 1501
rect 974 1505 980 1506
rect 974 1501 975 1505
rect 979 1501 980 1505
rect 974 1500 980 1501
rect 1046 1505 1052 1506
rect 1046 1501 1047 1505
rect 1051 1501 1052 1505
rect 1046 1500 1052 1501
rect 1118 1505 1124 1506
rect 1118 1501 1119 1505
rect 1123 1501 1124 1505
rect 1118 1500 1124 1501
rect 1190 1505 1196 1506
rect 1190 1501 1191 1505
rect 1195 1501 1196 1505
rect 1470 1505 1471 1509
rect 1475 1505 1476 1509
rect 1470 1504 1476 1505
rect 1622 1509 1628 1510
rect 1622 1505 1623 1509
rect 1627 1505 1628 1509
rect 1622 1504 1628 1505
rect 1758 1509 1764 1510
rect 1758 1505 1759 1509
rect 1763 1505 1764 1509
rect 1758 1504 1764 1505
rect 1870 1509 1876 1510
rect 1870 1505 1871 1509
rect 1875 1505 1876 1509
rect 1870 1504 1876 1505
rect 1966 1509 1972 1510
rect 1966 1505 1967 1509
rect 1971 1505 1972 1509
rect 1966 1504 1972 1505
rect 2054 1509 2060 1510
rect 2054 1505 2055 1509
rect 2059 1505 2060 1509
rect 2054 1504 2060 1505
rect 2126 1509 2132 1510
rect 2126 1505 2127 1509
rect 2131 1505 2132 1509
rect 2126 1504 2132 1505
rect 2190 1509 2196 1510
rect 2190 1505 2191 1509
rect 2195 1505 2196 1509
rect 2190 1504 2196 1505
rect 2254 1509 2260 1510
rect 2254 1505 2255 1509
rect 2259 1505 2260 1509
rect 2254 1504 2260 1505
rect 2318 1509 2324 1510
rect 2318 1505 2319 1509
rect 2323 1505 2324 1509
rect 2318 1504 2324 1505
rect 2358 1509 2364 1510
rect 2358 1505 2359 1509
rect 2363 1505 2364 1509
rect 2358 1504 2364 1505
rect 1190 1500 1196 1501
rect 1495 1503 1501 1504
rect 175 1499 181 1500
rect 175 1495 176 1499
rect 180 1498 181 1499
rect 206 1499 212 1500
rect 206 1498 207 1499
rect 180 1496 207 1498
rect 180 1495 181 1496
rect 175 1494 181 1495
rect 206 1495 207 1496
rect 211 1495 212 1499
rect 206 1494 212 1495
rect 223 1499 229 1500
rect 223 1495 224 1499
rect 228 1498 229 1499
rect 231 1499 237 1500
rect 231 1498 232 1499
rect 228 1496 232 1498
rect 228 1495 229 1496
rect 223 1494 229 1495
rect 231 1495 232 1496
rect 236 1495 237 1499
rect 231 1494 237 1495
rect 287 1499 293 1500
rect 287 1495 288 1499
rect 292 1498 293 1499
rect 295 1499 301 1500
rect 295 1498 296 1499
rect 292 1496 296 1498
rect 292 1495 293 1496
rect 287 1494 293 1495
rect 295 1495 296 1496
rect 300 1495 301 1499
rect 295 1494 301 1495
rect 367 1499 373 1500
rect 367 1495 368 1499
rect 372 1498 373 1499
rect 375 1499 381 1500
rect 375 1498 376 1499
rect 372 1496 376 1498
rect 372 1495 373 1496
rect 367 1494 373 1495
rect 375 1495 376 1496
rect 380 1495 381 1499
rect 375 1494 381 1495
rect 463 1499 469 1500
rect 463 1495 464 1499
rect 468 1498 469 1499
rect 471 1499 477 1500
rect 471 1498 472 1499
rect 468 1496 472 1498
rect 468 1495 469 1496
rect 463 1494 469 1495
rect 471 1495 472 1496
rect 476 1495 477 1499
rect 471 1494 477 1495
rect 559 1499 565 1500
rect 559 1495 560 1499
rect 564 1498 565 1499
rect 567 1499 573 1500
rect 567 1498 568 1499
rect 564 1496 568 1498
rect 564 1495 565 1496
rect 559 1494 565 1495
rect 567 1495 568 1496
rect 572 1495 573 1499
rect 567 1494 573 1495
rect 578 1499 584 1500
rect 578 1495 579 1499
rect 583 1498 584 1499
rect 663 1499 669 1500
rect 663 1498 664 1499
rect 583 1496 664 1498
rect 583 1495 584 1496
rect 578 1494 584 1495
rect 663 1495 664 1496
rect 668 1495 669 1499
rect 663 1494 669 1495
rect 759 1499 765 1500
rect 759 1495 760 1499
rect 764 1498 765 1499
rect 767 1499 773 1500
rect 767 1498 768 1499
rect 764 1496 768 1498
rect 764 1495 765 1496
rect 759 1494 765 1495
rect 767 1495 768 1496
rect 772 1495 773 1499
rect 767 1494 773 1495
rect 847 1499 853 1500
rect 847 1495 848 1499
rect 852 1498 853 1499
rect 855 1499 861 1500
rect 855 1498 856 1499
rect 852 1496 856 1498
rect 852 1495 853 1496
rect 847 1494 853 1495
rect 855 1495 856 1496
rect 860 1495 861 1499
rect 855 1494 861 1495
rect 927 1499 936 1500
rect 927 1495 928 1499
rect 935 1495 936 1499
rect 927 1494 936 1495
rect 998 1499 1005 1500
rect 998 1495 999 1499
rect 1004 1495 1005 1499
rect 998 1494 1005 1495
rect 1062 1499 1068 1500
rect 1062 1495 1063 1499
rect 1067 1498 1068 1499
rect 1071 1499 1077 1500
rect 1071 1498 1072 1499
rect 1067 1496 1072 1498
rect 1067 1495 1068 1496
rect 1062 1494 1068 1495
rect 1071 1495 1072 1496
rect 1076 1495 1077 1499
rect 1071 1494 1077 1495
rect 1134 1499 1140 1500
rect 1134 1495 1135 1499
rect 1139 1498 1140 1499
rect 1143 1499 1149 1500
rect 1143 1498 1144 1499
rect 1139 1496 1144 1498
rect 1139 1495 1140 1496
rect 1134 1494 1140 1495
rect 1143 1495 1144 1496
rect 1148 1495 1149 1499
rect 1143 1494 1149 1495
rect 1206 1499 1212 1500
rect 1206 1495 1207 1499
rect 1211 1498 1212 1499
rect 1215 1499 1221 1500
rect 1215 1498 1216 1499
rect 1211 1496 1216 1498
rect 1211 1495 1212 1496
rect 1206 1494 1212 1495
rect 1215 1495 1216 1496
rect 1220 1495 1221 1499
rect 1495 1499 1496 1503
rect 1500 1502 1501 1503
rect 1510 1503 1516 1504
rect 1510 1502 1511 1503
rect 1500 1500 1511 1502
rect 1500 1499 1501 1500
rect 1495 1498 1501 1499
rect 1510 1499 1511 1500
rect 1515 1499 1516 1503
rect 1510 1498 1516 1499
rect 1638 1503 1644 1504
rect 1638 1499 1639 1503
rect 1643 1502 1644 1503
rect 1647 1503 1653 1504
rect 1647 1502 1648 1503
rect 1643 1500 1648 1502
rect 1643 1499 1644 1500
rect 1638 1498 1644 1499
rect 1647 1499 1648 1500
rect 1652 1499 1653 1503
rect 1647 1498 1653 1499
rect 1783 1503 1789 1504
rect 1783 1499 1784 1503
rect 1788 1502 1789 1503
rect 1791 1503 1797 1504
rect 1791 1502 1792 1503
rect 1788 1500 1792 1502
rect 1788 1499 1789 1500
rect 1783 1498 1789 1499
rect 1791 1499 1792 1500
rect 1796 1499 1797 1503
rect 1791 1498 1797 1499
rect 1895 1503 1901 1504
rect 1895 1499 1896 1503
rect 1900 1502 1901 1503
rect 1903 1503 1909 1504
rect 1903 1502 1904 1503
rect 1900 1500 1904 1502
rect 1900 1499 1901 1500
rect 1895 1498 1901 1499
rect 1903 1499 1904 1500
rect 1908 1499 1909 1503
rect 1903 1498 1909 1499
rect 1991 1503 1997 1504
rect 1991 1499 1992 1503
rect 1996 1502 1997 1503
rect 2042 1503 2048 1504
rect 2042 1502 2043 1503
rect 1996 1500 2043 1502
rect 1996 1499 1997 1500
rect 1991 1498 1997 1499
rect 2042 1499 2043 1500
rect 2047 1499 2048 1503
rect 2042 1498 2048 1499
rect 2078 1503 2085 1504
rect 2078 1499 2079 1503
rect 2084 1499 2085 1503
rect 2078 1498 2085 1499
rect 2142 1503 2148 1504
rect 2142 1499 2143 1503
rect 2147 1502 2148 1503
rect 2151 1503 2157 1504
rect 2151 1502 2152 1503
rect 2147 1500 2152 1502
rect 2147 1499 2148 1500
rect 2142 1498 2148 1499
rect 2151 1499 2152 1500
rect 2156 1499 2157 1503
rect 2151 1498 2157 1499
rect 2206 1503 2212 1504
rect 2206 1499 2207 1503
rect 2211 1502 2212 1503
rect 2215 1503 2221 1504
rect 2215 1502 2216 1503
rect 2211 1500 2216 1502
rect 2211 1499 2212 1500
rect 2206 1498 2212 1499
rect 2215 1499 2216 1500
rect 2220 1499 2221 1503
rect 2215 1498 2221 1499
rect 2270 1503 2276 1504
rect 2270 1499 2271 1503
rect 2275 1502 2276 1503
rect 2279 1503 2285 1504
rect 2279 1502 2280 1503
rect 2275 1500 2280 1502
rect 2275 1499 2276 1500
rect 2270 1498 2276 1499
rect 2279 1499 2280 1500
rect 2284 1499 2285 1503
rect 2279 1498 2285 1499
rect 2343 1503 2352 1504
rect 2343 1499 2344 1503
rect 2351 1499 2352 1503
rect 2343 1498 2352 1499
rect 2374 1503 2380 1504
rect 2374 1499 2375 1503
rect 2379 1502 2380 1503
rect 2383 1503 2389 1504
rect 2383 1502 2384 1503
rect 2379 1500 2384 1502
rect 2379 1499 2380 1500
rect 2374 1498 2380 1499
rect 2383 1499 2384 1500
rect 2388 1499 2389 1503
rect 2383 1498 2389 1499
rect 1215 1494 1221 1495
rect 414 1479 420 1480
rect 414 1478 415 1479
rect 392 1476 415 1478
rect 343 1475 352 1476
rect 318 1471 324 1472
rect 318 1467 319 1471
rect 323 1467 324 1471
rect 343 1471 344 1475
rect 351 1471 352 1475
rect 383 1475 389 1476
rect 343 1470 352 1471
rect 358 1471 364 1472
rect 318 1466 324 1467
rect 358 1467 359 1471
rect 363 1467 364 1471
rect 383 1471 384 1475
rect 388 1474 389 1475
rect 392 1474 394 1476
rect 414 1475 415 1476
rect 419 1475 420 1479
rect 414 1474 420 1475
rect 423 1475 429 1476
rect 388 1472 394 1474
rect 388 1471 389 1472
rect 383 1470 389 1471
rect 398 1471 404 1472
rect 358 1466 364 1467
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 423 1471 424 1475
rect 428 1474 429 1475
rect 438 1475 444 1476
rect 438 1474 439 1475
rect 428 1472 439 1474
rect 428 1471 429 1472
rect 423 1470 429 1471
rect 438 1471 439 1472
rect 443 1471 444 1475
rect 471 1475 477 1476
rect 438 1470 444 1471
rect 446 1471 452 1472
rect 398 1466 404 1467
rect 446 1467 447 1471
rect 451 1467 452 1471
rect 471 1471 472 1475
rect 476 1474 477 1475
rect 494 1475 500 1476
rect 494 1474 495 1475
rect 476 1472 495 1474
rect 476 1471 477 1472
rect 471 1470 477 1471
rect 494 1471 495 1472
rect 499 1471 500 1475
rect 527 1475 533 1476
rect 494 1470 500 1471
rect 502 1471 508 1472
rect 446 1466 452 1467
rect 502 1467 503 1471
rect 507 1467 508 1471
rect 527 1471 528 1475
rect 532 1474 533 1475
rect 550 1475 556 1476
rect 550 1474 551 1475
rect 532 1472 551 1474
rect 532 1471 533 1472
rect 527 1470 533 1471
rect 550 1471 551 1472
rect 555 1471 556 1475
rect 583 1475 589 1476
rect 550 1470 556 1471
rect 558 1471 564 1472
rect 502 1466 508 1467
rect 558 1467 559 1471
rect 563 1467 564 1471
rect 583 1471 584 1475
rect 588 1474 589 1475
rect 606 1475 612 1476
rect 606 1474 607 1475
rect 588 1472 607 1474
rect 588 1471 589 1472
rect 583 1470 589 1471
rect 606 1471 607 1472
rect 611 1471 612 1475
rect 630 1475 636 1476
rect 606 1470 612 1471
rect 614 1471 620 1472
rect 558 1466 564 1467
rect 614 1467 615 1471
rect 619 1467 620 1471
rect 630 1471 631 1475
rect 635 1474 636 1475
rect 639 1475 645 1476
rect 639 1474 640 1475
rect 635 1472 640 1474
rect 635 1471 636 1472
rect 630 1470 636 1471
rect 639 1471 640 1472
rect 644 1471 645 1475
rect 695 1475 701 1476
rect 639 1470 645 1471
rect 670 1471 676 1472
rect 614 1466 620 1467
rect 670 1467 671 1471
rect 675 1467 676 1471
rect 695 1471 696 1475
rect 700 1474 701 1475
rect 726 1475 732 1476
rect 726 1474 727 1475
rect 700 1472 727 1474
rect 700 1471 701 1472
rect 695 1470 701 1471
rect 726 1471 727 1472
rect 731 1471 732 1475
rect 759 1475 765 1476
rect 726 1470 732 1471
rect 734 1471 740 1472
rect 670 1466 676 1467
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 759 1471 760 1475
rect 764 1474 765 1475
rect 790 1475 796 1476
rect 790 1474 791 1475
rect 764 1472 791 1474
rect 764 1471 765 1472
rect 759 1470 765 1471
rect 790 1471 791 1472
rect 795 1471 796 1475
rect 823 1475 829 1476
rect 790 1470 796 1471
rect 798 1471 804 1472
rect 734 1466 740 1467
rect 798 1467 799 1471
rect 803 1467 804 1471
rect 823 1471 824 1475
rect 828 1474 829 1475
rect 846 1475 852 1476
rect 846 1474 847 1475
rect 828 1472 847 1474
rect 828 1471 829 1472
rect 823 1470 829 1471
rect 846 1471 847 1472
rect 851 1471 852 1475
rect 879 1475 885 1476
rect 846 1470 852 1471
rect 854 1471 860 1472
rect 798 1466 804 1467
rect 854 1467 855 1471
rect 859 1467 860 1471
rect 879 1471 880 1475
rect 884 1474 885 1475
rect 902 1475 908 1476
rect 902 1474 903 1475
rect 884 1472 903 1474
rect 884 1471 885 1472
rect 879 1470 885 1471
rect 902 1471 903 1472
rect 907 1471 908 1475
rect 935 1475 941 1476
rect 902 1470 908 1471
rect 910 1471 916 1472
rect 854 1466 860 1467
rect 910 1467 911 1471
rect 915 1467 916 1471
rect 935 1471 936 1475
rect 940 1474 941 1475
rect 958 1475 964 1476
rect 958 1474 959 1475
rect 940 1472 959 1474
rect 940 1471 941 1472
rect 935 1470 941 1471
rect 958 1471 959 1472
rect 963 1471 964 1475
rect 991 1475 997 1476
rect 958 1470 964 1471
rect 966 1471 972 1472
rect 910 1466 916 1467
rect 966 1467 967 1471
rect 971 1467 972 1471
rect 991 1471 992 1475
rect 996 1474 997 1475
rect 1014 1475 1020 1476
rect 1014 1474 1015 1475
rect 996 1472 1015 1474
rect 996 1471 997 1472
rect 991 1470 997 1471
rect 1014 1471 1015 1472
rect 1019 1471 1020 1475
rect 1047 1475 1053 1476
rect 1014 1470 1020 1471
rect 1022 1471 1028 1472
rect 966 1466 972 1467
rect 1022 1467 1023 1471
rect 1027 1467 1028 1471
rect 1047 1471 1048 1475
rect 1052 1474 1053 1475
rect 1111 1475 1117 1476
rect 1052 1472 1082 1474
rect 1052 1471 1053 1472
rect 1047 1470 1053 1471
rect 1022 1466 1028 1467
rect 1080 1462 1082 1472
rect 1086 1471 1092 1472
rect 1086 1467 1087 1471
rect 1091 1467 1092 1471
rect 1111 1471 1112 1475
rect 1116 1474 1117 1475
rect 1135 1475 1141 1476
rect 1135 1474 1136 1475
rect 1116 1472 1136 1474
rect 1116 1471 1117 1472
rect 1111 1470 1117 1471
rect 1135 1471 1136 1472
rect 1140 1471 1141 1475
rect 1175 1475 1184 1476
rect 1135 1470 1141 1471
rect 1150 1471 1156 1472
rect 1086 1466 1092 1467
rect 1150 1467 1151 1471
rect 1155 1467 1156 1471
rect 1175 1471 1176 1475
rect 1183 1471 1184 1475
rect 1202 1475 1208 1476
rect 1175 1470 1184 1471
rect 1190 1471 1196 1472
rect 1150 1466 1156 1467
rect 1190 1467 1191 1471
rect 1195 1467 1196 1471
rect 1202 1471 1203 1475
rect 1207 1474 1208 1475
rect 1215 1475 1221 1476
rect 1215 1474 1216 1475
rect 1207 1472 1216 1474
rect 1207 1471 1208 1472
rect 1202 1470 1208 1471
rect 1215 1471 1216 1472
rect 1220 1471 1221 1475
rect 1215 1470 1221 1471
rect 1190 1466 1196 1467
rect 1218 1467 1224 1468
rect 1110 1463 1116 1464
rect 1110 1462 1111 1463
rect 1080 1460 1111 1462
rect 1110 1459 1111 1460
rect 1115 1459 1116 1463
rect 1218 1463 1219 1467
rect 1223 1466 1224 1467
rect 1223 1464 1314 1466
rect 1223 1463 1224 1464
rect 1218 1462 1224 1463
rect 1312 1462 1314 1464
rect 1327 1463 1333 1464
rect 1327 1462 1328 1463
rect 1312 1460 1328 1462
rect 1110 1458 1116 1459
rect 1302 1459 1308 1460
rect 1302 1455 1303 1459
rect 1307 1455 1308 1459
rect 1327 1459 1328 1460
rect 1332 1459 1333 1463
rect 1386 1463 1392 1464
rect 1327 1458 1333 1459
rect 1374 1459 1380 1460
rect 1302 1454 1308 1455
rect 1374 1455 1375 1459
rect 1379 1455 1380 1459
rect 1386 1459 1387 1463
rect 1391 1462 1392 1463
rect 1399 1463 1405 1464
rect 1399 1462 1400 1463
rect 1391 1460 1400 1462
rect 1391 1459 1392 1460
rect 1386 1458 1392 1459
rect 1399 1459 1400 1460
rect 1404 1459 1405 1463
rect 1503 1463 1509 1464
rect 1399 1458 1405 1459
rect 1478 1459 1484 1460
rect 1374 1454 1380 1455
rect 1478 1455 1479 1459
rect 1483 1455 1484 1459
rect 1503 1459 1504 1463
rect 1508 1462 1509 1463
rect 1574 1463 1580 1464
rect 1574 1462 1575 1463
rect 1508 1460 1575 1462
rect 1508 1459 1509 1460
rect 1503 1458 1509 1459
rect 1574 1459 1575 1460
rect 1579 1459 1580 1463
rect 1607 1463 1613 1464
rect 1574 1458 1580 1459
rect 1582 1459 1588 1460
rect 1478 1454 1484 1455
rect 1582 1455 1583 1459
rect 1587 1455 1588 1459
rect 1607 1459 1608 1463
rect 1612 1462 1613 1463
rect 1678 1463 1684 1464
rect 1678 1462 1679 1463
rect 1612 1460 1679 1462
rect 1612 1459 1613 1460
rect 1607 1458 1613 1459
rect 1678 1459 1679 1460
rect 1683 1459 1684 1463
rect 1698 1463 1704 1464
rect 1678 1458 1684 1459
rect 1686 1459 1692 1460
rect 1582 1454 1588 1455
rect 1686 1455 1687 1459
rect 1691 1455 1692 1459
rect 1698 1459 1699 1463
rect 1703 1462 1704 1463
rect 1711 1463 1717 1464
rect 1711 1462 1712 1463
rect 1703 1460 1712 1462
rect 1703 1459 1704 1460
rect 1698 1458 1704 1459
rect 1711 1459 1712 1460
rect 1716 1459 1717 1463
rect 1807 1463 1813 1464
rect 1711 1458 1717 1459
rect 1782 1459 1788 1460
rect 1686 1454 1692 1455
rect 1782 1455 1783 1459
rect 1787 1455 1788 1459
rect 1807 1459 1808 1463
rect 1812 1462 1813 1463
rect 1855 1463 1861 1464
rect 1855 1462 1856 1463
rect 1812 1460 1856 1462
rect 1812 1459 1813 1460
rect 1807 1458 1813 1459
rect 1855 1459 1856 1460
rect 1860 1459 1861 1463
rect 1895 1463 1901 1464
rect 1855 1458 1861 1459
rect 1870 1459 1876 1460
rect 1782 1454 1788 1455
rect 1870 1455 1871 1459
rect 1875 1455 1876 1459
rect 1895 1459 1896 1463
rect 1900 1462 1901 1463
rect 1942 1463 1948 1464
rect 1942 1462 1943 1463
rect 1900 1460 1943 1462
rect 1900 1459 1901 1460
rect 1895 1458 1901 1459
rect 1942 1459 1943 1460
rect 1947 1459 1948 1463
rect 1975 1463 1981 1464
rect 1942 1458 1948 1459
rect 1950 1459 1956 1460
rect 1870 1454 1876 1455
rect 1950 1455 1951 1459
rect 1955 1455 1956 1459
rect 1975 1459 1976 1463
rect 1980 1462 1981 1463
rect 2022 1463 2028 1464
rect 2022 1462 2023 1463
rect 1980 1460 2023 1462
rect 1980 1459 1981 1460
rect 1975 1458 1981 1459
rect 2022 1459 2023 1460
rect 2027 1459 2028 1463
rect 2055 1463 2061 1464
rect 2022 1458 2028 1459
rect 2030 1459 2036 1460
rect 1950 1454 1956 1455
rect 2030 1455 2031 1459
rect 2035 1455 2036 1459
rect 2055 1459 2056 1463
rect 2060 1462 2061 1463
rect 2094 1463 2100 1464
rect 2094 1462 2095 1463
rect 2060 1460 2095 1462
rect 2060 1459 2061 1460
rect 2055 1458 2061 1459
rect 2094 1459 2095 1460
rect 2099 1459 2100 1463
rect 2127 1463 2133 1464
rect 2094 1458 2100 1459
rect 2102 1459 2108 1460
rect 2030 1454 2036 1455
rect 2102 1455 2103 1459
rect 2107 1455 2108 1459
rect 2127 1459 2128 1463
rect 2132 1462 2133 1463
rect 2158 1463 2164 1464
rect 2158 1462 2159 1463
rect 2132 1460 2159 1462
rect 2132 1459 2133 1460
rect 2127 1458 2133 1459
rect 2158 1459 2159 1460
rect 2163 1459 2164 1463
rect 2191 1463 2197 1464
rect 2158 1458 2164 1459
rect 2166 1459 2172 1460
rect 2102 1454 2108 1455
rect 2166 1455 2167 1459
rect 2171 1455 2172 1459
rect 2191 1459 2192 1463
rect 2196 1462 2197 1463
rect 2230 1463 2236 1464
rect 2230 1462 2231 1463
rect 2196 1460 2231 1462
rect 2196 1459 2197 1460
rect 2191 1458 2197 1459
rect 2230 1459 2231 1460
rect 2235 1459 2236 1463
rect 2263 1463 2269 1464
rect 2230 1458 2236 1459
rect 2238 1459 2244 1460
rect 2166 1454 2172 1455
rect 2238 1455 2239 1459
rect 2243 1455 2244 1459
rect 2263 1459 2264 1463
rect 2268 1462 2269 1463
rect 2302 1463 2308 1464
rect 2302 1462 2303 1463
rect 2268 1460 2303 1462
rect 2268 1459 2269 1460
rect 2263 1458 2269 1459
rect 2302 1459 2303 1460
rect 2307 1459 2308 1463
rect 2322 1463 2328 1464
rect 2302 1458 2308 1459
rect 2310 1459 2316 1460
rect 2238 1454 2244 1455
rect 2310 1455 2311 1459
rect 2315 1455 2316 1459
rect 2322 1459 2323 1463
rect 2327 1462 2328 1463
rect 2335 1463 2341 1464
rect 2335 1462 2336 1463
rect 2327 1460 2336 1462
rect 2327 1459 2328 1460
rect 2322 1458 2328 1459
rect 2335 1459 2336 1460
rect 2340 1459 2341 1463
rect 2382 1463 2389 1464
rect 2335 1458 2341 1459
rect 2358 1459 2364 1460
rect 2310 1454 2316 1455
rect 2358 1455 2359 1459
rect 2363 1455 2364 1459
rect 2382 1459 2383 1463
rect 2388 1459 2389 1463
rect 2382 1458 2389 1459
rect 2358 1454 2364 1455
rect 346 1451 352 1452
rect 110 1448 116 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 346 1447 347 1451
rect 351 1450 352 1451
rect 1202 1451 1208 1452
rect 1202 1450 1203 1451
rect 351 1448 366 1450
rect 351 1447 352 1448
rect 346 1446 352 1447
rect 110 1443 116 1444
rect 343 1443 349 1444
rect 343 1439 344 1443
rect 348 1442 349 1443
rect 364 1442 366 1448
rect 1104 1448 1203 1450
rect 383 1443 389 1444
rect 383 1442 384 1443
rect 348 1440 362 1442
rect 364 1440 384 1442
rect 348 1439 349 1440
rect 343 1438 349 1439
rect 360 1434 362 1440
rect 383 1439 384 1440
rect 388 1439 389 1443
rect 383 1438 389 1439
rect 414 1443 420 1444
rect 414 1439 415 1443
rect 419 1442 420 1443
rect 423 1443 429 1444
rect 423 1442 424 1443
rect 419 1440 424 1442
rect 419 1439 420 1440
rect 414 1438 420 1439
rect 423 1439 424 1440
rect 428 1439 429 1443
rect 423 1438 429 1439
rect 438 1443 444 1444
rect 438 1439 439 1443
rect 443 1442 444 1443
rect 471 1443 477 1444
rect 471 1442 472 1443
rect 443 1440 472 1442
rect 443 1439 444 1440
rect 438 1438 444 1439
rect 471 1439 472 1440
rect 476 1439 477 1443
rect 471 1438 477 1439
rect 494 1443 500 1444
rect 494 1439 495 1443
rect 499 1442 500 1443
rect 527 1443 533 1444
rect 527 1442 528 1443
rect 499 1440 528 1442
rect 499 1439 500 1440
rect 494 1438 500 1439
rect 527 1439 528 1440
rect 532 1439 533 1443
rect 527 1438 533 1439
rect 550 1443 556 1444
rect 550 1439 551 1443
rect 555 1442 556 1443
rect 583 1443 589 1444
rect 583 1442 584 1443
rect 555 1440 584 1442
rect 555 1439 556 1440
rect 550 1438 556 1439
rect 583 1439 584 1440
rect 588 1439 589 1443
rect 583 1438 589 1439
rect 606 1443 612 1444
rect 606 1439 607 1443
rect 611 1442 612 1443
rect 639 1443 645 1444
rect 639 1442 640 1443
rect 611 1440 640 1442
rect 611 1439 612 1440
rect 606 1438 612 1439
rect 639 1439 640 1440
rect 644 1439 645 1443
rect 639 1438 645 1439
rect 695 1443 701 1444
rect 695 1439 696 1443
rect 700 1442 701 1443
rect 726 1443 732 1444
rect 700 1440 722 1442
rect 700 1439 701 1440
rect 695 1438 701 1439
rect 578 1435 584 1436
rect 578 1434 579 1435
rect 360 1432 579 1434
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 578 1431 579 1432
rect 583 1431 584 1435
rect 720 1434 722 1440
rect 726 1439 727 1443
rect 731 1442 732 1443
rect 759 1443 765 1444
rect 759 1442 760 1443
rect 731 1440 760 1442
rect 731 1439 732 1440
rect 726 1438 732 1439
rect 759 1439 760 1440
rect 764 1439 765 1443
rect 759 1438 765 1439
rect 790 1443 796 1444
rect 790 1439 791 1443
rect 795 1442 796 1443
rect 823 1443 829 1444
rect 823 1442 824 1443
rect 795 1440 824 1442
rect 795 1439 796 1440
rect 790 1438 796 1439
rect 823 1439 824 1440
rect 828 1439 829 1443
rect 823 1438 829 1439
rect 846 1443 852 1444
rect 846 1439 847 1443
rect 851 1442 852 1443
rect 879 1443 885 1444
rect 879 1442 880 1443
rect 851 1440 880 1442
rect 851 1439 852 1440
rect 846 1438 852 1439
rect 879 1439 880 1440
rect 884 1439 885 1443
rect 879 1438 885 1439
rect 902 1443 908 1444
rect 902 1439 903 1443
rect 907 1442 908 1443
rect 935 1443 941 1444
rect 935 1442 936 1443
rect 907 1440 936 1442
rect 907 1439 908 1440
rect 902 1438 908 1439
rect 935 1439 936 1440
rect 940 1439 941 1443
rect 935 1438 941 1439
rect 958 1443 964 1444
rect 958 1439 959 1443
rect 963 1442 964 1443
rect 991 1443 997 1444
rect 991 1442 992 1443
rect 963 1440 992 1442
rect 963 1439 964 1440
rect 958 1438 964 1439
rect 991 1439 992 1440
rect 996 1439 997 1443
rect 991 1438 997 1439
rect 1047 1443 1053 1444
rect 1047 1439 1048 1443
rect 1052 1442 1053 1443
rect 1104 1442 1106 1448
rect 1202 1447 1203 1448
rect 1207 1447 1208 1451
rect 1202 1446 1208 1447
rect 1238 1448 1244 1449
rect 1238 1444 1239 1448
rect 1243 1444 1244 1448
rect 1052 1440 1106 1442
rect 1110 1443 1117 1444
rect 1052 1439 1053 1440
rect 1047 1438 1053 1439
rect 1110 1439 1111 1443
rect 1116 1439 1117 1443
rect 1110 1438 1117 1439
rect 1135 1443 1141 1444
rect 1135 1439 1136 1443
rect 1140 1442 1141 1443
rect 1175 1443 1181 1444
rect 1175 1442 1176 1443
rect 1140 1440 1176 1442
rect 1140 1439 1141 1440
rect 1135 1438 1141 1439
rect 1175 1439 1176 1440
rect 1180 1439 1181 1443
rect 1175 1438 1181 1439
rect 1215 1443 1224 1444
rect 1238 1443 1244 1444
rect 1215 1439 1216 1443
rect 1223 1439 1224 1443
rect 1215 1438 1224 1439
rect 1698 1439 1704 1440
rect 1698 1438 1699 1439
rect 1278 1436 1284 1437
rect 838 1435 844 1436
rect 838 1434 839 1435
rect 720 1432 839 1434
rect 578 1430 584 1431
rect 838 1431 839 1432
rect 843 1431 844 1435
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1452 1436 1699 1438
rect 838 1430 844 1431
rect 1238 1431 1244 1432
rect 1278 1431 1284 1432
rect 1327 1431 1333 1432
rect 110 1426 116 1427
rect 1238 1427 1239 1431
rect 1243 1427 1244 1431
rect 1238 1426 1244 1427
rect 1327 1427 1328 1431
rect 1332 1430 1333 1431
rect 1386 1431 1392 1432
rect 1386 1430 1387 1431
rect 1332 1428 1387 1430
rect 1332 1427 1333 1428
rect 1327 1426 1333 1427
rect 1386 1427 1387 1428
rect 1391 1427 1392 1431
rect 1386 1426 1392 1427
rect 1399 1431 1405 1432
rect 1399 1427 1400 1431
rect 1404 1430 1405 1431
rect 1452 1430 1454 1436
rect 1698 1435 1699 1436
rect 1703 1435 1704 1439
rect 1698 1434 1704 1435
rect 1855 1439 1861 1440
rect 1855 1435 1856 1439
rect 1860 1438 1861 1439
rect 1860 1436 1898 1438
rect 1860 1435 1861 1436
rect 1855 1434 1861 1435
rect 1896 1434 1898 1436
rect 2406 1436 2412 1437
rect 1895 1433 1901 1434
rect 1404 1428 1454 1430
rect 1458 1431 1464 1432
rect 1404 1427 1405 1428
rect 1399 1426 1405 1427
rect 1458 1427 1459 1431
rect 1463 1430 1464 1431
rect 1503 1431 1509 1432
rect 1503 1430 1504 1431
rect 1463 1428 1504 1430
rect 1463 1427 1464 1428
rect 1458 1426 1464 1427
rect 1503 1427 1504 1428
rect 1508 1427 1509 1431
rect 1503 1426 1509 1427
rect 1574 1431 1580 1432
rect 1574 1427 1575 1431
rect 1579 1430 1580 1431
rect 1607 1431 1613 1432
rect 1607 1430 1608 1431
rect 1579 1428 1608 1430
rect 1579 1427 1580 1428
rect 1574 1426 1580 1427
rect 1607 1427 1608 1428
rect 1612 1427 1613 1431
rect 1607 1426 1613 1427
rect 1678 1431 1684 1432
rect 1678 1427 1679 1431
rect 1683 1430 1684 1431
rect 1711 1431 1717 1432
rect 1711 1430 1712 1431
rect 1683 1428 1712 1430
rect 1683 1427 1684 1428
rect 1678 1426 1684 1427
rect 1711 1427 1712 1428
rect 1716 1427 1717 1431
rect 1711 1426 1717 1427
rect 1807 1431 1813 1432
rect 1807 1427 1808 1431
rect 1812 1430 1813 1431
rect 1812 1428 1890 1430
rect 1895 1429 1896 1433
rect 1900 1429 1901 1433
rect 2406 1432 2407 1436
rect 2411 1432 2412 1436
rect 1895 1428 1901 1429
rect 1942 1431 1948 1432
rect 1812 1427 1813 1428
rect 1807 1426 1813 1427
rect 318 1424 324 1425
rect 318 1420 319 1424
rect 323 1420 324 1424
rect 318 1419 324 1420
rect 358 1424 364 1425
rect 358 1420 359 1424
rect 363 1420 364 1424
rect 358 1419 364 1420
rect 398 1424 404 1425
rect 398 1420 399 1424
rect 403 1420 404 1424
rect 398 1419 404 1420
rect 446 1424 452 1425
rect 446 1420 447 1424
rect 451 1420 452 1424
rect 446 1419 452 1420
rect 502 1424 508 1425
rect 502 1420 503 1424
rect 507 1420 508 1424
rect 502 1419 508 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 614 1424 620 1425
rect 614 1420 615 1424
rect 619 1420 620 1424
rect 614 1419 620 1420
rect 670 1424 676 1425
rect 670 1420 671 1424
rect 675 1420 676 1424
rect 670 1419 676 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 798 1424 804 1425
rect 798 1420 799 1424
rect 803 1420 804 1424
rect 798 1419 804 1420
rect 854 1424 860 1425
rect 854 1420 855 1424
rect 859 1420 860 1424
rect 854 1419 860 1420
rect 910 1424 916 1425
rect 910 1420 911 1424
rect 915 1420 916 1424
rect 910 1419 916 1420
rect 966 1424 972 1425
rect 966 1420 967 1424
rect 971 1420 972 1424
rect 966 1419 972 1420
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1086 1424 1092 1425
rect 1086 1420 1087 1424
rect 1091 1420 1092 1424
rect 1086 1419 1092 1420
rect 1150 1424 1156 1425
rect 1150 1420 1151 1424
rect 1155 1420 1156 1424
rect 1150 1419 1156 1420
rect 1190 1424 1196 1425
rect 1190 1420 1191 1424
rect 1195 1420 1196 1424
rect 1888 1422 1890 1428
rect 1942 1427 1943 1431
rect 1947 1430 1948 1431
rect 1975 1431 1981 1432
rect 1975 1430 1976 1431
rect 1947 1428 1976 1430
rect 1947 1427 1948 1428
rect 1942 1426 1948 1427
rect 1975 1427 1976 1428
rect 1980 1427 1981 1431
rect 1975 1426 1981 1427
rect 2022 1431 2028 1432
rect 2022 1427 2023 1431
rect 2027 1430 2028 1431
rect 2055 1431 2061 1432
rect 2055 1430 2056 1431
rect 2027 1428 2056 1430
rect 2027 1427 2028 1428
rect 2022 1426 2028 1427
rect 2055 1427 2056 1428
rect 2060 1427 2061 1431
rect 2055 1426 2061 1427
rect 2094 1431 2100 1432
rect 2094 1427 2095 1431
rect 2099 1430 2100 1431
rect 2127 1431 2133 1432
rect 2127 1430 2128 1431
rect 2099 1428 2128 1430
rect 2099 1427 2100 1428
rect 2094 1426 2100 1427
rect 2127 1427 2128 1428
rect 2132 1427 2133 1431
rect 2127 1426 2133 1427
rect 2158 1431 2164 1432
rect 2158 1427 2159 1431
rect 2163 1430 2164 1431
rect 2191 1431 2197 1432
rect 2191 1430 2192 1431
rect 2163 1428 2192 1430
rect 2163 1427 2164 1428
rect 2158 1426 2164 1427
rect 2191 1427 2192 1428
rect 2196 1427 2197 1431
rect 2191 1426 2197 1427
rect 2230 1431 2236 1432
rect 2230 1427 2231 1431
rect 2235 1430 2236 1431
rect 2263 1431 2269 1432
rect 2263 1430 2264 1431
rect 2235 1428 2264 1430
rect 2235 1427 2236 1428
rect 2230 1426 2236 1427
rect 2263 1427 2264 1428
rect 2268 1427 2269 1431
rect 2263 1426 2269 1427
rect 2302 1431 2308 1432
rect 2302 1427 2303 1431
rect 2307 1430 2308 1431
rect 2335 1431 2341 1432
rect 2335 1430 2336 1431
rect 2307 1428 2336 1430
rect 2307 1427 2308 1428
rect 2302 1426 2308 1427
rect 2335 1427 2336 1428
rect 2340 1427 2341 1431
rect 2335 1426 2341 1427
rect 2343 1431 2349 1432
rect 2343 1427 2344 1431
rect 2348 1430 2349 1431
rect 2383 1431 2389 1432
rect 2406 1431 2412 1432
rect 2383 1430 2384 1431
rect 2348 1428 2384 1430
rect 2348 1427 2349 1428
rect 2343 1426 2349 1427
rect 2383 1427 2384 1428
rect 2388 1427 2389 1431
rect 2383 1426 2389 1427
rect 2094 1423 2100 1424
rect 2094 1422 2095 1423
rect 1888 1420 2095 1422
rect 1190 1419 1196 1420
rect 1278 1419 1284 1420
rect 1278 1415 1279 1419
rect 1283 1415 1284 1419
rect 2094 1419 2095 1420
rect 2099 1419 2100 1423
rect 2094 1418 2100 1419
rect 2406 1419 2412 1420
rect 1278 1414 1284 1415
rect 2406 1415 2407 1419
rect 2411 1415 2412 1419
rect 2406 1414 2412 1415
rect 1302 1412 1308 1413
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 302 1408 308 1409
rect 302 1404 303 1408
rect 307 1404 308 1408
rect 302 1403 308 1404
rect 342 1408 348 1409
rect 342 1404 343 1408
rect 347 1404 348 1408
rect 342 1403 348 1404
rect 390 1408 396 1409
rect 390 1404 391 1408
rect 395 1404 396 1408
rect 390 1403 396 1404
rect 446 1408 452 1409
rect 446 1404 447 1408
rect 451 1404 452 1408
rect 446 1403 452 1404
rect 502 1408 508 1409
rect 502 1404 503 1408
rect 507 1404 508 1408
rect 502 1403 508 1404
rect 558 1408 564 1409
rect 558 1404 559 1408
rect 563 1404 564 1408
rect 558 1403 564 1404
rect 622 1408 628 1409
rect 622 1404 623 1408
rect 627 1404 628 1408
rect 622 1403 628 1404
rect 686 1408 692 1409
rect 686 1404 687 1408
rect 691 1404 692 1408
rect 686 1403 692 1404
rect 750 1408 756 1409
rect 750 1404 751 1408
rect 755 1404 756 1408
rect 750 1403 756 1404
rect 814 1408 820 1409
rect 814 1404 815 1408
rect 819 1404 820 1408
rect 814 1403 820 1404
rect 878 1408 884 1409
rect 878 1404 879 1408
rect 883 1404 884 1408
rect 878 1403 884 1404
rect 950 1408 956 1409
rect 950 1404 951 1408
rect 955 1404 956 1408
rect 950 1403 956 1404
rect 1022 1408 1028 1409
rect 1022 1404 1023 1408
rect 1027 1404 1028 1408
rect 1302 1408 1303 1412
rect 1307 1408 1308 1412
rect 1302 1407 1308 1408
rect 1374 1412 1380 1413
rect 1374 1408 1375 1412
rect 1379 1408 1380 1412
rect 1374 1407 1380 1408
rect 1478 1412 1484 1413
rect 1478 1408 1479 1412
rect 1483 1408 1484 1412
rect 1478 1407 1484 1408
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1582 1407 1588 1408
rect 1686 1412 1692 1413
rect 1686 1408 1687 1412
rect 1691 1408 1692 1412
rect 1686 1407 1692 1408
rect 1782 1412 1788 1413
rect 1782 1408 1783 1412
rect 1787 1408 1788 1412
rect 1782 1407 1788 1408
rect 1870 1412 1876 1413
rect 1870 1408 1871 1412
rect 1875 1408 1876 1412
rect 1870 1407 1876 1408
rect 1950 1412 1956 1413
rect 1950 1408 1951 1412
rect 1955 1408 1956 1412
rect 1950 1407 1956 1408
rect 2030 1412 2036 1413
rect 2030 1408 2031 1412
rect 2035 1408 2036 1412
rect 2030 1407 2036 1408
rect 2102 1412 2108 1413
rect 2102 1408 2103 1412
rect 2107 1408 2108 1412
rect 2102 1407 2108 1408
rect 2166 1412 2172 1413
rect 2166 1408 2167 1412
rect 2171 1408 2172 1412
rect 2166 1407 2172 1408
rect 2238 1412 2244 1413
rect 2238 1408 2239 1412
rect 2243 1408 2244 1412
rect 2238 1407 2244 1408
rect 2310 1412 2316 1413
rect 2310 1408 2311 1412
rect 2315 1408 2316 1412
rect 2310 1407 2316 1408
rect 2358 1412 2364 1413
rect 2358 1408 2359 1412
rect 2363 1408 2364 1412
rect 2358 1407 2364 1408
rect 1022 1403 1028 1404
rect 110 1401 116 1402
rect 110 1397 111 1401
rect 115 1397 116 1401
rect 110 1396 116 1397
rect 1238 1401 1244 1402
rect 1238 1397 1239 1401
rect 1243 1397 1244 1401
rect 1238 1396 1244 1397
rect 1302 1400 1308 1401
rect 1302 1396 1303 1400
rect 1307 1396 1308 1400
rect 1014 1395 1020 1396
rect 1302 1395 1308 1396
rect 1342 1400 1348 1401
rect 1342 1396 1343 1400
rect 1347 1396 1348 1400
rect 1342 1395 1348 1396
rect 1398 1400 1404 1401
rect 1398 1396 1399 1400
rect 1403 1396 1404 1400
rect 1398 1395 1404 1396
rect 1470 1400 1476 1401
rect 1470 1396 1471 1400
rect 1475 1396 1476 1400
rect 1470 1395 1476 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1814 1400 1820 1401
rect 1814 1396 1815 1400
rect 1819 1396 1820 1400
rect 1814 1395 1820 1396
rect 1902 1400 1908 1401
rect 1902 1396 1903 1400
rect 1907 1396 1908 1400
rect 1902 1395 1908 1396
rect 1990 1400 1996 1401
rect 1990 1396 1991 1400
rect 1995 1396 1996 1400
rect 1990 1395 1996 1396
rect 2070 1400 2076 1401
rect 2070 1396 2071 1400
rect 2075 1396 2076 1400
rect 2070 1395 2076 1396
rect 2150 1400 2156 1401
rect 2150 1396 2151 1400
rect 2155 1396 2156 1400
rect 2150 1395 2156 1396
rect 2222 1400 2228 1401
rect 2222 1396 2223 1400
rect 2227 1396 2228 1400
rect 2222 1395 2228 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 1014 1391 1015 1395
rect 1019 1394 1020 1395
rect 1019 1392 1050 1394
rect 1019 1391 1020 1392
rect 1014 1390 1020 1391
rect 1048 1388 1050 1392
rect 1278 1393 1284 1394
rect 1278 1389 1279 1393
rect 1283 1389 1284 1393
rect 1278 1388 1284 1389
rect 2406 1393 2412 1394
rect 2406 1389 2407 1393
rect 2411 1389 2412 1393
rect 2406 1388 2412 1389
rect 287 1387 293 1388
rect 110 1384 116 1385
rect 110 1380 111 1384
rect 115 1380 116 1384
rect 287 1383 288 1387
rect 292 1386 293 1387
rect 310 1387 316 1388
rect 292 1384 306 1386
rect 292 1383 293 1384
rect 287 1382 293 1383
rect 110 1379 116 1380
rect 304 1378 306 1384
rect 310 1383 311 1387
rect 315 1386 316 1387
rect 327 1387 333 1388
rect 327 1386 328 1387
rect 315 1384 328 1386
rect 315 1383 316 1384
rect 310 1382 316 1383
rect 327 1383 328 1384
rect 332 1383 333 1387
rect 327 1382 333 1383
rect 367 1387 373 1388
rect 367 1383 368 1387
rect 372 1386 373 1387
rect 406 1387 412 1388
rect 406 1386 407 1387
rect 372 1384 407 1386
rect 372 1383 373 1384
rect 367 1382 373 1383
rect 406 1383 407 1384
rect 411 1383 412 1387
rect 406 1382 412 1383
rect 415 1387 421 1388
rect 415 1383 416 1387
rect 420 1386 421 1387
rect 462 1387 468 1388
rect 462 1386 463 1387
rect 420 1384 463 1386
rect 420 1383 421 1384
rect 415 1382 421 1383
rect 462 1383 463 1384
rect 467 1383 468 1387
rect 462 1382 468 1383
rect 471 1387 477 1388
rect 471 1383 472 1387
rect 476 1386 477 1387
rect 518 1387 524 1388
rect 518 1386 519 1387
rect 476 1384 519 1386
rect 476 1383 477 1384
rect 471 1382 477 1383
rect 518 1383 519 1384
rect 523 1383 524 1387
rect 518 1382 524 1383
rect 527 1387 533 1388
rect 527 1383 528 1387
rect 532 1386 533 1387
rect 574 1387 580 1388
rect 574 1386 575 1387
rect 532 1384 575 1386
rect 532 1383 533 1384
rect 527 1382 533 1383
rect 574 1383 575 1384
rect 579 1383 580 1387
rect 574 1382 580 1383
rect 583 1387 589 1388
rect 583 1383 584 1387
rect 588 1386 589 1387
rect 630 1387 636 1388
rect 630 1386 631 1387
rect 588 1384 631 1386
rect 588 1383 589 1384
rect 583 1382 589 1383
rect 630 1383 631 1384
rect 635 1383 636 1387
rect 630 1382 636 1383
rect 647 1387 653 1388
rect 647 1383 648 1387
rect 652 1383 653 1387
rect 647 1382 653 1383
rect 655 1387 661 1388
rect 655 1383 656 1387
rect 660 1386 661 1387
rect 711 1387 717 1388
rect 711 1386 712 1387
rect 660 1384 712 1386
rect 660 1383 661 1384
rect 655 1382 661 1383
rect 711 1383 712 1384
rect 716 1383 717 1387
rect 711 1382 717 1383
rect 719 1387 725 1388
rect 719 1383 720 1387
rect 724 1386 725 1387
rect 775 1387 781 1388
rect 775 1386 776 1387
rect 724 1384 776 1386
rect 724 1383 725 1384
rect 719 1382 725 1383
rect 775 1383 776 1384
rect 780 1383 781 1387
rect 775 1382 781 1383
rect 783 1387 789 1388
rect 783 1383 784 1387
rect 788 1386 789 1387
rect 839 1387 845 1388
rect 839 1386 840 1387
rect 788 1384 840 1386
rect 788 1383 789 1384
rect 783 1382 789 1383
rect 839 1383 840 1384
rect 844 1383 845 1387
rect 839 1382 845 1383
rect 903 1387 909 1388
rect 903 1383 904 1387
rect 908 1386 909 1387
rect 966 1387 972 1388
rect 966 1386 967 1387
rect 908 1384 967 1386
rect 908 1383 909 1384
rect 903 1382 909 1383
rect 966 1383 967 1384
rect 971 1383 972 1387
rect 966 1382 972 1383
rect 975 1387 981 1388
rect 975 1383 976 1387
rect 980 1386 981 1387
rect 1038 1387 1044 1388
rect 1038 1386 1039 1387
rect 980 1384 1039 1386
rect 980 1383 981 1384
rect 975 1382 981 1383
rect 1038 1383 1039 1384
rect 1043 1383 1044 1387
rect 1038 1382 1044 1383
rect 1047 1387 1053 1388
rect 1047 1383 1048 1387
rect 1052 1383 1053 1387
rect 2322 1387 2328 1388
rect 2322 1386 2323 1387
rect 1047 1382 1053 1383
rect 1238 1384 1244 1385
rect 366 1379 372 1380
rect 366 1378 367 1379
rect 304 1376 367 1378
rect 366 1375 367 1376
rect 371 1375 372 1379
rect 648 1378 650 1382
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 2176 1384 2323 1386
rect 2176 1380 2178 1384
rect 2322 1383 2323 1384
rect 2327 1383 2328 1387
rect 2322 1382 2328 1383
rect 782 1379 788 1380
rect 1238 1379 1244 1380
rect 1327 1379 1333 1380
rect 782 1378 783 1379
rect 648 1376 783 1378
rect 366 1374 372 1375
rect 782 1375 783 1376
rect 787 1375 788 1379
rect 782 1374 788 1375
rect 1278 1376 1284 1377
rect 1278 1372 1279 1376
rect 1283 1372 1284 1376
rect 1327 1375 1328 1379
rect 1332 1378 1333 1379
rect 1350 1379 1356 1380
rect 1332 1376 1346 1378
rect 1332 1375 1333 1376
rect 1327 1374 1333 1375
rect 1278 1371 1284 1372
rect 1344 1370 1346 1376
rect 1350 1375 1351 1379
rect 1355 1378 1356 1379
rect 1367 1379 1373 1380
rect 1367 1378 1368 1379
rect 1355 1376 1368 1378
rect 1355 1375 1356 1376
rect 1350 1374 1356 1375
rect 1367 1375 1368 1376
rect 1372 1375 1373 1379
rect 1367 1374 1373 1375
rect 1375 1379 1381 1380
rect 1375 1375 1376 1379
rect 1380 1378 1381 1379
rect 1423 1379 1429 1380
rect 1423 1378 1424 1379
rect 1380 1376 1424 1378
rect 1380 1375 1381 1376
rect 1375 1374 1381 1375
rect 1423 1375 1424 1376
rect 1428 1375 1429 1379
rect 1423 1374 1429 1375
rect 1495 1379 1501 1380
rect 1495 1375 1496 1379
rect 1500 1378 1501 1379
rect 1574 1379 1581 1380
rect 1500 1376 1570 1378
rect 1500 1375 1501 1376
rect 1495 1374 1501 1375
rect 1494 1371 1500 1372
rect 1494 1370 1495 1371
rect 1344 1368 1495 1370
rect 1494 1367 1495 1368
rect 1499 1367 1500 1371
rect 1568 1370 1570 1376
rect 1574 1375 1575 1379
rect 1580 1375 1581 1379
rect 1574 1374 1581 1375
rect 1583 1379 1589 1380
rect 1583 1375 1584 1379
rect 1588 1378 1589 1379
rect 1663 1379 1669 1380
rect 1663 1378 1664 1379
rect 1588 1376 1664 1378
rect 1588 1375 1589 1376
rect 1583 1374 1589 1375
rect 1663 1375 1664 1376
rect 1668 1375 1669 1379
rect 1663 1374 1669 1375
rect 1671 1379 1677 1380
rect 1671 1375 1672 1379
rect 1676 1378 1677 1379
rect 1751 1379 1757 1380
rect 1751 1378 1752 1379
rect 1676 1376 1752 1378
rect 1676 1375 1677 1376
rect 1671 1374 1677 1375
rect 1751 1375 1752 1376
rect 1756 1375 1757 1379
rect 1751 1374 1757 1375
rect 1839 1379 1845 1380
rect 1839 1375 1840 1379
rect 1844 1378 1845 1379
rect 1926 1379 1933 1380
rect 1844 1376 1922 1378
rect 1844 1375 1845 1376
rect 1839 1374 1845 1375
rect 1746 1371 1752 1372
rect 1746 1370 1747 1371
rect 1568 1368 1747 1370
rect 1494 1366 1500 1367
rect 1746 1367 1747 1368
rect 1751 1367 1752 1371
rect 1920 1370 1922 1376
rect 1926 1375 1927 1379
rect 1932 1375 1933 1379
rect 1926 1374 1933 1375
rect 1935 1379 1941 1380
rect 1935 1375 1936 1379
rect 1940 1378 1941 1379
rect 2015 1379 2021 1380
rect 2015 1378 2016 1379
rect 1940 1376 2016 1378
rect 1940 1375 1941 1376
rect 1935 1374 1941 1375
rect 2015 1375 2016 1376
rect 2020 1375 2021 1379
rect 2015 1374 2021 1375
rect 2023 1379 2029 1380
rect 2023 1375 2024 1379
rect 2028 1378 2029 1379
rect 2095 1379 2101 1380
rect 2095 1378 2096 1379
rect 2028 1376 2096 1378
rect 2028 1375 2029 1376
rect 2023 1374 2029 1375
rect 2095 1375 2096 1376
rect 2100 1375 2101 1379
rect 2095 1374 2101 1375
rect 2175 1379 2181 1380
rect 2175 1375 2176 1379
rect 2180 1375 2181 1379
rect 2175 1374 2181 1375
rect 2183 1379 2189 1380
rect 2183 1375 2184 1379
rect 2188 1378 2189 1379
rect 2247 1379 2253 1380
rect 2247 1378 2248 1379
rect 2188 1376 2248 1378
rect 2188 1375 2189 1376
rect 2183 1374 2189 1375
rect 2247 1375 2248 1376
rect 2252 1375 2253 1379
rect 2247 1374 2253 1375
rect 2327 1379 2333 1380
rect 2327 1375 2328 1379
rect 2332 1378 2333 1379
rect 2374 1379 2380 1380
rect 2374 1378 2375 1379
rect 2332 1376 2375 1378
rect 2332 1375 2333 1376
rect 2327 1374 2333 1375
rect 2374 1375 2375 1376
rect 2379 1375 2380 1379
rect 2374 1374 2380 1375
rect 2382 1379 2389 1380
rect 2382 1375 2383 1379
rect 2388 1375 2389 1379
rect 2382 1374 2389 1375
rect 2406 1376 2412 1377
rect 2406 1372 2407 1376
rect 2411 1372 2412 1376
rect 2190 1371 2196 1372
rect 2406 1371 2412 1372
rect 2190 1370 2191 1371
rect 1920 1368 2191 1370
rect 1746 1366 1752 1367
rect 2190 1367 2191 1368
rect 2195 1367 2196 1371
rect 2190 1366 2196 1367
rect 262 1361 268 1362
rect 262 1357 263 1361
rect 267 1357 268 1361
rect 262 1356 268 1357
rect 302 1361 308 1362
rect 302 1357 303 1361
rect 307 1357 308 1361
rect 302 1356 308 1357
rect 342 1361 348 1362
rect 342 1357 343 1361
rect 347 1357 348 1361
rect 342 1356 348 1357
rect 390 1361 396 1362
rect 390 1357 391 1361
rect 395 1357 396 1361
rect 390 1356 396 1357
rect 446 1361 452 1362
rect 446 1357 447 1361
rect 451 1357 452 1361
rect 446 1356 452 1357
rect 502 1361 508 1362
rect 502 1357 503 1361
rect 507 1357 508 1361
rect 502 1356 508 1357
rect 558 1361 564 1362
rect 558 1357 559 1361
rect 563 1357 564 1361
rect 558 1356 564 1357
rect 622 1361 628 1362
rect 622 1357 623 1361
rect 627 1357 628 1361
rect 622 1356 628 1357
rect 686 1361 692 1362
rect 686 1357 687 1361
rect 691 1357 692 1361
rect 686 1356 692 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 814 1361 820 1362
rect 814 1357 815 1361
rect 819 1357 820 1361
rect 814 1356 820 1357
rect 878 1361 884 1362
rect 878 1357 879 1361
rect 883 1357 884 1361
rect 878 1356 884 1357
rect 950 1361 956 1362
rect 950 1357 951 1361
rect 955 1357 956 1361
rect 950 1356 956 1357
rect 1022 1361 1028 1362
rect 1022 1357 1023 1361
rect 1027 1357 1028 1361
rect 1022 1356 1028 1357
rect 287 1355 293 1356
rect 287 1351 288 1355
rect 292 1354 293 1355
rect 310 1355 316 1356
rect 310 1354 311 1355
rect 292 1352 311 1354
rect 292 1351 293 1352
rect 287 1350 293 1351
rect 310 1351 311 1352
rect 315 1351 316 1355
rect 310 1350 316 1351
rect 327 1355 333 1356
rect 327 1351 328 1355
rect 332 1354 333 1355
rect 350 1355 356 1356
rect 350 1354 351 1355
rect 332 1352 351 1354
rect 332 1351 333 1352
rect 327 1350 333 1351
rect 350 1351 351 1352
rect 355 1351 356 1355
rect 350 1350 356 1351
rect 366 1355 373 1356
rect 366 1351 367 1355
rect 372 1351 373 1355
rect 366 1350 373 1351
rect 406 1355 412 1356
rect 406 1351 407 1355
rect 411 1354 412 1355
rect 415 1355 421 1356
rect 415 1354 416 1355
rect 411 1352 416 1354
rect 411 1351 412 1352
rect 406 1350 412 1351
rect 415 1351 416 1352
rect 420 1351 421 1355
rect 415 1350 421 1351
rect 462 1355 468 1356
rect 462 1351 463 1355
rect 467 1354 468 1355
rect 471 1355 477 1356
rect 471 1354 472 1355
rect 467 1352 472 1354
rect 467 1351 468 1352
rect 462 1350 468 1351
rect 471 1351 472 1352
rect 476 1351 477 1355
rect 471 1350 477 1351
rect 518 1355 524 1356
rect 518 1351 519 1355
rect 523 1354 524 1355
rect 527 1355 533 1356
rect 527 1354 528 1355
rect 523 1352 528 1354
rect 523 1351 524 1352
rect 518 1350 524 1351
rect 527 1351 528 1352
rect 532 1351 533 1355
rect 527 1350 533 1351
rect 574 1355 580 1356
rect 574 1351 575 1355
rect 579 1354 580 1355
rect 583 1355 589 1356
rect 583 1354 584 1355
rect 579 1352 584 1354
rect 579 1351 580 1352
rect 574 1350 580 1351
rect 583 1351 584 1352
rect 588 1351 589 1355
rect 583 1350 589 1351
rect 647 1355 653 1356
rect 647 1351 648 1355
rect 652 1354 653 1355
rect 655 1355 661 1356
rect 655 1354 656 1355
rect 652 1352 656 1354
rect 652 1351 653 1352
rect 647 1350 653 1351
rect 655 1351 656 1352
rect 660 1351 661 1355
rect 655 1350 661 1351
rect 711 1355 717 1356
rect 711 1351 712 1355
rect 716 1354 717 1355
rect 719 1355 725 1356
rect 719 1354 720 1355
rect 716 1352 720 1354
rect 716 1351 717 1352
rect 711 1350 717 1351
rect 719 1351 720 1352
rect 724 1351 725 1355
rect 719 1350 725 1351
rect 775 1355 781 1356
rect 775 1351 776 1355
rect 780 1354 781 1355
rect 783 1355 789 1356
rect 783 1354 784 1355
rect 780 1352 784 1354
rect 780 1351 781 1352
rect 775 1350 781 1351
rect 783 1351 784 1352
rect 788 1351 789 1355
rect 783 1350 789 1351
rect 838 1355 845 1356
rect 838 1351 839 1355
rect 844 1351 845 1355
rect 838 1350 845 1351
rect 866 1355 872 1356
rect 866 1351 867 1355
rect 871 1354 872 1355
rect 903 1355 909 1356
rect 903 1354 904 1355
rect 871 1352 904 1354
rect 871 1351 872 1352
rect 866 1350 872 1351
rect 903 1351 904 1352
rect 908 1351 909 1355
rect 903 1350 909 1351
rect 966 1355 972 1356
rect 966 1351 967 1355
rect 971 1354 972 1355
rect 975 1355 981 1356
rect 975 1354 976 1355
rect 971 1352 976 1354
rect 971 1351 972 1352
rect 966 1350 972 1351
rect 975 1351 976 1352
rect 980 1351 981 1355
rect 975 1350 981 1351
rect 1038 1355 1044 1356
rect 1038 1351 1039 1355
rect 1043 1354 1044 1355
rect 1047 1355 1053 1356
rect 1047 1354 1048 1355
rect 1043 1352 1048 1354
rect 1043 1351 1044 1352
rect 1038 1350 1044 1351
rect 1047 1351 1048 1352
rect 1052 1351 1053 1355
rect 1926 1355 1932 1356
rect 1926 1354 1927 1355
rect 1047 1350 1053 1351
rect 1302 1353 1308 1354
rect 1302 1349 1303 1353
rect 1307 1349 1308 1353
rect 1302 1348 1308 1349
rect 1342 1353 1348 1354
rect 1342 1349 1343 1353
rect 1347 1349 1348 1353
rect 1342 1348 1348 1349
rect 1398 1353 1404 1354
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1470 1353 1476 1354
rect 1470 1349 1471 1353
rect 1475 1349 1476 1353
rect 1470 1348 1476 1349
rect 1550 1353 1556 1354
rect 1550 1349 1551 1353
rect 1555 1349 1556 1353
rect 1550 1348 1556 1349
rect 1638 1353 1644 1354
rect 1638 1349 1639 1353
rect 1643 1349 1644 1353
rect 1638 1348 1644 1349
rect 1726 1353 1732 1354
rect 1726 1349 1727 1353
rect 1731 1349 1732 1353
rect 1726 1348 1732 1349
rect 1814 1353 1820 1354
rect 1814 1349 1815 1353
rect 1819 1349 1820 1353
rect 1814 1348 1820 1349
rect 1902 1353 1908 1354
rect 1902 1349 1903 1353
rect 1907 1349 1908 1353
rect 1902 1348 1908 1349
rect 1912 1352 1927 1354
rect 1327 1347 1333 1348
rect 1327 1343 1328 1347
rect 1332 1346 1333 1347
rect 1350 1347 1356 1348
rect 1350 1346 1351 1347
rect 1332 1344 1351 1346
rect 1332 1343 1333 1344
rect 1327 1342 1333 1343
rect 1350 1343 1351 1344
rect 1355 1343 1356 1347
rect 1350 1342 1356 1343
rect 1367 1347 1373 1348
rect 1367 1343 1368 1347
rect 1372 1346 1373 1347
rect 1375 1347 1381 1348
rect 1375 1346 1376 1347
rect 1372 1344 1376 1346
rect 1372 1343 1373 1344
rect 1367 1342 1373 1343
rect 1375 1343 1376 1344
rect 1380 1343 1381 1347
rect 1375 1342 1381 1343
rect 1423 1347 1429 1348
rect 1423 1343 1424 1347
rect 1428 1346 1429 1347
rect 1458 1347 1464 1348
rect 1458 1346 1459 1347
rect 1428 1344 1459 1346
rect 1428 1343 1429 1344
rect 1423 1342 1429 1343
rect 1458 1343 1459 1344
rect 1463 1343 1464 1347
rect 1458 1342 1464 1343
rect 1494 1347 1501 1348
rect 1494 1343 1495 1347
rect 1500 1343 1501 1347
rect 1494 1342 1501 1343
rect 1575 1347 1581 1348
rect 1575 1343 1576 1347
rect 1580 1346 1581 1347
rect 1583 1347 1589 1348
rect 1583 1346 1584 1347
rect 1580 1344 1584 1346
rect 1580 1343 1581 1344
rect 1575 1342 1581 1343
rect 1583 1343 1584 1344
rect 1588 1343 1589 1347
rect 1583 1342 1589 1343
rect 1663 1347 1669 1348
rect 1663 1343 1664 1347
rect 1668 1346 1669 1347
rect 1671 1347 1677 1348
rect 1671 1346 1672 1347
rect 1668 1344 1672 1346
rect 1668 1343 1669 1344
rect 1663 1342 1669 1343
rect 1671 1343 1672 1344
rect 1676 1343 1677 1347
rect 1671 1342 1677 1343
rect 1746 1347 1757 1348
rect 1746 1343 1747 1347
rect 1751 1343 1752 1347
rect 1756 1343 1757 1347
rect 1746 1342 1757 1343
rect 1839 1347 1845 1348
rect 1839 1343 1840 1347
rect 1844 1346 1845 1347
rect 1912 1346 1914 1352
rect 1926 1351 1927 1352
rect 1931 1351 1932 1355
rect 1926 1350 1932 1351
rect 1990 1353 1996 1354
rect 1990 1349 1991 1353
rect 1995 1349 1996 1353
rect 1990 1348 1996 1349
rect 2070 1353 2076 1354
rect 2070 1349 2071 1353
rect 2075 1349 2076 1353
rect 2070 1348 2076 1349
rect 2150 1353 2156 1354
rect 2150 1349 2151 1353
rect 2155 1349 2156 1353
rect 2150 1348 2156 1349
rect 2222 1353 2228 1354
rect 2222 1349 2223 1353
rect 2227 1349 2228 1353
rect 2222 1348 2228 1349
rect 2302 1353 2308 1354
rect 2302 1349 2303 1353
rect 2307 1349 2308 1353
rect 2302 1348 2308 1349
rect 2358 1353 2364 1354
rect 2358 1349 2359 1353
rect 2363 1349 2364 1353
rect 2358 1348 2364 1349
rect 1844 1344 1914 1346
rect 1927 1347 1933 1348
rect 1844 1343 1845 1344
rect 1839 1342 1845 1343
rect 1927 1343 1928 1347
rect 1932 1346 1933 1347
rect 1935 1347 1941 1348
rect 1935 1346 1936 1347
rect 1932 1344 1936 1346
rect 1932 1343 1933 1344
rect 1927 1342 1933 1343
rect 1935 1343 1936 1344
rect 1940 1343 1941 1347
rect 1935 1342 1941 1343
rect 2015 1347 2021 1348
rect 2015 1343 2016 1347
rect 2020 1346 2021 1347
rect 2023 1347 2029 1348
rect 2023 1346 2024 1347
rect 2020 1344 2024 1346
rect 2020 1343 2021 1344
rect 2015 1342 2021 1343
rect 2023 1343 2024 1344
rect 2028 1343 2029 1347
rect 2023 1342 2029 1343
rect 2094 1347 2101 1348
rect 2094 1343 2095 1347
rect 2100 1343 2101 1347
rect 2094 1342 2101 1343
rect 2175 1347 2181 1348
rect 2175 1343 2176 1347
rect 2180 1346 2181 1347
rect 2183 1347 2189 1348
rect 2183 1346 2184 1347
rect 2180 1344 2184 1346
rect 2180 1343 2181 1344
rect 2175 1342 2181 1343
rect 2183 1343 2184 1344
rect 2188 1343 2189 1347
rect 2183 1342 2189 1343
rect 2247 1347 2253 1348
rect 2247 1343 2248 1347
rect 2252 1346 2253 1347
rect 2294 1347 2300 1348
rect 2294 1346 2295 1347
rect 2252 1344 2295 1346
rect 2252 1343 2253 1344
rect 2247 1342 2253 1343
rect 2294 1343 2295 1344
rect 2299 1343 2300 1347
rect 2294 1342 2300 1343
rect 2327 1347 2333 1348
rect 2327 1343 2328 1347
rect 2332 1346 2333 1347
rect 2343 1347 2349 1348
rect 2343 1346 2344 1347
rect 2332 1344 2344 1346
rect 2332 1343 2333 1344
rect 2327 1342 2333 1343
rect 2343 1343 2344 1344
rect 2348 1343 2349 1347
rect 2343 1342 2349 1343
rect 2374 1347 2380 1348
rect 2374 1343 2375 1347
rect 2379 1346 2380 1347
rect 2383 1347 2389 1348
rect 2383 1346 2384 1347
rect 2379 1344 2384 1346
rect 2379 1343 2380 1344
rect 2374 1342 2380 1343
rect 2383 1343 2384 1344
rect 2388 1343 2389 1347
rect 2383 1342 2389 1343
rect 190 1335 196 1336
rect 190 1334 191 1335
rect 161 1332 191 1334
rect 159 1331 165 1332
rect 134 1327 140 1328
rect 134 1323 135 1327
rect 139 1323 140 1327
rect 159 1327 160 1331
rect 164 1327 165 1331
rect 190 1331 191 1332
rect 195 1331 196 1335
rect 190 1330 196 1331
rect 199 1331 208 1332
rect 159 1326 165 1327
rect 174 1327 180 1328
rect 134 1322 140 1323
rect 174 1323 175 1327
rect 179 1323 180 1327
rect 199 1327 200 1331
rect 207 1327 208 1331
rect 238 1331 245 1332
rect 199 1326 208 1327
rect 214 1327 220 1328
rect 174 1322 180 1323
rect 214 1323 215 1327
rect 219 1323 220 1327
rect 238 1327 239 1331
rect 244 1327 245 1331
rect 279 1331 285 1332
rect 279 1330 280 1331
rect 264 1328 280 1330
rect 238 1326 245 1327
rect 254 1327 260 1328
rect 214 1322 220 1323
rect 254 1323 255 1327
rect 259 1323 260 1327
rect 254 1322 260 1323
rect 162 1319 168 1320
rect 162 1315 163 1319
rect 167 1318 168 1319
rect 264 1318 266 1328
rect 279 1327 280 1328
rect 284 1327 285 1331
rect 351 1331 357 1332
rect 279 1326 285 1327
rect 326 1327 332 1328
rect 326 1323 327 1327
rect 331 1323 332 1327
rect 351 1327 352 1331
rect 356 1330 357 1331
rect 398 1331 404 1332
rect 398 1330 399 1331
rect 356 1328 399 1330
rect 356 1327 357 1328
rect 351 1326 357 1327
rect 398 1327 399 1328
rect 403 1327 404 1331
rect 431 1331 437 1332
rect 398 1326 404 1327
rect 406 1327 412 1328
rect 326 1322 332 1323
rect 406 1323 407 1327
rect 411 1323 412 1327
rect 431 1327 432 1331
rect 436 1330 437 1331
rect 486 1331 492 1332
rect 486 1330 487 1331
rect 436 1328 487 1330
rect 436 1327 437 1328
rect 431 1326 437 1327
rect 486 1327 487 1328
rect 491 1327 492 1331
rect 506 1331 512 1332
rect 486 1326 492 1327
rect 494 1327 500 1328
rect 406 1322 412 1323
rect 494 1323 495 1327
rect 499 1323 500 1327
rect 506 1327 507 1331
rect 511 1330 512 1331
rect 519 1331 525 1332
rect 519 1330 520 1331
rect 511 1328 520 1330
rect 511 1327 512 1328
rect 506 1326 512 1327
rect 519 1327 520 1328
rect 524 1327 525 1331
rect 607 1331 613 1332
rect 519 1326 525 1327
rect 582 1327 588 1328
rect 494 1322 500 1323
rect 582 1323 583 1327
rect 587 1323 588 1327
rect 607 1327 608 1331
rect 612 1330 613 1331
rect 662 1331 668 1332
rect 662 1330 663 1331
rect 612 1328 663 1330
rect 612 1327 613 1328
rect 607 1326 613 1327
rect 662 1327 663 1328
rect 667 1327 668 1331
rect 695 1331 701 1332
rect 662 1326 668 1327
rect 670 1327 676 1328
rect 582 1322 588 1323
rect 670 1323 671 1327
rect 675 1323 676 1327
rect 695 1327 696 1331
rect 700 1330 701 1331
rect 750 1331 756 1332
rect 750 1330 751 1331
rect 700 1328 751 1330
rect 700 1327 701 1328
rect 695 1326 701 1327
rect 750 1327 751 1328
rect 755 1327 756 1331
rect 782 1331 789 1332
rect 750 1326 756 1327
rect 758 1327 764 1328
rect 670 1322 676 1323
rect 758 1323 759 1327
rect 763 1323 764 1327
rect 782 1327 783 1331
rect 788 1327 789 1331
rect 863 1331 869 1332
rect 782 1326 789 1327
rect 838 1327 844 1328
rect 758 1322 764 1323
rect 838 1323 839 1327
rect 843 1323 844 1327
rect 863 1327 864 1331
rect 868 1330 869 1331
rect 910 1331 916 1332
rect 910 1330 911 1331
rect 868 1328 911 1330
rect 868 1327 869 1328
rect 863 1326 869 1327
rect 910 1327 911 1328
rect 915 1327 916 1331
rect 943 1331 949 1332
rect 910 1326 916 1327
rect 918 1327 924 1328
rect 838 1322 844 1323
rect 918 1323 919 1327
rect 923 1323 924 1327
rect 943 1327 944 1331
rect 948 1330 949 1331
rect 998 1331 1004 1332
rect 998 1330 999 1331
rect 948 1328 999 1330
rect 948 1327 949 1328
rect 943 1326 949 1327
rect 998 1327 999 1328
rect 1003 1327 1004 1331
rect 1031 1331 1037 1332
rect 998 1326 1004 1327
rect 1006 1327 1012 1328
rect 918 1322 924 1323
rect 1006 1323 1007 1327
rect 1011 1323 1012 1327
rect 1031 1327 1032 1331
rect 1036 1330 1037 1331
rect 1086 1331 1092 1332
rect 1086 1330 1087 1331
rect 1036 1328 1087 1330
rect 1036 1327 1037 1328
rect 1031 1326 1037 1327
rect 1086 1327 1087 1328
rect 1091 1327 1092 1331
rect 1106 1331 1112 1332
rect 1086 1326 1092 1327
rect 1094 1327 1100 1328
rect 1006 1322 1012 1323
rect 1094 1323 1095 1327
rect 1099 1323 1100 1327
rect 1106 1327 1107 1331
rect 1111 1330 1112 1331
rect 1119 1331 1125 1332
rect 1119 1330 1120 1331
rect 1111 1328 1120 1330
rect 1111 1327 1112 1328
rect 1106 1326 1112 1327
rect 1119 1327 1120 1328
rect 1124 1327 1125 1331
rect 1119 1326 1125 1327
rect 1502 1327 1508 1328
rect 1502 1326 1503 1327
rect 1480 1324 1503 1326
rect 1094 1322 1100 1323
rect 1471 1323 1477 1324
rect 167 1316 266 1318
rect 1446 1319 1452 1320
rect 167 1315 168 1316
rect 162 1314 168 1315
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1471 1319 1472 1323
rect 1476 1322 1477 1323
rect 1480 1322 1482 1324
rect 1502 1323 1503 1324
rect 1507 1323 1508 1327
rect 1542 1327 1548 1328
rect 1542 1326 1543 1327
rect 1520 1324 1543 1326
rect 1502 1322 1508 1323
rect 1511 1323 1517 1324
rect 1476 1320 1482 1322
rect 1476 1319 1477 1320
rect 1471 1318 1477 1319
rect 1486 1319 1492 1320
rect 1446 1314 1452 1315
rect 1486 1315 1487 1319
rect 1491 1315 1492 1319
rect 1511 1319 1512 1323
rect 1516 1322 1517 1323
rect 1520 1322 1522 1324
rect 1542 1323 1543 1324
rect 1547 1323 1548 1327
rect 1574 1327 1580 1328
rect 1574 1326 1575 1327
rect 1542 1322 1548 1323
rect 1551 1325 1575 1326
rect 1516 1320 1522 1322
rect 1551 1321 1552 1325
rect 1556 1324 1575 1325
rect 1556 1321 1557 1324
rect 1574 1323 1575 1324
rect 1579 1323 1580 1327
rect 1574 1322 1580 1323
rect 1582 1323 1588 1324
rect 1551 1320 1557 1321
rect 1516 1319 1517 1320
rect 1511 1318 1517 1319
rect 1526 1319 1532 1320
rect 1486 1314 1492 1315
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1566 1319 1572 1320
rect 1566 1315 1567 1319
rect 1571 1315 1572 1319
rect 1582 1319 1583 1323
rect 1587 1322 1588 1323
rect 1591 1323 1597 1324
rect 1591 1322 1592 1323
rect 1587 1320 1592 1322
rect 1587 1319 1588 1320
rect 1582 1318 1588 1319
rect 1591 1319 1592 1320
rect 1596 1319 1597 1323
rect 1639 1323 1645 1324
rect 1591 1318 1597 1319
rect 1614 1319 1620 1320
rect 1566 1314 1572 1315
rect 1614 1315 1615 1319
rect 1619 1315 1620 1319
rect 1639 1319 1640 1323
rect 1644 1322 1645 1323
rect 1662 1323 1668 1324
rect 1662 1322 1663 1323
rect 1644 1320 1663 1322
rect 1644 1319 1645 1320
rect 1639 1318 1645 1319
rect 1662 1319 1663 1320
rect 1667 1319 1668 1323
rect 1695 1323 1701 1324
rect 1662 1318 1668 1319
rect 1670 1319 1676 1320
rect 1614 1314 1620 1315
rect 1670 1315 1671 1319
rect 1675 1315 1676 1319
rect 1695 1319 1696 1323
rect 1700 1322 1701 1323
rect 1710 1323 1716 1324
rect 1710 1322 1711 1323
rect 1700 1320 1711 1322
rect 1700 1319 1701 1320
rect 1695 1318 1701 1319
rect 1710 1319 1711 1320
rect 1715 1319 1716 1323
rect 1730 1323 1736 1324
rect 1710 1318 1716 1319
rect 1718 1319 1724 1320
rect 1670 1314 1676 1315
rect 1718 1315 1719 1319
rect 1723 1315 1724 1319
rect 1730 1319 1731 1323
rect 1735 1322 1736 1323
rect 1743 1323 1749 1324
rect 1743 1322 1744 1323
rect 1735 1320 1744 1322
rect 1735 1319 1736 1320
rect 1730 1318 1736 1319
rect 1743 1319 1744 1320
rect 1748 1319 1749 1323
rect 1799 1323 1805 1324
rect 1743 1318 1749 1319
rect 1774 1319 1780 1320
rect 1718 1314 1724 1315
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1799 1319 1800 1323
rect 1804 1322 1805 1323
rect 1822 1323 1828 1324
rect 1822 1322 1823 1323
rect 1804 1320 1823 1322
rect 1804 1319 1805 1320
rect 1799 1318 1805 1319
rect 1822 1319 1823 1320
rect 1827 1319 1828 1323
rect 1855 1323 1861 1324
rect 1822 1318 1828 1319
rect 1830 1319 1836 1320
rect 1774 1314 1780 1315
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1855 1319 1856 1323
rect 1860 1322 1861 1323
rect 1894 1323 1900 1324
rect 1894 1322 1895 1323
rect 1860 1320 1895 1322
rect 1860 1319 1861 1320
rect 1855 1318 1861 1319
rect 1894 1319 1895 1320
rect 1899 1319 1900 1323
rect 1927 1323 1933 1324
rect 1894 1318 1900 1319
rect 1902 1319 1908 1320
rect 1830 1314 1836 1315
rect 1902 1315 1903 1319
rect 1907 1315 1908 1319
rect 1927 1319 1928 1323
rect 1932 1322 1933 1323
rect 1962 1323 1968 1324
rect 1962 1322 1963 1323
rect 1932 1320 1963 1322
rect 1932 1319 1933 1320
rect 1927 1318 1933 1319
rect 1962 1319 1963 1320
rect 1967 1319 1968 1323
rect 2007 1323 2013 1324
rect 1962 1318 1968 1319
rect 1982 1319 1988 1320
rect 1902 1314 1908 1315
rect 1982 1315 1983 1319
rect 1987 1315 1988 1319
rect 2007 1319 2008 1323
rect 2012 1322 2013 1323
rect 2062 1323 2068 1324
rect 2062 1322 2063 1323
rect 2012 1320 2063 1322
rect 2012 1319 2013 1320
rect 2007 1318 2013 1319
rect 2062 1319 2063 1320
rect 2067 1319 2068 1323
rect 2095 1323 2101 1324
rect 2062 1318 2068 1319
rect 2070 1319 2076 1320
rect 1982 1314 1988 1315
rect 2070 1315 2071 1319
rect 2075 1315 2076 1319
rect 2095 1319 2096 1323
rect 2100 1322 2101 1323
rect 2158 1323 2164 1324
rect 2158 1322 2159 1323
rect 2100 1320 2159 1322
rect 2100 1319 2101 1320
rect 2095 1318 2101 1319
rect 2158 1319 2159 1320
rect 2163 1319 2164 1323
rect 2190 1323 2197 1324
rect 2158 1318 2164 1319
rect 2166 1319 2172 1320
rect 2070 1314 2076 1315
rect 2166 1315 2167 1319
rect 2171 1315 2172 1319
rect 2190 1319 2191 1323
rect 2196 1319 2197 1323
rect 2282 1323 2288 1324
rect 2190 1318 2197 1319
rect 2270 1319 2276 1320
rect 2166 1314 2172 1315
rect 2270 1315 2271 1319
rect 2275 1315 2276 1319
rect 2282 1319 2283 1323
rect 2287 1322 2288 1323
rect 2295 1323 2301 1324
rect 2295 1322 2296 1323
rect 2287 1320 2296 1322
rect 2287 1319 2288 1320
rect 2282 1318 2288 1319
rect 2295 1319 2296 1320
rect 2300 1319 2301 1323
rect 2382 1323 2389 1324
rect 2295 1318 2301 1319
rect 2358 1319 2364 1320
rect 2270 1314 2276 1315
rect 2358 1315 2359 1319
rect 2363 1315 2364 1319
rect 2382 1319 2383 1323
rect 2388 1319 2389 1323
rect 2382 1318 2389 1319
rect 2358 1314 2364 1315
rect 202 1307 208 1308
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 202 1303 203 1307
rect 207 1306 208 1307
rect 506 1307 512 1308
rect 506 1306 507 1307
rect 207 1304 243 1306
rect 207 1303 208 1304
rect 202 1302 208 1303
rect 241 1300 243 1304
rect 319 1304 507 1306
rect 110 1299 116 1300
rect 159 1299 168 1300
rect 159 1295 160 1299
rect 167 1295 168 1299
rect 159 1294 168 1295
rect 190 1299 196 1300
rect 190 1295 191 1299
rect 195 1298 196 1299
rect 199 1299 205 1300
rect 199 1298 200 1299
rect 195 1296 200 1298
rect 195 1295 196 1296
rect 190 1294 196 1295
rect 199 1295 200 1296
rect 204 1295 205 1299
rect 199 1294 205 1295
rect 239 1299 245 1300
rect 239 1295 240 1299
rect 244 1295 245 1299
rect 239 1294 245 1295
rect 279 1299 285 1300
rect 279 1295 280 1299
rect 284 1298 285 1299
rect 319 1298 321 1304
rect 506 1303 507 1304
rect 511 1303 512 1307
rect 506 1302 512 1303
rect 1238 1304 1244 1305
rect 1238 1300 1239 1304
rect 1243 1300 1244 1304
rect 284 1296 321 1298
rect 350 1299 357 1300
rect 284 1295 285 1296
rect 279 1294 285 1295
rect 350 1295 351 1299
rect 356 1295 357 1299
rect 350 1294 357 1295
rect 398 1299 404 1300
rect 398 1295 399 1299
rect 403 1298 404 1299
rect 431 1299 437 1300
rect 431 1298 432 1299
rect 403 1296 432 1298
rect 403 1295 404 1296
rect 398 1294 404 1295
rect 431 1295 432 1296
rect 436 1295 437 1299
rect 431 1294 437 1295
rect 486 1299 492 1300
rect 486 1295 487 1299
rect 491 1298 492 1299
rect 519 1299 525 1300
rect 519 1298 520 1299
rect 491 1296 520 1298
rect 491 1295 492 1296
rect 486 1294 492 1295
rect 519 1295 520 1296
rect 524 1295 525 1299
rect 519 1294 525 1295
rect 542 1299 548 1300
rect 542 1295 543 1299
rect 547 1298 548 1299
rect 607 1299 613 1300
rect 607 1298 608 1299
rect 547 1296 608 1298
rect 547 1295 548 1296
rect 542 1294 548 1295
rect 607 1295 608 1296
rect 612 1295 613 1299
rect 607 1294 613 1295
rect 662 1299 668 1300
rect 662 1295 663 1299
rect 667 1298 668 1299
rect 695 1299 701 1300
rect 695 1298 696 1299
rect 667 1296 696 1298
rect 667 1295 668 1296
rect 662 1294 668 1295
rect 695 1295 696 1296
rect 700 1295 701 1299
rect 695 1294 701 1295
rect 750 1299 756 1300
rect 750 1295 751 1299
rect 755 1298 756 1299
rect 783 1299 789 1300
rect 783 1298 784 1299
rect 755 1296 784 1298
rect 755 1295 756 1296
rect 750 1294 756 1295
rect 783 1295 784 1296
rect 788 1295 789 1299
rect 783 1294 789 1295
rect 863 1299 872 1300
rect 863 1295 864 1299
rect 871 1295 872 1299
rect 863 1294 872 1295
rect 910 1299 916 1300
rect 910 1295 911 1299
rect 915 1298 916 1299
rect 943 1299 949 1300
rect 943 1298 944 1299
rect 915 1296 944 1298
rect 915 1295 916 1296
rect 910 1294 916 1295
rect 943 1295 944 1296
rect 948 1295 949 1299
rect 943 1294 949 1295
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1298 1004 1299
rect 1031 1299 1037 1300
rect 1031 1298 1032 1299
rect 1003 1296 1032 1298
rect 1003 1295 1004 1296
rect 998 1294 1004 1295
rect 1031 1295 1032 1296
rect 1036 1295 1037 1299
rect 1031 1294 1037 1295
rect 1086 1299 1092 1300
rect 1086 1295 1087 1299
rect 1091 1298 1092 1299
rect 1119 1299 1125 1300
rect 1238 1299 1244 1300
rect 1582 1299 1588 1300
rect 1119 1298 1120 1299
rect 1091 1296 1120 1298
rect 1091 1295 1092 1296
rect 1086 1294 1092 1295
rect 1119 1295 1120 1296
rect 1124 1295 1125 1299
rect 1582 1298 1583 1299
rect 1119 1294 1125 1295
rect 1278 1296 1284 1297
rect 1278 1292 1279 1296
rect 1283 1292 1284 1296
rect 1496 1296 1583 1298
rect 1278 1291 1284 1292
rect 1471 1291 1477 1292
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 1238 1287 1244 1288
rect 1238 1283 1239 1287
rect 1243 1283 1244 1287
rect 1471 1287 1472 1291
rect 1476 1290 1477 1291
rect 1496 1290 1498 1296
rect 1582 1295 1583 1296
rect 1587 1295 1588 1299
rect 1730 1299 1736 1300
rect 1730 1298 1731 1299
rect 1582 1294 1588 1295
rect 1616 1296 1731 1298
rect 1476 1288 1498 1290
rect 1502 1291 1508 1292
rect 1476 1287 1477 1288
rect 1471 1286 1477 1287
rect 1502 1287 1503 1291
rect 1507 1290 1508 1291
rect 1511 1291 1517 1292
rect 1511 1290 1512 1291
rect 1507 1288 1512 1290
rect 1507 1287 1508 1288
rect 1502 1286 1508 1287
rect 1511 1287 1512 1288
rect 1516 1287 1517 1291
rect 1511 1286 1517 1287
rect 1542 1291 1548 1292
rect 1542 1287 1543 1291
rect 1547 1290 1548 1291
rect 1551 1291 1557 1292
rect 1551 1290 1552 1291
rect 1547 1288 1552 1290
rect 1547 1287 1548 1288
rect 1542 1286 1548 1287
rect 1551 1287 1552 1288
rect 1556 1287 1557 1291
rect 1551 1286 1557 1287
rect 1591 1291 1597 1292
rect 1591 1287 1592 1291
rect 1596 1290 1597 1291
rect 1616 1290 1618 1296
rect 1730 1295 1731 1296
rect 1735 1295 1736 1299
rect 1730 1294 1736 1295
rect 2406 1296 2412 1297
rect 2406 1292 2407 1296
rect 2411 1292 2412 1296
rect 1596 1288 1618 1290
rect 1622 1291 1628 1292
rect 1596 1287 1597 1288
rect 1591 1286 1597 1287
rect 1622 1287 1623 1291
rect 1627 1290 1628 1291
rect 1639 1291 1645 1292
rect 1639 1290 1640 1291
rect 1627 1288 1640 1290
rect 1627 1287 1628 1288
rect 1622 1286 1628 1287
rect 1639 1287 1640 1288
rect 1644 1287 1645 1291
rect 1639 1286 1645 1287
rect 1662 1291 1668 1292
rect 1662 1287 1663 1291
rect 1667 1290 1668 1291
rect 1695 1291 1701 1292
rect 1695 1290 1696 1291
rect 1667 1288 1696 1290
rect 1667 1287 1668 1288
rect 1662 1286 1668 1287
rect 1695 1287 1696 1288
rect 1700 1287 1701 1291
rect 1695 1286 1701 1287
rect 1710 1291 1716 1292
rect 1710 1287 1711 1291
rect 1715 1290 1716 1291
rect 1743 1291 1749 1292
rect 1743 1290 1744 1291
rect 1715 1288 1744 1290
rect 1715 1287 1716 1288
rect 1710 1286 1716 1287
rect 1743 1287 1744 1288
rect 1748 1287 1749 1291
rect 1743 1286 1749 1287
rect 1799 1291 1805 1292
rect 1799 1287 1800 1291
rect 1804 1290 1805 1291
rect 1822 1291 1828 1292
rect 1804 1288 1818 1290
rect 1804 1287 1805 1288
rect 1799 1286 1805 1287
rect 1238 1282 1244 1283
rect 1816 1282 1818 1288
rect 1822 1287 1823 1291
rect 1827 1290 1828 1291
rect 1855 1291 1861 1292
rect 1855 1290 1856 1291
rect 1827 1288 1856 1290
rect 1827 1287 1828 1288
rect 1822 1286 1828 1287
rect 1855 1287 1856 1288
rect 1860 1287 1861 1291
rect 1855 1286 1861 1287
rect 1894 1291 1900 1292
rect 1894 1287 1895 1291
rect 1899 1290 1900 1291
rect 1927 1291 1933 1292
rect 1927 1290 1928 1291
rect 1899 1288 1928 1290
rect 1899 1287 1900 1288
rect 1894 1286 1900 1287
rect 1927 1287 1928 1288
rect 1932 1287 1933 1291
rect 1927 1286 1933 1287
rect 1962 1291 1968 1292
rect 1962 1287 1963 1291
rect 1967 1290 1968 1291
rect 2007 1291 2013 1292
rect 2007 1290 2008 1291
rect 1967 1288 2008 1290
rect 1967 1287 1968 1288
rect 1962 1286 1968 1287
rect 2007 1287 2008 1288
rect 2012 1287 2013 1291
rect 2007 1286 2013 1287
rect 2062 1291 2068 1292
rect 2062 1287 2063 1291
rect 2067 1290 2068 1291
rect 2095 1291 2101 1292
rect 2095 1290 2096 1291
rect 2067 1288 2096 1290
rect 2067 1287 2068 1288
rect 2062 1286 2068 1287
rect 2095 1287 2096 1288
rect 2100 1287 2101 1291
rect 2095 1286 2101 1287
rect 2158 1291 2164 1292
rect 2158 1287 2159 1291
rect 2163 1290 2164 1291
rect 2191 1291 2197 1292
rect 2191 1290 2192 1291
rect 2163 1288 2192 1290
rect 2163 1287 2164 1288
rect 2158 1286 2164 1287
rect 2191 1287 2192 1288
rect 2196 1287 2197 1291
rect 2191 1286 2197 1287
rect 2294 1291 2301 1292
rect 2294 1287 2295 1291
rect 2300 1287 2301 1291
rect 2294 1286 2301 1287
rect 2382 1291 2389 1292
rect 2406 1291 2412 1292
rect 2382 1287 2383 1291
rect 2388 1287 2389 1291
rect 2382 1286 2389 1287
rect 2142 1283 2148 1284
rect 2142 1282 2143 1283
rect 134 1280 140 1281
rect 134 1276 135 1280
rect 139 1276 140 1280
rect 134 1275 140 1276
rect 174 1280 180 1281
rect 174 1276 175 1280
rect 179 1276 180 1280
rect 174 1275 180 1276
rect 214 1280 220 1281
rect 214 1276 215 1280
rect 219 1276 220 1280
rect 214 1275 220 1276
rect 254 1280 260 1281
rect 254 1276 255 1280
rect 259 1276 260 1280
rect 254 1275 260 1276
rect 326 1280 332 1281
rect 326 1276 327 1280
rect 331 1276 332 1280
rect 326 1275 332 1276
rect 406 1280 412 1281
rect 406 1276 407 1280
rect 411 1276 412 1280
rect 406 1275 412 1276
rect 494 1280 500 1281
rect 494 1276 495 1280
rect 499 1276 500 1280
rect 494 1275 500 1276
rect 582 1280 588 1281
rect 582 1276 583 1280
rect 587 1276 588 1280
rect 582 1275 588 1276
rect 670 1280 676 1281
rect 670 1276 671 1280
rect 675 1276 676 1280
rect 670 1275 676 1276
rect 758 1280 764 1281
rect 758 1276 759 1280
rect 763 1276 764 1280
rect 758 1275 764 1276
rect 838 1280 844 1281
rect 838 1276 839 1280
rect 843 1276 844 1280
rect 838 1275 844 1276
rect 918 1280 924 1281
rect 918 1276 919 1280
rect 923 1276 924 1280
rect 918 1275 924 1276
rect 1006 1280 1012 1281
rect 1006 1276 1007 1280
rect 1011 1276 1012 1280
rect 1006 1275 1012 1276
rect 1094 1280 1100 1281
rect 1816 1280 2143 1282
rect 1094 1276 1095 1280
rect 1099 1276 1100 1280
rect 1094 1275 1100 1276
rect 1278 1279 1284 1280
rect 1278 1275 1279 1279
rect 1283 1275 1284 1279
rect 2142 1279 2143 1280
rect 2147 1279 2148 1283
rect 2142 1278 2148 1279
rect 2406 1279 2412 1280
rect 1278 1274 1284 1275
rect 2406 1275 2407 1279
rect 2411 1275 2412 1279
rect 2406 1274 2412 1275
rect 1446 1272 1452 1273
rect 1446 1268 1447 1272
rect 1451 1268 1452 1272
rect 1446 1267 1452 1268
rect 1486 1272 1492 1273
rect 1486 1268 1487 1272
rect 1491 1268 1492 1272
rect 1486 1267 1492 1268
rect 1526 1272 1532 1273
rect 1526 1268 1527 1272
rect 1531 1268 1532 1272
rect 1526 1267 1532 1268
rect 1566 1272 1572 1273
rect 1566 1268 1567 1272
rect 1571 1268 1572 1272
rect 1566 1267 1572 1268
rect 1614 1272 1620 1273
rect 1614 1268 1615 1272
rect 1619 1268 1620 1272
rect 1614 1267 1620 1268
rect 1670 1272 1676 1273
rect 1670 1268 1671 1272
rect 1675 1268 1676 1272
rect 1670 1267 1676 1268
rect 1718 1272 1724 1273
rect 1718 1268 1719 1272
rect 1723 1268 1724 1272
rect 1718 1267 1724 1268
rect 1774 1272 1780 1273
rect 1774 1268 1775 1272
rect 1779 1268 1780 1272
rect 1774 1267 1780 1268
rect 1830 1272 1836 1273
rect 1830 1268 1831 1272
rect 1835 1268 1836 1272
rect 1830 1267 1836 1268
rect 1902 1272 1908 1273
rect 1902 1268 1903 1272
rect 1907 1268 1908 1272
rect 1902 1267 1908 1268
rect 1982 1272 1988 1273
rect 1982 1268 1983 1272
rect 1987 1268 1988 1272
rect 1982 1267 1988 1268
rect 2070 1272 2076 1273
rect 2070 1268 2071 1272
rect 2075 1268 2076 1272
rect 2070 1267 2076 1268
rect 2166 1272 2172 1273
rect 2166 1268 2167 1272
rect 2171 1268 2172 1272
rect 2166 1267 2172 1268
rect 2270 1272 2276 1273
rect 2270 1268 2271 1272
rect 2275 1268 2276 1272
rect 2270 1267 2276 1268
rect 2358 1272 2364 1273
rect 2358 1268 2359 1272
rect 2363 1268 2364 1272
rect 2358 1267 2364 1268
rect 134 1264 140 1265
rect 134 1260 135 1264
rect 139 1260 140 1264
rect 134 1259 140 1260
rect 174 1264 180 1265
rect 174 1260 175 1264
rect 179 1260 180 1264
rect 174 1259 180 1260
rect 246 1264 252 1265
rect 246 1260 247 1264
rect 251 1260 252 1264
rect 246 1259 252 1260
rect 326 1264 332 1265
rect 326 1260 327 1264
rect 331 1260 332 1264
rect 326 1259 332 1260
rect 414 1264 420 1265
rect 414 1260 415 1264
rect 419 1260 420 1264
rect 414 1259 420 1260
rect 502 1264 508 1265
rect 502 1260 503 1264
rect 507 1260 508 1264
rect 502 1259 508 1260
rect 590 1264 596 1265
rect 590 1260 591 1264
rect 595 1260 596 1264
rect 590 1259 596 1260
rect 670 1264 676 1265
rect 670 1260 671 1264
rect 675 1260 676 1264
rect 670 1259 676 1260
rect 742 1264 748 1265
rect 742 1260 743 1264
rect 747 1260 748 1264
rect 742 1259 748 1260
rect 814 1264 820 1265
rect 814 1260 815 1264
rect 819 1260 820 1264
rect 814 1259 820 1260
rect 878 1264 884 1265
rect 878 1260 879 1264
rect 883 1260 884 1264
rect 878 1259 884 1260
rect 942 1264 948 1265
rect 942 1260 943 1264
rect 947 1260 948 1264
rect 942 1259 948 1260
rect 1006 1264 1012 1265
rect 1006 1260 1007 1264
rect 1011 1260 1012 1264
rect 1006 1259 1012 1260
rect 1070 1264 1076 1265
rect 1070 1260 1071 1264
rect 1075 1260 1076 1264
rect 1070 1259 1076 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 1238 1257 1244 1258
rect 1238 1253 1239 1257
rect 1243 1253 1244 1257
rect 1238 1252 1244 1253
rect 1510 1256 1516 1257
rect 1510 1252 1511 1256
rect 1515 1252 1516 1256
rect 1510 1251 1516 1252
rect 1550 1256 1556 1257
rect 1550 1252 1551 1256
rect 1555 1252 1556 1256
rect 1550 1251 1556 1252
rect 1590 1256 1596 1257
rect 1590 1252 1591 1256
rect 1595 1252 1596 1256
rect 1590 1251 1596 1252
rect 1630 1256 1636 1257
rect 1630 1252 1631 1256
rect 1635 1252 1636 1256
rect 1630 1251 1636 1252
rect 1670 1256 1676 1257
rect 1670 1252 1671 1256
rect 1675 1252 1676 1256
rect 1670 1251 1676 1252
rect 1710 1256 1716 1257
rect 1710 1252 1711 1256
rect 1715 1252 1716 1256
rect 1710 1251 1716 1252
rect 1750 1256 1756 1257
rect 1750 1252 1751 1256
rect 1755 1252 1756 1256
rect 1750 1251 1756 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1838 1256 1844 1257
rect 1838 1252 1839 1256
rect 1843 1252 1844 1256
rect 1838 1251 1844 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 2206 1256 2212 1257
rect 2206 1252 2207 1256
rect 2211 1252 2212 1256
rect 2206 1251 2212 1252
rect 2294 1256 2300 1257
rect 2294 1252 2295 1256
rect 2299 1252 2300 1256
rect 2294 1251 2300 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 1278 1249 1284 1250
rect 1278 1245 1279 1249
rect 1283 1245 1284 1249
rect 1278 1244 1284 1245
rect 2406 1249 2412 1250
rect 2406 1245 2407 1249
rect 2411 1245 2412 1249
rect 2406 1244 2412 1245
rect 159 1243 165 1244
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 159 1239 160 1243
rect 164 1242 165 1243
rect 190 1243 196 1244
rect 190 1242 191 1243
rect 164 1240 191 1242
rect 164 1239 165 1240
rect 159 1238 165 1239
rect 190 1239 191 1240
rect 195 1239 196 1243
rect 190 1238 196 1239
rect 199 1243 205 1244
rect 199 1239 200 1243
rect 204 1239 205 1243
rect 199 1238 205 1239
rect 238 1243 244 1244
rect 238 1239 239 1243
rect 243 1242 244 1243
rect 271 1243 277 1244
rect 271 1242 272 1243
rect 243 1240 272 1242
rect 243 1239 244 1240
rect 238 1238 244 1239
rect 271 1239 272 1240
rect 276 1239 277 1243
rect 271 1238 277 1239
rect 295 1243 301 1244
rect 295 1239 296 1243
rect 300 1242 301 1243
rect 351 1243 357 1244
rect 351 1242 352 1243
rect 300 1240 352 1242
rect 300 1239 301 1240
rect 295 1238 301 1239
rect 351 1239 352 1240
rect 356 1239 357 1243
rect 351 1238 357 1239
rect 359 1243 365 1244
rect 359 1239 360 1243
rect 364 1242 365 1243
rect 439 1243 445 1244
rect 439 1242 440 1243
rect 364 1240 440 1242
rect 364 1239 365 1240
rect 359 1238 365 1239
rect 439 1239 440 1240
rect 444 1239 445 1243
rect 439 1238 445 1239
rect 527 1243 533 1244
rect 527 1239 528 1243
rect 532 1242 533 1243
rect 606 1243 612 1244
rect 606 1242 607 1243
rect 532 1240 607 1242
rect 532 1239 533 1240
rect 527 1238 533 1239
rect 606 1239 607 1240
rect 611 1239 612 1243
rect 606 1238 612 1239
rect 615 1243 621 1244
rect 615 1239 616 1243
rect 620 1242 621 1243
rect 662 1243 668 1244
rect 662 1242 663 1243
rect 620 1240 663 1242
rect 620 1239 621 1240
rect 615 1238 621 1239
rect 662 1239 663 1240
rect 667 1239 668 1243
rect 662 1238 668 1239
rect 678 1243 684 1244
rect 678 1239 679 1243
rect 683 1242 684 1243
rect 695 1243 701 1244
rect 695 1242 696 1243
rect 683 1240 696 1242
rect 683 1239 684 1240
rect 678 1238 684 1239
rect 695 1239 696 1240
rect 700 1239 701 1243
rect 695 1238 701 1239
rect 767 1243 773 1244
rect 767 1239 768 1243
rect 772 1239 773 1243
rect 767 1238 773 1239
rect 775 1243 781 1244
rect 775 1239 776 1243
rect 780 1242 781 1243
rect 839 1243 845 1244
rect 839 1242 840 1243
rect 780 1240 840 1242
rect 780 1239 781 1240
rect 775 1238 781 1239
rect 839 1239 840 1240
rect 844 1239 845 1243
rect 839 1238 845 1239
rect 903 1243 909 1244
rect 903 1239 904 1243
rect 908 1242 909 1243
rect 958 1243 964 1244
rect 958 1242 959 1243
rect 908 1240 959 1242
rect 908 1239 909 1240
rect 903 1238 909 1239
rect 958 1239 959 1240
rect 963 1239 964 1243
rect 958 1238 964 1239
rect 967 1243 973 1244
rect 967 1239 968 1243
rect 972 1242 973 1243
rect 1022 1243 1028 1244
rect 1022 1242 1023 1243
rect 972 1240 1023 1242
rect 972 1239 973 1240
rect 967 1238 973 1239
rect 1022 1239 1023 1240
rect 1027 1239 1028 1243
rect 1022 1238 1028 1239
rect 1031 1243 1037 1244
rect 1031 1239 1032 1243
rect 1036 1242 1037 1243
rect 1086 1243 1092 1244
rect 1086 1242 1087 1243
rect 1036 1240 1087 1242
rect 1036 1239 1037 1240
rect 1031 1238 1037 1239
rect 1086 1239 1087 1240
rect 1091 1239 1092 1243
rect 1086 1238 1092 1239
rect 1095 1243 1101 1244
rect 1095 1239 1096 1243
rect 1100 1242 1101 1243
rect 1106 1243 1112 1244
rect 1106 1242 1107 1243
rect 1100 1240 1107 1242
rect 1100 1239 1101 1240
rect 1095 1238 1101 1239
rect 1106 1239 1107 1240
rect 1111 1239 1112 1243
rect 1106 1238 1112 1239
rect 1238 1240 1244 1241
rect 110 1235 116 1236
rect 201 1234 203 1238
rect 422 1235 428 1236
rect 422 1234 423 1235
rect 201 1232 423 1234
rect 422 1231 423 1232
rect 427 1231 428 1235
rect 769 1234 771 1238
rect 1238 1236 1239 1240
rect 1243 1236 1244 1240
rect 902 1235 908 1236
rect 1238 1235 1244 1236
rect 1535 1235 1541 1236
rect 902 1234 903 1235
rect 769 1232 903 1234
rect 422 1230 428 1231
rect 902 1231 903 1232
rect 907 1231 908 1235
rect 902 1230 908 1231
rect 1278 1232 1284 1233
rect 1278 1228 1279 1232
rect 1283 1228 1284 1232
rect 1535 1231 1536 1235
rect 1540 1234 1541 1235
rect 1558 1235 1564 1236
rect 1540 1232 1554 1234
rect 1540 1231 1541 1232
rect 1535 1230 1541 1231
rect 1278 1227 1284 1228
rect 1552 1226 1554 1232
rect 1558 1231 1559 1235
rect 1563 1234 1564 1235
rect 1575 1235 1581 1236
rect 1575 1234 1576 1235
rect 1563 1232 1576 1234
rect 1563 1231 1564 1232
rect 1558 1230 1564 1231
rect 1575 1231 1576 1232
rect 1580 1231 1581 1235
rect 1575 1230 1581 1231
rect 1598 1235 1604 1236
rect 1598 1231 1599 1235
rect 1603 1234 1604 1235
rect 1615 1235 1621 1236
rect 1615 1234 1616 1235
rect 1603 1232 1616 1234
rect 1603 1231 1604 1232
rect 1598 1230 1604 1231
rect 1615 1231 1616 1232
rect 1620 1231 1621 1235
rect 1615 1230 1621 1231
rect 1655 1235 1661 1236
rect 1655 1231 1656 1235
rect 1660 1234 1661 1235
rect 1686 1235 1692 1236
rect 1686 1234 1687 1235
rect 1660 1232 1687 1234
rect 1660 1231 1661 1232
rect 1655 1230 1661 1231
rect 1686 1231 1687 1232
rect 1691 1231 1692 1235
rect 1686 1230 1692 1231
rect 1695 1235 1701 1236
rect 1695 1231 1696 1235
rect 1700 1234 1701 1235
rect 1726 1235 1732 1236
rect 1726 1234 1727 1235
rect 1700 1232 1727 1234
rect 1700 1231 1701 1232
rect 1695 1230 1701 1231
rect 1726 1231 1727 1232
rect 1731 1231 1732 1235
rect 1726 1230 1732 1231
rect 1735 1235 1741 1236
rect 1735 1231 1736 1235
rect 1740 1234 1741 1235
rect 1758 1235 1764 1236
rect 1758 1234 1759 1235
rect 1740 1232 1759 1234
rect 1740 1231 1741 1232
rect 1735 1230 1741 1231
rect 1758 1231 1759 1232
rect 1763 1231 1764 1235
rect 1758 1230 1764 1231
rect 1766 1235 1772 1236
rect 1766 1231 1767 1235
rect 1771 1234 1772 1235
rect 1775 1235 1781 1236
rect 1775 1234 1776 1235
rect 1771 1232 1776 1234
rect 1771 1231 1772 1232
rect 1766 1230 1772 1231
rect 1775 1231 1776 1232
rect 1780 1231 1781 1235
rect 1775 1230 1781 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1234 1812 1235
rect 1815 1235 1821 1236
rect 1815 1234 1816 1235
rect 1811 1232 1816 1234
rect 1811 1231 1812 1232
rect 1806 1230 1812 1231
rect 1815 1231 1816 1232
rect 1820 1231 1821 1235
rect 1815 1230 1821 1231
rect 1823 1235 1829 1236
rect 1823 1231 1824 1235
rect 1828 1234 1829 1235
rect 1863 1235 1869 1236
rect 1863 1234 1864 1235
rect 1828 1232 1864 1234
rect 1828 1231 1829 1232
rect 1823 1230 1829 1231
rect 1863 1231 1864 1232
rect 1868 1231 1869 1235
rect 1863 1230 1869 1231
rect 1871 1235 1877 1236
rect 1871 1231 1872 1235
rect 1876 1234 1877 1235
rect 1927 1235 1933 1236
rect 1927 1234 1928 1235
rect 1876 1232 1928 1234
rect 1876 1231 1877 1232
rect 1871 1230 1877 1231
rect 1927 1231 1928 1232
rect 1932 1231 1933 1235
rect 1927 1230 1933 1231
rect 1935 1235 1941 1236
rect 1935 1231 1936 1235
rect 1940 1234 1941 1235
rect 1991 1235 1997 1236
rect 1991 1234 1992 1235
rect 1940 1232 1992 1234
rect 1940 1231 1941 1232
rect 1935 1230 1941 1231
rect 1991 1231 1992 1232
rect 1996 1231 1997 1235
rect 1991 1230 1997 1231
rect 2030 1235 2036 1236
rect 2030 1231 2031 1235
rect 2035 1234 2036 1235
rect 2063 1235 2069 1236
rect 2063 1234 2064 1235
rect 2035 1232 2064 1234
rect 2035 1231 2036 1232
rect 2030 1230 2036 1231
rect 2063 1231 2064 1232
rect 2068 1231 2069 1235
rect 2063 1230 2069 1231
rect 2071 1235 2077 1236
rect 2071 1231 2072 1235
rect 2076 1234 2077 1235
rect 2143 1235 2149 1236
rect 2143 1234 2144 1235
rect 2076 1232 2144 1234
rect 2076 1231 2077 1232
rect 2071 1230 2077 1231
rect 2143 1231 2144 1232
rect 2148 1231 2149 1235
rect 2143 1230 2149 1231
rect 2231 1235 2237 1236
rect 2231 1231 2232 1235
rect 2236 1234 2237 1235
rect 2282 1235 2288 1236
rect 2282 1234 2283 1235
rect 2236 1232 2283 1234
rect 2236 1231 2237 1232
rect 2231 1230 2237 1231
rect 2282 1231 2283 1232
rect 2287 1231 2288 1235
rect 2282 1230 2288 1231
rect 2318 1235 2325 1236
rect 2318 1231 2319 1235
rect 2324 1231 2325 1235
rect 2318 1230 2325 1231
rect 2327 1235 2333 1236
rect 2327 1231 2328 1235
rect 2332 1234 2333 1235
rect 2383 1235 2389 1236
rect 2383 1234 2384 1235
rect 2332 1232 2384 1234
rect 2332 1231 2333 1232
rect 2327 1230 2333 1231
rect 2383 1231 2384 1232
rect 2388 1231 2389 1235
rect 2383 1230 2389 1231
rect 2406 1232 2412 1233
rect 2406 1228 2407 1232
rect 2411 1228 2412 1232
rect 1654 1227 1660 1228
rect 2406 1227 2412 1228
rect 1654 1226 1655 1227
rect 1552 1224 1655 1226
rect 1654 1223 1655 1224
rect 1659 1223 1660 1227
rect 1654 1222 1660 1223
rect 134 1217 140 1218
rect 134 1213 135 1217
rect 139 1213 140 1217
rect 134 1212 140 1213
rect 174 1217 180 1218
rect 174 1213 175 1217
rect 179 1213 180 1217
rect 174 1212 180 1213
rect 246 1217 252 1218
rect 246 1213 247 1217
rect 251 1213 252 1217
rect 246 1212 252 1213
rect 326 1217 332 1218
rect 326 1213 327 1217
rect 331 1213 332 1217
rect 326 1212 332 1213
rect 414 1217 420 1218
rect 414 1213 415 1217
rect 419 1213 420 1217
rect 414 1212 420 1213
rect 502 1217 508 1218
rect 502 1213 503 1217
rect 507 1213 508 1217
rect 502 1212 508 1213
rect 590 1217 596 1218
rect 590 1213 591 1217
rect 595 1213 596 1217
rect 590 1212 596 1213
rect 670 1217 676 1218
rect 670 1213 671 1217
rect 675 1213 676 1217
rect 670 1212 676 1213
rect 742 1217 748 1218
rect 742 1213 743 1217
rect 747 1213 748 1217
rect 742 1212 748 1213
rect 814 1217 820 1218
rect 814 1213 815 1217
rect 819 1213 820 1217
rect 814 1212 820 1213
rect 878 1217 884 1218
rect 878 1213 879 1217
rect 883 1213 884 1217
rect 878 1212 884 1213
rect 942 1217 948 1218
rect 942 1213 943 1217
rect 947 1213 948 1217
rect 942 1212 948 1213
rect 1006 1217 1012 1218
rect 1006 1213 1007 1217
rect 1011 1213 1012 1217
rect 1006 1212 1012 1213
rect 1070 1217 1076 1218
rect 1070 1213 1071 1217
rect 1075 1213 1076 1217
rect 1070 1212 1076 1213
rect 158 1211 165 1212
rect 158 1207 159 1211
rect 164 1207 165 1211
rect 158 1206 165 1207
rect 190 1211 196 1212
rect 190 1207 191 1211
rect 195 1210 196 1211
rect 199 1211 205 1212
rect 199 1210 200 1211
rect 195 1208 200 1210
rect 195 1207 196 1208
rect 190 1206 196 1207
rect 199 1207 200 1208
rect 204 1207 205 1211
rect 199 1206 205 1207
rect 271 1211 277 1212
rect 271 1207 272 1211
rect 276 1210 277 1211
rect 295 1211 301 1212
rect 295 1210 296 1211
rect 276 1208 296 1210
rect 276 1207 277 1208
rect 271 1206 277 1207
rect 295 1207 296 1208
rect 300 1207 301 1211
rect 295 1206 301 1207
rect 351 1211 357 1212
rect 351 1207 352 1211
rect 356 1210 357 1211
rect 359 1211 365 1212
rect 359 1210 360 1211
rect 356 1208 360 1210
rect 356 1207 357 1208
rect 351 1206 357 1207
rect 359 1207 360 1208
rect 364 1207 365 1211
rect 359 1206 365 1207
rect 422 1211 428 1212
rect 422 1207 423 1211
rect 427 1210 428 1211
rect 439 1211 445 1212
rect 439 1210 440 1211
rect 427 1208 440 1210
rect 427 1207 428 1208
rect 422 1206 428 1207
rect 439 1207 440 1208
rect 444 1207 445 1211
rect 439 1206 445 1207
rect 527 1211 533 1212
rect 527 1207 528 1211
rect 532 1210 533 1211
rect 542 1211 548 1212
rect 542 1210 543 1211
rect 532 1208 543 1210
rect 532 1207 533 1208
rect 527 1206 533 1207
rect 542 1207 543 1208
rect 547 1207 548 1211
rect 542 1206 548 1207
rect 606 1211 612 1212
rect 606 1207 607 1211
rect 611 1210 612 1211
rect 615 1211 621 1212
rect 615 1210 616 1211
rect 611 1208 616 1210
rect 611 1207 612 1208
rect 606 1206 612 1207
rect 615 1207 616 1208
rect 620 1207 621 1211
rect 615 1206 621 1207
rect 662 1211 668 1212
rect 662 1207 663 1211
rect 667 1210 668 1211
rect 695 1211 701 1212
rect 695 1210 696 1211
rect 667 1208 696 1210
rect 667 1207 668 1208
rect 662 1206 668 1207
rect 695 1207 696 1208
rect 700 1207 701 1211
rect 695 1206 701 1207
rect 767 1211 773 1212
rect 767 1207 768 1211
rect 772 1210 773 1211
rect 775 1211 781 1212
rect 775 1210 776 1211
rect 772 1208 776 1210
rect 772 1207 773 1208
rect 767 1206 773 1207
rect 775 1207 776 1208
rect 780 1207 781 1211
rect 775 1206 781 1207
rect 839 1211 845 1212
rect 839 1207 840 1211
rect 844 1210 845 1211
rect 894 1211 900 1212
rect 894 1210 895 1211
rect 844 1208 895 1210
rect 844 1207 845 1208
rect 839 1206 845 1207
rect 894 1207 895 1208
rect 899 1207 900 1211
rect 894 1206 900 1207
rect 902 1211 909 1212
rect 902 1207 903 1211
rect 908 1207 909 1211
rect 902 1206 909 1207
rect 958 1211 964 1212
rect 958 1207 959 1211
rect 963 1210 964 1211
rect 967 1211 973 1212
rect 967 1210 968 1211
rect 963 1208 968 1210
rect 963 1207 964 1208
rect 958 1206 964 1207
rect 967 1207 968 1208
rect 972 1207 973 1211
rect 967 1206 973 1207
rect 1022 1211 1028 1212
rect 1022 1207 1023 1211
rect 1027 1210 1028 1211
rect 1031 1211 1037 1212
rect 1031 1210 1032 1211
rect 1027 1208 1032 1210
rect 1027 1207 1028 1208
rect 1022 1206 1028 1207
rect 1031 1207 1032 1208
rect 1036 1207 1037 1211
rect 1031 1206 1037 1207
rect 1086 1211 1092 1212
rect 1086 1207 1087 1211
rect 1091 1210 1092 1211
rect 1095 1211 1101 1212
rect 1095 1210 1096 1211
rect 1091 1208 1096 1210
rect 1091 1207 1092 1208
rect 1086 1206 1092 1207
rect 1095 1207 1096 1208
rect 1100 1207 1101 1211
rect 1095 1206 1101 1207
rect 1510 1209 1516 1210
rect 1510 1205 1511 1209
rect 1515 1205 1516 1209
rect 1510 1204 1516 1205
rect 1550 1209 1556 1210
rect 1550 1205 1551 1209
rect 1555 1205 1556 1209
rect 1550 1204 1556 1205
rect 1590 1209 1596 1210
rect 1590 1205 1591 1209
rect 1595 1205 1596 1209
rect 1590 1204 1596 1205
rect 1630 1209 1636 1210
rect 1630 1205 1631 1209
rect 1635 1205 1636 1209
rect 1630 1204 1636 1205
rect 1670 1209 1676 1210
rect 1670 1205 1671 1209
rect 1675 1205 1676 1209
rect 1670 1204 1676 1205
rect 1710 1209 1716 1210
rect 1710 1205 1711 1209
rect 1715 1205 1716 1209
rect 1710 1204 1716 1205
rect 1750 1209 1756 1210
rect 1750 1205 1751 1209
rect 1755 1205 1756 1209
rect 1750 1204 1756 1205
rect 1790 1209 1796 1210
rect 1790 1205 1791 1209
rect 1795 1205 1796 1209
rect 1790 1204 1796 1205
rect 1838 1209 1844 1210
rect 1838 1205 1839 1209
rect 1843 1205 1844 1209
rect 1838 1204 1844 1205
rect 1902 1209 1908 1210
rect 1902 1205 1903 1209
rect 1907 1205 1908 1209
rect 1902 1204 1908 1205
rect 1966 1209 1972 1210
rect 1966 1205 1967 1209
rect 1971 1205 1972 1209
rect 1966 1204 1972 1205
rect 2038 1209 2044 1210
rect 2038 1205 2039 1209
rect 2043 1205 2044 1209
rect 2038 1204 2044 1205
rect 2118 1209 2124 1210
rect 2118 1205 2119 1209
rect 2123 1205 2124 1209
rect 2118 1204 2124 1205
rect 2206 1209 2212 1210
rect 2206 1205 2207 1209
rect 2211 1205 2212 1209
rect 2206 1204 2212 1205
rect 2294 1209 2300 1210
rect 2294 1205 2295 1209
rect 2299 1205 2300 1209
rect 2294 1204 2300 1205
rect 2358 1209 2364 1210
rect 2358 1205 2359 1209
rect 2363 1205 2364 1209
rect 2358 1204 2364 1205
rect 1535 1203 1541 1204
rect 1535 1199 1536 1203
rect 1540 1202 1541 1203
rect 1558 1203 1564 1204
rect 1558 1202 1559 1203
rect 1540 1200 1559 1202
rect 1540 1199 1541 1200
rect 1535 1198 1541 1199
rect 1558 1199 1559 1200
rect 1563 1199 1564 1203
rect 1558 1198 1564 1199
rect 1575 1203 1581 1204
rect 1575 1199 1576 1203
rect 1580 1202 1581 1203
rect 1598 1203 1604 1204
rect 1598 1202 1599 1203
rect 1580 1200 1599 1202
rect 1580 1199 1581 1200
rect 1575 1198 1581 1199
rect 1598 1199 1599 1200
rect 1603 1199 1604 1203
rect 1598 1198 1604 1199
rect 1615 1203 1621 1204
rect 1615 1199 1616 1203
rect 1620 1199 1621 1203
rect 1615 1198 1621 1199
rect 1654 1203 1661 1204
rect 1654 1199 1655 1203
rect 1660 1199 1661 1203
rect 1654 1198 1661 1199
rect 1686 1203 1692 1204
rect 1686 1199 1687 1203
rect 1691 1202 1692 1203
rect 1695 1203 1701 1204
rect 1695 1202 1696 1203
rect 1691 1200 1696 1202
rect 1691 1199 1692 1200
rect 1686 1198 1692 1199
rect 1695 1199 1696 1200
rect 1700 1199 1701 1203
rect 1695 1198 1701 1199
rect 1726 1203 1732 1204
rect 1726 1199 1727 1203
rect 1731 1202 1732 1203
rect 1735 1203 1741 1204
rect 1735 1202 1736 1203
rect 1731 1200 1736 1202
rect 1731 1199 1732 1200
rect 1726 1198 1732 1199
rect 1735 1199 1736 1200
rect 1740 1199 1741 1203
rect 1735 1198 1741 1199
rect 1758 1203 1764 1204
rect 1758 1199 1759 1203
rect 1763 1202 1764 1203
rect 1775 1203 1781 1204
rect 1775 1202 1776 1203
rect 1763 1200 1776 1202
rect 1763 1199 1764 1200
rect 1758 1198 1764 1199
rect 1775 1199 1776 1200
rect 1780 1199 1781 1203
rect 1775 1198 1781 1199
rect 1815 1203 1821 1204
rect 1815 1199 1816 1203
rect 1820 1202 1821 1203
rect 1823 1203 1829 1204
rect 1823 1202 1824 1203
rect 1820 1200 1824 1202
rect 1820 1199 1821 1200
rect 1815 1198 1821 1199
rect 1823 1199 1824 1200
rect 1828 1199 1829 1203
rect 1823 1198 1829 1199
rect 1863 1203 1869 1204
rect 1863 1199 1864 1203
rect 1868 1202 1869 1203
rect 1871 1203 1877 1204
rect 1871 1202 1872 1203
rect 1868 1200 1872 1202
rect 1868 1199 1869 1200
rect 1863 1198 1869 1199
rect 1871 1199 1872 1200
rect 1876 1199 1877 1203
rect 1871 1198 1877 1199
rect 1927 1203 1933 1204
rect 1927 1199 1928 1203
rect 1932 1202 1933 1203
rect 1935 1203 1941 1204
rect 1935 1202 1936 1203
rect 1932 1200 1936 1202
rect 1932 1199 1933 1200
rect 1927 1198 1933 1199
rect 1935 1199 1936 1200
rect 1940 1199 1941 1203
rect 1935 1198 1941 1199
rect 1991 1203 1997 1204
rect 1991 1199 1992 1203
rect 1996 1202 1997 1203
rect 2030 1203 2036 1204
rect 2030 1202 2031 1203
rect 1996 1200 2031 1202
rect 1996 1199 1997 1200
rect 1991 1198 1997 1199
rect 2030 1199 2031 1200
rect 2035 1199 2036 1203
rect 2030 1198 2036 1199
rect 2063 1203 2069 1204
rect 2063 1199 2064 1203
rect 2068 1202 2069 1203
rect 2071 1203 2077 1204
rect 2071 1202 2072 1203
rect 2068 1200 2072 1202
rect 2068 1199 2069 1200
rect 2063 1198 2069 1199
rect 2071 1199 2072 1200
rect 2076 1199 2077 1203
rect 2071 1198 2077 1199
rect 2142 1203 2149 1204
rect 2142 1199 2143 1203
rect 2148 1199 2149 1203
rect 2142 1198 2149 1199
rect 2218 1203 2224 1204
rect 2218 1199 2219 1203
rect 2223 1202 2224 1203
rect 2231 1203 2237 1204
rect 2231 1202 2232 1203
rect 2223 1200 2232 1202
rect 2223 1199 2224 1200
rect 2218 1198 2224 1199
rect 2231 1199 2232 1200
rect 2236 1199 2237 1203
rect 2231 1198 2237 1199
rect 2319 1203 2325 1204
rect 2319 1199 2320 1203
rect 2324 1202 2325 1203
rect 2327 1203 2333 1204
rect 2327 1202 2328 1203
rect 2324 1200 2328 1202
rect 2324 1199 2325 1200
rect 2319 1198 2325 1199
rect 2327 1199 2328 1200
rect 2332 1199 2333 1203
rect 2327 1198 2333 1199
rect 2382 1203 2389 1204
rect 2382 1199 2383 1203
rect 2388 1199 2389 1203
rect 2382 1198 2389 1199
rect 190 1187 196 1188
rect 190 1186 191 1187
rect 161 1184 191 1186
rect 159 1183 165 1184
rect 134 1179 140 1180
rect 134 1175 135 1179
rect 139 1175 140 1179
rect 159 1179 160 1183
rect 164 1179 165 1183
rect 190 1183 191 1184
rect 195 1183 196 1187
rect 1206 1187 1212 1188
rect 1206 1186 1207 1187
rect 1177 1184 1207 1186
rect 190 1182 196 1183
rect 199 1183 205 1184
rect 159 1178 165 1179
rect 174 1179 180 1180
rect 134 1174 140 1175
rect 174 1175 175 1179
rect 179 1175 180 1179
rect 199 1179 200 1183
rect 204 1182 205 1183
rect 222 1183 228 1184
rect 222 1182 223 1183
rect 204 1180 223 1182
rect 204 1179 205 1180
rect 199 1178 205 1179
rect 222 1179 223 1180
rect 227 1179 228 1183
rect 255 1183 261 1184
rect 222 1178 228 1179
rect 230 1179 236 1180
rect 174 1174 180 1175
rect 230 1175 231 1179
rect 235 1175 236 1179
rect 255 1179 256 1183
rect 260 1182 261 1183
rect 294 1183 300 1184
rect 294 1182 295 1183
rect 260 1180 295 1182
rect 260 1179 261 1180
rect 255 1178 261 1179
rect 294 1179 295 1180
rect 299 1179 300 1183
rect 327 1183 333 1184
rect 294 1178 300 1179
rect 302 1179 308 1180
rect 230 1174 236 1175
rect 302 1175 303 1179
rect 307 1175 308 1179
rect 327 1179 328 1183
rect 332 1182 333 1183
rect 374 1183 380 1184
rect 374 1182 375 1183
rect 332 1180 375 1182
rect 332 1179 333 1180
rect 327 1178 333 1179
rect 374 1179 375 1180
rect 379 1179 380 1183
rect 398 1183 404 1184
rect 374 1178 380 1179
rect 382 1179 388 1180
rect 302 1174 308 1175
rect 382 1175 383 1179
rect 387 1175 388 1179
rect 398 1179 399 1183
rect 403 1182 404 1183
rect 407 1183 413 1184
rect 407 1182 408 1183
rect 403 1180 408 1182
rect 403 1179 404 1180
rect 398 1178 404 1179
rect 407 1179 408 1180
rect 412 1179 413 1183
rect 495 1183 501 1184
rect 407 1178 413 1179
rect 470 1179 476 1180
rect 382 1174 388 1175
rect 470 1175 471 1179
rect 475 1175 476 1179
rect 495 1179 496 1183
rect 500 1182 501 1183
rect 550 1183 556 1184
rect 550 1182 551 1183
rect 500 1180 551 1182
rect 500 1179 501 1180
rect 495 1178 501 1179
rect 550 1179 551 1180
rect 555 1179 556 1183
rect 583 1183 589 1184
rect 550 1178 556 1179
rect 558 1179 564 1180
rect 470 1174 476 1175
rect 558 1175 559 1179
rect 563 1175 564 1179
rect 583 1179 584 1183
rect 588 1182 589 1183
rect 630 1183 636 1184
rect 630 1182 631 1183
rect 588 1180 631 1182
rect 588 1179 589 1180
rect 583 1178 589 1179
rect 630 1179 631 1180
rect 635 1179 636 1183
rect 663 1183 669 1184
rect 630 1178 636 1179
rect 638 1179 644 1180
rect 558 1174 564 1175
rect 638 1175 639 1179
rect 643 1175 644 1179
rect 663 1179 664 1183
rect 668 1182 669 1183
rect 678 1183 684 1184
rect 678 1182 679 1183
rect 668 1180 679 1182
rect 668 1179 669 1180
rect 663 1178 669 1179
rect 678 1179 679 1180
rect 683 1179 684 1183
rect 738 1183 749 1184
rect 678 1178 684 1179
rect 718 1179 724 1180
rect 638 1174 644 1175
rect 718 1175 719 1179
rect 723 1175 724 1179
rect 738 1179 739 1183
rect 743 1179 744 1183
rect 748 1179 749 1183
rect 810 1183 816 1184
rect 738 1178 749 1179
rect 798 1179 804 1180
rect 718 1174 724 1175
rect 798 1175 799 1179
rect 803 1175 804 1179
rect 810 1179 811 1183
rect 815 1182 816 1183
rect 823 1183 829 1184
rect 823 1182 824 1183
rect 815 1180 824 1182
rect 815 1179 816 1180
rect 810 1178 816 1179
rect 823 1179 824 1180
rect 828 1179 829 1183
rect 882 1183 888 1184
rect 823 1178 829 1179
rect 870 1179 876 1180
rect 798 1174 804 1175
rect 870 1175 871 1179
rect 875 1175 876 1179
rect 882 1179 883 1183
rect 887 1182 888 1183
rect 895 1183 901 1184
rect 895 1182 896 1183
rect 887 1180 896 1182
rect 887 1179 888 1180
rect 882 1178 888 1179
rect 895 1179 896 1180
rect 900 1179 901 1183
rect 959 1183 965 1184
rect 895 1178 901 1179
rect 934 1179 940 1180
rect 870 1174 876 1175
rect 934 1175 935 1179
rect 939 1175 940 1179
rect 959 1179 960 1183
rect 964 1182 965 1183
rect 982 1183 988 1184
rect 982 1182 983 1183
rect 964 1180 983 1182
rect 964 1179 965 1180
rect 959 1178 965 1179
rect 982 1179 983 1180
rect 987 1179 988 1183
rect 1015 1183 1021 1184
rect 982 1178 988 1179
rect 990 1179 996 1180
rect 934 1174 940 1175
rect 990 1175 991 1179
rect 995 1175 996 1179
rect 1015 1179 1016 1183
rect 1020 1182 1021 1183
rect 1038 1183 1044 1184
rect 1038 1182 1039 1183
rect 1020 1180 1039 1182
rect 1020 1179 1021 1180
rect 1015 1178 1021 1179
rect 1038 1179 1039 1180
rect 1043 1179 1044 1183
rect 1071 1183 1077 1184
rect 1038 1178 1044 1179
rect 1046 1179 1052 1180
rect 990 1174 996 1175
rect 1046 1175 1047 1179
rect 1051 1175 1052 1179
rect 1071 1179 1072 1183
rect 1076 1182 1077 1183
rect 1094 1183 1100 1184
rect 1094 1182 1095 1183
rect 1076 1180 1095 1182
rect 1076 1179 1077 1180
rect 1071 1178 1077 1179
rect 1094 1179 1095 1180
rect 1099 1179 1100 1183
rect 1127 1183 1133 1184
rect 1094 1178 1100 1179
rect 1102 1179 1108 1180
rect 1046 1174 1052 1175
rect 1102 1175 1103 1179
rect 1107 1175 1108 1179
rect 1127 1179 1128 1183
rect 1132 1182 1133 1183
rect 1142 1183 1148 1184
rect 1142 1182 1143 1183
rect 1132 1180 1143 1182
rect 1132 1179 1133 1180
rect 1127 1178 1133 1179
rect 1142 1179 1143 1180
rect 1147 1179 1148 1183
rect 1175 1183 1181 1184
rect 1142 1178 1148 1179
rect 1150 1179 1156 1180
rect 1102 1174 1108 1175
rect 1150 1175 1151 1179
rect 1155 1175 1156 1179
rect 1175 1179 1176 1183
rect 1180 1179 1181 1183
rect 1206 1183 1207 1184
rect 1211 1183 1212 1187
rect 1206 1182 1212 1183
rect 1214 1183 1221 1184
rect 1175 1178 1181 1179
rect 1190 1179 1196 1180
rect 1150 1174 1156 1175
rect 1190 1175 1191 1179
rect 1195 1175 1196 1179
rect 1214 1179 1215 1183
rect 1220 1179 1221 1183
rect 1614 1183 1620 1184
rect 1614 1182 1615 1183
rect 1585 1180 1615 1182
rect 1214 1178 1221 1179
rect 1583 1179 1589 1180
rect 1190 1174 1196 1175
rect 1558 1175 1564 1176
rect 1558 1171 1559 1175
rect 1563 1171 1564 1175
rect 1583 1175 1584 1179
rect 1588 1175 1589 1179
rect 1614 1179 1615 1180
rect 1619 1179 1620 1183
rect 1694 1183 1700 1184
rect 1694 1182 1695 1183
rect 1665 1180 1695 1182
rect 1614 1178 1620 1179
rect 1623 1179 1632 1180
rect 1583 1174 1589 1175
rect 1598 1175 1604 1176
rect 1558 1170 1564 1171
rect 1598 1171 1599 1175
rect 1603 1171 1604 1175
rect 1623 1175 1624 1179
rect 1631 1175 1632 1179
rect 1663 1179 1669 1180
rect 1623 1174 1632 1175
rect 1638 1175 1644 1176
rect 1598 1170 1604 1171
rect 1638 1171 1639 1175
rect 1643 1171 1644 1175
rect 1663 1175 1664 1179
rect 1668 1175 1669 1179
rect 1694 1179 1695 1180
rect 1699 1179 1700 1183
rect 1734 1183 1740 1184
rect 1734 1182 1735 1183
rect 1705 1180 1735 1182
rect 1694 1178 1700 1179
rect 1703 1179 1709 1180
rect 1663 1174 1669 1175
rect 1678 1175 1684 1176
rect 1638 1170 1644 1171
rect 1678 1171 1679 1175
rect 1683 1171 1684 1175
rect 1703 1175 1704 1179
rect 1708 1175 1709 1179
rect 1734 1179 1735 1180
rect 1739 1179 1740 1183
rect 1766 1183 1772 1184
rect 1766 1182 1767 1183
rect 1745 1180 1767 1182
rect 1734 1178 1740 1179
rect 1743 1179 1749 1180
rect 1703 1174 1709 1175
rect 1718 1175 1724 1176
rect 1678 1170 1684 1171
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1743 1175 1744 1179
rect 1748 1175 1749 1179
rect 1766 1179 1767 1180
rect 1771 1179 1772 1183
rect 1806 1183 1812 1184
rect 1806 1182 1807 1183
rect 1785 1180 1807 1182
rect 1766 1178 1772 1179
rect 1783 1179 1789 1180
rect 1743 1174 1749 1175
rect 1758 1175 1764 1176
rect 1718 1170 1724 1171
rect 1758 1171 1759 1175
rect 1763 1171 1764 1175
rect 1783 1175 1784 1179
rect 1788 1175 1789 1179
rect 1806 1179 1807 1180
rect 1811 1179 1812 1183
rect 2318 1183 2324 1184
rect 1806 1178 1812 1179
rect 1814 1179 1820 1180
rect 1783 1174 1789 1175
rect 1798 1175 1804 1176
rect 1758 1170 1764 1171
rect 1798 1171 1799 1175
rect 1803 1171 1804 1175
rect 1814 1175 1815 1179
rect 1819 1178 1820 1179
rect 1823 1179 1829 1180
rect 1823 1178 1824 1179
rect 1819 1176 1824 1178
rect 1819 1175 1820 1176
rect 1814 1174 1820 1175
rect 1823 1175 1824 1176
rect 1828 1175 1829 1179
rect 1866 1179 1872 1180
rect 1823 1174 1829 1175
rect 1854 1175 1860 1176
rect 1798 1170 1804 1171
rect 1854 1171 1855 1175
rect 1859 1171 1860 1175
rect 1866 1175 1867 1179
rect 1871 1178 1872 1179
rect 1879 1179 1885 1180
rect 1879 1178 1880 1179
rect 1871 1176 1880 1178
rect 1871 1175 1872 1176
rect 1866 1174 1872 1175
rect 1879 1175 1880 1176
rect 1884 1175 1885 1179
rect 1938 1179 1944 1180
rect 1879 1174 1885 1175
rect 1926 1175 1932 1176
rect 1854 1170 1860 1171
rect 1926 1171 1927 1175
rect 1931 1171 1932 1175
rect 1938 1175 1939 1179
rect 1943 1178 1944 1179
rect 1951 1179 1957 1180
rect 1951 1178 1952 1179
rect 1943 1176 1952 1178
rect 1943 1175 1944 1176
rect 1938 1174 1944 1175
rect 1951 1175 1952 1176
rect 1956 1175 1957 1179
rect 2047 1179 2053 1180
rect 1951 1174 1957 1175
rect 2022 1175 2028 1176
rect 1926 1170 1932 1171
rect 2022 1171 2023 1175
rect 2027 1171 2028 1175
rect 2047 1175 2048 1179
rect 2052 1178 2053 1179
rect 2126 1179 2132 1180
rect 2126 1178 2127 1179
rect 2052 1176 2127 1178
rect 2052 1175 2053 1176
rect 2047 1174 2053 1175
rect 2126 1175 2127 1176
rect 2131 1175 2132 1179
rect 2159 1179 2165 1180
rect 2126 1174 2132 1175
rect 2134 1175 2140 1176
rect 2022 1170 2028 1171
rect 2134 1171 2135 1175
rect 2139 1171 2140 1175
rect 2159 1175 2160 1179
rect 2164 1178 2165 1179
rect 2246 1179 2252 1180
rect 2246 1178 2247 1179
rect 2164 1176 2247 1178
rect 2164 1175 2165 1176
rect 2159 1174 2165 1175
rect 2246 1175 2247 1176
rect 2251 1175 2252 1179
rect 2266 1179 2272 1180
rect 2246 1174 2252 1175
rect 2254 1175 2260 1176
rect 2134 1170 2140 1171
rect 2254 1171 2255 1175
rect 2259 1171 2260 1175
rect 2266 1175 2267 1179
rect 2271 1178 2272 1179
rect 2279 1179 2285 1180
rect 2279 1178 2280 1179
rect 2271 1176 2280 1178
rect 2271 1175 2272 1176
rect 2266 1174 2272 1175
rect 2279 1175 2280 1176
rect 2284 1175 2285 1179
rect 2318 1179 2319 1183
rect 2323 1182 2324 1183
rect 2323 1180 2387 1182
rect 2323 1179 2324 1180
rect 2318 1178 2324 1179
rect 2383 1179 2389 1180
rect 2279 1174 2285 1175
rect 2358 1175 2364 1176
rect 2254 1170 2260 1171
rect 2358 1171 2359 1175
rect 2363 1171 2364 1175
rect 2383 1175 2384 1179
rect 2388 1175 2389 1179
rect 2383 1174 2389 1175
rect 2358 1170 2364 1171
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 1238 1156 1244 1157
rect 1238 1152 1239 1156
rect 1243 1152 1244 1156
rect 1626 1155 1632 1156
rect 110 1151 116 1152
rect 158 1151 165 1152
rect 158 1147 159 1151
rect 164 1147 165 1151
rect 158 1146 165 1147
rect 190 1151 196 1152
rect 190 1147 191 1151
rect 195 1150 196 1151
rect 199 1151 205 1152
rect 199 1150 200 1151
rect 195 1148 200 1150
rect 195 1147 196 1148
rect 190 1146 196 1147
rect 199 1147 200 1148
rect 204 1147 205 1151
rect 199 1146 205 1147
rect 222 1151 228 1152
rect 222 1147 223 1151
rect 227 1150 228 1151
rect 255 1151 261 1152
rect 255 1150 256 1151
rect 227 1148 256 1150
rect 227 1147 228 1148
rect 222 1146 228 1147
rect 255 1147 256 1148
rect 260 1147 261 1151
rect 255 1146 261 1147
rect 294 1151 300 1152
rect 294 1147 295 1151
rect 299 1150 300 1151
rect 327 1151 333 1152
rect 327 1150 328 1151
rect 299 1148 328 1150
rect 299 1147 300 1148
rect 294 1146 300 1147
rect 327 1147 328 1148
rect 332 1147 333 1151
rect 327 1146 333 1147
rect 374 1151 380 1152
rect 374 1147 375 1151
rect 379 1150 380 1151
rect 407 1151 413 1152
rect 407 1150 408 1151
rect 379 1148 408 1150
rect 379 1147 380 1148
rect 374 1146 380 1147
rect 407 1147 408 1148
rect 412 1147 413 1151
rect 407 1146 413 1147
rect 495 1151 504 1152
rect 495 1147 496 1151
rect 503 1147 504 1151
rect 495 1146 504 1147
rect 550 1151 556 1152
rect 550 1147 551 1151
rect 555 1150 556 1151
rect 583 1151 589 1152
rect 583 1150 584 1151
rect 555 1148 584 1150
rect 555 1147 556 1148
rect 550 1146 556 1147
rect 583 1147 584 1148
rect 588 1147 589 1151
rect 583 1146 589 1147
rect 630 1151 636 1152
rect 630 1147 631 1151
rect 635 1150 636 1151
rect 663 1151 669 1152
rect 663 1150 664 1151
rect 635 1148 664 1150
rect 635 1147 636 1148
rect 630 1146 636 1147
rect 663 1147 664 1148
rect 668 1147 669 1151
rect 663 1146 669 1147
rect 743 1151 749 1152
rect 743 1147 744 1151
rect 748 1150 749 1151
rect 810 1151 816 1152
rect 810 1150 811 1151
rect 748 1148 811 1150
rect 748 1147 749 1148
rect 743 1146 749 1147
rect 810 1147 811 1148
rect 815 1147 816 1151
rect 810 1146 816 1147
rect 823 1151 829 1152
rect 823 1147 824 1151
rect 828 1150 829 1151
rect 882 1151 888 1152
rect 882 1150 883 1151
rect 828 1148 883 1150
rect 828 1147 829 1148
rect 823 1146 829 1147
rect 882 1147 883 1148
rect 887 1147 888 1151
rect 882 1146 888 1147
rect 894 1151 901 1152
rect 894 1147 895 1151
rect 900 1147 901 1151
rect 894 1146 901 1147
rect 959 1151 965 1152
rect 959 1147 960 1151
rect 964 1150 965 1151
rect 982 1151 988 1152
rect 964 1148 978 1150
rect 964 1147 965 1148
rect 959 1146 965 1147
rect 976 1142 978 1148
rect 982 1147 983 1151
rect 987 1150 988 1151
rect 1015 1151 1021 1152
rect 1015 1150 1016 1151
rect 987 1148 1016 1150
rect 987 1147 988 1148
rect 982 1146 988 1147
rect 1015 1147 1016 1148
rect 1020 1147 1021 1151
rect 1015 1146 1021 1147
rect 1038 1151 1044 1152
rect 1038 1147 1039 1151
rect 1043 1150 1044 1151
rect 1071 1151 1077 1152
rect 1071 1150 1072 1151
rect 1043 1148 1072 1150
rect 1043 1147 1044 1148
rect 1038 1146 1044 1147
rect 1071 1147 1072 1148
rect 1076 1147 1077 1151
rect 1071 1146 1077 1147
rect 1094 1151 1100 1152
rect 1094 1147 1095 1151
rect 1099 1150 1100 1151
rect 1127 1151 1133 1152
rect 1127 1150 1128 1151
rect 1099 1148 1128 1150
rect 1099 1147 1100 1148
rect 1094 1146 1100 1147
rect 1127 1147 1128 1148
rect 1132 1147 1133 1151
rect 1127 1146 1133 1147
rect 1142 1151 1148 1152
rect 1142 1147 1143 1151
rect 1147 1150 1148 1151
rect 1175 1151 1181 1152
rect 1175 1150 1176 1151
rect 1147 1148 1176 1150
rect 1147 1147 1148 1148
rect 1142 1146 1148 1147
rect 1175 1147 1176 1148
rect 1180 1147 1181 1151
rect 1175 1146 1181 1147
rect 1206 1151 1212 1152
rect 1206 1147 1207 1151
rect 1211 1150 1212 1151
rect 1215 1151 1221 1152
rect 1238 1151 1244 1152
rect 1278 1152 1284 1153
rect 1215 1150 1216 1151
rect 1211 1148 1216 1150
rect 1211 1147 1212 1148
rect 1206 1146 1212 1147
rect 1215 1147 1216 1148
rect 1220 1147 1221 1151
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1626 1151 1627 1155
rect 1631 1154 1632 1155
rect 2266 1155 2272 1156
rect 2266 1154 2267 1155
rect 1631 1152 1667 1154
rect 1631 1151 1632 1152
rect 1626 1150 1632 1151
rect 1665 1148 1667 1152
rect 1968 1152 2267 1154
rect 1278 1147 1284 1148
rect 1583 1147 1589 1148
rect 1215 1146 1221 1147
rect 1014 1143 1020 1144
rect 1014 1142 1015 1143
rect 976 1140 1015 1142
rect 110 1139 116 1140
rect 110 1135 111 1139
rect 115 1135 116 1139
rect 1014 1139 1015 1140
rect 1019 1139 1020 1143
rect 1583 1143 1584 1147
rect 1588 1143 1589 1147
rect 1583 1142 1589 1143
rect 1614 1147 1620 1148
rect 1614 1143 1615 1147
rect 1619 1146 1620 1147
rect 1623 1147 1629 1148
rect 1623 1146 1624 1147
rect 1619 1144 1624 1146
rect 1619 1143 1620 1144
rect 1614 1142 1620 1143
rect 1623 1143 1624 1144
rect 1628 1143 1629 1147
rect 1623 1142 1629 1143
rect 1663 1147 1669 1148
rect 1663 1143 1664 1147
rect 1668 1143 1669 1147
rect 1663 1142 1669 1143
rect 1694 1147 1700 1148
rect 1694 1143 1695 1147
rect 1699 1146 1700 1147
rect 1703 1147 1709 1148
rect 1703 1146 1704 1147
rect 1699 1144 1704 1146
rect 1699 1143 1700 1144
rect 1694 1142 1700 1143
rect 1703 1143 1704 1144
rect 1708 1143 1709 1147
rect 1703 1142 1709 1143
rect 1734 1147 1740 1148
rect 1734 1143 1735 1147
rect 1739 1146 1740 1147
rect 1743 1147 1749 1148
rect 1743 1146 1744 1147
rect 1739 1144 1744 1146
rect 1739 1143 1740 1144
rect 1734 1142 1740 1143
rect 1743 1143 1744 1144
rect 1748 1143 1749 1147
rect 1743 1142 1749 1143
rect 1783 1147 1789 1148
rect 1783 1143 1784 1147
rect 1788 1146 1789 1147
rect 1814 1147 1820 1148
rect 1814 1146 1815 1147
rect 1788 1144 1815 1146
rect 1788 1143 1789 1144
rect 1783 1142 1789 1143
rect 1814 1143 1815 1144
rect 1819 1143 1820 1147
rect 1814 1142 1820 1143
rect 1823 1147 1829 1148
rect 1823 1143 1824 1147
rect 1828 1146 1829 1147
rect 1866 1147 1872 1148
rect 1866 1146 1867 1147
rect 1828 1144 1867 1146
rect 1828 1143 1829 1144
rect 1823 1142 1829 1143
rect 1866 1143 1867 1144
rect 1871 1143 1872 1147
rect 1866 1142 1872 1143
rect 1879 1147 1885 1148
rect 1879 1143 1880 1147
rect 1884 1146 1885 1147
rect 1938 1147 1944 1148
rect 1938 1146 1939 1147
rect 1884 1144 1939 1146
rect 1884 1143 1885 1144
rect 1879 1142 1885 1143
rect 1938 1143 1939 1144
rect 1943 1143 1944 1147
rect 1938 1142 1944 1143
rect 1951 1147 1957 1148
rect 1951 1143 1952 1147
rect 1956 1146 1957 1147
rect 1968 1146 1970 1152
rect 2266 1151 2267 1152
rect 2271 1151 2272 1155
rect 2266 1150 2272 1151
rect 2406 1152 2412 1153
rect 2406 1148 2407 1152
rect 2411 1148 2412 1152
rect 1956 1144 1970 1146
rect 1974 1147 1980 1148
rect 1956 1143 1957 1144
rect 1951 1142 1957 1143
rect 1974 1143 1975 1147
rect 1979 1146 1980 1147
rect 2047 1147 2053 1148
rect 2047 1146 2048 1147
rect 1979 1144 2048 1146
rect 1979 1143 1980 1144
rect 1974 1142 1980 1143
rect 2047 1143 2048 1144
rect 2052 1143 2053 1147
rect 2047 1142 2053 1143
rect 2126 1147 2132 1148
rect 2126 1143 2127 1147
rect 2131 1146 2132 1147
rect 2159 1147 2165 1148
rect 2159 1146 2160 1147
rect 2131 1144 2160 1146
rect 2131 1143 2132 1144
rect 2126 1142 2132 1143
rect 2159 1143 2160 1144
rect 2164 1143 2165 1147
rect 2159 1142 2165 1143
rect 2246 1147 2252 1148
rect 2246 1143 2247 1147
rect 2251 1146 2252 1147
rect 2279 1147 2285 1148
rect 2279 1146 2280 1147
rect 2251 1144 2280 1146
rect 2251 1143 2252 1144
rect 2246 1142 2252 1143
rect 2279 1143 2280 1144
rect 2284 1143 2285 1147
rect 2279 1142 2285 1143
rect 2382 1147 2389 1148
rect 2406 1147 2412 1148
rect 2382 1143 2383 1147
rect 2388 1143 2389 1147
rect 2382 1142 2389 1143
rect 1014 1138 1020 1139
rect 1238 1139 1244 1140
rect 110 1134 116 1135
rect 1238 1135 1239 1139
rect 1243 1135 1244 1139
rect 1585 1138 1587 1142
rect 1750 1139 1756 1140
rect 1750 1138 1751 1139
rect 1585 1136 1751 1138
rect 1238 1134 1244 1135
rect 1278 1135 1284 1136
rect 134 1132 140 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 134 1127 140 1128
rect 174 1132 180 1133
rect 174 1128 175 1132
rect 179 1128 180 1132
rect 174 1127 180 1128
rect 230 1132 236 1133
rect 230 1128 231 1132
rect 235 1128 236 1132
rect 230 1127 236 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 382 1132 388 1133
rect 382 1128 383 1132
rect 387 1128 388 1132
rect 382 1127 388 1128
rect 470 1132 476 1133
rect 470 1128 471 1132
rect 475 1128 476 1132
rect 470 1127 476 1128
rect 558 1132 564 1133
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 558 1127 564 1128
rect 638 1132 644 1133
rect 638 1128 639 1132
rect 643 1128 644 1132
rect 638 1127 644 1128
rect 718 1132 724 1133
rect 718 1128 719 1132
rect 723 1128 724 1132
rect 718 1127 724 1128
rect 798 1132 804 1133
rect 798 1128 799 1132
rect 803 1128 804 1132
rect 798 1127 804 1128
rect 870 1132 876 1133
rect 870 1128 871 1132
rect 875 1128 876 1132
rect 870 1127 876 1128
rect 934 1132 940 1133
rect 934 1128 935 1132
rect 939 1128 940 1132
rect 934 1127 940 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1046 1132 1052 1133
rect 1046 1128 1047 1132
rect 1051 1128 1052 1132
rect 1046 1127 1052 1128
rect 1102 1132 1108 1133
rect 1102 1128 1103 1132
rect 1107 1128 1108 1132
rect 1102 1127 1108 1128
rect 1150 1132 1156 1133
rect 1150 1128 1151 1132
rect 1155 1128 1156 1132
rect 1150 1127 1156 1128
rect 1190 1132 1196 1133
rect 1190 1128 1191 1132
rect 1195 1128 1196 1132
rect 1278 1131 1279 1135
rect 1283 1131 1284 1135
rect 1750 1135 1751 1136
rect 1755 1135 1756 1139
rect 1750 1134 1756 1135
rect 2406 1135 2412 1136
rect 1278 1130 1284 1131
rect 2406 1131 2407 1135
rect 2411 1131 2412 1135
rect 2406 1130 2412 1131
rect 1190 1127 1196 1128
rect 1558 1128 1564 1129
rect 1558 1124 1559 1128
rect 1563 1124 1564 1128
rect 1558 1123 1564 1124
rect 1598 1128 1604 1129
rect 1598 1124 1599 1128
rect 1603 1124 1604 1128
rect 1598 1123 1604 1124
rect 1638 1128 1644 1129
rect 1638 1124 1639 1128
rect 1643 1124 1644 1128
rect 1638 1123 1644 1124
rect 1678 1128 1684 1129
rect 1678 1124 1679 1128
rect 1683 1124 1684 1128
rect 1678 1123 1684 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1758 1128 1764 1129
rect 1758 1124 1759 1128
rect 1763 1124 1764 1128
rect 1758 1123 1764 1124
rect 1798 1128 1804 1129
rect 1798 1124 1799 1128
rect 1803 1124 1804 1128
rect 1798 1123 1804 1124
rect 1854 1128 1860 1129
rect 1854 1124 1855 1128
rect 1859 1124 1860 1128
rect 1854 1123 1860 1124
rect 1926 1128 1932 1129
rect 1926 1124 1927 1128
rect 1931 1124 1932 1128
rect 1926 1123 1932 1124
rect 2022 1128 2028 1129
rect 2022 1124 2023 1128
rect 2027 1124 2028 1128
rect 2022 1123 2028 1124
rect 2134 1128 2140 1129
rect 2134 1124 2135 1128
rect 2139 1124 2140 1128
rect 2134 1123 2140 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 134 1120 140 1121
rect 134 1116 135 1120
rect 139 1116 140 1120
rect 134 1115 140 1116
rect 214 1120 220 1121
rect 214 1116 215 1120
rect 219 1116 220 1120
rect 214 1115 220 1116
rect 302 1120 308 1121
rect 302 1116 303 1120
rect 307 1116 308 1120
rect 302 1115 308 1116
rect 390 1120 396 1121
rect 390 1116 391 1120
rect 395 1116 396 1120
rect 390 1115 396 1116
rect 478 1120 484 1121
rect 478 1116 479 1120
rect 483 1116 484 1120
rect 478 1115 484 1116
rect 558 1120 564 1121
rect 558 1116 559 1120
rect 563 1116 564 1120
rect 558 1115 564 1116
rect 638 1120 644 1121
rect 638 1116 639 1120
rect 643 1116 644 1120
rect 638 1115 644 1116
rect 710 1120 716 1121
rect 710 1116 711 1120
rect 715 1116 716 1120
rect 710 1115 716 1116
rect 774 1120 780 1121
rect 774 1116 775 1120
rect 779 1116 780 1120
rect 774 1115 780 1116
rect 838 1120 844 1121
rect 838 1116 839 1120
rect 843 1116 844 1120
rect 838 1115 844 1116
rect 902 1120 908 1121
rect 902 1116 903 1120
rect 907 1116 908 1120
rect 902 1115 908 1116
rect 958 1120 964 1121
rect 958 1116 959 1120
rect 963 1116 964 1120
rect 958 1115 964 1116
rect 1022 1120 1028 1121
rect 1022 1116 1023 1120
rect 1027 1116 1028 1120
rect 1022 1115 1028 1116
rect 1086 1120 1092 1121
rect 1086 1116 1087 1120
rect 1091 1116 1092 1120
rect 1086 1115 1092 1116
rect 1150 1120 1156 1121
rect 1150 1116 1151 1120
rect 1155 1116 1156 1120
rect 1150 1115 1156 1116
rect 1190 1120 1196 1121
rect 1190 1116 1191 1120
rect 1195 1116 1196 1120
rect 1190 1115 1196 1116
rect 110 1113 116 1114
rect 110 1109 111 1113
rect 115 1109 116 1113
rect 110 1108 116 1109
rect 1238 1113 1244 1114
rect 1238 1109 1239 1113
rect 1243 1109 1244 1113
rect 1238 1108 1244 1109
rect 1534 1108 1540 1109
rect 398 1107 404 1108
rect 398 1106 399 1107
rect 161 1104 399 1106
rect 161 1100 163 1104
rect 398 1103 399 1104
rect 403 1103 404 1107
rect 1214 1107 1220 1108
rect 1214 1106 1215 1107
rect 398 1102 404 1103
rect 1113 1104 1215 1106
rect 1113 1100 1115 1104
rect 1214 1103 1215 1104
rect 1219 1103 1220 1107
rect 1534 1104 1535 1108
rect 1539 1104 1540 1108
rect 1534 1103 1540 1104
rect 1598 1108 1604 1109
rect 1598 1104 1599 1108
rect 1603 1104 1604 1108
rect 1598 1103 1604 1104
rect 1662 1108 1668 1109
rect 1662 1104 1663 1108
rect 1667 1104 1668 1108
rect 1662 1103 1668 1104
rect 1726 1108 1732 1109
rect 1726 1104 1727 1108
rect 1731 1104 1732 1108
rect 1726 1103 1732 1104
rect 1790 1108 1796 1109
rect 1790 1104 1791 1108
rect 1795 1104 1796 1108
rect 1790 1103 1796 1104
rect 1854 1108 1860 1109
rect 1854 1104 1855 1108
rect 1859 1104 1860 1108
rect 1854 1103 1860 1104
rect 1910 1108 1916 1109
rect 1910 1104 1911 1108
rect 1915 1104 1916 1108
rect 1910 1103 1916 1104
rect 1966 1108 1972 1109
rect 1966 1104 1967 1108
rect 1971 1104 1972 1108
rect 1966 1103 1972 1104
rect 2022 1108 2028 1109
rect 2022 1104 2023 1108
rect 2027 1104 2028 1108
rect 2022 1103 2028 1104
rect 2078 1108 2084 1109
rect 2078 1104 2079 1108
rect 2083 1104 2084 1108
rect 2078 1103 2084 1104
rect 2134 1108 2140 1109
rect 2134 1104 2135 1108
rect 2139 1104 2140 1108
rect 2134 1103 2140 1104
rect 2190 1108 2196 1109
rect 2190 1104 2191 1108
rect 2195 1104 2196 1108
rect 2190 1103 2196 1104
rect 2254 1108 2260 1109
rect 2254 1104 2255 1108
rect 2259 1104 2260 1108
rect 2254 1103 2260 1104
rect 2318 1108 2324 1109
rect 2318 1104 2319 1108
rect 2323 1104 2324 1108
rect 2318 1103 2324 1104
rect 2358 1108 2364 1109
rect 2358 1104 2359 1108
rect 2363 1104 2364 1108
rect 2358 1103 2364 1104
rect 1214 1102 1220 1103
rect 1278 1101 1284 1102
rect 159 1099 165 1100
rect 110 1096 116 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 159 1095 160 1099
rect 164 1095 165 1099
rect 159 1094 165 1095
rect 167 1099 173 1100
rect 167 1095 168 1099
rect 172 1098 173 1099
rect 239 1099 245 1100
rect 239 1098 240 1099
rect 172 1096 240 1098
rect 172 1095 173 1096
rect 167 1094 173 1095
rect 239 1095 240 1096
rect 244 1095 245 1099
rect 239 1094 245 1095
rect 247 1099 253 1100
rect 247 1095 248 1099
rect 252 1098 253 1099
rect 327 1099 333 1100
rect 327 1098 328 1099
rect 252 1096 328 1098
rect 252 1095 253 1096
rect 247 1094 253 1095
rect 327 1095 328 1096
rect 332 1095 333 1099
rect 327 1094 333 1095
rect 335 1099 341 1100
rect 335 1095 336 1099
rect 340 1098 341 1099
rect 415 1099 421 1100
rect 415 1098 416 1099
rect 340 1096 416 1098
rect 340 1095 341 1096
rect 335 1094 341 1095
rect 415 1095 416 1096
rect 420 1095 421 1099
rect 415 1094 421 1095
rect 503 1099 509 1100
rect 503 1095 504 1099
rect 508 1098 509 1099
rect 566 1099 572 1100
rect 566 1098 567 1099
rect 508 1096 567 1098
rect 508 1095 509 1096
rect 503 1094 509 1095
rect 566 1095 567 1096
rect 571 1095 572 1099
rect 566 1094 572 1095
rect 574 1099 580 1100
rect 574 1095 575 1099
rect 579 1098 580 1099
rect 583 1099 589 1100
rect 583 1098 584 1099
rect 579 1096 584 1098
rect 579 1095 580 1096
rect 574 1094 580 1095
rect 583 1095 584 1096
rect 588 1095 589 1099
rect 583 1094 589 1095
rect 663 1099 669 1100
rect 663 1095 664 1099
rect 668 1098 669 1099
rect 726 1099 732 1100
rect 726 1098 727 1099
rect 668 1096 727 1098
rect 668 1095 669 1096
rect 663 1094 669 1095
rect 726 1095 727 1096
rect 731 1095 732 1099
rect 726 1094 732 1095
rect 735 1099 744 1100
rect 735 1095 736 1099
rect 743 1095 744 1099
rect 735 1094 744 1095
rect 799 1099 805 1100
rect 799 1095 800 1099
rect 804 1095 805 1099
rect 799 1094 805 1095
rect 807 1099 813 1100
rect 807 1095 808 1099
rect 812 1098 813 1099
rect 863 1099 869 1100
rect 863 1098 864 1099
rect 812 1096 864 1098
rect 812 1095 813 1096
rect 807 1094 813 1095
rect 863 1095 864 1096
rect 868 1095 869 1099
rect 863 1094 869 1095
rect 871 1099 877 1100
rect 871 1095 872 1099
rect 876 1098 877 1099
rect 927 1099 933 1100
rect 927 1098 928 1099
rect 876 1096 928 1098
rect 876 1095 877 1096
rect 871 1094 877 1095
rect 927 1095 928 1096
rect 932 1095 933 1099
rect 927 1094 933 1095
rect 935 1099 941 1100
rect 935 1095 936 1099
rect 940 1098 941 1099
rect 983 1099 989 1100
rect 983 1098 984 1099
rect 940 1096 984 1098
rect 940 1095 941 1096
rect 935 1094 941 1095
rect 983 1095 984 1096
rect 988 1095 989 1099
rect 983 1094 989 1095
rect 991 1099 997 1100
rect 991 1095 992 1099
rect 996 1098 997 1099
rect 1047 1099 1053 1100
rect 1047 1098 1048 1099
rect 996 1096 1048 1098
rect 996 1095 997 1096
rect 991 1094 997 1095
rect 1047 1095 1048 1096
rect 1052 1095 1053 1099
rect 1047 1094 1053 1095
rect 1111 1099 1117 1100
rect 1111 1095 1112 1099
rect 1116 1095 1117 1099
rect 1111 1094 1117 1095
rect 1119 1099 1125 1100
rect 1119 1095 1120 1099
rect 1124 1098 1125 1099
rect 1175 1099 1181 1100
rect 1175 1098 1176 1099
rect 1124 1096 1176 1098
rect 1124 1095 1125 1096
rect 1119 1094 1125 1095
rect 1175 1095 1176 1096
rect 1180 1095 1181 1099
rect 1175 1094 1181 1095
rect 1198 1099 1204 1100
rect 1198 1095 1199 1099
rect 1203 1098 1204 1099
rect 1215 1099 1221 1100
rect 1215 1098 1216 1099
rect 1203 1096 1216 1098
rect 1203 1095 1204 1096
rect 1198 1094 1204 1095
rect 1215 1095 1216 1096
rect 1220 1095 1221 1099
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1215 1094 1221 1095
rect 1238 1096 1244 1097
rect 1278 1096 1284 1097
rect 2406 1101 2412 1102
rect 2406 1097 2407 1101
rect 2411 1097 2412 1101
rect 2406 1096 2412 1097
rect 110 1091 116 1092
rect 801 1090 803 1094
rect 1238 1092 1239 1096
rect 1243 1092 1244 1096
rect 982 1091 988 1092
rect 1238 1091 1244 1092
rect 982 1090 983 1091
rect 801 1088 983 1090
rect 982 1087 983 1088
rect 987 1087 988 1091
rect 982 1086 988 1087
rect 1559 1087 1565 1088
rect 1278 1084 1284 1085
rect 1278 1080 1279 1084
rect 1283 1080 1284 1084
rect 1559 1083 1560 1087
rect 1564 1083 1565 1087
rect 1559 1082 1565 1083
rect 1567 1087 1573 1088
rect 1567 1083 1568 1087
rect 1572 1086 1573 1087
rect 1623 1087 1629 1088
rect 1623 1086 1624 1087
rect 1572 1084 1624 1086
rect 1572 1083 1573 1084
rect 1567 1082 1573 1083
rect 1623 1083 1624 1084
rect 1628 1083 1629 1087
rect 1623 1082 1629 1083
rect 1631 1087 1637 1088
rect 1631 1083 1632 1087
rect 1636 1086 1637 1087
rect 1687 1087 1693 1088
rect 1687 1086 1688 1087
rect 1636 1084 1688 1086
rect 1636 1083 1637 1084
rect 1631 1082 1637 1083
rect 1687 1083 1688 1084
rect 1692 1083 1693 1087
rect 1687 1082 1693 1083
rect 1695 1087 1701 1088
rect 1695 1083 1696 1087
rect 1700 1086 1701 1087
rect 1751 1087 1757 1088
rect 1751 1086 1752 1087
rect 1700 1084 1752 1086
rect 1700 1083 1701 1084
rect 1695 1082 1701 1083
rect 1751 1083 1752 1084
rect 1756 1083 1757 1087
rect 1751 1082 1757 1083
rect 1815 1087 1821 1088
rect 1815 1083 1816 1087
rect 1820 1083 1821 1087
rect 1815 1082 1821 1083
rect 1823 1087 1829 1088
rect 1823 1083 1824 1087
rect 1828 1086 1829 1087
rect 1879 1087 1885 1088
rect 1879 1086 1880 1087
rect 1828 1084 1880 1086
rect 1828 1083 1829 1084
rect 1823 1082 1829 1083
rect 1879 1083 1880 1084
rect 1884 1083 1885 1087
rect 1879 1082 1885 1083
rect 1887 1087 1893 1088
rect 1887 1083 1888 1087
rect 1892 1086 1893 1087
rect 1935 1087 1941 1088
rect 1935 1086 1936 1087
rect 1892 1084 1936 1086
rect 1892 1083 1893 1084
rect 1887 1082 1893 1083
rect 1935 1083 1936 1084
rect 1940 1083 1941 1087
rect 1935 1082 1941 1083
rect 1991 1087 1997 1088
rect 1991 1083 1992 1087
rect 1996 1086 1997 1087
rect 2038 1087 2044 1088
rect 1996 1084 2001 1086
rect 1996 1083 1997 1084
rect 1991 1082 1997 1083
rect 1278 1079 1284 1080
rect 1560 1078 1562 1082
rect 1758 1079 1764 1080
rect 1758 1078 1759 1079
rect 1560 1076 1759 1078
rect 1758 1075 1759 1076
rect 1763 1075 1764 1079
rect 1817 1078 1819 1082
rect 1990 1079 1996 1080
rect 1990 1078 1991 1079
rect 1817 1076 1991 1078
rect 1758 1074 1764 1075
rect 1990 1075 1991 1076
rect 1995 1075 1996 1079
rect 1999 1078 2001 1084
rect 2038 1083 2039 1087
rect 2043 1086 2044 1087
rect 2047 1087 2053 1088
rect 2047 1086 2048 1087
rect 2043 1084 2048 1086
rect 2043 1083 2044 1084
rect 2038 1082 2044 1083
rect 2047 1083 2048 1084
rect 2052 1083 2053 1087
rect 2047 1082 2053 1083
rect 2055 1087 2061 1088
rect 2055 1083 2056 1087
rect 2060 1086 2061 1087
rect 2103 1087 2109 1088
rect 2103 1086 2104 1087
rect 2060 1084 2104 1086
rect 2060 1083 2061 1084
rect 2055 1082 2061 1083
rect 2103 1083 2104 1084
rect 2108 1083 2109 1087
rect 2103 1082 2109 1083
rect 2111 1087 2117 1088
rect 2111 1083 2112 1087
rect 2116 1086 2117 1087
rect 2159 1087 2165 1088
rect 2159 1086 2160 1087
rect 2116 1084 2160 1086
rect 2116 1083 2117 1084
rect 2111 1082 2117 1083
rect 2159 1083 2160 1084
rect 2164 1083 2165 1087
rect 2159 1082 2165 1083
rect 2215 1087 2224 1088
rect 2215 1083 2216 1087
rect 2223 1083 2224 1087
rect 2215 1082 2224 1083
rect 2226 1087 2232 1088
rect 2226 1083 2227 1087
rect 2231 1086 2232 1087
rect 2279 1087 2285 1088
rect 2279 1086 2280 1087
rect 2231 1084 2280 1086
rect 2231 1083 2232 1084
rect 2226 1082 2232 1083
rect 2279 1083 2280 1084
rect 2284 1083 2285 1087
rect 2279 1082 2285 1083
rect 2287 1087 2293 1088
rect 2287 1083 2288 1087
rect 2292 1086 2293 1087
rect 2343 1087 2349 1088
rect 2343 1086 2344 1087
rect 2292 1084 2344 1086
rect 2292 1083 2293 1084
rect 2287 1082 2293 1083
rect 2343 1083 2344 1084
rect 2348 1083 2349 1087
rect 2343 1082 2349 1083
rect 2366 1087 2372 1088
rect 2366 1083 2367 1087
rect 2371 1086 2372 1087
rect 2383 1087 2389 1088
rect 2383 1086 2384 1087
rect 2371 1084 2384 1086
rect 2371 1083 2372 1084
rect 2366 1082 2372 1083
rect 2383 1083 2384 1084
rect 2388 1083 2389 1087
rect 2383 1082 2389 1083
rect 2406 1084 2412 1085
rect 2406 1080 2407 1084
rect 2411 1080 2412 1084
rect 2146 1079 2152 1080
rect 2406 1079 2412 1080
rect 2146 1078 2147 1079
rect 1999 1076 2147 1078
rect 1990 1074 1996 1075
rect 2146 1075 2147 1076
rect 2151 1075 2152 1079
rect 2146 1074 2152 1075
rect 134 1073 140 1074
rect 134 1069 135 1073
rect 139 1069 140 1073
rect 134 1068 140 1069
rect 214 1073 220 1074
rect 214 1069 215 1073
rect 219 1069 220 1073
rect 214 1068 220 1069
rect 302 1073 308 1074
rect 302 1069 303 1073
rect 307 1069 308 1073
rect 302 1068 308 1069
rect 390 1073 396 1074
rect 390 1069 391 1073
rect 395 1069 396 1073
rect 390 1068 396 1069
rect 478 1073 484 1074
rect 478 1069 479 1073
rect 483 1069 484 1073
rect 478 1068 484 1069
rect 558 1073 564 1074
rect 558 1069 559 1073
rect 563 1069 564 1073
rect 558 1068 564 1069
rect 638 1073 644 1074
rect 638 1069 639 1073
rect 643 1069 644 1073
rect 638 1068 644 1069
rect 710 1073 716 1074
rect 710 1069 711 1073
rect 715 1069 716 1073
rect 710 1068 716 1069
rect 774 1073 780 1074
rect 774 1069 775 1073
rect 779 1069 780 1073
rect 774 1068 780 1069
rect 838 1073 844 1074
rect 838 1069 839 1073
rect 843 1069 844 1073
rect 838 1068 844 1069
rect 902 1073 908 1074
rect 902 1069 903 1073
rect 907 1069 908 1073
rect 902 1068 908 1069
rect 958 1073 964 1074
rect 958 1069 959 1073
rect 963 1069 964 1073
rect 958 1068 964 1069
rect 1022 1073 1028 1074
rect 1022 1069 1023 1073
rect 1027 1069 1028 1073
rect 1022 1068 1028 1069
rect 1086 1073 1092 1074
rect 1086 1069 1087 1073
rect 1091 1069 1092 1073
rect 1086 1068 1092 1069
rect 1150 1073 1156 1074
rect 1150 1069 1151 1073
rect 1155 1069 1156 1073
rect 1150 1068 1156 1069
rect 1190 1073 1196 1074
rect 1190 1069 1191 1073
rect 1195 1069 1196 1073
rect 1190 1068 1196 1069
rect 159 1067 165 1068
rect 159 1063 160 1067
rect 164 1066 165 1067
rect 167 1067 173 1068
rect 167 1066 168 1067
rect 164 1064 168 1066
rect 164 1063 165 1064
rect 159 1062 165 1063
rect 167 1063 168 1064
rect 172 1063 173 1067
rect 167 1062 173 1063
rect 239 1067 245 1068
rect 239 1063 240 1067
rect 244 1066 245 1067
rect 247 1067 253 1068
rect 247 1066 248 1067
rect 244 1064 248 1066
rect 244 1063 245 1064
rect 239 1062 245 1063
rect 247 1063 248 1064
rect 252 1063 253 1067
rect 247 1062 253 1063
rect 327 1067 333 1068
rect 327 1063 328 1067
rect 332 1066 333 1067
rect 335 1067 341 1068
rect 335 1066 336 1067
rect 332 1064 336 1066
rect 332 1063 333 1064
rect 327 1062 333 1063
rect 335 1063 336 1064
rect 340 1063 341 1067
rect 415 1067 421 1068
rect 415 1066 416 1067
rect 335 1062 341 1063
rect 344 1064 416 1066
rect 266 1059 272 1060
rect 266 1055 267 1059
rect 271 1058 272 1059
rect 344 1058 346 1064
rect 415 1063 416 1064
rect 420 1063 421 1067
rect 415 1062 421 1063
rect 498 1067 509 1068
rect 498 1063 499 1067
rect 503 1063 504 1067
rect 508 1063 509 1067
rect 498 1062 509 1063
rect 566 1067 572 1068
rect 566 1063 567 1067
rect 571 1066 572 1067
rect 583 1067 589 1068
rect 583 1066 584 1067
rect 571 1064 584 1066
rect 571 1063 572 1064
rect 566 1062 572 1063
rect 583 1063 584 1064
rect 588 1063 589 1067
rect 583 1062 589 1063
rect 610 1067 616 1068
rect 610 1063 611 1067
rect 615 1066 616 1067
rect 663 1067 669 1068
rect 663 1066 664 1067
rect 615 1064 664 1066
rect 615 1063 616 1064
rect 610 1062 616 1063
rect 663 1063 664 1064
rect 668 1063 669 1067
rect 663 1062 669 1063
rect 726 1067 732 1068
rect 726 1063 727 1067
rect 731 1066 732 1067
rect 735 1067 741 1068
rect 735 1066 736 1067
rect 731 1064 736 1066
rect 731 1063 732 1064
rect 726 1062 732 1063
rect 735 1063 736 1064
rect 740 1063 741 1067
rect 735 1062 741 1063
rect 799 1067 805 1068
rect 799 1063 800 1067
rect 804 1066 805 1067
rect 807 1067 813 1068
rect 807 1066 808 1067
rect 804 1064 808 1066
rect 804 1063 805 1064
rect 799 1062 805 1063
rect 807 1063 808 1064
rect 812 1063 813 1067
rect 807 1062 813 1063
rect 863 1067 869 1068
rect 863 1063 864 1067
rect 868 1066 869 1067
rect 871 1067 877 1068
rect 871 1066 872 1067
rect 868 1064 872 1066
rect 868 1063 869 1064
rect 863 1062 869 1063
rect 871 1063 872 1064
rect 876 1063 877 1067
rect 871 1062 877 1063
rect 927 1067 933 1068
rect 927 1063 928 1067
rect 932 1066 933 1067
rect 935 1067 941 1068
rect 935 1066 936 1067
rect 932 1064 936 1066
rect 932 1063 933 1064
rect 927 1062 933 1063
rect 935 1063 936 1064
rect 940 1063 941 1067
rect 935 1062 941 1063
rect 983 1067 989 1068
rect 983 1063 984 1067
rect 988 1066 989 1067
rect 991 1067 997 1068
rect 991 1066 992 1067
rect 988 1064 992 1066
rect 988 1063 989 1064
rect 983 1062 989 1063
rect 991 1063 992 1064
rect 996 1063 997 1067
rect 991 1062 997 1063
rect 1014 1067 1020 1068
rect 1014 1063 1015 1067
rect 1019 1066 1020 1067
rect 1047 1067 1053 1068
rect 1047 1066 1048 1067
rect 1019 1064 1048 1066
rect 1019 1063 1020 1064
rect 1014 1062 1020 1063
rect 1047 1063 1048 1064
rect 1052 1063 1053 1067
rect 1047 1062 1053 1063
rect 1111 1067 1117 1068
rect 1111 1063 1112 1067
rect 1116 1066 1117 1067
rect 1119 1067 1125 1068
rect 1119 1066 1120 1067
rect 1116 1064 1120 1066
rect 1116 1063 1117 1064
rect 1111 1062 1117 1063
rect 1119 1063 1120 1064
rect 1124 1063 1125 1067
rect 1119 1062 1125 1063
rect 1175 1067 1181 1068
rect 1175 1063 1176 1067
rect 1180 1066 1181 1067
rect 1198 1067 1204 1068
rect 1198 1066 1199 1067
rect 1180 1064 1199 1066
rect 1180 1063 1181 1064
rect 1175 1062 1181 1063
rect 1198 1063 1199 1064
rect 1203 1063 1204 1067
rect 1198 1062 1204 1063
rect 1214 1067 1221 1068
rect 1214 1063 1215 1067
rect 1220 1063 1221 1067
rect 1214 1062 1221 1063
rect 271 1056 346 1058
rect 1534 1061 1540 1062
rect 1534 1057 1535 1061
rect 1539 1057 1540 1061
rect 1534 1056 1540 1057
rect 1598 1061 1604 1062
rect 1598 1057 1599 1061
rect 1603 1057 1604 1061
rect 1598 1056 1604 1057
rect 1662 1061 1668 1062
rect 1662 1057 1663 1061
rect 1667 1057 1668 1061
rect 1662 1056 1668 1057
rect 1726 1061 1732 1062
rect 1726 1057 1727 1061
rect 1731 1057 1732 1061
rect 1726 1056 1732 1057
rect 1790 1061 1796 1062
rect 1790 1057 1791 1061
rect 1795 1057 1796 1061
rect 1790 1056 1796 1057
rect 1854 1061 1860 1062
rect 1854 1057 1855 1061
rect 1859 1057 1860 1061
rect 1854 1056 1860 1057
rect 1910 1061 1916 1062
rect 1910 1057 1911 1061
rect 1915 1057 1916 1061
rect 1910 1056 1916 1057
rect 1966 1061 1972 1062
rect 1966 1057 1967 1061
rect 1971 1057 1972 1061
rect 1966 1056 1972 1057
rect 2022 1061 2028 1062
rect 2022 1057 2023 1061
rect 2027 1057 2028 1061
rect 2022 1056 2028 1057
rect 2078 1061 2084 1062
rect 2078 1057 2079 1061
rect 2083 1057 2084 1061
rect 2078 1056 2084 1057
rect 2134 1061 2140 1062
rect 2134 1057 2135 1061
rect 2139 1057 2140 1061
rect 2134 1056 2140 1057
rect 2190 1061 2196 1062
rect 2190 1057 2191 1061
rect 2195 1057 2196 1061
rect 2190 1056 2196 1057
rect 2254 1061 2260 1062
rect 2254 1057 2255 1061
rect 2259 1057 2260 1061
rect 2254 1056 2260 1057
rect 2318 1061 2324 1062
rect 2318 1057 2319 1061
rect 2323 1057 2324 1061
rect 2318 1056 2324 1057
rect 2358 1061 2364 1062
rect 2358 1057 2359 1061
rect 2363 1057 2364 1061
rect 2358 1056 2364 1057
rect 271 1055 272 1056
rect 266 1054 272 1055
rect 1559 1055 1565 1056
rect 1559 1051 1560 1055
rect 1564 1054 1565 1055
rect 1567 1055 1573 1056
rect 1567 1054 1568 1055
rect 1564 1052 1568 1054
rect 1564 1051 1565 1052
rect 1559 1050 1565 1051
rect 1567 1051 1568 1052
rect 1572 1051 1573 1055
rect 1567 1050 1573 1051
rect 1623 1055 1629 1056
rect 1623 1051 1624 1055
rect 1628 1054 1629 1055
rect 1631 1055 1637 1056
rect 1631 1054 1632 1055
rect 1628 1052 1632 1054
rect 1628 1051 1629 1052
rect 1623 1050 1629 1051
rect 1631 1051 1632 1052
rect 1636 1051 1637 1055
rect 1631 1050 1637 1051
rect 1687 1055 1693 1056
rect 1687 1051 1688 1055
rect 1692 1054 1693 1055
rect 1695 1055 1701 1056
rect 1695 1054 1696 1055
rect 1692 1052 1696 1054
rect 1692 1051 1693 1052
rect 1687 1050 1693 1051
rect 1695 1051 1696 1052
rect 1700 1051 1701 1055
rect 1695 1050 1701 1051
rect 1750 1055 1757 1056
rect 1750 1051 1751 1055
rect 1756 1051 1757 1055
rect 1750 1050 1757 1051
rect 1815 1055 1821 1056
rect 1815 1051 1816 1055
rect 1820 1054 1821 1055
rect 1823 1055 1829 1056
rect 1823 1054 1824 1055
rect 1820 1052 1824 1054
rect 1820 1051 1821 1052
rect 1815 1050 1821 1051
rect 1823 1051 1824 1052
rect 1828 1051 1829 1055
rect 1823 1050 1829 1051
rect 1879 1055 1885 1056
rect 1879 1051 1880 1055
rect 1884 1054 1885 1055
rect 1887 1055 1893 1056
rect 1887 1054 1888 1055
rect 1884 1052 1888 1054
rect 1884 1051 1885 1052
rect 1879 1050 1885 1051
rect 1887 1051 1888 1052
rect 1892 1051 1893 1055
rect 1887 1050 1893 1051
rect 1935 1055 1941 1056
rect 1935 1051 1936 1055
rect 1940 1054 1941 1055
rect 1974 1055 1980 1056
rect 1974 1054 1975 1055
rect 1940 1052 1975 1054
rect 1940 1051 1941 1052
rect 1935 1050 1941 1051
rect 1974 1051 1975 1052
rect 1979 1051 1980 1055
rect 1974 1050 1980 1051
rect 1990 1055 1997 1056
rect 1990 1051 1991 1055
rect 1996 1051 1997 1055
rect 1990 1050 1997 1051
rect 2047 1055 2053 1056
rect 2047 1051 2048 1055
rect 2052 1054 2053 1055
rect 2055 1055 2061 1056
rect 2055 1054 2056 1055
rect 2052 1052 2056 1054
rect 2052 1051 2053 1052
rect 2047 1050 2053 1051
rect 2055 1051 2056 1052
rect 2060 1051 2061 1055
rect 2055 1050 2061 1051
rect 2103 1055 2109 1056
rect 2103 1051 2104 1055
rect 2108 1054 2109 1055
rect 2111 1055 2117 1056
rect 2111 1054 2112 1055
rect 2108 1052 2112 1054
rect 2108 1051 2109 1052
rect 2103 1050 2109 1051
rect 2111 1051 2112 1052
rect 2116 1051 2117 1055
rect 2111 1050 2117 1051
rect 2146 1055 2152 1056
rect 2146 1051 2147 1055
rect 2151 1054 2152 1055
rect 2159 1055 2165 1056
rect 2159 1054 2160 1055
rect 2151 1052 2160 1054
rect 2151 1051 2152 1052
rect 2146 1050 2152 1051
rect 2159 1051 2160 1052
rect 2164 1051 2165 1055
rect 2159 1050 2165 1051
rect 2215 1055 2221 1056
rect 2215 1051 2216 1055
rect 2220 1054 2221 1055
rect 2226 1055 2232 1056
rect 2226 1054 2227 1055
rect 2220 1052 2227 1054
rect 2220 1051 2221 1052
rect 2215 1050 2221 1051
rect 2226 1051 2227 1052
rect 2231 1051 2232 1055
rect 2226 1050 2232 1051
rect 2279 1055 2285 1056
rect 2279 1051 2280 1055
rect 2284 1054 2285 1055
rect 2287 1055 2293 1056
rect 2287 1054 2288 1055
rect 2284 1052 2288 1054
rect 2284 1051 2285 1052
rect 2279 1050 2285 1051
rect 2287 1051 2288 1052
rect 2292 1051 2293 1055
rect 2287 1050 2293 1051
rect 2343 1055 2349 1056
rect 2343 1051 2344 1055
rect 2348 1054 2349 1055
rect 2366 1055 2372 1056
rect 2366 1054 2367 1055
rect 2348 1052 2367 1054
rect 2348 1051 2349 1052
rect 2343 1050 2349 1051
rect 2366 1051 2367 1052
rect 2371 1051 2372 1055
rect 2366 1050 2372 1051
rect 2382 1055 2389 1056
rect 2382 1051 2383 1055
rect 2388 1051 2389 1055
rect 2382 1050 2389 1051
rect 574 1047 580 1048
rect 574 1046 575 1047
rect 559 1045 575 1046
rect 223 1043 232 1044
rect 198 1039 204 1040
rect 198 1035 199 1039
rect 203 1035 204 1039
rect 223 1039 224 1043
rect 231 1039 232 1043
rect 263 1043 269 1044
rect 223 1038 232 1039
rect 238 1039 244 1040
rect 198 1034 204 1035
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 263 1039 264 1043
rect 268 1042 269 1043
rect 278 1043 284 1044
rect 278 1042 279 1043
rect 268 1040 279 1042
rect 268 1039 269 1040
rect 263 1038 269 1039
rect 278 1039 279 1040
rect 283 1039 284 1043
rect 311 1043 317 1044
rect 278 1038 284 1039
rect 286 1039 292 1040
rect 238 1034 244 1035
rect 286 1035 287 1039
rect 291 1035 292 1039
rect 311 1039 312 1043
rect 316 1042 317 1043
rect 334 1043 340 1044
rect 334 1042 335 1043
rect 316 1040 335 1042
rect 316 1039 317 1040
rect 311 1038 317 1039
rect 334 1039 335 1040
rect 339 1039 340 1043
rect 367 1043 373 1044
rect 334 1038 340 1039
rect 342 1039 348 1040
rect 286 1034 292 1035
rect 342 1035 343 1039
rect 347 1035 348 1039
rect 367 1039 368 1043
rect 372 1042 373 1043
rect 382 1043 388 1044
rect 382 1042 383 1043
rect 372 1040 383 1042
rect 372 1039 373 1040
rect 367 1038 373 1039
rect 382 1039 383 1040
rect 387 1039 388 1043
rect 406 1043 412 1044
rect 382 1038 388 1039
rect 390 1039 396 1040
rect 342 1034 348 1035
rect 390 1035 391 1039
rect 395 1035 396 1039
rect 406 1039 407 1043
rect 411 1042 412 1043
rect 415 1043 421 1044
rect 415 1042 416 1043
rect 411 1040 416 1042
rect 411 1039 412 1040
rect 406 1038 412 1039
rect 415 1039 416 1040
rect 420 1039 421 1043
rect 463 1043 469 1044
rect 415 1038 421 1039
rect 438 1039 444 1040
rect 390 1034 396 1035
rect 438 1035 439 1039
rect 443 1035 444 1039
rect 463 1039 464 1043
rect 468 1042 469 1043
rect 478 1043 484 1044
rect 478 1042 479 1043
rect 468 1040 479 1042
rect 468 1039 469 1040
rect 463 1038 469 1039
rect 478 1039 479 1040
rect 483 1039 484 1043
rect 511 1043 517 1044
rect 478 1038 484 1039
rect 486 1039 492 1040
rect 438 1034 444 1035
rect 486 1035 487 1039
rect 491 1035 492 1039
rect 511 1039 512 1043
rect 516 1042 517 1043
rect 526 1043 532 1044
rect 526 1042 527 1043
rect 516 1040 527 1042
rect 516 1039 517 1040
rect 511 1038 517 1039
rect 526 1039 527 1040
rect 531 1039 532 1043
rect 559 1041 560 1045
rect 564 1044 575 1045
rect 564 1041 565 1044
rect 574 1043 575 1044
rect 579 1043 580 1047
rect 574 1042 580 1043
rect 607 1043 613 1044
rect 559 1040 565 1041
rect 526 1038 532 1039
rect 534 1039 540 1040
rect 486 1034 492 1035
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 582 1039 588 1040
rect 582 1035 583 1039
rect 587 1035 588 1039
rect 607 1039 608 1043
rect 612 1042 613 1043
rect 622 1043 628 1044
rect 622 1042 623 1043
rect 612 1040 623 1042
rect 612 1039 613 1040
rect 607 1038 613 1039
rect 622 1039 623 1040
rect 627 1039 628 1043
rect 655 1043 661 1044
rect 622 1038 628 1039
rect 630 1039 636 1040
rect 582 1034 588 1035
rect 630 1035 631 1039
rect 635 1035 636 1039
rect 655 1039 656 1043
rect 660 1042 661 1043
rect 663 1043 669 1044
rect 663 1042 664 1043
rect 660 1040 664 1042
rect 660 1039 661 1040
rect 655 1038 661 1039
rect 663 1039 664 1040
rect 668 1039 669 1043
rect 703 1043 709 1044
rect 663 1038 669 1039
rect 678 1039 684 1040
rect 630 1034 636 1035
rect 678 1035 679 1039
rect 683 1035 684 1039
rect 703 1039 704 1043
rect 708 1042 709 1043
rect 718 1043 724 1044
rect 718 1042 719 1043
rect 708 1040 719 1042
rect 708 1039 709 1040
rect 703 1038 709 1039
rect 718 1039 719 1040
rect 723 1039 724 1043
rect 751 1043 757 1044
rect 718 1038 724 1039
rect 726 1039 732 1040
rect 678 1034 684 1035
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 751 1039 752 1043
rect 756 1042 757 1043
rect 774 1043 780 1044
rect 774 1042 775 1043
rect 756 1040 775 1042
rect 756 1039 757 1040
rect 751 1038 757 1039
rect 774 1039 775 1040
rect 779 1039 780 1043
rect 807 1043 813 1044
rect 774 1038 780 1039
rect 782 1039 788 1040
rect 726 1034 732 1035
rect 782 1035 783 1039
rect 787 1035 788 1039
rect 807 1039 808 1043
rect 812 1042 813 1043
rect 830 1043 836 1044
rect 830 1042 831 1043
rect 812 1040 831 1042
rect 812 1039 813 1040
rect 807 1038 813 1039
rect 830 1039 831 1040
rect 835 1039 836 1043
rect 863 1043 869 1044
rect 830 1038 836 1039
rect 838 1039 844 1040
rect 782 1034 788 1035
rect 838 1035 839 1039
rect 843 1035 844 1039
rect 863 1039 864 1043
rect 868 1042 869 1043
rect 886 1043 892 1044
rect 886 1042 887 1043
rect 868 1040 887 1042
rect 868 1039 869 1040
rect 863 1038 869 1039
rect 886 1039 887 1040
rect 891 1039 892 1043
rect 919 1043 925 1044
rect 886 1038 892 1039
rect 894 1039 900 1040
rect 838 1034 844 1035
rect 894 1035 895 1039
rect 899 1035 900 1039
rect 919 1039 920 1043
rect 924 1042 925 1043
rect 950 1043 956 1044
rect 950 1042 951 1043
rect 924 1040 951 1042
rect 924 1039 925 1040
rect 919 1038 925 1039
rect 950 1039 951 1040
rect 955 1039 956 1043
rect 982 1043 989 1044
rect 950 1038 956 1039
rect 958 1039 964 1040
rect 894 1034 900 1035
rect 958 1035 959 1039
rect 963 1035 964 1039
rect 982 1039 983 1043
rect 988 1039 989 1043
rect 1047 1043 1053 1044
rect 982 1038 989 1039
rect 1022 1039 1028 1040
rect 958 1034 964 1035
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1047 1039 1048 1043
rect 1052 1042 1053 1043
rect 1078 1043 1084 1044
rect 1078 1042 1079 1043
rect 1052 1040 1079 1042
rect 1052 1039 1053 1040
rect 1047 1038 1053 1039
rect 1078 1039 1079 1040
rect 1083 1039 1084 1043
rect 1110 1043 1117 1044
rect 1078 1038 1084 1039
rect 1086 1039 1092 1040
rect 1022 1034 1028 1035
rect 1086 1035 1087 1039
rect 1091 1035 1092 1039
rect 1110 1039 1111 1043
rect 1116 1039 1117 1043
rect 1166 1043 1172 1044
rect 1110 1038 1117 1039
rect 1150 1039 1156 1040
rect 1086 1034 1092 1035
rect 1150 1035 1151 1039
rect 1155 1035 1156 1039
rect 1166 1039 1167 1043
rect 1171 1042 1172 1043
rect 1175 1043 1181 1044
rect 1175 1042 1176 1043
rect 1171 1040 1176 1042
rect 1171 1039 1172 1040
rect 1166 1038 1172 1039
rect 1175 1039 1176 1040
rect 1180 1039 1181 1043
rect 1202 1043 1208 1044
rect 1175 1038 1181 1039
rect 1190 1039 1196 1040
rect 1150 1034 1156 1035
rect 1190 1035 1191 1039
rect 1195 1035 1196 1039
rect 1202 1039 1203 1043
rect 1207 1042 1208 1043
rect 1215 1043 1221 1044
rect 1215 1042 1216 1043
rect 1207 1040 1216 1042
rect 1207 1039 1208 1040
rect 1202 1038 1208 1039
rect 1215 1039 1216 1040
rect 1220 1039 1221 1043
rect 1215 1038 1221 1039
rect 1190 1034 1196 1035
rect 1934 1027 1940 1028
rect 1934 1026 1935 1027
rect 1912 1024 1935 1026
rect 1527 1023 1533 1024
rect 266 1019 272 1020
rect 266 1018 267 1019
rect 110 1016 116 1017
rect 110 1012 111 1016
rect 115 1012 116 1016
rect 228 1016 267 1018
rect 228 1012 230 1016
rect 266 1015 267 1016
rect 271 1015 272 1019
rect 1166 1019 1172 1020
rect 1166 1018 1167 1019
rect 266 1014 272 1015
rect 1049 1016 1167 1018
rect 1049 1012 1051 1016
rect 1166 1015 1167 1016
rect 1171 1015 1172 1019
rect 1502 1019 1508 1020
rect 1166 1014 1172 1015
rect 1238 1016 1244 1017
rect 1238 1012 1239 1016
rect 1243 1012 1244 1016
rect 1502 1015 1503 1019
rect 1507 1015 1508 1019
rect 1527 1019 1528 1023
rect 1532 1022 1533 1023
rect 1614 1023 1620 1024
rect 1614 1022 1615 1023
rect 1532 1020 1615 1022
rect 1532 1019 1533 1020
rect 1527 1018 1533 1019
rect 1614 1019 1615 1020
rect 1619 1019 1620 1023
rect 1647 1023 1653 1024
rect 1614 1018 1620 1019
rect 1622 1019 1628 1020
rect 1502 1014 1508 1015
rect 1622 1015 1623 1019
rect 1627 1015 1628 1019
rect 1647 1019 1648 1023
rect 1652 1022 1653 1023
rect 1726 1023 1732 1024
rect 1726 1022 1727 1023
rect 1652 1020 1727 1022
rect 1652 1019 1653 1020
rect 1647 1018 1653 1019
rect 1726 1019 1727 1020
rect 1731 1019 1732 1023
rect 1758 1023 1765 1024
rect 1726 1018 1732 1019
rect 1734 1019 1740 1020
rect 1622 1014 1628 1015
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1758 1019 1759 1023
rect 1764 1019 1765 1023
rect 1855 1023 1861 1024
rect 1758 1018 1765 1019
rect 1830 1019 1836 1020
rect 1734 1014 1740 1015
rect 1830 1015 1831 1019
rect 1835 1015 1836 1019
rect 1855 1019 1856 1023
rect 1860 1022 1861 1023
rect 1912 1022 1914 1024
rect 1934 1023 1935 1024
rect 1939 1023 1940 1027
rect 2038 1027 2044 1028
rect 2038 1026 2039 1027
rect 2023 1025 2039 1026
rect 1934 1022 1940 1023
rect 1943 1023 1949 1024
rect 1860 1020 1914 1022
rect 1860 1019 1861 1020
rect 1855 1018 1861 1019
rect 1918 1019 1924 1020
rect 1830 1014 1836 1015
rect 1918 1015 1919 1019
rect 1923 1015 1924 1019
rect 1943 1019 1944 1023
rect 1948 1022 1949 1023
rect 1967 1023 1973 1024
rect 1967 1022 1968 1023
rect 1948 1020 1968 1022
rect 1948 1019 1949 1020
rect 1943 1018 1949 1019
rect 1967 1019 1968 1020
rect 1972 1019 1973 1023
rect 2023 1021 2024 1025
rect 2028 1024 2039 1025
rect 2028 1021 2029 1024
rect 2038 1023 2039 1024
rect 2043 1023 2044 1027
rect 2038 1022 2044 1023
rect 2082 1023 2088 1024
rect 2023 1020 2029 1021
rect 1967 1018 1973 1019
rect 1998 1019 2004 1020
rect 1918 1014 1924 1015
rect 1998 1015 1999 1019
rect 2003 1015 2004 1019
rect 1998 1014 2004 1015
rect 2070 1019 2076 1020
rect 2070 1015 2071 1019
rect 2075 1015 2076 1019
rect 2082 1019 2083 1023
rect 2087 1022 2088 1023
rect 2095 1023 2101 1024
rect 2095 1022 2096 1023
rect 2087 1020 2096 1022
rect 2087 1019 2088 1020
rect 2082 1018 2088 1019
rect 2095 1019 2096 1020
rect 2100 1019 2101 1023
rect 2167 1023 2173 1024
rect 2095 1018 2101 1019
rect 2142 1019 2148 1020
rect 2070 1014 2076 1015
rect 2142 1015 2143 1019
rect 2147 1015 2148 1019
rect 2167 1019 2168 1023
rect 2172 1022 2173 1023
rect 2198 1023 2204 1024
rect 2198 1022 2199 1023
rect 2172 1020 2199 1022
rect 2172 1019 2173 1020
rect 2167 1018 2173 1019
rect 2198 1019 2199 1020
rect 2203 1019 2204 1023
rect 2231 1023 2237 1024
rect 2198 1018 2204 1019
rect 2206 1019 2212 1020
rect 2142 1014 2148 1015
rect 2206 1015 2207 1019
rect 2211 1015 2212 1019
rect 2231 1019 2232 1023
rect 2236 1022 2237 1023
rect 2270 1023 2276 1024
rect 2270 1022 2271 1023
rect 2236 1020 2271 1022
rect 2236 1019 2237 1020
rect 2231 1018 2237 1019
rect 2270 1019 2271 1020
rect 2275 1019 2276 1023
rect 2290 1023 2296 1024
rect 2270 1018 2276 1019
rect 2278 1019 2284 1020
rect 2206 1014 2212 1015
rect 2278 1015 2279 1019
rect 2283 1015 2284 1019
rect 2290 1019 2291 1023
rect 2295 1022 2296 1023
rect 2303 1023 2309 1024
rect 2303 1022 2304 1023
rect 2295 1020 2304 1022
rect 2295 1019 2296 1020
rect 2290 1018 2296 1019
rect 2303 1019 2304 1020
rect 2308 1019 2309 1023
rect 2303 1018 2309 1019
rect 2278 1014 2284 1015
rect 110 1011 116 1012
rect 223 1011 230 1012
rect 223 1007 224 1011
rect 228 1008 230 1011
rect 234 1011 240 1012
rect 228 1007 229 1008
rect 223 1006 229 1007
rect 234 1007 235 1011
rect 239 1010 240 1011
rect 263 1011 269 1012
rect 263 1010 264 1011
rect 239 1008 264 1010
rect 239 1007 240 1008
rect 234 1006 240 1007
rect 263 1007 264 1008
rect 268 1007 269 1011
rect 263 1006 269 1007
rect 278 1011 284 1012
rect 278 1007 279 1011
rect 283 1010 284 1011
rect 311 1011 317 1012
rect 311 1010 312 1011
rect 283 1008 312 1010
rect 283 1007 284 1008
rect 278 1006 284 1007
rect 311 1007 312 1008
rect 316 1007 317 1011
rect 311 1006 317 1007
rect 334 1011 340 1012
rect 334 1007 335 1011
rect 339 1010 340 1011
rect 367 1011 373 1012
rect 367 1010 368 1011
rect 339 1008 368 1010
rect 339 1007 340 1008
rect 334 1006 340 1007
rect 367 1007 368 1008
rect 372 1007 373 1011
rect 367 1006 373 1007
rect 382 1011 388 1012
rect 382 1007 383 1011
rect 387 1010 388 1011
rect 415 1011 421 1012
rect 415 1010 416 1011
rect 387 1008 416 1010
rect 387 1007 388 1008
rect 382 1006 388 1007
rect 415 1007 416 1008
rect 420 1007 421 1011
rect 415 1006 421 1007
rect 463 1011 469 1012
rect 463 1007 464 1011
rect 468 1007 469 1011
rect 463 1006 469 1007
rect 478 1011 484 1012
rect 478 1007 479 1011
rect 483 1010 484 1011
rect 511 1011 517 1012
rect 511 1010 512 1011
rect 483 1008 512 1010
rect 483 1007 484 1008
rect 478 1006 484 1007
rect 511 1007 512 1008
rect 516 1007 517 1011
rect 511 1006 517 1007
rect 526 1011 532 1012
rect 526 1007 527 1011
rect 531 1010 532 1011
rect 559 1011 565 1012
rect 559 1010 560 1011
rect 531 1008 560 1010
rect 531 1007 532 1008
rect 526 1006 532 1007
rect 559 1007 560 1008
rect 564 1007 565 1011
rect 559 1006 565 1007
rect 607 1011 616 1012
rect 607 1007 608 1011
rect 615 1007 616 1011
rect 607 1006 616 1007
rect 622 1011 628 1012
rect 622 1007 623 1011
rect 627 1010 628 1011
rect 655 1011 661 1012
rect 655 1010 656 1011
rect 627 1008 656 1010
rect 627 1007 628 1008
rect 622 1006 628 1007
rect 655 1007 656 1008
rect 660 1007 661 1011
rect 655 1006 661 1007
rect 663 1011 669 1012
rect 663 1007 664 1011
rect 668 1010 669 1011
rect 703 1011 709 1012
rect 703 1010 704 1011
rect 668 1008 704 1010
rect 668 1007 669 1008
rect 663 1006 669 1007
rect 703 1007 704 1008
rect 708 1007 709 1011
rect 703 1006 709 1007
rect 718 1011 724 1012
rect 718 1007 719 1011
rect 723 1010 724 1011
rect 751 1011 757 1012
rect 751 1010 752 1011
rect 723 1008 752 1010
rect 723 1007 724 1008
rect 718 1006 724 1007
rect 751 1007 752 1008
rect 756 1007 757 1011
rect 751 1006 757 1007
rect 774 1011 780 1012
rect 774 1007 775 1011
rect 779 1010 780 1011
rect 807 1011 813 1012
rect 807 1010 808 1011
rect 779 1008 808 1010
rect 779 1007 780 1008
rect 774 1006 780 1007
rect 807 1007 808 1008
rect 812 1007 813 1011
rect 807 1006 813 1007
rect 830 1011 836 1012
rect 830 1007 831 1011
rect 835 1010 836 1011
rect 863 1011 869 1012
rect 863 1010 864 1011
rect 835 1008 864 1010
rect 835 1007 836 1008
rect 830 1006 836 1007
rect 863 1007 864 1008
rect 868 1007 869 1011
rect 863 1006 869 1007
rect 886 1011 892 1012
rect 886 1007 887 1011
rect 891 1010 892 1011
rect 919 1011 925 1012
rect 919 1010 920 1011
rect 891 1008 920 1010
rect 891 1007 892 1008
rect 886 1006 892 1007
rect 919 1007 920 1008
rect 924 1007 925 1011
rect 919 1006 925 1007
rect 950 1011 956 1012
rect 950 1007 951 1011
rect 955 1010 956 1011
rect 983 1011 989 1012
rect 983 1010 984 1011
rect 955 1008 984 1010
rect 955 1007 956 1008
rect 950 1006 956 1007
rect 983 1007 984 1008
rect 988 1007 989 1011
rect 983 1006 989 1007
rect 1047 1011 1053 1012
rect 1047 1007 1048 1011
rect 1052 1007 1053 1011
rect 1047 1006 1053 1007
rect 1078 1011 1084 1012
rect 1078 1007 1079 1011
rect 1083 1010 1084 1011
rect 1111 1011 1117 1012
rect 1111 1010 1112 1011
rect 1083 1008 1112 1010
rect 1083 1007 1084 1008
rect 1078 1006 1084 1007
rect 1111 1007 1112 1008
rect 1116 1007 1117 1011
rect 1111 1006 1117 1007
rect 1175 1011 1181 1012
rect 1175 1007 1176 1011
rect 1180 1010 1181 1011
rect 1202 1011 1208 1012
rect 1202 1010 1203 1011
rect 1180 1008 1203 1010
rect 1180 1007 1181 1008
rect 1175 1006 1181 1007
rect 1202 1007 1203 1008
rect 1207 1007 1208 1011
rect 1202 1006 1208 1007
rect 1214 1011 1221 1012
rect 1238 1011 1244 1012
rect 1214 1007 1215 1011
rect 1220 1007 1221 1011
rect 1214 1006 1221 1007
rect 465 1002 467 1006
rect 574 1003 580 1004
rect 574 1002 575 1003
rect 465 1000 575 1002
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 574 999 575 1000
rect 579 999 580 1003
rect 574 998 580 999
rect 1238 999 1244 1000
rect 110 994 116 995
rect 1238 995 1239 999
rect 1243 995 1244 999
rect 2082 999 2088 1000
rect 2082 998 2083 999
rect 1238 994 1244 995
rect 1278 996 1284 997
rect 198 992 204 993
rect 198 988 199 992
rect 203 988 204 992
rect 198 987 204 988
rect 238 992 244 993
rect 238 988 239 992
rect 243 988 244 992
rect 238 987 244 988
rect 286 992 292 993
rect 286 988 287 992
rect 291 988 292 992
rect 286 987 292 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 390 992 396 993
rect 390 988 391 992
rect 395 988 396 992
rect 390 987 396 988
rect 438 992 444 993
rect 438 988 439 992
rect 443 988 444 992
rect 438 987 444 988
rect 486 992 492 993
rect 486 988 487 992
rect 491 988 492 992
rect 486 987 492 988
rect 534 992 540 993
rect 534 988 535 992
rect 539 988 540 992
rect 534 987 540 988
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 678 992 684 993
rect 678 988 679 992
rect 683 988 684 992
rect 678 987 684 988
rect 726 992 732 993
rect 726 988 727 992
rect 731 988 732 992
rect 726 987 732 988
rect 782 992 788 993
rect 782 988 783 992
rect 787 988 788 992
rect 782 987 788 988
rect 838 992 844 993
rect 838 988 839 992
rect 843 988 844 992
rect 838 987 844 988
rect 894 992 900 993
rect 894 988 895 992
rect 899 988 900 992
rect 894 987 900 988
rect 958 992 964 993
rect 958 988 959 992
rect 963 988 964 992
rect 958 987 964 988
rect 1022 992 1028 993
rect 1022 988 1023 992
rect 1027 988 1028 992
rect 1022 987 1028 988
rect 1086 992 1092 993
rect 1086 988 1087 992
rect 1091 988 1092 992
rect 1086 987 1092 988
rect 1150 992 1156 993
rect 1150 988 1151 992
rect 1155 988 1156 992
rect 1150 987 1156 988
rect 1190 992 1196 993
rect 1190 988 1191 992
rect 1195 988 1196 992
rect 1278 992 1279 996
rect 1283 992 1284 996
rect 1928 996 2083 998
rect 1278 991 1284 992
rect 1495 991 1501 992
rect 1190 987 1196 988
rect 1495 987 1496 991
rect 1500 990 1501 991
rect 1527 991 1533 992
rect 1527 990 1528 991
rect 1500 988 1528 990
rect 1500 987 1501 988
rect 1495 986 1501 987
rect 1527 987 1528 988
rect 1532 987 1533 991
rect 1527 986 1533 987
rect 1614 991 1620 992
rect 1614 987 1615 991
rect 1619 990 1620 991
rect 1647 991 1653 992
rect 1647 990 1648 991
rect 1619 988 1648 990
rect 1619 987 1620 988
rect 1614 986 1620 987
rect 1647 987 1648 988
rect 1652 987 1653 991
rect 1647 986 1653 987
rect 1726 991 1732 992
rect 1726 987 1727 991
rect 1731 990 1732 991
rect 1759 991 1765 992
rect 1759 990 1760 991
rect 1731 988 1760 990
rect 1731 987 1732 988
rect 1726 986 1732 987
rect 1759 987 1760 988
rect 1764 987 1765 991
rect 1759 986 1765 987
rect 1855 991 1861 992
rect 1855 987 1856 991
rect 1860 990 1861 991
rect 1928 990 1930 996
rect 2082 995 2083 996
rect 2087 995 2088 999
rect 2290 999 2296 1000
rect 2290 998 2291 999
rect 2082 994 2088 995
rect 2124 996 2291 998
rect 1860 988 1930 990
rect 1934 991 1940 992
rect 1860 987 1861 988
rect 1855 986 1861 987
rect 1934 987 1935 991
rect 1939 990 1940 991
rect 1943 991 1949 992
rect 1943 990 1944 991
rect 1939 988 1944 990
rect 1939 987 1940 988
rect 1934 986 1940 987
rect 1943 987 1944 988
rect 1948 987 1949 991
rect 1943 986 1949 987
rect 1967 991 1973 992
rect 1967 987 1968 991
rect 1972 990 1973 991
rect 2023 991 2029 992
rect 2023 990 2024 991
rect 1972 988 2024 990
rect 1972 987 1973 988
rect 1967 986 1973 987
rect 2023 987 2024 988
rect 2028 987 2029 991
rect 2023 986 2029 987
rect 2095 991 2101 992
rect 2095 987 2096 991
rect 2100 990 2101 991
rect 2124 990 2126 996
rect 2290 995 2291 996
rect 2295 995 2296 999
rect 2290 994 2296 995
rect 2406 996 2412 997
rect 2406 992 2407 996
rect 2411 992 2412 996
rect 2100 988 2126 990
rect 2130 991 2136 992
rect 2100 987 2101 988
rect 2095 986 2101 987
rect 2130 987 2131 991
rect 2135 990 2136 991
rect 2167 991 2173 992
rect 2167 990 2168 991
rect 2135 988 2168 990
rect 2135 987 2136 988
rect 2130 986 2136 987
rect 2167 987 2168 988
rect 2172 987 2173 991
rect 2167 986 2173 987
rect 2198 991 2204 992
rect 2198 987 2199 991
rect 2203 990 2204 991
rect 2231 991 2237 992
rect 2231 990 2232 991
rect 2203 988 2232 990
rect 2203 987 2204 988
rect 2198 986 2204 987
rect 2231 987 2232 988
rect 2236 987 2237 991
rect 2231 986 2237 987
rect 2270 991 2276 992
rect 2270 987 2271 991
rect 2275 990 2276 991
rect 2303 991 2309 992
rect 2406 991 2412 992
rect 2303 990 2304 991
rect 2275 988 2304 990
rect 2275 987 2276 988
rect 2270 986 2276 987
rect 2303 987 2304 988
rect 2308 987 2309 991
rect 2303 986 2309 987
rect 1278 979 1284 980
rect 1278 975 1279 979
rect 1283 975 1284 979
rect 1278 974 1284 975
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 1502 972 1508 973
rect 294 968 300 969
rect 294 964 295 968
rect 299 964 300 968
rect 294 963 300 964
rect 342 968 348 969
rect 342 964 343 968
rect 347 964 348 968
rect 342 963 348 964
rect 398 968 404 969
rect 398 964 399 968
rect 403 964 404 968
rect 398 963 404 964
rect 470 968 476 969
rect 470 964 471 968
rect 475 964 476 968
rect 470 963 476 964
rect 550 968 556 969
rect 550 964 551 968
rect 555 964 556 968
rect 550 963 556 964
rect 638 968 644 969
rect 638 964 639 968
rect 643 964 644 968
rect 638 963 644 964
rect 726 968 732 969
rect 726 964 727 968
rect 731 964 732 968
rect 726 963 732 964
rect 806 968 812 969
rect 806 964 807 968
rect 811 964 812 968
rect 806 963 812 964
rect 886 968 892 969
rect 886 964 887 968
rect 891 964 892 968
rect 886 963 892 964
rect 958 968 964 969
rect 958 964 959 968
rect 963 964 964 968
rect 958 963 964 964
rect 1022 968 1028 969
rect 1022 964 1023 968
rect 1027 964 1028 968
rect 1022 963 1028 964
rect 1086 968 1092 969
rect 1086 964 1087 968
rect 1091 964 1092 968
rect 1086 963 1092 964
rect 1150 968 1156 969
rect 1150 964 1151 968
rect 1155 964 1156 968
rect 1150 963 1156 964
rect 1190 968 1196 969
rect 1190 964 1191 968
rect 1195 964 1196 968
rect 1502 968 1503 972
rect 1507 968 1508 972
rect 1502 967 1508 968
rect 1622 972 1628 973
rect 1622 968 1623 972
rect 1627 968 1628 972
rect 1622 967 1628 968
rect 1734 972 1740 973
rect 1734 968 1735 972
rect 1739 968 1740 972
rect 1734 967 1740 968
rect 1830 972 1836 973
rect 1830 968 1831 972
rect 1835 968 1836 972
rect 1830 967 1836 968
rect 1918 972 1924 973
rect 1918 968 1919 972
rect 1923 968 1924 972
rect 1918 967 1924 968
rect 1998 972 2004 973
rect 1998 968 1999 972
rect 2003 968 2004 972
rect 1998 967 2004 968
rect 2070 972 2076 973
rect 2070 968 2071 972
rect 2075 968 2076 972
rect 2070 967 2076 968
rect 2142 972 2148 973
rect 2142 968 2143 972
rect 2147 968 2148 972
rect 2142 967 2148 968
rect 2206 972 2212 973
rect 2206 968 2207 972
rect 2211 968 2212 972
rect 2206 967 2212 968
rect 2278 972 2284 973
rect 2278 968 2279 972
rect 2283 968 2284 972
rect 2278 967 2284 968
rect 1190 963 1196 964
rect 110 961 116 962
rect 110 957 111 961
rect 115 957 116 961
rect 110 956 116 957
rect 1238 961 1244 962
rect 1238 957 1239 961
rect 1243 957 1244 961
rect 1238 956 1244 957
rect 406 955 412 956
rect 406 954 407 955
rect 320 952 407 954
rect 320 948 322 952
rect 406 951 407 952
rect 411 951 412 955
rect 406 950 412 951
rect 1318 952 1324 953
rect 1318 948 1319 952
rect 1323 948 1324 952
rect 319 947 325 948
rect 110 944 116 945
rect 110 940 111 944
rect 115 940 116 944
rect 319 943 320 947
rect 324 943 325 947
rect 319 942 325 943
rect 327 947 333 948
rect 327 943 328 947
rect 332 946 333 947
rect 367 947 373 948
rect 367 946 368 947
rect 332 944 368 946
rect 332 943 333 944
rect 327 942 333 943
rect 367 943 368 944
rect 372 943 373 947
rect 367 942 373 943
rect 375 947 381 948
rect 375 943 376 947
rect 380 946 381 947
rect 423 947 429 948
rect 423 946 424 947
rect 380 944 424 946
rect 380 943 381 944
rect 375 942 381 943
rect 423 943 424 944
rect 428 943 429 947
rect 423 942 429 943
rect 431 947 437 948
rect 431 943 432 947
rect 436 946 437 947
rect 495 947 501 948
rect 495 946 496 947
rect 436 944 496 946
rect 436 943 437 944
rect 431 942 437 943
rect 495 943 496 944
rect 500 943 501 947
rect 495 942 501 943
rect 575 947 581 948
rect 575 943 576 947
rect 580 946 581 947
rect 654 947 660 948
rect 654 946 655 947
rect 580 944 655 946
rect 580 943 581 944
rect 575 942 581 943
rect 654 943 655 944
rect 659 943 660 947
rect 654 942 660 943
rect 663 947 669 948
rect 663 943 664 947
rect 668 946 669 947
rect 718 947 724 948
rect 718 946 719 947
rect 668 944 719 946
rect 668 943 669 944
rect 663 942 669 943
rect 718 943 719 944
rect 723 943 724 947
rect 718 942 724 943
rect 738 947 744 948
rect 738 943 739 947
rect 743 946 744 947
rect 751 947 757 948
rect 751 946 752 947
rect 743 944 752 946
rect 743 943 744 944
rect 738 942 744 943
rect 751 943 752 944
rect 756 943 757 947
rect 751 942 757 943
rect 831 947 837 948
rect 831 943 832 947
rect 836 943 837 947
rect 831 942 837 943
rect 839 947 845 948
rect 839 943 840 947
rect 844 946 845 947
rect 911 947 917 948
rect 911 946 912 947
rect 844 944 912 946
rect 844 943 845 944
rect 839 942 845 943
rect 911 943 912 944
rect 916 943 917 947
rect 911 942 917 943
rect 919 947 925 948
rect 919 943 920 947
rect 924 946 925 947
rect 983 947 989 948
rect 983 946 984 947
rect 924 944 984 946
rect 924 943 925 944
rect 919 942 925 943
rect 983 943 984 944
rect 988 943 989 947
rect 983 942 989 943
rect 991 947 997 948
rect 991 943 992 947
rect 996 946 997 947
rect 1047 947 1053 948
rect 1047 946 1048 947
rect 996 944 1048 946
rect 996 943 997 944
rect 991 942 997 943
rect 1047 943 1048 944
rect 1052 943 1053 947
rect 1047 942 1053 943
rect 1110 947 1117 948
rect 1110 943 1111 947
rect 1116 943 1117 947
rect 1110 942 1117 943
rect 1119 947 1125 948
rect 1119 943 1120 947
rect 1124 946 1125 947
rect 1175 947 1181 948
rect 1175 946 1176 947
rect 1124 944 1176 946
rect 1124 943 1125 944
rect 1119 942 1125 943
rect 1175 943 1176 944
rect 1180 943 1181 947
rect 1175 942 1181 943
rect 1198 947 1204 948
rect 1198 943 1199 947
rect 1203 946 1204 947
rect 1215 947 1221 948
rect 1318 947 1324 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1398 952 1404 953
rect 1398 948 1399 952
rect 1403 948 1404 952
rect 1398 947 1404 948
rect 1462 952 1468 953
rect 1462 948 1463 952
rect 1467 948 1468 952
rect 1462 947 1468 948
rect 1542 952 1548 953
rect 1542 948 1543 952
rect 1547 948 1548 952
rect 1542 947 1548 948
rect 1638 952 1644 953
rect 1638 948 1639 952
rect 1643 948 1644 952
rect 1638 947 1644 948
rect 1734 952 1740 953
rect 1734 948 1735 952
rect 1739 948 1740 952
rect 1734 947 1740 948
rect 1838 952 1844 953
rect 1838 948 1839 952
rect 1843 948 1844 952
rect 1838 947 1844 948
rect 1934 952 1940 953
rect 1934 948 1935 952
rect 1939 948 1940 952
rect 1934 947 1940 948
rect 2022 952 2028 953
rect 2022 948 2023 952
rect 2027 948 2028 952
rect 2022 947 2028 948
rect 2102 952 2108 953
rect 2102 948 2103 952
rect 2107 948 2108 952
rect 2102 947 2108 948
rect 2174 952 2180 953
rect 2174 948 2175 952
rect 2179 948 2180 952
rect 2174 947 2180 948
rect 2238 952 2244 953
rect 2238 948 2239 952
rect 2243 948 2244 952
rect 2238 947 2244 948
rect 2310 952 2316 953
rect 2310 948 2311 952
rect 2315 948 2316 952
rect 2310 947 2316 948
rect 2358 952 2364 953
rect 2358 948 2359 952
rect 2363 948 2364 952
rect 2358 947 2364 948
rect 1215 946 1216 947
rect 1203 944 1216 946
rect 1203 943 1204 944
rect 1198 942 1204 943
rect 1215 943 1216 944
rect 1220 943 1221 947
rect 1278 945 1284 946
rect 1215 942 1221 943
rect 1238 944 1244 945
rect 110 939 116 940
rect 832 938 834 942
rect 1238 940 1239 944
rect 1243 940 1244 944
rect 1278 941 1279 945
rect 1283 941 1284 945
rect 1278 940 1284 941
rect 2406 945 2412 946
rect 2406 941 2407 945
rect 2411 941 2412 945
rect 2406 940 2412 941
rect 1214 939 1220 940
rect 1238 939 1244 940
rect 1214 938 1215 939
rect 832 936 1215 938
rect 1214 935 1215 936
rect 1219 935 1220 939
rect 1214 934 1220 935
rect 1343 931 1352 932
rect 1278 928 1284 929
rect 1278 924 1279 928
rect 1283 924 1284 928
rect 1343 927 1344 931
rect 1351 927 1352 931
rect 1343 926 1352 927
rect 1366 931 1372 932
rect 1366 927 1367 931
rect 1371 930 1372 931
rect 1383 931 1389 932
rect 1383 930 1384 931
rect 1371 928 1384 930
rect 1371 927 1372 928
rect 1366 926 1372 927
rect 1383 927 1384 928
rect 1388 927 1389 931
rect 1383 926 1389 927
rect 1406 931 1412 932
rect 1406 927 1407 931
rect 1411 930 1412 931
rect 1423 931 1429 932
rect 1423 930 1424 931
rect 1411 928 1424 930
rect 1411 927 1412 928
rect 1406 926 1412 927
rect 1423 927 1424 928
rect 1428 927 1429 931
rect 1423 926 1429 927
rect 1487 931 1496 932
rect 1487 927 1488 931
rect 1495 927 1496 931
rect 1567 931 1573 932
rect 1567 930 1568 931
rect 1487 926 1496 927
rect 1500 928 1568 930
rect 1278 923 1284 924
rect 1426 923 1432 924
rect 294 921 300 922
rect 294 917 295 921
rect 299 917 300 921
rect 294 916 300 917
rect 342 921 348 922
rect 342 917 343 921
rect 347 917 348 921
rect 342 916 348 917
rect 398 921 404 922
rect 398 917 399 921
rect 403 917 404 921
rect 398 916 404 917
rect 470 921 476 922
rect 470 917 471 921
rect 475 917 476 921
rect 470 916 476 917
rect 550 921 556 922
rect 550 917 551 921
rect 555 917 556 921
rect 550 916 556 917
rect 638 921 644 922
rect 638 917 639 921
rect 643 917 644 921
rect 638 916 644 917
rect 726 921 732 922
rect 726 917 727 921
rect 731 917 732 921
rect 726 916 732 917
rect 806 921 812 922
rect 806 917 807 921
rect 811 917 812 921
rect 806 916 812 917
rect 886 921 892 922
rect 886 917 887 921
rect 891 917 892 921
rect 886 916 892 917
rect 958 921 964 922
rect 958 917 959 921
rect 963 917 964 921
rect 958 916 964 917
rect 1022 921 1028 922
rect 1022 917 1023 921
rect 1027 917 1028 921
rect 1022 916 1028 917
rect 1086 921 1092 922
rect 1086 917 1087 921
rect 1091 917 1092 921
rect 1086 916 1092 917
rect 1150 921 1156 922
rect 1150 917 1151 921
rect 1155 917 1156 921
rect 1150 916 1156 917
rect 1190 921 1196 922
rect 1190 917 1191 921
rect 1195 917 1196 921
rect 1426 919 1427 923
rect 1431 922 1432 923
rect 1500 922 1502 928
rect 1567 927 1568 928
rect 1572 927 1573 931
rect 1567 926 1573 927
rect 1575 931 1581 932
rect 1575 927 1576 931
rect 1580 930 1581 931
rect 1663 931 1669 932
rect 1663 930 1664 931
rect 1580 928 1664 930
rect 1580 927 1581 928
rect 1575 926 1581 927
rect 1663 927 1664 928
rect 1668 927 1669 931
rect 1663 926 1669 927
rect 1671 931 1677 932
rect 1671 927 1672 931
rect 1676 930 1677 931
rect 1759 931 1765 932
rect 1759 930 1760 931
rect 1676 928 1760 930
rect 1676 927 1677 928
rect 1671 926 1677 927
rect 1759 927 1760 928
rect 1764 927 1765 931
rect 1759 926 1765 927
rect 1767 931 1773 932
rect 1767 927 1768 931
rect 1772 930 1773 931
rect 1863 931 1869 932
rect 1863 930 1864 931
rect 1772 928 1864 930
rect 1772 927 1773 928
rect 1767 926 1773 927
rect 1863 927 1864 928
rect 1868 927 1869 931
rect 1863 926 1869 927
rect 1959 931 1965 932
rect 1959 927 1960 931
rect 1964 930 1965 931
rect 1986 931 1992 932
rect 1964 928 1982 930
rect 1964 927 1965 928
rect 1959 926 1965 927
rect 1431 920 1502 922
rect 1980 922 1982 928
rect 1986 927 1987 931
rect 1991 930 1992 931
rect 2047 931 2053 932
rect 2047 930 2048 931
rect 1991 928 2048 930
rect 1991 927 1992 928
rect 1986 926 1992 927
rect 2047 927 2048 928
rect 2052 927 2053 931
rect 2047 926 2053 927
rect 2055 931 2061 932
rect 2055 927 2056 931
rect 2060 930 2061 931
rect 2127 931 2133 932
rect 2127 930 2128 931
rect 2060 928 2128 930
rect 2060 927 2061 928
rect 2055 926 2061 927
rect 2127 927 2128 928
rect 2132 927 2133 931
rect 2127 926 2133 927
rect 2199 931 2205 932
rect 2199 927 2200 931
rect 2204 930 2205 931
rect 2254 931 2260 932
rect 2254 930 2255 931
rect 2204 928 2255 930
rect 2204 927 2205 928
rect 2199 926 2205 927
rect 2254 927 2255 928
rect 2259 927 2260 931
rect 2254 926 2260 927
rect 2263 931 2269 932
rect 2263 927 2264 931
rect 2268 930 2269 931
rect 2326 931 2332 932
rect 2326 930 2327 931
rect 2268 928 2327 930
rect 2268 927 2269 928
rect 2263 926 2269 927
rect 2326 927 2327 928
rect 2331 927 2332 931
rect 2326 926 2332 927
rect 2335 931 2341 932
rect 2335 927 2336 931
rect 2340 930 2341 931
rect 2374 931 2380 932
rect 2374 930 2375 931
rect 2340 928 2375 930
rect 2340 927 2341 928
rect 2335 926 2341 927
rect 2374 927 2375 928
rect 2379 927 2380 931
rect 2374 926 2380 927
rect 2382 931 2389 932
rect 2382 927 2383 931
rect 2388 927 2389 931
rect 2382 926 2389 927
rect 2406 928 2412 929
rect 2406 924 2407 928
rect 2411 924 2412 928
rect 2198 923 2204 924
rect 2406 923 2412 924
rect 2198 922 2199 923
rect 1980 920 2199 922
rect 1431 919 1432 920
rect 1426 918 1432 919
rect 2198 919 2199 920
rect 2203 919 2204 923
rect 2198 918 2204 919
rect 1190 916 1196 917
rect 319 915 325 916
rect 319 911 320 915
rect 324 914 325 915
rect 327 915 333 916
rect 327 914 328 915
rect 324 912 328 914
rect 324 911 325 912
rect 319 910 325 911
rect 327 911 328 912
rect 332 911 333 915
rect 327 910 333 911
rect 367 915 373 916
rect 367 911 368 915
rect 372 914 373 915
rect 375 915 381 916
rect 375 914 376 915
rect 372 912 376 914
rect 372 911 373 912
rect 367 910 373 911
rect 375 911 376 912
rect 380 911 381 915
rect 375 910 381 911
rect 423 915 429 916
rect 423 911 424 915
rect 428 914 429 915
rect 431 915 437 916
rect 431 914 432 915
rect 428 912 432 914
rect 428 911 429 912
rect 423 910 429 911
rect 431 911 432 912
rect 436 911 437 915
rect 431 910 437 911
rect 495 915 501 916
rect 495 911 496 915
rect 500 914 501 915
rect 558 915 564 916
rect 558 914 559 915
rect 500 912 559 914
rect 500 911 501 912
rect 495 910 501 911
rect 558 911 559 912
rect 563 911 564 915
rect 558 910 564 911
rect 574 915 581 916
rect 574 911 575 915
rect 580 911 581 915
rect 574 910 581 911
rect 654 915 660 916
rect 654 911 655 915
rect 659 914 660 915
rect 663 915 669 916
rect 663 914 664 915
rect 659 912 664 914
rect 659 911 660 912
rect 654 910 660 911
rect 663 911 664 912
rect 668 911 669 915
rect 663 910 669 911
rect 718 915 724 916
rect 718 911 719 915
rect 723 914 724 915
rect 751 915 757 916
rect 751 914 752 915
rect 723 912 752 914
rect 723 911 724 912
rect 718 910 724 911
rect 751 911 752 912
rect 756 911 757 915
rect 751 910 757 911
rect 831 915 837 916
rect 831 911 832 915
rect 836 914 837 915
rect 839 915 845 916
rect 839 914 840 915
rect 836 912 840 914
rect 836 911 837 912
rect 831 910 837 911
rect 839 911 840 912
rect 844 911 845 915
rect 839 910 845 911
rect 911 915 917 916
rect 911 911 912 915
rect 916 914 917 915
rect 919 915 925 916
rect 919 914 920 915
rect 916 912 920 914
rect 916 911 917 912
rect 911 910 917 911
rect 919 911 920 912
rect 924 911 925 915
rect 919 910 925 911
rect 983 915 989 916
rect 983 911 984 915
rect 988 914 989 915
rect 991 915 997 916
rect 991 914 992 915
rect 988 912 992 914
rect 988 911 989 912
rect 983 910 989 911
rect 991 911 992 912
rect 996 911 997 915
rect 991 910 997 911
rect 1047 915 1053 916
rect 1047 911 1048 915
rect 1052 914 1053 915
rect 1078 915 1084 916
rect 1078 914 1079 915
rect 1052 912 1079 914
rect 1052 911 1053 912
rect 1047 910 1053 911
rect 1078 911 1079 912
rect 1083 911 1084 915
rect 1078 910 1084 911
rect 1111 915 1117 916
rect 1111 911 1112 915
rect 1116 914 1117 915
rect 1119 915 1125 916
rect 1119 914 1120 915
rect 1116 912 1120 914
rect 1116 911 1117 912
rect 1111 910 1117 911
rect 1119 911 1120 912
rect 1124 911 1125 915
rect 1119 910 1125 911
rect 1175 915 1181 916
rect 1175 911 1176 915
rect 1180 914 1181 915
rect 1198 915 1204 916
rect 1198 914 1199 915
rect 1180 912 1199 914
rect 1180 911 1181 912
rect 1175 910 1181 911
rect 1198 911 1199 912
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1214 915 1221 916
rect 1214 911 1215 915
rect 1220 911 1221 915
rect 1214 910 1221 911
rect 1318 905 1324 906
rect 1318 901 1319 905
rect 1323 901 1324 905
rect 1318 900 1324 901
rect 1358 905 1364 906
rect 1358 901 1359 905
rect 1363 901 1364 905
rect 1358 900 1364 901
rect 1398 905 1404 906
rect 1398 901 1399 905
rect 1403 901 1404 905
rect 1398 900 1404 901
rect 1462 905 1468 906
rect 1462 901 1463 905
rect 1467 901 1468 905
rect 1462 900 1468 901
rect 1542 905 1548 906
rect 1542 901 1543 905
rect 1547 901 1548 905
rect 1542 900 1548 901
rect 1638 905 1644 906
rect 1638 901 1639 905
rect 1643 901 1644 905
rect 1638 900 1644 901
rect 1734 905 1740 906
rect 1734 901 1735 905
rect 1739 901 1740 905
rect 1734 900 1740 901
rect 1838 905 1844 906
rect 1838 901 1839 905
rect 1843 901 1844 905
rect 1838 900 1844 901
rect 1934 905 1940 906
rect 1934 901 1935 905
rect 1939 901 1940 905
rect 1934 900 1940 901
rect 2022 905 2028 906
rect 2022 901 2023 905
rect 2027 901 2028 905
rect 2022 900 2028 901
rect 2102 905 2108 906
rect 2102 901 2103 905
rect 2107 901 2108 905
rect 2102 900 2108 901
rect 2174 905 2180 906
rect 2174 901 2175 905
rect 2179 901 2180 905
rect 2174 900 2180 901
rect 2238 905 2244 906
rect 2238 901 2239 905
rect 2243 901 2244 905
rect 2238 900 2244 901
rect 2310 905 2316 906
rect 2310 901 2311 905
rect 2315 901 2316 905
rect 2310 900 2316 901
rect 2358 905 2364 906
rect 2358 901 2359 905
rect 2363 901 2364 905
rect 2358 900 2364 901
rect 1343 899 1349 900
rect 1343 895 1344 899
rect 1348 898 1349 899
rect 1366 899 1372 900
rect 1366 898 1367 899
rect 1348 896 1367 898
rect 1348 895 1349 896
rect 1343 894 1349 895
rect 1366 895 1367 896
rect 1371 895 1372 899
rect 1366 894 1372 895
rect 1383 899 1389 900
rect 1383 895 1384 899
rect 1388 898 1389 899
rect 1406 899 1412 900
rect 1406 898 1407 899
rect 1388 896 1407 898
rect 1388 895 1389 896
rect 1383 894 1389 895
rect 1406 895 1407 896
rect 1411 895 1412 899
rect 1406 894 1412 895
rect 1423 899 1432 900
rect 1423 895 1424 899
rect 1431 895 1432 899
rect 1423 894 1432 895
rect 1487 899 1493 900
rect 1487 895 1488 899
rect 1492 898 1493 899
rect 1495 899 1501 900
rect 1495 898 1496 899
rect 1492 896 1496 898
rect 1492 895 1493 896
rect 1487 894 1493 895
rect 1495 895 1496 896
rect 1500 895 1501 899
rect 1495 894 1501 895
rect 1567 899 1573 900
rect 1567 895 1568 899
rect 1572 898 1573 899
rect 1575 899 1581 900
rect 1575 898 1576 899
rect 1572 896 1576 898
rect 1572 895 1573 896
rect 1567 894 1573 895
rect 1575 895 1576 896
rect 1580 895 1581 899
rect 1575 894 1581 895
rect 1663 899 1669 900
rect 1663 895 1664 899
rect 1668 898 1669 899
rect 1671 899 1677 900
rect 1671 898 1672 899
rect 1668 896 1672 898
rect 1668 895 1669 896
rect 1663 894 1669 895
rect 1671 895 1672 896
rect 1676 895 1677 899
rect 1671 894 1677 895
rect 1759 899 1765 900
rect 1759 895 1760 899
rect 1764 898 1765 899
rect 1767 899 1773 900
rect 1767 898 1768 899
rect 1764 896 1768 898
rect 1764 895 1765 896
rect 1759 894 1765 895
rect 1767 895 1768 896
rect 1772 895 1773 899
rect 1767 894 1773 895
rect 1778 899 1784 900
rect 1778 895 1779 899
rect 1783 898 1784 899
rect 1863 899 1869 900
rect 1863 898 1864 899
rect 1783 896 1864 898
rect 1783 895 1784 896
rect 1778 894 1784 895
rect 1863 895 1864 896
rect 1868 895 1869 899
rect 1863 894 1869 895
rect 1959 899 1965 900
rect 1959 895 1960 899
rect 1964 898 1965 899
rect 1986 899 1992 900
rect 1986 898 1987 899
rect 1964 896 1987 898
rect 1964 895 1965 896
rect 1959 894 1965 895
rect 1986 895 1987 896
rect 1991 895 1992 899
rect 1986 894 1992 895
rect 2047 899 2053 900
rect 2047 895 2048 899
rect 2052 898 2053 899
rect 2055 899 2061 900
rect 2055 898 2056 899
rect 2052 896 2056 898
rect 2052 895 2053 896
rect 2047 894 2053 895
rect 2055 895 2056 896
rect 2060 895 2061 899
rect 2055 894 2061 895
rect 2127 899 2136 900
rect 2127 895 2128 899
rect 2135 895 2136 899
rect 2127 894 2136 895
rect 2198 899 2205 900
rect 2198 895 2199 899
rect 2204 895 2205 899
rect 2198 894 2205 895
rect 2254 899 2260 900
rect 2254 895 2255 899
rect 2259 898 2260 899
rect 2263 899 2269 900
rect 2263 898 2264 899
rect 2259 896 2264 898
rect 2259 895 2260 896
rect 2254 894 2260 895
rect 2263 895 2264 896
rect 2268 895 2269 899
rect 2263 894 2269 895
rect 2326 899 2332 900
rect 2326 895 2327 899
rect 2331 898 2332 899
rect 2335 899 2341 900
rect 2335 898 2336 899
rect 2331 896 2336 898
rect 2331 895 2332 896
rect 2326 894 2332 895
rect 2335 895 2336 896
rect 2340 895 2341 899
rect 2335 894 2341 895
rect 2374 899 2380 900
rect 2374 895 2375 899
rect 2379 898 2380 899
rect 2383 899 2389 900
rect 2383 898 2384 899
rect 2379 896 2384 898
rect 2379 895 2380 896
rect 2374 894 2380 895
rect 2383 895 2384 896
rect 2388 895 2389 899
rect 2383 894 2389 895
rect 279 887 285 888
rect 254 883 260 884
rect 254 879 255 883
rect 259 879 260 883
rect 279 883 280 887
rect 284 886 285 887
rect 295 887 301 888
rect 295 886 296 887
rect 284 884 296 886
rect 284 883 285 884
rect 279 882 285 883
rect 295 883 296 884
rect 300 883 301 887
rect 334 887 341 888
rect 295 882 301 883
rect 310 883 316 884
rect 254 878 260 879
rect 310 879 311 883
rect 315 879 316 883
rect 334 883 335 887
rect 340 883 341 887
rect 386 887 392 888
rect 334 882 341 883
rect 374 883 380 884
rect 310 878 316 879
rect 374 879 375 883
rect 379 879 380 883
rect 386 883 387 887
rect 391 886 392 887
rect 399 887 405 888
rect 399 886 400 887
rect 391 884 400 886
rect 391 883 392 884
rect 386 882 392 883
rect 399 883 400 884
rect 404 883 405 887
rect 466 887 472 888
rect 399 882 405 883
rect 454 883 460 884
rect 374 878 380 879
rect 454 879 455 883
rect 459 879 460 883
rect 466 883 467 887
rect 471 886 472 887
rect 479 887 485 888
rect 479 886 480 887
rect 471 884 480 886
rect 471 883 472 884
rect 466 882 472 883
rect 479 883 480 884
rect 484 883 485 887
rect 546 887 552 888
rect 479 882 485 883
rect 534 883 540 884
rect 454 878 460 879
rect 534 879 535 883
rect 539 879 540 883
rect 546 883 547 887
rect 551 886 552 887
rect 559 887 565 888
rect 559 886 560 887
rect 551 884 560 886
rect 551 883 552 884
rect 546 882 552 883
rect 559 883 560 884
rect 564 883 565 887
rect 647 887 653 888
rect 559 882 565 883
rect 622 883 628 884
rect 534 878 540 879
rect 622 879 623 883
rect 627 879 628 883
rect 647 883 648 887
rect 652 886 653 887
rect 702 887 708 888
rect 702 886 703 887
rect 652 884 703 886
rect 652 883 653 884
rect 647 882 653 883
rect 702 883 703 884
rect 707 883 708 887
rect 735 887 744 888
rect 702 882 708 883
rect 710 883 716 884
rect 622 878 628 879
rect 710 879 711 883
rect 715 879 716 883
rect 735 883 736 887
rect 743 883 744 887
rect 815 887 821 888
rect 735 882 744 883
rect 790 883 796 884
rect 710 878 716 879
rect 790 879 791 883
rect 795 879 796 883
rect 815 883 816 887
rect 820 886 821 887
rect 854 887 860 888
rect 854 886 855 887
rect 820 884 855 886
rect 820 883 821 884
rect 815 882 821 883
rect 854 883 855 884
rect 859 883 860 887
rect 887 887 893 888
rect 854 882 860 883
rect 862 883 868 884
rect 790 878 796 879
rect 862 879 863 883
rect 867 879 868 883
rect 887 883 888 887
rect 892 886 893 887
rect 918 887 924 888
rect 918 886 919 887
rect 892 884 919 886
rect 892 883 893 884
rect 887 882 893 883
rect 918 883 919 884
rect 923 883 924 887
rect 946 887 952 888
rect 918 882 924 883
rect 934 883 940 884
rect 862 878 868 879
rect 934 879 935 883
rect 939 879 940 883
rect 946 883 947 887
rect 951 886 952 887
rect 959 887 965 888
rect 959 886 960 887
rect 951 884 960 886
rect 951 883 952 884
rect 946 882 952 883
rect 959 883 960 884
rect 964 883 965 887
rect 1010 887 1016 888
rect 959 882 965 883
rect 998 883 1004 884
rect 934 878 940 879
rect 998 879 999 883
rect 1003 879 1004 883
rect 1010 883 1011 887
rect 1015 886 1016 887
rect 1023 887 1029 888
rect 1023 886 1024 887
rect 1015 884 1024 886
rect 1015 883 1016 884
rect 1010 882 1016 883
rect 1023 883 1024 884
rect 1028 883 1029 887
rect 1079 887 1085 888
rect 1023 882 1029 883
rect 1054 883 1060 884
rect 998 878 1004 879
rect 1054 879 1055 883
rect 1059 879 1060 883
rect 1079 883 1080 887
rect 1084 886 1085 887
rect 1110 887 1116 888
rect 1110 886 1111 887
rect 1084 884 1111 886
rect 1084 883 1085 884
rect 1079 882 1085 883
rect 1110 883 1111 884
rect 1115 883 1116 887
rect 1143 887 1149 888
rect 1110 882 1116 883
rect 1118 883 1124 884
rect 1054 878 1060 879
rect 1118 879 1119 883
rect 1123 879 1124 883
rect 1143 883 1144 887
rect 1148 886 1149 887
rect 1174 887 1180 888
rect 1174 886 1175 887
rect 1148 884 1175 886
rect 1148 883 1149 884
rect 1143 882 1149 883
rect 1174 883 1175 884
rect 1179 883 1180 887
rect 1194 887 1200 888
rect 1174 882 1180 883
rect 1182 883 1188 884
rect 1118 878 1124 879
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1194 883 1195 887
rect 1199 886 1200 887
rect 1207 887 1213 888
rect 1207 886 1208 887
rect 1199 884 1208 886
rect 1199 883 1200 884
rect 1194 882 1200 883
rect 1207 883 1208 884
rect 1212 883 1213 887
rect 1207 882 1213 883
rect 1182 878 1188 879
rect 1346 879 1352 880
rect 1346 875 1347 879
rect 1351 878 1352 879
rect 1351 876 1426 878
rect 1351 875 1352 876
rect 1346 874 1352 875
rect 1359 871 1368 872
rect 1334 867 1340 868
rect 386 863 392 864
rect 386 862 387 863
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 319 860 387 862
rect 319 858 321 860
rect 386 859 387 860
rect 391 859 392 863
rect 946 863 952 864
rect 946 862 947 863
rect 386 858 392 859
rect 849 860 947 862
rect 281 856 321 858
rect 110 855 116 856
rect 279 855 285 856
rect 279 851 280 855
rect 284 851 285 855
rect 335 855 341 856
rect 335 854 336 855
rect 319 852 336 854
rect 279 850 285 851
rect 295 851 301 852
rect 295 847 296 851
rect 300 850 301 851
rect 319 850 321 852
rect 335 851 336 852
rect 340 851 341 855
rect 335 850 341 851
rect 399 855 405 856
rect 399 851 400 855
rect 404 854 405 855
rect 466 855 472 856
rect 466 854 467 855
rect 404 852 467 854
rect 404 851 405 852
rect 399 850 405 851
rect 466 851 467 852
rect 471 851 472 855
rect 466 850 472 851
rect 479 855 485 856
rect 479 851 480 855
rect 484 854 485 855
rect 546 855 552 856
rect 546 854 547 855
rect 484 852 547 854
rect 484 851 485 852
rect 479 850 485 851
rect 546 851 547 852
rect 551 851 552 855
rect 546 850 552 851
rect 558 855 565 856
rect 558 851 559 855
rect 564 851 565 855
rect 558 850 565 851
rect 638 855 644 856
rect 638 851 639 855
rect 643 854 644 855
rect 647 855 653 856
rect 647 854 648 855
rect 643 852 648 854
rect 643 851 644 852
rect 638 850 644 851
rect 647 851 648 852
rect 652 851 653 855
rect 647 850 653 851
rect 702 855 708 856
rect 702 851 703 855
rect 707 854 708 855
rect 735 855 741 856
rect 735 854 736 855
rect 707 852 736 854
rect 707 851 708 852
rect 702 850 708 851
rect 735 851 736 852
rect 740 851 741 855
rect 735 850 741 851
rect 815 855 821 856
rect 815 851 816 855
rect 820 854 821 855
rect 849 854 851 860
rect 946 859 947 860
rect 951 859 952 863
rect 1194 863 1200 864
rect 1194 862 1195 863
rect 946 858 952 859
rect 1073 860 1195 862
rect 820 852 851 854
rect 854 855 860 856
rect 820 851 821 852
rect 815 850 821 851
rect 854 851 855 855
rect 859 854 860 855
rect 887 855 893 856
rect 887 854 888 855
rect 859 852 888 854
rect 859 851 860 852
rect 854 850 860 851
rect 887 851 888 852
rect 892 851 893 855
rect 887 850 893 851
rect 959 855 965 856
rect 959 851 960 855
rect 964 854 965 855
rect 1010 855 1016 856
rect 1010 854 1011 855
rect 964 852 1011 854
rect 964 851 965 852
rect 959 850 965 851
rect 1010 851 1011 852
rect 1015 851 1016 855
rect 1010 850 1016 851
rect 1023 855 1029 856
rect 1023 851 1024 855
rect 1028 854 1029 855
rect 1073 854 1075 860
rect 1194 859 1195 860
rect 1199 859 1200 863
rect 1334 863 1335 867
rect 1339 863 1340 867
rect 1359 867 1360 871
rect 1367 867 1368 871
rect 1399 871 1408 872
rect 1359 866 1368 867
rect 1374 867 1380 868
rect 1334 862 1340 863
rect 1374 863 1375 867
rect 1379 863 1380 867
rect 1399 867 1400 871
rect 1407 867 1408 871
rect 1424 870 1426 876
rect 1439 871 1445 872
rect 1439 870 1440 871
rect 1424 868 1440 870
rect 1399 866 1408 867
rect 1414 867 1420 868
rect 1374 862 1380 863
rect 1414 863 1415 867
rect 1419 863 1420 867
rect 1439 867 1440 868
rect 1444 867 1445 871
rect 1490 871 1501 872
rect 1439 866 1445 867
rect 1470 867 1476 868
rect 1414 862 1420 863
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 1490 867 1491 871
rect 1495 867 1496 871
rect 1500 867 1501 871
rect 1546 871 1552 872
rect 1490 866 1501 867
rect 1534 867 1540 868
rect 1470 862 1476 863
rect 1534 863 1535 867
rect 1539 863 1540 867
rect 1546 867 1547 871
rect 1551 870 1552 871
rect 1559 871 1565 872
rect 1559 870 1560 871
rect 1551 868 1560 870
rect 1551 867 1552 868
rect 1546 866 1552 867
rect 1559 867 1560 868
rect 1564 867 1565 871
rect 1631 871 1637 872
rect 1559 866 1565 867
rect 1606 867 1612 868
rect 1534 862 1540 863
rect 1606 863 1607 867
rect 1611 863 1612 867
rect 1631 867 1632 871
rect 1636 870 1637 871
rect 1646 871 1652 872
rect 1646 870 1647 871
rect 1636 868 1647 870
rect 1636 867 1637 868
rect 1631 866 1637 867
rect 1646 867 1647 868
rect 1651 867 1652 871
rect 1690 871 1696 872
rect 1646 866 1652 867
rect 1678 867 1684 868
rect 1606 862 1612 863
rect 1678 863 1679 867
rect 1683 863 1684 867
rect 1690 867 1691 871
rect 1695 870 1696 871
rect 1703 871 1709 872
rect 1703 870 1704 871
rect 1695 868 1704 870
rect 1695 867 1696 868
rect 1690 866 1696 867
rect 1703 867 1704 868
rect 1708 867 1709 871
rect 1762 871 1768 872
rect 1703 866 1709 867
rect 1750 867 1756 868
rect 1678 862 1684 863
rect 1750 863 1751 867
rect 1755 863 1756 867
rect 1762 867 1763 871
rect 1767 870 1768 871
rect 1775 871 1781 872
rect 1775 870 1776 871
rect 1767 868 1776 870
rect 1767 867 1768 868
rect 1762 866 1768 867
rect 1775 867 1776 868
rect 1780 867 1781 871
rect 1847 871 1853 872
rect 1775 866 1781 867
rect 1822 867 1828 868
rect 1750 862 1756 863
rect 1822 863 1823 867
rect 1827 863 1828 867
rect 1847 867 1848 871
rect 1852 870 1853 871
rect 1886 871 1892 872
rect 1886 870 1887 871
rect 1852 868 1887 870
rect 1852 867 1853 868
rect 1847 866 1853 867
rect 1886 867 1887 868
rect 1891 867 1892 871
rect 1919 871 1925 872
rect 1886 866 1892 867
rect 1894 867 1900 868
rect 1822 862 1828 863
rect 1894 863 1895 867
rect 1899 863 1900 867
rect 1919 867 1920 871
rect 1924 870 1925 871
rect 1950 871 1956 872
rect 1950 870 1951 871
rect 1924 868 1951 870
rect 1924 867 1925 868
rect 1919 866 1925 867
rect 1950 867 1951 868
rect 1955 867 1956 871
rect 1983 871 1989 872
rect 1950 866 1956 867
rect 1958 867 1964 868
rect 1894 862 1900 863
rect 1958 863 1959 867
rect 1963 863 1964 867
rect 1983 867 1984 871
rect 1988 870 1989 871
rect 2014 871 2020 872
rect 2014 870 2015 871
rect 1988 868 2015 870
rect 1988 867 1989 868
rect 1983 866 1989 867
rect 2014 867 2015 868
rect 2019 867 2020 871
rect 2047 871 2053 872
rect 2014 866 2020 867
rect 2022 867 2028 868
rect 1958 862 1964 863
rect 2022 863 2023 867
rect 2027 863 2028 867
rect 2047 867 2048 871
rect 2052 870 2053 871
rect 2078 871 2084 872
rect 2078 870 2079 871
rect 2052 868 2079 870
rect 2052 867 2053 868
rect 2047 866 2053 867
rect 2078 867 2079 868
rect 2083 867 2084 871
rect 2111 871 2117 872
rect 2078 866 2084 867
rect 2086 867 2092 868
rect 2022 862 2028 863
rect 2086 863 2087 867
rect 2091 863 2092 867
rect 2111 867 2112 871
rect 2116 870 2117 871
rect 2134 871 2140 872
rect 2134 870 2135 871
rect 2116 868 2135 870
rect 2116 867 2117 868
rect 2111 866 2117 867
rect 2134 867 2135 868
rect 2139 867 2140 871
rect 2167 871 2173 872
rect 2134 866 2140 867
rect 2142 867 2148 868
rect 2086 862 2092 863
rect 2142 863 2143 867
rect 2147 863 2148 867
rect 2167 867 2168 871
rect 2172 870 2173 871
rect 2183 871 2189 872
rect 2183 870 2184 871
rect 2172 868 2184 870
rect 2172 867 2173 868
rect 2167 866 2173 867
rect 2183 867 2184 868
rect 2188 867 2189 871
rect 2223 871 2229 872
rect 2183 866 2189 867
rect 2198 867 2204 868
rect 2142 862 2148 863
rect 2198 863 2199 867
rect 2203 863 2204 867
rect 2223 867 2224 871
rect 2228 870 2229 871
rect 2246 871 2252 872
rect 2246 870 2247 871
rect 2228 868 2247 870
rect 2228 867 2229 868
rect 2223 866 2229 867
rect 2246 867 2247 868
rect 2251 867 2252 871
rect 2279 871 2285 872
rect 2246 866 2252 867
rect 2254 867 2260 868
rect 2198 862 2204 863
rect 2254 863 2255 867
rect 2259 863 2260 867
rect 2279 867 2280 871
rect 2284 870 2285 871
rect 2310 871 2316 872
rect 2310 870 2311 871
rect 2284 868 2311 870
rect 2284 867 2285 868
rect 2279 866 2285 867
rect 2310 867 2311 868
rect 2315 867 2316 871
rect 2343 871 2352 872
rect 2310 866 2316 867
rect 2318 867 2324 868
rect 2254 862 2260 863
rect 2318 863 2319 867
rect 2323 863 2324 867
rect 2343 867 2344 871
rect 2351 867 2352 871
rect 2382 871 2389 872
rect 2343 866 2352 867
rect 2358 867 2364 868
rect 2318 862 2324 863
rect 2358 863 2359 867
rect 2363 863 2364 867
rect 2382 867 2383 871
rect 2388 867 2389 871
rect 2382 866 2389 867
rect 2358 862 2364 863
rect 1194 858 1200 859
rect 1238 860 1244 861
rect 1238 856 1239 860
rect 1243 856 1244 860
rect 1028 852 1075 854
rect 1078 855 1085 856
rect 1028 851 1029 852
rect 1023 850 1029 851
rect 1078 851 1079 855
rect 1084 851 1085 855
rect 1078 850 1085 851
rect 1110 855 1116 856
rect 1110 851 1111 855
rect 1115 854 1116 855
rect 1143 855 1149 856
rect 1143 854 1144 855
rect 1115 852 1144 854
rect 1115 851 1116 852
rect 1110 850 1116 851
rect 1143 851 1144 852
rect 1148 851 1149 855
rect 1143 850 1149 851
rect 1174 855 1180 856
rect 1174 851 1175 855
rect 1179 854 1180 855
rect 1207 855 1213 856
rect 1238 855 1244 856
rect 1207 854 1208 855
rect 1179 852 1208 854
rect 1179 851 1180 852
rect 1174 850 1180 851
rect 1207 851 1208 852
rect 1212 851 1213 855
rect 1207 850 1213 851
rect 300 848 321 850
rect 300 847 301 848
rect 295 846 301 847
rect 1886 847 1892 848
rect 1278 844 1284 845
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1278 840 1279 844
rect 1283 840 1284 844
rect 1886 843 1887 847
rect 1891 846 1892 847
rect 2346 847 2352 848
rect 1891 844 1922 846
rect 1891 843 1892 844
rect 1886 842 1892 843
rect 1920 842 1922 844
rect 2346 843 2347 847
rect 2351 846 2352 847
rect 2351 844 2387 846
rect 2351 843 2352 844
rect 2346 842 2352 843
rect 1919 841 1925 842
rect 1278 839 1284 840
rect 1350 839 1356 840
rect 1238 838 1244 839
rect 254 836 260 837
rect 254 832 255 836
rect 259 832 260 836
rect 254 831 260 832
rect 310 836 316 837
rect 310 832 311 836
rect 315 832 316 836
rect 310 831 316 832
rect 374 836 380 837
rect 374 832 375 836
rect 379 832 380 836
rect 374 831 380 832
rect 454 836 460 837
rect 454 832 455 836
rect 459 832 460 836
rect 454 831 460 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 790 836 796 837
rect 790 832 791 836
rect 795 832 796 836
rect 790 831 796 832
rect 862 836 868 837
rect 862 832 863 836
rect 867 832 868 836
rect 862 831 868 832
rect 934 836 940 837
rect 934 832 935 836
rect 939 832 940 836
rect 934 831 940 832
rect 998 836 1004 837
rect 998 832 999 836
rect 1003 832 1004 836
rect 998 831 1004 832
rect 1054 836 1060 837
rect 1054 832 1055 836
rect 1059 832 1060 836
rect 1054 831 1060 832
rect 1118 836 1124 837
rect 1118 832 1119 836
rect 1123 832 1124 836
rect 1118 831 1124 832
rect 1182 836 1188 837
rect 1182 832 1183 836
rect 1187 832 1188 836
rect 1350 835 1351 839
rect 1355 838 1356 839
rect 1359 839 1365 840
rect 1359 838 1360 839
rect 1355 836 1360 838
rect 1355 835 1356 836
rect 1350 834 1356 835
rect 1359 835 1360 836
rect 1364 835 1365 839
rect 1359 834 1365 835
rect 1370 839 1376 840
rect 1370 835 1371 839
rect 1375 838 1376 839
rect 1399 839 1405 840
rect 1399 838 1400 839
rect 1375 836 1400 838
rect 1375 835 1376 836
rect 1370 834 1376 835
rect 1399 835 1400 836
rect 1404 835 1405 839
rect 1399 834 1405 835
rect 1410 839 1416 840
rect 1410 835 1411 839
rect 1415 838 1416 839
rect 1439 839 1445 840
rect 1439 838 1440 839
rect 1415 836 1440 838
rect 1415 835 1416 836
rect 1410 834 1416 835
rect 1439 835 1440 836
rect 1444 835 1445 839
rect 1439 834 1445 835
rect 1495 839 1501 840
rect 1495 835 1496 839
rect 1500 838 1501 839
rect 1546 839 1552 840
rect 1546 838 1547 839
rect 1500 836 1547 838
rect 1500 835 1501 836
rect 1495 834 1501 835
rect 1546 835 1547 836
rect 1551 835 1552 839
rect 1546 834 1552 835
rect 1559 839 1565 840
rect 1559 835 1560 839
rect 1564 838 1565 839
rect 1574 839 1580 840
rect 1574 838 1575 839
rect 1564 836 1575 838
rect 1564 835 1565 836
rect 1559 834 1565 835
rect 1574 835 1575 836
rect 1579 835 1580 839
rect 1574 834 1580 835
rect 1631 839 1637 840
rect 1631 835 1632 839
rect 1636 838 1637 839
rect 1690 839 1696 840
rect 1690 838 1691 839
rect 1636 836 1691 838
rect 1636 835 1637 836
rect 1631 834 1637 835
rect 1690 835 1691 836
rect 1695 835 1696 839
rect 1690 834 1696 835
rect 1703 839 1709 840
rect 1703 835 1704 839
rect 1708 838 1709 839
rect 1762 839 1768 840
rect 1762 838 1763 839
rect 1708 836 1763 838
rect 1708 835 1709 836
rect 1703 834 1709 835
rect 1762 835 1763 836
rect 1767 835 1768 839
rect 1762 834 1768 835
rect 1775 839 1784 840
rect 1775 835 1776 839
rect 1783 835 1784 839
rect 1775 834 1784 835
rect 1847 839 1853 840
rect 1847 835 1848 839
rect 1852 838 1853 839
rect 1852 836 1914 838
rect 1919 837 1920 841
rect 1924 837 1925 841
rect 2385 840 2387 844
rect 2406 844 2412 845
rect 2406 840 2407 844
rect 2411 840 2412 844
rect 1919 836 1925 837
rect 1950 839 1956 840
rect 1852 835 1853 836
rect 1847 834 1853 835
rect 1182 831 1188 832
rect 1912 830 1914 836
rect 1950 835 1951 839
rect 1955 838 1956 839
rect 1983 839 1989 840
rect 1983 838 1984 839
rect 1955 836 1984 838
rect 1955 835 1956 836
rect 1950 834 1956 835
rect 1983 835 1984 836
rect 1988 835 1989 839
rect 1983 834 1989 835
rect 2014 839 2020 840
rect 2014 835 2015 839
rect 2019 838 2020 839
rect 2047 839 2053 840
rect 2047 838 2048 839
rect 2019 836 2048 838
rect 2019 835 2020 836
rect 2014 834 2020 835
rect 2047 835 2048 836
rect 2052 835 2053 839
rect 2047 834 2053 835
rect 2078 839 2084 840
rect 2078 835 2079 839
rect 2083 838 2084 839
rect 2111 839 2117 840
rect 2111 838 2112 839
rect 2083 836 2112 838
rect 2083 835 2084 836
rect 2078 834 2084 835
rect 2111 835 2112 836
rect 2116 835 2117 839
rect 2111 834 2117 835
rect 2134 839 2140 840
rect 2134 835 2135 839
rect 2139 838 2140 839
rect 2167 839 2173 840
rect 2167 838 2168 839
rect 2139 836 2168 838
rect 2139 835 2140 836
rect 2134 834 2140 835
rect 2167 835 2168 836
rect 2172 835 2173 839
rect 2167 834 2173 835
rect 2223 839 2229 840
rect 2223 835 2224 839
rect 2228 835 2229 839
rect 2223 834 2229 835
rect 2246 839 2252 840
rect 2246 835 2247 839
rect 2251 838 2252 839
rect 2279 839 2285 840
rect 2279 838 2280 839
rect 2251 836 2280 838
rect 2251 835 2252 836
rect 2246 834 2252 835
rect 2279 835 2280 836
rect 2284 835 2285 839
rect 2279 834 2285 835
rect 2310 839 2316 840
rect 2310 835 2311 839
rect 2315 838 2316 839
rect 2343 839 2349 840
rect 2343 838 2344 839
rect 2315 836 2344 838
rect 2315 835 2316 836
rect 2310 834 2316 835
rect 2343 835 2344 836
rect 2348 835 2349 839
rect 2343 834 2349 835
rect 2383 839 2389 840
rect 2406 839 2412 840
rect 2383 835 2384 839
rect 2388 835 2389 839
rect 2383 834 2389 835
rect 2046 831 2052 832
rect 2046 830 2047 831
rect 1912 828 2047 830
rect 1278 827 1284 828
rect 190 824 196 825
rect 190 820 191 824
rect 195 820 196 824
rect 190 819 196 820
rect 246 824 252 825
rect 246 820 247 824
rect 251 820 252 824
rect 246 819 252 820
rect 310 824 316 825
rect 310 820 311 824
rect 315 820 316 824
rect 310 819 316 820
rect 382 824 388 825
rect 382 820 383 824
rect 387 820 388 824
rect 382 819 388 820
rect 462 824 468 825
rect 462 820 463 824
rect 467 820 468 824
rect 462 819 468 820
rect 542 824 548 825
rect 542 820 543 824
rect 547 820 548 824
rect 542 819 548 820
rect 614 824 620 825
rect 614 820 615 824
rect 619 820 620 824
rect 614 819 620 820
rect 686 824 692 825
rect 686 820 687 824
rect 691 820 692 824
rect 686 819 692 820
rect 750 824 756 825
rect 750 820 751 824
rect 755 820 756 824
rect 750 819 756 820
rect 814 824 820 825
rect 814 820 815 824
rect 819 820 820 824
rect 814 819 820 820
rect 870 824 876 825
rect 870 820 871 824
rect 875 820 876 824
rect 870 819 876 820
rect 926 824 932 825
rect 926 820 927 824
rect 931 820 932 824
rect 926 819 932 820
rect 982 824 988 825
rect 982 820 983 824
rect 987 820 988 824
rect 982 819 988 820
rect 1046 824 1052 825
rect 1046 820 1047 824
rect 1051 820 1052 824
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 2046 827 2047 828
rect 2051 827 2052 831
rect 2225 830 2227 834
rect 2382 831 2388 832
rect 2382 830 2383 831
rect 2225 828 2383 830
rect 2046 826 2052 827
rect 2382 827 2383 828
rect 2387 827 2388 831
rect 2382 826 2388 827
rect 2406 827 2412 828
rect 1278 822 1284 823
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 1046 819 1052 820
rect 1334 820 1340 821
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 110 812 116 813
rect 1238 817 1244 818
rect 1238 813 1239 817
rect 1243 813 1244 817
rect 1334 816 1335 820
rect 1339 816 1340 820
rect 1334 815 1340 816
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1414 815 1420 816
rect 1470 820 1476 821
rect 1470 816 1471 820
rect 1475 816 1476 820
rect 1470 815 1476 816
rect 1534 820 1540 821
rect 1534 816 1535 820
rect 1539 816 1540 820
rect 1534 815 1540 816
rect 1606 820 1612 821
rect 1606 816 1607 820
rect 1611 816 1612 820
rect 1606 815 1612 816
rect 1678 820 1684 821
rect 1678 816 1679 820
rect 1683 816 1684 820
rect 1678 815 1684 816
rect 1750 820 1756 821
rect 1750 816 1751 820
rect 1755 816 1756 820
rect 1750 815 1756 816
rect 1822 820 1828 821
rect 1822 816 1823 820
rect 1827 816 1828 820
rect 1822 815 1828 816
rect 1894 820 1900 821
rect 1894 816 1895 820
rect 1899 816 1900 820
rect 1894 815 1900 816
rect 1958 820 1964 821
rect 1958 816 1959 820
rect 1963 816 1964 820
rect 1958 815 1964 816
rect 2022 820 2028 821
rect 2022 816 2023 820
rect 2027 816 2028 820
rect 2022 815 2028 816
rect 2086 820 2092 821
rect 2086 816 2087 820
rect 2091 816 2092 820
rect 2086 815 2092 816
rect 2142 820 2148 821
rect 2142 816 2143 820
rect 2147 816 2148 820
rect 2142 815 2148 816
rect 2198 820 2204 821
rect 2198 816 2199 820
rect 2203 816 2204 820
rect 2198 815 2204 816
rect 2254 820 2260 821
rect 2254 816 2255 820
rect 2259 816 2260 820
rect 2254 815 2260 816
rect 2318 820 2324 821
rect 2318 816 2319 820
rect 2323 816 2324 820
rect 2318 815 2324 816
rect 2358 820 2364 821
rect 2358 816 2359 820
rect 2363 816 2364 820
rect 2358 815 2364 816
rect 1238 812 1244 813
rect 1302 804 1308 805
rect 215 803 221 804
rect 110 800 116 801
rect 110 796 111 800
rect 115 796 116 800
rect 215 799 216 803
rect 220 802 221 803
rect 270 803 277 804
rect 220 800 266 802
rect 220 799 221 800
rect 215 798 221 799
rect 110 795 116 796
rect 264 794 266 800
rect 270 799 271 803
rect 276 799 277 803
rect 270 798 277 799
rect 334 803 341 804
rect 334 799 335 803
rect 340 799 341 803
rect 334 798 341 799
rect 346 803 352 804
rect 346 799 347 803
rect 351 802 352 803
rect 407 803 413 804
rect 407 802 408 803
rect 351 800 408 802
rect 351 799 352 800
rect 346 798 352 799
rect 407 799 408 800
rect 412 799 413 803
rect 407 798 413 799
rect 487 803 493 804
rect 487 799 488 803
rect 492 802 493 803
rect 518 803 524 804
rect 518 802 519 803
rect 492 800 519 802
rect 492 799 493 800
rect 487 798 493 799
rect 518 799 519 800
rect 523 799 524 803
rect 518 798 524 799
rect 526 803 532 804
rect 526 799 527 803
rect 531 802 532 803
rect 567 803 573 804
rect 567 802 568 803
rect 531 800 568 802
rect 531 799 532 800
rect 526 798 532 799
rect 567 799 568 800
rect 572 799 573 803
rect 567 798 573 799
rect 575 803 581 804
rect 575 799 576 803
rect 580 802 581 803
rect 639 803 645 804
rect 639 802 640 803
rect 580 800 640 802
rect 580 799 581 800
rect 575 798 581 799
rect 639 799 640 800
rect 644 799 645 803
rect 639 798 645 799
rect 711 803 717 804
rect 711 799 712 803
rect 716 799 717 803
rect 711 798 717 799
rect 719 803 725 804
rect 719 799 720 803
rect 724 802 725 803
rect 775 803 781 804
rect 775 802 776 803
rect 724 800 776 802
rect 724 799 725 800
rect 719 798 725 799
rect 775 799 776 800
rect 780 799 781 803
rect 775 798 781 799
rect 783 803 789 804
rect 783 799 784 803
rect 788 802 789 803
rect 839 803 845 804
rect 839 802 840 803
rect 788 800 840 802
rect 788 799 789 800
rect 783 798 789 799
rect 839 799 840 800
rect 844 799 845 803
rect 839 798 845 799
rect 895 803 901 804
rect 895 799 896 803
rect 900 802 901 803
rect 918 803 924 804
rect 900 800 914 802
rect 900 799 901 800
rect 895 798 901 799
rect 406 795 412 796
rect 406 794 407 795
rect 264 792 407 794
rect 406 791 407 792
rect 411 791 412 795
rect 712 794 714 798
rect 894 795 900 796
rect 894 794 895 795
rect 712 792 895 794
rect 406 790 412 791
rect 894 791 895 792
rect 899 791 900 795
rect 912 794 914 800
rect 918 799 919 803
rect 923 802 924 803
rect 951 803 957 804
rect 951 802 952 803
rect 923 800 952 802
rect 923 799 924 800
rect 918 798 924 799
rect 951 799 952 800
rect 956 799 957 803
rect 951 798 957 799
rect 959 803 965 804
rect 959 799 960 803
rect 964 802 965 803
rect 1007 803 1013 804
rect 1007 802 1008 803
rect 964 800 1008 802
rect 964 799 965 800
rect 959 798 965 799
rect 1007 799 1008 800
rect 1012 799 1013 803
rect 1007 798 1013 799
rect 1015 803 1021 804
rect 1015 799 1016 803
rect 1020 802 1021 803
rect 1071 803 1077 804
rect 1071 802 1072 803
rect 1020 800 1072 802
rect 1020 799 1021 800
rect 1015 798 1021 799
rect 1071 799 1072 800
rect 1076 799 1077 803
rect 1071 798 1077 799
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1302 800 1303 804
rect 1307 800 1308 804
rect 1302 799 1308 800
rect 1342 804 1348 805
rect 1342 800 1343 804
rect 1347 800 1348 804
rect 1342 799 1348 800
rect 1406 804 1412 805
rect 1406 800 1407 804
rect 1411 800 1412 804
rect 1406 799 1412 800
rect 1478 804 1484 805
rect 1478 800 1479 804
rect 1483 800 1484 804
rect 1478 799 1484 800
rect 1550 804 1556 805
rect 1550 800 1551 804
rect 1555 800 1556 804
rect 1550 799 1556 800
rect 1622 804 1628 805
rect 1622 800 1623 804
rect 1627 800 1628 804
rect 1622 799 1628 800
rect 1694 804 1700 805
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1758 804 1764 805
rect 1758 800 1759 804
rect 1763 800 1764 804
rect 1758 799 1764 800
rect 1822 804 1828 805
rect 1822 800 1823 804
rect 1827 800 1828 804
rect 1822 799 1828 800
rect 1886 804 1892 805
rect 1886 800 1887 804
rect 1891 800 1892 804
rect 1886 799 1892 800
rect 1950 804 1956 805
rect 1950 800 1951 804
rect 1955 800 1956 804
rect 1950 799 1956 800
rect 2022 804 2028 805
rect 2022 800 2023 804
rect 2027 800 2028 804
rect 2022 799 2028 800
rect 2102 804 2108 805
rect 2102 800 2103 804
rect 2107 800 2108 804
rect 2102 799 2108 800
rect 2190 804 2196 805
rect 2190 800 2191 804
rect 2195 800 2196 804
rect 2190 799 2196 800
rect 2278 804 2284 805
rect 2278 800 2279 804
rect 2283 800 2284 804
rect 2278 799 2284 800
rect 2358 804 2364 805
rect 2358 800 2359 804
rect 2363 800 2364 804
rect 2358 799 2364 800
rect 1070 795 1076 796
rect 1238 795 1244 796
rect 1278 797 1284 798
rect 1070 794 1071 795
rect 912 792 1071 794
rect 894 790 900 791
rect 1070 791 1071 792
rect 1075 791 1076 795
rect 1278 793 1279 797
rect 1283 793 1284 797
rect 1278 792 1284 793
rect 2406 797 2412 798
rect 2406 793 2407 797
rect 2411 793 2412 797
rect 2406 792 2412 793
rect 1070 790 1076 791
rect 1327 783 1333 784
rect 1278 780 1284 781
rect 190 777 196 778
rect 190 773 191 777
rect 195 773 196 777
rect 190 772 196 773
rect 246 777 252 778
rect 246 773 247 777
rect 251 773 252 777
rect 246 772 252 773
rect 310 777 316 778
rect 310 773 311 777
rect 315 773 316 777
rect 310 772 316 773
rect 382 777 388 778
rect 382 773 383 777
rect 387 773 388 777
rect 382 772 388 773
rect 462 777 468 778
rect 462 773 463 777
rect 467 773 468 777
rect 462 772 468 773
rect 542 777 548 778
rect 542 773 543 777
rect 547 773 548 777
rect 542 772 548 773
rect 614 777 620 778
rect 614 773 615 777
rect 619 773 620 777
rect 614 772 620 773
rect 686 777 692 778
rect 686 773 687 777
rect 691 773 692 777
rect 686 772 692 773
rect 750 777 756 778
rect 750 773 751 777
rect 755 773 756 777
rect 750 772 756 773
rect 814 777 820 778
rect 814 773 815 777
rect 819 773 820 777
rect 814 772 820 773
rect 870 777 876 778
rect 870 773 871 777
rect 875 773 876 777
rect 870 772 876 773
rect 926 777 932 778
rect 926 773 927 777
rect 931 773 932 777
rect 926 772 932 773
rect 982 777 988 778
rect 982 773 983 777
rect 987 773 988 777
rect 982 772 988 773
rect 1046 777 1052 778
rect 1046 773 1047 777
rect 1051 773 1052 777
rect 1278 776 1279 780
rect 1283 776 1284 780
rect 1327 779 1328 783
rect 1332 782 1333 783
rect 1358 783 1364 784
rect 1358 782 1359 783
rect 1332 780 1359 782
rect 1332 779 1333 780
rect 1327 778 1333 779
rect 1358 779 1359 780
rect 1363 779 1364 783
rect 1358 778 1364 779
rect 1367 783 1373 784
rect 1367 779 1368 783
rect 1372 782 1373 783
rect 1386 783 1392 784
rect 1386 782 1387 783
rect 1372 780 1387 782
rect 1372 779 1373 780
rect 1367 778 1373 779
rect 1386 779 1387 780
rect 1391 779 1392 783
rect 1386 778 1392 779
rect 1394 783 1400 784
rect 1394 779 1395 783
rect 1399 782 1400 783
rect 1431 783 1437 784
rect 1431 782 1432 783
rect 1399 780 1432 782
rect 1399 779 1400 780
rect 1394 778 1400 779
rect 1431 779 1432 780
rect 1436 779 1437 783
rect 1431 778 1437 779
rect 1490 783 1496 784
rect 1490 779 1491 783
rect 1495 782 1496 783
rect 1503 783 1509 784
rect 1503 782 1504 783
rect 1495 780 1504 782
rect 1495 779 1496 780
rect 1490 778 1496 779
rect 1503 779 1504 780
rect 1508 779 1509 783
rect 1503 778 1509 779
rect 1511 783 1517 784
rect 1511 779 1512 783
rect 1516 782 1517 783
rect 1575 783 1581 784
rect 1575 782 1576 783
rect 1516 780 1576 782
rect 1516 779 1517 780
rect 1511 778 1517 779
rect 1575 779 1576 780
rect 1580 779 1581 783
rect 1575 778 1581 779
rect 1646 783 1653 784
rect 1646 779 1647 783
rect 1652 779 1653 783
rect 1646 778 1653 779
rect 1655 783 1661 784
rect 1655 779 1656 783
rect 1660 782 1661 783
rect 1719 783 1725 784
rect 1719 782 1720 783
rect 1660 780 1720 782
rect 1660 779 1661 780
rect 1655 778 1661 779
rect 1719 779 1720 780
rect 1724 779 1725 783
rect 1719 778 1725 779
rect 1783 783 1789 784
rect 1783 779 1784 783
rect 1788 782 1789 783
rect 1798 783 1804 784
rect 1798 782 1799 783
rect 1788 780 1799 782
rect 1788 779 1789 780
rect 1783 778 1789 779
rect 1798 779 1799 780
rect 1803 779 1804 783
rect 1798 778 1804 779
rect 1807 783 1813 784
rect 1807 779 1808 783
rect 1812 782 1813 783
rect 1847 783 1853 784
rect 1847 782 1848 783
rect 1812 780 1848 782
rect 1812 779 1813 780
rect 1807 778 1813 779
rect 1847 779 1848 780
rect 1852 779 1853 783
rect 1847 778 1853 779
rect 1855 783 1861 784
rect 1855 779 1856 783
rect 1860 782 1861 783
rect 1911 783 1917 784
rect 1911 782 1912 783
rect 1860 780 1912 782
rect 1860 779 1861 780
rect 1855 778 1861 779
rect 1911 779 1912 780
rect 1916 779 1917 783
rect 1911 778 1917 779
rect 1919 783 1925 784
rect 1919 779 1920 783
rect 1924 782 1925 783
rect 1975 783 1981 784
rect 1975 782 1976 783
rect 1924 780 1976 782
rect 1924 779 1925 780
rect 1919 778 1925 779
rect 1975 779 1976 780
rect 1980 779 1981 783
rect 1975 778 1981 779
rect 1983 783 1989 784
rect 1983 779 1984 783
rect 1988 782 1989 783
rect 2047 783 2053 784
rect 2047 782 2048 783
rect 1988 780 2048 782
rect 1988 779 1989 780
rect 1983 778 1989 779
rect 2047 779 2048 780
rect 2052 779 2053 783
rect 2047 778 2053 779
rect 2127 783 2133 784
rect 2127 779 2128 783
rect 2132 782 2133 783
rect 2183 783 2189 784
rect 2132 780 2178 782
rect 2132 779 2133 780
rect 2127 778 2133 779
rect 1278 775 1284 776
rect 1046 772 1052 773
rect 2176 774 2178 780
rect 2183 779 2184 783
rect 2188 782 2189 783
rect 2215 783 2221 784
rect 2215 782 2216 783
rect 2188 780 2216 782
rect 2188 779 2189 780
rect 2183 778 2189 779
rect 2215 779 2216 780
rect 2220 779 2221 783
rect 2215 778 2221 779
rect 2223 783 2229 784
rect 2223 779 2224 783
rect 2228 782 2229 783
rect 2303 783 2309 784
rect 2303 782 2304 783
rect 2228 780 2304 782
rect 2228 779 2229 780
rect 2223 778 2229 779
rect 2303 779 2304 780
rect 2308 779 2309 783
rect 2303 778 2309 779
rect 2322 783 2328 784
rect 2322 779 2323 783
rect 2327 782 2328 783
rect 2383 783 2389 784
rect 2383 782 2384 783
rect 2327 780 2384 782
rect 2327 779 2328 780
rect 2322 778 2328 779
rect 2383 779 2384 780
rect 2388 779 2389 783
rect 2383 778 2389 779
rect 2406 780 2412 781
rect 2406 776 2407 780
rect 2411 776 2412 780
rect 2302 775 2308 776
rect 2406 775 2412 776
rect 2302 774 2303 775
rect 2176 772 2303 774
rect 215 771 221 772
rect 215 767 216 771
rect 220 770 221 771
rect 262 771 268 772
rect 262 770 263 771
rect 220 768 263 770
rect 220 767 221 768
rect 215 766 221 767
rect 262 767 263 768
rect 267 767 268 771
rect 262 766 268 767
rect 271 771 277 772
rect 271 767 272 771
rect 276 770 277 771
rect 302 771 308 772
rect 302 770 303 771
rect 276 768 303 770
rect 276 767 277 768
rect 271 766 277 767
rect 302 767 303 768
rect 307 767 308 771
rect 302 766 308 767
rect 335 771 341 772
rect 335 767 336 771
rect 340 770 341 771
rect 346 771 352 772
rect 346 770 347 771
rect 340 768 347 770
rect 340 767 341 768
rect 335 766 341 767
rect 346 767 347 768
rect 351 767 352 771
rect 346 766 352 767
rect 406 771 413 772
rect 406 767 407 771
rect 412 767 413 771
rect 406 766 413 767
rect 487 771 493 772
rect 487 767 488 771
rect 492 770 493 771
rect 526 771 532 772
rect 526 770 527 771
rect 492 768 527 770
rect 492 767 493 768
rect 487 766 493 767
rect 526 767 527 768
rect 531 767 532 771
rect 526 766 532 767
rect 567 771 573 772
rect 567 767 568 771
rect 572 770 573 771
rect 575 771 581 772
rect 575 770 576 771
rect 572 768 576 770
rect 572 767 573 768
rect 567 766 573 767
rect 575 767 576 768
rect 580 767 581 771
rect 575 766 581 767
rect 638 771 645 772
rect 638 767 639 771
rect 644 767 645 771
rect 638 766 645 767
rect 711 771 717 772
rect 711 767 712 771
rect 716 770 717 771
rect 719 771 725 772
rect 719 770 720 771
rect 716 768 720 770
rect 716 767 717 768
rect 711 766 717 767
rect 719 767 720 768
rect 724 767 725 771
rect 719 766 725 767
rect 775 771 781 772
rect 775 767 776 771
rect 780 770 781 771
rect 783 771 789 772
rect 783 770 784 771
rect 780 768 784 770
rect 780 767 781 768
rect 775 766 781 767
rect 783 767 784 768
rect 788 767 789 771
rect 783 766 789 767
rect 839 771 845 772
rect 839 767 840 771
rect 844 770 845 771
rect 886 771 892 772
rect 886 770 887 771
rect 844 768 887 770
rect 844 767 845 768
rect 839 766 845 767
rect 886 767 887 768
rect 891 767 892 771
rect 886 766 892 767
rect 894 771 901 772
rect 894 767 895 771
rect 900 767 901 771
rect 894 766 901 767
rect 951 771 957 772
rect 951 767 952 771
rect 956 770 957 771
rect 959 771 965 772
rect 959 770 960 771
rect 956 768 960 770
rect 956 767 957 768
rect 951 766 957 767
rect 959 767 960 768
rect 964 767 965 771
rect 959 766 965 767
rect 1007 771 1013 772
rect 1007 767 1008 771
rect 1012 770 1013 771
rect 1015 771 1021 772
rect 1015 770 1016 771
rect 1012 768 1016 770
rect 1012 767 1013 768
rect 1007 766 1013 767
rect 1015 767 1016 768
rect 1020 767 1021 771
rect 1015 766 1021 767
rect 1070 771 1077 772
rect 1070 767 1071 771
rect 1076 767 1077 771
rect 2302 771 2303 772
rect 2307 771 2308 775
rect 2302 770 2308 771
rect 1070 766 1077 767
rect 1302 757 1308 758
rect 1302 753 1303 757
rect 1307 753 1308 757
rect 1302 752 1308 753
rect 1342 757 1348 758
rect 1342 753 1343 757
rect 1347 753 1348 757
rect 1342 752 1348 753
rect 1406 757 1412 758
rect 1406 753 1407 757
rect 1411 753 1412 757
rect 1406 752 1412 753
rect 1478 757 1484 758
rect 1478 753 1479 757
rect 1483 753 1484 757
rect 1478 752 1484 753
rect 1550 757 1556 758
rect 1550 753 1551 757
rect 1555 753 1556 757
rect 1550 752 1556 753
rect 1622 757 1628 758
rect 1622 753 1623 757
rect 1627 753 1628 757
rect 1622 752 1628 753
rect 1694 757 1700 758
rect 1694 753 1695 757
rect 1699 753 1700 757
rect 1694 752 1700 753
rect 1758 757 1764 758
rect 1758 753 1759 757
rect 1763 753 1764 757
rect 1758 752 1764 753
rect 1822 757 1828 758
rect 1822 753 1823 757
rect 1827 753 1828 757
rect 1822 752 1828 753
rect 1886 757 1892 758
rect 1886 753 1887 757
rect 1891 753 1892 757
rect 1886 752 1892 753
rect 1950 757 1956 758
rect 1950 753 1951 757
rect 1955 753 1956 757
rect 1950 752 1956 753
rect 2022 757 2028 758
rect 2022 753 2023 757
rect 2027 753 2028 757
rect 2022 752 2028 753
rect 2102 757 2108 758
rect 2102 753 2103 757
rect 2107 753 2108 757
rect 2102 752 2108 753
rect 2190 757 2196 758
rect 2190 753 2191 757
rect 2195 753 2196 757
rect 2190 752 2196 753
rect 2278 757 2284 758
rect 2278 753 2279 757
rect 2283 753 2284 757
rect 2278 752 2284 753
rect 2358 757 2364 758
rect 2358 753 2359 757
rect 2363 753 2364 757
rect 2358 752 2364 753
rect 159 751 168 752
rect 134 747 140 748
rect 134 743 135 747
rect 139 743 140 747
rect 159 747 160 751
rect 167 747 168 751
rect 198 751 205 752
rect 159 746 168 747
rect 174 747 180 748
rect 134 742 140 743
rect 174 743 175 747
rect 179 743 180 747
rect 198 747 199 751
rect 204 747 205 751
rect 239 751 245 752
rect 198 746 205 747
rect 214 747 220 748
rect 174 742 180 743
rect 214 743 215 747
rect 219 743 220 747
rect 239 747 240 751
rect 244 747 245 751
rect 303 751 309 752
rect 239 746 245 747
rect 278 747 284 748
rect 214 742 220 743
rect 167 739 173 740
rect 167 735 168 739
rect 172 738 173 739
rect 241 738 243 746
rect 278 743 279 747
rect 283 743 284 747
rect 303 747 304 751
rect 308 750 309 751
rect 342 751 348 752
rect 342 750 343 751
rect 308 748 343 750
rect 308 747 309 748
rect 303 746 309 747
rect 342 747 343 748
rect 347 747 348 751
rect 362 751 368 752
rect 342 746 348 747
rect 350 747 356 748
rect 278 742 284 743
rect 350 743 351 747
rect 355 743 356 747
rect 362 747 363 751
rect 367 750 368 751
rect 375 751 381 752
rect 375 750 376 751
rect 367 748 376 750
rect 367 747 368 748
rect 362 746 368 747
rect 375 747 376 748
rect 380 747 381 751
rect 447 751 453 752
rect 375 746 381 747
rect 422 747 428 748
rect 350 742 356 743
rect 422 743 423 747
rect 427 743 428 747
rect 447 747 448 751
rect 452 750 453 751
rect 486 751 492 752
rect 486 750 487 751
rect 452 748 487 750
rect 452 747 453 748
rect 447 746 453 747
rect 486 747 487 748
rect 491 747 492 751
rect 518 751 525 752
rect 486 746 492 747
rect 494 747 500 748
rect 422 742 428 743
rect 494 743 495 747
rect 499 743 500 747
rect 518 747 519 751
rect 524 747 525 751
rect 583 751 589 752
rect 518 746 525 747
rect 558 747 564 748
rect 494 742 500 743
rect 558 743 559 747
rect 563 743 564 747
rect 583 747 584 751
rect 588 750 589 751
rect 614 751 620 752
rect 614 750 615 751
rect 588 748 615 750
rect 588 747 589 748
rect 583 746 589 747
rect 614 747 615 748
rect 619 747 620 751
rect 647 751 653 752
rect 614 746 620 747
rect 622 747 628 748
rect 558 742 564 743
rect 622 743 623 747
rect 627 743 628 747
rect 647 747 648 751
rect 652 750 653 751
rect 686 751 692 752
rect 686 750 687 751
rect 652 748 687 750
rect 652 747 653 748
rect 647 746 653 747
rect 686 747 687 748
rect 691 747 692 751
rect 719 751 725 752
rect 686 746 692 747
rect 694 747 700 748
rect 622 742 628 743
rect 694 743 695 747
rect 699 743 700 747
rect 719 747 720 751
rect 724 750 725 751
rect 758 751 764 752
rect 758 750 759 751
rect 724 748 759 750
rect 724 747 725 748
rect 719 746 725 747
rect 758 747 759 748
rect 763 747 764 751
rect 794 751 800 752
rect 758 746 764 747
rect 782 747 788 748
rect 694 742 700 743
rect 782 743 783 747
rect 787 743 788 747
rect 794 747 795 751
rect 799 750 800 751
rect 807 751 813 752
rect 807 750 808 751
rect 799 748 808 750
rect 799 747 800 748
rect 794 746 800 747
rect 807 747 808 748
rect 812 747 813 751
rect 903 751 909 752
rect 807 746 813 747
rect 878 747 884 748
rect 782 742 788 743
rect 878 743 879 747
rect 883 743 884 747
rect 903 747 904 751
rect 908 750 909 751
rect 974 751 980 752
rect 974 750 975 751
rect 908 748 975 750
rect 908 747 909 748
rect 903 746 909 747
rect 974 747 975 748
rect 979 747 980 751
rect 1007 751 1013 752
rect 974 746 980 747
rect 982 747 988 748
rect 878 742 884 743
rect 982 743 983 747
rect 987 743 988 747
rect 1007 747 1008 751
rect 1012 750 1013 751
rect 1086 751 1092 752
rect 1086 750 1087 751
rect 1012 748 1087 750
rect 1012 747 1013 748
rect 1007 746 1013 747
rect 1086 747 1087 748
rect 1091 747 1092 751
rect 1106 751 1112 752
rect 1086 746 1092 747
rect 1094 747 1100 748
rect 982 742 988 743
rect 1094 743 1095 747
rect 1099 743 1100 747
rect 1106 747 1107 751
rect 1111 750 1112 751
rect 1119 751 1125 752
rect 1119 750 1120 751
rect 1111 748 1120 750
rect 1111 747 1112 748
rect 1106 746 1112 747
rect 1119 747 1120 748
rect 1124 747 1125 751
rect 1215 751 1221 752
rect 1119 746 1125 747
rect 1190 747 1196 748
rect 1094 742 1100 743
rect 1190 743 1191 747
rect 1195 743 1196 747
rect 1215 747 1216 751
rect 1220 750 1221 751
rect 1318 751 1324 752
rect 1318 750 1319 751
rect 1220 748 1319 750
rect 1220 747 1221 748
rect 1215 746 1221 747
rect 1318 747 1319 748
rect 1323 747 1324 751
rect 1318 746 1324 747
rect 1327 751 1333 752
rect 1327 747 1328 751
rect 1332 750 1333 751
rect 1350 751 1356 752
rect 1350 750 1351 751
rect 1332 748 1351 750
rect 1332 747 1333 748
rect 1327 746 1333 747
rect 1350 747 1351 748
rect 1355 747 1356 751
rect 1350 746 1356 747
rect 1358 751 1364 752
rect 1358 747 1359 751
rect 1363 750 1364 751
rect 1367 751 1373 752
rect 1367 750 1368 751
rect 1363 748 1368 750
rect 1363 747 1364 748
rect 1358 746 1364 747
rect 1367 747 1368 748
rect 1372 747 1373 751
rect 1367 746 1373 747
rect 1386 751 1392 752
rect 1386 747 1387 751
rect 1391 750 1392 751
rect 1431 751 1437 752
rect 1431 750 1432 751
rect 1391 748 1432 750
rect 1391 747 1392 748
rect 1386 746 1392 747
rect 1431 747 1432 748
rect 1436 747 1437 751
rect 1431 746 1437 747
rect 1503 751 1509 752
rect 1503 747 1504 751
rect 1508 750 1509 751
rect 1511 751 1517 752
rect 1511 750 1512 751
rect 1508 748 1512 750
rect 1508 747 1509 748
rect 1503 746 1509 747
rect 1511 747 1512 748
rect 1516 747 1517 751
rect 1511 746 1517 747
rect 1574 751 1581 752
rect 1574 747 1575 751
rect 1580 747 1581 751
rect 1574 746 1581 747
rect 1647 751 1653 752
rect 1647 747 1648 751
rect 1652 750 1653 751
rect 1655 751 1661 752
rect 1655 750 1656 751
rect 1652 748 1656 750
rect 1652 747 1653 748
rect 1647 746 1653 747
rect 1655 747 1656 748
rect 1660 747 1661 751
rect 1655 746 1661 747
rect 1718 751 1725 752
rect 1718 747 1719 751
rect 1724 747 1725 751
rect 1718 746 1725 747
rect 1783 751 1789 752
rect 1783 747 1784 751
rect 1788 750 1789 751
rect 1807 751 1813 752
rect 1807 750 1808 751
rect 1788 748 1808 750
rect 1788 747 1789 748
rect 1783 746 1789 747
rect 1807 747 1808 748
rect 1812 747 1813 751
rect 1807 746 1813 747
rect 1847 751 1853 752
rect 1847 747 1848 751
rect 1852 750 1853 751
rect 1855 751 1861 752
rect 1855 750 1856 751
rect 1852 748 1856 750
rect 1852 747 1853 748
rect 1847 746 1853 747
rect 1855 747 1856 748
rect 1860 747 1861 751
rect 1855 746 1861 747
rect 1911 751 1917 752
rect 1911 747 1912 751
rect 1916 750 1917 751
rect 1919 751 1925 752
rect 1919 750 1920 751
rect 1916 748 1920 750
rect 1916 747 1917 748
rect 1911 746 1917 747
rect 1919 747 1920 748
rect 1924 747 1925 751
rect 1919 746 1925 747
rect 1975 751 1981 752
rect 1975 747 1976 751
rect 1980 750 1981 751
rect 1983 751 1989 752
rect 1983 750 1984 751
rect 1980 748 1984 750
rect 1980 747 1981 748
rect 1975 746 1981 747
rect 1983 747 1984 748
rect 1988 747 1989 751
rect 1983 746 1989 747
rect 2046 751 2053 752
rect 2046 747 2047 751
rect 2052 747 2053 751
rect 2046 746 2053 747
rect 2127 751 2133 752
rect 2127 747 2128 751
rect 2132 750 2133 751
rect 2142 751 2148 752
rect 2142 750 2143 751
rect 2132 748 2143 750
rect 2132 747 2133 748
rect 2127 746 2133 747
rect 2142 747 2143 748
rect 2147 747 2148 751
rect 2142 746 2148 747
rect 2215 751 2221 752
rect 2215 747 2216 751
rect 2220 750 2221 751
rect 2223 751 2229 752
rect 2223 750 2224 751
rect 2220 748 2224 750
rect 2220 747 2221 748
rect 2215 746 2221 747
rect 2223 747 2224 748
rect 2228 747 2229 751
rect 2223 746 2229 747
rect 2302 751 2309 752
rect 2302 747 2303 751
rect 2308 747 2309 751
rect 2302 746 2309 747
rect 2382 751 2389 752
rect 2382 747 2383 751
rect 2388 747 2389 751
rect 2382 746 2389 747
rect 1190 742 1196 743
rect 172 736 243 738
rect 172 735 173 736
rect 167 734 173 735
rect 1327 731 1333 732
rect 162 727 168 728
rect 110 724 116 725
rect 110 720 111 724
rect 115 720 116 724
rect 162 723 163 727
rect 167 726 168 727
rect 362 727 368 728
rect 362 726 363 727
rect 167 724 203 726
rect 167 723 168 724
rect 162 722 168 723
rect 201 720 203 724
rect 241 724 363 726
rect 241 720 243 724
rect 362 723 363 724
rect 367 723 368 727
rect 794 727 800 728
rect 794 726 795 727
rect 362 722 368 723
rect 585 724 795 726
rect 585 720 587 724
rect 794 723 795 724
rect 799 723 800 727
rect 1106 727 1112 728
rect 1106 726 1107 727
rect 794 722 800 723
rect 880 724 1107 726
rect 110 719 116 720
rect 159 719 165 720
rect 159 715 160 719
rect 164 718 165 719
rect 167 719 173 720
rect 167 718 168 719
rect 164 716 168 718
rect 164 715 165 716
rect 159 714 165 715
rect 167 715 168 716
rect 172 715 173 719
rect 167 714 173 715
rect 199 719 205 720
rect 199 715 200 719
rect 204 715 205 719
rect 199 714 205 715
rect 239 719 245 720
rect 239 715 240 719
rect 244 715 245 719
rect 239 714 245 715
rect 302 719 309 720
rect 302 715 303 719
rect 308 715 309 719
rect 302 714 309 715
rect 342 719 348 720
rect 342 715 343 719
rect 347 718 348 719
rect 375 719 381 720
rect 375 718 376 719
rect 347 716 376 718
rect 347 715 348 716
rect 342 714 348 715
rect 375 715 376 716
rect 380 715 381 719
rect 375 714 381 715
rect 438 719 444 720
rect 438 715 439 719
rect 443 718 444 719
rect 447 719 453 720
rect 447 718 448 719
rect 443 716 448 718
rect 443 715 444 716
rect 438 714 444 715
rect 447 715 448 716
rect 452 715 453 719
rect 447 714 453 715
rect 486 719 492 720
rect 486 715 487 719
rect 491 718 492 719
rect 519 719 525 720
rect 519 718 520 719
rect 491 716 520 718
rect 491 715 492 716
rect 486 714 492 715
rect 519 715 520 716
rect 524 715 525 719
rect 519 714 525 715
rect 583 719 589 720
rect 583 715 584 719
rect 588 715 589 719
rect 583 714 589 715
rect 614 719 620 720
rect 614 715 615 719
rect 619 718 620 719
rect 647 719 653 720
rect 647 718 648 719
rect 619 716 648 718
rect 619 715 620 716
rect 614 714 620 715
rect 647 715 648 716
rect 652 715 653 719
rect 647 714 653 715
rect 686 719 692 720
rect 686 715 687 719
rect 691 718 692 719
rect 719 719 725 720
rect 719 718 720 719
rect 691 716 720 718
rect 691 715 692 716
rect 686 714 692 715
rect 719 715 720 716
rect 724 715 725 719
rect 719 714 725 715
rect 807 719 813 720
rect 807 715 808 719
rect 812 718 813 719
rect 880 718 882 724
rect 1106 723 1107 724
rect 1111 723 1112 727
rect 1302 727 1308 728
rect 1106 722 1112 723
rect 1238 724 1244 725
rect 1238 720 1239 724
rect 1243 720 1244 724
rect 1302 723 1303 727
rect 1307 723 1308 727
rect 1327 727 1328 731
rect 1332 730 1333 731
rect 1358 731 1364 732
rect 1358 730 1359 731
rect 1332 728 1359 730
rect 1332 727 1333 728
rect 1327 726 1333 727
rect 1358 727 1359 728
rect 1363 727 1364 731
rect 1391 731 1400 732
rect 1358 726 1364 727
rect 1366 727 1372 728
rect 1302 722 1308 723
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 1391 727 1392 731
rect 1399 727 1400 731
rect 1479 731 1485 732
rect 1391 726 1400 727
rect 1454 727 1460 728
rect 1366 722 1372 723
rect 1454 723 1455 727
rect 1459 723 1460 727
rect 1479 727 1480 731
rect 1484 730 1485 731
rect 1490 731 1496 732
rect 1490 730 1491 731
rect 1484 728 1491 730
rect 1484 727 1485 728
rect 1479 726 1485 727
rect 1490 727 1491 728
rect 1495 727 1496 731
rect 1546 731 1552 732
rect 1490 726 1496 727
rect 1534 727 1540 728
rect 1454 722 1460 723
rect 1534 723 1535 727
rect 1539 723 1540 727
rect 1546 727 1547 731
rect 1551 730 1552 731
rect 1559 731 1565 732
rect 1559 730 1560 731
rect 1551 728 1560 730
rect 1551 727 1552 728
rect 1546 726 1552 727
rect 1559 727 1560 728
rect 1564 727 1565 731
rect 1639 731 1645 732
rect 1559 726 1565 727
rect 1614 727 1620 728
rect 1534 722 1540 723
rect 1614 723 1615 727
rect 1619 723 1620 727
rect 1639 727 1640 731
rect 1644 730 1645 731
rect 1662 731 1668 732
rect 1662 730 1663 731
rect 1644 728 1663 730
rect 1644 727 1645 728
rect 1639 726 1645 727
rect 1662 727 1663 728
rect 1667 727 1668 731
rect 1706 731 1712 732
rect 1662 726 1668 727
rect 1694 727 1700 728
rect 1614 722 1620 723
rect 1694 723 1695 727
rect 1699 723 1700 727
rect 1706 727 1707 731
rect 1711 730 1712 731
rect 1719 731 1725 732
rect 1719 730 1720 731
rect 1711 728 1720 730
rect 1711 727 1712 728
rect 1706 726 1712 727
rect 1719 727 1720 728
rect 1724 727 1725 731
rect 1798 731 1805 732
rect 1719 726 1725 727
rect 1774 727 1780 728
rect 1694 722 1700 723
rect 1774 723 1775 727
rect 1779 723 1780 727
rect 1798 727 1799 731
rect 1804 727 1805 731
rect 1866 731 1872 732
rect 1798 726 1805 727
rect 1854 727 1860 728
rect 1774 722 1780 723
rect 1854 723 1855 727
rect 1859 723 1860 727
rect 1866 727 1867 731
rect 1871 730 1872 731
rect 1879 731 1885 732
rect 1879 730 1880 731
rect 1871 728 1880 730
rect 1871 727 1872 728
rect 1866 726 1872 727
rect 1879 727 1880 728
rect 1884 727 1885 731
rect 1954 731 1960 732
rect 1879 726 1885 727
rect 1942 727 1948 728
rect 1854 722 1860 723
rect 1942 723 1943 727
rect 1947 723 1948 727
rect 1954 727 1955 731
rect 1959 730 1960 731
rect 1967 731 1973 732
rect 1967 730 1968 731
rect 1959 728 1968 730
rect 1959 727 1960 728
rect 1954 726 1960 727
rect 1967 727 1968 728
rect 1972 727 1973 731
rect 2042 731 2048 732
rect 1967 726 1973 727
rect 2030 727 2036 728
rect 1942 722 1948 723
rect 2030 723 2031 727
rect 2035 723 2036 727
rect 2042 727 2043 731
rect 2047 730 2048 731
rect 2055 731 2061 732
rect 2055 730 2056 731
rect 2047 728 2056 730
rect 2047 727 2048 728
rect 2042 726 2048 727
rect 2055 727 2056 728
rect 2060 727 2061 731
rect 2143 731 2149 732
rect 2055 726 2061 727
rect 2118 727 2124 728
rect 2030 722 2036 723
rect 2118 723 2119 727
rect 2123 723 2124 727
rect 2143 727 2144 731
rect 2148 730 2149 731
rect 2198 731 2204 732
rect 2198 730 2199 731
rect 2148 728 2199 730
rect 2148 727 2149 728
rect 2143 726 2149 727
rect 2198 727 2199 728
rect 2203 727 2204 731
rect 2231 731 2237 732
rect 2198 726 2204 727
rect 2206 727 2212 728
rect 2118 722 2124 723
rect 2206 723 2207 727
rect 2211 723 2212 727
rect 2231 727 2232 731
rect 2236 730 2237 731
rect 2286 731 2292 732
rect 2286 730 2287 731
rect 2236 728 2287 730
rect 2236 727 2237 728
rect 2231 726 2237 727
rect 2286 727 2287 728
rect 2291 727 2292 731
rect 2319 731 2328 732
rect 2286 726 2292 727
rect 2294 727 2300 728
rect 2206 722 2212 723
rect 2294 723 2295 727
rect 2299 723 2300 727
rect 2319 727 2320 731
rect 2327 727 2328 731
rect 2370 731 2376 732
rect 2319 726 2328 727
rect 2358 727 2364 728
rect 2294 722 2300 723
rect 2358 723 2359 727
rect 2363 723 2364 727
rect 2370 727 2371 731
rect 2375 730 2376 731
rect 2383 731 2389 732
rect 2383 730 2384 731
rect 2375 728 2384 730
rect 2375 727 2376 728
rect 2370 726 2376 727
rect 2383 727 2384 728
rect 2388 727 2389 731
rect 2383 726 2389 727
rect 2358 722 2364 723
rect 812 716 882 718
rect 886 719 892 720
rect 812 715 813 716
rect 807 714 813 715
rect 886 715 887 719
rect 891 718 892 719
rect 903 719 909 720
rect 903 718 904 719
rect 891 716 904 718
rect 891 715 892 716
rect 886 714 892 715
rect 903 715 904 716
rect 908 715 909 719
rect 903 714 909 715
rect 974 719 980 720
rect 974 715 975 719
rect 979 718 980 719
rect 1007 719 1013 720
rect 1007 718 1008 719
rect 979 716 1008 718
rect 979 715 980 716
rect 974 714 980 715
rect 1007 715 1008 716
rect 1012 715 1013 719
rect 1007 714 1013 715
rect 1086 719 1092 720
rect 1086 715 1087 719
rect 1091 718 1092 719
rect 1119 719 1125 720
rect 1119 718 1120 719
rect 1091 716 1120 718
rect 1091 715 1092 716
rect 1086 714 1092 715
rect 1119 715 1120 716
rect 1124 715 1125 719
rect 1119 714 1125 715
rect 1174 719 1180 720
rect 1174 715 1175 719
rect 1179 718 1180 719
rect 1215 719 1221 720
rect 1238 719 1244 720
rect 1215 718 1216 719
rect 1179 716 1216 718
rect 1179 715 1180 716
rect 1174 714 1180 715
rect 1215 715 1216 716
rect 1220 715 1221 719
rect 1215 714 1221 715
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 1238 707 1244 708
rect 1238 703 1239 707
rect 1243 703 1244 707
rect 1238 702 1244 703
rect 1278 704 1284 705
rect 134 700 140 701
rect 134 696 135 700
rect 139 696 140 700
rect 134 695 140 696
rect 174 700 180 701
rect 174 696 175 700
rect 179 696 180 700
rect 174 695 180 696
rect 214 700 220 701
rect 214 696 215 700
rect 219 696 220 700
rect 214 695 220 696
rect 278 700 284 701
rect 278 696 279 700
rect 283 696 284 700
rect 278 695 284 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 422 700 428 701
rect 422 696 423 700
rect 427 696 428 700
rect 422 695 428 696
rect 494 700 500 701
rect 494 696 495 700
rect 499 696 500 700
rect 494 695 500 696
rect 558 700 564 701
rect 558 696 559 700
rect 563 696 564 700
rect 558 695 564 696
rect 622 700 628 701
rect 622 696 623 700
rect 627 696 628 700
rect 622 695 628 696
rect 694 700 700 701
rect 694 696 695 700
rect 699 696 700 700
rect 694 695 700 696
rect 782 700 788 701
rect 782 696 783 700
rect 787 696 788 700
rect 782 695 788 696
rect 878 700 884 701
rect 878 696 879 700
rect 883 696 884 700
rect 878 695 884 696
rect 982 700 988 701
rect 982 696 983 700
rect 987 696 988 700
rect 982 695 988 696
rect 1094 700 1100 701
rect 1094 696 1095 700
rect 1099 696 1100 700
rect 1094 695 1100 696
rect 1190 700 1196 701
rect 1190 696 1191 700
rect 1195 696 1196 700
rect 1278 700 1279 704
rect 1283 700 1284 704
rect 2406 704 2412 705
rect 2406 700 2407 704
rect 2411 700 2412 704
rect 1278 699 1284 700
rect 1318 699 1324 700
rect 1190 695 1196 696
rect 1318 695 1319 699
rect 1323 698 1324 699
rect 1327 699 1333 700
rect 1327 698 1328 699
rect 1323 696 1328 698
rect 1323 695 1324 696
rect 1318 694 1324 695
rect 1327 695 1328 696
rect 1332 695 1333 699
rect 1327 694 1333 695
rect 1358 699 1364 700
rect 1358 695 1359 699
rect 1363 698 1364 699
rect 1391 699 1397 700
rect 1391 698 1392 699
rect 1363 696 1392 698
rect 1363 695 1364 696
rect 1358 694 1364 695
rect 1391 695 1392 696
rect 1396 695 1397 699
rect 1391 694 1397 695
rect 1479 699 1485 700
rect 1479 695 1480 699
rect 1484 698 1485 699
rect 1546 699 1552 700
rect 1546 698 1547 699
rect 1484 696 1547 698
rect 1484 695 1485 696
rect 1479 694 1485 695
rect 1546 695 1547 696
rect 1551 695 1552 699
rect 1546 694 1552 695
rect 1559 699 1565 700
rect 1559 695 1560 699
rect 1564 698 1565 699
rect 1606 699 1612 700
rect 1606 698 1607 699
rect 1564 696 1607 698
rect 1564 695 1565 696
rect 1559 694 1565 695
rect 1606 695 1607 696
rect 1611 695 1612 699
rect 1606 694 1612 695
rect 1639 699 1645 700
rect 1639 695 1640 699
rect 1644 698 1645 699
rect 1706 699 1712 700
rect 1706 698 1707 699
rect 1644 696 1707 698
rect 1644 695 1645 696
rect 1639 694 1645 695
rect 1706 695 1707 696
rect 1711 695 1712 699
rect 1706 694 1712 695
rect 1718 699 1725 700
rect 1718 695 1719 699
rect 1724 695 1725 699
rect 1718 694 1725 695
rect 1799 699 1805 700
rect 1799 695 1800 699
rect 1804 698 1805 699
rect 1866 699 1872 700
rect 1866 698 1867 699
rect 1804 696 1867 698
rect 1804 695 1805 696
rect 1799 694 1805 695
rect 1866 695 1867 696
rect 1871 695 1872 699
rect 1866 694 1872 695
rect 1879 699 1885 700
rect 1879 695 1880 699
rect 1884 698 1885 699
rect 1954 699 1960 700
rect 1954 698 1955 699
rect 1884 696 1955 698
rect 1884 695 1885 696
rect 1879 694 1885 695
rect 1954 695 1955 696
rect 1959 695 1960 699
rect 1954 694 1960 695
rect 1967 699 1973 700
rect 1967 695 1968 699
rect 1972 698 1973 699
rect 2042 699 2048 700
rect 2042 698 2043 699
rect 1972 696 2043 698
rect 1972 695 1973 696
rect 1967 694 1973 695
rect 2042 695 2043 696
rect 2047 695 2048 699
rect 2042 694 2048 695
rect 2055 699 2061 700
rect 2055 695 2056 699
rect 2060 698 2061 699
rect 2134 699 2140 700
rect 2134 698 2135 699
rect 2060 696 2135 698
rect 2060 695 2061 696
rect 2055 694 2061 695
rect 2134 695 2135 696
rect 2139 695 2140 699
rect 2134 694 2140 695
rect 2142 699 2149 700
rect 2142 695 2143 699
rect 2148 695 2149 699
rect 2142 694 2149 695
rect 2198 699 2204 700
rect 2198 695 2199 699
rect 2203 698 2204 699
rect 2231 699 2237 700
rect 2231 698 2232 699
rect 2203 696 2232 698
rect 2203 695 2204 696
rect 2198 694 2204 695
rect 2231 695 2232 696
rect 2236 695 2237 699
rect 2231 694 2237 695
rect 2319 699 2325 700
rect 2319 695 2320 699
rect 2324 698 2325 699
rect 2370 699 2376 700
rect 2370 698 2371 699
rect 2324 696 2371 698
rect 2324 695 2325 696
rect 2319 694 2325 695
rect 2370 695 2371 696
rect 2375 695 2376 699
rect 2370 694 2376 695
rect 2382 699 2389 700
rect 2406 699 2412 700
rect 2382 695 2383 699
rect 2388 695 2389 699
rect 2382 694 2389 695
rect 1278 687 1284 688
rect 1278 683 1279 687
rect 1283 683 1284 687
rect 1278 682 1284 683
rect 2406 687 2412 688
rect 2406 683 2407 687
rect 2411 683 2412 687
rect 2406 682 2412 683
rect 134 680 140 681
rect 134 676 135 680
rect 139 676 140 680
rect 134 675 140 676
rect 174 680 180 681
rect 174 676 175 680
rect 179 676 180 680
rect 174 675 180 676
rect 230 680 236 681
rect 230 676 231 680
rect 235 676 236 680
rect 230 675 236 676
rect 286 680 292 681
rect 286 676 287 680
rect 291 676 292 680
rect 286 675 292 676
rect 342 680 348 681
rect 342 676 343 680
rect 347 676 348 680
rect 342 675 348 676
rect 398 680 404 681
rect 398 676 399 680
rect 403 676 404 680
rect 398 675 404 676
rect 454 680 460 681
rect 454 676 455 680
rect 459 676 460 680
rect 454 675 460 676
rect 502 680 508 681
rect 502 676 503 680
rect 507 676 508 680
rect 502 675 508 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 694 680 700 681
rect 694 676 695 680
rect 699 676 700 680
rect 694 675 700 676
rect 766 680 772 681
rect 766 676 767 680
rect 771 676 772 680
rect 766 675 772 676
rect 838 680 844 681
rect 838 676 839 680
rect 843 676 844 680
rect 838 675 844 676
rect 902 680 908 681
rect 902 676 903 680
rect 907 676 908 680
rect 902 675 908 676
rect 966 680 972 681
rect 966 676 967 680
rect 971 676 972 680
rect 966 675 972 676
rect 1022 680 1028 681
rect 1022 676 1023 680
rect 1027 676 1028 680
rect 1022 675 1028 676
rect 1086 680 1092 681
rect 1086 676 1087 680
rect 1091 676 1092 680
rect 1086 675 1092 676
rect 1150 680 1156 681
rect 1150 676 1151 680
rect 1155 676 1156 680
rect 1150 675 1156 676
rect 1190 680 1196 681
rect 1190 676 1191 680
rect 1195 676 1196 680
rect 1190 675 1196 676
rect 1302 680 1308 681
rect 1302 676 1303 680
rect 1307 676 1308 680
rect 1302 675 1308 676
rect 1366 680 1372 681
rect 1366 676 1367 680
rect 1371 676 1372 680
rect 1366 675 1372 676
rect 1454 680 1460 681
rect 1454 676 1455 680
rect 1459 676 1460 680
rect 1454 675 1460 676
rect 1534 680 1540 681
rect 1534 676 1535 680
rect 1539 676 1540 680
rect 1534 675 1540 676
rect 1614 680 1620 681
rect 1614 676 1615 680
rect 1619 676 1620 680
rect 1614 675 1620 676
rect 1694 680 1700 681
rect 1694 676 1695 680
rect 1699 676 1700 680
rect 1694 675 1700 676
rect 1774 680 1780 681
rect 1774 676 1775 680
rect 1779 676 1780 680
rect 1774 675 1780 676
rect 1854 680 1860 681
rect 1854 676 1855 680
rect 1859 676 1860 680
rect 1854 675 1860 676
rect 1942 680 1948 681
rect 1942 676 1943 680
rect 1947 676 1948 680
rect 1942 675 1948 676
rect 2030 680 2036 681
rect 2030 676 2031 680
rect 2035 676 2036 680
rect 2030 675 2036 676
rect 2118 680 2124 681
rect 2118 676 2119 680
rect 2123 676 2124 680
rect 2118 675 2124 676
rect 2206 680 2212 681
rect 2206 676 2207 680
rect 2211 676 2212 680
rect 2206 675 2212 676
rect 2294 680 2300 681
rect 2294 676 2295 680
rect 2299 676 2300 680
rect 2294 675 2300 676
rect 2358 680 2364 681
rect 2358 676 2359 680
rect 2363 676 2364 680
rect 2358 675 2364 676
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 1238 673 1244 674
rect 1238 669 1239 673
rect 1243 669 1244 673
rect 1238 668 1244 669
rect 1590 668 1596 669
rect 1590 664 1591 668
rect 1595 664 1596 668
rect 1590 663 1596 664
rect 1638 668 1644 669
rect 1638 664 1639 668
rect 1643 664 1644 668
rect 1638 663 1644 664
rect 1686 668 1692 669
rect 1686 664 1687 668
rect 1691 664 1692 668
rect 1686 663 1692 664
rect 1742 668 1748 669
rect 1742 664 1743 668
rect 1747 664 1748 668
rect 1742 663 1748 664
rect 1798 668 1804 669
rect 1798 664 1799 668
rect 1803 664 1804 668
rect 1798 663 1804 664
rect 1870 668 1876 669
rect 1870 664 1871 668
rect 1875 664 1876 668
rect 1870 663 1876 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2150 668 2156 669
rect 2150 664 2151 668
rect 2155 664 2156 668
rect 2150 663 2156 664
rect 2262 668 2268 669
rect 2262 664 2263 668
rect 2267 664 2268 668
rect 2262 663 2268 664
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 1278 661 1284 662
rect 159 659 165 660
rect 110 656 116 657
rect 110 652 111 656
rect 115 652 116 656
rect 159 655 160 659
rect 164 655 165 659
rect 159 654 165 655
rect 198 659 205 660
rect 198 655 199 659
rect 204 655 205 659
rect 198 654 205 655
rect 210 659 216 660
rect 210 655 211 659
rect 215 658 216 659
rect 255 659 261 660
rect 255 658 256 659
rect 215 656 256 658
rect 215 655 216 656
rect 210 654 216 655
rect 255 655 256 656
rect 260 655 261 659
rect 255 654 261 655
rect 263 659 269 660
rect 263 655 264 659
rect 268 658 269 659
rect 311 659 317 660
rect 311 658 312 659
rect 268 656 312 658
rect 268 655 269 656
rect 263 654 269 655
rect 311 655 312 656
rect 316 655 317 659
rect 311 654 317 655
rect 367 659 373 660
rect 367 655 368 659
rect 372 655 373 659
rect 367 654 373 655
rect 375 659 381 660
rect 375 655 376 659
rect 380 658 381 659
rect 423 659 429 660
rect 423 658 424 659
rect 380 656 424 658
rect 380 655 381 656
rect 375 654 381 655
rect 423 655 424 656
rect 428 655 429 659
rect 423 654 429 655
rect 479 659 485 660
rect 479 655 480 659
rect 484 658 485 659
rect 494 659 500 660
rect 494 658 495 659
rect 484 656 495 658
rect 484 655 485 656
rect 479 654 485 655
rect 494 655 495 656
rect 499 655 500 659
rect 494 654 500 655
rect 514 659 520 660
rect 514 655 515 659
rect 519 658 520 659
rect 527 659 533 660
rect 527 658 528 659
rect 519 656 528 658
rect 519 655 520 656
rect 514 654 520 655
rect 527 655 528 656
rect 532 655 533 659
rect 527 654 533 655
rect 583 659 589 660
rect 583 655 584 659
rect 588 658 589 659
rect 638 659 644 660
rect 588 656 634 658
rect 588 655 589 656
rect 583 654 589 655
rect 110 651 116 652
rect 161 650 163 654
rect 310 651 316 652
rect 310 650 311 651
rect 161 648 311 650
rect 310 647 311 648
rect 315 647 316 651
rect 368 650 370 654
rect 478 651 484 652
rect 478 650 479 651
rect 368 648 479 650
rect 310 646 316 647
rect 478 647 479 648
rect 483 647 484 651
rect 632 650 634 656
rect 638 655 639 659
rect 643 658 644 659
rect 647 659 653 660
rect 647 658 648 659
rect 643 656 648 658
rect 643 655 644 656
rect 638 654 644 655
rect 647 655 648 656
rect 652 655 653 659
rect 647 654 653 655
rect 719 659 725 660
rect 719 655 720 659
rect 724 658 725 659
rect 758 659 764 660
rect 724 656 754 658
rect 724 655 725 656
rect 719 654 725 655
rect 718 651 724 652
rect 718 650 719 651
rect 632 648 719 650
rect 478 646 484 647
rect 718 647 719 648
rect 723 647 724 651
rect 752 650 754 656
rect 758 655 759 659
rect 763 658 764 659
rect 791 659 797 660
rect 791 658 792 659
rect 763 656 792 658
rect 763 655 764 656
rect 758 654 764 655
rect 791 655 792 656
rect 796 655 797 659
rect 791 654 797 655
rect 799 659 805 660
rect 799 655 800 659
rect 804 658 805 659
rect 863 659 869 660
rect 863 658 864 659
rect 804 656 864 658
rect 804 655 805 656
rect 799 654 805 655
rect 863 655 864 656
rect 868 655 869 659
rect 863 654 869 655
rect 914 659 920 660
rect 914 655 915 659
rect 919 658 920 659
rect 927 659 933 660
rect 927 658 928 659
rect 919 656 928 658
rect 919 655 920 656
rect 914 654 920 655
rect 927 655 928 656
rect 932 655 933 659
rect 927 654 933 655
rect 935 659 941 660
rect 935 655 936 659
rect 940 658 941 659
rect 991 659 997 660
rect 991 658 992 659
rect 940 656 992 658
rect 940 655 941 656
rect 935 654 941 655
rect 991 655 992 656
rect 996 655 997 659
rect 991 654 997 655
rect 999 659 1005 660
rect 999 655 1000 659
rect 1004 658 1005 659
rect 1047 659 1053 660
rect 1047 658 1048 659
rect 1004 656 1048 658
rect 1004 655 1005 656
rect 999 654 1005 655
rect 1047 655 1048 656
rect 1052 655 1053 659
rect 1047 654 1053 655
rect 1111 659 1117 660
rect 1111 655 1112 659
rect 1116 655 1117 659
rect 1111 654 1117 655
rect 1119 659 1125 660
rect 1119 655 1120 659
rect 1124 658 1125 659
rect 1175 659 1181 660
rect 1175 658 1176 659
rect 1124 656 1176 658
rect 1124 655 1125 656
rect 1119 654 1125 655
rect 1175 655 1176 656
rect 1180 655 1181 659
rect 1175 654 1181 655
rect 1214 659 1221 660
rect 1214 655 1215 659
rect 1220 655 1221 659
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1214 654 1221 655
rect 1238 656 1244 657
rect 1278 656 1284 657
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 862 651 868 652
rect 862 650 863 651
rect 752 648 863 650
rect 718 646 724 647
rect 862 647 863 648
rect 867 647 868 651
rect 1112 650 1114 654
rect 1238 652 1239 656
rect 1243 652 1244 656
rect 1198 651 1204 652
rect 1238 651 1244 652
rect 1198 650 1199 651
rect 1112 648 1199 650
rect 862 646 868 647
rect 1198 647 1199 648
rect 1203 647 1204 651
rect 1198 646 1204 647
rect 1582 647 1588 648
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1582 643 1583 647
rect 1587 646 1588 647
rect 1615 647 1621 648
rect 1615 646 1616 647
rect 1587 644 1616 646
rect 1587 643 1588 644
rect 1582 642 1588 643
rect 1615 643 1616 644
rect 1620 643 1621 647
rect 1615 642 1621 643
rect 1662 647 1669 648
rect 1662 643 1663 647
rect 1668 643 1669 647
rect 1662 642 1669 643
rect 1671 647 1677 648
rect 1671 643 1672 647
rect 1676 646 1677 647
rect 1711 647 1717 648
rect 1711 646 1712 647
rect 1676 644 1712 646
rect 1676 643 1677 644
rect 1671 642 1677 643
rect 1711 643 1712 644
rect 1716 643 1717 647
rect 1711 642 1717 643
rect 1719 647 1725 648
rect 1719 643 1720 647
rect 1724 646 1725 647
rect 1767 647 1773 648
rect 1767 646 1768 647
rect 1724 644 1768 646
rect 1724 643 1725 644
rect 1719 642 1725 643
rect 1767 643 1768 644
rect 1772 643 1773 647
rect 1767 642 1773 643
rect 1775 647 1781 648
rect 1775 643 1776 647
rect 1780 646 1781 647
rect 1823 647 1829 648
rect 1823 646 1824 647
rect 1780 644 1824 646
rect 1780 643 1781 644
rect 1775 642 1781 643
rect 1823 643 1824 644
rect 1828 643 1829 647
rect 1823 642 1829 643
rect 1831 647 1837 648
rect 1831 643 1832 647
rect 1836 646 1837 647
rect 1895 647 1901 648
rect 1895 646 1896 647
rect 1836 644 1896 646
rect 1836 643 1837 644
rect 1831 642 1837 643
rect 1895 643 1896 644
rect 1900 643 1901 647
rect 1895 642 1901 643
rect 1974 647 1981 648
rect 1974 643 1975 647
rect 1980 643 1981 647
rect 1974 642 1981 643
rect 1983 647 1989 648
rect 1983 643 1984 647
rect 1988 646 1989 647
rect 2071 647 2077 648
rect 2071 646 2072 647
rect 1988 644 2072 646
rect 1988 643 1989 644
rect 1983 642 1989 643
rect 2071 643 2072 644
rect 2076 643 2077 647
rect 2071 642 2077 643
rect 2082 647 2088 648
rect 2082 643 2083 647
rect 2087 646 2088 647
rect 2175 647 2181 648
rect 2175 646 2176 647
rect 2087 644 2176 646
rect 2087 643 2088 644
rect 2082 642 2088 643
rect 2175 643 2176 644
rect 2180 643 2181 647
rect 2175 642 2181 643
rect 2286 647 2293 648
rect 2286 643 2287 647
rect 2292 643 2293 647
rect 2286 642 2293 643
rect 2383 647 2389 648
rect 2383 643 2384 647
rect 2388 646 2389 647
rect 2391 647 2397 648
rect 2391 646 2392 647
rect 2388 644 2392 646
rect 2388 643 2389 644
rect 2383 642 2389 643
rect 2391 643 2392 644
rect 2396 643 2397 647
rect 2391 642 2397 643
rect 2406 644 2412 645
rect 1278 639 1284 640
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 134 633 140 634
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 230 633 236 634
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 286 633 292 634
rect 286 629 287 633
rect 291 629 292 633
rect 286 628 292 629
rect 342 633 348 634
rect 342 629 343 633
rect 347 629 348 633
rect 342 628 348 629
rect 398 633 404 634
rect 398 629 399 633
rect 403 629 404 633
rect 398 628 404 629
rect 454 633 460 634
rect 454 629 455 633
rect 459 629 460 633
rect 454 628 460 629
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 558 633 564 634
rect 558 629 559 633
rect 563 629 564 633
rect 558 628 564 629
rect 622 633 628 634
rect 622 629 623 633
rect 627 629 628 633
rect 622 628 628 629
rect 694 633 700 634
rect 694 629 695 633
rect 699 629 700 633
rect 694 628 700 629
rect 766 633 772 634
rect 766 629 767 633
rect 771 629 772 633
rect 766 628 772 629
rect 838 633 844 634
rect 838 629 839 633
rect 843 629 844 633
rect 838 628 844 629
rect 902 633 908 634
rect 902 629 903 633
rect 907 629 908 633
rect 902 628 908 629
rect 966 633 972 634
rect 966 629 967 633
rect 971 629 972 633
rect 966 628 972 629
rect 1022 633 1028 634
rect 1022 629 1023 633
rect 1027 629 1028 633
rect 1022 628 1028 629
rect 1086 633 1092 634
rect 1086 629 1087 633
rect 1091 629 1092 633
rect 1086 628 1092 629
rect 1150 633 1156 634
rect 1150 629 1151 633
rect 1155 629 1156 633
rect 1150 628 1156 629
rect 1190 633 1196 634
rect 1190 629 1191 633
rect 1195 629 1196 633
rect 1190 628 1196 629
rect 158 627 165 628
rect 158 623 159 627
rect 164 623 165 627
rect 158 622 165 623
rect 199 627 205 628
rect 199 623 200 627
rect 204 626 205 627
rect 210 627 216 628
rect 210 626 211 627
rect 204 624 211 626
rect 204 623 205 624
rect 199 622 205 623
rect 210 623 211 624
rect 215 623 216 627
rect 210 622 216 623
rect 255 627 261 628
rect 255 623 256 627
rect 260 626 261 627
rect 263 627 269 628
rect 263 626 264 627
rect 260 624 264 626
rect 260 623 261 624
rect 255 622 261 623
rect 263 623 264 624
rect 268 623 269 627
rect 263 622 269 623
rect 310 627 317 628
rect 310 623 311 627
rect 316 623 317 627
rect 310 622 317 623
rect 367 627 373 628
rect 367 623 368 627
rect 372 626 373 627
rect 375 627 381 628
rect 375 626 376 627
rect 372 624 376 626
rect 372 623 373 624
rect 367 622 373 623
rect 375 623 376 624
rect 380 623 381 627
rect 375 622 381 623
rect 423 627 429 628
rect 423 623 424 627
rect 428 626 429 627
rect 438 627 444 628
rect 438 626 439 627
rect 428 624 439 626
rect 428 623 429 624
rect 423 622 429 623
rect 438 623 439 624
rect 443 623 444 627
rect 438 622 444 623
rect 478 627 485 628
rect 478 623 479 627
rect 484 623 485 627
rect 478 622 485 623
rect 494 627 500 628
rect 494 623 495 627
rect 499 626 500 627
rect 527 627 533 628
rect 527 626 528 627
rect 499 624 528 626
rect 499 623 500 624
rect 494 622 500 623
rect 527 623 528 624
rect 532 623 533 627
rect 527 622 533 623
rect 583 627 589 628
rect 583 623 584 627
rect 588 626 589 627
rect 638 627 644 628
rect 638 626 639 627
rect 588 624 639 626
rect 588 623 589 624
rect 583 622 589 623
rect 638 623 639 624
rect 643 623 644 627
rect 638 622 644 623
rect 647 627 653 628
rect 647 623 648 627
rect 652 626 653 627
rect 662 627 668 628
rect 662 626 663 627
rect 652 624 663 626
rect 652 623 653 624
rect 647 622 653 623
rect 662 623 663 624
rect 667 623 668 627
rect 662 622 668 623
rect 718 627 725 628
rect 718 623 719 627
rect 724 623 725 627
rect 718 622 725 623
rect 791 627 797 628
rect 791 623 792 627
rect 796 626 797 627
rect 799 627 805 628
rect 799 626 800 627
rect 796 624 800 626
rect 796 623 797 624
rect 791 622 797 623
rect 799 623 800 624
rect 804 623 805 627
rect 799 622 805 623
rect 862 627 869 628
rect 862 623 863 627
rect 868 623 869 627
rect 862 622 869 623
rect 927 627 933 628
rect 927 623 928 627
rect 932 626 933 627
rect 935 627 941 628
rect 935 626 936 627
rect 932 624 936 626
rect 932 623 933 624
rect 927 622 933 623
rect 935 623 936 624
rect 940 623 941 627
rect 935 622 941 623
rect 991 627 997 628
rect 991 623 992 627
rect 996 626 997 627
rect 999 627 1005 628
rect 999 626 1000 627
rect 996 624 1000 626
rect 996 623 997 624
rect 991 622 997 623
rect 999 623 1000 624
rect 1004 623 1005 627
rect 999 622 1005 623
rect 1047 627 1053 628
rect 1047 623 1048 627
rect 1052 626 1053 627
rect 1102 627 1108 628
rect 1102 626 1103 627
rect 1052 624 1103 626
rect 1052 623 1053 624
rect 1047 622 1053 623
rect 1102 623 1103 624
rect 1107 623 1108 627
rect 1102 622 1108 623
rect 1111 627 1117 628
rect 1111 623 1112 627
rect 1116 626 1117 627
rect 1119 627 1125 628
rect 1119 626 1120 627
rect 1116 624 1120 626
rect 1116 623 1117 624
rect 1111 622 1117 623
rect 1119 623 1120 624
rect 1124 623 1125 627
rect 1119 622 1125 623
rect 1174 627 1181 628
rect 1174 623 1175 627
rect 1180 623 1181 627
rect 1174 622 1181 623
rect 1198 627 1204 628
rect 1198 623 1199 627
rect 1203 626 1204 627
rect 1215 627 1221 628
rect 1215 626 1216 627
rect 1203 624 1216 626
rect 1203 623 1204 624
rect 1198 622 1204 623
rect 1215 623 1216 624
rect 1220 623 1221 627
rect 1215 622 1221 623
rect 1590 621 1596 622
rect 1590 617 1591 621
rect 1595 617 1596 621
rect 1590 616 1596 617
rect 1638 621 1644 622
rect 1638 617 1639 621
rect 1643 617 1644 621
rect 1638 616 1644 617
rect 1686 621 1692 622
rect 1686 617 1687 621
rect 1691 617 1692 621
rect 1686 616 1692 617
rect 1742 621 1748 622
rect 1742 617 1743 621
rect 1747 617 1748 621
rect 1742 616 1748 617
rect 1798 621 1804 622
rect 1798 617 1799 621
rect 1803 617 1804 621
rect 1798 616 1804 617
rect 1870 621 1876 622
rect 1870 617 1871 621
rect 1875 617 1876 621
rect 1870 616 1876 617
rect 1950 621 1956 622
rect 1950 617 1951 621
rect 1955 617 1956 621
rect 1950 616 1956 617
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2150 621 2156 622
rect 2150 617 2151 621
rect 2155 617 2156 621
rect 2150 616 2156 617
rect 2262 621 2268 622
rect 2262 617 2263 621
rect 2267 617 2268 621
rect 2262 616 2268 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 1606 615 1612 616
rect 1606 611 1607 615
rect 1611 614 1612 615
rect 1615 615 1621 616
rect 1615 614 1616 615
rect 1611 612 1616 614
rect 1611 611 1612 612
rect 1606 610 1612 611
rect 1615 611 1616 612
rect 1620 611 1621 615
rect 1615 610 1621 611
rect 1663 615 1669 616
rect 1663 611 1664 615
rect 1668 614 1669 615
rect 1671 615 1677 616
rect 1671 614 1672 615
rect 1668 612 1672 614
rect 1668 611 1669 612
rect 1663 610 1669 611
rect 1671 611 1672 612
rect 1676 611 1677 615
rect 1671 610 1677 611
rect 1711 615 1717 616
rect 1711 611 1712 615
rect 1716 614 1717 615
rect 1719 615 1725 616
rect 1719 614 1720 615
rect 1716 612 1720 614
rect 1716 611 1717 612
rect 1711 610 1717 611
rect 1719 611 1720 612
rect 1724 611 1725 615
rect 1719 610 1725 611
rect 1767 615 1773 616
rect 1767 611 1768 615
rect 1772 614 1773 615
rect 1775 615 1781 616
rect 1775 614 1776 615
rect 1772 612 1776 614
rect 1772 611 1773 612
rect 1767 610 1773 611
rect 1775 611 1776 612
rect 1780 611 1781 615
rect 1775 610 1781 611
rect 1823 615 1829 616
rect 1823 611 1824 615
rect 1828 614 1829 615
rect 1831 615 1837 616
rect 1831 614 1832 615
rect 1828 612 1832 614
rect 1828 611 1829 612
rect 1823 610 1829 611
rect 1831 611 1832 612
rect 1836 611 1837 615
rect 1831 610 1837 611
rect 1890 615 1901 616
rect 1890 611 1891 615
rect 1895 611 1896 615
rect 1900 611 1901 615
rect 1890 610 1901 611
rect 1975 615 1981 616
rect 1975 611 1976 615
rect 1980 614 1981 615
rect 1983 615 1989 616
rect 1983 614 1984 615
rect 1980 612 1984 614
rect 1980 611 1981 612
rect 1975 610 1981 611
rect 1983 611 1984 612
rect 1988 611 1989 615
rect 1983 610 1989 611
rect 2071 615 2077 616
rect 2071 611 2072 615
rect 2076 614 2077 615
rect 2082 615 2088 616
rect 2082 614 2083 615
rect 2076 612 2083 614
rect 2076 611 2077 612
rect 2071 610 2077 611
rect 2082 611 2083 612
rect 2087 611 2088 615
rect 2082 610 2088 611
rect 2134 615 2140 616
rect 2134 611 2135 615
rect 2139 614 2140 615
rect 2175 615 2181 616
rect 2175 614 2176 615
rect 2139 612 2176 614
rect 2139 611 2140 612
rect 2134 610 2140 611
rect 2175 611 2176 612
rect 2180 611 2181 615
rect 2175 610 2181 611
rect 2215 615 2221 616
rect 2215 611 2216 615
rect 2220 614 2221 615
rect 2287 615 2293 616
rect 2287 614 2288 615
rect 2220 612 2288 614
rect 2220 611 2221 612
rect 2215 610 2221 611
rect 2287 611 2288 612
rect 2292 611 2293 615
rect 2287 610 2293 611
rect 2382 615 2389 616
rect 2382 611 2383 615
rect 2388 611 2389 615
rect 2382 610 2389 611
rect 159 607 165 608
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 159 603 160 607
rect 164 606 165 607
rect 174 607 180 608
rect 174 606 175 607
rect 164 604 175 606
rect 164 603 165 604
rect 159 602 165 603
rect 174 603 175 604
rect 179 603 180 607
rect 207 607 213 608
rect 174 602 180 603
rect 182 603 188 604
rect 134 598 140 599
rect 182 599 183 603
rect 187 599 188 603
rect 207 603 208 607
rect 212 606 213 607
rect 246 607 252 608
rect 246 606 247 607
rect 212 604 247 606
rect 212 603 213 604
rect 207 602 213 603
rect 246 603 247 604
rect 251 603 252 607
rect 279 607 285 608
rect 246 602 252 603
rect 254 603 260 604
rect 182 598 188 599
rect 254 599 255 603
rect 259 599 260 603
rect 279 603 280 607
rect 284 606 285 607
rect 318 607 324 608
rect 318 606 319 607
rect 284 604 319 606
rect 284 603 285 604
rect 279 602 285 603
rect 318 603 319 604
rect 323 603 324 607
rect 338 607 344 608
rect 318 602 324 603
rect 326 603 332 604
rect 254 598 260 599
rect 326 599 327 603
rect 331 599 332 603
rect 338 603 339 607
rect 343 606 344 607
rect 351 607 357 608
rect 351 606 352 607
rect 343 604 352 606
rect 343 603 344 604
rect 338 602 344 603
rect 351 603 352 604
rect 356 603 357 607
rect 423 607 429 608
rect 351 602 357 603
rect 398 603 404 604
rect 326 598 332 599
rect 398 599 399 603
rect 403 599 404 603
rect 423 603 424 607
rect 428 606 429 607
rect 470 607 476 608
rect 470 606 471 607
rect 428 604 471 606
rect 428 603 429 604
rect 423 602 429 603
rect 470 603 471 604
rect 475 603 476 607
rect 503 607 509 608
rect 470 602 476 603
rect 478 603 484 604
rect 398 598 404 599
rect 478 599 479 603
rect 483 599 484 603
rect 503 603 504 607
rect 508 606 509 607
rect 514 607 520 608
rect 514 606 515 607
rect 508 604 515 606
rect 508 603 509 604
rect 503 602 509 603
rect 514 603 515 604
rect 519 603 520 607
rect 570 607 576 608
rect 514 602 520 603
rect 558 603 564 604
rect 478 598 484 599
rect 558 599 559 603
rect 563 599 564 603
rect 570 603 571 607
rect 575 606 576 607
rect 583 607 589 608
rect 583 606 584 607
rect 575 604 584 606
rect 575 603 576 604
rect 570 602 576 603
rect 583 603 584 604
rect 588 603 589 607
rect 663 607 669 608
rect 583 602 589 603
rect 638 603 644 604
rect 558 598 564 599
rect 638 599 639 603
rect 643 599 644 603
rect 663 603 664 607
rect 668 606 669 607
rect 710 607 716 608
rect 710 606 711 607
rect 668 604 711 606
rect 668 603 669 604
rect 663 602 669 603
rect 710 603 711 604
rect 715 603 716 607
rect 743 607 749 608
rect 710 602 716 603
rect 718 603 724 604
rect 638 598 644 599
rect 718 599 719 603
rect 723 599 724 603
rect 743 603 744 607
rect 748 606 749 607
rect 790 607 796 608
rect 790 606 791 607
rect 748 604 791 606
rect 748 603 749 604
rect 743 602 749 603
rect 790 603 791 604
rect 795 603 796 607
rect 810 607 816 608
rect 790 602 796 603
rect 798 603 804 604
rect 718 598 724 599
rect 798 599 799 603
rect 803 599 804 603
rect 810 603 811 607
rect 815 606 816 607
rect 823 607 829 608
rect 823 606 824 607
rect 815 604 824 606
rect 815 603 816 604
rect 810 602 816 603
rect 823 603 824 604
rect 828 603 829 607
rect 903 607 909 608
rect 823 602 829 603
rect 878 603 884 604
rect 798 598 804 599
rect 878 599 879 603
rect 883 599 884 603
rect 903 603 904 607
rect 908 606 909 607
rect 914 607 920 608
rect 914 606 915 607
rect 908 604 915 606
rect 908 603 909 604
rect 903 602 909 603
rect 914 603 915 604
rect 919 603 920 607
rect 962 607 968 608
rect 914 602 920 603
rect 950 603 956 604
rect 878 598 884 599
rect 950 599 951 603
rect 955 599 956 603
rect 962 603 963 607
rect 967 606 968 607
rect 975 607 981 608
rect 975 606 976 607
rect 967 604 976 606
rect 967 603 968 604
rect 962 602 968 603
rect 975 603 976 604
rect 980 603 981 607
rect 1026 607 1032 608
rect 975 602 981 603
rect 1014 603 1020 604
rect 950 598 956 599
rect 1014 599 1015 603
rect 1019 599 1020 603
rect 1026 603 1027 607
rect 1031 606 1032 607
rect 1039 607 1045 608
rect 1039 606 1040 607
rect 1031 604 1040 606
rect 1031 603 1032 604
rect 1026 602 1032 603
rect 1039 603 1040 604
rect 1044 603 1045 607
rect 1103 607 1109 608
rect 1039 602 1045 603
rect 1078 603 1084 604
rect 1014 598 1020 599
rect 1078 599 1079 603
rect 1083 599 1084 603
rect 1103 603 1104 607
rect 1108 606 1109 607
rect 1134 607 1140 608
rect 1134 606 1135 607
rect 1108 604 1135 606
rect 1108 603 1109 604
rect 1103 602 1109 603
rect 1134 603 1135 604
rect 1139 603 1140 607
rect 1167 607 1173 608
rect 1134 602 1140 603
rect 1142 603 1148 604
rect 1078 598 1084 599
rect 1142 599 1143 603
rect 1147 599 1148 603
rect 1167 603 1168 607
rect 1172 606 1173 607
rect 1182 607 1188 608
rect 1182 606 1183 607
rect 1172 604 1183 606
rect 1172 603 1173 604
rect 1167 602 1173 603
rect 1182 603 1183 604
rect 1187 603 1188 607
rect 1214 607 1221 608
rect 1182 602 1188 603
rect 1190 603 1196 604
rect 1142 598 1148 599
rect 1190 599 1191 603
rect 1195 599 1196 603
rect 1214 603 1215 607
rect 1220 603 1221 607
rect 1214 602 1221 603
rect 1190 598 1196 599
rect 1974 591 1980 592
rect 1582 587 1589 588
rect 570 583 576 584
rect 570 582 571 583
rect 110 580 116 581
rect 110 576 111 580
rect 115 576 116 580
rect 464 580 571 582
rect 110 575 116 576
rect 158 575 165 576
rect 158 571 159 575
rect 164 571 165 575
rect 158 570 165 571
rect 174 575 180 576
rect 174 571 175 575
rect 179 574 180 575
rect 207 575 213 576
rect 207 574 208 575
rect 179 572 208 574
rect 179 571 180 572
rect 174 570 180 571
rect 207 571 208 572
rect 212 571 213 575
rect 207 570 213 571
rect 246 575 252 576
rect 246 571 247 575
rect 251 574 252 575
rect 279 575 285 576
rect 279 574 280 575
rect 251 572 280 574
rect 251 571 252 572
rect 246 570 252 571
rect 279 571 280 572
rect 284 571 285 575
rect 279 570 285 571
rect 318 575 324 576
rect 318 571 319 575
rect 323 574 324 575
rect 351 575 357 576
rect 351 574 352 575
rect 323 572 352 574
rect 323 571 324 572
rect 318 570 324 571
rect 351 571 352 572
rect 356 571 357 575
rect 351 570 357 571
rect 423 575 429 576
rect 423 571 424 575
rect 428 574 429 575
rect 464 574 466 580
rect 570 579 571 580
rect 575 579 576 583
rect 1558 583 1564 584
rect 570 578 576 579
rect 1238 580 1244 581
rect 1238 576 1239 580
rect 1243 576 1244 580
rect 1558 579 1559 583
rect 1563 579 1564 583
rect 1582 583 1583 587
rect 1588 583 1589 587
rect 1610 587 1616 588
rect 1582 582 1589 583
rect 1598 583 1604 584
rect 1558 578 1564 579
rect 1598 579 1599 583
rect 1603 579 1604 583
rect 1610 583 1611 587
rect 1615 586 1616 587
rect 1623 587 1629 588
rect 1623 586 1624 587
rect 1615 584 1624 586
rect 1615 583 1616 584
rect 1610 582 1616 583
rect 1623 583 1624 584
rect 1628 583 1629 587
rect 1650 587 1656 588
rect 1623 582 1629 583
rect 1638 583 1644 584
rect 1598 578 1604 579
rect 1638 579 1639 583
rect 1643 579 1644 583
rect 1650 583 1651 587
rect 1655 586 1656 587
rect 1663 587 1669 588
rect 1663 586 1664 587
rect 1655 584 1664 586
rect 1655 583 1656 584
rect 1650 582 1656 583
rect 1663 583 1664 584
rect 1668 583 1669 587
rect 1703 587 1712 588
rect 1663 582 1669 583
rect 1678 583 1684 584
rect 1638 578 1644 579
rect 1678 579 1679 583
rect 1683 579 1684 583
rect 1703 583 1704 587
rect 1711 583 1712 587
rect 1743 587 1752 588
rect 1703 582 1712 583
rect 1718 583 1724 584
rect 1678 578 1684 579
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1743 583 1744 587
rect 1751 583 1752 587
rect 1783 587 1789 588
rect 1743 582 1752 583
rect 1758 583 1764 584
rect 1718 578 1724 579
rect 1758 579 1759 583
rect 1763 579 1764 583
rect 1783 583 1784 587
rect 1788 586 1789 587
rect 1798 587 1804 588
rect 1798 586 1799 587
rect 1788 584 1799 586
rect 1788 583 1789 584
rect 1783 582 1789 583
rect 1798 583 1799 584
rect 1803 583 1804 587
rect 1831 587 1837 588
rect 1831 586 1832 587
rect 1816 584 1832 586
rect 1798 582 1804 583
rect 1806 583 1812 584
rect 1758 578 1764 579
rect 1806 579 1807 583
rect 1811 579 1812 583
rect 1806 578 1812 579
rect 428 572 466 574
rect 470 575 476 576
rect 428 571 429 572
rect 423 570 429 571
rect 470 571 471 575
rect 475 574 476 575
rect 503 575 509 576
rect 503 574 504 575
rect 475 572 504 574
rect 475 571 476 572
rect 470 570 476 571
rect 503 571 504 572
rect 508 571 509 575
rect 503 570 509 571
rect 578 575 589 576
rect 578 571 579 575
rect 583 571 584 575
rect 588 571 589 575
rect 578 570 589 571
rect 662 575 669 576
rect 662 571 663 575
rect 668 571 669 575
rect 662 570 669 571
rect 710 575 716 576
rect 710 571 711 575
rect 715 574 716 575
rect 743 575 749 576
rect 743 574 744 575
rect 715 572 744 574
rect 715 571 716 572
rect 710 570 716 571
rect 743 571 744 572
rect 748 571 749 575
rect 743 570 749 571
rect 790 575 796 576
rect 790 571 791 575
rect 795 574 796 575
rect 823 575 829 576
rect 823 574 824 575
rect 795 572 824 574
rect 795 571 796 572
rect 790 570 796 571
rect 823 571 824 572
rect 828 571 829 575
rect 823 570 829 571
rect 903 575 909 576
rect 903 571 904 575
rect 908 574 909 575
rect 962 575 968 576
rect 962 574 963 575
rect 908 572 963 574
rect 908 571 909 572
rect 903 570 909 571
rect 962 571 963 572
rect 967 571 968 575
rect 962 570 968 571
rect 975 575 981 576
rect 975 571 976 575
rect 980 574 981 575
rect 1026 575 1032 576
rect 1026 574 1027 575
rect 980 572 1027 574
rect 980 571 981 572
rect 975 570 981 571
rect 1026 571 1027 572
rect 1031 571 1032 575
rect 1026 570 1032 571
rect 1039 575 1045 576
rect 1039 571 1040 575
rect 1044 574 1045 575
rect 1094 575 1100 576
rect 1094 574 1095 575
rect 1044 572 1095 574
rect 1044 571 1045 572
rect 1039 570 1045 571
rect 1094 571 1095 572
rect 1099 571 1100 575
rect 1094 570 1100 571
rect 1102 575 1109 576
rect 1102 571 1103 575
rect 1108 571 1109 575
rect 1102 570 1109 571
rect 1134 575 1140 576
rect 1134 571 1135 575
rect 1139 574 1140 575
rect 1167 575 1173 576
rect 1167 574 1168 575
rect 1139 572 1168 574
rect 1139 571 1140 572
rect 1134 570 1140 571
rect 1167 571 1168 572
rect 1172 571 1173 575
rect 1167 570 1173 571
rect 1182 575 1188 576
rect 1182 571 1183 575
rect 1187 574 1188 575
rect 1215 575 1221 576
rect 1238 575 1244 576
rect 1666 575 1672 576
rect 1215 574 1216 575
rect 1187 572 1216 574
rect 1187 571 1188 572
rect 1182 570 1188 571
rect 1215 571 1216 572
rect 1220 571 1221 575
rect 1215 570 1221 571
rect 1666 571 1667 575
rect 1671 574 1672 575
rect 1816 574 1818 584
rect 1831 583 1832 584
rect 1836 583 1837 587
rect 1879 587 1885 588
rect 1831 582 1837 583
rect 1854 583 1860 584
rect 1854 579 1855 583
rect 1859 579 1860 583
rect 1879 583 1880 587
rect 1884 586 1885 587
rect 1902 587 1908 588
rect 1902 586 1903 587
rect 1884 584 1903 586
rect 1884 583 1885 584
rect 1879 582 1885 583
rect 1902 583 1903 584
rect 1907 583 1908 587
rect 1935 587 1941 588
rect 1902 582 1908 583
rect 1910 583 1916 584
rect 1854 578 1860 579
rect 1910 579 1911 583
rect 1915 579 1916 583
rect 1935 583 1936 587
rect 1940 586 1941 587
rect 1958 587 1964 588
rect 1958 586 1959 587
rect 1940 584 1959 586
rect 1940 583 1941 584
rect 1935 582 1941 583
rect 1958 583 1959 584
rect 1963 583 1964 587
rect 1974 587 1975 591
rect 1979 590 1980 591
rect 1979 588 1995 590
rect 1979 587 1980 588
rect 1974 586 1980 587
rect 1991 587 1997 588
rect 1958 582 1964 583
rect 1966 583 1972 584
rect 1910 578 1916 579
rect 1966 579 1967 583
rect 1971 579 1972 583
rect 1991 583 1992 587
rect 1996 583 1997 587
rect 2042 587 2048 588
rect 1991 582 1997 583
rect 2030 583 2036 584
rect 1966 578 1972 579
rect 2030 579 2031 583
rect 2035 579 2036 583
rect 2042 583 2043 587
rect 2047 586 2048 587
rect 2055 587 2061 588
rect 2055 586 2056 587
rect 2047 584 2056 586
rect 2047 583 2048 584
rect 2042 582 2048 583
rect 2055 583 2056 584
rect 2060 583 2061 587
rect 2106 587 2112 588
rect 2055 582 2061 583
rect 2094 583 2100 584
rect 2030 578 2036 579
rect 2094 579 2095 583
rect 2099 579 2100 583
rect 2106 583 2107 587
rect 2111 586 2112 587
rect 2119 587 2125 588
rect 2119 586 2120 587
rect 2111 584 2120 586
rect 2111 583 2112 584
rect 2106 582 2112 583
rect 2119 583 2120 584
rect 2124 583 2125 587
rect 2191 587 2197 588
rect 2119 582 2125 583
rect 2166 583 2172 584
rect 2094 578 2100 579
rect 2166 579 2167 583
rect 2171 579 2172 583
rect 2191 583 2192 587
rect 2196 586 2197 587
rect 2230 587 2236 588
rect 2230 586 2231 587
rect 2196 584 2231 586
rect 2196 583 2197 584
rect 2191 582 2197 583
rect 2230 583 2231 584
rect 2235 583 2236 587
rect 2263 587 2269 588
rect 2230 582 2236 583
rect 2238 583 2244 584
rect 2166 578 2172 579
rect 2238 579 2239 583
rect 2243 579 2244 583
rect 2263 583 2264 587
rect 2268 586 2269 587
rect 2302 587 2308 588
rect 2302 586 2303 587
rect 2268 584 2303 586
rect 2268 583 2269 584
rect 2263 582 2269 583
rect 2302 583 2303 584
rect 2307 583 2308 587
rect 2335 587 2341 588
rect 2302 582 2308 583
rect 2310 583 2316 584
rect 2238 578 2244 579
rect 2310 579 2311 583
rect 2315 579 2316 583
rect 2335 583 2336 587
rect 2340 586 2341 587
rect 2350 587 2356 588
rect 2350 586 2351 587
rect 2340 584 2351 586
rect 2340 583 2341 584
rect 2335 582 2341 583
rect 2350 583 2351 584
rect 2355 583 2356 587
rect 2383 587 2389 588
rect 2350 582 2356 583
rect 2358 583 2364 584
rect 2310 578 2316 579
rect 2358 579 2359 583
rect 2363 579 2364 583
rect 2383 583 2384 587
rect 2388 586 2389 587
rect 2391 587 2397 588
rect 2391 586 2392 587
rect 2388 584 2392 586
rect 2388 583 2389 584
rect 2383 582 2389 583
rect 2391 583 2392 584
rect 2396 583 2397 587
rect 2391 582 2397 583
rect 2358 578 2364 579
rect 1671 572 1818 574
rect 1671 571 1672 572
rect 1666 570 1672 571
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 110 558 116 559
rect 1238 563 1244 564
rect 1238 559 1239 563
rect 1243 559 1244 563
rect 1746 563 1752 564
rect 1238 558 1244 559
rect 1278 560 1284 561
rect 134 556 140 557
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 182 556 188 557
rect 182 552 183 556
rect 187 552 188 556
rect 182 551 188 552
rect 254 556 260 557
rect 254 552 255 556
rect 259 552 260 556
rect 254 551 260 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 398 556 404 557
rect 398 552 399 556
rect 403 552 404 556
rect 398 551 404 552
rect 478 556 484 557
rect 478 552 479 556
rect 483 552 484 556
rect 478 551 484 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 638 556 644 557
rect 638 552 639 556
rect 643 552 644 556
rect 638 551 644 552
rect 718 556 724 557
rect 718 552 719 556
rect 723 552 724 556
rect 718 551 724 552
rect 798 556 804 557
rect 798 552 799 556
rect 803 552 804 556
rect 798 551 804 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 950 556 956 557
rect 950 552 951 556
rect 955 552 956 556
rect 950 551 956 552
rect 1014 556 1020 557
rect 1014 552 1015 556
rect 1019 552 1020 556
rect 1014 551 1020 552
rect 1078 556 1084 557
rect 1078 552 1079 556
rect 1083 552 1084 556
rect 1078 551 1084 552
rect 1142 556 1148 557
rect 1142 552 1143 556
rect 1147 552 1148 556
rect 1142 551 1148 552
rect 1190 556 1196 557
rect 1190 552 1191 556
rect 1195 552 1196 556
rect 1278 556 1279 560
rect 1283 556 1284 560
rect 1746 559 1747 563
rect 1751 562 1752 563
rect 1751 560 1787 562
rect 1751 559 1752 560
rect 1746 558 1752 559
rect 1785 556 1787 560
rect 2406 560 2412 561
rect 2406 556 2407 560
rect 2411 556 2412 560
rect 1278 555 1284 556
rect 1583 555 1589 556
rect 1190 551 1196 552
rect 1583 551 1584 555
rect 1588 554 1589 555
rect 1610 555 1616 556
rect 1610 554 1611 555
rect 1588 552 1611 554
rect 1588 551 1589 552
rect 1583 550 1589 551
rect 1610 551 1611 552
rect 1615 551 1616 555
rect 1610 550 1616 551
rect 1623 555 1629 556
rect 1623 551 1624 555
rect 1628 554 1629 555
rect 1650 555 1656 556
rect 1650 554 1651 555
rect 1628 552 1651 554
rect 1628 551 1629 552
rect 1623 550 1629 551
rect 1650 551 1651 552
rect 1655 551 1656 555
rect 1650 550 1656 551
rect 1663 555 1672 556
rect 1663 551 1664 555
rect 1671 551 1672 555
rect 1663 550 1672 551
rect 1703 555 1709 556
rect 1703 551 1704 555
rect 1708 554 1709 555
rect 1734 555 1740 556
rect 1734 554 1735 555
rect 1708 552 1735 554
rect 1708 551 1709 552
rect 1703 550 1709 551
rect 1734 551 1735 552
rect 1739 551 1740 555
rect 1734 550 1740 551
rect 1743 555 1749 556
rect 1743 551 1744 555
rect 1748 551 1749 555
rect 1743 550 1749 551
rect 1783 555 1789 556
rect 1783 551 1784 555
rect 1788 551 1789 555
rect 1783 550 1789 551
rect 1798 555 1804 556
rect 1798 551 1799 555
rect 1803 554 1804 555
rect 1831 555 1837 556
rect 1831 554 1832 555
rect 1803 552 1832 554
rect 1803 551 1804 552
rect 1798 550 1804 551
rect 1831 551 1832 552
rect 1836 551 1837 555
rect 1831 550 1837 551
rect 1879 555 1885 556
rect 1879 551 1880 555
rect 1884 554 1885 555
rect 1890 555 1896 556
rect 1890 554 1891 555
rect 1884 552 1891 554
rect 1884 551 1885 552
rect 1879 550 1885 551
rect 1890 551 1891 552
rect 1895 551 1896 555
rect 1890 550 1896 551
rect 1902 555 1908 556
rect 1902 551 1903 555
rect 1907 554 1908 555
rect 1935 555 1941 556
rect 1935 554 1936 555
rect 1907 552 1936 554
rect 1907 551 1908 552
rect 1902 550 1908 551
rect 1935 551 1936 552
rect 1940 551 1941 555
rect 1935 550 1941 551
rect 1991 555 1997 556
rect 1991 551 1992 555
rect 1996 554 1997 555
rect 2042 555 2048 556
rect 2042 554 2043 555
rect 1996 552 2043 554
rect 1996 551 1997 552
rect 1991 550 1997 551
rect 2042 551 2043 552
rect 2047 551 2048 555
rect 2042 550 2048 551
rect 2055 555 2061 556
rect 2055 551 2056 555
rect 2060 554 2061 555
rect 2106 555 2112 556
rect 2106 554 2107 555
rect 2060 552 2107 554
rect 2060 551 2061 552
rect 2055 550 2061 551
rect 2106 551 2107 552
rect 2111 551 2112 555
rect 2106 550 2112 551
rect 2119 555 2128 556
rect 2119 551 2120 555
rect 2127 551 2128 555
rect 2119 550 2128 551
rect 2191 555 2197 556
rect 2191 551 2192 555
rect 2196 554 2197 555
rect 2215 555 2221 556
rect 2215 554 2216 555
rect 2196 552 2216 554
rect 2196 551 2197 552
rect 2191 550 2197 551
rect 2215 551 2216 552
rect 2220 551 2221 555
rect 2215 550 2221 551
rect 2230 555 2236 556
rect 2230 551 2231 555
rect 2235 554 2236 555
rect 2263 555 2269 556
rect 2263 554 2264 555
rect 2235 552 2264 554
rect 2235 551 2236 552
rect 2230 550 2236 551
rect 2263 551 2264 552
rect 2268 551 2269 555
rect 2263 550 2269 551
rect 2335 555 2344 556
rect 2335 551 2336 555
rect 2343 551 2344 555
rect 2335 550 2344 551
rect 2350 555 2356 556
rect 2350 551 2351 555
rect 2355 554 2356 555
rect 2383 555 2389 556
rect 2406 555 2412 556
rect 2383 554 2384 555
rect 2355 552 2384 554
rect 2355 551 2356 552
rect 2350 550 2356 551
rect 2383 551 2384 552
rect 2388 551 2389 555
rect 2383 550 2389 551
rect 1706 547 1712 548
rect 1278 543 1284 544
rect 150 540 156 541
rect 150 536 151 540
rect 155 536 156 540
rect 150 535 156 536
rect 222 540 228 541
rect 222 536 223 540
rect 227 536 228 540
rect 222 535 228 536
rect 286 540 292 541
rect 286 536 287 540
rect 291 536 292 540
rect 286 535 292 536
rect 350 540 356 541
rect 350 536 351 540
rect 355 536 356 540
rect 350 535 356 536
rect 414 540 420 541
rect 414 536 415 540
rect 419 536 420 540
rect 414 535 420 536
rect 478 540 484 541
rect 478 536 479 540
rect 483 536 484 540
rect 478 535 484 536
rect 550 540 556 541
rect 550 536 551 540
rect 555 536 556 540
rect 550 535 556 536
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 694 540 700 541
rect 694 536 695 540
rect 699 536 700 540
rect 694 535 700 536
rect 766 540 772 541
rect 766 536 767 540
rect 771 536 772 540
rect 766 535 772 536
rect 838 540 844 541
rect 838 536 839 540
rect 843 536 844 540
rect 838 535 844 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 998 540 1004 541
rect 998 536 999 540
rect 1003 536 1004 540
rect 998 535 1004 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1278 539 1279 543
rect 1283 539 1284 543
rect 1706 543 1707 547
rect 1711 546 1712 547
rect 1745 546 1747 550
rect 1711 544 1747 546
rect 1711 543 1712 544
rect 1706 542 1712 543
rect 2406 543 2412 544
rect 1278 538 1284 539
rect 2406 539 2407 543
rect 2411 539 2412 543
rect 2406 538 2412 539
rect 1078 535 1084 536
rect 1558 536 1564 537
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 1238 533 1244 534
rect 1238 529 1239 533
rect 1243 529 1244 533
rect 1558 532 1559 536
rect 1563 532 1564 536
rect 1558 531 1564 532
rect 1598 536 1604 537
rect 1598 532 1599 536
rect 1603 532 1604 536
rect 1598 531 1604 532
rect 1638 536 1644 537
rect 1638 532 1639 536
rect 1643 532 1644 536
rect 1638 531 1644 532
rect 1678 536 1684 537
rect 1678 532 1679 536
rect 1683 532 1684 536
rect 1678 531 1684 532
rect 1718 536 1724 537
rect 1718 532 1719 536
rect 1723 532 1724 536
rect 1718 531 1724 532
rect 1758 536 1764 537
rect 1758 532 1759 536
rect 1763 532 1764 536
rect 1758 531 1764 532
rect 1806 536 1812 537
rect 1806 532 1807 536
rect 1811 532 1812 536
rect 1806 531 1812 532
rect 1854 536 1860 537
rect 1854 532 1855 536
rect 1859 532 1860 536
rect 1854 531 1860 532
rect 1910 536 1916 537
rect 1910 532 1911 536
rect 1915 532 1916 536
rect 1910 531 1916 532
rect 1966 536 1972 537
rect 1966 532 1967 536
rect 1971 532 1972 536
rect 1966 531 1972 532
rect 2030 536 2036 537
rect 2030 532 2031 536
rect 2035 532 2036 536
rect 2030 531 2036 532
rect 2094 536 2100 537
rect 2094 532 2095 536
rect 2099 532 2100 536
rect 2094 531 2100 532
rect 2166 536 2172 537
rect 2166 532 2167 536
rect 2171 532 2172 536
rect 2166 531 2172 532
rect 2238 536 2244 537
rect 2238 532 2239 536
rect 2243 532 2244 536
rect 2238 531 2244 532
rect 2310 536 2316 537
rect 2310 532 2311 536
rect 2315 532 2316 536
rect 2310 531 2316 532
rect 2358 536 2364 537
rect 2358 532 2359 536
rect 2363 532 2364 536
rect 2358 531 2364 532
rect 1238 528 1244 529
rect 810 527 816 528
rect 810 526 811 527
rect 679 524 811 526
rect 679 522 681 524
rect 810 523 811 524
rect 815 523 816 527
rect 810 522 816 523
rect 1406 524 1412 525
rect 664 520 681 522
rect 1406 520 1407 524
rect 1411 520 1412 524
rect 175 519 181 520
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 175 515 176 519
rect 180 515 181 519
rect 175 514 181 515
rect 183 519 189 520
rect 183 515 184 519
rect 188 518 189 519
rect 247 519 253 520
rect 247 518 248 519
rect 188 516 248 518
rect 188 515 189 516
rect 183 514 189 515
rect 247 515 248 516
rect 252 515 253 519
rect 247 514 253 515
rect 311 519 317 520
rect 311 515 312 519
rect 316 518 317 519
rect 338 519 344 520
rect 338 518 339 519
rect 316 516 339 518
rect 316 515 317 516
rect 311 514 317 515
rect 338 515 339 516
rect 343 515 344 519
rect 338 514 344 515
rect 375 519 381 520
rect 375 515 376 519
rect 380 515 381 519
rect 375 514 381 515
rect 383 519 389 520
rect 383 515 384 519
rect 388 518 389 519
rect 439 519 445 520
rect 439 518 440 519
rect 388 516 440 518
rect 388 515 389 516
rect 383 514 389 515
rect 439 515 440 516
rect 444 515 445 519
rect 439 514 445 515
rect 447 519 453 520
rect 447 515 448 519
rect 452 518 453 519
rect 503 519 509 520
rect 503 518 504 519
rect 452 516 504 518
rect 452 515 453 516
rect 447 514 453 515
rect 503 515 504 516
rect 508 515 509 519
rect 503 514 509 515
rect 511 519 517 520
rect 511 515 512 519
rect 516 518 517 519
rect 575 519 581 520
rect 575 518 576 519
rect 516 516 576 518
rect 516 515 517 516
rect 511 514 517 515
rect 575 515 576 516
rect 580 515 581 519
rect 575 514 581 515
rect 647 519 653 520
rect 647 515 648 519
rect 652 518 653 519
rect 664 518 666 520
rect 719 519 725 520
rect 719 518 720 519
rect 652 516 666 518
rect 679 516 720 518
rect 652 515 653 516
rect 647 514 653 515
rect 670 515 676 516
rect 110 511 116 512
rect 176 510 178 514
rect 310 511 316 512
rect 310 510 311 511
rect 176 508 311 510
rect 310 507 311 508
rect 315 507 316 511
rect 376 510 378 514
rect 462 511 468 512
rect 462 510 463 511
rect 376 508 463 510
rect 310 506 316 507
rect 462 507 463 508
rect 467 507 468 511
rect 670 511 671 515
rect 675 514 676 515
rect 679 514 681 516
rect 719 515 720 516
rect 724 515 725 519
rect 719 514 725 515
rect 727 519 733 520
rect 727 515 728 519
rect 732 518 733 519
rect 791 519 797 520
rect 791 518 792 519
rect 732 516 792 518
rect 732 515 733 516
rect 727 514 733 515
rect 791 515 792 516
rect 796 515 797 519
rect 791 514 797 515
rect 830 519 836 520
rect 830 515 831 519
rect 835 518 836 519
rect 863 519 869 520
rect 863 518 864 519
rect 835 516 864 518
rect 835 515 836 516
rect 830 514 836 515
rect 863 515 864 516
rect 868 515 869 519
rect 863 514 869 515
rect 943 519 949 520
rect 943 515 944 519
rect 948 518 949 519
rect 974 519 980 520
rect 974 518 975 519
rect 948 516 975 518
rect 948 515 949 516
rect 943 514 949 515
rect 974 515 975 516
rect 979 515 980 519
rect 974 514 980 515
rect 982 519 988 520
rect 982 515 983 519
rect 987 518 988 519
rect 1023 519 1029 520
rect 1023 518 1024 519
rect 987 516 1024 518
rect 987 515 988 516
rect 982 514 988 515
rect 1023 515 1024 516
rect 1028 515 1029 519
rect 1023 514 1029 515
rect 1031 519 1037 520
rect 1031 515 1032 519
rect 1036 518 1037 519
rect 1103 519 1109 520
rect 1406 519 1412 520
rect 1446 524 1452 525
rect 1446 520 1447 524
rect 1451 520 1452 524
rect 1446 519 1452 520
rect 1486 524 1492 525
rect 1486 520 1487 524
rect 1491 520 1492 524
rect 1486 519 1492 520
rect 1534 524 1540 525
rect 1534 520 1535 524
rect 1539 520 1540 524
rect 1534 519 1540 520
rect 1590 524 1596 525
rect 1590 520 1591 524
rect 1595 520 1596 524
rect 1590 519 1596 520
rect 1646 524 1652 525
rect 1646 520 1647 524
rect 1651 520 1652 524
rect 1646 519 1652 520
rect 1710 524 1716 525
rect 1710 520 1711 524
rect 1715 520 1716 524
rect 1710 519 1716 520
rect 1782 524 1788 525
rect 1782 520 1783 524
rect 1787 520 1788 524
rect 1782 519 1788 520
rect 1862 524 1868 525
rect 1862 520 1863 524
rect 1867 520 1868 524
rect 1862 519 1868 520
rect 1942 524 1948 525
rect 1942 520 1943 524
rect 1947 520 1948 524
rect 1942 519 1948 520
rect 2022 524 2028 525
rect 2022 520 2023 524
rect 2027 520 2028 524
rect 2022 519 2028 520
rect 2102 524 2108 525
rect 2102 520 2103 524
rect 2107 520 2108 524
rect 2102 519 2108 520
rect 2190 524 2196 525
rect 2190 520 2191 524
rect 2195 520 2196 524
rect 2190 519 2196 520
rect 2286 524 2292 525
rect 2286 520 2287 524
rect 2291 520 2292 524
rect 2286 519 2292 520
rect 2358 524 2364 525
rect 2358 520 2359 524
rect 2363 520 2364 524
rect 2358 519 2364 520
rect 1103 518 1104 519
rect 1036 516 1104 518
rect 1036 515 1037 516
rect 1031 514 1037 515
rect 1103 515 1104 516
rect 1108 515 1109 519
rect 1278 517 1284 518
rect 1103 514 1109 515
rect 1238 516 1244 517
rect 675 512 681 514
rect 1238 512 1239 516
rect 1243 512 1244 516
rect 1278 513 1279 517
rect 1283 513 1284 517
rect 1278 512 1284 513
rect 2406 517 2412 518
rect 2406 513 2407 517
rect 2411 513 2412 517
rect 2406 512 2412 513
rect 675 511 676 512
rect 1238 511 1244 512
rect 670 510 676 511
rect 462 506 468 507
rect 1431 503 1437 504
rect 1278 500 1284 501
rect 1278 496 1279 500
rect 1283 496 1284 500
rect 1431 499 1432 503
rect 1436 502 1437 503
rect 1454 503 1460 504
rect 1436 500 1450 502
rect 1436 499 1437 500
rect 1431 498 1437 499
rect 830 495 836 496
rect 1278 495 1284 496
rect 150 493 156 494
rect 150 489 151 493
rect 155 489 156 493
rect 150 488 156 489
rect 222 493 228 494
rect 222 489 223 493
rect 227 489 228 493
rect 222 488 228 489
rect 286 493 292 494
rect 286 489 287 493
rect 291 489 292 493
rect 286 488 292 489
rect 350 493 356 494
rect 350 489 351 493
rect 355 489 356 493
rect 350 488 356 489
rect 414 493 420 494
rect 414 489 415 493
rect 419 489 420 493
rect 414 488 420 489
rect 478 493 484 494
rect 478 489 479 493
rect 483 489 484 493
rect 478 488 484 489
rect 550 493 556 494
rect 550 489 551 493
rect 555 489 556 493
rect 550 488 556 489
rect 622 493 628 494
rect 622 489 623 493
rect 627 489 628 493
rect 622 488 628 489
rect 694 493 700 494
rect 694 489 695 493
rect 699 489 700 493
rect 694 488 700 489
rect 766 493 772 494
rect 766 489 767 493
rect 771 489 772 493
rect 830 491 831 495
rect 835 491 836 495
rect 1448 494 1450 500
rect 1454 499 1455 503
rect 1459 502 1460 503
rect 1471 503 1477 504
rect 1471 502 1472 503
rect 1459 500 1472 502
rect 1459 499 1460 500
rect 1454 498 1460 499
rect 1471 499 1472 500
rect 1476 499 1477 503
rect 1471 498 1477 499
rect 1494 503 1500 504
rect 1494 499 1495 503
rect 1499 502 1500 503
rect 1511 503 1517 504
rect 1511 502 1512 503
rect 1499 500 1512 502
rect 1499 499 1500 500
rect 1494 498 1500 499
rect 1511 499 1512 500
rect 1516 499 1517 503
rect 1511 498 1517 499
rect 1519 503 1525 504
rect 1519 499 1520 503
rect 1524 502 1525 503
rect 1559 503 1565 504
rect 1559 502 1560 503
rect 1524 500 1560 502
rect 1524 499 1525 500
rect 1519 498 1525 499
rect 1559 499 1560 500
rect 1564 499 1565 503
rect 1559 498 1565 499
rect 1567 503 1573 504
rect 1567 499 1568 503
rect 1572 502 1573 503
rect 1615 503 1621 504
rect 1615 502 1616 503
rect 1572 500 1616 502
rect 1572 499 1573 500
rect 1567 498 1573 499
rect 1615 499 1616 500
rect 1620 499 1621 503
rect 1615 498 1621 499
rect 1623 503 1629 504
rect 1623 499 1624 503
rect 1628 502 1629 503
rect 1671 503 1677 504
rect 1671 502 1672 503
rect 1628 500 1672 502
rect 1628 499 1629 500
rect 1623 498 1629 499
rect 1671 499 1672 500
rect 1676 499 1677 503
rect 1671 498 1677 499
rect 1679 503 1685 504
rect 1679 499 1680 503
rect 1684 502 1685 503
rect 1735 503 1741 504
rect 1735 502 1736 503
rect 1684 500 1736 502
rect 1684 499 1685 500
rect 1679 498 1685 499
rect 1735 499 1736 500
rect 1740 499 1741 503
rect 1735 498 1741 499
rect 1807 503 1813 504
rect 1807 499 1808 503
rect 1812 502 1813 503
rect 1878 503 1884 504
rect 1878 502 1879 503
rect 1812 500 1879 502
rect 1812 499 1813 500
rect 1807 498 1813 499
rect 1878 499 1879 500
rect 1883 499 1884 503
rect 1878 498 1884 499
rect 1887 503 1893 504
rect 1887 499 1888 503
rect 1892 502 1893 503
rect 1950 503 1956 504
rect 1950 502 1951 503
rect 1892 500 1951 502
rect 1892 499 1893 500
rect 1887 498 1893 499
rect 1950 499 1951 500
rect 1955 499 1956 503
rect 1950 498 1956 499
rect 1958 503 1964 504
rect 1958 499 1959 503
rect 1963 502 1964 503
rect 1967 503 1973 504
rect 1967 502 1968 503
rect 1963 500 1968 502
rect 1963 499 1964 500
rect 1958 498 1964 499
rect 1967 499 1968 500
rect 1972 499 1973 503
rect 1967 498 1973 499
rect 2038 503 2044 504
rect 2038 499 2039 503
rect 2043 502 2044 503
rect 2047 503 2053 504
rect 2047 502 2048 503
rect 2043 500 2048 502
rect 2043 499 2044 500
rect 2038 498 2044 499
rect 2047 499 2048 500
rect 2052 499 2053 503
rect 2047 498 2053 499
rect 2055 503 2061 504
rect 2055 499 2056 503
rect 2060 502 2061 503
rect 2127 503 2133 504
rect 2127 502 2128 503
rect 2060 500 2128 502
rect 2060 499 2061 500
rect 2055 498 2061 499
rect 2127 499 2128 500
rect 2132 499 2133 503
rect 2127 498 2133 499
rect 2215 503 2221 504
rect 2215 499 2216 503
rect 2220 502 2221 503
rect 2294 503 2300 504
rect 2294 502 2295 503
rect 2220 500 2295 502
rect 2220 499 2221 500
rect 2215 498 2221 499
rect 2294 499 2295 500
rect 2299 499 2300 503
rect 2294 498 2300 499
rect 2302 503 2308 504
rect 2302 499 2303 503
rect 2307 502 2308 503
rect 2311 503 2317 504
rect 2311 502 2312 503
rect 2307 500 2312 502
rect 2307 499 2308 500
rect 2302 498 2308 499
rect 2311 499 2312 500
rect 2316 499 2317 503
rect 2311 498 2317 499
rect 2382 503 2389 504
rect 2382 499 2383 503
rect 2388 499 2389 503
rect 2382 498 2389 499
rect 2406 500 2412 501
rect 2406 496 2407 500
rect 2411 496 2412 500
rect 1758 495 1764 496
rect 2406 495 2412 496
rect 1758 494 1759 495
rect 830 490 836 491
rect 838 493 844 494
rect 766 488 772 489
rect 796 488 834 490
rect 838 489 839 493
rect 843 489 844 493
rect 838 488 844 489
rect 918 493 924 494
rect 918 489 919 493
rect 923 489 924 493
rect 918 488 924 489
rect 998 493 1004 494
rect 998 489 999 493
rect 1003 489 1004 493
rect 998 488 1004 489
rect 1078 493 1084 494
rect 1078 489 1079 493
rect 1083 489 1084 493
rect 1448 492 1759 494
rect 1758 491 1759 492
rect 1763 491 1764 495
rect 1758 490 1764 491
rect 1078 488 1084 489
rect 175 487 181 488
rect 175 483 176 487
rect 180 486 181 487
rect 183 487 189 488
rect 183 486 184 487
rect 180 484 184 486
rect 180 483 181 484
rect 175 482 181 483
rect 183 483 184 484
rect 188 483 189 487
rect 183 482 189 483
rect 247 487 253 488
rect 247 483 248 487
rect 252 486 253 487
rect 262 487 268 488
rect 262 486 263 487
rect 252 484 263 486
rect 252 483 253 484
rect 247 482 253 483
rect 262 483 263 484
rect 267 483 268 487
rect 262 482 268 483
rect 310 487 317 488
rect 310 483 311 487
rect 316 483 317 487
rect 310 482 317 483
rect 375 487 381 488
rect 375 483 376 487
rect 380 486 381 487
rect 383 487 389 488
rect 383 486 384 487
rect 380 484 384 486
rect 380 483 381 484
rect 375 482 381 483
rect 383 483 384 484
rect 388 483 389 487
rect 383 482 389 483
rect 439 487 445 488
rect 439 483 440 487
rect 444 486 445 487
rect 447 487 453 488
rect 447 486 448 487
rect 444 484 448 486
rect 444 483 445 484
rect 439 482 445 483
rect 447 483 448 484
rect 452 483 453 487
rect 447 482 453 483
rect 503 487 509 488
rect 503 483 504 487
rect 508 486 509 487
rect 511 487 517 488
rect 511 486 512 487
rect 508 484 512 486
rect 508 483 509 484
rect 503 482 509 483
rect 511 483 512 484
rect 516 483 517 487
rect 511 482 517 483
rect 575 487 584 488
rect 575 483 576 487
rect 583 483 584 487
rect 575 482 584 483
rect 647 487 653 488
rect 647 483 648 487
rect 652 486 653 487
rect 670 487 676 488
rect 670 486 671 487
rect 652 484 671 486
rect 652 483 653 484
rect 647 482 653 483
rect 670 483 671 484
rect 675 483 676 487
rect 670 482 676 483
rect 719 487 725 488
rect 719 483 720 487
rect 724 486 725 487
rect 727 487 733 488
rect 727 486 728 487
rect 724 484 728 486
rect 724 483 725 484
rect 719 482 725 483
rect 727 483 728 484
rect 732 483 733 487
rect 727 482 733 483
rect 791 487 798 488
rect 791 483 792 487
rect 796 484 798 487
rect 863 487 869 488
rect 863 486 864 487
rect 800 484 864 486
rect 796 483 797 484
rect 791 482 797 483
rect 658 479 664 480
rect 658 475 659 479
rect 663 478 664 479
rect 800 478 802 484
rect 863 483 864 484
rect 868 483 869 487
rect 863 482 869 483
rect 943 487 949 488
rect 943 483 944 487
rect 948 486 949 487
rect 982 487 988 488
rect 982 486 983 487
rect 948 484 983 486
rect 948 483 949 484
rect 943 482 949 483
rect 982 483 983 484
rect 987 483 988 487
rect 982 482 988 483
rect 1023 487 1029 488
rect 1023 483 1024 487
rect 1028 486 1029 487
rect 1031 487 1037 488
rect 1031 486 1032 487
rect 1028 484 1032 486
rect 1028 483 1029 484
rect 1023 482 1029 483
rect 1031 483 1032 484
rect 1036 483 1037 487
rect 1031 482 1037 483
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 486 1100 487
rect 1103 487 1109 488
rect 1103 486 1104 487
rect 1099 484 1104 486
rect 1099 483 1100 484
rect 1094 482 1100 483
rect 1103 483 1104 484
rect 1108 483 1109 487
rect 1103 482 1109 483
rect 663 476 802 478
rect 1406 477 1412 478
rect 663 475 664 476
rect 658 474 664 475
rect 1406 473 1407 477
rect 1411 473 1412 477
rect 1406 472 1412 473
rect 1446 477 1452 478
rect 1446 473 1447 477
rect 1451 473 1452 477
rect 1446 472 1452 473
rect 1486 477 1492 478
rect 1486 473 1487 477
rect 1491 473 1492 477
rect 1486 472 1492 473
rect 1534 477 1540 478
rect 1534 473 1535 477
rect 1539 473 1540 477
rect 1534 472 1540 473
rect 1590 477 1596 478
rect 1590 473 1591 477
rect 1595 473 1596 477
rect 1590 472 1596 473
rect 1646 477 1652 478
rect 1646 473 1647 477
rect 1651 473 1652 477
rect 1646 472 1652 473
rect 1710 477 1716 478
rect 1710 473 1711 477
rect 1715 473 1716 477
rect 1710 472 1716 473
rect 1782 477 1788 478
rect 1782 473 1783 477
rect 1787 473 1788 477
rect 1782 472 1788 473
rect 1862 477 1868 478
rect 1862 473 1863 477
rect 1867 473 1868 477
rect 1862 472 1868 473
rect 1942 477 1948 478
rect 1942 473 1943 477
rect 1947 473 1948 477
rect 1942 472 1948 473
rect 2022 477 2028 478
rect 2022 473 2023 477
rect 2027 473 2028 477
rect 2022 472 2028 473
rect 2102 477 2108 478
rect 2102 473 2103 477
rect 2107 473 2108 477
rect 2102 472 2108 473
rect 2190 477 2196 478
rect 2190 473 2191 477
rect 2195 473 2196 477
rect 2190 472 2196 473
rect 2286 477 2292 478
rect 2286 473 2287 477
rect 2291 473 2292 477
rect 2286 472 2292 473
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 294 471 300 472
rect 294 470 295 471
rect 263 469 295 470
rect 263 465 264 469
rect 268 468 295 469
rect 268 465 269 468
rect 294 467 295 468
rect 299 467 300 471
rect 1431 471 1437 472
rect 294 466 300 467
rect 303 467 309 468
rect 263 464 269 465
rect 238 463 244 464
rect 238 459 239 463
rect 243 459 244 463
rect 238 458 244 459
rect 278 463 284 464
rect 278 459 279 463
rect 283 459 284 463
rect 303 463 304 467
rect 308 466 309 467
rect 318 467 324 468
rect 318 466 319 467
rect 308 464 319 466
rect 308 463 309 464
rect 303 462 309 463
rect 318 463 319 464
rect 323 463 324 467
rect 351 467 357 468
rect 318 462 324 463
rect 326 463 332 464
rect 278 458 284 459
rect 326 459 327 463
rect 331 459 332 463
rect 351 463 352 467
rect 356 466 357 467
rect 374 467 380 468
rect 374 466 375 467
rect 356 464 375 466
rect 356 463 357 464
rect 351 462 357 463
rect 374 463 375 464
rect 379 463 380 467
rect 406 467 413 468
rect 374 462 380 463
rect 382 463 388 464
rect 326 458 332 459
rect 382 459 383 463
rect 387 459 388 463
rect 406 463 407 467
rect 412 463 413 467
rect 462 467 469 468
rect 406 462 413 463
rect 438 463 444 464
rect 382 458 388 459
rect 438 459 439 463
rect 443 459 444 463
rect 462 463 463 467
rect 468 463 469 467
rect 514 467 520 468
rect 462 462 469 463
rect 502 463 508 464
rect 438 458 444 459
rect 502 459 503 463
rect 507 459 508 463
rect 514 463 515 467
rect 519 466 520 467
rect 527 467 533 468
rect 527 466 528 467
rect 519 464 528 466
rect 519 463 520 464
rect 514 462 520 463
rect 527 463 528 464
rect 532 463 533 467
rect 578 467 584 468
rect 527 462 533 463
rect 566 463 572 464
rect 502 458 508 459
rect 566 459 567 463
rect 571 459 572 463
rect 578 463 579 467
rect 583 466 584 467
rect 591 467 597 468
rect 591 466 592 467
rect 583 464 592 466
rect 583 463 584 464
rect 578 462 584 463
rect 591 463 592 464
rect 596 463 597 467
rect 655 467 661 468
rect 591 462 597 463
rect 630 463 636 464
rect 566 458 572 459
rect 630 459 631 463
rect 635 459 636 463
rect 655 463 656 467
rect 660 466 661 467
rect 686 467 692 468
rect 686 466 687 467
rect 660 464 687 466
rect 660 463 661 464
rect 655 462 661 463
rect 686 463 687 464
rect 691 463 692 467
rect 719 467 725 468
rect 686 462 692 463
rect 694 463 700 464
rect 630 458 636 459
rect 694 459 695 463
rect 699 459 700 463
rect 719 463 720 467
rect 724 466 725 467
rect 750 467 756 468
rect 750 466 751 467
rect 724 464 751 466
rect 724 463 725 464
rect 719 462 725 463
rect 750 463 751 464
rect 755 463 756 467
rect 783 467 789 468
rect 750 462 756 463
rect 758 463 764 464
rect 694 458 700 459
rect 758 459 759 463
rect 763 459 764 463
rect 783 463 784 467
rect 788 466 789 467
rect 814 467 820 468
rect 814 466 815 467
rect 788 464 815 466
rect 788 463 789 464
rect 783 462 789 463
rect 814 463 815 464
rect 819 463 820 467
rect 847 467 853 468
rect 814 462 820 463
rect 822 463 828 464
rect 758 458 764 459
rect 822 459 823 463
rect 827 459 828 463
rect 847 463 848 467
rect 852 466 853 467
rect 878 467 884 468
rect 878 466 879 467
rect 852 464 879 466
rect 852 463 853 464
rect 847 462 853 463
rect 878 463 879 464
rect 883 463 884 467
rect 898 467 904 468
rect 878 462 884 463
rect 886 463 892 464
rect 822 458 828 459
rect 886 459 887 463
rect 891 459 892 463
rect 898 463 899 467
rect 903 466 904 467
rect 911 467 917 468
rect 911 466 912 467
rect 903 464 912 466
rect 903 463 904 464
rect 898 462 904 463
rect 911 463 912 464
rect 916 463 917 467
rect 974 467 981 468
rect 911 462 917 463
rect 950 463 956 464
rect 886 458 892 459
rect 950 459 951 463
rect 955 459 956 463
rect 974 463 975 467
rect 980 463 981 467
rect 1026 467 1032 468
rect 974 462 981 463
rect 1014 463 1020 464
rect 950 458 956 459
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1026 463 1027 467
rect 1031 466 1032 467
rect 1039 467 1045 468
rect 1039 466 1040 467
rect 1031 464 1040 466
rect 1031 463 1032 464
rect 1026 462 1032 463
rect 1039 463 1040 464
rect 1044 463 1045 467
rect 1431 467 1432 471
rect 1436 470 1437 471
rect 1454 471 1460 472
rect 1454 470 1455 471
rect 1436 468 1455 470
rect 1436 467 1437 468
rect 1431 466 1437 467
rect 1454 467 1455 468
rect 1459 467 1460 471
rect 1454 466 1460 467
rect 1471 471 1477 472
rect 1471 467 1472 471
rect 1476 470 1477 471
rect 1494 471 1500 472
rect 1494 470 1495 471
rect 1476 468 1495 470
rect 1476 467 1477 468
rect 1471 466 1477 467
rect 1494 467 1495 468
rect 1499 467 1500 471
rect 1494 466 1500 467
rect 1511 471 1517 472
rect 1511 467 1512 471
rect 1516 470 1517 471
rect 1519 471 1525 472
rect 1519 470 1520 471
rect 1516 468 1520 470
rect 1516 467 1517 468
rect 1511 466 1517 467
rect 1519 467 1520 468
rect 1524 467 1525 471
rect 1519 466 1525 467
rect 1559 471 1565 472
rect 1559 467 1560 471
rect 1564 470 1565 471
rect 1567 471 1573 472
rect 1567 470 1568 471
rect 1564 468 1568 470
rect 1564 467 1565 468
rect 1559 466 1565 467
rect 1567 467 1568 468
rect 1572 467 1573 471
rect 1567 466 1573 467
rect 1615 471 1621 472
rect 1615 467 1616 471
rect 1620 470 1621 471
rect 1623 471 1629 472
rect 1623 470 1624 471
rect 1620 468 1624 470
rect 1620 467 1621 468
rect 1615 466 1621 467
rect 1623 467 1624 468
rect 1628 467 1629 471
rect 1623 466 1629 467
rect 1671 471 1677 472
rect 1671 467 1672 471
rect 1676 470 1677 471
rect 1679 471 1685 472
rect 1679 470 1680 471
rect 1676 468 1680 470
rect 1676 467 1677 468
rect 1671 466 1677 467
rect 1679 467 1680 468
rect 1684 467 1685 471
rect 1679 466 1685 467
rect 1734 471 1741 472
rect 1734 467 1735 471
rect 1740 467 1741 471
rect 1734 466 1741 467
rect 1807 471 1813 472
rect 1807 467 1808 471
rect 1812 470 1813 471
rect 1854 471 1860 472
rect 1854 470 1855 471
rect 1812 468 1855 470
rect 1812 467 1813 468
rect 1807 466 1813 467
rect 1854 467 1855 468
rect 1859 467 1860 471
rect 1854 466 1860 467
rect 1878 471 1884 472
rect 1878 467 1879 471
rect 1883 470 1884 471
rect 1887 471 1893 472
rect 1887 470 1888 471
rect 1883 468 1888 470
rect 1883 467 1884 468
rect 1878 466 1884 467
rect 1887 467 1888 468
rect 1892 467 1893 471
rect 1887 466 1893 467
rect 1950 471 1956 472
rect 1950 467 1951 471
rect 1955 470 1956 471
rect 1967 471 1973 472
rect 1967 470 1968 471
rect 1955 468 1968 470
rect 1955 467 1956 468
rect 1950 466 1956 467
rect 1967 467 1968 468
rect 1972 467 1973 471
rect 1967 466 1973 467
rect 2047 471 2053 472
rect 2047 467 2048 471
rect 2052 470 2053 471
rect 2055 471 2061 472
rect 2055 470 2056 471
rect 2052 468 2056 470
rect 2052 467 2053 468
rect 2047 466 2053 467
rect 2055 467 2056 468
rect 2060 467 2061 471
rect 2055 466 2061 467
rect 2122 471 2133 472
rect 2122 467 2123 471
rect 2127 467 2128 471
rect 2132 467 2133 471
rect 2215 471 2221 472
rect 2215 470 2216 471
rect 2122 466 2133 467
rect 2136 468 2216 470
rect 1039 462 1045 463
rect 2110 463 2116 464
rect 1014 458 1020 459
rect 2110 459 2111 463
rect 2115 462 2116 463
rect 2136 462 2138 468
rect 2215 467 2216 468
rect 2220 467 2221 471
rect 2215 466 2221 467
rect 2294 471 2300 472
rect 2294 467 2295 471
rect 2299 470 2300 471
rect 2311 471 2317 472
rect 2311 470 2312 471
rect 2299 468 2312 470
rect 2299 467 2300 468
rect 2294 466 2300 467
rect 2311 467 2312 468
rect 2316 467 2317 471
rect 2311 466 2317 467
rect 2338 471 2344 472
rect 2338 467 2339 471
rect 2343 470 2344 471
rect 2383 471 2389 472
rect 2383 470 2384 471
rect 2343 468 2384 470
rect 2343 467 2344 468
rect 2338 466 2344 467
rect 2383 467 2384 468
rect 2388 467 2389 471
rect 2383 466 2389 467
rect 2115 460 2138 462
rect 2115 459 2116 460
rect 2110 458 2116 459
rect 1358 455 1364 456
rect 1358 454 1359 455
rect 1336 452 1359 454
rect 1327 451 1333 452
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1327 447 1328 451
rect 1332 450 1333 451
rect 1336 450 1338 452
rect 1358 451 1359 452
rect 1363 451 1364 455
rect 1398 455 1404 456
rect 1398 454 1399 455
rect 1376 452 1399 454
rect 1358 450 1364 451
rect 1367 451 1373 452
rect 1332 448 1338 450
rect 1332 447 1333 448
rect 1327 446 1333 447
rect 1342 447 1348 448
rect 1302 442 1308 443
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1367 447 1368 451
rect 1372 450 1373 451
rect 1376 450 1378 452
rect 1398 451 1399 452
rect 1403 451 1404 455
rect 2038 455 2044 456
rect 2038 454 2039 455
rect 2023 453 2039 454
rect 1398 450 1404 451
rect 1407 451 1413 452
rect 1372 448 1378 450
rect 1372 447 1373 448
rect 1367 446 1373 447
rect 1382 447 1388 448
rect 1342 442 1348 443
rect 1382 443 1383 447
rect 1387 443 1388 447
rect 1407 447 1408 451
rect 1412 450 1413 451
rect 1438 451 1444 452
rect 1438 450 1439 451
rect 1412 448 1439 450
rect 1412 447 1413 448
rect 1407 446 1413 447
rect 1438 447 1439 448
rect 1443 447 1444 451
rect 1471 451 1477 452
rect 1438 446 1444 447
rect 1446 447 1452 448
rect 1382 442 1388 443
rect 1446 443 1447 447
rect 1451 443 1452 447
rect 1471 447 1472 451
rect 1476 450 1477 451
rect 1526 451 1532 452
rect 1526 450 1527 451
rect 1476 448 1527 450
rect 1476 447 1477 448
rect 1471 446 1477 447
rect 1526 447 1527 448
rect 1531 447 1532 451
rect 1559 451 1565 452
rect 1526 446 1532 447
rect 1534 447 1540 448
rect 1446 442 1452 443
rect 1534 443 1535 447
rect 1539 443 1540 447
rect 1559 447 1560 451
rect 1564 450 1565 451
rect 1606 451 1612 452
rect 1606 450 1607 451
rect 1564 448 1607 450
rect 1564 447 1565 448
rect 1559 446 1565 447
rect 1606 447 1607 448
rect 1611 447 1612 451
rect 1655 451 1661 452
rect 1606 446 1612 447
rect 1630 447 1636 448
rect 1534 442 1540 443
rect 1630 443 1631 447
rect 1635 443 1636 447
rect 1655 447 1656 451
rect 1660 450 1661 451
rect 1726 451 1732 452
rect 1726 450 1727 451
rect 1660 448 1727 450
rect 1660 447 1661 448
rect 1655 446 1661 447
rect 1726 447 1727 448
rect 1731 447 1732 451
rect 1758 451 1765 452
rect 1726 446 1732 447
rect 1734 447 1740 448
rect 1630 442 1636 443
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1758 447 1759 451
rect 1764 447 1765 451
rect 1855 451 1861 452
rect 1758 446 1765 447
rect 1830 447 1836 448
rect 1734 442 1740 443
rect 1830 443 1831 447
rect 1835 443 1836 447
rect 1855 447 1856 451
rect 1860 450 1861 451
rect 1910 451 1916 452
rect 1910 450 1911 451
rect 1860 448 1911 450
rect 1860 447 1861 448
rect 1855 446 1861 447
rect 1910 447 1911 448
rect 1915 447 1916 451
rect 1943 451 1949 452
rect 1910 446 1916 447
rect 1918 447 1924 448
rect 1830 442 1836 443
rect 1918 443 1919 447
rect 1923 443 1924 447
rect 1943 447 1944 451
rect 1948 450 1949 451
rect 1978 451 1984 452
rect 1978 450 1979 451
rect 1948 448 1979 450
rect 1948 447 1949 448
rect 1943 446 1949 447
rect 1978 447 1979 448
rect 1983 447 1984 451
rect 2023 449 2024 453
rect 2028 452 2039 453
rect 2028 449 2029 452
rect 2038 451 2039 452
rect 2043 451 2044 455
rect 2038 450 2044 451
rect 2095 451 2101 452
rect 2023 448 2029 449
rect 1978 446 1984 447
rect 1998 447 2004 448
rect 1918 442 1924 443
rect 1998 443 1999 447
rect 2003 443 2004 447
rect 1998 442 2004 443
rect 2070 447 2076 448
rect 2070 443 2071 447
rect 2075 443 2076 447
rect 2095 447 2096 451
rect 2100 450 2101 451
rect 2126 451 2132 452
rect 2126 450 2127 451
rect 2100 448 2127 450
rect 2100 447 2101 448
rect 2095 446 2101 447
rect 2126 447 2127 448
rect 2131 447 2132 451
rect 2159 451 2165 452
rect 2126 446 2132 447
rect 2134 447 2140 448
rect 2070 442 2076 443
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2159 447 2160 451
rect 2164 450 2165 451
rect 2190 451 2196 452
rect 2190 450 2191 451
rect 2164 448 2191 450
rect 2164 447 2165 448
rect 2159 446 2165 447
rect 2190 447 2191 448
rect 2195 447 2196 451
rect 2223 451 2229 452
rect 2190 446 2196 447
rect 2198 447 2204 448
rect 2134 442 2140 443
rect 2198 443 2199 447
rect 2203 443 2204 447
rect 2223 447 2224 451
rect 2228 450 2229 451
rect 2246 451 2252 452
rect 2246 450 2247 451
rect 2228 448 2247 450
rect 2228 447 2229 448
rect 2223 446 2229 447
rect 2246 447 2247 448
rect 2251 447 2252 451
rect 2279 451 2285 452
rect 2246 446 2252 447
rect 2254 447 2260 448
rect 2198 442 2204 443
rect 2254 443 2255 447
rect 2259 443 2260 447
rect 2279 447 2280 451
rect 2284 450 2285 451
rect 2310 451 2316 452
rect 2310 450 2311 451
rect 2284 448 2311 450
rect 2284 447 2285 448
rect 2279 446 2285 447
rect 2310 447 2311 448
rect 2315 447 2316 451
rect 2343 451 2352 452
rect 2310 446 2316 447
rect 2318 447 2324 448
rect 2254 442 2260 443
rect 2318 443 2319 447
rect 2323 443 2324 447
rect 2343 447 2344 451
rect 2351 447 2352 451
rect 2382 451 2389 452
rect 2343 446 2352 447
rect 2358 447 2364 448
rect 2318 442 2324 443
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2382 447 2383 451
rect 2388 447 2389 451
rect 2382 446 2389 447
rect 2358 442 2364 443
rect 110 440 116 441
rect 110 436 111 440
rect 115 436 116 440
rect 1238 440 1244 441
rect 1238 436 1239 440
rect 1243 436 1244 440
rect 110 435 116 436
rect 262 435 269 436
rect 262 431 263 435
rect 268 431 269 435
rect 262 430 269 431
rect 294 435 300 436
rect 294 431 295 435
rect 299 434 300 435
rect 303 435 309 436
rect 303 434 304 435
rect 299 432 304 434
rect 299 431 300 432
rect 294 430 300 431
rect 303 431 304 432
rect 308 431 309 435
rect 303 430 309 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 434 324 435
rect 351 435 357 436
rect 351 434 352 435
rect 323 432 352 434
rect 323 431 324 432
rect 318 430 324 431
rect 351 431 352 432
rect 356 431 357 435
rect 351 430 357 431
rect 374 435 380 436
rect 374 431 375 435
rect 379 434 380 435
rect 407 435 413 436
rect 407 434 408 435
rect 379 432 408 434
rect 379 431 380 432
rect 374 430 380 431
rect 407 431 408 432
rect 412 431 413 435
rect 407 430 413 431
rect 463 435 469 436
rect 463 431 464 435
rect 468 434 469 435
rect 514 435 520 436
rect 514 434 515 435
rect 468 432 515 434
rect 468 431 469 432
rect 463 430 469 431
rect 514 431 515 432
rect 519 431 520 435
rect 514 430 520 431
rect 527 435 533 436
rect 527 431 528 435
rect 532 434 533 435
rect 574 435 580 436
rect 574 434 575 435
rect 532 432 575 434
rect 532 431 533 432
rect 527 430 533 431
rect 574 431 575 432
rect 579 431 580 435
rect 574 430 580 431
rect 582 435 588 436
rect 582 431 583 435
rect 587 434 588 435
rect 591 435 597 436
rect 591 434 592 435
rect 587 432 592 434
rect 587 431 588 432
rect 582 430 588 431
rect 591 431 592 432
rect 596 431 597 435
rect 591 430 597 431
rect 655 435 664 436
rect 655 431 656 435
rect 663 431 664 435
rect 655 430 664 431
rect 686 435 692 436
rect 686 431 687 435
rect 691 434 692 435
rect 719 435 725 436
rect 719 434 720 435
rect 691 432 720 434
rect 691 431 692 432
rect 686 430 692 431
rect 719 431 720 432
rect 724 431 725 435
rect 719 430 725 431
rect 750 435 756 436
rect 750 431 751 435
rect 755 434 756 435
rect 783 435 789 436
rect 783 434 784 435
rect 755 432 784 434
rect 755 431 756 432
rect 750 430 756 431
rect 783 431 784 432
rect 788 431 789 435
rect 783 430 789 431
rect 814 435 820 436
rect 814 431 815 435
rect 819 434 820 435
rect 847 435 853 436
rect 847 434 848 435
rect 819 432 848 434
rect 819 431 820 432
rect 814 430 820 431
rect 847 431 848 432
rect 852 431 853 435
rect 847 430 853 431
rect 878 435 884 436
rect 878 431 879 435
rect 883 434 884 435
rect 911 435 917 436
rect 911 434 912 435
rect 883 432 912 434
rect 883 431 884 432
rect 878 430 884 431
rect 911 431 912 432
rect 916 431 917 435
rect 911 430 917 431
rect 975 435 981 436
rect 975 431 976 435
rect 980 434 981 435
rect 1026 435 1032 436
rect 1026 434 1027 435
rect 980 432 1027 434
rect 980 431 981 432
rect 975 430 981 431
rect 1026 431 1027 432
rect 1031 431 1032 435
rect 1026 430 1032 431
rect 1039 435 1045 436
rect 1039 431 1040 435
rect 1044 434 1045 435
rect 1054 435 1060 436
rect 1238 435 1244 436
rect 1054 434 1055 435
rect 1044 432 1055 434
rect 1044 431 1045 432
rect 1039 430 1045 431
rect 1054 431 1055 432
rect 1059 431 1060 435
rect 1054 430 1060 431
rect 2346 427 2352 428
rect 1278 424 1284 425
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 2346 423 2347 427
rect 2351 426 2352 427
rect 2351 424 2387 426
rect 2351 423 2352 424
rect 2346 422 2352 423
rect 2385 420 2387 424
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 1278 419 1284 420
rect 1327 419 1333 420
rect 1238 418 1244 419
rect 238 416 244 417
rect 238 412 239 416
rect 243 412 244 416
rect 238 411 244 412
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 382 416 388 417
rect 382 412 383 416
rect 387 412 388 416
rect 382 411 388 412
rect 438 416 444 417
rect 438 412 439 416
rect 443 412 444 416
rect 438 411 444 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 566 416 572 417
rect 566 412 567 416
rect 571 412 572 416
rect 566 411 572 412
rect 630 416 636 417
rect 630 412 631 416
rect 635 412 636 416
rect 630 411 636 412
rect 694 416 700 417
rect 694 412 695 416
rect 699 412 700 416
rect 694 411 700 412
rect 758 416 764 417
rect 758 412 759 416
rect 763 412 764 416
rect 758 411 764 412
rect 822 416 828 417
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 886 416 892 417
rect 886 412 887 416
rect 891 412 892 416
rect 886 411 892 412
rect 950 416 956 417
rect 950 412 951 416
rect 955 412 956 416
rect 950 411 956 412
rect 1014 416 1020 417
rect 1014 412 1015 416
rect 1019 412 1020 416
rect 1327 415 1328 419
rect 1332 418 1333 419
rect 1350 419 1356 420
rect 1350 418 1351 419
rect 1332 416 1351 418
rect 1332 415 1333 416
rect 1327 414 1333 415
rect 1350 415 1351 416
rect 1355 415 1356 419
rect 1350 414 1356 415
rect 1358 419 1364 420
rect 1358 415 1359 419
rect 1363 418 1364 419
rect 1367 419 1373 420
rect 1367 418 1368 419
rect 1363 416 1368 418
rect 1363 415 1364 416
rect 1358 414 1364 415
rect 1367 415 1368 416
rect 1372 415 1373 419
rect 1367 414 1373 415
rect 1398 419 1404 420
rect 1398 415 1399 419
rect 1403 418 1404 419
rect 1407 419 1413 420
rect 1407 418 1408 419
rect 1403 416 1408 418
rect 1403 415 1404 416
rect 1398 414 1404 415
rect 1407 415 1408 416
rect 1412 415 1413 419
rect 1407 414 1413 415
rect 1438 419 1444 420
rect 1438 415 1439 419
rect 1443 418 1444 419
rect 1471 419 1477 420
rect 1471 418 1472 419
rect 1443 416 1472 418
rect 1443 415 1444 416
rect 1438 414 1444 415
rect 1471 415 1472 416
rect 1476 415 1477 419
rect 1471 414 1477 415
rect 1526 419 1532 420
rect 1526 415 1527 419
rect 1531 418 1532 419
rect 1559 419 1565 420
rect 1559 418 1560 419
rect 1531 416 1560 418
rect 1531 415 1532 416
rect 1526 414 1532 415
rect 1559 415 1560 416
rect 1564 415 1565 419
rect 1559 414 1565 415
rect 1606 419 1612 420
rect 1606 415 1607 419
rect 1611 418 1612 419
rect 1655 419 1661 420
rect 1655 418 1656 419
rect 1611 416 1656 418
rect 1611 415 1612 416
rect 1606 414 1612 415
rect 1655 415 1656 416
rect 1660 415 1661 419
rect 1655 414 1661 415
rect 1726 419 1732 420
rect 1726 415 1727 419
rect 1731 418 1732 419
rect 1759 419 1765 420
rect 1759 418 1760 419
rect 1731 416 1760 418
rect 1731 415 1732 416
rect 1726 414 1732 415
rect 1759 415 1760 416
rect 1764 415 1765 419
rect 1759 414 1765 415
rect 1854 419 1861 420
rect 1854 415 1855 419
rect 1860 415 1861 419
rect 1854 414 1861 415
rect 1943 419 1949 420
rect 1943 415 1944 419
rect 1948 418 1949 419
rect 1978 419 1984 420
rect 1948 416 1974 418
rect 1948 415 1949 416
rect 1943 414 1949 415
rect 1014 411 1020 412
rect 1972 410 1974 416
rect 1978 415 1979 419
rect 1983 418 1984 419
rect 2023 419 2029 420
rect 2023 418 2024 419
rect 1983 416 2024 418
rect 1983 415 1984 416
rect 1978 414 1984 415
rect 2023 415 2024 416
rect 2028 415 2029 419
rect 2023 414 2029 415
rect 2095 419 2101 420
rect 2095 415 2096 419
rect 2100 418 2101 419
rect 2110 419 2116 420
rect 2110 418 2111 419
rect 2100 416 2111 418
rect 2100 415 2101 416
rect 2095 414 2101 415
rect 2110 415 2111 416
rect 2115 415 2116 419
rect 2110 414 2116 415
rect 2126 419 2132 420
rect 2126 415 2127 419
rect 2131 418 2132 419
rect 2159 419 2165 420
rect 2159 418 2160 419
rect 2131 416 2160 418
rect 2131 415 2132 416
rect 2126 414 2132 415
rect 2159 415 2160 416
rect 2164 415 2165 419
rect 2159 414 2165 415
rect 2190 419 2196 420
rect 2190 415 2191 419
rect 2195 418 2196 419
rect 2223 419 2229 420
rect 2223 418 2224 419
rect 2195 416 2224 418
rect 2195 415 2196 416
rect 2190 414 2196 415
rect 2223 415 2224 416
rect 2228 415 2229 419
rect 2223 414 2229 415
rect 2246 419 2252 420
rect 2246 415 2247 419
rect 2251 418 2252 419
rect 2279 419 2285 420
rect 2279 418 2280 419
rect 2251 416 2280 418
rect 2251 415 2252 416
rect 2246 414 2252 415
rect 2279 415 2280 416
rect 2284 415 2285 419
rect 2279 414 2285 415
rect 2343 419 2352 420
rect 2343 415 2344 419
rect 2351 415 2352 419
rect 2343 414 2352 415
rect 2383 419 2389 420
rect 2406 419 2412 420
rect 2383 415 2384 419
rect 2388 415 2389 419
rect 2383 414 2389 415
rect 2098 411 2104 412
rect 2098 410 2099 411
rect 1972 408 2099 410
rect 1278 407 1284 408
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 2098 407 2099 408
rect 2103 407 2104 411
rect 2098 406 2104 407
rect 2406 407 2412 408
rect 1278 402 1284 403
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 142 400 148 401
rect 142 396 143 400
rect 147 396 148 400
rect 142 395 148 396
rect 182 400 188 401
rect 182 396 183 400
rect 187 396 188 400
rect 182 395 188 396
rect 222 400 228 401
rect 222 396 223 400
rect 227 396 228 400
rect 222 395 228 396
rect 270 400 276 401
rect 270 396 271 400
rect 275 396 276 400
rect 270 395 276 396
rect 334 400 340 401
rect 334 396 335 400
rect 339 396 340 400
rect 334 395 340 396
rect 398 400 404 401
rect 398 396 399 400
rect 403 396 404 400
rect 398 395 404 396
rect 470 400 476 401
rect 470 396 471 400
rect 475 396 476 400
rect 470 395 476 396
rect 542 400 548 401
rect 542 396 543 400
rect 547 396 548 400
rect 542 395 548 396
rect 614 400 620 401
rect 614 396 615 400
rect 619 396 620 400
rect 614 395 620 396
rect 686 400 692 401
rect 686 396 687 400
rect 691 396 692 400
rect 686 395 692 396
rect 750 400 756 401
rect 750 396 751 400
rect 755 396 756 400
rect 750 395 756 396
rect 806 400 812 401
rect 806 396 807 400
rect 811 396 812 400
rect 806 395 812 396
rect 862 400 868 401
rect 862 396 863 400
rect 867 396 868 400
rect 862 395 868 396
rect 918 400 924 401
rect 918 396 919 400
rect 923 396 924 400
rect 918 395 924 396
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 1030 400 1036 401
rect 1030 396 1031 400
rect 1035 396 1036 400
rect 1030 395 1036 396
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1382 400 1388 401
rect 1382 396 1383 400
rect 1387 396 1388 400
rect 1382 395 1388 396
rect 1446 400 1452 401
rect 1446 396 1447 400
rect 1451 396 1452 400
rect 1446 395 1452 396
rect 1534 400 1540 401
rect 1534 396 1535 400
rect 1539 396 1540 400
rect 1534 395 1540 396
rect 1630 400 1636 401
rect 1630 396 1631 400
rect 1635 396 1636 400
rect 1630 395 1636 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1830 400 1836 401
rect 1830 396 1831 400
rect 1835 396 1836 400
rect 1830 395 1836 396
rect 1918 400 1924 401
rect 1918 396 1919 400
rect 1923 396 1924 400
rect 1918 395 1924 396
rect 1998 400 2004 401
rect 1998 396 1999 400
rect 2003 396 2004 400
rect 1998 395 2004 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2198 400 2204 401
rect 2198 396 2199 400
rect 2203 396 2204 400
rect 2198 395 2204 396
rect 2254 400 2260 401
rect 2254 396 2255 400
rect 2259 396 2260 400
rect 2254 395 2260 396
rect 2318 400 2324 401
rect 2318 396 2319 400
rect 2323 396 2324 400
rect 2318 395 2324 396
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 1238 393 1244 394
rect 1238 389 1239 393
rect 1243 389 1244 393
rect 1238 388 1244 389
rect 1358 388 1364 389
rect 406 387 412 388
rect 406 386 407 387
rect 352 384 407 386
rect 167 379 173 380
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 167 375 168 379
rect 172 378 173 379
rect 198 379 204 380
rect 198 378 199 379
rect 172 376 199 378
rect 172 375 173 376
rect 167 374 173 375
rect 198 375 199 376
rect 203 375 204 379
rect 198 374 204 375
rect 207 379 213 380
rect 207 375 208 379
rect 212 378 213 379
rect 238 379 244 380
rect 238 378 239 379
rect 212 376 239 378
rect 212 375 213 376
rect 207 374 213 375
rect 238 375 239 376
rect 243 375 244 379
rect 238 374 244 375
rect 247 379 253 380
rect 247 375 248 379
rect 252 378 253 379
rect 286 379 292 380
rect 286 378 287 379
rect 252 376 287 378
rect 252 375 253 376
rect 247 374 253 375
rect 286 375 287 376
rect 291 375 292 379
rect 286 374 292 375
rect 295 379 301 380
rect 295 375 296 379
rect 300 378 301 379
rect 352 378 354 384
rect 406 383 407 384
rect 411 383 412 387
rect 1358 384 1359 388
rect 1363 384 1364 388
rect 1358 383 1364 384
rect 1398 388 1404 389
rect 1398 384 1399 388
rect 1403 384 1404 388
rect 1398 383 1404 384
rect 1438 388 1444 389
rect 1438 384 1439 388
rect 1443 384 1444 388
rect 1438 383 1444 384
rect 1486 388 1492 389
rect 1486 384 1487 388
rect 1491 384 1492 388
rect 1486 383 1492 384
rect 1542 388 1548 389
rect 1542 384 1543 388
rect 1547 384 1548 388
rect 1542 383 1548 384
rect 1606 388 1612 389
rect 1606 384 1607 388
rect 1611 384 1612 388
rect 1606 383 1612 384
rect 1678 388 1684 389
rect 1678 384 1679 388
rect 1683 384 1684 388
rect 1678 383 1684 384
rect 1758 388 1764 389
rect 1758 384 1759 388
rect 1763 384 1764 388
rect 1758 383 1764 384
rect 1838 388 1844 389
rect 1838 384 1839 388
rect 1843 384 1844 388
rect 1838 383 1844 384
rect 1918 388 1924 389
rect 1918 384 1919 388
rect 1923 384 1924 388
rect 1918 383 1924 384
rect 1998 388 2004 389
rect 1998 384 1999 388
rect 2003 384 2004 388
rect 1998 383 2004 384
rect 2078 388 2084 389
rect 2078 384 2079 388
rect 2083 384 2084 388
rect 2078 383 2084 384
rect 2158 388 2164 389
rect 2158 384 2159 388
rect 2163 384 2164 388
rect 2158 383 2164 384
rect 2246 388 2252 389
rect 2246 384 2247 388
rect 2251 384 2252 388
rect 2246 383 2252 384
rect 2334 388 2340 389
rect 2334 384 2335 388
rect 2339 384 2340 388
rect 2334 383 2340 384
rect 406 382 412 383
rect 1278 381 1284 382
rect 300 376 354 378
rect 359 379 365 380
rect 300 375 301 376
rect 295 374 301 375
rect 359 375 360 379
rect 364 375 365 379
rect 359 374 365 375
rect 367 379 373 380
rect 367 375 368 379
rect 372 378 373 379
rect 423 379 429 380
rect 423 378 424 379
rect 372 376 424 378
rect 372 375 373 376
rect 367 374 373 375
rect 423 375 424 376
rect 428 375 429 379
rect 423 374 429 375
rect 431 379 437 380
rect 431 375 432 379
rect 436 378 437 379
rect 495 379 501 380
rect 495 378 496 379
rect 436 376 496 378
rect 436 375 437 376
rect 431 374 437 375
rect 495 375 496 376
rect 500 375 501 379
rect 495 374 501 375
rect 506 379 512 380
rect 506 375 507 379
rect 511 378 512 379
rect 567 379 573 380
rect 567 378 568 379
rect 511 376 568 378
rect 511 375 512 376
rect 506 374 512 375
rect 567 375 568 376
rect 572 375 573 379
rect 567 374 573 375
rect 639 379 645 380
rect 639 375 640 379
rect 644 378 645 379
rect 702 379 708 380
rect 702 378 703 379
rect 644 376 703 378
rect 644 375 645 376
rect 639 374 645 375
rect 702 375 703 376
rect 707 375 708 379
rect 702 374 708 375
rect 711 379 717 380
rect 711 375 712 379
rect 716 378 717 379
rect 766 379 772 380
rect 766 378 767 379
rect 716 376 767 378
rect 716 375 717 376
rect 711 374 717 375
rect 766 375 767 376
rect 771 375 772 379
rect 766 374 772 375
rect 775 379 781 380
rect 775 375 776 379
rect 780 378 781 379
rect 822 379 828 380
rect 822 378 823 379
rect 780 376 823 378
rect 780 375 781 376
rect 775 374 781 375
rect 822 375 823 376
rect 827 375 828 379
rect 822 374 828 375
rect 831 379 837 380
rect 831 375 832 379
rect 836 378 837 379
rect 878 379 884 380
rect 878 378 879 379
rect 836 376 879 378
rect 836 375 837 376
rect 831 374 837 375
rect 878 375 879 376
rect 883 375 884 379
rect 878 374 884 375
rect 887 379 893 380
rect 887 375 888 379
rect 892 378 893 379
rect 898 379 904 380
rect 898 378 899 379
rect 892 376 899 378
rect 892 375 893 376
rect 887 374 893 375
rect 898 375 899 376
rect 903 375 904 379
rect 898 374 904 375
rect 906 379 912 380
rect 906 375 907 379
rect 911 378 912 379
rect 943 379 949 380
rect 943 378 944 379
rect 911 376 944 378
rect 911 375 912 376
rect 906 374 912 375
rect 943 375 944 376
rect 948 375 949 379
rect 943 374 949 375
rect 951 379 957 380
rect 951 375 952 379
rect 956 378 957 379
rect 999 379 1005 380
rect 999 378 1000 379
rect 956 376 1000 378
rect 956 375 957 376
rect 951 374 957 375
rect 999 375 1000 376
rect 1004 375 1005 379
rect 999 374 1005 375
rect 1007 379 1013 380
rect 1007 375 1008 379
rect 1012 378 1013 379
rect 1055 379 1061 380
rect 1055 378 1056 379
rect 1012 376 1056 378
rect 1012 375 1013 376
rect 1007 374 1013 375
rect 1055 375 1056 376
rect 1060 375 1061 379
rect 1278 377 1279 381
rect 1283 377 1284 381
rect 1055 374 1061 375
rect 1238 376 1244 377
rect 1278 376 1284 377
rect 2406 381 2412 382
rect 2406 377 2407 381
rect 2411 377 2412 381
rect 2406 376 2412 377
rect 110 371 116 372
rect 360 370 362 374
rect 1238 372 1239 376
rect 1243 372 1244 376
rect 462 371 468 372
rect 1238 371 1244 372
rect 462 370 463 371
rect 360 368 463 370
rect 462 367 463 368
rect 467 367 468 371
rect 462 366 468 367
rect 1383 367 1389 368
rect 1278 364 1284 365
rect 1278 360 1279 364
rect 1283 360 1284 364
rect 1383 363 1384 367
rect 1388 366 1389 367
rect 1414 367 1420 368
rect 1414 366 1415 367
rect 1388 364 1415 366
rect 1388 363 1389 364
rect 1383 362 1389 363
rect 1414 363 1415 364
rect 1419 363 1420 367
rect 1414 362 1420 363
rect 1423 367 1429 368
rect 1423 363 1424 367
rect 1428 366 1429 367
rect 1454 367 1460 368
rect 1454 366 1455 367
rect 1428 364 1455 366
rect 1428 363 1429 364
rect 1423 362 1429 363
rect 1454 363 1455 364
rect 1459 363 1460 367
rect 1454 362 1460 363
rect 1463 367 1469 368
rect 1463 363 1464 367
rect 1468 366 1469 367
rect 1502 367 1508 368
rect 1502 366 1503 367
rect 1468 364 1503 366
rect 1468 363 1469 364
rect 1463 362 1469 363
rect 1502 363 1503 364
rect 1507 363 1508 367
rect 1502 362 1508 363
rect 1511 367 1517 368
rect 1511 363 1512 367
rect 1516 366 1517 367
rect 1558 367 1564 368
rect 1558 366 1559 367
rect 1516 364 1559 366
rect 1516 363 1517 364
rect 1511 362 1517 363
rect 1558 363 1559 364
rect 1563 363 1564 367
rect 1558 362 1564 363
rect 1567 367 1573 368
rect 1567 363 1568 367
rect 1572 366 1573 367
rect 1614 367 1620 368
rect 1572 364 1610 366
rect 1572 363 1573 364
rect 1567 362 1573 363
rect 1278 359 1284 360
rect 1608 358 1610 364
rect 1614 363 1615 367
rect 1619 366 1620 367
rect 1631 367 1637 368
rect 1631 366 1632 367
rect 1619 364 1632 366
rect 1619 363 1620 364
rect 1614 362 1620 363
rect 1631 363 1632 364
rect 1636 363 1637 367
rect 1631 362 1637 363
rect 1639 367 1645 368
rect 1639 363 1640 367
rect 1644 366 1645 367
rect 1703 367 1709 368
rect 1703 366 1704 367
rect 1644 364 1704 366
rect 1644 363 1645 364
rect 1639 362 1645 363
rect 1703 363 1704 364
rect 1708 363 1709 367
rect 1703 362 1709 363
rect 1783 367 1789 368
rect 1783 363 1784 367
rect 1788 366 1789 367
rect 1854 367 1860 368
rect 1854 366 1855 367
rect 1788 364 1855 366
rect 1788 363 1789 364
rect 1783 362 1789 363
rect 1854 363 1855 364
rect 1859 363 1860 367
rect 1854 362 1860 363
rect 1863 367 1869 368
rect 1863 363 1864 367
rect 1868 363 1869 367
rect 1863 362 1869 363
rect 1910 367 1916 368
rect 1910 363 1911 367
rect 1915 366 1916 367
rect 1943 367 1949 368
rect 1943 366 1944 367
rect 1915 364 1944 366
rect 1915 363 1916 364
rect 1910 362 1916 363
rect 1943 363 1944 364
rect 1948 363 1949 367
rect 1943 362 1949 363
rect 1951 367 1957 368
rect 1951 363 1952 367
rect 1956 366 1957 367
rect 2023 367 2029 368
rect 2023 366 2024 367
rect 1956 364 2024 366
rect 1956 363 1957 364
rect 1951 362 1957 363
rect 2023 363 2024 364
rect 2028 363 2029 367
rect 2023 362 2029 363
rect 2103 367 2109 368
rect 2103 363 2104 367
rect 2108 366 2109 367
rect 2174 367 2180 368
rect 2174 366 2175 367
rect 2108 364 2175 366
rect 2108 363 2109 364
rect 2103 362 2109 363
rect 2174 363 2175 364
rect 2179 363 2180 367
rect 2174 362 2180 363
rect 2183 367 2189 368
rect 2183 363 2184 367
rect 2188 366 2189 367
rect 2218 367 2224 368
rect 2218 366 2219 367
rect 2188 364 2219 366
rect 2188 363 2189 364
rect 2183 362 2189 363
rect 2218 363 2219 364
rect 2223 363 2224 367
rect 2218 362 2224 363
rect 2226 367 2232 368
rect 2226 363 2227 367
rect 2231 366 2232 367
rect 2271 367 2277 368
rect 2271 366 2272 367
rect 2231 364 2272 366
rect 2231 363 2232 364
rect 2226 362 2232 363
rect 2271 363 2272 364
rect 2276 363 2277 367
rect 2271 362 2277 363
rect 2310 367 2316 368
rect 2310 363 2311 367
rect 2315 366 2316 367
rect 2359 367 2365 368
rect 2359 366 2360 367
rect 2315 364 2360 366
rect 2315 363 2316 364
rect 2310 362 2316 363
rect 2359 363 2360 364
rect 2364 363 2365 367
rect 2359 362 2365 363
rect 2406 364 2412 365
rect 1702 359 1708 360
rect 1702 358 1703 359
rect 1608 356 1703 358
rect 1702 355 1703 356
rect 1707 355 1708 359
rect 1865 358 1867 362
rect 2406 360 2407 364
rect 2411 360 2412 364
rect 2022 359 2028 360
rect 2406 359 2412 360
rect 2022 358 2023 359
rect 1865 356 2023 358
rect 1702 354 1708 355
rect 2022 355 2023 356
rect 2027 355 2028 359
rect 2022 354 2028 355
rect 142 353 148 354
rect 142 349 143 353
rect 147 349 148 353
rect 142 348 148 349
rect 182 353 188 354
rect 182 349 183 353
rect 187 349 188 353
rect 182 348 188 349
rect 222 353 228 354
rect 222 349 223 353
rect 227 349 228 353
rect 222 348 228 349
rect 270 353 276 354
rect 270 349 271 353
rect 275 349 276 353
rect 270 348 276 349
rect 334 353 340 354
rect 334 349 335 353
rect 339 349 340 353
rect 334 348 340 349
rect 398 353 404 354
rect 398 349 399 353
rect 403 349 404 353
rect 398 348 404 349
rect 470 353 476 354
rect 470 349 471 353
rect 475 349 476 353
rect 470 348 476 349
rect 542 353 548 354
rect 542 349 543 353
rect 547 349 548 353
rect 614 353 620 354
rect 582 351 588 352
rect 582 350 583 351
rect 542 348 548 349
rect 567 349 583 350
rect 167 347 173 348
rect 167 343 168 347
rect 172 346 173 347
rect 198 347 204 348
rect 198 346 199 347
rect 172 344 199 346
rect 172 343 173 344
rect 167 342 173 343
rect 198 343 199 344
rect 203 343 204 347
rect 198 342 204 343
rect 206 347 213 348
rect 206 343 207 347
rect 212 343 213 347
rect 206 342 213 343
rect 238 347 244 348
rect 238 343 239 347
rect 243 346 244 347
rect 247 347 253 348
rect 247 346 248 347
rect 243 344 248 346
rect 243 343 244 344
rect 238 342 244 343
rect 247 343 248 344
rect 252 343 253 347
rect 247 342 253 343
rect 286 347 292 348
rect 286 343 287 347
rect 291 346 292 347
rect 295 347 301 348
rect 295 346 296 347
rect 291 344 296 346
rect 291 343 292 344
rect 286 342 292 343
rect 295 343 296 344
rect 300 343 301 347
rect 295 342 301 343
rect 359 347 365 348
rect 359 343 360 347
rect 364 346 365 347
rect 367 347 373 348
rect 367 346 368 347
rect 364 344 368 346
rect 364 343 365 344
rect 359 342 365 343
rect 367 343 368 344
rect 372 343 373 347
rect 367 342 373 343
rect 423 347 429 348
rect 423 343 424 347
rect 428 346 429 347
rect 431 347 437 348
rect 431 346 432 347
rect 428 344 432 346
rect 428 343 429 344
rect 423 342 429 343
rect 431 343 432 344
rect 436 343 437 347
rect 431 342 437 343
rect 495 347 501 348
rect 495 343 496 347
rect 500 346 501 347
rect 506 347 512 348
rect 506 346 507 347
rect 500 344 507 346
rect 500 343 501 344
rect 495 342 501 343
rect 506 343 507 344
rect 511 343 512 347
rect 567 345 568 349
rect 572 348 583 349
rect 572 345 573 348
rect 582 347 583 348
rect 587 347 588 351
rect 614 349 615 353
rect 619 349 620 353
rect 614 348 620 349
rect 686 353 692 354
rect 686 349 687 353
rect 691 349 692 353
rect 686 348 692 349
rect 750 353 756 354
rect 750 349 751 353
rect 755 349 756 353
rect 750 348 756 349
rect 806 353 812 354
rect 806 349 807 353
rect 811 349 812 353
rect 806 348 812 349
rect 862 353 868 354
rect 862 349 863 353
rect 867 349 868 353
rect 862 348 868 349
rect 918 353 924 354
rect 918 349 919 353
rect 923 349 924 353
rect 918 348 924 349
rect 974 353 980 354
rect 974 349 975 353
rect 979 349 980 353
rect 974 348 980 349
rect 1030 353 1036 354
rect 1030 349 1031 353
rect 1035 349 1036 353
rect 1030 348 1036 349
rect 582 346 588 347
rect 630 347 636 348
rect 567 344 573 345
rect 506 342 512 343
rect 630 343 631 347
rect 635 346 636 347
rect 639 347 645 348
rect 639 346 640 347
rect 635 344 640 346
rect 635 343 636 344
rect 630 342 636 343
rect 639 343 640 344
rect 644 343 645 347
rect 639 342 645 343
rect 702 347 708 348
rect 702 343 703 347
rect 707 346 708 347
rect 711 347 717 348
rect 711 346 712 347
rect 707 344 712 346
rect 707 343 708 344
rect 702 342 708 343
rect 711 343 712 344
rect 716 343 717 347
rect 711 342 717 343
rect 766 347 772 348
rect 766 343 767 347
rect 771 346 772 347
rect 775 347 781 348
rect 775 346 776 347
rect 771 344 776 346
rect 771 343 772 344
rect 766 342 772 343
rect 775 343 776 344
rect 780 343 781 347
rect 775 342 781 343
rect 822 347 828 348
rect 822 343 823 347
rect 827 346 828 347
rect 831 347 837 348
rect 831 346 832 347
rect 827 344 832 346
rect 827 343 828 344
rect 822 342 828 343
rect 831 343 832 344
rect 836 343 837 347
rect 831 342 837 343
rect 878 347 884 348
rect 878 343 879 347
rect 883 346 884 347
rect 887 347 893 348
rect 887 346 888 347
rect 883 344 888 346
rect 883 343 884 344
rect 878 342 884 343
rect 887 343 888 344
rect 892 343 893 347
rect 887 342 893 343
rect 943 347 949 348
rect 943 343 944 347
rect 948 346 949 347
rect 951 347 957 348
rect 951 346 952 347
rect 948 344 952 346
rect 948 343 949 344
rect 943 342 949 343
rect 951 343 952 344
rect 956 343 957 347
rect 951 342 957 343
rect 999 347 1005 348
rect 999 343 1000 347
rect 1004 346 1005 347
rect 1007 347 1013 348
rect 1007 346 1008 347
rect 1004 344 1008 346
rect 1004 343 1005 344
rect 999 342 1005 343
rect 1007 343 1008 344
rect 1012 343 1013 347
rect 1007 342 1013 343
rect 1054 347 1061 348
rect 1054 343 1055 347
rect 1060 343 1061 347
rect 1054 342 1061 343
rect 1358 341 1364 342
rect 1358 337 1359 341
rect 1363 337 1364 341
rect 1358 336 1364 337
rect 1398 341 1404 342
rect 1398 337 1399 341
rect 1403 337 1404 341
rect 1398 336 1404 337
rect 1438 341 1444 342
rect 1438 337 1439 341
rect 1443 337 1444 341
rect 1438 336 1444 337
rect 1486 341 1492 342
rect 1486 337 1487 341
rect 1491 337 1492 341
rect 1486 336 1492 337
rect 1542 341 1548 342
rect 1542 337 1543 341
rect 1547 337 1548 341
rect 1542 336 1548 337
rect 1606 341 1612 342
rect 1606 337 1607 341
rect 1611 337 1612 341
rect 1606 336 1612 337
rect 1678 341 1684 342
rect 1678 337 1679 341
rect 1683 337 1684 341
rect 1678 336 1684 337
rect 1758 341 1764 342
rect 1758 337 1759 341
rect 1763 337 1764 341
rect 1758 336 1764 337
rect 1838 341 1844 342
rect 1838 337 1839 341
rect 1843 337 1844 341
rect 1838 336 1844 337
rect 1918 341 1924 342
rect 1918 337 1919 341
rect 1923 337 1924 341
rect 1918 336 1924 337
rect 1998 341 2004 342
rect 1998 337 1999 341
rect 2003 337 2004 341
rect 1998 336 2004 337
rect 2078 341 2084 342
rect 2078 337 2079 341
rect 2083 337 2084 341
rect 2078 336 2084 337
rect 2158 341 2164 342
rect 2158 337 2159 341
rect 2163 337 2164 341
rect 2158 336 2164 337
rect 2246 341 2252 342
rect 2246 337 2247 341
rect 2251 337 2252 341
rect 2246 336 2252 337
rect 2334 341 2340 342
rect 2334 337 2335 341
rect 2339 337 2340 341
rect 2334 336 2340 337
rect 1350 335 1356 336
rect 1350 331 1351 335
rect 1355 334 1356 335
rect 1383 335 1389 336
rect 1383 334 1384 335
rect 1355 332 1384 334
rect 1355 331 1356 332
rect 1350 330 1356 331
rect 1383 331 1384 332
rect 1388 331 1389 335
rect 1383 330 1389 331
rect 1414 335 1420 336
rect 1414 331 1415 335
rect 1419 334 1420 335
rect 1423 335 1429 336
rect 1423 334 1424 335
rect 1419 332 1424 334
rect 1419 331 1420 332
rect 1414 330 1420 331
rect 1423 331 1424 332
rect 1428 331 1429 335
rect 1423 330 1429 331
rect 1454 335 1460 336
rect 1454 331 1455 335
rect 1459 334 1460 335
rect 1463 335 1469 336
rect 1463 334 1464 335
rect 1459 332 1464 334
rect 1459 331 1460 332
rect 1454 330 1460 331
rect 1463 331 1464 332
rect 1468 331 1469 335
rect 1463 330 1469 331
rect 1502 335 1508 336
rect 1502 331 1503 335
rect 1507 334 1508 335
rect 1511 335 1517 336
rect 1511 334 1512 335
rect 1507 332 1512 334
rect 1507 331 1508 332
rect 1502 330 1508 331
rect 1511 331 1512 332
rect 1516 331 1517 335
rect 1511 330 1517 331
rect 1558 335 1564 336
rect 1558 331 1559 335
rect 1563 334 1564 335
rect 1567 335 1573 336
rect 1567 334 1568 335
rect 1563 332 1568 334
rect 1563 331 1564 332
rect 1558 330 1564 331
rect 1567 331 1568 332
rect 1572 331 1573 335
rect 1567 330 1573 331
rect 1631 335 1637 336
rect 1631 331 1632 335
rect 1636 334 1637 335
rect 1639 335 1645 336
rect 1639 334 1640 335
rect 1636 332 1640 334
rect 1636 331 1637 332
rect 1631 330 1637 331
rect 1639 331 1640 332
rect 1644 331 1645 335
rect 1639 330 1645 331
rect 1702 335 1709 336
rect 1702 331 1703 335
rect 1708 331 1709 335
rect 1702 330 1709 331
rect 1783 335 1789 336
rect 1783 331 1784 335
rect 1788 334 1789 335
rect 1846 335 1852 336
rect 1846 334 1847 335
rect 1788 332 1847 334
rect 1788 331 1789 332
rect 1783 330 1789 331
rect 1846 331 1847 332
rect 1851 331 1852 335
rect 1846 330 1852 331
rect 1854 335 1860 336
rect 1854 331 1855 335
rect 1859 334 1860 335
rect 1863 335 1869 336
rect 1863 334 1864 335
rect 1859 332 1864 334
rect 1859 331 1860 332
rect 1854 330 1860 331
rect 1863 331 1864 332
rect 1868 331 1869 335
rect 1863 330 1869 331
rect 1943 335 1949 336
rect 1943 331 1944 335
rect 1948 334 1949 335
rect 1951 335 1957 336
rect 1951 334 1952 335
rect 1948 332 1952 334
rect 1948 331 1949 332
rect 1943 330 1949 331
rect 1951 331 1952 332
rect 1956 331 1957 335
rect 1951 330 1957 331
rect 2022 335 2029 336
rect 2022 331 2023 335
rect 2028 331 2029 335
rect 2022 330 2029 331
rect 2098 335 2109 336
rect 2098 331 2099 335
rect 2103 331 2104 335
rect 2108 331 2109 335
rect 2098 330 2109 331
rect 2174 335 2180 336
rect 2174 331 2175 335
rect 2179 334 2180 335
rect 2183 335 2189 336
rect 2183 334 2184 335
rect 2179 332 2184 334
rect 2179 331 2180 332
rect 2174 330 2180 331
rect 2183 331 2184 332
rect 2188 331 2189 335
rect 2183 330 2189 331
rect 2218 335 2224 336
rect 2218 331 2219 335
rect 2223 334 2224 335
rect 2271 335 2277 336
rect 2271 334 2272 335
rect 2223 332 2272 334
rect 2223 331 2224 332
rect 2218 330 2224 331
rect 2271 331 2272 332
rect 2276 331 2277 335
rect 2271 330 2277 331
rect 2346 335 2352 336
rect 2346 331 2347 335
rect 2351 334 2352 335
rect 2359 335 2365 336
rect 2359 334 2360 335
rect 2351 332 2360 334
rect 2351 331 2352 332
rect 2346 330 2352 331
rect 2359 331 2360 332
rect 2364 331 2365 335
rect 2359 330 2365 331
rect 230 323 236 324
rect 230 322 231 323
rect 201 320 231 322
rect 158 319 165 320
rect 134 315 140 316
rect 134 311 135 315
rect 139 311 140 315
rect 158 315 159 319
rect 164 315 165 319
rect 199 319 205 320
rect 158 314 165 315
rect 174 315 180 316
rect 134 310 140 311
rect 174 311 175 315
rect 179 311 180 315
rect 199 315 200 319
rect 204 315 205 319
rect 230 319 231 320
rect 235 319 236 323
rect 654 323 660 324
rect 654 322 655 323
rect 632 320 655 322
rect 230 318 236 319
rect 239 319 248 320
rect 199 314 205 315
rect 214 315 220 316
rect 174 310 180 311
rect 214 311 215 315
rect 219 311 220 315
rect 239 315 240 319
rect 247 315 248 319
rect 266 319 272 320
rect 239 314 248 315
rect 254 315 260 316
rect 214 310 220 311
rect 254 311 255 315
rect 259 311 260 315
rect 266 315 267 319
rect 271 318 272 319
rect 279 319 285 320
rect 279 318 280 319
rect 271 316 280 318
rect 271 315 272 316
rect 266 314 272 315
rect 279 315 280 316
rect 284 315 285 319
rect 319 319 328 320
rect 279 314 285 315
rect 294 315 300 316
rect 254 310 260 311
rect 294 311 295 315
rect 299 311 300 315
rect 319 315 320 319
rect 327 315 328 319
rect 359 319 365 320
rect 319 314 328 315
rect 334 315 340 316
rect 294 310 300 311
rect 334 311 335 315
rect 339 311 340 315
rect 359 315 360 319
rect 364 318 365 319
rect 382 319 388 320
rect 382 318 383 319
rect 364 316 383 318
rect 364 315 365 316
rect 359 314 365 315
rect 382 315 383 316
rect 387 315 388 319
rect 415 319 421 320
rect 382 314 388 315
rect 390 315 396 316
rect 334 310 340 311
rect 390 311 391 315
rect 395 311 396 315
rect 415 315 416 319
rect 420 318 421 319
rect 438 319 444 320
rect 438 318 439 319
rect 420 316 439 318
rect 420 315 421 316
rect 415 314 421 315
rect 438 315 439 316
rect 443 315 444 319
rect 462 319 468 320
rect 438 314 444 315
rect 446 315 452 316
rect 390 310 396 311
rect 446 311 447 315
rect 451 311 452 315
rect 462 315 463 319
rect 467 318 468 319
rect 471 319 477 320
rect 471 318 472 319
rect 467 316 472 318
rect 467 315 468 316
rect 462 314 468 315
rect 471 315 472 316
rect 476 315 477 319
rect 519 319 525 320
rect 471 314 477 315
rect 494 315 500 316
rect 446 310 452 311
rect 494 311 495 315
rect 499 311 500 315
rect 519 315 520 319
rect 524 318 525 319
rect 534 319 540 320
rect 534 318 535 319
rect 524 316 535 318
rect 524 315 525 316
rect 519 314 525 315
rect 534 315 535 316
rect 539 315 540 319
rect 567 319 573 320
rect 534 314 540 315
rect 542 315 548 316
rect 494 310 500 311
rect 542 311 543 315
rect 547 311 548 315
rect 567 315 568 319
rect 572 318 573 319
rect 615 319 621 320
rect 572 316 586 318
rect 572 315 573 316
rect 567 314 573 315
rect 542 310 548 311
rect 584 306 586 316
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 615 315 616 319
rect 620 318 621 319
rect 632 318 634 320
rect 654 319 655 320
rect 659 319 660 323
rect 654 318 660 319
rect 663 319 669 320
rect 620 316 634 318
rect 620 315 621 316
rect 615 314 621 315
rect 638 315 644 316
rect 590 310 596 311
rect 638 311 639 315
rect 643 311 644 315
rect 663 315 664 319
rect 668 318 669 319
rect 678 319 684 320
rect 678 318 679 319
rect 668 316 679 318
rect 668 315 669 316
rect 663 314 669 315
rect 678 315 679 316
rect 683 315 684 319
rect 711 319 717 320
rect 678 314 684 315
rect 686 315 692 316
rect 638 310 644 311
rect 686 311 687 315
rect 691 311 692 315
rect 711 315 712 319
rect 716 318 717 319
rect 726 319 732 320
rect 726 318 727 319
rect 716 316 727 318
rect 716 315 717 316
rect 711 314 717 315
rect 726 315 727 316
rect 731 315 732 319
rect 759 319 765 320
rect 726 314 732 315
rect 734 315 740 316
rect 686 310 692 311
rect 734 311 735 315
rect 739 311 740 315
rect 759 315 760 319
rect 764 318 765 319
rect 774 319 780 320
rect 774 318 775 319
rect 764 316 775 318
rect 764 315 765 316
rect 759 314 765 315
rect 774 315 775 316
rect 779 315 780 319
rect 794 319 800 320
rect 774 314 780 315
rect 782 315 788 316
rect 734 310 740 311
rect 782 311 783 315
rect 787 311 788 315
rect 794 315 795 319
rect 799 318 800 319
rect 807 319 813 320
rect 807 318 808 319
rect 799 316 808 318
rect 799 315 800 316
rect 794 314 800 315
rect 807 315 808 316
rect 812 315 813 319
rect 863 319 869 320
rect 807 314 813 315
rect 838 315 844 316
rect 782 310 788 311
rect 838 311 839 315
rect 843 311 844 315
rect 863 315 864 319
rect 868 318 869 319
rect 906 319 912 320
rect 906 318 907 319
rect 868 316 907 318
rect 868 315 869 316
rect 863 314 869 315
rect 906 315 907 316
rect 911 315 912 319
rect 906 314 912 315
rect 838 310 844 311
rect 1598 311 1604 312
rect 1598 310 1599 311
rect 1584 308 1599 310
rect 862 307 868 308
rect 862 306 863 307
rect 584 304 863 306
rect 862 303 863 304
rect 867 303 868 307
rect 1535 307 1544 308
rect 862 302 868 303
rect 1510 303 1516 304
rect 1510 299 1511 303
rect 1515 299 1516 303
rect 1535 303 1536 307
rect 1543 303 1544 307
rect 1575 307 1581 308
rect 1535 302 1544 303
rect 1550 303 1556 304
rect 1510 298 1516 299
rect 1550 299 1551 303
rect 1555 299 1556 303
rect 1575 303 1576 307
rect 1580 306 1581 307
rect 1584 306 1586 308
rect 1598 307 1599 308
rect 1603 307 1604 311
rect 1686 311 1692 312
rect 1686 310 1687 311
rect 1664 308 1687 310
rect 1598 306 1604 307
rect 1614 307 1621 308
rect 1580 304 1586 306
rect 1580 303 1581 304
rect 1575 302 1581 303
rect 1590 303 1596 304
rect 1550 298 1556 299
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1614 303 1615 307
rect 1620 303 1621 307
rect 1655 307 1661 308
rect 1614 302 1621 303
rect 1630 303 1636 304
rect 1590 298 1596 299
rect 1630 299 1631 303
rect 1635 299 1636 303
rect 1655 303 1656 307
rect 1660 306 1661 307
rect 1664 306 1666 308
rect 1686 307 1687 308
rect 1691 307 1692 311
rect 1766 311 1772 312
rect 1766 310 1767 311
rect 1744 308 1767 310
rect 1686 306 1692 307
rect 1695 307 1704 308
rect 1660 304 1666 306
rect 1660 303 1661 304
rect 1655 302 1661 303
rect 1670 303 1676 304
rect 1630 298 1636 299
rect 1670 299 1671 303
rect 1675 299 1676 303
rect 1695 303 1696 307
rect 1703 303 1704 307
rect 1735 307 1741 308
rect 1695 302 1704 303
rect 1710 303 1716 304
rect 1670 298 1676 299
rect 1710 299 1711 303
rect 1715 299 1716 303
rect 1735 303 1736 307
rect 1740 306 1741 307
rect 1744 306 1746 308
rect 1766 307 1767 308
rect 1771 307 1772 311
rect 1766 306 1772 307
rect 1775 307 1784 308
rect 1740 304 1746 306
rect 1740 303 1741 304
rect 1735 302 1741 303
rect 1750 303 1756 304
rect 1710 298 1716 299
rect 1750 299 1751 303
rect 1755 299 1756 303
rect 1775 303 1776 307
rect 1783 303 1784 307
rect 1815 307 1821 308
rect 1815 306 1816 307
rect 1800 304 1816 306
rect 1775 302 1784 303
rect 1790 303 1796 304
rect 1750 298 1756 299
rect 1790 299 1791 303
rect 1795 299 1796 303
rect 1790 298 1796 299
rect 266 295 272 296
rect 266 294 267 295
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 161 292 267 294
rect 161 288 163 292
rect 266 291 267 292
rect 271 291 272 295
rect 266 290 272 291
rect 322 295 328 296
rect 322 291 323 295
rect 327 294 328 295
rect 1543 295 1549 296
rect 327 292 363 294
rect 327 291 328 292
rect 322 290 328 291
rect 361 288 363 292
rect 1238 292 1244 293
rect 1238 288 1239 292
rect 1243 288 1244 292
rect 1543 291 1544 295
rect 1548 294 1549 295
rect 1800 294 1802 304
rect 1815 303 1816 304
rect 1820 303 1821 307
rect 1863 307 1869 308
rect 1815 302 1821 303
rect 1838 303 1844 304
rect 1838 299 1839 303
rect 1843 299 1844 303
rect 1863 303 1864 307
rect 1868 306 1869 307
rect 1894 307 1900 308
rect 1894 306 1895 307
rect 1868 304 1895 306
rect 1868 303 1869 304
rect 1863 302 1869 303
rect 1894 303 1895 304
rect 1899 303 1900 307
rect 1927 307 1933 308
rect 1894 302 1900 303
rect 1902 303 1908 304
rect 1838 298 1844 299
rect 1902 299 1903 303
rect 1907 299 1908 303
rect 1927 303 1928 307
rect 1932 306 1933 307
rect 1958 307 1964 308
rect 1958 306 1959 307
rect 1932 304 1959 306
rect 1932 303 1933 304
rect 1927 302 1933 303
rect 1958 303 1959 304
rect 1963 303 1964 307
rect 1991 307 1997 308
rect 1958 302 1964 303
rect 1966 303 1972 304
rect 1902 298 1908 299
rect 1966 299 1967 303
rect 1971 299 1972 303
rect 1991 303 1992 307
rect 1996 306 1997 307
rect 2026 307 2032 308
rect 2026 306 2027 307
rect 1996 304 2027 306
rect 1996 303 1997 304
rect 1991 302 1997 303
rect 2026 303 2027 304
rect 2031 303 2032 307
rect 2063 307 2069 308
rect 2026 302 2032 303
rect 2038 303 2044 304
rect 1966 298 1972 299
rect 2038 299 2039 303
rect 2043 299 2044 303
rect 2063 303 2064 307
rect 2068 306 2069 307
rect 2110 307 2116 308
rect 2110 306 2111 307
rect 2068 304 2111 306
rect 2068 303 2069 304
rect 2063 302 2069 303
rect 2110 303 2111 304
rect 2115 303 2116 307
rect 2130 307 2136 308
rect 2110 302 2116 303
rect 2118 303 2124 304
rect 2038 298 2044 299
rect 2118 299 2119 303
rect 2123 299 2124 303
rect 2130 303 2131 307
rect 2135 306 2136 307
rect 2143 307 2149 308
rect 2143 306 2144 307
rect 2135 304 2144 306
rect 2135 303 2136 304
rect 2130 302 2136 303
rect 2143 303 2144 304
rect 2148 303 2149 307
rect 2223 307 2232 308
rect 2143 302 2149 303
rect 2198 303 2204 304
rect 2118 298 2124 299
rect 2198 299 2199 303
rect 2203 299 2204 303
rect 2223 303 2224 307
rect 2231 303 2232 307
rect 2290 307 2296 308
rect 2223 302 2232 303
rect 2278 303 2284 304
rect 2198 298 2204 299
rect 2278 299 2279 303
rect 2283 299 2284 303
rect 2290 303 2291 307
rect 2295 306 2296 307
rect 2303 307 2309 308
rect 2303 306 2304 307
rect 2295 304 2304 306
rect 2295 303 2296 304
rect 2290 302 2296 303
rect 2303 303 2304 304
rect 2308 303 2309 307
rect 2370 307 2376 308
rect 2303 302 2309 303
rect 2358 303 2364 304
rect 2278 298 2284 299
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2370 303 2371 307
rect 2375 306 2376 307
rect 2383 307 2389 308
rect 2383 306 2384 307
rect 2375 304 2384 306
rect 2375 303 2376 304
rect 2370 302 2376 303
rect 2383 303 2384 304
rect 2388 303 2389 307
rect 2383 302 2389 303
rect 2358 298 2364 299
rect 1548 292 1802 294
rect 1548 291 1549 292
rect 1543 290 1549 291
rect 110 287 116 288
rect 159 287 165 288
rect 159 283 160 287
rect 164 283 165 287
rect 159 282 165 283
rect 198 287 205 288
rect 198 283 199 287
rect 204 283 205 287
rect 198 282 205 283
rect 230 287 236 288
rect 230 283 231 287
rect 235 286 236 287
rect 239 287 245 288
rect 239 286 240 287
rect 235 284 240 286
rect 235 283 236 284
rect 230 282 236 283
rect 239 283 240 284
rect 244 283 245 287
rect 239 282 245 283
rect 250 287 256 288
rect 250 283 251 287
rect 255 286 256 287
rect 279 287 285 288
rect 279 286 280 287
rect 255 284 280 286
rect 255 283 256 284
rect 250 282 256 283
rect 279 283 280 284
rect 284 283 285 287
rect 279 282 285 283
rect 319 287 325 288
rect 319 283 320 287
rect 324 283 325 287
rect 319 282 325 283
rect 359 287 365 288
rect 359 283 360 287
rect 364 283 365 287
rect 359 282 365 283
rect 382 287 388 288
rect 382 283 383 287
rect 387 286 388 287
rect 415 287 421 288
rect 415 286 416 287
rect 387 284 416 286
rect 387 283 388 284
rect 382 282 388 283
rect 415 283 416 284
rect 420 283 421 287
rect 415 282 421 283
rect 438 287 444 288
rect 438 283 439 287
rect 443 286 444 287
rect 471 287 477 288
rect 471 286 472 287
rect 443 284 472 286
rect 443 283 444 284
rect 438 282 444 283
rect 471 283 472 284
rect 476 283 477 287
rect 471 282 477 283
rect 519 287 525 288
rect 519 283 520 287
rect 524 283 525 287
rect 519 282 525 283
rect 534 287 540 288
rect 534 283 535 287
rect 539 286 540 287
rect 567 287 573 288
rect 567 286 568 287
rect 539 284 568 286
rect 539 283 540 284
rect 534 282 540 283
rect 567 283 568 284
rect 572 283 573 287
rect 567 282 573 283
rect 615 287 621 288
rect 615 283 616 287
rect 620 286 621 287
rect 630 287 636 288
rect 630 286 631 287
rect 620 284 631 286
rect 620 283 621 284
rect 615 282 621 283
rect 630 283 631 284
rect 635 283 636 287
rect 630 282 636 283
rect 654 287 660 288
rect 654 283 655 287
rect 659 286 660 287
rect 663 287 669 288
rect 663 286 664 287
rect 659 284 664 286
rect 659 283 660 284
rect 654 282 660 283
rect 663 283 664 284
rect 668 283 669 287
rect 663 282 669 283
rect 678 287 684 288
rect 678 283 679 287
rect 683 286 684 287
rect 711 287 717 288
rect 711 286 712 287
rect 683 284 712 286
rect 683 283 684 284
rect 678 282 684 283
rect 711 283 712 284
rect 716 283 717 287
rect 711 282 717 283
rect 726 287 732 288
rect 726 283 727 287
rect 731 286 732 287
rect 759 287 765 288
rect 759 286 760 287
rect 731 284 760 286
rect 731 283 732 284
rect 726 282 732 283
rect 759 283 760 284
rect 764 283 765 287
rect 759 282 765 283
rect 774 287 780 288
rect 774 283 775 287
rect 779 286 780 287
rect 807 287 813 288
rect 807 286 808 287
rect 779 284 808 286
rect 779 283 780 284
rect 774 282 780 283
rect 807 283 808 284
rect 812 283 813 287
rect 807 282 813 283
rect 862 287 869 288
rect 1238 287 1244 288
rect 862 283 863 287
rect 868 283 869 287
rect 862 282 869 283
rect 1538 283 1544 284
rect 150 279 156 280
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 150 275 151 279
rect 155 278 156 279
rect 319 278 321 282
rect 155 276 321 278
rect 521 278 523 282
rect 1278 280 1284 281
rect 670 279 676 280
rect 670 278 671 279
rect 521 276 671 278
rect 155 275 156 276
rect 150 274 156 275
rect 670 275 671 276
rect 675 275 676 279
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 1538 279 1539 283
rect 1543 282 1544 283
rect 1698 283 1704 284
rect 1543 280 1558 282
rect 1543 279 1544 280
rect 1538 278 1544 279
rect 670 274 676 275
rect 1238 275 1244 276
rect 1278 275 1284 276
rect 1535 275 1541 276
rect 110 270 116 271
rect 1238 271 1239 275
rect 1243 271 1244 275
rect 1238 270 1244 271
rect 1535 271 1536 275
rect 1540 274 1541 275
rect 1543 275 1549 276
rect 1543 274 1544 275
rect 1540 272 1544 274
rect 1540 271 1541 272
rect 1535 270 1541 271
rect 1543 271 1544 272
rect 1548 271 1549 275
rect 1556 274 1558 280
rect 1698 279 1699 283
rect 1703 282 1704 283
rect 1778 283 1784 284
rect 1703 280 1718 282
rect 1703 279 1704 280
rect 1698 278 1704 279
rect 1575 275 1581 276
rect 1575 274 1576 275
rect 1556 272 1576 274
rect 1543 270 1549 271
rect 1575 271 1576 272
rect 1580 271 1581 275
rect 1575 270 1581 271
rect 1598 275 1604 276
rect 1598 271 1599 275
rect 1603 274 1604 275
rect 1615 275 1621 276
rect 1615 274 1616 275
rect 1603 272 1616 274
rect 1603 271 1604 272
rect 1598 270 1604 271
rect 1615 271 1616 272
rect 1620 271 1621 275
rect 1615 270 1621 271
rect 1655 275 1661 276
rect 1655 271 1656 275
rect 1660 274 1661 275
rect 1678 275 1684 276
rect 1678 274 1679 275
rect 1660 272 1679 274
rect 1660 271 1661 272
rect 1655 270 1661 271
rect 1678 271 1679 272
rect 1683 271 1684 275
rect 1678 270 1684 271
rect 1686 275 1692 276
rect 1686 271 1687 275
rect 1691 274 1692 275
rect 1695 275 1701 276
rect 1695 274 1696 275
rect 1691 272 1696 274
rect 1691 271 1692 272
rect 1686 270 1692 271
rect 1695 271 1696 272
rect 1700 271 1701 275
rect 1716 274 1718 280
rect 1778 279 1779 283
rect 1783 282 1784 283
rect 1783 280 1798 282
rect 1783 279 1784 280
rect 1778 278 1784 279
rect 1735 275 1741 276
rect 1735 274 1736 275
rect 1716 272 1736 274
rect 1695 270 1701 271
rect 1735 271 1736 272
rect 1740 271 1741 275
rect 1735 270 1741 271
rect 1766 275 1772 276
rect 1766 271 1767 275
rect 1771 274 1772 275
rect 1775 275 1781 276
rect 1775 274 1776 275
rect 1771 272 1776 274
rect 1771 271 1772 272
rect 1766 270 1772 271
rect 1775 271 1776 272
rect 1780 271 1781 275
rect 1796 274 1798 280
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 1815 275 1821 276
rect 1815 274 1816 275
rect 1796 272 1816 274
rect 1775 270 1781 271
rect 1815 271 1816 272
rect 1820 271 1821 275
rect 1815 270 1821 271
rect 1846 275 1852 276
rect 1846 271 1847 275
rect 1851 274 1852 275
rect 1863 275 1869 276
rect 1863 274 1864 275
rect 1851 272 1864 274
rect 1851 271 1852 272
rect 1846 270 1852 271
rect 1863 271 1864 272
rect 1868 271 1869 275
rect 1863 270 1869 271
rect 1894 275 1900 276
rect 1894 271 1895 275
rect 1899 274 1900 275
rect 1927 275 1933 276
rect 1927 274 1928 275
rect 1899 272 1928 274
rect 1899 271 1900 272
rect 1894 270 1900 271
rect 1927 271 1928 272
rect 1932 271 1933 275
rect 1927 270 1933 271
rect 1958 275 1964 276
rect 1958 271 1959 275
rect 1963 274 1964 275
rect 1991 275 1997 276
rect 1991 274 1992 275
rect 1963 272 1992 274
rect 1963 271 1964 272
rect 1958 270 1964 271
rect 1991 271 1992 272
rect 1996 271 1997 275
rect 1991 270 1997 271
rect 2026 275 2032 276
rect 2026 271 2027 275
rect 2031 274 2032 275
rect 2063 275 2069 276
rect 2063 274 2064 275
rect 2031 272 2064 274
rect 2031 271 2032 272
rect 2026 270 2032 271
rect 2063 271 2064 272
rect 2068 271 2069 275
rect 2063 270 2069 271
rect 2110 275 2116 276
rect 2110 271 2111 275
rect 2115 274 2116 275
rect 2143 275 2149 276
rect 2143 274 2144 275
rect 2115 272 2144 274
rect 2115 271 2116 272
rect 2110 270 2116 271
rect 2143 271 2144 272
rect 2148 271 2149 275
rect 2143 270 2149 271
rect 2223 275 2229 276
rect 2223 271 2224 275
rect 2228 274 2229 275
rect 2290 275 2296 276
rect 2290 274 2291 275
rect 2228 272 2291 274
rect 2228 271 2229 272
rect 2223 270 2229 271
rect 2290 271 2291 272
rect 2295 271 2296 275
rect 2290 270 2296 271
rect 2303 275 2309 276
rect 2303 271 2304 275
rect 2308 274 2309 275
rect 2370 275 2376 276
rect 2370 274 2371 275
rect 2308 272 2371 274
rect 2308 271 2309 272
rect 2303 270 2309 271
rect 2370 271 2371 272
rect 2375 271 2376 275
rect 2370 270 2376 271
rect 2383 275 2389 276
rect 2406 275 2412 276
rect 2383 271 2384 275
rect 2388 271 2389 275
rect 2383 270 2389 271
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 174 268 180 269
rect 174 264 175 268
rect 179 264 180 268
rect 174 263 180 264
rect 214 268 220 269
rect 214 264 215 268
rect 219 264 220 268
rect 214 263 220 264
rect 254 268 260 269
rect 254 264 255 268
rect 259 264 260 268
rect 254 263 260 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 334 268 340 269
rect 334 264 335 268
rect 339 264 340 268
rect 334 263 340 264
rect 390 268 396 269
rect 390 264 391 268
rect 395 264 396 268
rect 390 263 396 264
rect 446 268 452 269
rect 446 264 447 268
rect 451 264 452 268
rect 446 263 452 264
rect 494 268 500 269
rect 494 264 495 268
rect 499 264 500 268
rect 494 263 500 264
rect 542 268 548 269
rect 542 264 543 268
rect 547 264 548 268
rect 542 263 548 264
rect 590 268 596 269
rect 590 264 591 268
rect 595 264 596 268
rect 590 263 596 264
rect 638 268 644 269
rect 638 264 639 268
rect 643 264 644 268
rect 638 263 644 264
rect 686 268 692 269
rect 686 264 687 268
rect 691 264 692 268
rect 686 263 692 264
rect 734 268 740 269
rect 734 264 735 268
rect 739 264 740 268
rect 734 263 740 264
rect 782 268 788 269
rect 782 264 783 268
rect 787 264 788 268
rect 782 263 788 264
rect 838 268 844 269
rect 838 264 839 268
rect 843 264 844 268
rect 2322 267 2328 268
rect 838 263 844 264
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 2322 263 2323 267
rect 2327 266 2328 267
rect 2384 266 2386 270
rect 2327 264 2386 266
rect 2327 263 2328 264
rect 2322 262 2328 263
rect 2406 263 2412 264
rect 1278 258 1284 259
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 1510 256 1516 257
rect 1510 252 1511 256
rect 1515 252 1516 256
rect 1510 251 1516 252
rect 1550 256 1556 257
rect 1550 252 1551 256
rect 1555 252 1556 256
rect 1550 251 1556 252
rect 1590 256 1596 257
rect 1590 252 1591 256
rect 1595 252 1596 256
rect 1590 251 1596 252
rect 1630 256 1636 257
rect 1630 252 1631 256
rect 1635 252 1636 256
rect 1630 251 1636 252
rect 1670 256 1676 257
rect 1670 252 1671 256
rect 1675 252 1676 256
rect 1670 251 1676 252
rect 1710 256 1716 257
rect 1710 252 1711 256
rect 1715 252 1716 256
rect 1710 251 1716 252
rect 1750 256 1756 257
rect 1750 252 1751 256
rect 1755 252 1756 256
rect 1750 251 1756 252
rect 1790 256 1796 257
rect 1790 252 1791 256
rect 1795 252 1796 256
rect 1790 251 1796 252
rect 1838 256 1844 257
rect 1838 252 1839 256
rect 1843 252 1844 256
rect 1838 251 1844 252
rect 1902 256 1908 257
rect 1902 252 1903 256
rect 1907 252 1908 256
rect 1902 251 1908 252
rect 1966 256 1972 257
rect 1966 252 1967 256
rect 1971 252 1972 256
rect 1966 251 1972 252
rect 2038 256 2044 257
rect 2038 252 2039 256
rect 2043 252 2044 256
rect 2038 251 2044 252
rect 2118 256 2124 257
rect 2118 252 2119 256
rect 2123 252 2124 256
rect 2118 251 2124 252
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2278 256 2284 257
rect 2278 252 2279 256
rect 2283 252 2284 256
rect 2278 251 2284 252
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 134 248 140 249
rect 134 244 135 248
rect 139 244 140 248
rect 134 243 140 244
rect 222 248 228 249
rect 222 244 223 248
rect 227 244 228 248
rect 222 243 228 244
rect 310 248 316 249
rect 310 244 311 248
rect 315 244 316 248
rect 310 243 316 244
rect 390 248 396 249
rect 390 244 391 248
rect 395 244 396 248
rect 390 243 396 244
rect 462 248 468 249
rect 462 244 463 248
rect 467 244 468 248
rect 462 243 468 244
rect 526 248 532 249
rect 526 244 527 248
rect 531 244 532 248
rect 526 243 532 244
rect 590 248 596 249
rect 590 244 591 248
rect 595 244 596 248
rect 590 243 596 244
rect 646 248 652 249
rect 646 244 647 248
rect 651 244 652 248
rect 646 243 652 244
rect 694 248 700 249
rect 694 244 695 248
rect 699 244 700 248
rect 694 243 700 244
rect 734 248 740 249
rect 734 244 735 248
rect 739 244 740 248
rect 734 243 740 244
rect 782 248 788 249
rect 782 244 783 248
rect 787 244 788 248
rect 782 243 788 244
rect 830 248 836 249
rect 830 244 831 248
rect 835 244 836 248
rect 830 243 836 244
rect 878 248 884 249
rect 878 244 879 248
rect 883 244 884 248
rect 878 243 884 244
rect 926 248 932 249
rect 926 244 927 248
rect 931 244 932 248
rect 926 243 932 244
rect 974 248 980 249
rect 974 244 975 248
rect 979 244 980 248
rect 974 243 980 244
rect 1022 248 1028 249
rect 1022 244 1023 248
rect 1027 244 1028 248
rect 1022 243 1028 244
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 1238 241 1244 242
rect 1238 237 1239 241
rect 1243 237 1244 241
rect 1238 236 1244 237
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 794 235 800 236
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1454 240 1460 241
rect 1454 236 1455 240
rect 1459 236 1460 240
rect 1454 235 1460 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1566 240 1572 241
rect 1566 236 1567 240
rect 1571 236 1572 240
rect 1566 235 1572 236
rect 1630 240 1636 241
rect 1630 236 1631 240
rect 1635 236 1636 240
rect 1630 235 1636 236
rect 1702 240 1708 241
rect 1702 236 1703 240
rect 1707 236 1708 240
rect 1702 235 1708 236
rect 1774 240 1780 241
rect 1774 236 1775 240
rect 1779 236 1780 240
rect 1774 235 1780 236
rect 1854 240 1860 241
rect 1854 236 1855 240
rect 1859 236 1860 240
rect 1854 235 1860 236
rect 1942 240 1948 241
rect 1942 236 1943 240
rect 1947 236 1948 240
rect 1942 235 1948 236
rect 2030 240 2036 241
rect 2030 236 2031 240
rect 2035 236 2036 240
rect 2030 235 2036 236
rect 2118 240 2124 241
rect 2118 236 2119 240
rect 2123 236 2124 240
rect 2118 235 2124 236
rect 2206 240 2212 241
rect 2206 236 2207 240
rect 2211 236 2212 240
rect 2206 235 2212 236
rect 2294 240 2300 241
rect 2294 236 2295 240
rect 2299 236 2300 240
rect 2294 235 2300 236
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 794 234 795 235
rect 736 232 795 234
rect 158 227 165 228
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 158 223 159 227
rect 164 223 165 227
rect 158 222 165 223
rect 247 227 253 228
rect 247 223 248 227
rect 252 226 253 227
rect 286 227 292 228
rect 252 224 283 226
rect 252 223 253 224
rect 247 222 253 223
rect 110 219 116 220
rect 281 218 283 224
rect 286 223 287 227
rect 291 226 292 227
rect 335 227 341 228
rect 335 226 336 227
rect 291 224 336 226
rect 291 223 292 224
rect 286 222 292 223
rect 335 223 336 224
rect 340 223 341 227
rect 335 222 341 223
rect 343 227 349 228
rect 343 223 344 227
rect 348 226 349 227
rect 415 227 421 228
rect 415 226 416 227
rect 348 224 416 226
rect 348 223 349 224
rect 343 222 349 223
rect 415 223 416 224
rect 420 223 421 227
rect 415 222 421 223
rect 423 227 429 228
rect 423 223 424 227
rect 428 226 429 227
rect 487 227 493 228
rect 487 226 488 227
rect 428 224 488 226
rect 428 223 429 224
rect 423 222 429 223
rect 487 223 488 224
rect 492 223 493 227
rect 487 222 493 223
rect 495 227 501 228
rect 495 223 496 227
rect 500 226 501 227
rect 551 227 557 228
rect 551 226 552 227
rect 500 224 552 226
rect 500 223 501 224
rect 495 222 501 223
rect 551 223 552 224
rect 556 223 557 227
rect 551 222 557 223
rect 559 227 565 228
rect 559 223 560 227
rect 564 226 565 227
rect 615 227 621 228
rect 615 226 616 227
rect 564 224 616 226
rect 564 223 565 224
rect 559 222 565 223
rect 615 223 616 224
rect 620 223 621 227
rect 615 222 621 223
rect 623 227 629 228
rect 623 223 624 227
rect 628 226 629 227
rect 671 227 677 228
rect 671 226 672 227
rect 628 224 672 226
rect 628 223 629 224
rect 623 222 629 223
rect 671 223 672 224
rect 676 223 677 227
rect 671 222 677 223
rect 719 227 725 228
rect 719 223 720 227
rect 724 226 725 227
rect 736 226 738 232
rect 794 231 795 232
rect 799 231 800 235
rect 794 230 800 231
rect 1278 233 1284 234
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 724 224 738 226
rect 742 227 748 228
rect 724 223 725 224
rect 719 222 725 223
rect 742 223 743 227
rect 747 226 748 227
rect 759 227 765 228
rect 759 226 760 227
rect 747 224 760 226
rect 747 223 748 224
rect 742 222 748 223
rect 759 223 760 224
rect 764 223 765 227
rect 759 222 765 223
rect 767 227 773 228
rect 767 223 768 227
rect 772 226 773 227
rect 807 227 813 228
rect 807 226 808 227
rect 772 224 808 226
rect 772 223 773 224
rect 767 222 773 223
rect 807 223 808 224
rect 812 223 813 227
rect 807 222 813 223
rect 815 227 821 228
rect 815 223 816 227
rect 820 226 821 227
rect 855 227 861 228
rect 855 226 856 227
rect 820 224 856 226
rect 820 223 821 224
rect 815 222 821 223
rect 855 223 856 224
rect 860 223 861 227
rect 855 222 861 223
rect 863 227 869 228
rect 863 223 864 227
rect 868 226 869 227
rect 903 227 909 228
rect 903 226 904 227
rect 868 224 904 226
rect 868 223 869 224
rect 863 222 869 223
rect 903 223 904 224
rect 908 223 909 227
rect 903 222 909 223
rect 911 227 917 228
rect 911 223 912 227
rect 916 226 917 227
rect 951 227 957 228
rect 951 226 952 227
rect 916 224 952 226
rect 916 223 917 224
rect 911 222 917 223
rect 951 223 952 224
rect 956 223 957 227
rect 951 222 957 223
rect 959 227 965 228
rect 959 223 960 227
rect 964 226 965 227
rect 999 227 1005 228
rect 999 226 1000 227
rect 964 224 1000 226
rect 964 223 965 224
rect 959 222 965 223
rect 999 223 1000 224
rect 1004 223 1005 227
rect 999 222 1005 223
rect 1007 227 1013 228
rect 1007 223 1008 227
rect 1012 226 1013 227
rect 1047 227 1053 228
rect 1047 226 1048 227
rect 1012 224 1048 226
rect 1012 223 1013 224
rect 1007 222 1013 223
rect 1047 223 1048 224
rect 1052 223 1053 227
rect 2130 227 2136 228
rect 2130 226 2131 227
rect 1047 222 1053 223
rect 1238 224 1244 225
rect 1238 220 1239 224
rect 1243 220 1244 224
rect 1800 224 2131 226
rect 1800 220 1802 224
rect 2130 223 2131 224
rect 2135 223 2136 227
rect 2130 222 2136 223
rect 614 219 620 220
rect 1238 219 1244 220
rect 1391 219 1397 220
rect 614 218 615 219
rect 281 216 615 218
rect 614 215 615 216
rect 619 215 620 219
rect 614 214 620 215
rect 1278 216 1284 217
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1391 215 1392 219
rect 1396 218 1397 219
rect 1414 219 1420 220
rect 1396 216 1410 218
rect 1396 215 1397 216
rect 1391 214 1397 215
rect 1278 211 1284 212
rect 1408 210 1410 216
rect 1414 215 1415 219
rect 1419 218 1420 219
rect 1431 219 1437 220
rect 1431 218 1432 219
rect 1419 216 1432 218
rect 1419 215 1420 216
rect 1414 214 1420 215
rect 1431 215 1432 216
rect 1436 215 1437 219
rect 1431 214 1437 215
rect 1439 219 1445 220
rect 1439 215 1440 219
rect 1444 218 1445 219
rect 1479 219 1485 220
rect 1479 218 1480 219
rect 1444 216 1480 218
rect 1444 215 1445 216
rect 1439 214 1445 215
rect 1479 215 1480 216
rect 1484 215 1485 219
rect 1479 214 1485 215
rect 1487 219 1493 220
rect 1487 215 1488 219
rect 1492 218 1493 219
rect 1535 219 1541 220
rect 1535 218 1536 219
rect 1492 216 1536 218
rect 1492 215 1493 216
rect 1487 214 1493 215
rect 1535 215 1536 216
rect 1540 215 1541 219
rect 1535 214 1541 215
rect 1543 219 1549 220
rect 1543 215 1544 219
rect 1548 218 1549 219
rect 1591 219 1597 220
rect 1591 218 1592 219
rect 1548 216 1592 218
rect 1548 215 1549 216
rect 1543 214 1549 215
rect 1591 215 1592 216
rect 1596 215 1597 219
rect 1591 214 1597 215
rect 1599 219 1605 220
rect 1599 215 1600 219
rect 1604 218 1605 219
rect 1655 219 1661 220
rect 1655 218 1656 219
rect 1604 216 1656 218
rect 1604 215 1605 216
rect 1599 214 1605 215
rect 1655 215 1656 216
rect 1660 215 1661 219
rect 1655 214 1661 215
rect 1663 219 1669 220
rect 1663 215 1664 219
rect 1668 218 1669 219
rect 1727 219 1733 220
rect 1727 218 1728 219
rect 1668 216 1728 218
rect 1668 215 1669 216
rect 1663 214 1669 215
rect 1727 215 1728 216
rect 1732 215 1733 219
rect 1727 214 1733 215
rect 1799 219 1805 220
rect 1799 215 1800 219
rect 1804 215 1805 219
rect 1799 214 1805 215
rect 1807 219 1813 220
rect 1807 215 1808 219
rect 1812 218 1813 219
rect 1879 219 1885 220
rect 1879 218 1880 219
rect 1812 216 1880 218
rect 1812 215 1813 216
rect 1807 214 1813 215
rect 1879 215 1880 216
rect 1884 215 1885 219
rect 1879 214 1885 215
rect 1887 219 1893 220
rect 1887 215 1888 219
rect 1892 218 1893 219
rect 1967 219 1973 220
rect 1967 218 1968 219
rect 1892 216 1968 218
rect 1892 215 1893 216
rect 1887 214 1893 215
rect 1967 215 1968 216
rect 1972 215 1973 219
rect 1967 214 1973 215
rect 1975 219 1981 220
rect 1975 215 1976 219
rect 1980 218 1981 219
rect 2055 219 2061 220
rect 2055 218 2056 219
rect 1980 216 2056 218
rect 1980 215 1981 216
rect 1975 214 1981 215
rect 2055 215 2056 216
rect 2060 215 2061 219
rect 2055 214 2061 215
rect 2063 219 2069 220
rect 2063 215 2064 219
rect 2068 218 2069 219
rect 2143 219 2149 220
rect 2143 218 2144 219
rect 2068 216 2144 218
rect 2068 215 2069 216
rect 2063 214 2069 215
rect 2143 215 2144 216
rect 2148 215 2149 219
rect 2143 214 2149 215
rect 2226 219 2237 220
rect 2226 215 2227 219
rect 2231 215 2232 219
rect 2236 215 2237 219
rect 2226 214 2237 215
rect 2319 219 2325 220
rect 2319 215 2320 219
rect 2324 218 2325 219
rect 2374 219 2380 220
rect 2374 218 2375 219
rect 2324 216 2375 218
rect 2324 215 2325 216
rect 2319 214 2325 215
rect 2374 215 2375 216
rect 2379 215 2380 219
rect 2374 214 2380 215
rect 2382 219 2389 220
rect 2382 215 2383 219
rect 2388 215 2389 219
rect 2382 214 2389 215
rect 2406 216 2412 217
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 1670 211 1676 212
rect 2406 211 2412 212
rect 1670 210 1671 211
rect 1408 208 1671 210
rect 1670 207 1671 208
rect 1675 207 1676 211
rect 1670 206 1676 207
rect 134 201 140 202
rect 134 197 135 201
rect 139 197 140 201
rect 134 196 140 197
rect 222 201 228 202
rect 222 197 223 201
rect 227 197 228 201
rect 222 196 228 197
rect 310 201 316 202
rect 310 197 311 201
rect 315 197 316 201
rect 310 196 316 197
rect 390 201 396 202
rect 390 197 391 201
rect 395 197 396 201
rect 390 196 396 197
rect 462 201 468 202
rect 462 197 463 201
rect 467 197 468 201
rect 462 196 468 197
rect 526 201 532 202
rect 526 197 527 201
rect 531 197 532 201
rect 526 196 532 197
rect 590 201 596 202
rect 590 197 591 201
rect 595 197 596 201
rect 590 196 596 197
rect 646 201 652 202
rect 646 197 647 201
rect 651 197 652 201
rect 646 196 652 197
rect 694 201 700 202
rect 694 197 695 201
rect 699 197 700 201
rect 694 196 700 197
rect 734 201 740 202
rect 734 197 735 201
rect 739 197 740 201
rect 734 196 740 197
rect 782 201 788 202
rect 782 197 783 201
rect 787 197 788 201
rect 782 196 788 197
rect 830 201 836 202
rect 830 197 831 201
rect 835 197 836 201
rect 830 196 836 197
rect 878 201 884 202
rect 878 197 879 201
rect 883 197 884 201
rect 878 196 884 197
rect 926 201 932 202
rect 926 197 927 201
rect 931 197 932 201
rect 926 196 932 197
rect 974 201 980 202
rect 974 197 975 201
rect 979 197 980 201
rect 974 196 980 197
rect 1022 201 1028 202
rect 1022 197 1023 201
rect 1027 197 1028 201
rect 1022 196 1028 197
rect 150 195 156 196
rect 150 191 151 195
rect 155 194 156 195
rect 159 195 165 196
rect 159 194 160 195
rect 155 192 160 194
rect 155 191 156 192
rect 150 190 156 191
rect 159 191 160 192
rect 164 191 165 195
rect 159 190 165 191
rect 247 195 253 196
rect 247 191 248 195
rect 252 194 253 195
rect 286 195 292 196
rect 286 194 287 195
rect 252 192 287 194
rect 252 191 253 192
rect 247 190 253 191
rect 286 191 287 192
rect 291 191 292 195
rect 286 190 292 191
rect 335 195 341 196
rect 335 191 336 195
rect 340 194 341 195
rect 343 195 349 196
rect 343 194 344 195
rect 340 192 344 194
rect 340 191 341 192
rect 335 190 341 191
rect 343 191 344 192
rect 348 191 349 195
rect 343 190 349 191
rect 415 195 421 196
rect 415 191 416 195
rect 420 194 421 195
rect 423 195 429 196
rect 423 194 424 195
rect 420 192 424 194
rect 420 191 421 192
rect 415 190 421 191
rect 423 191 424 192
rect 428 191 429 195
rect 423 190 429 191
rect 487 195 493 196
rect 487 191 488 195
rect 492 194 493 195
rect 495 195 501 196
rect 495 194 496 195
rect 492 192 496 194
rect 492 191 493 192
rect 487 190 493 191
rect 495 191 496 192
rect 500 191 501 195
rect 495 190 501 191
rect 551 195 557 196
rect 551 191 552 195
rect 556 194 557 195
rect 559 195 565 196
rect 559 194 560 195
rect 556 192 560 194
rect 556 191 557 192
rect 551 190 557 191
rect 559 191 560 192
rect 564 191 565 195
rect 559 190 565 191
rect 615 195 621 196
rect 615 191 616 195
rect 620 194 621 195
rect 623 195 629 196
rect 623 194 624 195
rect 620 192 624 194
rect 620 191 621 192
rect 615 190 621 191
rect 623 191 624 192
rect 628 191 629 195
rect 623 190 629 191
rect 670 195 677 196
rect 670 191 671 195
rect 676 191 677 195
rect 670 190 677 191
rect 719 195 725 196
rect 719 191 720 195
rect 724 194 725 195
rect 742 195 748 196
rect 742 194 743 195
rect 724 192 743 194
rect 724 191 725 192
rect 719 190 725 191
rect 742 191 743 192
rect 747 191 748 195
rect 742 190 748 191
rect 759 195 765 196
rect 759 191 760 195
rect 764 194 765 195
rect 767 195 773 196
rect 767 194 768 195
rect 764 192 768 194
rect 764 191 765 192
rect 759 190 765 191
rect 767 191 768 192
rect 772 191 773 195
rect 767 190 773 191
rect 807 195 813 196
rect 807 191 808 195
rect 812 194 813 195
rect 815 195 821 196
rect 815 194 816 195
rect 812 192 816 194
rect 812 191 813 192
rect 807 190 813 191
rect 815 191 816 192
rect 820 191 821 195
rect 815 190 821 191
rect 855 195 861 196
rect 855 191 856 195
rect 860 194 861 195
rect 863 195 869 196
rect 863 194 864 195
rect 860 192 864 194
rect 860 191 861 192
rect 855 190 861 191
rect 863 191 864 192
rect 868 191 869 195
rect 863 190 869 191
rect 903 195 909 196
rect 903 191 904 195
rect 908 194 909 195
rect 911 195 917 196
rect 911 194 912 195
rect 908 192 912 194
rect 908 191 909 192
rect 903 190 909 191
rect 911 191 912 192
rect 916 191 917 195
rect 911 190 917 191
rect 951 195 957 196
rect 951 191 952 195
rect 956 194 957 195
rect 959 195 965 196
rect 959 194 960 195
rect 956 192 960 194
rect 956 191 957 192
rect 951 190 957 191
rect 959 191 960 192
rect 964 191 965 195
rect 959 190 965 191
rect 999 195 1005 196
rect 999 191 1000 195
rect 1004 194 1005 195
rect 1007 195 1013 196
rect 1007 194 1008 195
rect 1004 192 1008 194
rect 1004 191 1005 192
rect 999 190 1005 191
rect 1007 191 1008 192
rect 1012 191 1013 195
rect 1007 190 1013 191
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 194 1044 195
rect 1047 195 1053 196
rect 1047 194 1048 195
rect 1043 192 1048 194
rect 1043 191 1044 192
rect 1038 190 1044 191
rect 1047 191 1048 192
rect 1052 191 1053 195
rect 1047 190 1053 191
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1454 193 1460 194
rect 1454 189 1455 193
rect 1459 189 1460 193
rect 1454 188 1460 189
rect 1510 193 1516 194
rect 1510 189 1511 193
rect 1515 189 1516 193
rect 1510 188 1516 189
rect 1566 193 1572 194
rect 1566 189 1567 193
rect 1571 189 1572 193
rect 1566 188 1572 189
rect 1630 193 1636 194
rect 1630 189 1631 193
rect 1635 189 1636 193
rect 1630 188 1636 189
rect 1702 193 1708 194
rect 1702 189 1703 193
rect 1707 189 1708 193
rect 1702 188 1708 189
rect 1774 193 1780 194
rect 1774 189 1775 193
rect 1779 189 1780 193
rect 1774 188 1780 189
rect 1854 193 1860 194
rect 1854 189 1855 193
rect 1859 189 1860 193
rect 1854 188 1860 189
rect 1942 193 1948 194
rect 1942 189 1943 193
rect 1947 189 1948 193
rect 1942 188 1948 189
rect 2030 193 2036 194
rect 2030 189 2031 193
rect 2035 189 2036 193
rect 2030 188 2036 189
rect 2118 193 2124 194
rect 2118 189 2119 193
rect 2123 189 2124 193
rect 2118 188 2124 189
rect 2206 193 2212 194
rect 2206 189 2207 193
rect 2211 189 2212 193
rect 2206 188 2212 189
rect 2294 193 2300 194
rect 2294 189 2295 193
rect 2299 189 2300 193
rect 2294 188 2300 189
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 1391 187 1397 188
rect 1391 183 1392 187
rect 1396 186 1397 187
rect 1414 187 1420 188
rect 1414 186 1415 187
rect 1396 184 1415 186
rect 1396 183 1397 184
rect 1391 182 1397 183
rect 1414 183 1415 184
rect 1419 183 1420 187
rect 1414 182 1420 183
rect 1431 187 1437 188
rect 1431 183 1432 187
rect 1436 186 1437 187
rect 1439 187 1445 188
rect 1439 186 1440 187
rect 1436 184 1440 186
rect 1436 183 1437 184
rect 1431 182 1437 183
rect 1439 183 1440 184
rect 1444 183 1445 187
rect 1439 182 1445 183
rect 1479 187 1485 188
rect 1479 183 1480 187
rect 1484 186 1485 187
rect 1487 187 1493 188
rect 1487 186 1488 187
rect 1484 184 1488 186
rect 1484 183 1485 184
rect 1479 182 1485 183
rect 1487 183 1488 184
rect 1492 183 1493 187
rect 1487 182 1493 183
rect 1535 187 1541 188
rect 1535 183 1536 187
rect 1540 186 1541 187
rect 1543 187 1549 188
rect 1543 186 1544 187
rect 1540 184 1544 186
rect 1540 183 1541 184
rect 1535 182 1541 183
rect 1543 183 1544 184
rect 1548 183 1549 187
rect 1543 182 1549 183
rect 1591 187 1597 188
rect 1591 183 1592 187
rect 1596 186 1597 187
rect 1599 187 1605 188
rect 1599 186 1600 187
rect 1596 184 1600 186
rect 1596 183 1597 184
rect 1591 182 1597 183
rect 1599 183 1600 184
rect 1604 183 1605 187
rect 1599 182 1605 183
rect 1655 187 1661 188
rect 1655 183 1656 187
rect 1660 186 1661 187
rect 1663 187 1669 188
rect 1663 186 1664 187
rect 1660 184 1664 186
rect 1660 183 1661 184
rect 1655 182 1661 183
rect 1663 183 1664 184
rect 1668 183 1669 187
rect 1663 182 1669 183
rect 1678 187 1684 188
rect 1678 183 1679 187
rect 1683 186 1684 187
rect 1727 187 1733 188
rect 1727 186 1728 187
rect 1683 184 1728 186
rect 1683 183 1684 184
rect 1678 182 1684 183
rect 1727 183 1728 184
rect 1732 183 1733 187
rect 1727 182 1733 183
rect 1799 187 1805 188
rect 1799 183 1800 187
rect 1804 186 1805 187
rect 1807 187 1813 188
rect 1807 186 1808 187
rect 1804 184 1808 186
rect 1804 183 1805 184
rect 1799 182 1805 183
rect 1807 183 1808 184
rect 1812 183 1813 187
rect 1807 182 1813 183
rect 1879 187 1885 188
rect 1879 183 1880 187
rect 1884 186 1885 187
rect 1887 187 1893 188
rect 1887 186 1888 187
rect 1884 184 1888 186
rect 1884 183 1885 184
rect 1879 182 1885 183
rect 1887 183 1888 184
rect 1892 183 1893 187
rect 1887 182 1893 183
rect 1967 187 1973 188
rect 1967 183 1968 187
rect 1972 186 1973 187
rect 1975 187 1981 188
rect 1975 186 1976 187
rect 1972 184 1976 186
rect 1972 183 1973 184
rect 1967 182 1973 183
rect 1975 183 1976 184
rect 1980 183 1981 187
rect 1975 182 1981 183
rect 2055 187 2061 188
rect 2055 183 2056 187
rect 2060 186 2061 187
rect 2063 187 2069 188
rect 2063 186 2064 187
rect 2060 184 2064 186
rect 2060 183 2061 184
rect 2055 182 2061 183
rect 2063 183 2064 184
rect 2068 183 2069 187
rect 2143 187 2149 188
rect 2143 186 2144 187
rect 2063 182 2069 183
rect 2072 184 2144 186
rect 1738 179 1744 180
rect 1738 175 1739 179
rect 1743 178 1744 179
rect 2072 178 2074 184
rect 2143 183 2144 184
rect 2148 183 2149 187
rect 2143 182 2149 183
rect 2231 187 2237 188
rect 2231 183 2232 187
rect 2236 186 2237 187
rect 2262 187 2268 188
rect 2262 186 2263 187
rect 2236 184 2263 186
rect 2236 183 2237 184
rect 2231 182 2237 183
rect 2262 183 2263 184
rect 2267 183 2268 187
rect 2262 182 2268 183
rect 2319 187 2328 188
rect 2319 183 2320 187
rect 2327 183 2328 187
rect 2319 182 2328 183
rect 2374 187 2380 188
rect 2374 183 2375 187
rect 2379 186 2380 187
rect 2383 187 2389 188
rect 2383 186 2384 187
rect 2379 184 2384 186
rect 2379 183 2380 184
rect 2374 182 2380 183
rect 2383 183 2384 184
rect 2388 183 2389 187
rect 2383 182 2389 183
rect 1743 176 2074 178
rect 1743 175 1744 176
rect 1738 174 1744 175
rect 2022 163 2028 164
rect 2022 162 2023 163
rect 2008 160 2023 162
rect 1327 159 1336 160
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1327 155 1328 159
rect 1335 155 1336 159
rect 1367 159 1376 160
rect 1327 154 1336 155
rect 1342 155 1348 156
rect 1302 150 1308 151
rect 1342 151 1343 155
rect 1347 151 1348 155
rect 1367 155 1368 159
rect 1375 155 1376 159
rect 1407 159 1416 160
rect 1367 154 1376 155
rect 1382 155 1388 156
rect 1342 150 1348 151
rect 1382 151 1383 155
rect 1387 151 1388 155
rect 1407 155 1408 159
rect 1415 155 1416 159
rect 1447 159 1456 160
rect 1407 154 1416 155
rect 1422 155 1428 156
rect 1382 150 1388 151
rect 1422 151 1423 155
rect 1427 151 1428 155
rect 1447 155 1448 159
rect 1455 155 1456 159
rect 1487 159 1493 160
rect 1447 154 1456 155
rect 1462 155 1468 156
rect 1422 150 1428 151
rect 1462 151 1463 155
rect 1467 151 1468 155
rect 1487 155 1488 159
rect 1492 158 1493 159
rect 1510 159 1516 160
rect 1510 158 1511 159
rect 1492 156 1511 158
rect 1492 155 1493 156
rect 1487 154 1493 155
rect 1510 155 1511 156
rect 1515 155 1516 159
rect 1543 159 1549 160
rect 1510 154 1516 155
rect 1518 155 1524 156
rect 1462 150 1468 151
rect 1518 151 1519 155
rect 1523 151 1524 155
rect 1543 155 1544 159
rect 1548 158 1549 159
rect 1574 159 1580 160
rect 1574 158 1575 159
rect 1548 156 1575 158
rect 1548 155 1549 156
rect 1543 154 1549 155
rect 1574 155 1575 156
rect 1579 155 1580 159
rect 1607 159 1613 160
rect 1574 154 1580 155
rect 1582 155 1588 156
rect 1518 150 1524 151
rect 1582 151 1583 155
rect 1587 151 1588 155
rect 1607 155 1608 159
rect 1612 158 1613 159
rect 1638 159 1644 160
rect 1638 158 1639 159
rect 1612 156 1639 158
rect 1612 155 1613 156
rect 1607 154 1613 155
rect 1638 155 1639 156
rect 1643 155 1644 159
rect 1670 159 1677 160
rect 1638 154 1644 155
rect 1646 155 1652 156
rect 1582 150 1588 151
rect 1646 151 1647 155
rect 1651 151 1652 155
rect 1670 155 1671 159
rect 1676 155 1677 159
rect 1735 159 1741 160
rect 1670 154 1677 155
rect 1710 155 1716 156
rect 1646 150 1652 151
rect 1710 151 1711 155
rect 1715 151 1716 155
rect 1735 155 1736 159
rect 1740 158 1741 159
rect 1766 159 1772 160
rect 1766 158 1767 159
rect 1740 156 1767 158
rect 1740 155 1741 156
rect 1735 154 1741 155
rect 1766 155 1767 156
rect 1771 155 1772 159
rect 1799 159 1805 160
rect 1766 154 1772 155
rect 1774 155 1780 156
rect 1710 150 1716 151
rect 1774 151 1775 155
rect 1779 151 1780 155
rect 1799 155 1800 159
rect 1804 158 1805 159
rect 1822 159 1828 160
rect 1822 158 1823 159
rect 1804 156 1823 158
rect 1804 155 1805 156
rect 1799 154 1805 155
rect 1822 155 1823 156
rect 1827 155 1828 159
rect 1855 159 1861 160
rect 1822 154 1828 155
rect 1830 155 1836 156
rect 1774 150 1780 151
rect 1830 151 1831 155
rect 1835 151 1836 155
rect 1855 155 1856 159
rect 1860 158 1861 159
rect 1878 159 1884 160
rect 1878 158 1879 159
rect 1860 156 1879 158
rect 1860 155 1861 156
rect 1855 154 1861 155
rect 1878 155 1879 156
rect 1883 155 1884 159
rect 1911 159 1917 160
rect 1878 154 1884 155
rect 1886 155 1892 156
rect 1830 150 1836 151
rect 1886 151 1887 155
rect 1891 151 1892 155
rect 1911 155 1912 159
rect 1916 158 1917 159
rect 1926 159 1932 160
rect 1926 158 1927 159
rect 1916 156 1927 158
rect 1916 155 1917 156
rect 1911 154 1917 155
rect 1926 155 1927 156
rect 1931 155 1932 159
rect 1959 159 1968 160
rect 1926 154 1932 155
rect 1934 155 1940 156
rect 1886 150 1892 151
rect 1934 151 1935 155
rect 1939 151 1940 155
rect 1959 155 1960 159
rect 1967 155 1968 159
rect 1999 159 2005 160
rect 1959 154 1968 155
rect 1974 155 1980 156
rect 1934 150 1940 151
rect 1974 151 1975 155
rect 1979 151 1980 155
rect 1999 155 2000 159
rect 2004 158 2005 159
rect 2008 158 2010 160
rect 2022 159 2023 160
rect 2027 159 2028 163
rect 2070 163 2076 164
rect 2070 162 2071 163
rect 2048 160 2071 162
rect 2022 158 2028 159
rect 2039 159 2045 160
rect 2004 156 2010 158
rect 2004 155 2005 156
rect 1999 154 2005 155
rect 2014 155 2020 156
rect 1974 150 1980 151
rect 2014 151 2015 155
rect 2019 151 2020 155
rect 2039 155 2040 159
rect 2044 158 2045 159
rect 2048 158 2050 160
rect 2070 159 2071 160
rect 2075 159 2076 163
rect 2102 163 2108 164
rect 2102 162 2103 163
rect 2088 160 2103 162
rect 2070 158 2076 159
rect 2079 159 2085 160
rect 2044 156 2050 158
rect 2044 155 2045 156
rect 2039 154 2045 155
rect 2054 155 2060 156
rect 2014 150 2020 151
rect 2054 151 2055 155
rect 2059 151 2060 155
rect 2079 155 2080 159
rect 2084 158 2085 159
rect 2088 158 2090 160
rect 2102 159 2103 160
rect 2107 159 2108 163
rect 2286 163 2292 164
rect 2286 162 2287 163
rect 2273 160 2287 162
rect 2102 158 2108 159
rect 2119 159 2125 160
rect 2084 156 2090 158
rect 2084 155 2085 156
rect 2079 154 2085 155
rect 2094 155 2100 156
rect 2054 150 2060 151
rect 2094 151 2095 155
rect 2099 151 2100 155
rect 2119 155 2120 159
rect 2124 158 2125 159
rect 2134 159 2140 160
rect 2134 158 2135 159
rect 2124 156 2135 158
rect 2124 155 2125 156
rect 2119 154 2125 155
rect 2134 155 2135 156
rect 2139 155 2140 159
rect 2167 159 2173 160
rect 2134 154 2140 155
rect 2142 155 2148 156
rect 2094 150 2100 151
rect 2142 151 2143 155
rect 2147 151 2148 155
rect 2167 155 2168 159
rect 2172 158 2173 159
rect 2182 159 2188 160
rect 2182 158 2183 159
rect 2172 156 2183 158
rect 2172 155 2173 156
rect 2167 154 2173 155
rect 2182 155 2183 156
rect 2187 155 2188 159
rect 2215 159 2221 160
rect 2182 154 2188 155
rect 2190 155 2196 156
rect 2142 150 2148 151
rect 2190 151 2191 155
rect 2195 151 2196 155
rect 2215 155 2216 159
rect 2220 158 2221 159
rect 2226 159 2232 160
rect 2226 158 2227 159
rect 2220 156 2227 158
rect 2220 155 2221 156
rect 2215 154 2221 155
rect 2226 155 2227 156
rect 2231 155 2232 159
rect 2263 159 2269 160
rect 2226 154 2232 155
rect 2238 155 2244 156
rect 2190 150 2196 151
rect 2238 151 2239 155
rect 2243 151 2244 155
rect 2263 155 2264 159
rect 2268 158 2269 159
rect 2273 158 2275 160
rect 2286 159 2287 160
rect 2291 159 2292 163
rect 2334 163 2340 164
rect 2334 162 2335 163
rect 2312 160 2335 162
rect 2286 158 2292 159
rect 2303 159 2309 160
rect 2268 156 2275 158
rect 2268 155 2269 156
rect 2263 154 2269 155
rect 2278 155 2284 156
rect 2238 150 2244 151
rect 2278 151 2279 155
rect 2283 151 2284 155
rect 2303 155 2304 159
rect 2308 158 2309 159
rect 2312 158 2314 160
rect 2334 159 2335 160
rect 2339 159 2340 163
rect 2366 163 2372 164
rect 2366 162 2367 163
rect 2352 160 2367 162
rect 2334 158 2340 159
rect 2343 159 2349 160
rect 2308 156 2314 158
rect 2308 155 2309 156
rect 2303 154 2309 155
rect 2318 155 2324 156
rect 2278 150 2284 151
rect 2318 151 2319 155
rect 2323 151 2324 155
rect 2343 155 2344 159
rect 2348 158 2349 159
rect 2352 158 2354 160
rect 2366 159 2367 160
rect 2371 159 2372 163
rect 2366 158 2372 159
rect 2382 159 2389 160
rect 2348 156 2354 158
rect 2348 155 2349 156
rect 2343 154 2349 155
rect 2358 155 2364 156
rect 2318 150 2324 151
rect 2358 151 2359 155
rect 2363 151 2364 155
rect 2382 155 2383 159
rect 2388 155 2389 159
rect 2382 154 2389 155
rect 2358 150 2364 151
rect 446 147 452 148
rect 446 146 447 147
rect 417 144 447 146
rect 175 143 184 144
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 175 139 176 143
rect 183 139 184 143
rect 215 143 224 144
rect 175 138 184 139
rect 190 139 196 140
rect 150 134 156 135
rect 190 135 191 139
rect 195 135 196 139
rect 215 139 216 143
rect 223 139 224 143
rect 255 143 264 144
rect 215 138 224 139
rect 230 139 236 140
rect 190 134 196 135
rect 230 135 231 139
rect 235 135 236 139
rect 255 139 256 143
rect 263 139 264 143
rect 295 143 304 144
rect 255 138 264 139
rect 270 139 276 140
rect 230 134 236 135
rect 270 135 271 139
rect 275 135 276 139
rect 295 139 296 143
rect 303 139 304 143
rect 335 143 344 144
rect 295 138 304 139
rect 310 139 316 140
rect 270 134 276 135
rect 310 135 311 139
rect 315 135 316 139
rect 335 139 336 143
rect 343 139 344 143
rect 375 143 384 144
rect 335 138 344 139
rect 350 139 356 140
rect 310 134 316 135
rect 350 135 351 139
rect 355 135 356 139
rect 375 139 376 143
rect 383 139 384 143
rect 415 143 421 144
rect 375 138 384 139
rect 390 139 396 140
rect 350 134 356 135
rect 390 135 391 139
rect 395 135 396 139
rect 415 139 416 143
rect 420 139 421 143
rect 446 143 447 144
rect 451 143 452 147
rect 1166 147 1172 148
rect 1166 146 1167 147
rect 1144 144 1167 146
rect 446 142 452 143
rect 455 143 464 144
rect 415 138 421 139
rect 430 139 436 140
rect 390 134 396 135
rect 430 135 431 139
rect 435 135 436 139
rect 455 139 456 143
rect 463 139 464 143
rect 495 143 504 144
rect 455 138 464 139
rect 470 139 476 140
rect 430 134 436 135
rect 470 135 471 139
rect 475 135 476 139
rect 495 139 496 143
rect 503 139 504 143
rect 535 143 544 144
rect 495 138 504 139
rect 510 139 516 140
rect 470 134 476 135
rect 510 135 511 139
rect 515 135 516 139
rect 535 139 536 143
rect 543 139 544 143
rect 575 143 584 144
rect 535 138 544 139
rect 550 139 556 140
rect 510 134 516 135
rect 550 135 551 139
rect 555 135 556 139
rect 575 139 576 143
rect 583 139 584 143
rect 614 143 621 144
rect 575 138 584 139
rect 590 139 596 140
rect 550 134 556 135
rect 590 135 591 139
rect 595 135 596 139
rect 614 139 615 143
rect 620 139 621 143
rect 655 143 664 144
rect 614 138 621 139
rect 630 139 636 140
rect 590 134 596 135
rect 630 135 631 139
rect 635 135 636 139
rect 655 139 656 143
rect 663 139 664 143
rect 695 143 704 144
rect 655 138 664 139
rect 670 139 676 140
rect 630 134 636 135
rect 670 135 671 139
rect 675 135 676 139
rect 695 139 696 143
rect 703 139 704 143
rect 735 143 744 144
rect 695 138 704 139
rect 710 139 716 140
rect 670 134 676 135
rect 710 135 711 139
rect 715 135 716 139
rect 735 139 736 143
rect 743 139 744 143
rect 775 143 784 144
rect 735 138 744 139
rect 750 139 756 140
rect 710 134 716 135
rect 750 135 751 139
rect 755 135 756 139
rect 775 139 776 143
rect 783 139 784 143
rect 815 143 824 144
rect 775 138 784 139
rect 790 139 796 140
rect 750 134 756 135
rect 790 135 791 139
rect 795 135 796 139
rect 815 139 816 143
rect 823 139 824 143
rect 855 143 864 144
rect 815 138 824 139
rect 830 139 836 140
rect 790 134 796 135
rect 830 135 831 139
rect 835 135 836 139
rect 855 139 856 143
rect 863 139 864 143
rect 895 143 904 144
rect 855 138 864 139
rect 870 139 876 140
rect 830 134 836 135
rect 870 135 871 139
rect 875 135 876 139
rect 895 139 896 143
rect 903 139 904 143
rect 935 143 944 144
rect 895 138 904 139
rect 910 139 916 140
rect 870 134 876 135
rect 910 135 911 139
rect 915 135 916 139
rect 935 139 936 143
rect 943 139 944 143
rect 975 143 984 144
rect 935 138 944 139
rect 950 139 956 140
rect 910 134 916 135
rect 950 135 951 139
rect 955 135 956 139
rect 975 139 976 143
rect 983 139 984 143
rect 1015 143 1024 144
rect 975 138 984 139
rect 990 139 996 140
rect 950 134 956 135
rect 990 135 991 139
rect 995 135 996 139
rect 1015 139 1016 143
rect 1023 139 1024 143
rect 1055 143 1064 144
rect 1015 138 1024 139
rect 1030 139 1036 140
rect 990 134 996 135
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1055 139 1056 143
rect 1063 139 1064 143
rect 1095 143 1104 144
rect 1055 138 1064 139
rect 1070 139 1076 140
rect 1030 134 1036 135
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1095 139 1096 143
rect 1103 139 1104 143
rect 1135 143 1141 144
rect 1095 138 1104 139
rect 1110 139 1116 140
rect 1070 134 1076 135
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1135 139 1136 143
rect 1140 142 1141 143
rect 1144 142 1146 144
rect 1166 143 1167 144
rect 1171 143 1172 147
rect 1198 147 1204 148
rect 1198 146 1199 147
rect 1184 144 1199 146
rect 1166 142 1172 143
rect 1175 143 1181 144
rect 1140 140 1146 142
rect 1140 139 1141 140
rect 1135 138 1141 139
rect 1150 139 1156 140
rect 1110 134 1116 135
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1175 139 1176 143
rect 1180 142 1181 143
rect 1184 142 1186 144
rect 1198 143 1199 144
rect 1203 143 1204 147
rect 1198 142 1204 143
rect 1215 143 1221 144
rect 1180 140 1186 142
rect 1180 139 1181 140
rect 1175 138 1181 139
rect 1190 139 1196 140
rect 1150 134 1156 135
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1215 139 1216 143
rect 1220 142 1221 143
rect 1220 140 1290 142
rect 1220 139 1221 140
rect 1215 138 1221 139
rect 1190 134 1196 135
rect 1278 132 1284 133
rect 1278 128 1279 132
rect 1283 128 1284 132
rect 1278 127 1284 128
rect 1288 126 1290 140
rect 1962 135 1968 136
rect 1962 131 1963 135
rect 1967 134 1968 135
rect 1967 132 2001 134
rect 1967 131 1968 132
rect 1962 130 1968 131
rect 1999 128 2001 132
rect 2406 132 2412 133
rect 2406 128 2407 132
rect 2411 128 2412 132
rect 1327 127 1333 128
rect 1327 126 1328 127
rect 1288 124 1328 126
rect 1327 123 1328 124
rect 1332 123 1333 127
rect 1327 122 1333 123
rect 1338 127 1344 128
rect 1338 123 1339 127
rect 1343 126 1344 127
rect 1367 127 1373 128
rect 1367 126 1368 127
rect 1343 124 1368 126
rect 1343 123 1344 124
rect 1338 122 1344 123
rect 1367 123 1368 124
rect 1372 123 1373 127
rect 1367 122 1373 123
rect 1378 127 1384 128
rect 1378 123 1379 127
rect 1383 126 1384 127
rect 1407 127 1413 128
rect 1407 126 1408 127
rect 1383 124 1408 126
rect 1383 123 1384 124
rect 1378 122 1384 123
rect 1407 123 1408 124
rect 1412 123 1413 127
rect 1407 122 1413 123
rect 1418 127 1424 128
rect 1418 123 1419 127
rect 1423 126 1424 127
rect 1447 127 1453 128
rect 1447 126 1448 127
rect 1423 124 1448 126
rect 1423 123 1424 124
rect 1418 122 1424 123
rect 1447 123 1448 124
rect 1452 123 1453 127
rect 1447 122 1453 123
rect 1458 127 1464 128
rect 1458 123 1459 127
rect 1463 126 1464 127
rect 1487 127 1493 128
rect 1487 126 1488 127
rect 1463 124 1488 126
rect 1463 123 1464 124
rect 1458 122 1464 123
rect 1487 123 1488 124
rect 1492 123 1493 127
rect 1487 122 1493 123
rect 1510 127 1516 128
rect 1510 123 1511 127
rect 1515 126 1516 127
rect 1543 127 1549 128
rect 1543 126 1544 127
rect 1515 124 1544 126
rect 1515 123 1516 124
rect 1510 122 1516 123
rect 1543 123 1544 124
rect 1548 123 1549 127
rect 1543 122 1549 123
rect 1574 127 1580 128
rect 1574 123 1575 127
rect 1579 126 1580 127
rect 1607 127 1613 128
rect 1607 126 1608 127
rect 1579 124 1608 126
rect 1579 123 1580 124
rect 1574 122 1580 123
rect 1607 123 1608 124
rect 1612 123 1613 127
rect 1607 122 1613 123
rect 1638 127 1644 128
rect 1638 123 1639 127
rect 1643 126 1644 127
rect 1671 127 1677 128
rect 1671 126 1672 127
rect 1643 124 1672 126
rect 1643 123 1644 124
rect 1638 122 1644 123
rect 1671 123 1672 124
rect 1676 123 1677 127
rect 1671 122 1677 123
rect 1735 127 1744 128
rect 1735 123 1736 127
rect 1743 123 1744 127
rect 1735 122 1744 123
rect 1766 127 1772 128
rect 1766 123 1767 127
rect 1771 126 1772 127
rect 1799 127 1805 128
rect 1799 126 1800 127
rect 1771 124 1800 126
rect 1771 123 1772 124
rect 1766 122 1772 123
rect 1799 123 1800 124
rect 1804 123 1805 127
rect 1799 122 1805 123
rect 1822 127 1828 128
rect 1822 123 1823 127
rect 1827 126 1828 127
rect 1855 127 1861 128
rect 1855 126 1856 127
rect 1827 124 1856 126
rect 1827 123 1828 124
rect 1822 122 1828 123
rect 1855 123 1856 124
rect 1860 123 1861 127
rect 1855 122 1861 123
rect 1878 127 1884 128
rect 1878 123 1879 127
rect 1883 126 1884 127
rect 1911 127 1917 128
rect 1911 126 1912 127
rect 1883 124 1912 126
rect 1883 123 1884 124
rect 1878 122 1884 123
rect 1911 123 1912 124
rect 1916 123 1917 127
rect 1911 122 1917 123
rect 1926 127 1932 128
rect 1926 123 1927 127
rect 1931 126 1932 127
rect 1959 127 1965 128
rect 1959 126 1960 127
rect 1931 124 1960 126
rect 1931 123 1932 124
rect 1926 122 1932 123
rect 1959 123 1960 124
rect 1964 123 1965 127
rect 1959 122 1965 123
rect 1999 127 2005 128
rect 1999 123 2000 127
rect 2004 123 2005 127
rect 1999 122 2005 123
rect 2022 127 2028 128
rect 2022 123 2023 127
rect 2027 126 2028 127
rect 2039 127 2045 128
rect 2039 126 2040 127
rect 2027 124 2040 126
rect 2027 123 2028 124
rect 2022 122 2028 123
rect 2039 123 2040 124
rect 2044 123 2045 127
rect 2039 122 2045 123
rect 2070 127 2076 128
rect 2070 123 2071 127
rect 2075 126 2076 127
rect 2079 127 2085 128
rect 2079 126 2080 127
rect 2075 124 2080 126
rect 2075 123 2076 124
rect 2070 122 2076 123
rect 2079 123 2080 124
rect 2084 123 2085 127
rect 2079 122 2085 123
rect 2102 127 2108 128
rect 2102 123 2103 127
rect 2107 126 2108 127
rect 2119 127 2125 128
rect 2119 126 2120 127
rect 2107 124 2120 126
rect 2107 123 2108 124
rect 2102 122 2108 123
rect 2119 123 2120 124
rect 2124 123 2125 127
rect 2119 122 2125 123
rect 2134 127 2140 128
rect 2134 123 2135 127
rect 2139 126 2140 127
rect 2167 127 2173 128
rect 2167 126 2168 127
rect 2139 124 2168 126
rect 2139 123 2140 124
rect 2134 122 2140 123
rect 2167 123 2168 124
rect 2172 123 2173 127
rect 2167 122 2173 123
rect 2182 127 2188 128
rect 2182 123 2183 127
rect 2187 126 2188 127
rect 2215 127 2221 128
rect 2215 126 2216 127
rect 2187 124 2216 126
rect 2187 123 2188 124
rect 2182 122 2188 123
rect 2215 123 2216 124
rect 2220 123 2221 127
rect 2215 122 2221 123
rect 2262 127 2269 128
rect 2262 123 2263 127
rect 2268 123 2269 127
rect 2262 122 2269 123
rect 2286 127 2292 128
rect 2286 123 2287 127
rect 2291 126 2292 127
rect 2303 127 2309 128
rect 2303 126 2304 127
rect 2291 124 2304 126
rect 2291 123 2292 124
rect 2286 122 2292 123
rect 2303 123 2304 124
rect 2308 123 2309 127
rect 2303 122 2309 123
rect 2334 127 2340 128
rect 2334 123 2335 127
rect 2339 126 2340 127
rect 2343 127 2349 128
rect 2343 126 2344 127
rect 2339 124 2344 126
rect 2339 123 2340 124
rect 2334 122 2340 123
rect 2343 123 2344 124
rect 2348 123 2349 127
rect 2343 122 2349 123
rect 2366 127 2372 128
rect 2366 123 2367 127
rect 2371 126 2372 127
rect 2383 127 2389 128
rect 2406 127 2412 128
rect 2383 126 2384 127
rect 2371 124 2384 126
rect 2371 123 2372 124
rect 2366 122 2372 123
rect 2383 123 2384 124
rect 2388 123 2389 127
rect 2383 122 2389 123
rect 298 119 304 120
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 298 115 299 119
rect 303 118 304 119
rect 303 116 321 118
rect 303 115 304 116
rect 298 114 304 115
rect 110 111 116 112
rect 178 111 184 112
rect 178 107 179 111
rect 183 110 184 111
rect 215 111 221 112
rect 215 110 216 111
rect 183 108 216 110
rect 183 107 184 108
rect 178 106 184 107
rect 215 107 216 108
rect 220 107 221 111
rect 215 106 221 107
rect 226 111 232 112
rect 226 107 227 111
rect 231 110 232 111
rect 255 111 261 112
rect 255 110 256 111
rect 231 108 256 110
rect 231 107 232 108
rect 226 106 232 107
rect 255 107 256 108
rect 260 107 261 111
rect 255 106 261 107
rect 266 111 272 112
rect 266 107 267 111
rect 271 110 272 111
rect 295 111 301 112
rect 295 110 296 111
rect 271 108 296 110
rect 271 107 272 108
rect 266 106 272 107
rect 295 107 296 108
rect 300 107 301 111
rect 319 110 321 116
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 335 111 341 112
rect 335 110 336 111
rect 319 108 336 110
rect 295 106 301 107
rect 335 107 336 108
rect 340 107 341 111
rect 335 106 341 107
rect 346 111 352 112
rect 346 107 347 111
rect 351 110 352 111
rect 375 111 381 112
rect 375 110 376 111
rect 351 108 376 110
rect 351 107 352 108
rect 346 106 352 107
rect 375 107 376 108
rect 380 107 381 111
rect 375 106 381 107
rect 386 111 392 112
rect 386 107 387 111
rect 391 110 392 111
rect 415 111 421 112
rect 415 110 416 111
rect 391 108 416 110
rect 391 107 392 108
rect 386 106 392 107
rect 415 107 416 108
rect 420 107 421 111
rect 415 106 421 107
rect 446 111 452 112
rect 446 107 447 111
rect 451 110 452 111
rect 455 111 461 112
rect 455 110 456 111
rect 451 108 456 110
rect 451 107 452 108
rect 446 106 452 107
rect 455 107 456 108
rect 460 107 461 111
rect 455 106 461 107
rect 466 111 472 112
rect 466 107 467 111
rect 471 110 472 111
rect 495 111 501 112
rect 495 110 496 111
rect 471 108 496 110
rect 471 107 472 108
rect 466 106 472 107
rect 495 107 496 108
rect 500 107 501 111
rect 495 106 501 107
rect 506 111 512 112
rect 506 107 507 111
rect 511 110 512 111
rect 535 111 541 112
rect 535 110 536 111
rect 511 108 536 110
rect 511 107 512 108
rect 506 106 512 107
rect 535 107 536 108
rect 540 107 541 111
rect 535 106 541 107
rect 546 111 552 112
rect 546 107 547 111
rect 551 110 552 111
rect 575 111 581 112
rect 575 110 576 111
rect 551 108 576 110
rect 551 107 552 108
rect 546 106 552 107
rect 575 107 576 108
rect 580 107 581 111
rect 575 106 581 107
rect 586 111 592 112
rect 586 107 587 111
rect 591 110 592 111
rect 615 111 621 112
rect 615 110 616 111
rect 591 108 616 110
rect 591 107 592 108
rect 586 106 592 107
rect 615 107 616 108
rect 620 107 621 111
rect 615 106 621 107
rect 650 111 661 112
rect 650 107 651 111
rect 655 107 656 111
rect 660 107 661 111
rect 650 106 661 107
rect 666 111 672 112
rect 666 107 667 111
rect 671 110 672 111
rect 695 111 701 112
rect 695 110 696 111
rect 671 108 696 110
rect 671 107 672 108
rect 666 106 672 107
rect 695 107 696 108
rect 700 107 701 111
rect 695 106 701 107
rect 706 111 712 112
rect 706 107 707 111
rect 711 110 712 111
rect 735 111 741 112
rect 735 110 736 111
rect 711 108 736 110
rect 711 107 712 108
rect 706 106 712 107
rect 735 107 736 108
rect 740 107 741 111
rect 735 106 741 107
rect 746 111 752 112
rect 746 107 747 111
rect 751 110 752 111
rect 775 111 781 112
rect 775 110 776 111
rect 751 108 776 110
rect 751 107 752 108
rect 746 106 752 107
rect 775 107 776 108
rect 780 107 781 111
rect 775 106 781 107
rect 786 111 792 112
rect 786 107 787 111
rect 791 110 792 111
rect 815 111 821 112
rect 815 110 816 111
rect 791 108 816 110
rect 791 107 792 108
rect 786 106 792 107
rect 815 107 816 108
rect 820 107 821 111
rect 815 106 821 107
rect 826 111 832 112
rect 826 107 827 111
rect 831 110 832 111
rect 855 111 861 112
rect 855 110 856 111
rect 831 108 856 110
rect 831 107 832 108
rect 826 106 832 107
rect 855 107 856 108
rect 860 107 861 111
rect 855 106 861 107
rect 866 111 872 112
rect 866 107 867 111
rect 871 110 872 111
rect 895 111 901 112
rect 895 110 896 111
rect 871 108 896 110
rect 871 107 872 108
rect 866 106 872 107
rect 895 107 896 108
rect 900 107 901 111
rect 895 106 901 107
rect 906 111 912 112
rect 906 107 907 111
rect 911 110 912 111
rect 935 111 941 112
rect 935 110 936 111
rect 911 108 936 110
rect 911 107 912 108
rect 906 106 912 107
rect 935 107 936 108
rect 940 107 941 111
rect 935 106 941 107
rect 946 111 952 112
rect 946 107 947 111
rect 951 110 952 111
rect 975 111 981 112
rect 975 110 976 111
rect 951 108 976 110
rect 951 107 952 108
rect 946 106 952 107
rect 975 107 976 108
rect 980 107 981 111
rect 975 106 981 107
rect 986 111 992 112
rect 986 107 987 111
rect 991 110 992 111
rect 1015 111 1021 112
rect 1015 110 1016 111
rect 991 108 1016 110
rect 991 107 992 108
rect 986 106 992 107
rect 1015 107 1016 108
rect 1020 107 1021 111
rect 1015 106 1021 107
rect 1026 111 1032 112
rect 1026 107 1027 111
rect 1031 110 1032 111
rect 1055 111 1061 112
rect 1055 110 1056 111
rect 1031 108 1056 110
rect 1031 107 1032 108
rect 1026 106 1032 107
rect 1055 107 1056 108
rect 1060 107 1061 111
rect 1055 106 1061 107
rect 1066 111 1072 112
rect 1066 107 1067 111
rect 1071 110 1072 111
rect 1095 111 1101 112
rect 1095 110 1096 111
rect 1071 108 1096 110
rect 1071 107 1072 108
rect 1066 106 1072 107
rect 1095 107 1096 108
rect 1100 107 1101 111
rect 1095 106 1101 107
rect 1106 111 1112 112
rect 1106 107 1107 111
rect 1111 110 1112 111
rect 1135 111 1141 112
rect 1135 110 1136 111
rect 1111 108 1136 110
rect 1111 107 1112 108
rect 1106 106 1112 107
rect 1135 107 1136 108
rect 1140 107 1141 111
rect 1135 106 1141 107
rect 1166 111 1172 112
rect 1166 107 1167 111
rect 1171 110 1172 111
rect 1175 111 1181 112
rect 1175 110 1176 111
rect 1171 108 1176 110
rect 1171 107 1172 108
rect 1166 106 1172 107
rect 1175 107 1176 108
rect 1180 107 1181 111
rect 1175 106 1181 107
rect 1198 111 1204 112
rect 1198 107 1199 111
rect 1203 110 1204 111
rect 1215 111 1221 112
rect 1238 111 1244 112
rect 1278 115 1284 116
rect 1278 111 1279 115
rect 1283 111 1284 115
rect 1215 110 1216 111
rect 1203 108 1216 110
rect 1203 107 1204 108
rect 1198 106 1204 107
rect 1215 107 1216 108
rect 1220 107 1221 111
rect 1278 110 1284 111
rect 2406 115 2412 116
rect 2406 111 2407 115
rect 2411 111 2412 115
rect 2406 110 2412 111
rect 1215 106 1221 107
rect 1302 108 1308 109
rect 1302 104 1303 108
rect 1307 104 1308 108
rect 1302 103 1308 104
rect 1342 108 1348 109
rect 1342 104 1343 108
rect 1347 104 1348 108
rect 1342 103 1348 104
rect 1382 108 1388 109
rect 1382 104 1383 108
rect 1387 104 1388 108
rect 1382 103 1388 104
rect 1422 108 1428 109
rect 1422 104 1423 108
rect 1427 104 1428 108
rect 1422 103 1428 104
rect 1462 108 1468 109
rect 1462 104 1463 108
rect 1467 104 1468 108
rect 1462 103 1468 104
rect 1518 108 1524 109
rect 1518 104 1519 108
rect 1523 104 1524 108
rect 1518 103 1524 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1646 108 1652 109
rect 1646 104 1647 108
rect 1651 104 1652 108
rect 1646 103 1652 104
rect 1710 108 1716 109
rect 1710 104 1711 108
rect 1715 104 1716 108
rect 1710 103 1716 104
rect 1774 108 1780 109
rect 1774 104 1775 108
rect 1779 104 1780 108
rect 1774 103 1780 104
rect 1830 108 1836 109
rect 1830 104 1831 108
rect 1835 104 1836 108
rect 1830 103 1836 104
rect 1886 108 1892 109
rect 1886 104 1887 108
rect 1891 104 1892 108
rect 1886 103 1892 104
rect 1934 108 1940 109
rect 1934 104 1935 108
rect 1939 104 1940 108
rect 1934 103 1940 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2014 108 2020 109
rect 2014 104 2015 108
rect 2019 104 2020 108
rect 2014 103 2020 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2094 108 2100 109
rect 2094 104 2095 108
rect 2099 104 2100 108
rect 2094 103 2100 104
rect 2142 108 2148 109
rect 2142 104 2143 108
rect 2147 104 2148 108
rect 2142 103 2148 104
rect 2190 108 2196 109
rect 2190 104 2191 108
rect 2195 104 2196 108
rect 2190 103 2196 104
rect 2238 108 2244 109
rect 2238 104 2239 108
rect 2243 104 2244 108
rect 2238 103 2244 104
rect 2278 108 2284 109
rect 2278 104 2279 108
rect 2283 104 2284 108
rect 2278 103 2284 104
rect 2318 108 2324 109
rect 2318 104 2319 108
rect 2323 104 2324 108
rect 2318 103 2324 104
rect 2358 108 2364 109
rect 2358 104 2359 108
rect 2363 104 2364 108
rect 2358 103 2364 104
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1238 94 1244 95
rect 150 92 156 93
rect 150 88 151 92
rect 155 88 156 92
rect 150 87 156 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 270 92 276 93
rect 270 88 271 92
rect 275 88 276 92
rect 270 87 276 88
rect 310 92 316 93
rect 310 88 311 92
rect 315 88 316 92
rect 310 87 316 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 390 92 396 93
rect 390 88 391 92
rect 395 88 396 92
rect 390 87 396 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 510 87 516 88
rect 550 92 556 93
rect 550 88 551 92
rect 555 88 556 92
rect 550 87 556 88
rect 590 92 596 93
rect 590 88 591 92
rect 595 88 596 92
rect 590 87 596 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 710 92 716 93
rect 710 88 711 92
rect 715 88 716 92
rect 710 87 716 88
rect 750 92 756 93
rect 750 88 751 92
rect 755 88 756 92
rect 750 87 756 88
rect 790 92 796 93
rect 790 88 791 92
rect 795 88 796 92
rect 790 87 796 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 910 92 916 93
rect 910 88 911 92
rect 915 88 916 92
rect 910 87 916 88
rect 950 92 956 93
rect 950 88 951 92
rect 955 88 956 92
rect 950 87 956 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1030 92 1036 93
rect 1030 88 1031 92
rect 1035 88 1036 92
rect 1030 87 1036 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
<< m3c >>
rect 231 2475 235 2479
rect 259 2479 260 2483
rect 260 2479 263 2483
rect 271 2475 275 2479
rect 327 2483 331 2487
rect 311 2475 315 2479
rect 359 2483 363 2487
rect 351 2475 355 2479
rect 391 2479 395 2483
rect 399 2475 403 2479
rect 447 2479 451 2483
rect 455 2475 459 2479
rect 503 2479 507 2483
rect 511 2475 515 2479
rect 567 2479 571 2483
rect 575 2475 579 2479
rect 631 2479 635 2483
rect 639 2475 643 2479
rect 651 2479 655 2483
rect 703 2475 707 2479
rect 783 2483 787 2487
rect 767 2475 771 2479
rect 815 2479 819 2483
rect 823 2475 827 2479
rect 871 2479 875 2483
rect 879 2475 883 2479
rect 919 2479 923 2483
rect 927 2475 931 2479
rect 967 2479 971 2483
rect 975 2475 979 2479
rect 1015 2479 1019 2483
rect 1023 2475 1027 2479
rect 1063 2479 1067 2483
rect 1071 2475 1075 2479
rect 1127 2483 1131 2487
rect 1111 2475 1115 2479
rect 1167 2483 1171 2487
rect 1151 2475 1155 2479
rect 1203 2483 1207 2487
rect 1191 2475 1195 2479
rect 1319 2479 1323 2483
rect 1303 2471 1307 2475
rect 1359 2479 1363 2483
rect 1343 2471 1347 2475
rect 1399 2479 1403 2483
rect 1383 2471 1387 2475
rect 1431 2475 1435 2479
rect 1439 2471 1443 2475
rect 1503 2475 1507 2479
rect 1511 2471 1515 2475
rect 1575 2475 1579 2479
rect 1583 2471 1587 2475
rect 1655 2475 1659 2479
rect 1663 2471 1667 2475
rect 1687 2475 1688 2479
rect 1688 2475 1691 2479
rect 1735 2471 1739 2475
rect 1799 2475 1803 2479
rect 1807 2471 1811 2475
rect 1879 2475 1883 2479
rect 1887 2471 1891 2475
rect 1959 2475 1963 2479
rect 1967 2471 1971 2475
rect 2063 2471 2067 2475
rect 2159 2475 2163 2479
rect 2167 2471 2171 2475
rect 2263 2475 2267 2479
rect 2271 2471 2275 2475
rect 2287 2475 2291 2479
rect 2359 2471 2363 2475
rect 111 2452 115 2456
rect 1239 2452 1243 2456
rect 243 2447 247 2451
rect 267 2447 271 2451
rect 327 2447 331 2451
rect 359 2447 363 2451
rect 391 2447 395 2451
rect 447 2447 451 2451
rect 503 2447 507 2451
rect 567 2447 571 2451
rect 631 2447 635 2451
rect 775 2447 779 2451
rect 783 2447 787 2451
rect 815 2447 819 2451
rect 871 2447 875 2451
rect 919 2447 923 2451
rect 967 2447 971 2451
rect 1015 2447 1019 2451
rect 1063 2447 1067 2451
rect 1127 2447 1131 2451
rect 1167 2447 1171 2451
rect 1203 2447 1207 2451
rect 1279 2448 1283 2452
rect 2407 2448 2411 2452
rect 1319 2443 1323 2447
rect 1359 2443 1363 2447
rect 1399 2443 1403 2447
rect 1431 2443 1435 2447
rect 1503 2443 1507 2447
rect 1575 2443 1579 2447
rect 1655 2443 1659 2447
rect 111 2435 115 2439
rect 1239 2435 1243 2439
rect 1799 2443 1803 2447
rect 1879 2443 1883 2447
rect 1959 2443 1963 2447
rect 2159 2443 2163 2447
rect 2263 2443 2267 2447
rect 2383 2443 2384 2447
rect 2384 2443 2387 2447
rect 231 2428 235 2432
rect 271 2428 275 2432
rect 311 2428 315 2432
rect 351 2428 355 2432
rect 399 2428 403 2432
rect 455 2428 459 2432
rect 511 2428 515 2432
rect 575 2428 579 2432
rect 639 2428 643 2432
rect 703 2428 707 2432
rect 767 2428 771 2432
rect 823 2428 827 2432
rect 879 2428 883 2432
rect 927 2428 931 2432
rect 975 2428 979 2432
rect 1023 2428 1027 2432
rect 1071 2428 1075 2432
rect 1111 2428 1115 2432
rect 1151 2428 1155 2432
rect 1191 2428 1195 2432
rect 1279 2431 1283 2435
rect 1975 2435 1979 2439
rect 2407 2431 2411 2435
rect 1303 2424 1307 2428
rect 1343 2424 1347 2428
rect 1383 2424 1387 2428
rect 1439 2424 1443 2428
rect 1511 2424 1515 2428
rect 1583 2424 1587 2428
rect 1663 2424 1667 2428
rect 1735 2424 1739 2428
rect 1807 2424 1811 2428
rect 1887 2424 1891 2428
rect 1967 2424 1971 2428
rect 2063 2424 2067 2428
rect 2167 2424 2171 2428
rect 2271 2424 2275 2428
rect 2359 2424 2363 2428
rect 199 2408 203 2412
rect 263 2408 267 2412
rect 327 2408 331 2412
rect 399 2408 403 2412
rect 471 2408 475 2412
rect 543 2408 547 2412
rect 615 2408 619 2412
rect 687 2408 691 2412
rect 751 2408 755 2412
rect 823 2408 827 2412
rect 895 2408 899 2412
rect 967 2408 971 2412
rect 1375 2412 1379 2416
rect 1415 2412 1419 2416
rect 1455 2412 1459 2416
rect 1503 2412 1507 2416
rect 1559 2412 1563 2416
rect 1615 2412 1619 2416
rect 1679 2412 1683 2416
rect 1735 2412 1739 2416
rect 1799 2412 1803 2416
rect 1871 2412 1875 2416
rect 1951 2412 1955 2416
rect 2047 2412 2051 2416
rect 2151 2412 2155 2416
rect 2263 2412 2267 2416
rect 2359 2412 2363 2416
rect 111 2401 115 2405
rect 1239 2401 1243 2405
rect 1279 2405 1283 2409
rect 2407 2405 2411 2409
rect 651 2395 655 2399
rect 111 2384 115 2388
rect 279 2387 283 2391
rect 343 2387 347 2391
rect 415 2387 419 2391
rect 423 2387 424 2391
rect 424 2387 427 2391
rect 839 2387 843 2391
rect 907 2387 911 2391
rect 1239 2384 1243 2388
rect 1279 2388 1283 2392
rect 1687 2399 1691 2403
rect 1423 2391 1427 2395
rect 1463 2391 1467 2395
rect 2287 2391 2288 2395
rect 2288 2391 2291 2395
rect 1903 2383 1907 2387
rect 2407 2388 2411 2392
rect 991 2379 995 2383
rect 2287 2383 2291 2387
rect 199 2361 203 2365
rect 263 2361 267 2365
rect 327 2361 331 2365
rect 399 2361 403 2365
rect 471 2361 475 2365
rect 543 2361 547 2365
rect 615 2361 619 2365
rect 687 2361 691 2365
rect 751 2361 755 2365
rect 823 2361 827 2365
rect 895 2361 899 2365
rect 967 2361 971 2365
rect 1375 2365 1379 2369
rect 1415 2365 1419 2369
rect 1455 2365 1459 2369
rect 1503 2365 1507 2369
rect 1559 2365 1563 2369
rect 1615 2365 1619 2369
rect 1679 2365 1683 2369
rect 1735 2365 1739 2369
rect 1799 2365 1803 2369
rect 1871 2365 1875 2369
rect 1951 2365 1955 2369
rect 2047 2365 2051 2369
rect 2151 2365 2155 2369
rect 2263 2365 2267 2369
rect 2359 2365 2363 2369
rect 243 2355 247 2359
rect 279 2355 283 2359
rect 343 2355 347 2359
rect 415 2355 419 2359
rect 735 2355 739 2359
rect 775 2355 776 2359
rect 776 2355 779 2359
rect 839 2355 843 2359
rect 991 2355 992 2359
rect 992 2355 995 2359
rect 1423 2359 1427 2363
rect 1463 2359 1467 2363
rect 1659 2359 1663 2363
rect 1975 2359 1976 2363
rect 1976 2359 1979 2363
rect 2187 2359 2191 2363
rect 2287 2359 2288 2363
rect 2288 2359 2291 2363
rect 2383 2359 2384 2363
rect 2384 2359 2387 2363
rect 271 2327 275 2331
rect 319 2331 323 2335
rect 327 2327 331 2331
rect 391 2331 395 2335
rect 399 2327 403 2331
rect 423 2331 424 2335
rect 424 2331 427 2335
rect 471 2327 475 2331
rect 483 2331 487 2335
rect 551 2327 555 2331
rect 563 2331 567 2335
rect 631 2327 635 2331
rect 671 2331 675 2335
rect 711 2327 715 2331
rect 723 2331 727 2335
rect 783 2327 787 2331
rect 847 2331 851 2335
rect 855 2327 859 2331
rect 907 2331 911 2335
rect 919 2327 923 2331
rect 931 2331 935 2335
rect 991 2327 995 2331
rect 1055 2331 1059 2335
rect 1063 2327 1067 2331
rect 1075 2331 1079 2335
rect 1327 2331 1331 2335
rect 1355 2335 1356 2339
rect 1356 2335 1359 2339
rect 1383 2331 1387 2335
rect 1395 2335 1399 2339
rect 1439 2331 1443 2335
rect 1451 2335 1455 2339
rect 1503 2331 1507 2335
rect 1515 2335 1519 2339
rect 1575 2331 1579 2335
rect 1587 2335 1591 2339
rect 1647 2331 1651 2335
rect 1711 2335 1715 2339
rect 1719 2331 1723 2335
rect 1791 2335 1795 2339
rect 1799 2331 1803 2335
rect 1871 2335 1875 2339
rect 1879 2331 1883 2335
rect 1903 2335 1904 2339
rect 1904 2335 1907 2339
rect 1967 2331 1971 2335
rect 1979 2335 1983 2339
rect 2063 2331 2067 2335
rect 2075 2335 2079 2339
rect 2167 2331 2171 2335
rect 2179 2335 2183 2339
rect 2271 2331 2275 2335
rect 2351 2335 2355 2339
rect 2359 2331 2363 2335
rect 111 2304 115 2308
rect 483 2307 487 2311
rect 319 2299 323 2303
rect 391 2299 395 2303
rect 563 2299 567 2303
rect 579 2299 580 2303
rect 580 2299 583 2303
rect 723 2299 727 2303
rect 735 2299 736 2303
rect 736 2299 739 2303
rect 931 2307 935 2311
rect 847 2299 851 2303
rect 1075 2307 1079 2311
rect 1239 2304 1243 2308
rect 1279 2308 1283 2312
rect 2407 2308 2411 2312
rect 1007 2299 1011 2303
rect 1055 2299 1059 2303
rect 1395 2303 1399 2307
rect 1451 2303 1455 2307
rect 1515 2303 1519 2307
rect 1587 2303 1591 2307
rect 1659 2303 1663 2307
rect 1711 2303 1715 2307
rect 1791 2303 1795 2307
rect 1871 2303 1875 2307
rect 2075 2303 2079 2307
rect 2179 2303 2183 2307
rect 2187 2303 2191 2307
rect 2343 2303 2347 2307
rect 2351 2303 2355 2307
rect 111 2287 115 2291
rect 1239 2287 1243 2291
rect 1279 2291 1283 2295
rect 1791 2295 1795 2299
rect 2407 2291 2411 2295
rect 271 2280 275 2284
rect 327 2280 331 2284
rect 399 2280 403 2284
rect 471 2280 475 2284
rect 551 2280 555 2284
rect 631 2280 635 2284
rect 711 2280 715 2284
rect 783 2280 787 2284
rect 855 2280 859 2284
rect 919 2280 923 2284
rect 991 2280 995 2284
rect 1063 2280 1067 2284
rect 1327 2284 1331 2288
rect 1383 2284 1387 2288
rect 1439 2284 1443 2288
rect 1503 2284 1507 2288
rect 1575 2284 1579 2288
rect 1647 2284 1651 2288
rect 1719 2284 1723 2288
rect 1799 2284 1803 2288
rect 1879 2284 1883 2288
rect 1967 2284 1971 2288
rect 2063 2284 2067 2288
rect 2167 2284 2171 2288
rect 2271 2284 2275 2288
rect 2359 2284 2363 2288
rect 1335 2272 1339 2276
rect 1407 2272 1411 2276
rect 1487 2272 1491 2276
rect 1559 2272 1563 2276
rect 1631 2272 1635 2276
rect 1703 2272 1707 2276
rect 1775 2272 1779 2276
rect 1839 2272 1843 2276
rect 1911 2272 1915 2276
rect 1991 2272 1995 2276
rect 2079 2272 2083 2276
rect 2175 2272 2179 2276
rect 2279 2272 2283 2276
rect 2359 2272 2363 2276
rect 1279 2265 1283 2269
rect 143 2260 147 2264
rect 183 2260 187 2264
rect 223 2260 227 2264
rect 279 2260 283 2264
rect 335 2260 339 2264
rect 407 2260 411 2264
rect 479 2260 483 2264
rect 559 2260 563 2264
rect 647 2260 651 2264
rect 727 2260 731 2264
rect 807 2260 811 2264
rect 887 2260 891 2264
rect 967 2260 971 2264
rect 1047 2260 1051 2264
rect 2407 2265 2411 2269
rect 1127 2260 1131 2264
rect 111 2253 115 2257
rect 1239 2253 1243 2257
rect 1979 2259 1983 2263
rect 1279 2248 1283 2252
rect 1355 2251 1359 2255
rect 1615 2251 1619 2255
rect 1623 2251 1627 2255
rect 2383 2251 2384 2255
rect 2384 2251 2387 2255
rect 2407 2248 2411 2252
rect 111 2236 115 2240
rect 199 2239 203 2243
rect 239 2239 243 2243
rect 295 2239 299 2243
rect 351 2239 355 2243
rect 379 2239 383 2243
rect 387 2239 391 2243
rect 543 2239 547 2243
rect 551 2239 555 2243
rect 671 2239 672 2243
rect 672 2239 675 2243
rect 687 2239 691 2243
rect 1135 2239 1139 2243
rect 1143 2239 1147 2243
rect 1239 2236 1243 2240
rect 1071 2231 1075 2235
rect 1335 2225 1339 2229
rect 1407 2225 1411 2229
rect 1487 2225 1491 2229
rect 1559 2225 1563 2229
rect 1631 2225 1635 2229
rect 1703 2225 1707 2229
rect 1775 2225 1779 2229
rect 1839 2225 1843 2229
rect 1911 2225 1915 2229
rect 1991 2225 1995 2229
rect 2079 2225 2083 2229
rect 2175 2225 2179 2229
rect 2279 2225 2283 2229
rect 2359 2225 2363 2229
rect 1535 2219 1539 2223
rect 1623 2219 1627 2223
rect 1791 2219 1795 2223
rect 2343 2219 2347 2223
rect 143 2213 147 2217
rect 183 2213 187 2217
rect 223 2213 227 2217
rect 279 2213 283 2217
rect 335 2213 339 2217
rect 407 2213 411 2217
rect 479 2213 483 2217
rect 559 2213 563 2217
rect 647 2213 651 2217
rect 727 2213 731 2217
rect 807 2213 811 2217
rect 887 2213 891 2217
rect 967 2213 971 2217
rect 163 2207 167 2211
rect 199 2207 203 2211
rect 239 2207 243 2211
rect 295 2207 299 2211
rect 351 2207 355 2211
rect 379 2207 383 2211
rect 551 2207 555 2211
rect 579 2207 583 2211
rect 687 2207 691 2211
rect 855 2207 859 2211
rect 1007 2211 1011 2215
rect 1047 2213 1051 2217
rect 1127 2213 1131 2217
rect 1071 2207 1072 2211
rect 1072 2207 1075 2211
rect 1135 2207 1139 2211
rect 1859 2211 1863 2215
rect 135 2183 139 2187
rect 199 2187 203 2191
rect 207 2183 211 2187
rect 279 2183 283 2187
rect 351 2187 355 2191
rect 359 2183 363 2187
rect 387 2187 388 2191
rect 388 2187 391 2191
rect 439 2183 443 2187
rect 451 2187 455 2191
rect 519 2183 523 2187
rect 543 2187 544 2191
rect 544 2187 547 2191
rect 599 2183 603 2187
rect 679 2183 683 2187
rect 747 2187 751 2191
rect 759 2183 763 2187
rect 771 2187 775 2191
rect 831 2183 835 2187
rect 843 2187 847 2191
rect 903 2183 907 2187
rect 967 2187 971 2191
rect 975 2183 979 2187
rect 1039 2187 1043 2191
rect 1047 2183 1051 2187
rect 1111 2187 1115 2191
rect 1119 2183 1123 2187
rect 1143 2187 1144 2191
rect 1144 2187 1147 2191
rect 1375 2187 1379 2191
rect 1423 2191 1427 2195
rect 1439 2187 1443 2191
rect 1451 2191 1455 2195
rect 1511 2187 1515 2191
rect 1523 2191 1527 2195
rect 1591 2187 1595 2191
rect 1615 2191 1616 2195
rect 1616 2191 1619 2195
rect 1671 2187 1675 2191
rect 1683 2191 1687 2195
rect 1751 2187 1755 2191
rect 1763 2191 1767 2195
rect 1831 2187 1835 2191
rect 1895 2191 1899 2195
rect 1903 2187 1907 2191
rect 1959 2191 1963 2195
rect 1967 2187 1971 2191
rect 2023 2191 2027 2195
rect 2031 2187 2035 2191
rect 2087 2191 2091 2195
rect 2095 2187 2099 2191
rect 2159 2191 2163 2195
rect 2167 2187 2171 2191
rect 2231 2191 2235 2195
rect 2239 2187 2243 2191
rect 2251 2191 2255 2195
rect 2311 2187 2315 2191
rect 2351 2191 2355 2195
rect 2359 2187 2363 2191
rect 2383 2191 2384 2195
rect 2384 2191 2387 2195
rect 111 2160 115 2164
rect 163 2155 164 2159
rect 164 2155 167 2159
rect 199 2155 203 2159
rect 451 2163 455 2167
rect 1239 2160 1243 2164
rect 1279 2164 1283 2168
rect 2407 2164 2411 2168
rect 351 2155 355 2159
rect 451 2155 455 2159
rect 771 2155 775 2159
rect 843 2155 847 2159
rect 855 2155 856 2159
rect 856 2155 859 2159
rect 967 2155 971 2159
rect 1039 2155 1043 2159
rect 1111 2155 1115 2159
rect 1451 2159 1455 2163
rect 1523 2159 1527 2163
rect 1535 2159 1536 2163
rect 1536 2159 1539 2163
rect 1683 2159 1687 2163
rect 1763 2159 1767 2163
rect 1847 2159 1851 2163
rect 1859 2159 1860 2163
rect 1860 2159 1863 2163
rect 1895 2159 1899 2163
rect 1959 2159 1963 2163
rect 2023 2159 2027 2163
rect 2087 2159 2091 2163
rect 2159 2159 2163 2163
rect 2231 2159 2235 2163
rect 2339 2159 2340 2163
rect 2340 2159 2343 2163
rect 2351 2159 2355 2163
rect 111 2143 115 2147
rect 1071 2147 1075 2151
rect 1239 2143 1243 2147
rect 1279 2147 1283 2151
rect 2407 2147 2411 2151
rect 135 2136 139 2140
rect 207 2136 211 2140
rect 279 2136 283 2140
rect 359 2136 363 2140
rect 439 2136 443 2140
rect 519 2136 523 2140
rect 599 2136 603 2140
rect 679 2136 683 2140
rect 759 2136 763 2140
rect 831 2136 835 2140
rect 903 2136 907 2140
rect 975 2136 979 2140
rect 1047 2136 1051 2140
rect 1119 2136 1123 2140
rect 1375 2140 1379 2144
rect 1439 2140 1443 2144
rect 1511 2140 1515 2144
rect 1591 2140 1595 2144
rect 1671 2140 1675 2144
rect 1751 2140 1755 2144
rect 1831 2140 1835 2144
rect 1903 2140 1907 2144
rect 1967 2140 1971 2144
rect 2031 2140 2035 2144
rect 2095 2140 2099 2144
rect 2167 2140 2171 2144
rect 2239 2140 2243 2144
rect 2311 2140 2315 2144
rect 2359 2140 2363 2144
rect 1399 2128 1403 2132
rect 1439 2128 1443 2132
rect 1495 2128 1499 2132
rect 1567 2128 1571 2132
rect 1647 2128 1651 2132
rect 1735 2128 1739 2132
rect 1823 2128 1827 2132
rect 1911 2128 1915 2132
rect 1999 2128 2003 2132
rect 2087 2128 2091 2132
rect 2175 2128 2179 2132
rect 2271 2128 2275 2132
rect 2359 2128 2363 2132
rect 1279 2121 1283 2125
rect 135 2116 139 2120
rect 191 2116 195 2120
rect 271 2116 275 2120
rect 343 2116 347 2120
rect 415 2116 419 2120
rect 479 2116 483 2120
rect 543 2116 547 2120
rect 607 2116 611 2120
rect 671 2116 675 2120
rect 735 2116 739 2120
rect 791 2116 795 2120
rect 839 2116 843 2120
rect 887 2116 891 2120
rect 935 2116 939 2120
rect 991 2116 995 2120
rect 2407 2121 2411 2125
rect 1047 2116 1051 2120
rect 111 2109 115 2113
rect 1239 2109 1243 2113
rect 1279 2104 1283 2108
rect 1423 2107 1424 2111
rect 1424 2107 1427 2111
rect 1447 2107 1451 2111
rect 1939 2107 1940 2111
rect 1940 2107 1943 2111
rect 1947 2107 1951 2111
rect 2347 2107 2351 2111
rect 2407 2104 2411 2108
rect 111 2092 115 2096
rect 207 2095 211 2099
rect 507 2095 508 2099
rect 508 2095 511 2099
rect 623 2095 627 2099
rect 687 2095 691 2099
rect 699 2095 700 2099
rect 700 2095 703 2099
rect 747 2095 751 2099
rect 1239 2092 1243 2096
rect 499 2087 503 2091
rect 1399 2081 1403 2085
rect 1439 2081 1443 2085
rect 1495 2081 1499 2085
rect 1567 2081 1571 2085
rect 1647 2081 1651 2085
rect 1735 2081 1739 2085
rect 1823 2081 1827 2085
rect 1911 2081 1915 2085
rect 1999 2081 2003 2085
rect 2087 2081 2091 2085
rect 2175 2081 2179 2085
rect 2271 2081 2275 2085
rect 2359 2081 2363 2085
rect 1447 2075 1451 2079
rect 1847 2075 1848 2079
rect 1848 2075 1851 2079
rect 1947 2075 1951 2079
rect 135 2069 139 2073
rect 191 2069 195 2073
rect 271 2069 275 2073
rect 343 2069 347 2073
rect 415 2069 419 2073
rect 159 2063 160 2067
rect 160 2063 163 2067
rect 207 2063 211 2067
rect 451 2067 455 2071
rect 479 2069 483 2073
rect 543 2069 547 2073
rect 607 2069 611 2073
rect 671 2069 675 2073
rect 735 2069 739 2073
rect 791 2069 795 2073
rect 839 2069 843 2073
rect 887 2069 891 2073
rect 935 2069 939 2073
rect 991 2069 995 2073
rect 1047 2069 1051 2073
rect 499 2063 503 2067
rect 623 2063 627 2067
rect 687 2063 691 2067
rect 1071 2063 1072 2067
rect 1072 2063 1075 2067
rect 2107 2067 2111 2071
rect 2339 2075 2343 2079
rect 1943 2059 1947 2063
rect 2039 2051 2043 2055
rect 2079 2051 2083 2055
rect 2091 2055 2095 2059
rect 2119 2051 2123 2055
rect 2147 2055 2148 2059
rect 2148 2055 2151 2059
rect 2159 2051 2163 2055
rect 2207 2059 2211 2063
rect 2199 2051 2203 2055
rect 2255 2059 2259 2063
rect 2239 2051 2243 2055
rect 2267 2055 2268 2059
rect 2268 2055 2271 2059
rect 2279 2051 2283 2055
rect 2295 2055 2299 2059
rect 2319 2051 2323 2055
rect 2347 2055 2348 2059
rect 2348 2055 2351 2059
rect 2359 2051 2363 2055
rect 2371 2055 2375 2059
rect 135 2035 139 2039
rect 183 2043 187 2047
rect 175 2035 179 2039
rect 203 2039 204 2043
rect 204 2039 207 2043
rect 215 2035 219 2039
rect 271 2039 275 2043
rect 279 2035 283 2039
rect 343 2039 347 2043
rect 351 2035 355 2039
rect 415 2039 419 2043
rect 423 2035 427 2039
rect 435 2039 439 2043
rect 487 2035 491 2039
rect 507 2039 511 2043
rect 551 2035 555 2039
rect 563 2039 567 2043
rect 615 2035 619 2039
rect 679 2035 683 2039
rect 699 2039 703 2043
rect 743 2035 747 2039
rect 755 2039 759 2043
rect 815 2035 819 2039
rect 827 2039 831 2043
rect 1279 2028 1283 2032
rect 2147 2031 2151 2035
rect 2267 2031 2271 2035
rect 2407 2028 2411 2032
rect 2091 2023 2095 2027
rect 2107 2023 2108 2027
rect 2108 2023 2111 2027
rect 111 2012 115 2016
rect 755 2015 759 2019
rect 2207 2023 2211 2027
rect 2255 2023 2259 2027
rect 2371 2023 2375 2027
rect 2383 2023 2384 2027
rect 2384 2023 2387 2027
rect 1239 2012 1243 2016
rect 159 2007 160 2011
rect 160 2007 163 2011
rect 183 2007 187 2011
rect 211 2007 215 2011
rect 271 2007 275 2011
rect 343 2007 347 2011
rect 415 2007 419 2011
rect 563 2007 567 2011
rect 603 2007 607 2011
rect 823 2007 827 2011
rect 831 2007 835 2011
rect 1279 2011 1283 2015
rect 2215 2015 2219 2019
rect 2407 2011 2411 2015
rect 2039 2004 2043 2008
rect 2079 2004 2083 2008
rect 2119 2004 2123 2008
rect 2159 2004 2163 2008
rect 2199 2004 2203 2008
rect 2239 2004 2243 2008
rect 2279 2004 2283 2008
rect 2319 2004 2323 2008
rect 2359 2004 2363 2008
rect 111 1995 115 1999
rect 1239 1995 1243 1999
rect 135 1988 139 1992
rect 175 1988 179 1992
rect 215 1988 219 1992
rect 279 1988 283 1992
rect 351 1988 355 1992
rect 423 1988 427 1992
rect 487 1988 491 1992
rect 551 1988 555 1992
rect 615 1988 619 1992
rect 679 1988 683 1992
rect 743 1988 747 1992
rect 815 1988 819 1992
rect 1399 1992 1403 1996
rect 1439 1992 1443 1996
rect 1479 1992 1483 1996
rect 1519 1992 1523 1996
rect 1559 1992 1563 1996
rect 1599 1992 1603 1996
rect 1639 1992 1643 1996
rect 1679 1992 1683 1996
rect 1719 1992 1723 1996
rect 1767 1992 1771 1996
rect 1823 1992 1827 1996
rect 1871 1992 1875 1996
rect 1919 1992 1923 1996
rect 1967 1992 1971 1996
rect 2015 1992 2019 1996
rect 2055 1992 2059 1996
rect 2095 1992 2099 1996
rect 2143 1992 2147 1996
rect 2191 1992 2195 1996
rect 2239 1992 2243 1996
rect 2279 1992 2283 1996
rect 2319 1992 2323 1996
rect 2359 1992 2363 1996
rect 1279 1985 1283 1989
rect 2407 1985 2411 1989
rect 135 1976 139 1980
rect 175 1976 179 1980
rect 215 1976 219 1980
rect 271 1976 275 1980
rect 343 1976 347 1980
rect 415 1976 419 1980
rect 495 1976 499 1980
rect 575 1976 579 1980
rect 647 1976 651 1980
rect 719 1976 723 1980
rect 791 1976 795 1980
rect 863 1976 867 1980
rect 935 1976 939 1980
rect 1007 1976 1011 1980
rect 111 1969 115 1973
rect 1239 1969 1243 1973
rect 1279 1968 1283 1972
rect 435 1963 439 1967
rect 1447 1971 1451 1975
rect 1487 1971 1491 1975
rect 1575 1971 1579 1975
rect 1615 1971 1619 1975
rect 1655 1971 1659 1975
rect 1695 1971 1699 1975
rect 1735 1971 1739 1975
rect 1783 1971 1787 1975
rect 1839 1971 1843 1975
rect 1879 1971 1883 1975
rect 1543 1963 1547 1967
rect 1943 1971 1944 1975
rect 1944 1971 1947 1975
rect 2023 1971 2027 1975
rect 2083 1971 2084 1975
rect 2084 1971 2087 1975
rect 2103 1971 2107 1975
rect 2295 1971 2299 1975
rect 2327 1971 2331 1975
rect 2367 1971 2371 1975
rect 2047 1963 2051 1967
rect 2287 1963 2291 1967
rect 2407 1968 2411 1972
rect 111 1952 115 1956
rect 183 1955 187 1959
rect 223 1955 227 1959
rect 439 1947 443 1951
rect 663 1955 667 1959
rect 683 1955 687 1959
rect 691 1955 695 1959
rect 879 1955 883 1959
rect 951 1955 955 1959
rect 1015 1955 1019 1959
rect 1023 1955 1027 1959
rect 1239 1952 1243 1956
rect 1399 1945 1403 1949
rect 1439 1945 1443 1949
rect 1479 1945 1483 1949
rect 1519 1945 1523 1949
rect 1559 1945 1563 1949
rect 1599 1945 1603 1949
rect 1639 1945 1643 1949
rect 1679 1945 1683 1949
rect 1719 1945 1723 1949
rect 1767 1945 1771 1949
rect 1823 1945 1827 1949
rect 1871 1945 1875 1949
rect 1919 1945 1923 1949
rect 1967 1945 1971 1949
rect 2015 1945 2019 1949
rect 2055 1945 2059 1949
rect 2095 1945 2099 1949
rect 2143 1945 2147 1949
rect 2191 1945 2195 1949
rect 2239 1945 2243 1949
rect 2279 1945 2283 1949
rect 2319 1945 2323 1949
rect 2359 1945 2363 1949
rect 1447 1939 1451 1943
rect 1487 1939 1491 1943
rect 1535 1939 1539 1943
rect 1543 1939 1544 1943
rect 1544 1939 1547 1943
rect 1575 1939 1579 1943
rect 1615 1939 1619 1943
rect 1655 1939 1659 1943
rect 1695 1939 1699 1943
rect 1735 1939 1739 1943
rect 1783 1939 1787 1943
rect 1839 1939 1843 1943
rect 1879 1939 1883 1943
rect 2023 1939 2027 1943
rect 2071 1939 2075 1943
rect 2103 1939 2107 1943
rect 2215 1939 2216 1943
rect 2216 1939 2219 1943
rect 2287 1939 2291 1943
rect 2327 1939 2331 1943
rect 2367 1939 2371 1943
rect 2383 1939 2384 1943
rect 2384 1939 2387 1943
rect 135 1929 139 1933
rect 175 1929 179 1933
rect 215 1929 219 1933
rect 271 1929 275 1933
rect 343 1929 347 1933
rect 415 1929 419 1933
rect 495 1929 499 1933
rect 575 1929 579 1933
rect 647 1929 651 1933
rect 719 1929 723 1933
rect 791 1929 795 1933
rect 863 1929 867 1933
rect 935 1929 939 1933
rect 1007 1929 1011 1933
rect 183 1923 187 1927
rect 223 1923 227 1927
rect 439 1923 440 1927
rect 440 1923 443 1927
rect 295 1915 299 1919
rect 603 1923 604 1927
rect 604 1923 607 1927
rect 663 1923 667 1927
rect 683 1923 687 1927
rect 831 1923 835 1927
rect 879 1923 883 1927
rect 951 1923 955 1927
rect 1015 1923 1019 1927
rect 1343 1911 1347 1915
rect 1371 1915 1372 1919
rect 1372 1915 1375 1919
rect 1383 1911 1387 1915
rect 1395 1915 1399 1919
rect 1423 1911 1427 1915
rect 1435 1915 1439 1919
rect 1463 1911 1467 1915
rect 1475 1915 1479 1919
rect 1511 1911 1515 1915
rect 1559 1915 1563 1919
rect 1567 1911 1571 1915
rect 1623 1915 1627 1919
rect 1631 1911 1635 1915
rect 1643 1915 1647 1919
rect 1711 1911 1715 1915
rect 1799 1915 1803 1919
rect 1807 1911 1811 1915
rect 1911 1915 1915 1919
rect 1919 1911 1923 1915
rect 2023 1915 2027 1919
rect 2031 1911 2035 1915
rect 2047 1915 2051 1919
rect 2083 1919 2087 1923
rect 2151 1911 2155 1915
rect 247 1895 251 1899
rect 303 1903 307 1907
rect 287 1895 291 1899
rect 315 1899 316 1903
rect 316 1899 319 1903
rect 327 1895 331 1899
rect 355 1899 356 1903
rect 356 1899 359 1903
rect 367 1895 371 1899
rect 407 1899 411 1903
rect 415 1895 419 1899
rect 463 1899 467 1903
rect 471 1895 475 1899
rect 527 1899 531 1903
rect 535 1895 539 1899
rect 591 1899 595 1903
rect 599 1895 603 1899
rect 611 1899 615 1903
rect 663 1895 667 1899
rect 691 1899 692 1903
rect 692 1899 695 1903
rect 727 1895 731 1899
rect 739 1899 743 1903
rect 791 1895 795 1899
rect 803 1899 807 1903
rect 855 1895 859 1899
rect 867 1899 871 1903
rect 919 1895 923 1899
rect 975 1899 979 1903
rect 1023 1903 1027 1907
rect 983 1895 987 1899
rect 1055 1895 1059 1899
rect 1119 1899 1123 1903
rect 1127 1895 1131 1899
rect 1139 1899 1143 1903
rect 1279 1888 1283 1892
rect 1395 1883 1399 1887
rect 1435 1883 1439 1887
rect 1475 1883 1479 1887
rect 1643 1891 1647 1895
rect 2407 1888 2411 1892
rect 1535 1883 1536 1887
rect 1536 1883 1539 1887
rect 1559 1883 1563 1887
rect 1623 1883 1627 1887
rect 1799 1883 1803 1887
rect 1911 1883 1915 1887
rect 2023 1883 2027 1887
rect 2071 1883 2075 1887
rect 111 1872 115 1876
rect 295 1871 299 1875
rect 315 1875 319 1879
rect 303 1867 307 1871
rect 363 1867 367 1871
rect 407 1867 411 1871
rect 463 1867 467 1871
rect 527 1867 531 1871
rect 591 1867 595 1871
rect 739 1867 743 1871
rect 803 1867 807 1871
rect 863 1867 867 1871
rect 871 1867 875 1871
rect 1139 1875 1143 1879
rect 1239 1872 1243 1876
rect 975 1867 979 1871
rect 1071 1867 1075 1871
rect 1119 1867 1123 1871
rect 1279 1871 1283 1875
rect 2407 1871 2411 1875
rect 1343 1864 1347 1868
rect 1383 1864 1387 1868
rect 1423 1864 1427 1868
rect 1463 1864 1467 1868
rect 1511 1864 1515 1868
rect 1567 1864 1571 1868
rect 1631 1864 1635 1868
rect 1711 1864 1715 1868
rect 1807 1864 1811 1868
rect 1919 1864 1923 1868
rect 2031 1864 2035 1868
rect 2151 1864 2155 1868
rect 111 1855 115 1859
rect 1239 1855 1243 1859
rect 247 1848 251 1852
rect 287 1848 291 1852
rect 327 1848 331 1852
rect 367 1848 371 1852
rect 415 1848 419 1852
rect 471 1848 475 1852
rect 535 1848 539 1852
rect 599 1848 603 1852
rect 663 1848 667 1852
rect 727 1848 731 1852
rect 791 1848 795 1852
rect 855 1848 859 1852
rect 919 1848 923 1852
rect 983 1848 987 1852
rect 1055 1848 1059 1852
rect 1127 1848 1131 1852
rect 1359 1844 1363 1848
rect 1399 1844 1403 1848
rect 1447 1844 1451 1848
rect 1503 1844 1507 1848
rect 1559 1844 1563 1848
rect 1615 1844 1619 1848
rect 1671 1844 1675 1848
rect 1727 1844 1731 1848
rect 1783 1844 1787 1848
rect 1839 1844 1843 1848
rect 1895 1844 1899 1848
rect 1951 1844 1955 1848
rect 1279 1837 1283 1841
rect 399 1832 403 1836
rect 439 1832 443 1836
rect 479 1832 483 1836
rect 519 1832 523 1836
rect 567 1832 571 1836
rect 623 1832 627 1836
rect 687 1832 691 1836
rect 759 1832 763 1836
rect 831 1832 835 1836
rect 903 1832 907 1836
rect 975 1832 979 1836
rect 1047 1832 1051 1836
rect 1127 1832 1131 1836
rect 2407 1837 2411 1841
rect 1191 1832 1195 1836
rect 111 1825 115 1829
rect 1239 1825 1243 1829
rect 111 1808 115 1812
rect 611 1819 615 1823
rect 1279 1820 1283 1824
rect 1371 1823 1375 1827
rect 1407 1823 1411 1827
rect 1743 1823 1747 1827
rect 1799 1823 1803 1827
rect 1855 1823 1859 1827
rect 1903 1823 1907 1827
rect 2407 1820 2411 1824
rect 447 1811 451 1815
rect 487 1811 491 1815
rect 527 1811 531 1815
rect 959 1811 963 1815
rect 1207 1811 1211 1815
rect 1975 1815 1979 1819
rect 927 1803 931 1807
rect 1151 1803 1155 1807
rect 1171 1803 1175 1807
rect 1239 1808 1243 1812
rect 1359 1797 1363 1801
rect 1399 1797 1403 1801
rect 1447 1797 1451 1801
rect 1503 1797 1507 1801
rect 1559 1797 1563 1801
rect 1615 1797 1619 1801
rect 1671 1797 1675 1801
rect 1727 1797 1731 1801
rect 1783 1797 1787 1801
rect 1839 1797 1843 1801
rect 1895 1797 1899 1801
rect 1951 1797 1955 1801
rect 1407 1791 1411 1795
rect 1603 1791 1607 1795
rect 1743 1791 1747 1795
rect 1799 1791 1803 1795
rect 1855 1791 1859 1795
rect 1975 1791 1976 1795
rect 1976 1791 1979 1795
rect 399 1785 403 1789
rect 439 1785 443 1789
rect 479 1785 483 1789
rect 519 1785 523 1789
rect 567 1785 571 1789
rect 623 1785 627 1789
rect 687 1785 691 1789
rect 759 1785 763 1789
rect 831 1785 835 1789
rect 447 1779 451 1783
rect 487 1779 491 1783
rect 527 1779 531 1783
rect 675 1779 679 1783
rect 871 1783 875 1787
rect 903 1785 907 1789
rect 975 1785 979 1789
rect 1047 1785 1051 1789
rect 1127 1785 1131 1789
rect 1191 1785 1195 1789
rect 927 1779 928 1783
rect 928 1779 931 1783
rect 1071 1779 1072 1783
rect 1072 1779 1075 1783
rect 1151 1779 1152 1783
rect 1152 1779 1155 1783
rect 1207 1779 1211 1783
rect 407 1755 411 1759
rect 435 1759 436 1763
rect 436 1759 439 1763
rect 447 1755 451 1759
rect 459 1759 463 1763
rect 487 1755 491 1759
rect 499 1759 503 1763
rect 527 1755 531 1759
rect 539 1759 543 1763
rect 567 1755 571 1759
rect 579 1759 583 1763
rect 607 1755 611 1759
rect 619 1759 623 1763
rect 647 1755 651 1759
rect 659 1759 663 1763
rect 695 1755 699 1759
rect 743 1759 747 1763
rect 751 1755 755 1759
rect 799 1759 803 1763
rect 807 1755 811 1759
rect 863 1759 867 1763
rect 871 1755 875 1759
rect 927 1759 931 1763
rect 935 1755 939 1759
rect 959 1759 960 1763
rect 960 1759 963 1763
rect 999 1755 1003 1759
rect 1071 1755 1075 1759
rect 1127 1759 1131 1763
rect 1143 1755 1147 1759
rect 1171 1759 1172 1763
rect 1172 1759 1175 1763
rect 1191 1755 1195 1759
rect 1203 1759 1207 1763
rect 1303 1755 1307 1759
rect 1315 1759 1319 1763
rect 1343 1755 1347 1759
rect 1355 1759 1359 1763
rect 1391 1755 1395 1759
rect 1447 1759 1451 1763
rect 1455 1755 1459 1759
rect 1511 1759 1515 1763
rect 1519 1755 1523 1759
rect 1575 1759 1579 1763
rect 1583 1755 1587 1759
rect 1595 1759 1599 1763
rect 1647 1755 1651 1759
rect 1695 1759 1699 1763
rect 1703 1755 1707 1759
rect 1751 1759 1755 1763
rect 1759 1755 1763 1759
rect 1799 1759 1803 1763
rect 1807 1755 1811 1759
rect 1095 1747 1099 1751
rect 1675 1747 1679 1751
rect 1863 1755 1867 1759
rect 1903 1759 1907 1763
rect 1919 1755 1923 1759
rect 1967 1759 1971 1763
rect 1975 1755 1979 1759
rect 1831 1747 1835 1751
rect 111 1732 115 1736
rect 459 1727 463 1731
rect 499 1727 503 1731
rect 539 1727 543 1731
rect 579 1727 583 1731
rect 619 1727 623 1731
rect 659 1727 663 1731
rect 675 1727 676 1731
rect 676 1727 679 1731
rect 703 1727 707 1731
rect 743 1727 747 1731
rect 799 1727 803 1731
rect 863 1727 867 1731
rect 927 1727 931 1731
rect 1203 1735 1207 1739
rect 1239 1732 1243 1736
rect 1095 1727 1096 1731
rect 1096 1727 1099 1731
rect 1127 1727 1131 1731
rect 1279 1732 1283 1736
rect 1315 1723 1319 1727
rect 1355 1727 1359 1731
rect 1367 1727 1368 1731
rect 1368 1727 1371 1731
rect 1603 1735 1607 1739
rect 1799 1735 1803 1739
rect 1447 1727 1451 1731
rect 1511 1727 1515 1731
rect 1575 1727 1579 1731
rect 1675 1727 1676 1731
rect 1676 1727 1679 1731
rect 1695 1727 1699 1731
rect 1751 1727 1755 1731
rect 1831 1727 1832 1731
rect 1832 1727 1835 1731
rect 2407 1732 2411 1736
rect 1967 1727 1971 1731
rect 111 1715 115 1719
rect 1239 1715 1243 1719
rect 1279 1715 1283 1719
rect 2407 1715 2411 1719
rect 407 1708 411 1712
rect 447 1708 451 1712
rect 487 1708 491 1712
rect 527 1708 531 1712
rect 567 1708 571 1712
rect 607 1708 611 1712
rect 647 1708 651 1712
rect 695 1708 699 1712
rect 751 1708 755 1712
rect 807 1708 811 1712
rect 871 1708 875 1712
rect 935 1708 939 1712
rect 999 1708 1003 1712
rect 1071 1708 1075 1712
rect 1143 1708 1147 1712
rect 1191 1708 1195 1712
rect 1303 1708 1307 1712
rect 1343 1708 1347 1712
rect 1391 1708 1395 1712
rect 1455 1708 1459 1712
rect 1519 1708 1523 1712
rect 1583 1708 1587 1712
rect 1647 1708 1651 1712
rect 1703 1708 1707 1712
rect 1759 1708 1763 1712
rect 1807 1708 1811 1712
rect 1863 1708 1867 1712
rect 1919 1708 1923 1712
rect 1975 1708 1979 1712
rect 279 1692 283 1696
rect 319 1692 323 1696
rect 359 1692 363 1696
rect 399 1692 403 1696
rect 447 1692 451 1696
rect 495 1692 499 1696
rect 543 1692 547 1696
rect 591 1692 595 1696
rect 639 1692 643 1696
rect 687 1692 691 1696
rect 735 1692 739 1696
rect 783 1692 787 1696
rect 839 1692 843 1696
rect 895 1692 899 1696
rect 1303 1692 1307 1696
rect 1343 1692 1347 1696
rect 1383 1692 1387 1696
rect 1423 1692 1427 1696
rect 1463 1692 1467 1696
rect 1503 1692 1507 1696
rect 1559 1692 1563 1696
rect 1623 1692 1627 1696
rect 1687 1692 1691 1696
rect 1751 1692 1755 1696
rect 1807 1692 1811 1696
rect 1863 1692 1867 1696
rect 1919 1692 1923 1696
rect 1975 1692 1979 1696
rect 2031 1692 2035 1696
rect 2087 1692 2091 1696
rect 111 1685 115 1689
rect 1239 1685 1243 1689
rect 1279 1685 1283 1689
rect 2407 1685 2411 1689
rect 567 1679 571 1683
rect 1595 1679 1599 1683
rect 2111 1679 2115 1683
rect 111 1668 115 1672
rect 331 1671 335 1675
rect 367 1671 371 1675
rect 435 1671 439 1675
rect 751 1671 755 1675
rect 799 1671 803 1675
rect 819 1671 823 1675
rect 423 1663 427 1667
rect 711 1663 715 1667
rect 1239 1668 1243 1672
rect 1279 1668 1283 1672
rect 919 1663 923 1667
rect 1351 1671 1355 1675
rect 1407 1663 1411 1667
rect 1431 1671 1435 1675
rect 1471 1671 1475 1675
rect 1787 1671 1791 1675
rect 1955 1671 1959 1675
rect 1487 1663 1491 1667
rect 2407 1668 2411 1672
rect 1943 1663 1947 1667
rect 279 1645 283 1649
rect 319 1645 323 1649
rect 359 1645 363 1649
rect 399 1645 403 1649
rect 447 1645 451 1649
rect 495 1645 499 1649
rect 543 1645 547 1649
rect 591 1645 595 1649
rect 639 1645 643 1649
rect 687 1645 691 1649
rect 735 1645 739 1649
rect 783 1645 787 1649
rect 839 1645 843 1649
rect 895 1645 899 1649
rect 1303 1645 1307 1649
rect 1343 1645 1347 1649
rect 1383 1645 1387 1649
rect 1423 1645 1427 1649
rect 1463 1645 1467 1649
rect 1503 1645 1507 1649
rect 1559 1645 1563 1649
rect 1623 1645 1627 1649
rect 1687 1645 1691 1649
rect 1751 1645 1755 1649
rect 1807 1645 1811 1649
rect 1863 1645 1867 1649
rect 1919 1645 1923 1649
rect 1975 1645 1979 1649
rect 2031 1645 2035 1649
rect 2087 1645 2091 1649
rect 331 1639 335 1643
rect 367 1639 371 1643
rect 407 1639 411 1643
rect 423 1639 424 1643
rect 424 1639 427 1643
rect 567 1639 568 1643
rect 568 1639 571 1643
rect 703 1639 707 1643
rect 711 1639 712 1643
rect 712 1639 715 1643
rect 751 1639 755 1643
rect 799 1639 803 1643
rect 919 1639 920 1643
rect 920 1639 923 1643
rect 1351 1639 1355 1643
rect 1367 1639 1368 1643
rect 1368 1639 1371 1643
rect 1407 1639 1408 1643
rect 1408 1639 1411 1643
rect 1471 1639 1475 1643
rect 1487 1639 1488 1643
rect 1488 1639 1491 1643
rect 1787 1639 1791 1643
rect 1943 1639 1944 1643
rect 1944 1639 1947 1643
rect 2111 1639 2112 1643
rect 2112 1639 2115 1643
rect 135 1611 139 1615
rect 163 1615 164 1619
rect 164 1615 167 1619
rect 175 1611 179 1615
rect 187 1615 191 1619
rect 215 1611 219 1615
rect 255 1611 259 1615
rect 267 1615 271 1619
rect 311 1611 315 1615
rect 327 1615 331 1619
rect 391 1611 395 1615
rect 463 1615 467 1619
rect 471 1611 475 1615
rect 551 1615 555 1619
rect 559 1611 563 1615
rect 571 1615 575 1619
rect 639 1611 643 1615
rect 711 1615 715 1619
rect 719 1611 723 1615
rect 783 1615 787 1619
rect 791 1611 795 1615
rect 819 1615 820 1619
rect 820 1615 823 1619
rect 855 1611 859 1615
rect 867 1615 871 1619
rect 919 1611 923 1615
rect 975 1615 979 1619
rect 983 1611 987 1615
rect 1039 1615 1043 1619
rect 1047 1611 1051 1615
rect 1059 1615 1063 1619
rect 1303 1611 1307 1615
rect 1359 1619 1363 1623
rect 1343 1611 1347 1615
rect 1399 1619 1403 1623
rect 1431 1619 1435 1623
rect 1383 1611 1387 1615
rect 1423 1611 1427 1615
rect 1439 1615 1443 1619
rect 1463 1611 1467 1615
rect 1475 1615 1479 1619
rect 1503 1611 1507 1615
rect 1515 1615 1519 1619
rect 1559 1611 1563 1615
rect 1623 1615 1627 1619
rect 1631 1611 1635 1615
rect 1695 1615 1699 1619
rect 1703 1611 1707 1615
rect 1775 1615 1779 1619
rect 1783 1611 1787 1615
rect 1795 1615 1799 1619
rect 1855 1611 1859 1615
rect 1919 1615 1923 1619
rect 1927 1611 1931 1615
rect 1955 1615 1956 1619
rect 1956 1615 1959 1619
rect 1999 1611 2003 1615
rect 2011 1615 2015 1619
rect 2063 1611 2067 1615
rect 2119 1615 2123 1619
rect 2127 1611 2131 1615
rect 2183 1615 2187 1619
rect 2191 1611 2195 1615
rect 2203 1615 2207 1619
rect 2255 1611 2259 1615
rect 2279 1615 2280 1619
rect 2280 1615 2283 1619
rect 2319 1611 2323 1615
rect 2331 1615 2335 1619
rect 2359 1611 2363 1615
rect 2371 1615 2375 1619
rect 111 1588 115 1592
rect 163 1591 167 1595
rect 267 1583 271 1587
rect 327 1583 331 1587
rect 571 1591 575 1595
rect 867 1591 871 1595
rect 407 1583 411 1587
rect 463 1583 467 1587
rect 551 1583 555 1587
rect 711 1583 715 1587
rect 783 1583 787 1587
rect 1059 1591 1063 1595
rect 1239 1588 1243 1592
rect 931 1583 935 1587
rect 975 1583 979 1587
rect 1039 1583 1043 1587
rect 1279 1588 1283 1592
rect 1439 1591 1443 1595
rect 1359 1583 1363 1587
rect 1399 1583 1403 1587
rect 1475 1583 1479 1587
rect 1515 1591 1519 1595
rect 2011 1591 2015 1595
rect 1511 1583 1515 1587
rect 1623 1583 1627 1587
rect 1695 1583 1699 1587
rect 1775 1583 1779 1587
rect 1919 1583 1923 1587
rect 2203 1591 2207 1595
rect 2407 1588 2411 1592
rect 2043 1583 2047 1587
rect 2119 1583 2123 1587
rect 2183 1583 2187 1587
rect 2331 1583 2335 1587
rect 2371 1583 2375 1587
rect 111 1571 115 1575
rect 1239 1571 1243 1575
rect 1279 1571 1283 1575
rect 2347 1575 2351 1579
rect 2407 1571 2411 1575
rect 135 1564 139 1568
rect 175 1564 179 1568
rect 215 1564 219 1568
rect 255 1564 259 1568
rect 311 1564 315 1568
rect 391 1564 395 1568
rect 471 1564 475 1568
rect 559 1564 563 1568
rect 639 1564 643 1568
rect 719 1564 723 1568
rect 791 1564 795 1568
rect 855 1564 859 1568
rect 919 1564 923 1568
rect 983 1564 987 1568
rect 1047 1564 1051 1568
rect 1303 1564 1307 1568
rect 1343 1564 1347 1568
rect 1383 1564 1387 1568
rect 1423 1564 1427 1568
rect 1463 1564 1467 1568
rect 1503 1564 1507 1568
rect 1559 1564 1563 1568
rect 1631 1564 1635 1568
rect 1703 1564 1707 1568
rect 1783 1564 1787 1568
rect 1855 1564 1859 1568
rect 1927 1564 1931 1568
rect 1999 1564 2003 1568
rect 2063 1564 2067 1568
rect 2127 1564 2131 1568
rect 2191 1564 2195 1568
rect 2255 1564 2259 1568
rect 2319 1564 2323 1568
rect 2359 1564 2363 1568
rect 151 1548 155 1552
rect 199 1548 203 1552
rect 263 1548 267 1552
rect 343 1548 347 1552
rect 439 1548 443 1552
rect 535 1548 539 1552
rect 639 1548 643 1552
rect 735 1548 739 1552
rect 823 1548 827 1552
rect 903 1548 907 1552
rect 975 1548 979 1552
rect 1047 1548 1051 1552
rect 1119 1548 1123 1552
rect 1191 1548 1195 1552
rect 1471 1552 1475 1556
rect 1623 1552 1627 1556
rect 1759 1552 1763 1556
rect 1871 1552 1875 1556
rect 1967 1552 1971 1556
rect 2055 1552 2059 1556
rect 2127 1552 2131 1556
rect 2191 1552 2195 1556
rect 2255 1552 2259 1556
rect 2319 1552 2323 1556
rect 2359 1552 2363 1556
rect 111 1541 115 1545
rect 1239 1541 1243 1545
rect 1279 1545 1283 1549
rect 2407 1545 2411 1549
rect 111 1524 115 1528
rect 187 1527 191 1531
rect 207 1527 211 1531
rect 1063 1527 1067 1531
rect 1135 1527 1139 1531
rect 1207 1527 1211 1531
rect 999 1519 1003 1523
rect 1179 1519 1183 1523
rect 1239 1524 1243 1528
rect 1279 1528 1283 1532
rect 1639 1531 1643 1535
rect 1795 1539 1799 1543
rect 2143 1531 2147 1535
rect 2207 1531 2211 1535
rect 2271 1531 2275 1535
rect 2279 1531 2280 1535
rect 2280 1531 2283 1535
rect 2375 1531 2379 1535
rect 2383 1531 2384 1535
rect 2384 1531 2387 1535
rect 2407 1528 2411 1532
rect 2079 1523 2083 1527
rect 151 1501 155 1505
rect 199 1501 203 1505
rect 263 1501 267 1505
rect 343 1501 347 1505
rect 439 1501 443 1505
rect 535 1501 539 1505
rect 639 1501 643 1505
rect 735 1501 739 1505
rect 823 1501 827 1505
rect 903 1501 907 1505
rect 975 1501 979 1505
rect 1047 1501 1051 1505
rect 1119 1501 1123 1505
rect 1191 1501 1195 1505
rect 1471 1505 1475 1509
rect 1623 1505 1627 1509
rect 1759 1505 1763 1509
rect 1871 1505 1875 1509
rect 1967 1505 1971 1509
rect 2055 1505 2059 1509
rect 2127 1505 2131 1509
rect 2191 1505 2195 1509
rect 2255 1505 2259 1509
rect 2319 1505 2323 1509
rect 2359 1505 2363 1509
rect 207 1495 211 1499
rect 579 1495 583 1499
rect 931 1495 932 1499
rect 932 1495 935 1499
rect 999 1495 1000 1499
rect 1000 1495 1003 1499
rect 1063 1495 1067 1499
rect 1135 1495 1139 1499
rect 1207 1495 1211 1499
rect 1511 1499 1515 1503
rect 1639 1499 1643 1503
rect 2043 1499 2047 1503
rect 2079 1499 2080 1503
rect 2080 1499 2083 1503
rect 2143 1499 2147 1503
rect 2207 1499 2211 1503
rect 2271 1499 2275 1503
rect 2347 1499 2348 1503
rect 2348 1499 2351 1503
rect 2375 1499 2379 1503
rect 319 1467 323 1471
rect 347 1471 348 1475
rect 348 1471 351 1475
rect 359 1467 363 1471
rect 415 1475 419 1479
rect 399 1467 403 1471
rect 439 1471 443 1475
rect 447 1467 451 1471
rect 495 1471 499 1475
rect 503 1467 507 1471
rect 551 1471 555 1475
rect 559 1467 563 1471
rect 607 1471 611 1475
rect 615 1467 619 1471
rect 631 1471 635 1475
rect 671 1467 675 1471
rect 727 1471 731 1475
rect 735 1467 739 1471
rect 791 1471 795 1475
rect 799 1467 803 1471
rect 847 1471 851 1475
rect 855 1467 859 1471
rect 903 1471 907 1475
rect 911 1467 915 1471
rect 959 1471 963 1475
rect 967 1467 971 1471
rect 1015 1471 1019 1475
rect 1023 1467 1027 1471
rect 1087 1467 1091 1471
rect 1151 1467 1155 1471
rect 1179 1471 1180 1475
rect 1180 1471 1183 1475
rect 1191 1467 1195 1471
rect 1203 1471 1207 1475
rect 1111 1459 1115 1463
rect 1219 1463 1223 1467
rect 1303 1455 1307 1459
rect 1375 1455 1379 1459
rect 1387 1459 1391 1463
rect 1479 1455 1483 1459
rect 1575 1459 1579 1463
rect 1583 1455 1587 1459
rect 1679 1459 1683 1463
rect 1687 1455 1691 1459
rect 1699 1459 1703 1463
rect 1783 1455 1787 1459
rect 1871 1455 1875 1459
rect 1943 1459 1947 1463
rect 1951 1455 1955 1459
rect 2023 1459 2027 1463
rect 2031 1455 2035 1459
rect 2095 1459 2099 1463
rect 2103 1455 2107 1459
rect 2159 1459 2163 1463
rect 2167 1455 2171 1459
rect 2231 1459 2235 1463
rect 2239 1455 2243 1459
rect 2303 1459 2307 1463
rect 2311 1455 2315 1459
rect 2323 1459 2327 1463
rect 2359 1455 2363 1459
rect 2383 1459 2384 1463
rect 2384 1459 2387 1463
rect 111 1444 115 1448
rect 347 1447 351 1451
rect 415 1439 419 1443
rect 439 1439 443 1443
rect 495 1439 499 1443
rect 551 1439 555 1443
rect 607 1439 611 1443
rect 111 1427 115 1431
rect 579 1431 583 1435
rect 727 1439 731 1443
rect 791 1439 795 1443
rect 847 1439 851 1443
rect 903 1439 907 1443
rect 959 1439 963 1443
rect 1203 1447 1207 1451
rect 1239 1444 1243 1448
rect 1111 1439 1112 1443
rect 1112 1439 1115 1443
rect 1219 1439 1220 1443
rect 1220 1439 1223 1443
rect 839 1431 843 1435
rect 1279 1432 1283 1436
rect 1239 1427 1243 1431
rect 1387 1427 1391 1431
rect 1699 1435 1703 1439
rect 1459 1427 1463 1431
rect 1575 1427 1579 1431
rect 1679 1427 1683 1431
rect 2407 1432 2411 1436
rect 319 1420 323 1424
rect 359 1420 363 1424
rect 399 1420 403 1424
rect 447 1420 451 1424
rect 503 1420 507 1424
rect 559 1420 563 1424
rect 615 1420 619 1424
rect 671 1420 675 1424
rect 735 1420 739 1424
rect 799 1420 803 1424
rect 855 1420 859 1424
rect 911 1420 915 1424
rect 967 1420 971 1424
rect 1023 1420 1027 1424
rect 1087 1420 1091 1424
rect 1151 1420 1155 1424
rect 1191 1420 1195 1424
rect 1943 1427 1947 1431
rect 2023 1427 2027 1431
rect 2095 1427 2099 1431
rect 2159 1427 2163 1431
rect 2231 1427 2235 1431
rect 2303 1427 2307 1431
rect 1279 1415 1283 1419
rect 2095 1419 2099 1423
rect 2407 1415 2411 1419
rect 263 1404 267 1408
rect 303 1404 307 1408
rect 343 1404 347 1408
rect 391 1404 395 1408
rect 447 1404 451 1408
rect 503 1404 507 1408
rect 559 1404 563 1408
rect 623 1404 627 1408
rect 687 1404 691 1408
rect 751 1404 755 1408
rect 815 1404 819 1408
rect 879 1404 883 1408
rect 951 1404 955 1408
rect 1023 1404 1027 1408
rect 1303 1408 1307 1412
rect 1375 1408 1379 1412
rect 1479 1408 1483 1412
rect 1583 1408 1587 1412
rect 1687 1408 1691 1412
rect 1783 1408 1787 1412
rect 1871 1408 1875 1412
rect 1951 1408 1955 1412
rect 2031 1408 2035 1412
rect 2103 1408 2107 1412
rect 2167 1408 2171 1412
rect 2239 1408 2243 1412
rect 2311 1408 2315 1412
rect 2359 1408 2363 1412
rect 111 1397 115 1401
rect 1239 1397 1243 1401
rect 1303 1396 1307 1400
rect 1343 1396 1347 1400
rect 1399 1396 1403 1400
rect 1471 1396 1475 1400
rect 1551 1396 1555 1400
rect 1639 1396 1643 1400
rect 1727 1396 1731 1400
rect 1815 1396 1819 1400
rect 1903 1396 1907 1400
rect 1991 1396 1995 1400
rect 2071 1396 2075 1400
rect 2151 1396 2155 1400
rect 2223 1396 2227 1400
rect 2303 1396 2307 1400
rect 2359 1396 2363 1400
rect 1015 1391 1019 1395
rect 1279 1389 1283 1393
rect 2407 1389 2411 1393
rect 111 1380 115 1384
rect 311 1383 315 1387
rect 407 1383 411 1387
rect 463 1383 467 1387
rect 519 1383 523 1387
rect 575 1383 579 1387
rect 631 1383 635 1387
rect 967 1383 971 1387
rect 1039 1383 1043 1387
rect 367 1375 371 1379
rect 1239 1380 1243 1384
rect 2323 1383 2327 1387
rect 783 1375 787 1379
rect 1279 1372 1283 1376
rect 1351 1375 1355 1379
rect 1495 1367 1499 1371
rect 1575 1375 1576 1379
rect 1576 1375 1579 1379
rect 1747 1367 1751 1371
rect 1927 1375 1928 1379
rect 1928 1375 1931 1379
rect 2375 1375 2379 1379
rect 2383 1375 2384 1379
rect 2384 1375 2387 1379
rect 2407 1372 2411 1376
rect 2191 1367 2195 1371
rect 263 1357 267 1361
rect 303 1357 307 1361
rect 343 1357 347 1361
rect 391 1357 395 1361
rect 447 1357 451 1361
rect 503 1357 507 1361
rect 559 1357 563 1361
rect 623 1357 627 1361
rect 687 1357 691 1361
rect 751 1357 755 1361
rect 815 1357 819 1361
rect 879 1357 883 1361
rect 951 1357 955 1361
rect 1023 1357 1027 1361
rect 311 1351 315 1355
rect 351 1351 355 1355
rect 367 1351 368 1355
rect 368 1351 371 1355
rect 407 1351 411 1355
rect 463 1351 467 1355
rect 519 1351 523 1355
rect 575 1351 579 1355
rect 839 1351 840 1355
rect 840 1351 843 1355
rect 867 1351 871 1355
rect 967 1351 971 1355
rect 1039 1351 1043 1355
rect 1303 1349 1307 1353
rect 1343 1349 1347 1353
rect 1399 1349 1403 1353
rect 1471 1349 1475 1353
rect 1551 1349 1555 1353
rect 1639 1349 1643 1353
rect 1727 1349 1731 1353
rect 1815 1349 1819 1353
rect 1903 1349 1907 1353
rect 1351 1343 1355 1347
rect 1459 1343 1463 1347
rect 1495 1343 1496 1347
rect 1496 1343 1499 1347
rect 1747 1343 1751 1347
rect 1927 1351 1931 1355
rect 1991 1349 1995 1353
rect 2071 1349 2075 1353
rect 2151 1349 2155 1353
rect 2223 1349 2227 1353
rect 2303 1349 2307 1353
rect 2359 1349 2363 1353
rect 2095 1343 2096 1347
rect 2096 1343 2099 1347
rect 2295 1343 2299 1347
rect 2375 1343 2379 1347
rect 135 1323 139 1327
rect 191 1331 195 1335
rect 175 1323 179 1327
rect 203 1327 204 1331
rect 204 1327 207 1331
rect 215 1323 219 1327
rect 239 1327 240 1331
rect 240 1327 243 1331
rect 255 1323 259 1327
rect 163 1315 167 1319
rect 327 1323 331 1327
rect 399 1327 403 1331
rect 407 1323 411 1327
rect 487 1327 491 1331
rect 495 1323 499 1327
rect 507 1327 511 1331
rect 583 1323 587 1327
rect 663 1327 667 1331
rect 671 1323 675 1327
rect 751 1327 755 1331
rect 759 1323 763 1327
rect 783 1327 784 1331
rect 784 1327 787 1331
rect 839 1323 843 1327
rect 911 1327 915 1331
rect 919 1323 923 1327
rect 999 1327 1003 1331
rect 1007 1323 1011 1327
rect 1087 1327 1091 1331
rect 1095 1323 1099 1327
rect 1107 1327 1111 1331
rect 1447 1315 1451 1319
rect 1503 1323 1507 1327
rect 1487 1315 1491 1319
rect 1543 1323 1547 1327
rect 1575 1323 1579 1327
rect 1527 1315 1531 1319
rect 1567 1315 1571 1319
rect 1583 1319 1587 1323
rect 1615 1315 1619 1319
rect 1663 1319 1667 1323
rect 1671 1315 1675 1319
rect 1711 1319 1715 1323
rect 1719 1315 1723 1319
rect 1731 1319 1735 1323
rect 1775 1315 1779 1319
rect 1823 1319 1827 1323
rect 1831 1315 1835 1319
rect 1895 1319 1899 1323
rect 1903 1315 1907 1319
rect 1963 1319 1967 1323
rect 1983 1315 1987 1319
rect 2063 1319 2067 1323
rect 2071 1315 2075 1319
rect 2159 1319 2163 1323
rect 2167 1315 2171 1319
rect 2191 1319 2192 1323
rect 2192 1319 2195 1323
rect 2271 1315 2275 1319
rect 2283 1319 2287 1323
rect 2359 1315 2363 1319
rect 2383 1319 2384 1323
rect 2384 1319 2387 1323
rect 111 1300 115 1304
rect 203 1303 207 1307
rect 163 1295 164 1299
rect 164 1295 167 1299
rect 191 1295 195 1299
rect 507 1303 511 1307
rect 1239 1300 1243 1304
rect 351 1295 352 1299
rect 352 1295 355 1299
rect 399 1295 403 1299
rect 487 1295 491 1299
rect 543 1295 547 1299
rect 663 1295 667 1299
rect 751 1295 755 1299
rect 867 1295 868 1299
rect 868 1295 871 1299
rect 911 1295 915 1299
rect 999 1295 1003 1299
rect 1087 1295 1091 1299
rect 1279 1292 1283 1296
rect 111 1283 115 1287
rect 1239 1283 1243 1287
rect 1583 1295 1587 1299
rect 1503 1287 1507 1291
rect 1543 1287 1547 1291
rect 1731 1295 1735 1299
rect 2407 1292 2411 1296
rect 1623 1287 1627 1291
rect 1663 1287 1667 1291
rect 1711 1287 1715 1291
rect 1823 1287 1827 1291
rect 1895 1287 1899 1291
rect 1963 1287 1967 1291
rect 2063 1287 2067 1291
rect 2159 1287 2163 1291
rect 2295 1287 2296 1291
rect 2296 1287 2299 1291
rect 2383 1287 2384 1291
rect 2384 1287 2387 1291
rect 135 1276 139 1280
rect 175 1276 179 1280
rect 215 1276 219 1280
rect 255 1276 259 1280
rect 327 1276 331 1280
rect 407 1276 411 1280
rect 495 1276 499 1280
rect 583 1276 587 1280
rect 671 1276 675 1280
rect 759 1276 763 1280
rect 839 1276 843 1280
rect 919 1276 923 1280
rect 1007 1276 1011 1280
rect 1095 1276 1099 1280
rect 1279 1275 1283 1279
rect 2143 1279 2147 1283
rect 2407 1275 2411 1279
rect 1447 1268 1451 1272
rect 1487 1268 1491 1272
rect 1527 1268 1531 1272
rect 1567 1268 1571 1272
rect 1615 1268 1619 1272
rect 1671 1268 1675 1272
rect 1719 1268 1723 1272
rect 1775 1268 1779 1272
rect 1831 1268 1835 1272
rect 1903 1268 1907 1272
rect 1983 1268 1987 1272
rect 2071 1268 2075 1272
rect 2167 1268 2171 1272
rect 2271 1268 2275 1272
rect 2359 1268 2363 1272
rect 135 1260 139 1264
rect 175 1260 179 1264
rect 247 1260 251 1264
rect 327 1260 331 1264
rect 415 1260 419 1264
rect 503 1260 507 1264
rect 591 1260 595 1264
rect 671 1260 675 1264
rect 743 1260 747 1264
rect 815 1260 819 1264
rect 879 1260 883 1264
rect 943 1260 947 1264
rect 1007 1260 1011 1264
rect 1071 1260 1075 1264
rect 111 1253 115 1257
rect 1239 1253 1243 1257
rect 1511 1252 1515 1256
rect 1551 1252 1555 1256
rect 1591 1252 1595 1256
rect 1631 1252 1635 1256
rect 1671 1252 1675 1256
rect 1711 1252 1715 1256
rect 1751 1252 1755 1256
rect 1791 1252 1795 1256
rect 1839 1252 1843 1256
rect 1903 1252 1907 1256
rect 1967 1252 1971 1256
rect 2039 1252 2043 1256
rect 2119 1252 2123 1256
rect 2207 1252 2211 1256
rect 2295 1252 2299 1256
rect 2359 1252 2363 1256
rect 1279 1245 1283 1249
rect 2407 1245 2411 1249
rect 111 1236 115 1240
rect 191 1239 195 1243
rect 239 1239 243 1243
rect 607 1239 611 1243
rect 663 1239 667 1243
rect 679 1239 683 1243
rect 959 1239 963 1243
rect 1023 1239 1027 1243
rect 1087 1239 1091 1243
rect 1107 1239 1111 1243
rect 423 1231 427 1235
rect 1239 1236 1243 1240
rect 903 1231 907 1235
rect 1279 1228 1283 1232
rect 1559 1231 1563 1235
rect 1599 1231 1603 1235
rect 1687 1231 1691 1235
rect 1727 1231 1731 1235
rect 1759 1231 1763 1235
rect 1767 1231 1771 1235
rect 1807 1231 1811 1235
rect 2031 1231 2035 1235
rect 2283 1231 2287 1235
rect 2319 1231 2320 1235
rect 2320 1231 2323 1235
rect 2407 1228 2411 1232
rect 1655 1223 1659 1227
rect 135 1213 139 1217
rect 175 1213 179 1217
rect 247 1213 251 1217
rect 327 1213 331 1217
rect 415 1213 419 1217
rect 503 1213 507 1217
rect 591 1213 595 1217
rect 671 1213 675 1217
rect 743 1213 747 1217
rect 815 1213 819 1217
rect 879 1213 883 1217
rect 943 1213 947 1217
rect 1007 1213 1011 1217
rect 1071 1213 1075 1217
rect 159 1207 160 1211
rect 160 1207 163 1211
rect 191 1207 195 1211
rect 423 1207 427 1211
rect 543 1207 547 1211
rect 607 1207 611 1211
rect 663 1207 667 1211
rect 895 1207 899 1211
rect 903 1207 904 1211
rect 904 1207 907 1211
rect 959 1207 963 1211
rect 1023 1207 1027 1211
rect 1087 1207 1091 1211
rect 1511 1205 1515 1209
rect 1551 1205 1555 1209
rect 1591 1205 1595 1209
rect 1631 1205 1635 1209
rect 1671 1205 1675 1209
rect 1711 1205 1715 1209
rect 1751 1205 1755 1209
rect 1791 1205 1795 1209
rect 1839 1205 1843 1209
rect 1903 1205 1907 1209
rect 1967 1205 1971 1209
rect 2039 1205 2043 1209
rect 2119 1205 2123 1209
rect 2207 1205 2211 1209
rect 2295 1205 2299 1209
rect 2359 1205 2363 1209
rect 1559 1199 1563 1203
rect 1599 1199 1603 1203
rect 1616 1199 1620 1203
rect 1655 1199 1656 1203
rect 1656 1199 1659 1203
rect 1687 1199 1691 1203
rect 1727 1199 1731 1203
rect 1759 1199 1763 1203
rect 2031 1199 2035 1203
rect 2143 1199 2144 1203
rect 2144 1199 2147 1203
rect 2219 1199 2223 1203
rect 2383 1199 2384 1203
rect 2384 1199 2387 1203
rect 135 1175 139 1179
rect 191 1183 195 1187
rect 175 1175 179 1179
rect 223 1179 227 1183
rect 231 1175 235 1179
rect 295 1179 299 1183
rect 303 1175 307 1179
rect 375 1179 379 1183
rect 383 1175 387 1179
rect 399 1179 403 1183
rect 471 1175 475 1179
rect 551 1179 555 1183
rect 559 1175 563 1179
rect 631 1179 635 1183
rect 639 1175 643 1179
rect 679 1179 683 1183
rect 719 1175 723 1179
rect 739 1179 743 1183
rect 799 1175 803 1179
rect 811 1179 815 1183
rect 871 1175 875 1179
rect 883 1179 887 1183
rect 935 1175 939 1179
rect 983 1179 987 1183
rect 991 1175 995 1179
rect 1039 1179 1043 1183
rect 1047 1175 1051 1179
rect 1095 1179 1099 1183
rect 1103 1175 1107 1179
rect 1143 1179 1147 1183
rect 1151 1175 1155 1179
rect 1207 1183 1211 1187
rect 1191 1175 1195 1179
rect 1215 1179 1216 1183
rect 1216 1179 1219 1183
rect 1559 1171 1563 1175
rect 1615 1179 1619 1183
rect 1599 1171 1603 1175
rect 1627 1175 1628 1179
rect 1628 1175 1631 1179
rect 1639 1171 1643 1175
rect 1695 1179 1699 1183
rect 1679 1171 1683 1175
rect 1735 1179 1739 1183
rect 1719 1171 1723 1175
rect 1767 1179 1771 1183
rect 1759 1171 1763 1175
rect 1807 1179 1811 1183
rect 1799 1171 1803 1175
rect 1815 1175 1819 1179
rect 1855 1171 1859 1175
rect 1867 1175 1871 1179
rect 1927 1171 1931 1175
rect 1939 1175 1943 1179
rect 2023 1171 2027 1175
rect 2127 1175 2131 1179
rect 2135 1171 2139 1175
rect 2247 1175 2251 1179
rect 2255 1171 2259 1175
rect 2267 1175 2271 1179
rect 2319 1179 2323 1183
rect 2359 1171 2363 1175
rect 111 1152 115 1156
rect 1239 1152 1243 1156
rect 159 1147 160 1151
rect 160 1147 163 1151
rect 191 1147 195 1151
rect 223 1147 227 1151
rect 295 1147 299 1151
rect 375 1147 379 1151
rect 499 1147 500 1151
rect 500 1147 503 1151
rect 551 1147 555 1151
rect 631 1147 635 1151
rect 811 1147 815 1151
rect 883 1147 887 1151
rect 895 1147 896 1151
rect 896 1147 899 1151
rect 983 1147 987 1151
rect 1039 1147 1043 1151
rect 1095 1147 1099 1151
rect 1143 1147 1147 1151
rect 1207 1147 1211 1151
rect 1279 1148 1283 1152
rect 1627 1151 1631 1155
rect 111 1135 115 1139
rect 1015 1139 1019 1143
rect 1615 1143 1619 1147
rect 1695 1143 1699 1147
rect 1735 1143 1739 1147
rect 1815 1143 1819 1147
rect 1867 1143 1871 1147
rect 1939 1143 1943 1147
rect 2267 1151 2271 1155
rect 2407 1148 2411 1152
rect 1975 1143 1979 1147
rect 2127 1143 2131 1147
rect 2247 1143 2251 1147
rect 2383 1143 2384 1147
rect 2384 1143 2387 1147
rect 1239 1135 1243 1139
rect 135 1128 139 1132
rect 175 1128 179 1132
rect 231 1128 235 1132
rect 303 1128 307 1132
rect 383 1128 387 1132
rect 471 1128 475 1132
rect 559 1128 563 1132
rect 639 1128 643 1132
rect 719 1128 723 1132
rect 799 1128 803 1132
rect 871 1128 875 1132
rect 935 1128 939 1132
rect 991 1128 995 1132
rect 1047 1128 1051 1132
rect 1103 1128 1107 1132
rect 1151 1128 1155 1132
rect 1191 1128 1195 1132
rect 1279 1131 1283 1135
rect 1751 1135 1755 1139
rect 2407 1131 2411 1135
rect 1559 1124 1563 1128
rect 1599 1124 1603 1128
rect 1639 1124 1643 1128
rect 1679 1124 1683 1128
rect 1719 1124 1723 1128
rect 1759 1124 1763 1128
rect 1799 1124 1803 1128
rect 1855 1124 1859 1128
rect 1927 1124 1931 1128
rect 2023 1124 2027 1128
rect 2135 1124 2139 1128
rect 2255 1124 2259 1128
rect 2359 1124 2363 1128
rect 135 1116 139 1120
rect 215 1116 219 1120
rect 303 1116 307 1120
rect 391 1116 395 1120
rect 479 1116 483 1120
rect 559 1116 563 1120
rect 639 1116 643 1120
rect 711 1116 715 1120
rect 775 1116 779 1120
rect 839 1116 843 1120
rect 903 1116 907 1120
rect 959 1116 963 1120
rect 1023 1116 1027 1120
rect 1087 1116 1091 1120
rect 1151 1116 1155 1120
rect 1191 1116 1195 1120
rect 111 1109 115 1113
rect 1239 1109 1243 1113
rect 399 1103 403 1107
rect 1215 1103 1219 1107
rect 1535 1104 1539 1108
rect 1599 1104 1603 1108
rect 1663 1104 1667 1108
rect 1727 1104 1731 1108
rect 1791 1104 1795 1108
rect 1855 1104 1859 1108
rect 1911 1104 1915 1108
rect 1967 1104 1971 1108
rect 2023 1104 2027 1108
rect 2079 1104 2083 1108
rect 2135 1104 2139 1108
rect 2191 1104 2195 1108
rect 2255 1104 2259 1108
rect 2319 1104 2323 1108
rect 2359 1104 2363 1108
rect 111 1092 115 1096
rect 567 1095 571 1099
rect 575 1095 579 1099
rect 727 1095 731 1099
rect 739 1095 740 1099
rect 740 1095 743 1099
rect 1199 1095 1203 1099
rect 1279 1097 1283 1101
rect 2407 1097 2411 1101
rect 1239 1092 1243 1096
rect 983 1087 987 1091
rect 1279 1080 1283 1084
rect 1759 1075 1763 1079
rect 1991 1075 1995 1079
rect 2039 1083 2043 1087
rect 2219 1083 2220 1087
rect 2220 1083 2223 1087
rect 2227 1083 2231 1087
rect 2367 1083 2371 1087
rect 2407 1080 2411 1084
rect 2147 1075 2151 1079
rect 135 1069 139 1073
rect 215 1069 219 1073
rect 303 1069 307 1073
rect 391 1069 395 1073
rect 479 1069 483 1073
rect 559 1069 563 1073
rect 639 1069 643 1073
rect 711 1069 715 1073
rect 775 1069 779 1073
rect 839 1069 843 1073
rect 903 1069 907 1073
rect 959 1069 963 1073
rect 1023 1069 1027 1073
rect 1087 1069 1091 1073
rect 1151 1069 1155 1073
rect 1191 1069 1195 1073
rect 267 1055 271 1059
rect 499 1063 503 1067
rect 567 1063 571 1067
rect 611 1063 615 1067
rect 727 1063 731 1067
rect 1015 1063 1019 1067
rect 1199 1063 1203 1067
rect 1215 1063 1216 1067
rect 1216 1063 1219 1067
rect 1535 1057 1539 1061
rect 1599 1057 1603 1061
rect 1663 1057 1667 1061
rect 1727 1057 1731 1061
rect 1791 1057 1795 1061
rect 1855 1057 1859 1061
rect 1911 1057 1915 1061
rect 1967 1057 1971 1061
rect 2023 1057 2027 1061
rect 2079 1057 2083 1061
rect 2135 1057 2139 1061
rect 2191 1057 2195 1061
rect 2255 1057 2259 1061
rect 2319 1057 2323 1061
rect 2359 1057 2363 1061
rect 1751 1051 1752 1055
rect 1752 1051 1755 1055
rect 1975 1051 1979 1055
rect 1991 1051 1992 1055
rect 1992 1051 1995 1055
rect 2147 1051 2151 1055
rect 2227 1051 2231 1055
rect 2367 1051 2371 1055
rect 2383 1051 2384 1055
rect 2384 1051 2387 1055
rect 199 1035 203 1039
rect 227 1039 228 1043
rect 228 1039 231 1043
rect 239 1035 243 1039
rect 279 1039 283 1043
rect 287 1035 291 1039
rect 335 1039 339 1043
rect 343 1035 347 1039
rect 383 1039 387 1043
rect 391 1035 395 1039
rect 407 1039 411 1043
rect 439 1035 443 1039
rect 479 1039 483 1043
rect 487 1035 491 1039
rect 527 1039 531 1043
rect 575 1043 579 1047
rect 535 1035 539 1039
rect 583 1035 587 1039
rect 623 1039 627 1043
rect 631 1035 635 1039
rect 679 1035 683 1039
rect 719 1039 723 1043
rect 727 1035 731 1039
rect 775 1039 779 1043
rect 783 1035 787 1039
rect 831 1039 835 1043
rect 839 1035 843 1039
rect 887 1039 891 1043
rect 895 1035 899 1039
rect 951 1039 955 1043
rect 959 1035 963 1039
rect 983 1039 984 1043
rect 984 1039 987 1043
rect 1023 1035 1027 1039
rect 1079 1039 1083 1043
rect 1087 1035 1091 1039
rect 1111 1039 1112 1043
rect 1112 1039 1115 1043
rect 1151 1035 1155 1039
rect 1167 1039 1171 1043
rect 1191 1035 1195 1039
rect 1203 1039 1207 1043
rect 111 1012 115 1016
rect 267 1015 271 1019
rect 1167 1015 1171 1019
rect 1239 1012 1243 1016
rect 1503 1015 1507 1019
rect 1615 1019 1619 1023
rect 1623 1015 1627 1019
rect 1727 1019 1731 1023
rect 1735 1015 1739 1019
rect 1759 1019 1760 1023
rect 1760 1019 1763 1023
rect 1831 1015 1835 1019
rect 1935 1023 1939 1027
rect 1919 1015 1923 1019
rect 2039 1023 2043 1027
rect 1999 1015 2003 1019
rect 2071 1015 2075 1019
rect 2083 1019 2087 1023
rect 2143 1015 2147 1019
rect 2199 1019 2203 1023
rect 2207 1015 2211 1019
rect 2271 1019 2275 1023
rect 2279 1015 2283 1019
rect 2291 1019 2295 1023
rect 235 1007 239 1011
rect 279 1007 283 1011
rect 335 1007 339 1011
rect 383 1007 387 1011
rect 479 1007 483 1011
rect 527 1007 531 1011
rect 611 1007 612 1011
rect 612 1007 615 1011
rect 623 1007 627 1011
rect 719 1007 723 1011
rect 775 1007 779 1011
rect 831 1007 835 1011
rect 887 1007 891 1011
rect 951 1007 955 1011
rect 1079 1007 1083 1011
rect 1203 1007 1207 1011
rect 1215 1007 1216 1011
rect 1216 1007 1219 1011
rect 111 995 115 999
rect 575 999 579 1003
rect 1239 995 1243 999
rect 199 988 203 992
rect 239 988 243 992
rect 287 988 291 992
rect 343 988 347 992
rect 391 988 395 992
rect 439 988 443 992
rect 487 988 491 992
rect 535 988 539 992
rect 583 988 587 992
rect 631 988 635 992
rect 679 988 683 992
rect 727 988 731 992
rect 783 988 787 992
rect 839 988 843 992
rect 895 988 899 992
rect 959 988 963 992
rect 1023 988 1027 992
rect 1087 988 1091 992
rect 1151 988 1155 992
rect 1191 988 1195 992
rect 1279 992 1283 996
rect 1615 987 1619 991
rect 1727 987 1731 991
rect 2083 995 2087 999
rect 1935 987 1939 991
rect 2291 995 2295 999
rect 2407 992 2411 996
rect 2131 987 2135 991
rect 2199 987 2203 991
rect 2271 987 2275 991
rect 1279 975 1283 979
rect 2407 975 2411 979
rect 295 964 299 968
rect 343 964 347 968
rect 399 964 403 968
rect 471 964 475 968
rect 551 964 555 968
rect 639 964 643 968
rect 727 964 731 968
rect 807 964 811 968
rect 887 964 891 968
rect 959 964 963 968
rect 1023 964 1027 968
rect 1087 964 1091 968
rect 1151 964 1155 968
rect 1191 964 1195 968
rect 1503 968 1507 972
rect 1623 968 1627 972
rect 1735 968 1739 972
rect 1831 968 1835 972
rect 1919 968 1923 972
rect 1999 968 2003 972
rect 2071 968 2075 972
rect 2143 968 2147 972
rect 2207 968 2211 972
rect 2279 968 2283 972
rect 111 957 115 961
rect 1239 957 1243 961
rect 407 951 411 955
rect 1319 948 1323 952
rect 111 940 115 944
rect 655 943 659 947
rect 719 943 723 947
rect 739 943 743 947
rect 1111 943 1112 947
rect 1112 943 1115 947
rect 1199 943 1203 947
rect 1359 948 1363 952
rect 1399 948 1403 952
rect 1463 948 1467 952
rect 1543 948 1547 952
rect 1639 948 1643 952
rect 1735 948 1739 952
rect 1839 948 1843 952
rect 1935 948 1939 952
rect 2023 948 2027 952
rect 2103 948 2107 952
rect 2175 948 2179 952
rect 2239 948 2243 952
rect 2311 948 2315 952
rect 2359 948 2363 952
rect 1239 940 1243 944
rect 1279 941 1283 945
rect 2407 941 2411 945
rect 1215 935 1219 939
rect 1279 924 1283 928
rect 1347 927 1348 931
rect 1348 927 1351 931
rect 1367 927 1371 931
rect 1407 927 1411 931
rect 1491 927 1492 931
rect 1492 927 1495 931
rect 295 917 299 921
rect 343 917 347 921
rect 399 917 403 921
rect 471 917 475 921
rect 551 917 555 921
rect 639 917 643 921
rect 727 917 731 921
rect 807 917 811 921
rect 887 917 891 921
rect 959 917 963 921
rect 1023 917 1027 921
rect 1087 917 1091 921
rect 1151 917 1155 921
rect 1191 917 1195 921
rect 1427 919 1431 923
rect 1987 927 1991 931
rect 2255 927 2259 931
rect 2327 927 2331 931
rect 2375 927 2379 931
rect 2383 927 2384 931
rect 2384 927 2387 931
rect 2407 924 2411 928
rect 2199 919 2203 923
rect 559 911 563 915
rect 575 911 576 915
rect 576 911 579 915
rect 655 911 659 915
rect 719 911 723 915
rect 1079 911 1083 915
rect 1199 911 1203 915
rect 1215 911 1216 915
rect 1216 911 1219 915
rect 1319 901 1323 905
rect 1359 901 1363 905
rect 1399 901 1403 905
rect 1463 901 1467 905
rect 1543 901 1547 905
rect 1639 901 1643 905
rect 1735 901 1739 905
rect 1839 901 1843 905
rect 1935 901 1939 905
rect 2023 901 2027 905
rect 2103 901 2107 905
rect 2175 901 2179 905
rect 2239 901 2243 905
rect 2311 901 2315 905
rect 2359 901 2363 905
rect 1367 895 1371 899
rect 1407 895 1411 899
rect 1427 895 1428 899
rect 1428 895 1431 899
rect 1779 895 1783 899
rect 1987 895 1991 899
rect 2131 895 2132 899
rect 2132 895 2135 899
rect 2199 895 2200 899
rect 2200 895 2203 899
rect 2255 895 2259 899
rect 2327 895 2331 899
rect 2375 895 2379 899
rect 255 879 259 883
rect 311 879 315 883
rect 335 883 336 887
rect 336 883 339 887
rect 375 879 379 883
rect 387 883 391 887
rect 455 879 459 883
rect 467 883 471 887
rect 535 879 539 883
rect 547 883 551 887
rect 623 879 627 883
rect 703 883 707 887
rect 711 879 715 883
rect 739 883 740 887
rect 740 883 743 887
rect 791 879 795 883
rect 855 883 859 887
rect 863 879 867 883
rect 919 883 923 887
rect 935 879 939 883
rect 947 883 951 887
rect 999 879 1003 883
rect 1011 883 1015 887
rect 1055 879 1059 883
rect 1111 883 1115 887
rect 1119 879 1123 883
rect 1175 883 1179 887
rect 1183 879 1187 883
rect 1195 883 1199 887
rect 1347 875 1351 879
rect 111 856 115 860
rect 387 859 391 863
rect 467 851 471 855
rect 547 851 551 855
rect 559 851 560 855
rect 560 851 563 855
rect 639 851 643 855
rect 703 851 707 855
rect 947 859 951 863
rect 855 851 859 855
rect 1011 851 1015 855
rect 1195 859 1199 863
rect 1335 863 1339 867
rect 1363 867 1364 871
rect 1364 867 1367 871
rect 1375 863 1379 867
rect 1403 867 1404 871
rect 1404 867 1407 871
rect 1415 863 1419 867
rect 1471 863 1475 867
rect 1491 867 1495 871
rect 1535 863 1539 867
rect 1547 867 1551 871
rect 1607 863 1611 867
rect 1647 867 1651 871
rect 1679 863 1683 867
rect 1691 867 1695 871
rect 1751 863 1755 867
rect 1763 867 1767 871
rect 1823 863 1827 867
rect 1887 867 1891 871
rect 1895 863 1899 867
rect 1951 867 1955 871
rect 1959 863 1963 867
rect 2015 867 2019 871
rect 2023 863 2027 867
rect 2079 867 2083 871
rect 2087 863 2091 867
rect 2135 867 2139 871
rect 2143 863 2147 867
rect 2199 863 2203 867
rect 2247 867 2251 871
rect 2255 863 2259 867
rect 2311 867 2315 871
rect 2319 863 2323 867
rect 2347 867 2348 871
rect 2348 867 2351 871
rect 2359 863 2363 867
rect 2383 867 2384 871
rect 2384 867 2387 871
rect 1239 856 1243 860
rect 1079 851 1080 855
rect 1080 851 1083 855
rect 1111 851 1115 855
rect 1175 851 1179 855
rect 111 839 115 843
rect 1239 839 1243 843
rect 1279 840 1283 844
rect 1887 843 1891 847
rect 2347 843 2351 847
rect 255 832 259 836
rect 311 832 315 836
rect 375 832 379 836
rect 455 832 459 836
rect 535 832 539 836
rect 623 832 627 836
rect 711 832 715 836
rect 791 832 795 836
rect 863 832 867 836
rect 935 832 939 836
rect 999 832 1003 836
rect 1055 832 1059 836
rect 1119 832 1123 836
rect 1183 832 1187 836
rect 1351 835 1355 839
rect 1371 835 1375 839
rect 1411 835 1415 839
rect 1547 835 1551 839
rect 1575 835 1579 839
rect 1691 835 1695 839
rect 1763 835 1767 839
rect 1779 835 1780 839
rect 1780 835 1783 839
rect 2407 840 2411 844
rect 1951 835 1955 839
rect 2015 835 2019 839
rect 2079 835 2083 839
rect 2135 835 2139 839
rect 2247 835 2251 839
rect 2311 835 2315 839
rect 191 820 195 824
rect 247 820 251 824
rect 311 820 315 824
rect 383 820 387 824
rect 463 820 467 824
rect 543 820 547 824
rect 615 820 619 824
rect 687 820 691 824
rect 751 820 755 824
rect 815 820 819 824
rect 871 820 875 824
rect 927 820 931 824
rect 983 820 987 824
rect 1047 820 1051 824
rect 1279 823 1283 827
rect 2047 827 2051 831
rect 2383 827 2387 831
rect 2407 823 2411 827
rect 111 813 115 817
rect 1239 813 1243 817
rect 1335 816 1339 820
rect 1375 816 1379 820
rect 1415 816 1419 820
rect 1471 816 1475 820
rect 1535 816 1539 820
rect 1607 816 1611 820
rect 1679 816 1683 820
rect 1751 816 1755 820
rect 1823 816 1827 820
rect 1895 816 1899 820
rect 1959 816 1963 820
rect 2023 816 2027 820
rect 2087 816 2091 820
rect 2143 816 2147 820
rect 2199 816 2203 820
rect 2255 816 2259 820
rect 2319 816 2323 820
rect 2359 816 2363 820
rect 111 796 115 800
rect 271 799 272 803
rect 272 799 275 803
rect 335 799 336 803
rect 336 799 339 803
rect 347 799 351 803
rect 519 799 523 803
rect 527 799 531 803
rect 407 791 411 795
rect 895 791 899 795
rect 919 799 923 803
rect 1239 796 1243 800
rect 1303 800 1307 804
rect 1343 800 1347 804
rect 1407 800 1411 804
rect 1479 800 1483 804
rect 1551 800 1555 804
rect 1623 800 1627 804
rect 1695 800 1699 804
rect 1759 800 1763 804
rect 1823 800 1827 804
rect 1887 800 1891 804
rect 1951 800 1955 804
rect 2023 800 2027 804
rect 2103 800 2107 804
rect 2191 800 2195 804
rect 2279 800 2283 804
rect 2359 800 2363 804
rect 1071 791 1075 795
rect 1279 793 1283 797
rect 2407 793 2411 797
rect 191 773 195 777
rect 247 773 251 777
rect 311 773 315 777
rect 383 773 387 777
rect 463 773 467 777
rect 543 773 547 777
rect 615 773 619 777
rect 687 773 691 777
rect 751 773 755 777
rect 815 773 819 777
rect 871 773 875 777
rect 927 773 931 777
rect 983 773 987 777
rect 1047 773 1051 777
rect 1279 776 1283 780
rect 1359 779 1363 783
rect 1387 779 1391 783
rect 1395 779 1399 783
rect 1491 779 1495 783
rect 1647 779 1648 783
rect 1648 779 1651 783
rect 1799 779 1803 783
rect 2323 779 2327 783
rect 2407 776 2411 780
rect 263 767 267 771
rect 303 767 307 771
rect 347 767 351 771
rect 407 767 408 771
rect 408 767 411 771
rect 527 767 531 771
rect 639 767 640 771
rect 640 767 643 771
rect 887 767 891 771
rect 895 767 896 771
rect 896 767 899 771
rect 1071 767 1072 771
rect 1072 767 1075 771
rect 2303 771 2307 775
rect 1303 753 1307 757
rect 1343 753 1347 757
rect 1407 753 1411 757
rect 1479 753 1483 757
rect 1551 753 1555 757
rect 1623 753 1627 757
rect 1695 753 1699 757
rect 1759 753 1763 757
rect 1823 753 1827 757
rect 1887 753 1891 757
rect 1951 753 1955 757
rect 2023 753 2027 757
rect 2103 753 2107 757
rect 2191 753 2195 757
rect 2279 753 2283 757
rect 2359 753 2363 757
rect 135 743 139 747
rect 163 747 164 751
rect 164 747 167 751
rect 175 743 179 747
rect 199 747 200 751
rect 200 747 203 751
rect 215 743 219 747
rect 279 743 283 747
rect 343 747 347 751
rect 351 743 355 747
rect 363 747 367 751
rect 423 743 427 747
rect 487 747 491 751
rect 495 743 499 747
rect 519 747 520 751
rect 520 747 523 751
rect 559 743 563 747
rect 615 747 619 751
rect 623 743 627 747
rect 687 747 691 751
rect 695 743 699 747
rect 759 747 763 751
rect 783 743 787 747
rect 795 747 799 751
rect 879 743 883 747
rect 975 747 979 751
rect 983 743 987 747
rect 1087 747 1091 751
rect 1095 743 1099 747
rect 1107 747 1111 751
rect 1191 743 1195 747
rect 1319 747 1323 751
rect 1351 747 1355 751
rect 1359 747 1363 751
rect 1387 747 1391 751
rect 1575 747 1576 751
rect 1576 747 1579 751
rect 1719 747 1720 751
rect 1720 747 1723 751
rect 2047 747 2048 751
rect 2048 747 2051 751
rect 2143 747 2147 751
rect 2303 747 2304 751
rect 2304 747 2307 751
rect 2383 747 2384 751
rect 2384 747 2387 751
rect 111 720 115 724
rect 163 723 167 727
rect 363 723 367 727
rect 795 723 799 727
rect 303 715 304 719
rect 304 715 307 719
rect 343 715 347 719
rect 439 715 443 719
rect 487 715 491 719
rect 615 715 619 719
rect 687 715 691 719
rect 1107 723 1111 727
rect 1239 720 1243 724
rect 1303 723 1307 727
rect 1359 727 1363 731
rect 1367 723 1371 727
rect 1395 727 1396 731
rect 1396 727 1399 731
rect 1455 723 1459 727
rect 1491 727 1495 731
rect 1535 723 1539 727
rect 1547 727 1551 731
rect 1615 723 1619 727
rect 1663 727 1667 731
rect 1695 723 1699 727
rect 1707 727 1711 731
rect 1775 723 1779 727
rect 1799 727 1800 731
rect 1800 727 1803 731
rect 1855 723 1859 727
rect 1867 727 1871 731
rect 1943 723 1947 727
rect 1955 727 1959 731
rect 2031 723 2035 727
rect 2043 727 2047 731
rect 2119 723 2123 727
rect 2199 727 2203 731
rect 2207 723 2211 727
rect 2287 727 2291 731
rect 2295 723 2299 727
rect 2323 727 2324 731
rect 2324 727 2327 731
rect 2359 723 2363 727
rect 2371 727 2375 731
rect 887 715 891 719
rect 975 715 979 719
rect 1087 715 1091 719
rect 1175 715 1179 719
rect 111 703 115 707
rect 1239 703 1243 707
rect 135 696 139 700
rect 175 696 179 700
rect 215 696 219 700
rect 279 696 283 700
rect 351 696 355 700
rect 423 696 427 700
rect 495 696 499 700
rect 559 696 563 700
rect 623 696 627 700
rect 695 696 699 700
rect 783 696 787 700
rect 879 696 883 700
rect 983 696 987 700
rect 1095 696 1099 700
rect 1191 696 1195 700
rect 1279 700 1283 704
rect 2407 700 2411 704
rect 1319 695 1323 699
rect 1359 695 1363 699
rect 1547 695 1551 699
rect 1607 695 1611 699
rect 1707 695 1711 699
rect 1719 695 1720 699
rect 1720 695 1723 699
rect 1867 695 1871 699
rect 1955 695 1959 699
rect 2043 695 2047 699
rect 2135 695 2139 699
rect 2143 695 2144 699
rect 2144 695 2147 699
rect 2199 695 2203 699
rect 2371 695 2375 699
rect 2383 695 2384 699
rect 2384 695 2387 699
rect 1279 683 1283 687
rect 2407 683 2411 687
rect 135 676 139 680
rect 175 676 179 680
rect 231 676 235 680
rect 287 676 291 680
rect 343 676 347 680
rect 399 676 403 680
rect 455 676 459 680
rect 503 676 507 680
rect 559 676 563 680
rect 623 676 627 680
rect 695 676 699 680
rect 767 676 771 680
rect 839 676 843 680
rect 903 676 907 680
rect 967 676 971 680
rect 1023 676 1027 680
rect 1087 676 1091 680
rect 1151 676 1155 680
rect 1191 676 1195 680
rect 1303 676 1307 680
rect 1367 676 1371 680
rect 1455 676 1459 680
rect 1535 676 1539 680
rect 1615 676 1619 680
rect 1695 676 1699 680
rect 1775 676 1779 680
rect 1855 676 1859 680
rect 1943 676 1947 680
rect 2031 676 2035 680
rect 2119 676 2123 680
rect 2207 676 2211 680
rect 2295 676 2299 680
rect 2359 676 2363 680
rect 111 669 115 673
rect 1239 669 1243 673
rect 1591 664 1595 668
rect 1639 664 1643 668
rect 1687 664 1691 668
rect 1743 664 1747 668
rect 1799 664 1803 668
rect 1871 664 1875 668
rect 1951 664 1955 668
rect 2047 664 2051 668
rect 2151 664 2155 668
rect 2263 664 2267 668
rect 2359 664 2363 668
rect 111 652 115 656
rect 199 655 200 659
rect 200 655 203 659
rect 211 655 215 659
rect 495 655 499 659
rect 515 655 519 659
rect 311 647 315 651
rect 479 647 483 651
rect 639 655 643 659
rect 719 647 723 651
rect 759 655 763 659
rect 915 655 919 659
rect 1215 655 1216 659
rect 1216 655 1219 659
rect 1279 657 1283 661
rect 2407 657 2411 661
rect 863 647 867 651
rect 1239 652 1243 656
rect 1199 647 1203 651
rect 1279 640 1283 644
rect 1583 643 1587 647
rect 1663 643 1664 647
rect 1664 643 1667 647
rect 1975 643 1976 647
rect 1976 643 1979 647
rect 2083 643 2087 647
rect 2287 643 2288 647
rect 2288 643 2291 647
rect 2407 640 2411 644
rect 135 629 139 633
rect 175 629 179 633
rect 231 629 235 633
rect 287 629 291 633
rect 343 629 347 633
rect 399 629 403 633
rect 455 629 459 633
rect 503 629 507 633
rect 559 629 563 633
rect 623 629 627 633
rect 695 629 699 633
rect 767 629 771 633
rect 839 629 843 633
rect 903 629 907 633
rect 967 629 971 633
rect 1023 629 1027 633
rect 1087 629 1091 633
rect 1151 629 1155 633
rect 1191 629 1195 633
rect 159 623 160 627
rect 160 623 163 627
rect 211 623 215 627
rect 311 623 312 627
rect 312 623 315 627
rect 439 623 443 627
rect 479 623 480 627
rect 480 623 483 627
rect 495 623 499 627
rect 639 623 643 627
rect 663 623 667 627
rect 719 623 720 627
rect 720 623 723 627
rect 863 623 864 627
rect 864 623 867 627
rect 1103 623 1107 627
rect 1175 623 1176 627
rect 1176 623 1179 627
rect 1199 623 1203 627
rect 1591 617 1595 621
rect 1639 617 1643 621
rect 1687 617 1691 621
rect 1743 617 1747 621
rect 1799 617 1803 621
rect 1871 617 1875 621
rect 1951 617 1955 621
rect 2047 617 2051 621
rect 2151 617 2155 621
rect 2263 617 2267 621
rect 2359 617 2363 621
rect 1607 611 1611 615
rect 1891 611 1895 615
rect 2083 611 2087 615
rect 2135 611 2139 615
rect 2383 611 2384 615
rect 2384 611 2387 615
rect 135 599 139 603
rect 175 603 179 607
rect 183 599 187 603
rect 247 603 251 607
rect 255 599 259 603
rect 319 603 323 607
rect 327 599 331 603
rect 339 603 343 607
rect 399 599 403 603
rect 471 603 475 607
rect 479 599 483 603
rect 515 603 519 607
rect 559 599 563 603
rect 571 603 575 607
rect 639 599 643 603
rect 711 603 715 607
rect 719 599 723 603
rect 791 603 795 607
rect 799 599 803 603
rect 811 603 815 607
rect 879 599 883 603
rect 915 603 919 607
rect 951 599 955 603
rect 963 603 967 607
rect 1015 599 1019 603
rect 1027 603 1031 607
rect 1079 599 1083 603
rect 1135 603 1139 607
rect 1143 599 1147 603
rect 1183 603 1187 607
rect 1191 599 1195 603
rect 1215 603 1216 607
rect 1216 603 1219 607
rect 111 576 115 580
rect 159 571 160 575
rect 160 571 163 575
rect 175 571 179 575
rect 247 571 251 575
rect 319 571 323 575
rect 571 579 575 583
rect 1239 576 1243 580
rect 1559 579 1563 583
rect 1583 583 1584 587
rect 1584 583 1587 587
rect 1599 579 1603 583
rect 1611 583 1615 587
rect 1639 579 1643 583
rect 1651 583 1655 587
rect 1679 579 1683 583
rect 1707 583 1708 587
rect 1708 583 1711 587
rect 1719 579 1723 583
rect 1747 583 1748 587
rect 1748 583 1751 587
rect 1759 579 1763 583
rect 1799 583 1803 587
rect 1807 579 1811 583
rect 471 571 475 575
rect 579 571 583 575
rect 663 571 664 575
rect 664 571 667 575
rect 711 571 715 575
rect 791 571 795 575
rect 963 571 967 575
rect 1027 571 1031 575
rect 1095 571 1099 575
rect 1103 571 1104 575
rect 1104 571 1107 575
rect 1135 571 1139 575
rect 1183 571 1187 575
rect 1667 571 1671 575
rect 1855 579 1859 583
rect 1903 583 1907 587
rect 1911 579 1915 583
rect 1959 583 1963 587
rect 1975 587 1979 591
rect 1967 579 1971 583
rect 2031 579 2035 583
rect 2043 583 2047 587
rect 2095 579 2099 583
rect 2107 583 2111 587
rect 2167 579 2171 583
rect 2231 583 2235 587
rect 2239 579 2243 583
rect 2303 583 2307 587
rect 2311 579 2315 583
rect 2351 583 2355 587
rect 2359 579 2363 583
rect 111 559 115 563
rect 1239 559 1243 563
rect 135 552 139 556
rect 183 552 187 556
rect 255 552 259 556
rect 327 552 331 556
rect 399 552 403 556
rect 479 552 483 556
rect 559 552 563 556
rect 639 552 643 556
rect 719 552 723 556
rect 799 552 803 556
rect 879 552 883 556
rect 951 552 955 556
rect 1015 552 1019 556
rect 1079 552 1083 556
rect 1143 552 1147 556
rect 1191 552 1195 556
rect 1279 556 1283 560
rect 1747 559 1751 563
rect 2407 556 2411 560
rect 1611 551 1615 555
rect 1651 551 1655 555
rect 1667 551 1668 555
rect 1668 551 1671 555
rect 1735 551 1739 555
rect 1799 551 1803 555
rect 1891 551 1895 555
rect 1903 551 1907 555
rect 2043 551 2047 555
rect 2107 551 2111 555
rect 2123 551 2124 555
rect 2124 551 2127 555
rect 2231 551 2235 555
rect 2339 551 2340 555
rect 2340 551 2343 555
rect 2351 551 2355 555
rect 151 536 155 540
rect 223 536 227 540
rect 287 536 291 540
rect 351 536 355 540
rect 415 536 419 540
rect 479 536 483 540
rect 551 536 555 540
rect 623 536 627 540
rect 695 536 699 540
rect 767 536 771 540
rect 839 536 843 540
rect 919 536 923 540
rect 999 536 1003 540
rect 1079 536 1083 540
rect 1279 539 1283 543
rect 1707 543 1711 547
rect 2407 539 2411 543
rect 111 529 115 533
rect 1239 529 1243 533
rect 1559 532 1563 536
rect 1599 532 1603 536
rect 1639 532 1643 536
rect 1679 532 1683 536
rect 1719 532 1723 536
rect 1759 532 1763 536
rect 1807 532 1811 536
rect 1855 532 1859 536
rect 1911 532 1915 536
rect 1967 532 1971 536
rect 2031 532 2035 536
rect 2095 532 2099 536
rect 2167 532 2171 536
rect 2239 532 2243 536
rect 2311 532 2315 536
rect 2359 532 2363 536
rect 811 523 815 527
rect 1407 520 1411 524
rect 111 512 115 516
rect 339 515 343 519
rect 311 507 315 511
rect 463 507 467 511
rect 671 511 675 515
rect 831 515 835 519
rect 975 515 979 519
rect 983 515 987 519
rect 1447 520 1451 524
rect 1487 520 1491 524
rect 1535 520 1539 524
rect 1591 520 1595 524
rect 1647 520 1651 524
rect 1711 520 1715 524
rect 1783 520 1787 524
rect 1863 520 1867 524
rect 1943 520 1947 524
rect 2023 520 2027 524
rect 2103 520 2107 524
rect 2191 520 2195 524
rect 2287 520 2291 524
rect 2359 520 2363 524
rect 1239 512 1243 516
rect 1279 513 1283 517
rect 2407 513 2411 517
rect 1279 496 1283 500
rect 151 489 155 493
rect 223 489 227 493
rect 287 489 291 493
rect 351 489 355 493
rect 415 489 419 493
rect 479 489 483 493
rect 551 489 555 493
rect 623 489 627 493
rect 695 489 699 493
rect 767 489 771 493
rect 831 491 835 495
rect 1455 499 1459 503
rect 1495 499 1499 503
rect 1879 499 1883 503
rect 1951 499 1955 503
rect 1959 499 1963 503
rect 2039 499 2043 503
rect 2295 499 2299 503
rect 2303 499 2307 503
rect 2383 499 2384 503
rect 2384 499 2387 503
rect 2407 496 2411 500
rect 839 489 843 493
rect 919 489 923 493
rect 999 489 1003 493
rect 1079 489 1083 493
rect 1759 491 1763 495
rect 263 483 267 487
rect 311 483 312 487
rect 312 483 315 487
rect 579 483 580 487
rect 580 483 583 487
rect 671 483 675 487
rect 659 475 663 479
rect 983 483 987 487
rect 1095 483 1099 487
rect 1407 473 1411 477
rect 1447 473 1451 477
rect 1487 473 1491 477
rect 1535 473 1539 477
rect 1591 473 1595 477
rect 1647 473 1651 477
rect 1711 473 1715 477
rect 1783 473 1787 477
rect 1863 473 1867 477
rect 1943 473 1947 477
rect 2023 473 2027 477
rect 2103 473 2107 477
rect 2191 473 2195 477
rect 2287 473 2291 477
rect 2359 473 2363 477
rect 295 467 299 471
rect 239 459 243 463
rect 279 459 283 463
rect 319 463 323 467
rect 327 459 331 463
rect 375 463 379 467
rect 383 459 387 463
rect 407 463 408 467
rect 408 463 411 467
rect 439 459 443 463
rect 463 463 464 467
rect 464 463 467 467
rect 503 459 507 463
rect 515 463 519 467
rect 567 459 571 463
rect 579 463 583 467
rect 631 459 635 463
rect 687 463 691 467
rect 695 459 699 463
rect 751 463 755 467
rect 759 459 763 463
rect 815 463 819 467
rect 823 459 827 463
rect 879 463 883 467
rect 887 459 891 463
rect 899 463 903 467
rect 951 459 955 463
rect 975 463 976 467
rect 976 463 979 467
rect 1015 459 1019 463
rect 1027 463 1031 467
rect 1455 467 1459 471
rect 1495 467 1499 471
rect 1735 467 1736 471
rect 1736 467 1739 471
rect 1855 467 1859 471
rect 1879 467 1883 471
rect 1951 467 1955 471
rect 2123 467 2127 471
rect 2111 459 2115 463
rect 2295 467 2299 471
rect 2339 467 2343 471
rect 1303 443 1307 447
rect 1359 451 1363 455
rect 1343 443 1347 447
rect 1399 451 1403 455
rect 1383 443 1387 447
rect 1439 447 1443 451
rect 1447 443 1451 447
rect 1527 447 1531 451
rect 1535 443 1539 447
rect 1607 447 1611 451
rect 1631 443 1635 447
rect 1727 447 1731 451
rect 1735 443 1739 447
rect 1759 447 1760 451
rect 1760 447 1763 451
rect 1831 443 1835 447
rect 1911 447 1915 451
rect 1919 443 1923 447
rect 1979 447 1983 451
rect 2039 451 2043 455
rect 1999 443 2003 447
rect 2071 443 2075 447
rect 2127 447 2131 451
rect 2135 443 2139 447
rect 2191 447 2195 451
rect 2199 443 2203 447
rect 2247 447 2251 451
rect 2255 443 2259 447
rect 2311 447 2315 451
rect 2319 443 2323 447
rect 2347 447 2348 451
rect 2348 447 2351 451
rect 2359 443 2363 447
rect 2383 447 2384 451
rect 2384 447 2387 451
rect 111 436 115 440
rect 1239 436 1243 440
rect 263 431 264 435
rect 264 431 267 435
rect 295 431 299 435
rect 319 431 323 435
rect 375 431 379 435
rect 515 431 519 435
rect 575 431 579 435
rect 583 431 587 435
rect 659 431 660 435
rect 660 431 663 435
rect 687 431 691 435
rect 751 431 755 435
rect 815 431 819 435
rect 879 431 883 435
rect 1027 431 1031 435
rect 1055 431 1059 435
rect 111 419 115 423
rect 1239 419 1243 423
rect 1279 420 1283 424
rect 2347 423 2351 427
rect 2407 420 2411 424
rect 239 412 243 416
rect 279 412 283 416
rect 327 412 331 416
rect 383 412 387 416
rect 439 412 443 416
rect 503 412 507 416
rect 567 412 571 416
rect 631 412 635 416
rect 695 412 699 416
rect 759 412 763 416
rect 823 412 827 416
rect 887 412 891 416
rect 951 412 955 416
rect 1015 412 1019 416
rect 1351 415 1355 419
rect 1359 415 1363 419
rect 1399 415 1403 419
rect 1439 415 1443 419
rect 1527 415 1531 419
rect 1607 415 1611 419
rect 1727 415 1731 419
rect 1855 415 1856 419
rect 1856 415 1859 419
rect 1979 415 1983 419
rect 2111 415 2115 419
rect 2127 415 2131 419
rect 2191 415 2195 419
rect 2247 415 2251 419
rect 2347 415 2348 419
rect 2348 415 2351 419
rect 1279 403 1283 407
rect 2099 407 2103 411
rect 2407 403 2411 407
rect 143 396 147 400
rect 183 396 187 400
rect 223 396 227 400
rect 271 396 275 400
rect 335 396 339 400
rect 399 396 403 400
rect 471 396 475 400
rect 543 396 547 400
rect 615 396 619 400
rect 687 396 691 400
rect 751 396 755 400
rect 807 396 811 400
rect 863 396 867 400
rect 919 396 923 400
rect 975 396 979 400
rect 1031 396 1035 400
rect 1303 396 1307 400
rect 1343 396 1347 400
rect 1383 396 1387 400
rect 1447 396 1451 400
rect 1535 396 1539 400
rect 1631 396 1635 400
rect 1735 396 1739 400
rect 1831 396 1835 400
rect 1919 396 1923 400
rect 1999 396 2003 400
rect 2071 396 2075 400
rect 2135 396 2139 400
rect 2199 396 2203 400
rect 2255 396 2259 400
rect 2319 396 2323 400
rect 2359 396 2363 400
rect 111 389 115 393
rect 1239 389 1243 393
rect 111 372 115 376
rect 199 375 203 379
rect 239 375 243 379
rect 287 375 291 379
rect 407 383 411 387
rect 1359 384 1363 388
rect 1399 384 1403 388
rect 1439 384 1443 388
rect 1487 384 1491 388
rect 1543 384 1547 388
rect 1607 384 1611 388
rect 1679 384 1683 388
rect 1759 384 1763 388
rect 1839 384 1843 388
rect 1919 384 1923 388
rect 1999 384 2003 388
rect 2079 384 2083 388
rect 2159 384 2163 388
rect 2247 384 2251 388
rect 2335 384 2339 388
rect 507 375 511 379
rect 703 375 707 379
rect 767 375 771 379
rect 823 375 827 379
rect 879 375 883 379
rect 899 375 903 379
rect 907 375 911 379
rect 1279 377 1283 381
rect 2407 377 2411 381
rect 1239 372 1243 376
rect 463 367 467 371
rect 1279 360 1283 364
rect 1415 363 1419 367
rect 1455 363 1459 367
rect 1503 363 1507 367
rect 1559 363 1563 367
rect 1615 363 1619 367
rect 1855 363 1859 367
rect 1911 363 1915 367
rect 2175 363 2179 367
rect 2219 363 2223 367
rect 2227 363 2231 367
rect 2311 363 2315 367
rect 1703 355 1707 359
rect 2407 360 2411 364
rect 2023 355 2027 359
rect 143 349 147 353
rect 183 349 187 353
rect 223 349 227 353
rect 271 349 275 353
rect 335 349 339 353
rect 399 349 403 353
rect 471 349 475 353
rect 543 349 547 353
rect 199 343 203 347
rect 207 343 208 347
rect 208 343 211 347
rect 239 343 243 347
rect 287 343 291 347
rect 507 343 511 347
rect 583 347 587 351
rect 615 349 619 353
rect 687 349 691 353
rect 751 349 755 353
rect 807 349 811 353
rect 863 349 867 353
rect 919 349 923 353
rect 975 349 979 353
rect 1031 349 1035 353
rect 631 343 635 347
rect 703 343 707 347
rect 767 343 771 347
rect 823 343 827 347
rect 879 343 883 347
rect 1055 343 1056 347
rect 1056 343 1059 347
rect 1359 337 1363 341
rect 1399 337 1403 341
rect 1439 337 1443 341
rect 1487 337 1491 341
rect 1543 337 1547 341
rect 1607 337 1611 341
rect 1679 337 1683 341
rect 1759 337 1763 341
rect 1839 337 1843 341
rect 1919 337 1923 341
rect 1999 337 2003 341
rect 2079 337 2083 341
rect 2159 337 2163 341
rect 2247 337 2251 341
rect 2335 337 2339 341
rect 1351 331 1355 335
rect 1415 331 1419 335
rect 1455 331 1459 335
rect 1503 331 1507 335
rect 1559 331 1563 335
rect 1703 331 1704 335
rect 1704 331 1707 335
rect 1847 331 1851 335
rect 1855 331 1859 335
rect 2023 331 2024 335
rect 2024 331 2027 335
rect 2099 331 2103 335
rect 2175 331 2179 335
rect 2219 331 2223 335
rect 2347 331 2351 335
rect 135 311 139 315
rect 159 315 160 319
rect 160 315 163 319
rect 175 311 179 315
rect 231 319 235 323
rect 215 311 219 315
rect 243 315 244 319
rect 244 315 247 319
rect 255 311 259 315
rect 267 315 271 319
rect 295 311 299 315
rect 323 315 324 319
rect 324 315 327 319
rect 335 311 339 315
rect 383 315 387 319
rect 391 311 395 315
rect 439 315 443 319
rect 447 311 451 315
rect 463 315 467 319
rect 495 311 499 315
rect 535 315 539 319
rect 543 311 547 315
rect 591 311 595 315
rect 655 319 659 323
rect 639 311 643 315
rect 679 315 683 319
rect 687 311 691 315
rect 727 315 731 319
rect 735 311 739 315
rect 775 315 779 319
rect 783 311 787 315
rect 795 315 799 319
rect 839 311 843 315
rect 907 315 911 319
rect 863 303 867 307
rect 1511 299 1515 303
rect 1539 303 1540 307
rect 1540 303 1543 307
rect 1551 299 1555 303
rect 1599 307 1603 311
rect 1591 299 1595 303
rect 1615 303 1616 307
rect 1616 303 1619 307
rect 1631 299 1635 303
rect 1687 307 1691 311
rect 1671 299 1675 303
rect 1699 303 1700 307
rect 1700 303 1703 307
rect 1711 299 1715 303
rect 1767 307 1771 311
rect 1751 299 1755 303
rect 1779 303 1780 307
rect 1780 303 1783 307
rect 1791 299 1795 303
rect 111 288 115 292
rect 267 291 271 295
rect 323 291 327 295
rect 1239 288 1243 292
rect 1839 299 1843 303
rect 1895 303 1899 307
rect 1903 299 1907 303
rect 1959 303 1963 307
rect 1967 299 1971 303
rect 2027 303 2031 307
rect 2039 299 2043 303
rect 2111 303 2115 307
rect 2119 299 2123 303
rect 2131 303 2135 307
rect 2199 299 2203 303
rect 2227 303 2228 307
rect 2228 303 2231 307
rect 2279 299 2283 303
rect 2291 303 2295 307
rect 2359 299 2363 303
rect 2371 303 2375 307
rect 199 283 200 287
rect 200 283 203 287
rect 231 283 235 287
rect 251 283 255 287
rect 383 283 387 287
rect 439 283 443 287
rect 535 283 539 287
rect 631 283 635 287
rect 655 283 659 287
rect 679 283 683 287
rect 727 283 731 287
rect 775 283 779 287
rect 863 283 864 287
rect 864 283 867 287
rect 111 271 115 275
rect 151 275 155 279
rect 671 275 675 279
rect 1279 276 1283 280
rect 1539 279 1543 283
rect 1239 271 1243 275
rect 1699 279 1703 283
rect 1599 271 1603 275
rect 1679 271 1683 275
rect 1687 271 1691 275
rect 1779 279 1783 283
rect 1767 271 1771 275
rect 2407 276 2411 280
rect 1847 271 1851 275
rect 1895 271 1899 275
rect 1959 271 1963 275
rect 2027 271 2031 275
rect 2111 271 2115 275
rect 2291 271 2295 275
rect 2371 271 2375 275
rect 135 264 139 268
rect 175 264 179 268
rect 215 264 219 268
rect 255 264 259 268
rect 295 264 299 268
rect 335 264 339 268
rect 391 264 395 268
rect 447 264 451 268
rect 495 264 499 268
rect 543 264 547 268
rect 591 264 595 268
rect 639 264 643 268
rect 687 264 691 268
rect 735 264 739 268
rect 783 264 787 268
rect 839 264 843 268
rect 1279 259 1283 263
rect 2323 263 2327 267
rect 2407 259 2411 263
rect 1511 252 1515 256
rect 1551 252 1555 256
rect 1591 252 1595 256
rect 1631 252 1635 256
rect 1671 252 1675 256
rect 1711 252 1715 256
rect 1751 252 1755 256
rect 1791 252 1795 256
rect 1839 252 1843 256
rect 1903 252 1907 256
rect 1967 252 1971 256
rect 2039 252 2043 256
rect 2119 252 2123 256
rect 2199 252 2203 256
rect 2279 252 2283 256
rect 2359 252 2363 256
rect 135 244 139 248
rect 223 244 227 248
rect 311 244 315 248
rect 391 244 395 248
rect 463 244 467 248
rect 527 244 531 248
rect 591 244 595 248
rect 647 244 651 248
rect 695 244 699 248
rect 735 244 739 248
rect 783 244 787 248
rect 831 244 835 248
rect 879 244 883 248
rect 927 244 931 248
rect 975 244 979 248
rect 1023 244 1027 248
rect 111 237 115 241
rect 1239 237 1243 241
rect 1367 236 1371 240
rect 1407 236 1411 240
rect 1455 236 1459 240
rect 1511 236 1515 240
rect 1567 236 1571 240
rect 1631 236 1635 240
rect 1703 236 1707 240
rect 1775 236 1779 240
rect 1855 236 1859 240
rect 1943 236 1947 240
rect 2031 236 2035 240
rect 2119 236 2123 240
rect 2207 236 2211 240
rect 2295 236 2299 240
rect 2359 236 2363 240
rect 111 220 115 224
rect 159 223 160 227
rect 160 223 163 227
rect 287 223 291 227
rect 795 231 799 235
rect 1279 229 1283 233
rect 2407 229 2411 233
rect 743 223 747 227
rect 1239 220 1243 224
rect 2131 223 2135 227
rect 615 215 619 219
rect 1279 212 1283 216
rect 1415 215 1419 219
rect 2227 215 2231 219
rect 2375 215 2379 219
rect 2383 215 2384 219
rect 2384 215 2387 219
rect 2407 212 2411 216
rect 1671 207 1675 211
rect 135 197 139 201
rect 223 197 227 201
rect 311 197 315 201
rect 391 197 395 201
rect 463 197 467 201
rect 527 197 531 201
rect 591 197 595 201
rect 647 197 651 201
rect 695 197 699 201
rect 735 197 739 201
rect 783 197 787 201
rect 831 197 835 201
rect 879 197 883 201
rect 927 197 931 201
rect 975 197 979 201
rect 1023 197 1027 201
rect 151 191 155 195
rect 287 191 291 195
rect 671 191 672 195
rect 672 191 675 195
rect 743 191 747 195
rect 1039 191 1043 195
rect 1367 189 1371 193
rect 1407 189 1411 193
rect 1455 189 1459 193
rect 1511 189 1515 193
rect 1567 189 1571 193
rect 1631 189 1635 193
rect 1703 189 1707 193
rect 1775 189 1779 193
rect 1855 189 1859 193
rect 1943 189 1947 193
rect 2031 189 2035 193
rect 2119 189 2123 193
rect 2207 189 2211 193
rect 2295 189 2299 193
rect 2359 189 2363 193
rect 1415 183 1419 187
rect 1679 183 1683 187
rect 1739 175 1743 179
rect 2263 183 2267 187
rect 2323 183 2324 187
rect 2324 183 2327 187
rect 2375 183 2379 187
rect 1303 151 1307 155
rect 1331 155 1332 159
rect 1332 155 1335 159
rect 1343 151 1347 155
rect 1371 155 1372 159
rect 1372 155 1375 159
rect 1383 151 1387 155
rect 1411 155 1412 159
rect 1412 155 1415 159
rect 1423 151 1427 155
rect 1451 155 1452 159
rect 1452 155 1455 159
rect 1463 151 1467 155
rect 1511 155 1515 159
rect 1519 151 1523 155
rect 1575 155 1579 159
rect 1583 151 1587 155
rect 1639 155 1643 159
rect 1647 151 1651 155
rect 1671 155 1672 159
rect 1672 155 1675 159
rect 1711 151 1715 155
rect 1767 155 1771 159
rect 1775 151 1779 155
rect 1823 155 1827 159
rect 1831 151 1835 155
rect 1879 155 1883 159
rect 1887 151 1891 155
rect 1927 155 1931 159
rect 1935 151 1939 155
rect 1963 155 1964 159
rect 1964 155 1967 159
rect 1975 151 1979 155
rect 2023 159 2027 163
rect 2015 151 2019 155
rect 2071 159 2075 163
rect 2055 151 2059 155
rect 2103 159 2107 163
rect 2095 151 2099 155
rect 2135 155 2139 159
rect 2143 151 2147 155
rect 2183 155 2187 159
rect 2191 151 2195 155
rect 2227 155 2231 159
rect 2239 151 2243 155
rect 2287 159 2291 163
rect 2279 151 2283 155
rect 2335 159 2339 163
rect 2319 151 2323 155
rect 2367 159 2371 163
rect 2359 151 2363 155
rect 2383 155 2384 159
rect 2384 155 2387 159
rect 151 135 155 139
rect 179 139 180 143
rect 180 139 183 143
rect 191 135 195 139
rect 219 139 220 143
rect 220 139 223 143
rect 231 135 235 139
rect 259 139 260 143
rect 260 139 263 143
rect 271 135 275 139
rect 299 139 300 143
rect 300 139 303 143
rect 311 135 315 139
rect 339 139 340 143
rect 340 139 343 143
rect 351 135 355 139
rect 379 139 380 143
rect 380 139 383 143
rect 391 135 395 139
rect 447 143 451 147
rect 431 135 435 139
rect 459 139 460 143
rect 460 139 463 143
rect 471 135 475 139
rect 499 139 500 143
rect 500 139 503 143
rect 511 135 515 139
rect 539 139 540 143
rect 540 139 543 143
rect 551 135 555 139
rect 579 139 580 143
rect 580 139 583 143
rect 591 135 595 139
rect 615 139 616 143
rect 616 139 619 143
rect 631 135 635 139
rect 659 139 660 143
rect 660 139 663 143
rect 671 135 675 139
rect 699 139 700 143
rect 700 139 703 143
rect 711 135 715 139
rect 739 139 740 143
rect 740 139 743 143
rect 751 135 755 139
rect 779 139 780 143
rect 780 139 783 143
rect 791 135 795 139
rect 819 139 820 143
rect 820 139 823 143
rect 831 135 835 139
rect 859 139 860 143
rect 860 139 863 143
rect 871 135 875 139
rect 899 139 900 143
rect 900 139 903 143
rect 911 135 915 139
rect 939 139 940 143
rect 940 139 943 143
rect 951 135 955 139
rect 979 139 980 143
rect 980 139 983 143
rect 991 135 995 139
rect 1019 139 1020 143
rect 1020 139 1023 143
rect 1031 135 1035 139
rect 1059 139 1060 143
rect 1060 139 1063 143
rect 1071 135 1075 139
rect 1099 139 1100 143
rect 1100 139 1103 143
rect 1111 135 1115 139
rect 1167 143 1171 147
rect 1151 135 1155 139
rect 1199 143 1203 147
rect 1191 135 1195 139
rect 1279 128 1283 132
rect 1963 131 1967 135
rect 2407 128 2411 132
rect 1339 123 1343 127
rect 1379 123 1383 127
rect 1419 123 1423 127
rect 1459 123 1463 127
rect 1511 123 1515 127
rect 1575 123 1579 127
rect 1639 123 1643 127
rect 1739 123 1740 127
rect 1740 123 1743 127
rect 1767 123 1771 127
rect 1823 123 1827 127
rect 1879 123 1883 127
rect 1927 123 1931 127
rect 2023 123 2027 127
rect 2071 123 2075 127
rect 2103 123 2107 127
rect 2135 123 2139 127
rect 2183 123 2187 127
rect 2263 123 2264 127
rect 2264 123 2267 127
rect 2287 123 2291 127
rect 2335 123 2339 127
rect 2367 123 2371 127
rect 111 112 115 116
rect 299 115 303 119
rect 179 107 183 111
rect 227 107 231 111
rect 267 107 271 111
rect 1239 112 1243 116
rect 347 107 351 111
rect 387 107 391 111
rect 447 107 451 111
rect 467 107 471 111
rect 507 107 511 111
rect 547 107 551 111
rect 587 107 591 111
rect 651 107 655 111
rect 667 107 671 111
rect 707 107 711 111
rect 747 107 751 111
rect 787 107 791 111
rect 827 107 831 111
rect 867 107 871 111
rect 907 107 911 111
rect 947 107 951 111
rect 987 107 991 111
rect 1027 107 1031 111
rect 1067 107 1071 111
rect 1107 107 1111 111
rect 1167 107 1171 111
rect 1199 107 1203 111
rect 1279 111 1283 115
rect 2407 111 2411 115
rect 1303 104 1307 108
rect 1343 104 1347 108
rect 1383 104 1387 108
rect 1423 104 1427 108
rect 1463 104 1467 108
rect 1519 104 1523 108
rect 1583 104 1587 108
rect 1647 104 1651 108
rect 1711 104 1715 108
rect 1775 104 1779 108
rect 1831 104 1835 108
rect 1887 104 1891 108
rect 1935 104 1939 108
rect 1975 104 1979 108
rect 2015 104 2019 108
rect 2055 104 2059 108
rect 2095 104 2099 108
rect 2143 104 2147 108
rect 2191 104 2195 108
rect 2239 104 2243 108
rect 2279 104 2283 108
rect 2319 104 2323 108
rect 2359 104 2363 108
rect 111 95 115 99
rect 1239 95 1243 99
rect 151 88 155 92
rect 191 88 195 92
rect 231 88 235 92
rect 271 88 275 92
rect 311 88 315 92
rect 351 88 355 92
rect 391 88 395 92
rect 431 88 435 92
rect 471 88 475 92
rect 511 88 515 92
rect 551 88 555 92
rect 591 88 595 92
rect 631 88 635 92
rect 671 88 675 92
rect 711 88 715 92
rect 751 88 755 92
rect 791 88 795 92
rect 831 88 835 92
rect 871 88 875 92
rect 911 88 915 92
rect 951 88 955 92
rect 991 88 995 92
rect 1031 88 1035 92
rect 1071 88 1075 92
rect 1111 88 1115 92
rect 1151 88 1155 92
rect 1191 88 1195 92
<< m3 >>
rect 111 2494 115 2495
rect 111 2489 115 2490
rect 231 2494 235 2495
rect 231 2489 235 2490
rect 271 2494 275 2495
rect 271 2489 275 2490
rect 311 2494 315 2495
rect 311 2489 315 2490
rect 351 2494 355 2495
rect 351 2489 355 2490
rect 399 2494 403 2495
rect 399 2489 403 2490
rect 455 2494 459 2495
rect 455 2489 459 2490
rect 511 2494 515 2495
rect 511 2489 515 2490
rect 575 2494 579 2495
rect 575 2489 579 2490
rect 639 2494 643 2495
rect 639 2489 643 2490
rect 703 2494 707 2495
rect 703 2489 707 2490
rect 767 2494 771 2495
rect 767 2489 771 2490
rect 823 2494 827 2495
rect 823 2489 827 2490
rect 879 2494 883 2495
rect 879 2489 883 2490
rect 927 2494 931 2495
rect 927 2489 931 2490
rect 975 2494 979 2495
rect 975 2489 979 2490
rect 1023 2494 1027 2495
rect 1023 2489 1027 2490
rect 1071 2494 1075 2495
rect 1071 2489 1075 2490
rect 1111 2494 1115 2495
rect 1111 2489 1115 2490
rect 1151 2494 1155 2495
rect 1151 2489 1155 2490
rect 1191 2494 1195 2495
rect 1191 2489 1195 2490
rect 1239 2494 1243 2495
rect 1239 2489 1243 2490
rect 1279 2490 1283 2491
rect 112 2457 114 2489
rect 232 2480 234 2489
rect 258 2483 264 2484
rect 230 2479 236 2480
rect 230 2475 231 2479
rect 235 2475 236 2479
rect 258 2479 259 2483
rect 263 2479 264 2483
rect 272 2480 274 2489
rect 312 2480 314 2489
rect 326 2487 332 2488
rect 326 2483 327 2487
rect 331 2483 332 2487
rect 326 2482 332 2483
rect 258 2478 264 2479
rect 270 2479 276 2480
rect 230 2474 236 2475
rect 110 2456 116 2457
rect 110 2452 111 2456
rect 115 2452 116 2456
rect 110 2451 116 2452
rect 242 2451 248 2452
rect 242 2447 243 2451
rect 247 2447 248 2451
rect 260 2450 262 2478
rect 270 2475 271 2479
rect 275 2475 276 2479
rect 270 2474 276 2475
rect 310 2479 316 2480
rect 310 2475 311 2479
rect 315 2475 316 2479
rect 310 2474 316 2475
rect 328 2452 330 2482
rect 352 2480 354 2489
rect 358 2487 364 2488
rect 358 2483 359 2487
rect 363 2483 364 2487
rect 358 2482 364 2483
rect 390 2483 396 2484
rect 350 2479 356 2480
rect 350 2475 351 2479
rect 355 2475 356 2479
rect 350 2474 356 2475
rect 360 2452 362 2482
rect 390 2479 391 2483
rect 395 2479 396 2483
rect 400 2480 402 2489
rect 446 2483 452 2484
rect 390 2478 396 2479
rect 398 2479 404 2480
rect 392 2452 394 2478
rect 398 2475 399 2479
rect 403 2475 404 2479
rect 446 2479 447 2483
rect 451 2479 452 2483
rect 456 2480 458 2489
rect 502 2483 508 2484
rect 446 2478 452 2479
rect 454 2479 460 2480
rect 398 2474 404 2475
rect 448 2452 450 2478
rect 454 2475 455 2479
rect 459 2475 460 2479
rect 502 2479 503 2483
rect 507 2479 508 2483
rect 512 2480 514 2489
rect 566 2483 572 2484
rect 502 2478 508 2479
rect 510 2479 516 2480
rect 454 2474 460 2475
rect 504 2452 506 2478
rect 510 2475 511 2479
rect 515 2475 516 2479
rect 566 2479 567 2483
rect 571 2479 572 2483
rect 576 2480 578 2489
rect 630 2483 636 2484
rect 566 2478 572 2479
rect 574 2479 580 2480
rect 510 2474 516 2475
rect 568 2452 570 2478
rect 574 2475 575 2479
rect 579 2475 580 2479
rect 630 2479 631 2483
rect 635 2479 636 2483
rect 640 2480 642 2489
rect 650 2483 656 2484
rect 630 2478 636 2479
rect 638 2479 644 2480
rect 574 2474 580 2475
rect 632 2452 634 2478
rect 638 2475 639 2479
rect 643 2475 644 2479
rect 650 2479 651 2483
rect 655 2479 656 2483
rect 704 2480 706 2489
rect 768 2480 770 2489
rect 782 2487 788 2488
rect 782 2483 783 2487
rect 787 2483 788 2487
rect 782 2482 788 2483
rect 814 2483 820 2484
rect 650 2478 656 2479
rect 702 2479 708 2480
rect 638 2474 644 2475
rect 266 2451 272 2452
rect 266 2450 267 2451
rect 260 2448 267 2450
rect 242 2446 248 2447
rect 266 2447 267 2448
rect 271 2447 272 2451
rect 266 2446 272 2447
rect 326 2451 332 2452
rect 326 2447 327 2451
rect 331 2447 332 2451
rect 326 2446 332 2447
rect 358 2451 364 2452
rect 358 2447 359 2451
rect 363 2447 364 2451
rect 358 2446 364 2447
rect 390 2451 396 2452
rect 390 2447 391 2451
rect 395 2447 396 2451
rect 390 2446 396 2447
rect 446 2451 452 2452
rect 446 2447 447 2451
rect 451 2447 452 2451
rect 446 2446 452 2447
rect 502 2451 508 2452
rect 502 2447 503 2451
rect 507 2447 508 2451
rect 502 2446 508 2447
rect 566 2451 572 2452
rect 566 2447 567 2451
rect 571 2447 572 2451
rect 566 2446 572 2447
rect 630 2451 636 2452
rect 630 2447 631 2451
rect 635 2447 636 2451
rect 630 2446 636 2447
rect 110 2439 116 2440
rect 110 2435 111 2439
rect 115 2435 116 2439
rect 110 2434 116 2435
rect 112 2419 114 2434
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 232 2419 234 2427
rect 111 2418 115 2419
rect 111 2413 115 2414
rect 199 2418 203 2419
rect 199 2413 203 2414
rect 231 2418 235 2419
rect 231 2413 235 2414
rect 112 2406 114 2413
rect 198 2412 204 2413
rect 198 2408 199 2412
rect 203 2408 204 2412
rect 198 2407 204 2408
rect 110 2405 116 2406
rect 110 2401 111 2405
rect 115 2401 116 2405
rect 110 2400 116 2401
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 112 2347 114 2383
rect 198 2365 204 2366
rect 198 2361 199 2365
rect 203 2361 204 2365
rect 198 2360 204 2361
rect 244 2360 246 2446
rect 270 2432 276 2433
rect 270 2428 271 2432
rect 275 2428 276 2432
rect 270 2427 276 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 350 2432 356 2433
rect 350 2428 351 2432
rect 355 2428 356 2432
rect 350 2427 356 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 454 2432 460 2433
rect 454 2428 455 2432
rect 459 2428 460 2432
rect 454 2427 460 2428
rect 510 2432 516 2433
rect 510 2428 511 2432
rect 515 2428 516 2432
rect 510 2427 516 2428
rect 574 2432 580 2433
rect 574 2428 575 2432
rect 579 2428 580 2432
rect 574 2427 580 2428
rect 638 2432 644 2433
rect 638 2428 639 2432
rect 643 2428 644 2432
rect 638 2427 644 2428
rect 272 2419 274 2427
rect 312 2419 314 2427
rect 352 2419 354 2427
rect 400 2419 402 2427
rect 456 2419 458 2427
rect 512 2419 514 2427
rect 576 2419 578 2427
rect 640 2419 642 2427
rect 263 2418 267 2419
rect 263 2413 267 2414
rect 271 2418 275 2419
rect 271 2413 275 2414
rect 311 2418 315 2419
rect 311 2413 315 2414
rect 327 2418 331 2419
rect 327 2413 331 2414
rect 351 2418 355 2419
rect 351 2413 355 2414
rect 399 2418 403 2419
rect 399 2413 403 2414
rect 455 2418 459 2419
rect 455 2413 459 2414
rect 471 2418 475 2419
rect 471 2413 475 2414
rect 511 2418 515 2419
rect 511 2413 515 2414
rect 543 2418 547 2419
rect 543 2413 547 2414
rect 575 2418 579 2419
rect 575 2413 579 2414
rect 615 2418 619 2419
rect 615 2413 619 2414
rect 639 2418 643 2419
rect 639 2413 643 2414
rect 262 2412 268 2413
rect 262 2408 263 2412
rect 267 2408 268 2412
rect 262 2407 268 2408
rect 326 2412 332 2413
rect 326 2408 327 2412
rect 331 2408 332 2412
rect 326 2407 332 2408
rect 398 2412 404 2413
rect 398 2408 399 2412
rect 403 2408 404 2412
rect 398 2407 404 2408
rect 470 2412 476 2413
rect 470 2408 471 2412
rect 475 2408 476 2412
rect 470 2407 476 2408
rect 542 2412 548 2413
rect 542 2408 543 2412
rect 547 2408 548 2412
rect 542 2407 548 2408
rect 614 2412 620 2413
rect 614 2408 615 2412
rect 619 2408 620 2412
rect 614 2407 620 2408
rect 652 2400 654 2478
rect 702 2475 703 2479
rect 707 2475 708 2479
rect 702 2474 708 2475
rect 766 2479 772 2480
rect 766 2475 767 2479
rect 771 2475 772 2479
rect 766 2474 772 2475
rect 784 2452 786 2482
rect 814 2479 815 2483
rect 819 2479 820 2483
rect 824 2480 826 2489
rect 870 2483 876 2484
rect 814 2478 820 2479
rect 822 2479 828 2480
rect 816 2452 818 2478
rect 822 2475 823 2479
rect 827 2475 828 2479
rect 870 2479 871 2483
rect 875 2479 876 2483
rect 880 2480 882 2489
rect 918 2483 924 2484
rect 870 2478 876 2479
rect 878 2479 884 2480
rect 822 2474 828 2475
rect 872 2452 874 2478
rect 878 2475 879 2479
rect 883 2475 884 2479
rect 918 2479 919 2483
rect 923 2479 924 2483
rect 928 2480 930 2489
rect 966 2483 972 2484
rect 918 2478 924 2479
rect 926 2479 932 2480
rect 878 2474 884 2475
rect 920 2452 922 2478
rect 926 2475 927 2479
rect 931 2475 932 2479
rect 966 2479 967 2483
rect 971 2479 972 2483
rect 976 2480 978 2489
rect 1014 2483 1020 2484
rect 966 2478 972 2479
rect 974 2479 980 2480
rect 926 2474 932 2475
rect 968 2452 970 2478
rect 974 2475 975 2479
rect 979 2475 980 2479
rect 1014 2479 1015 2483
rect 1019 2479 1020 2483
rect 1024 2480 1026 2489
rect 1062 2483 1068 2484
rect 1014 2478 1020 2479
rect 1022 2479 1028 2480
rect 974 2474 980 2475
rect 1016 2452 1018 2478
rect 1022 2475 1023 2479
rect 1027 2475 1028 2479
rect 1062 2479 1063 2483
rect 1067 2479 1068 2483
rect 1072 2480 1074 2489
rect 1112 2480 1114 2489
rect 1126 2487 1132 2488
rect 1126 2483 1127 2487
rect 1131 2483 1132 2487
rect 1126 2482 1132 2483
rect 1062 2478 1068 2479
rect 1070 2479 1076 2480
rect 1022 2474 1028 2475
rect 1064 2452 1066 2478
rect 1070 2475 1071 2479
rect 1075 2475 1076 2479
rect 1070 2474 1076 2475
rect 1110 2479 1116 2480
rect 1110 2475 1111 2479
rect 1115 2475 1116 2479
rect 1110 2474 1116 2475
rect 1128 2452 1130 2482
rect 1152 2480 1154 2489
rect 1166 2487 1172 2488
rect 1166 2483 1167 2487
rect 1171 2483 1172 2487
rect 1166 2482 1172 2483
rect 1150 2479 1156 2480
rect 1150 2475 1151 2479
rect 1155 2475 1156 2479
rect 1150 2474 1156 2475
rect 1168 2452 1170 2482
rect 1192 2480 1194 2489
rect 1202 2487 1208 2488
rect 1202 2483 1203 2487
rect 1207 2483 1208 2487
rect 1202 2482 1208 2483
rect 1190 2479 1196 2480
rect 1190 2475 1191 2479
rect 1195 2475 1196 2479
rect 1190 2474 1196 2475
rect 1204 2452 1206 2482
rect 1240 2457 1242 2489
rect 1279 2485 1283 2486
rect 1303 2490 1307 2491
rect 1303 2485 1307 2486
rect 1343 2490 1347 2491
rect 1343 2485 1347 2486
rect 1383 2490 1387 2491
rect 1383 2485 1387 2486
rect 1439 2490 1443 2491
rect 1439 2485 1443 2486
rect 1511 2490 1515 2491
rect 1511 2485 1515 2486
rect 1583 2490 1587 2491
rect 1583 2485 1587 2486
rect 1663 2490 1667 2491
rect 1663 2485 1667 2486
rect 1735 2490 1739 2491
rect 1735 2485 1739 2486
rect 1807 2490 1811 2491
rect 1807 2485 1811 2486
rect 1887 2490 1891 2491
rect 1887 2485 1891 2486
rect 1967 2490 1971 2491
rect 1967 2485 1971 2486
rect 2063 2490 2067 2491
rect 2063 2485 2067 2486
rect 2167 2490 2171 2491
rect 2167 2485 2171 2486
rect 2271 2490 2275 2491
rect 2271 2485 2275 2486
rect 2359 2490 2363 2491
rect 2359 2485 2363 2486
rect 2407 2490 2411 2491
rect 2407 2485 2411 2486
rect 1238 2456 1244 2457
rect 1238 2452 1239 2456
rect 1243 2452 1244 2456
rect 1280 2453 1282 2485
rect 1304 2476 1306 2485
rect 1318 2483 1324 2484
rect 1318 2479 1319 2483
rect 1323 2479 1324 2483
rect 1318 2478 1324 2479
rect 1302 2475 1308 2476
rect 1302 2471 1303 2475
rect 1307 2471 1308 2475
rect 1302 2470 1308 2471
rect 774 2451 780 2452
rect 774 2447 775 2451
rect 779 2447 780 2451
rect 774 2446 780 2447
rect 782 2451 788 2452
rect 782 2447 783 2451
rect 787 2447 788 2451
rect 782 2446 788 2447
rect 814 2451 820 2452
rect 814 2447 815 2451
rect 819 2447 820 2451
rect 814 2446 820 2447
rect 870 2451 876 2452
rect 870 2447 871 2451
rect 875 2447 876 2451
rect 870 2446 876 2447
rect 918 2451 924 2452
rect 918 2447 919 2451
rect 923 2447 924 2451
rect 918 2446 924 2447
rect 966 2451 972 2452
rect 966 2447 967 2451
rect 971 2447 972 2451
rect 966 2446 972 2447
rect 1014 2451 1020 2452
rect 1014 2447 1015 2451
rect 1019 2447 1020 2451
rect 1014 2446 1020 2447
rect 1062 2451 1068 2452
rect 1062 2447 1063 2451
rect 1067 2447 1068 2451
rect 1062 2446 1068 2447
rect 1126 2451 1132 2452
rect 1126 2447 1127 2451
rect 1131 2447 1132 2451
rect 1126 2446 1132 2447
rect 1166 2451 1172 2452
rect 1166 2447 1167 2451
rect 1171 2447 1172 2451
rect 1166 2446 1172 2447
rect 1202 2451 1208 2452
rect 1238 2451 1244 2452
rect 1278 2452 1284 2453
rect 1202 2447 1203 2451
rect 1207 2447 1208 2451
rect 1278 2448 1279 2452
rect 1283 2448 1284 2452
rect 1320 2448 1322 2478
rect 1344 2476 1346 2485
rect 1358 2483 1364 2484
rect 1358 2479 1359 2483
rect 1363 2479 1364 2483
rect 1358 2478 1364 2479
rect 1342 2475 1348 2476
rect 1342 2471 1343 2475
rect 1347 2471 1348 2475
rect 1342 2470 1348 2471
rect 1360 2448 1362 2478
rect 1384 2476 1386 2485
rect 1398 2483 1404 2484
rect 1398 2479 1399 2483
rect 1403 2479 1404 2483
rect 1398 2478 1404 2479
rect 1430 2479 1436 2480
rect 1382 2475 1388 2476
rect 1382 2471 1383 2475
rect 1387 2471 1388 2475
rect 1382 2470 1388 2471
rect 1400 2448 1402 2478
rect 1430 2475 1431 2479
rect 1435 2475 1436 2479
rect 1440 2476 1442 2485
rect 1502 2479 1508 2480
rect 1430 2474 1436 2475
rect 1438 2475 1444 2476
rect 1432 2448 1434 2474
rect 1438 2471 1439 2475
rect 1443 2471 1444 2475
rect 1502 2475 1503 2479
rect 1507 2475 1508 2479
rect 1512 2476 1514 2485
rect 1574 2479 1580 2480
rect 1502 2474 1508 2475
rect 1510 2475 1516 2476
rect 1438 2470 1444 2471
rect 1504 2448 1506 2474
rect 1510 2471 1511 2475
rect 1515 2471 1516 2475
rect 1574 2475 1575 2479
rect 1579 2475 1580 2479
rect 1584 2476 1586 2485
rect 1654 2479 1660 2480
rect 1574 2474 1580 2475
rect 1582 2475 1588 2476
rect 1510 2470 1516 2471
rect 1576 2448 1578 2474
rect 1582 2471 1583 2475
rect 1587 2471 1588 2475
rect 1654 2475 1655 2479
rect 1659 2475 1660 2479
rect 1664 2476 1666 2485
rect 1686 2479 1692 2480
rect 1654 2474 1660 2475
rect 1662 2475 1668 2476
rect 1582 2470 1588 2471
rect 1656 2448 1658 2474
rect 1662 2471 1663 2475
rect 1667 2471 1668 2475
rect 1686 2475 1687 2479
rect 1691 2475 1692 2479
rect 1736 2476 1738 2485
rect 1798 2479 1804 2480
rect 1686 2474 1692 2475
rect 1734 2475 1740 2476
rect 1662 2470 1668 2471
rect 1278 2447 1284 2448
rect 1318 2447 1324 2448
rect 1202 2446 1208 2447
rect 702 2432 708 2433
rect 702 2428 703 2432
rect 707 2428 708 2432
rect 702 2427 708 2428
rect 766 2432 772 2433
rect 766 2428 767 2432
rect 771 2428 772 2432
rect 766 2427 772 2428
rect 704 2419 706 2427
rect 768 2419 770 2427
rect 687 2418 691 2419
rect 687 2413 691 2414
rect 703 2418 707 2419
rect 703 2413 707 2414
rect 751 2418 755 2419
rect 751 2413 755 2414
rect 767 2418 771 2419
rect 767 2413 771 2414
rect 686 2412 692 2413
rect 686 2408 687 2412
rect 691 2408 692 2412
rect 686 2407 692 2408
rect 750 2412 756 2413
rect 750 2408 751 2412
rect 755 2408 756 2412
rect 750 2407 756 2408
rect 650 2399 656 2400
rect 650 2395 651 2399
rect 655 2395 656 2399
rect 650 2394 656 2395
rect 278 2391 284 2392
rect 278 2387 279 2391
rect 283 2387 284 2391
rect 278 2386 284 2387
rect 342 2391 348 2392
rect 342 2387 343 2391
rect 347 2387 348 2391
rect 342 2386 348 2387
rect 414 2391 420 2392
rect 414 2387 415 2391
rect 419 2387 420 2391
rect 414 2386 420 2387
rect 422 2391 428 2392
rect 422 2387 423 2391
rect 427 2387 428 2391
rect 422 2386 428 2387
rect 262 2365 268 2366
rect 262 2361 263 2365
rect 267 2361 268 2365
rect 262 2360 268 2361
rect 280 2360 282 2386
rect 326 2365 332 2366
rect 326 2361 327 2365
rect 331 2361 332 2365
rect 326 2360 332 2361
rect 344 2360 346 2386
rect 398 2365 404 2366
rect 398 2361 399 2365
rect 403 2361 404 2365
rect 398 2360 404 2361
rect 416 2360 418 2386
rect 200 2347 202 2360
rect 242 2359 248 2360
rect 242 2355 243 2359
rect 247 2355 248 2359
rect 242 2354 248 2355
rect 264 2347 266 2360
rect 278 2359 284 2360
rect 278 2355 279 2359
rect 283 2355 284 2359
rect 278 2354 284 2355
rect 328 2347 330 2360
rect 342 2359 348 2360
rect 342 2355 343 2359
rect 347 2355 348 2359
rect 342 2354 348 2355
rect 400 2347 402 2360
rect 414 2359 420 2360
rect 414 2355 415 2359
rect 419 2355 420 2359
rect 414 2354 420 2355
rect 111 2346 115 2347
rect 111 2341 115 2342
rect 199 2346 203 2347
rect 199 2341 203 2342
rect 263 2346 267 2347
rect 263 2341 267 2342
rect 271 2346 275 2347
rect 271 2341 275 2342
rect 327 2346 331 2347
rect 327 2341 331 2342
rect 399 2346 403 2347
rect 399 2341 403 2342
rect 112 2309 114 2341
rect 272 2332 274 2341
rect 318 2335 324 2336
rect 270 2331 276 2332
rect 270 2327 271 2331
rect 275 2327 276 2331
rect 318 2331 319 2335
rect 323 2331 324 2335
rect 328 2332 330 2341
rect 390 2335 396 2336
rect 318 2330 324 2331
rect 326 2331 332 2332
rect 270 2326 276 2327
rect 110 2308 116 2309
rect 110 2304 111 2308
rect 115 2304 116 2308
rect 320 2304 322 2330
rect 326 2327 327 2331
rect 331 2327 332 2331
rect 390 2331 391 2335
rect 395 2331 396 2335
rect 400 2332 402 2341
rect 424 2336 426 2386
rect 470 2365 476 2366
rect 470 2361 471 2365
rect 475 2361 476 2365
rect 470 2360 476 2361
rect 542 2365 548 2366
rect 542 2361 543 2365
rect 547 2361 548 2365
rect 542 2360 548 2361
rect 614 2365 620 2366
rect 614 2361 615 2365
rect 619 2361 620 2365
rect 614 2360 620 2361
rect 686 2365 692 2366
rect 686 2361 687 2365
rect 691 2361 692 2365
rect 686 2360 692 2361
rect 750 2365 756 2366
rect 750 2361 751 2365
rect 755 2361 756 2365
rect 750 2360 756 2361
rect 776 2360 778 2446
rect 1318 2443 1319 2447
rect 1323 2443 1324 2447
rect 1318 2442 1324 2443
rect 1358 2447 1364 2448
rect 1358 2443 1359 2447
rect 1363 2443 1364 2447
rect 1358 2442 1364 2443
rect 1398 2447 1404 2448
rect 1398 2443 1399 2447
rect 1403 2443 1404 2447
rect 1398 2442 1404 2443
rect 1430 2447 1436 2448
rect 1430 2443 1431 2447
rect 1435 2443 1436 2447
rect 1430 2442 1436 2443
rect 1502 2447 1508 2448
rect 1502 2443 1503 2447
rect 1507 2443 1508 2447
rect 1502 2442 1508 2443
rect 1574 2447 1580 2448
rect 1574 2443 1575 2447
rect 1579 2443 1580 2447
rect 1574 2442 1580 2443
rect 1654 2447 1660 2448
rect 1654 2443 1655 2447
rect 1659 2443 1660 2447
rect 1654 2442 1660 2443
rect 1238 2439 1244 2440
rect 1238 2435 1239 2439
rect 1243 2435 1244 2439
rect 1238 2434 1244 2435
rect 1278 2435 1284 2436
rect 822 2432 828 2433
rect 822 2428 823 2432
rect 827 2428 828 2432
rect 822 2427 828 2428
rect 878 2432 884 2433
rect 878 2428 879 2432
rect 883 2428 884 2432
rect 878 2427 884 2428
rect 926 2432 932 2433
rect 926 2428 927 2432
rect 931 2428 932 2432
rect 926 2427 932 2428
rect 974 2432 980 2433
rect 974 2428 975 2432
rect 979 2428 980 2432
rect 974 2427 980 2428
rect 1022 2432 1028 2433
rect 1022 2428 1023 2432
rect 1027 2428 1028 2432
rect 1022 2427 1028 2428
rect 1070 2432 1076 2433
rect 1070 2428 1071 2432
rect 1075 2428 1076 2432
rect 1070 2427 1076 2428
rect 1110 2432 1116 2433
rect 1110 2428 1111 2432
rect 1115 2428 1116 2432
rect 1110 2427 1116 2428
rect 1150 2432 1156 2433
rect 1150 2428 1151 2432
rect 1155 2428 1156 2432
rect 1150 2427 1156 2428
rect 1190 2432 1196 2433
rect 1190 2428 1191 2432
rect 1195 2428 1196 2432
rect 1190 2427 1196 2428
rect 824 2419 826 2427
rect 880 2419 882 2427
rect 928 2419 930 2427
rect 976 2419 978 2427
rect 1024 2419 1026 2427
rect 1072 2419 1074 2427
rect 1112 2419 1114 2427
rect 1152 2419 1154 2427
rect 1192 2419 1194 2427
rect 1240 2419 1242 2434
rect 1278 2431 1279 2435
rect 1283 2431 1284 2435
rect 1278 2430 1284 2431
rect 1280 2423 1282 2430
rect 1302 2428 1308 2429
rect 1302 2424 1303 2428
rect 1307 2424 1308 2428
rect 1302 2423 1308 2424
rect 1342 2428 1348 2429
rect 1342 2424 1343 2428
rect 1347 2424 1348 2428
rect 1342 2423 1348 2424
rect 1382 2428 1388 2429
rect 1382 2424 1383 2428
rect 1387 2424 1388 2428
rect 1382 2423 1388 2424
rect 1438 2428 1444 2429
rect 1438 2424 1439 2428
rect 1443 2424 1444 2428
rect 1438 2423 1444 2424
rect 1510 2428 1516 2429
rect 1510 2424 1511 2428
rect 1515 2424 1516 2428
rect 1510 2423 1516 2424
rect 1582 2428 1588 2429
rect 1582 2424 1583 2428
rect 1587 2424 1588 2428
rect 1582 2423 1588 2424
rect 1662 2428 1668 2429
rect 1662 2424 1663 2428
rect 1667 2424 1668 2428
rect 1662 2423 1668 2424
rect 1279 2422 1283 2423
rect 823 2418 827 2419
rect 823 2413 827 2414
rect 879 2418 883 2419
rect 879 2413 883 2414
rect 895 2418 899 2419
rect 895 2413 899 2414
rect 927 2418 931 2419
rect 927 2413 931 2414
rect 967 2418 971 2419
rect 967 2413 971 2414
rect 975 2418 979 2419
rect 975 2413 979 2414
rect 1023 2418 1027 2419
rect 1023 2413 1027 2414
rect 1071 2418 1075 2419
rect 1071 2413 1075 2414
rect 1111 2418 1115 2419
rect 1111 2413 1115 2414
rect 1151 2418 1155 2419
rect 1151 2413 1155 2414
rect 1191 2418 1195 2419
rect 1191 2413 1195 2414
rect 1239 2418 1243 2419
rect 1279 2417 1283 2418
rect 1303 2422 1307 2423
rect 1303 2417 1307 2418
rect 1343 2422 1347 2423
rect 1343 2417 1347 2418
rect 1375 2422 1379 2423
rect 1375 2417 1379 2418
rect 1383 2422 1387 2423
rect 1383 2417 1387 2418
rect 1415 2422 1419 2423
rect 1415 2417 1419 2418
rect 1439 2422 1443 2423
rect 1439 2417 1443 2418
rect 1455 2422 1459 2423
rect 1455 2417 1459 2418
rect 1503 2422 1507 2423
rect 1503 2417 1507 2418
rect 1511 2422 1515 2423
rect 1511 2417 1515 2418
rect 1559 2422 1563 2423
rect 1559 2417 1563 2418
rect 1583 2422 1587 2423
rect 1583 2417 1587 2418
rect 1615 2422 1619 2423
rect 1615 2417 1619 2418
rect 1663 2422 1667 2423
rect 1663 2417 1667 2418
rect 1679 2422 1683 2423
rect 1679 2417 1683 2418
rect 1239 2413 1243 2414
rect 822 2412 828 2413
rect 822 2408 823 2412
rect 827 2408 828 2412
rect 822 2407 828 2408
rect 894 2412 900 2413
rect 894 2408 895 2412
rect 899 2408 900 2412
rect 894 2407 900 2408
rect 966 2412 972 2413
rect 966 2408 967 2412
rect 971 2408 972 2412
rect 966 2407 972 2408
rect 1240 2406 1242 2413
rect 1280 2410 1282 2417
rect 1374 2416 1380 2417
rect 1374 2412 1375 2416
rect 1379 2412 1380 2416
rect 1374 2411 1380 2412
rect 1414 2416 1420 2417
rect 1414 2412 1415 2416
rect 1419 2412 1420 2416
rect 1414 2411 1420 2412
rect 1454 2416 1460 2417
rect 1454 2412 1455 2416
rect 1459 2412 1460 2416
rect 1454 2411 1460 2412
rect 1502 2416 1508 2417
rect 1502 2412 1503 2416
rect 1507 2412 1508 2416
rect 1502 2411 1508 2412
rect 1558 2416 1564 2417
rect 1558 2412 1559 2416
rect 1563 2412 1564 2416
rect 1558 2411 1564 2412
rect 1614 2416 1620 2417
rect 1614 2412 1615 2416
rect 1619 2412 1620 2416
rect 1614 2411 1620 2412
rect 1678 2416 1684 2417
rect 1678 2412 1679 2416
rect 1683 2412 1684 2416
rect 1678 2411 1684 2412
rect 1278 2409 1284 2410
rect 1238 2405 1244 2406
rect 1238 2401 1239 2405
rect 1243 2401 1244 2405
rect 1278 2405 1279 2409
rect 1283 2405 1284 2409
rect 1278 2404 1284 2405
rect 1688 2404 1690 2474
rect 1734 2471 1735 2475
rect 1739 2471 1740 2475
rect 1798 2475 1799 2479
rect 1803 2475 1804 2479
rect 1808 2476 1810 2485
rect 1878 2479 1884 2480
rect 1798 2474 1804 2475
rect 1806 2475 1812 2476
rect 1734 2470 1740 2471
rect 1800 2448 1802 2474
rect 1806 2471 1807 2475
rect 1811 2471 1812 2475
rect 1878 2475 1879 2479
rect 1883 2475 1884 2479
rect 1888 2476 1890 2485
rect 1958 2479 1964 2480
rect 1878 2474 1884 2475
rect 1886 2475 1892 2476
rect 1806 2470 1812 2471
rect 1880 2448 1882 2474
rect 1886 2471 1887 2475
rect 1891 2471 1892 2475
rect 1958 2475 1959 2479
rect 1963 2475 1964 2479
rect 1968 2476 1970 2485
rect 2064 2476 2066 2485
rect 2158 2479 2164 2480
rect 1958 2474 1964 2475
rect 1966 2475 1972 2476
rect 1886 2470 1892 2471
rect 1960 2448 1962 2474
rect 1966 2471 1967 2475
rect 1971 2471 1972 2475
rect 1966 2470 1972 2471
rect 2062 2475 2068 2476
rect 2062 2471 2063 2475
rect 2067 2471 2068 2475
rect 2158 2475 2159 2479
rect 2163 2475 2164 2479
rect 2168 2476 2170 2485
rect 2262 2479 2268 2480
rect 2158 2474 2164 2475
rect 2166 2475 2172 2476
rect 2062 2470 2068 2471
rect 2160 2448 2162 2474
rect 2166 2471 2167 2475
rect 2171 2471 2172 2475
rect 2262 2475 2263 2479
rect 2267 2475 2268 2479
rect 2272 2476 2274 2485
rect 2286 2479 2292 2480
rect 2262 2474 2268 2475
rect 2270 2475 2276 2476
rect 2166 2470 2172 2471
rect 2264 2448 2266 2474
rect 2270 2471 2271 2475
rect 2275 2471 2276 2475
rect 2286 2475 2287 2479
rect 2291 2475 2292 2479
rect 2360 2476 2362 2485
rect 2286 2474 2292 2475
rect 2358 2475 2364 2476
rect 2270 2470 2276 2471
rect 1798 2447 1804 2448
rect 1798 2443 1799 2447
rect 1803 2443 1804 2447
rect 1798 2442 1804 2443
rect 1878 2447 1884 2448
rect 1878 2443 1879 2447
rect 1883 2443 1884 2447
rect 1878 2442 1884 2443
rect 1958 2447 1964 2448
rect 1958 2443 1959 2447
rect 1963 2443 1964 2447
rect 1958 2442 1964 2443
rect 2158 2447 2164 2448
rect 2158 2443 2159 2447
rect 2163 2443 2164 2447
rect 2158 2442 2164 2443
rect 2262 2447 2268 2448
rect 2262 2443 2263 2447
rect 2267 2443 2268 2447
rect 2262 2442 2268 2443
rect 1974 2439 1980 2440
rect 1974 2435 1975 2439
rect 1979 2435 1980 2439
rect 1974 2434 1980 2435
rect 1734 2428 1740 2429
rect 1734 2424 1735 2428
rect 1739 2424 1740 2428
rect 1734 2423 1740 2424
rect 1806 2428 1812 2429
rect 1806 2424 1807 2428
rect 1811 2424 1812 2428
rect 1806 2423 1812 2424
rect 1886 2428 1892 2429
rect 1886 2424 1887 2428
rect 1891 2424 1892 2428
rect 1886 2423 1892 2424
rect 1966 2428 1972 2429
rect 1966 2424 1967 2428
rect 1971 2424 1972 2428
rect 1966 2423 1972 2424
rect 1735 2422 1739 2423
rect 1735 2417 1739 2418
rect 1799 2422 1803 2423
rect 1799 2417 1803 2418
rect 1807 2422 1811 2423
rect 1807 2417 1811 2418
rect 1871 2422 1875 2423
rect 1871 2417 1875 2418
rect 1887 2422 1891 2423
rect 1887 2417 1891 2418
rect 1951 2422 1955 2423
rect 1951 2417 1955 2418
rect 1967 2422 1971 2423
rect 1967 2417 1971 2418
rect 1734 2416 1740 2417
rect 1734 2412 1735 2416
rect 1739 2412 1740 2416
rect 1734 2411 1740 2412
rect 1798 2416 1804 2417
rect 1798 2412 1799 2416
rect 1803 2412 1804 2416
rect 1798 2411 1804 2412
rect 1870 2416 1876 2417
rect 1870 2412 1871 2416
rect 1875 2412 1876 2416
rect 1870 2411 1876 2412
rect 1950 2416 1956 2417
rect 1950 2412 1951 2416
rect 1955 2412 1956 2416
rect 1950 2411 1956 2412
rect 1238 2400 1244 2401
rect 1686 2403 1692 2404
rect 1686 2399 1687 2403
rect 1691 2399 1692 2403
rect 1686 2398 1692 2399
rect 1422 2395 1428 2396
rect 1278 2392 1284 2393
rect 838 2391 844 2392
rect 838 2387 839 2391
rect 843 2387 844 2391
rect 838 2386 844 2387
rect 906 2391 912 2392
rect 906 2387 907 2391
rect 911 2387 912 2391
rect 906 2386 912 2387
rect 1238 2388 1244 2389
rect 822 2365 828 2366
rect 822 2361 823 2365
rect 827 2361 828 2365
rect 822 2360 828 2361
rect 840 2360 842 2386
rect 894 2365 900 2366
rect 894 2361 895 2365
rect 899 2361 900 2365
rect 894 2360 900 2361
rect 472 2347 474 2360
rect 544 2347 546 2360
rect 616 2347 618 2360
rect 688 2347 690 2360
rect 734 2359 740 2360
rect 734 2355 735 2359
rect 739 2355 740 2359
rect 734 2354 740 2355
rect 471 2346 475 2347
rect 471 2341 475 2342
rect 543 2346 547 2347
rect 543 2341 547 2342
rect 551 2346 555 2347
rect 551 2341 555 2342
rect 615 2346 619 2347
rect 615 2341 619 2342
rect 631 2346 635 2347
rect 631 2341 635 2342
rect 687 2346 691 2347
rect 687 2341 691 2342
rect 711 2346 715 2347
rect 711 2341 715 2342
rect 422 2335 428 2336
rect 390 2330 396 2331
rect 398 2331 404 2332
rect 326 2326 332 2327
rect 392 2304 394 2330
rect 398 2327 399 2331
rect 403 2327 404 2331
rect 422 2331 423 2335
rect 427 2331 428 2335
rect 472 2332 474 2341
rect 482 2335 488 2336
rect 422 2330 428 2331
rect 470 2331 476 2332
rect 398 2326 404 2327
rect 470 2327 471 2331
rect 475 2327 476 2331
rect 482 2331 483 2335
rect 487 2331 488 2335
rect 552 2332 554 2341
rect 562 2335 568 2336
rect 482 2330 488 2331
rect 550 2331 556 2332
rect 470 2326 476 2327
rect 484 2312 486 2330
rect 550 2327 551 2331
rect 555 2327 556 2331
rect 562 2331 563 2335
rect 567 2331 568 2335
rect 632 2332 634 2341
rect 670 2335 676 2336
rect 562 2330 568 2331
rect 630 2331 636 2332
rect 550 2326 556 2327
rect 482 2311 488 2312
rect 482 2307 483 2311
rect 487 2307 488 2311
rect 482 2306 488 2307
rect 564 2304 566 2330
rect 630 2327 631 2331
rect 635 2327 636 2331
rect 670 2331 671 2335
rect 675 2331 676 2335
rect 712 2332 714 2341
rect 722 2335 728 2336
rect 670 2330 676 2331
rect 710 2331 716 2332
rect 630 2326 636 2327
rect 110 2303 116 2304
rect 318 2303 324 2304
rect 318 2299 319 2303
rect 323 2299 324 2303
rect 318 2298 324 2299
rect 390 2303 396 2304
rect 390 2299 391 2303
rect 395 2299 396 2303
rect 390 2298 396 2299
rect 562 2303 568 2304
rect 562 2299 563 2303
rect 567 2299 568 2303
rect 562 2298 568 2299
rect 578 2303 584 2304
rect 578 2299 579 2303
rect 583 2299 584 2303
rect 578 2298 584 2299
rect 110 2291 116 2292
rect 110 2287 111 2291
rect 115 2287 116 2291
rect 110 2286 116 2287
rect 112 2271 114 2286
rect 270 2284 276 2285
rect 270 2280 271 2284
rect 275 2280 276 2284
rect 270 2279 276 2280
rect 326 2284 332 2285
rect 326 2280 327 2284
rect 331 2280 332 2284
rect 326 2279 332 2280
rect 398 2284 404 2285
rect 398 2280 399 2284
rect 403 2280 404 2284
rect 398 2279 404 2280
rect 470 2284 476 2285
rect 470 2280 471 2284
rect 475 2280 476 2284
rect 470 2279 476 2280
rect 550 2284 556 2285
rect 550 2280 551 2284
rect 555 2280 556 2284
rect 550 2279 556 2280
rect 272 2271 274 2279
rect 328 2271 330 2279
rect 400 2271 402 2279
rect 472 2271 474 2279
rect 552 2271 554 2279
rect 111 2270 115 2271
rect 111 2265 115 2266
rect 143 2270 147 2271
rect 143 2265 147 2266
rect 183 2270 187 2271
rect 183 2265 187 2266
rect 223 2270 227 2271
rect 223 2265 227 2266
rect 271 2270 275 2271
rect 271 2265 275 2266
rect 279 2270 283 2271
rect 279 2265 283 2266
rect 327 2270 331 2271
rect 327 2265 331 2266
rect 335 2270 339 2271
rect 335 2265 339 2266
rect 399 2270 403 2271
rect 399 2265 403 2266
rect 407 2270 411 2271
rect 407 2265 411 2266
rect 471 2270 475 2271
rect 471 2265 475 2266
rect 479 2270 483 2271
rect 479 2265 483 2266
rect 551 2270 555 2271
rect 551 2265 555 2266
rect 559 2270 563 2271
rect 559 2265 563 2266
rect 112 2258 114 2265
rect 142 2264 148 2265
rect 142 2260 143 2264
rect 147 2260 148 2264
rect 142 2259 148 2260
rect 182 2264 188 2265
rect 182 2260 183 2264
rect 187 2260 188 2264
rect 182 2259 188 2260
rect 222 2264 228 2265
rect 222 2260 223 2264
rect 227 2260 228 2264
rect 222 2259 228 2260
rect 278 2264 284 2265
rect 278 2260 279 2264
rect 283 2260 284 2264
rect 278 2259 284 2260
rect 334 2264 340 2265
rect 334 2260 335 2264
rect 339 2260 340 2264
rect 334 2259 340 2260
rect 406 2264 412 2265
rect 406 2260 407 2264
rect 411 2260 412 2264
rect 406 2259 412 2260
rect 478 2264 484 2265
rect 478 2260 479 2264
rect 483 2260 484 2264
rect 478 2259 484 2260
rect 558 2264 564 2265
rect 558 2260 559 2264
rect 563 2260 564 2264
rect 558 2259 564 2260
rect 110 2257 116 2258
rect 110 2253 111 2257
rect 115 2253 116 2257
rect 110 2252 116 2253
rect 198 2243 204 2244
rect 110 2240 116 2241
rect 110 2236 111 2240
rect 115 2236 116 2240
rect 198 2239 199 2243
rect 203 2239 204 2243
rect 198 2238 204 2239
rect 238 2243 244 2244
rect 238 2239 239 2243
rect 243 2239 244 2243
rect 238 2238 244 2239
rect 294 2243 300 2244
rect 294 2239 295 2243
rect 299 2239 300 2243
rect 294 2238 300 2239
rect 350 2243 356 2244
rect 350 2239 351 2243
rect 355 2239 356 2243
rect 350 2238 356 2239
rect 378 2243 384 2244
rect 378 2239 379 2243
rect 383 2239 384 2243
rect 378 2238 384 2239
rect 386 2243 392 2244
rect 386 2239 387 2243
rect 391 2239 392 2243
rect 386 2238 392 2239
rect 542 2243 548 2244
rect 542 2239 543 2243
rect 547 2239 548 2243
rect 542 2238 548 2239
rect 550 2243 556 2244
rect 550 2239 551 2243
rect 555 2239 556 2243
rect 550 2238 556 2239
rect 110 2235 116 2236
rect 112 2203 114 2235
rect 142 2217 148 2218
rect 142 2213 143 2217
rect 147 2213 148 2217
rect 142 2212 148 2213
rect 182 2217 188 2218
rect 182 2213 183 2217
rect 187 2213 188 2217
rect 182 2212 188 2213
rect 200 2212 202 2238
rect 222 2217 228 2218
rect 222 2213 223 2217
rect 227 2213 228 2217
rect 222 2212 228 2213
rect 240 2212 242 2238
rect 278 2217 284 2218
rect 278 2213 279 2217
rect 283 2213 284 2217
rect 278 2212 284 2213
rect 296 2212 298 2238
rect 334 2217 340 2218
rect 334 2213 335 2217
rect 339 2213 340 2217
rect 334 2212 340 2213
rect 352 2212 354 2238
rect 380 2212 382 2238
rect 144 2203 146 2212
rect 162 2211 168 2212
rect 162 2207 163 2211
rect 167 2207 168 2211
rect 162 2206 168 2207
rect 111 2202 115 2203
rect 111 2197 115 2198
rect 135 2202 139 2203
rect 135 2197 139 2198
rect 143 2202 147 2203
rect 143 2197 147 2198
rect 112 2165 114 2197
rect 136 2188 138 2197
rect 134 2187 140 2188
rect 134 2183 135 2187
rect 139 2183 140 2187
rect 134 2182 140 2183
rect 110 2164 116 2165
rect 110 2160 111 2164
rect 115 2160 116 2164
rect 164 2160 166 2206
rect 184 2203 186 2212
rect 198 2211 204 2212
rect 198 2207 199 2211
rect 203 2207 204 2211
rect 198 2206 204 2207
rect 224 2203 226 2212
rect 238 2211 244 2212
rect 238 2207 239 2211
rect 243 2207 244 2211
rect 238 2206 244 2207
rect 280 2203 282 2212
rect 294 2211 300 2212
rect 294 2207 295 2211
rect 299 2207 300 2211
rect 294 2206 300 2207
rect 336 2203 338 2212
rect 350 2211 356 2212
rect 350 2207 351 2211
rect 355 2207 356 2211
rect 350 2206 356 2207
rect 378 2211 384 2212
rect 378 2207 379 2211
rect 383 2207 384 2211
rect 378 2206 384 2207
rect 183 2202 187 2203
rect 183 2197 187 2198
rect 207 2202 211 2203
rect 207 2197 211 2198
rect 223 2202 227 2203
rect 223 2197 227 2198
rect 279 2202 283 2203
rect 279 2197 283 2198
rect 335 2202 339 2203
rect 335 2197 339 2198
rect 359 2202 363 2203
rect 359 2197 363 2198
rect 198 2191 204 2192
rect 198 2187 199 2191
rect 203 2187 204 2191
rect 208 2188 210 2197
rect 280 2188 282 2197
rect 350 2191 356 2192
rect 198 2186 204 2187
rect 206 2187 212 2188
rect 200 2160 202 2186
rect 206 2183 207 2187
rect 211 2183 212 2187
rect 206 2182 212 2183
rect 278 2187 284 2188
rect 278 2183 279 2187
rect 283 2183 284 2187
rect 350 2187 351 2191
rect 355 2187 356 2191
rect 360 2188 362 2197
rect 388 2192 390 2238
rect 406 2217 412 2218
rect 406 2213 407 2217
rect 411 2213 412 2217
rect 406 2212 412 2213
rect 478 2217 484 2218
rect 478 2213 479 2217
rect 483 2213 484 2217
rect 478 2212 484 2213
rect 408 2203 410 2212
rect 480 2203 482 2212
rect 407 2202 411 2203
rect 407 2197 411 2198
rect 439 2202 443 2203
rect 439 2197 443 2198
rect 479 2202 483 2203
rect 479 2197 483 2198
rect 519 2202 523 2203
rect 519 2197 523 2198
rect 386 2191 392 2192
rect 350 2186 356 2187
rect 358 2187 364 2188
rect 278 2182 284 2183
rect 352 2160 354 2186
rect 358 2183 359 2187
rect 363 2183 364 2187
rect 386 2187 387 2191
rect 391 2187 392 2191
rect 440 2188 442 2197
rect 450 2191 456 2192
rect 386 2186 392 2187
rect 438 2187 444 2188
rect 358 2182 364 2183
rect 438 2183 439 2187
rect 443 2183 444 2187
rect 450 2187 451 2191
rect 455 2187 456 2191
rect 520 2188 522 2197
rect 544 2192 546 2238
rect 552 2212 554 2238
rect 558 2217 564 2218
rect 558 2213 559 2217
rect 563 2213 564 2217
rect 558 2212 564 2213
rect 580 2212 582 2298
rect 630 2284 636 2285
rect 630 2280 631 2284
rect 635 2280 636 2284
rect 630 2279 636 2280
rect 632 2271 634 2279
rect 631 2270 635 2271
rect 631 2265 635 2266
rect 647 2270 651 2271
rect 647 2265 651 2266
rect 646 2264 652 2265
rect 646 2260 647 2264
rect 651 2260 652 2264
rect 646 2259 652 2260
rect 672 2244 674 2330
rect 710 2327 711 2331
rect 715 2327 716 2331
rect 722 2331 723 2335
rect 727 2331 728 2335
rect 722 2330 728 2331
rect 710 2326 716 2327
rect 724 2304 726 2330
rect 736 2304 738 2354
rect 752 2347 754 2360
rect 774 2359 780 2360
rect 774 2355 775 2359
rect 779 2355 780 2359
rect 774 2354 780 2355
rect 824 2347 826 2360
rect 838 2359 844 2360
rect 838 2355 839 2359
rect 843 2355 844 2359
rect 838 2354 844 2355
rect 896 2347 898 2360
rect 751 2346 755 2347
rect 751 2341 755 2342
rect 783 2346 787 2347
rect 783 2341 787 2342
rect 823 2346 827 2347
rect 823 2341 827 2342
rect 855 2346 859 2347
rect 855 2341 859 2342
rect 895 2346 899 2347
rect 895 2341 899 2342
rect 784 2332 786 2341
rect 846 2335 852 2336
rect 782 2331 788 2332
rect 782 2327 783 2331
rect 787 2327 788 2331
rect 846 2331 847 2335
rect 851 2331 852 2335
rect 856 2332 858 2341
rect 908 2336 910 2386
rect 1238 2384 1239 2388
rect 1243 2384 1244 2388
rect 1278 2388 1279 2392
rect 1283 2388 1284 2392
rect 1422 2391 1423 2395
rect 1427 2391 1428 2395
rect 1422 2390 1428 2391
rect 1462 2395 1468 2396
rect 1462 2391 1463 2395
rect 1467 2391 1468 2395
rect 1462 2390 1468 2391
rect 1278 2387 1284 2388
rect 990 2383 996 2384
rect 1238 2383 1244 2384
rect 990 2379 991 2383
rect 995 2379 996 2383
rect 990 2378 996 2379
rect 966 2365 972 2366
rect 966 2361 967 2365
rect 971 2361 972 2365
rect 966 2360 972 2361
rect 992 2360 994 2378
rect 968 2347 970 2360
rect 990 2359 996 2360
rect 990 2355 991 2359
rect 995 2355 996 2359
rect 990 2354 996 2355
rect 1240 2347 1242 2383
rect 1280 2351 1282 2387
rect 1374 2369 1380 2370
rect 1374 2365 1375 2369
rect 1379 2365 1380 2369
rect 1374 2364 1380 2365
rect 1414 2369 1420 2370
rect 1414 2365 1415 2369
rect 1419 2365 1420 2369
rect 1414 2364 1420 2365
rect 1424 2364 1426 2390
rect 1454 2369 1460 2370
rect 1454 2365 1455 2369
rect 1459 2365 1460 2369
rect 1454 2364 1460 2365
rect 1464 2364 1466 2390
rect 1902 2387 1908 2388
rect 1902 2383 1903 2387
rect 1907 2383 1908 2387
rect 1902 2382 1908 2383
rect 1502 2369 1508 2370
rect 1502 2365 1503 2369
rect 1507 2365 1508 2369
rect 1502 2364 1508 2365
rect 1558 2369 1564 2370
rect 1558 2365 1559 2369
rect 1563 2365 1564 2369
rect 1558 2364 1564 2365
rect 1614 2369 1620 2370
rect 1614 2365 1615 2369
rect 1619 2365 1620 2369
rect 1614 2364 1620 2365
rect 1678 2369 1684 2370
rect 1678 2365 1679 2369
rect 1683 2365 1684 2369
rect 1678 2364 1684 2365
rect 1734 2369 1740 2370
rect 1734 2365 1735 2369
rect 1739 2365 1740 2369
rect 1734 2364 1740 2365
rect 1798 2369 1804 2370
rect 1798 2365 1799 2369
rect 1803 2365 1804 2369
rect 1798 2364 1804 2365
rect 1870 2369 1876 2370
rect 1870 2365 1871 2369
rect 1875 2365 1876 2369
rect 1870 2364 1876 2365
rect 1376 2351 1378 2364
rect 1416 2351 1418 2364
rect 1422 2363 1428 2364
rect 1422 2359 1423 2363
rect 1427 2359 1428 2363
rect 1422 2358 1428 2359
rect 1456 2351 1458 2364
rect 1462 2363 1468 2364
rect 1462 2359 1463 2363
rect 1467 2359 1468 2363
rect 1462 2358 1468 2359
rect 1504 2351 1506 2364
rect 1560 2351 1562 2364
rect 1616 2351 1618 2364
rect 1658 2363 1664 2364
rect 1658 2359 1659 2363
rect 1663 2359 1664 2363
rect 1658 2358 1664 2359
rect 1279 2350 1283 2351
rect 919 2346 923 2347
rect 919 2341 923 2342
rect 967 2346 971 2347
rect 967 2341 971 2342
rect 991 2346 995 2347
rect 991 2341 995 2342
rect 1063 2346 1067 2347
rect 1063 2341 1067 2342
rect 1239 2346 1243 2347
rect 1279 2345 1283 2346
rect 1327 2350 1331 2351
rect 1327 2345 1331 2346
rect 1375 2350 1379 2351
rect 1375 2345 1379 2346
rect 1383 2350 1387 2351
rect 1383 2345 1387 2346
rect 1415 2350 1419 2351
rect 1415 2345 1419 2346
rect 1439 2350 1443 2351
rect 1439 2345 1443 2346
rect 1455 2350 1459 2351
rect 1455 2345 1459 2346
rect 1503 2350 1507 2351
rect 1503 2345 1507 2346
rect 1559 2350 1563 2351
rect 1559 2345 1563 2346
rect 1575 2350 1579 2351
rect 1575 2345 1579 2346
rect 1615 2350 1619 2351
rect 1615 2345 1619 2346
rect 1647 2350 1651 2351
rect 1647 2345 1651 2346
rect 1239 2341 1243 2342
rect 906 2335 912 2336
rect 846 2330 852 2331
rect 854 2331 860 2332
rect 782 2326 788 2327
rect 848 2304 850 2330
rect 854 2327 855 2331
rect 859 2327 860 2331
rect 906 2331 907 2335
rect 911 2331 912 2335
rect 920 2332 922 2341
rect 930 2335 936 2336
rect 906 2330 912 2331
rect 918 2331 924 2332
rect 854 2326 860 2327
rect 918 2327 919 2331
rect 923 2327 924 2331
rect 930 2331 931 2335
rect 935 2331 936 2335
rect 992 2332 994 2341
rect 1054 2335 1060 2336
rect 930 2330 936 2331
rect 990 2331 996 2332
rect 918 2326 924 2327
rect 932 2312 934 2330
rect 990 2327 991 2331
rect 995 2327 996 2331
rect 1054 2331 1055 2335
rect 1059 2331 1060 2335
rect 1064 2332 1066 2341
rect 1074 2335 1080 2336
rect 1054 2330 1060 2331
rect 1062 2331 1068 2332
rect 990 2326 996 2327
rect 930 2311 936 2312
rect 930 2307 931 2311
rect 935 2307 936 2311
rect 930 2306 936 2307
rect 1056 2304 1058 2330
rect 1062 2327 1063 2331
rect 1067 2327 1068 2331
rect 1074 2331 1075 2335
rect 1079 2331 1080 2335
rect 1074 2330 1080 2331
rect 1062 2326 1068 2327
rect 1076 2312 1078 2330
rect 1074 2311 1080 2312
rect 1074 2307 1075 2311
rect 1079 2307 1080 2311
rect 1240 2309 1242 2341
rect 1280 2313 1282 2345
rect 1328 2336 1330 2345
rect 1354 2339 1360 2340
rect 1326 2335 1332 2336
rect 1326 2331 1327 2335
rect 1331 2331 1332 2335
rect 1354 2335 1355 2339
rect 1359 2335 1360 2339
rect 1384 2336 1386 2345
rect 1394 2339 1400 2340
rect 1354 2334 1360 2335
rect 1382 2335 1388 2336
rect 1326 2330 1332 2331
rect 1278 2312 1284 2313
rect 1074 2306 1080 2307
rect 1238 2308 1244 2309
rect 1238 2304 1239 2308
rect 1243 2304 1244 2308
rect 1278 2308 1279 2312
rect 1283 2308 1284 2312
rect 1278 2307 1284 2308
rect 722 2303 728 2304
rect 722 2299 723 2303
rect 727 2299 728 2303
rect 722 2298 728 2299
rect 734 2303 740 2304
rect 734 2299 735 2303
rect 739 2299 740 2303
rect 734 2298 740 2299
rect 846 2303 852 2304
rect 846 2299 847 2303
rect 851 2299 852 2303
rect 846 2298 852 2299
rect 1006 2303 1012 2304
rect 1006 2299 1007 2303
rect 1011 2299 1012 2303
rect 1006 2298 1012 2299
rect 1054 2303 1060 2304
rect 1238 2303 1244 2304
rect 1054 2299 1055 2303
rect 1059 2299 1060 2303
rect 1054 2298 1060 2299
rect 710 2284 716 2285
rect 710 2280 711 2284
rect 715 2280 716 2284
rect 710 2279 716 2280
rect 782 2284 788 2285
rect 782 2280 783 2284
rect 787 2280 788 2284
rect 782 2279 788 2280
rect 854 2284 860 2285
rect 854 2280 855 2284
rect 859 2280 860 2284
rect 854 2279 860 2280
rect 918 2284 924 2285
rect 918 2280 919 2284
rect 923 2280 924 2284
rect 918 2279 924 2280
rect 990 2284 996 2285
rect 990 2280 991 2284
rect 995 2280 996 2284
rect 990 2279 996 2280
rect 712 2271 714 2279
rect 784 2271 786 2279
rect 856 2271 858 2279
rect 920 2271 922 2279
rect 992 2271 994 2279
rect 711 2270 715 2271
rect 711 2265 715 2266
rect 727 2270 731 2271
rect 727 2265 731 2266
rect 783 2270 787 2271
rect 783 2265 787 2266
rect 807 2270 811 2271
rect 807 2265 811 2266
rect 855 2270 859 2271
rect 855 2265 859 2266
rect 887 2270 891 2271
rect 887 2265 891 2266
rect 919 2270 923 2271
rect 919 2265 923 2266
rect 967 2270 971 2271
rect 967 2265 971 2266
rect 991 2270 995 2271
rect 991 2265 995 2266
rect 726 2264 732 2265
rect 726 2260 727 2264
rect 731 2260 732 2264
rect 726 2259 732 2260
rect 806 2264 812 2265
rect 806 2260 807 2264
rect 811 2260 812 2264
rect 806 2259 812 2260
rect 886 2264 892 2265
rect 886 2260 887 2264
rect 891 2260 892 2264
rect 886 2259 892 2260
rect 966 2264 972 2265
rect 966 2260 967 2264
rect 971 2260 972 2264
rect 966 2259 972 2260
rect 670 2243 676 2244
rect 670 2239 671 2243
rect 675 2239 676 2243
rect 670 2238 676 2239
rect 686 2243 692 2244
rect 686 2239 687 2243
rect 691 2239 692 2243
rect 686 2238 692 2239
rect 646 2217 652 2218
rect 646 2213 647 2217
rect 651 2213 652 2217
rect 646 2212 652 2213
rect 688 2212 690 2238
rect 726 2217 732 2218
rect 726 2213 727 2217
rect 731 2213 732 2217
rect 726 2212 732 2213
rect 806 2217 812 2218
rect 806 2213 807 2217
rect 811 2213 812 2217
rect 806 2212 812 2213
rect 886 2217 892 2218
rect 886 2213 887 2217
rect 891 2213 892 2217
rect 886 2212 892 2213
rect 966 2217 972 2218
rect 966 2213 967 2217
rect 971 2213 972 2217
rect 1008 2216 1010 2298
rect 1278 2295 1284 2296
rect 1238 2291 1244 2292
rect 1238 2287 1239 2291
rect 1243 2287 1244 2291
rect 1278 2291 1279 2295
rect 1283 2291 1284 2295
rect 1278 2290 1284 2291
rect 1238 2286 1244 2287
rect 1062 2284 1068 2285
rect 1062 2280 1063 2284
rect 1067 2280 1068 2284
rect 1062 2279 1068 2280
rect 1064 2271 1066 2279
rect 1240 2271 1242 2286
rect 1280 2283 1282 2290
rect 1326 2288 1332 2289
rect 1326 2284 1327 2288
rect 1331 2284 1332 2288
rect 1326 2283 1332 2284
rect 1279 2282 1283 2283
rect 1279 2277 1283 2278
rect 1327 2282 1331 2283
rect 1327 2277 1331 2278
rect 1335 2282 1339 2283
rect 1335 2277 1339 2278
rect 1047 2270 1051 2271
rect 1047 2265 1051 2266
rect 1063 2270 1067 2271
rect 1063 2265 1067 2266
rect 1127 2270 1131 2271
rect 1127 2265 1131 2266
rect 1239 2270 1243 2271
rect 1280 2270 1282 2277
rect 1334 2276 1340 2277
rect 1334 2272 1335 2276
rect 1339 2272 1340 2276
rect 1334 2271 1340 2272
rect 1239 2265 1243 2266
rect 1278 2269 1284 2270
rect 1278 2265 1279 2269
rect 1283 2265 1284 2269
rect 1046 2264 1052 2265
rect 1046 2260 1047 2264
rect 1051 2260 1052 2264
rect 1046 2259 1052 2260
rect 1126 2264 1132 2265
rect 1126 2260 1127 2264
rect 1131 2260 1132 2264
rect 1126 2259 1132 2260
rect 1240 2258 1242 2265
rect 1278 2264 1284 2265
rect 1238 2257 1244 2258
rect 1238 2253 1239 2257
rect 1243 2253 1244 2257
rect 1356 2256 1358 2334
rect 1382 2331 1383 2335
rect 1387 2331 1388 2335
rect 1394 2335 1395 2339
rect 1399 2335 1400 2339
rect 1440 2336 1442 2345
rect 1450 2339 1456 2340
rect 1394 2334 1400 2335
rect 1438 2335 1444 2336
rect 1382 2330 1388 2331
rect 1396 2308 1398 2334
rect 1438 2331 1439 2335
rect 1443 2331 1444 2335
rect 1450 2335 1451 2339
rect 1455 2335 1456 2339
rect 1504 2336 1506 2345
rect 1514 2339 1520 2340
rect 1450 2334 1456 2335
rect 1502 2335 1508 2336
rect 1438 2330 1444 2331
rect 1452 2308 1454 2334
rect 1502 2331 1503 2335
rect 1507 2331 1508 2335
rect 1514 2335 1515 2339
rect 1519 2335 1520 2339
rect 1576 2336 1578 2345
rect 1586 2339 1592 2340
rect 1514 2334 1520 2335
rect 1574 2335 1580 2336
rect 1502 2330 1508 2331
rect 1516 2308 1518 2334
rect 1574 2331 1575 2335
rect 1579 2331 1580 2335
rect 1586 2335 1587 2339
rect 1591 2335 1592 2339
rect 1648 2336 1650 2345
rect 1586 2334 1592 2335
rect 1646 2335 1652 2336
rect 1574 2330 1580 2331
rect 1588 2308 1590 2334
rect 1646 2331 1647 2335
rect 1651 2331 1652 2335
rect 1646 2330 1652 2331
rect 1660 2308 1662 2358
rect 1680 2351 1682 2364
rect 1736 2351 1738 2364
rect 1800 2351 1802 2364
rect 1872 2351 1874 2364
rect 1679 2350 1683 2351
rect 1679 2345 1683 2346
rect 1719 2350 1723 2351
rect 1719 2345 1723 2346
rect 1735 2350 1739 2351
rect 1735 2345 1739 2346
rect 1799 2350 1803 2351
rect 1799 2345 1803 2346
rect 1871 2350 1875 2351
rect 1871 2345 1875 2346
rect 1879 2350 1883 2351
rect 1879 2345 1883 2346
rect 1710 2339 1716 2340
rect 1710 2335 1711 2339
rect 1715 2335 1716 2339
rect 1720 2336 1722 2345
rect 1790 2339 1796 2340
rect 1710 2334 1716 2335
rect 1718 2335 1724 2336
rect 1712 2308 1714 2334
rect 1718 2331 1719 2335
rect 1723 2331 1724 2335
rect 1790 2335 1791 2339
rect 1795 2335 1796 2339
rect 1800 2336 1802 2345
rect 1870 2339 1876 2340
rect 1790 2334 1796 2335
rect 1798 2335 1804 2336
rect 1718 2330 1724 2331
rect 1792 2308 1794 2334
rect 1798 2331 1799 2335
rect 1803 2331 1804 2335
rect 1870 2335 1871 2339
rect 1875 2335 1876 2339
rect 1880 2336 1882 2345
rect 1904 2340 1906 2382
rect 1950 2369 1956 2370
rect 1950 2365 1951 2369
rect 1955 2365 1956 2369
rect 1950 2364 1956 2365
rect 1976 2364 1978 2434
rect 2062 2428 2068 2429
rect 2062 2424 2063 2428
rect 2067 2424 2068 2428
rect 2062 2423 2068 2424
rect 2166 2428 2172 2429
rect 2166 2424 2167 2428
rect 2171 2424 2172 2428
rect 2166 2423 2172 2424
rect 2270 2428 2276 2429
rect 2270 2424 2271 2428
rect 2275 2424 2276 2428
rect 2270 2423 2276 2424
rect 2047 2422 2051 2423
rect 2047 2417 2051 2418
rect 2063 2422 2067 2423
rect 2063 2417 2067 2418
rect 2151 2422 2155 2423
rect 2151 2417 2155 2418
rect 2167 2422 2171 2423
rect 2167 2417 2171 2418
rect 2263 2422 2267 2423
rect 2263 2417 2267 2418
rect 2271 2422 2275 2423
rect 2271 2417 2275 2418
rect 2046 2416 2052 2417
rect 2046 2412 2047 2416
rect 2051 2412 2052 2416
rect 2046 2411 2052 2412
rect 2150 2416 2156 2417
rect 2150 2412 2151 2416
rect 2155 2412 2156 2416
rect 2150 2411 2156 2412
rect 2262 2416 2268 2417
rect 2262 2412 2263 2416
rect 2267 2412 2268 2416
rect 2262 2411 2268 2412
rect 2288 2396 2290 2474
rect 2358 2471 2359 2475
rect 2363 2471 2364 2475
rect 2358 2470 2364 2471
rect 2408 2453 2410 2485
rect 2406 2452 2412 2453
rect 2406 2448 2407 2452
rect 2411 2448 2412 2452
rect 2382 2447 2388 2448
rect 2406 2447 2412 2448
rect 2382 2443 2383 2447
rect 2387 2443 2388 2447
rect 2382 2442 2388 2443
rect 2358 2428 2364 2429
rect 2358 2424 2359 2428
rect 2363 2424 2364 2428
rect 2358 2423 2364 2424
rect 2359 2422 2363 2423
rect 2359 2417 2363 2418
rect 2358 2416 2364 2417
rect 2358 2412 2359 2416
rect 2363 2412 2364 2416
rect 2358 2411 2364 2412
rect 2286 2395 2292 2396
rect 2286 2391 2287 2395
rect 2291 2391 2292 2395
rect 2286 2390 2292 2391
rect 2286 2387 2292 2388
rect 2286 2383 2287 2387
rect 2291 2383 2292 2387
rect 2286 2382 2292 2383
rect 2046 2369 2052 2370
rect 2046 2365 2047 2369
rect 2051 2365 2052 2369
rect 2046 2364 2052 2365
rect 2150 2369 2156 2370
rect 2150 2365 2151 2369
rect 2155 2365 2156 2369
rect 2150 2364 2156 2365
rect 2262 2369 2268 2370
rect 2262 2365 2263 2369
rect 2267 2365 2268 2369
rect 2262 2364 2268 2365
rect 2288 2364 2290 2382
rect 2358 2369 2364 2370
rect 2358 2365 2359 2369
rect 2363 2365 2364 2369
rect 2358 2364 2364 2365
rect 2384 2364 2386 2442
rect 2406 2435 2412 2436
rect 2406 2431 2407 2435
rect 2411 2431 2412 2435
rect 2406 2430 2412 2431
rect 2408 2423 2410 2430
rect 2407 2422 2411 2423
rect 2407 2417 2411 2418
rect 2408 2410 2410 2417
rect 2406 2409 2412 2410
rect 2406 2405 2407 2409
rect 2411 2405 2412 2409
rect 2406 2404 2412 2405
rect 2406 2392 2412 2393
rect 2406 2388 2407 2392
rect 2411 2388 2412 2392
rect 2406 2387 2412 2388
rect 1952 2351 1954 2364
rect 1974 2363 1980 2364
rect 1974 2359 1975 2363
rect 1979 2359 1980 2363
rect 1974 2358 1980 2359
rect 2048 2351 2050 2364
rect 2152 2351 2154 2364
rect 2186 2363 2192 2364
rect 2186 2359 2187 2363
rect 2191 2359 2192 2363
rect 2186 2358 2192 2359
rect 1951 2350 1955 2351
rect 1951 2345 1955 2346
rect 1967 2350 1971 2351
rect 1967 2345 1971 2346
rect 2047 2350 2051 2351
rect 2047 2345 2051 2346
rect 2063 2350 2067 2351
rect 2063 2345 2067 2346
rect 2151 2350 2155 2351
rect 2151 2345 2155 2346
rect 2167 2350 2171 2351
rect 2167 2345 2171 2346
rect 1902 2339 1908 2340
rect 1870 2334 1876 2335
rect 1878 2335 1884 2336
rect 1798 2330 1804 2331
rect 1872 2308 1874 2334
rect 1878 2331 1879 2335
rect 1883 2331 1884 2335
rect 1902 2335 1903 2339
rect 1907 2335 1908 2339
rect 1968 2336 1970 2345
rect 1978 2339 1984 2340
rect 1902 2334 1908 2335
rect 1966 2335 1972 2336
rect 1878 2330 1884 2331
rect 1966 2331 1967 2335
rect 1971 2331 1972 2335
rect 1978 2335 1979 2339
rect 1983 2335 1984 2339
rect 2064 2336 2066 2345
rect 2074 2339 2080 2340
rect 1978 2334 1984 2335
rect 2062 2335 2068 2336
rect 1966 2330 1972 2331
rect 1394 2307 1400 2308
rect 1394 2303 1395 2307
rect 1399 2303 1400 2307
rect 1394 2302 1400 2303
rect 1450 2307 1456 2308
rect 1450 2303 1451 2307
rect 1455 2303 1456 2307
rect 1450 2302 1456 2303
rect 1514 2307 1520 2308
rect 1514 2303 1515 2307
rect 1519 2303 1520 2307
rect 1514 2302 1520 2303
rect 1586 2307 1592 2308
rect 1586 2303 1587 2307
rect 1591 2303 1592 2307
rect 1586 2302 1592 2303
rect 1658 2307 1664 2308
rect 1658 2303 1659 2307
rect 1663 2303 1664 2307
rect 1658 2302 1664 2303
rect 1710 2307 1716 2308
rect 1710 2303 1711 2307
rect 1715 2303 1716 2307
rect 1710 2302 1716 2303
rect 1790 2307 1796 2308
rect 1790 2303 1791 2307
rect 1795 2303 1796 2307
rect 1790 2302 1796 2303
rect 1870 2307 1876 2308
rect 1870 2303 1871 2307
rect 1875 2303 1876 2307
rect 1870 2302 1876 2303
rect 1790 2299 1796 2300
rect 1790 2295 1791 2299
rect 1795 2295 1796 2299
rect 1790 2294 1796 2295
rect 1382 2288 1388 2289
rect 1382 2284 1383 2288
rect 1387 2284 1388 2288
rect 1382 2283 1388 2284
rect 1438 2288 1444 2289
rect 1438 2284 1439 2288
rect 1443 2284 1444 2288
rect 1438 2283 1444 2284
rect 1502 2288 1508 2289
rect 1502 2284 1503 2288
rect 1507 2284 1508 2288
rect 1502 2283 1508 2284
rect 1574 2288 1580 2289
rect 1574 2284 1575 2288
rect 1579 2284 1580 2288
rect 1574 2283 1580 2284
rect 1646 2288 1652 2289
rect 1646 2284 1647 2288
rect 1651 2284 1652 2288
rect 1646 2283 1652 2284
rect 1718 2288 1724 2289
rect 1718 2284 1719 2288
rect 1723 2284 1724 2288
rect 1718 2283 1724 2284
rect 1383 2282 1387 2283
rect 1383 2277 1387 2278
rect 1407 2282 1411 2283
rect 1407 2277 1411 2278
rect 1439 2282 1443 2283
rect 1439 2277 1443 2278
rect 1487 2282 1491 2283
rect 1487 2277 1491 2278
rect 1503 2282 1507 2283
rect 1503 2277 1507 2278
rect 1559 2282 1563 2283
rect 1559 2277 1563 2278
rect 1575 2282 1579 2283
rect 1575 2277 1579 2278
rect 1631 2282 1635 2283
rect 1631 2277 1635 2278
rect 1647 2282 1651 2283
rect 1647 2277 1651 2278
rect 1703 2282 1707 2283
rect 1703 2277 1707 2278
rect 1719 2282 1723 2283
rect 1719 2277 1723 2278
rect 1775 2282 1779 2283
rect 1775 2277 1779 2278
rect 1406 2276 1412 2277
rect 1406 2272 1407 2276
rect 1411 2272 1412 2276
rect 1406 2271 1412 2272
rect 1486 2276 1492 2277
rect 1486 2272 1487 2276
rect 1491 2272 1492 2276
rect 1486 2271 1492 2272
rect 1558 2276 1564 2277
rect 1558 2272 1559 2276
rect 1563 2272 1564 2276
rect 1558 2271 1564 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1702 2276 1708 2277
rect 1702 2272 1703 2276
rect 1707 2272 1708 2276
rect 1702 2271 1708 2272
rect 1774 2276 1780 2277
rect 1774 2272 1775 2276
rect 1779 2272 1780 2276
rect 1774 2271 1780 2272
rect 1354 2255 1360 2256
rect 1238 2252 1244 2253
rect 1278 2252 1284 2253
rect 1278 2248 1279 2252
rect 1283 2248 1284 2252
rect 1354 2251 1355 2255
rect 1359 2251 1360 2255
rect 1354 2250 1360 2251
rect 1614 2255 1620 2256
rect 1614 2251 1615 2255
rect 1619 2251 1620 2255
rect 1614 2250 1620 2251
rect 1622 2255 1628 2256
rect 1622 2251 1623 2255
rect 1627 2251 1628 2255
rect 1622 2250 1628 2251
rect 1278 2247 1284 2248
rect 1134 2243 1140 2244
rect 1134 2239 1135 2243
rect 1139 2239 1140 2243
rect 1134 2238 1140 2239
rect 1142 2243 1148 2244
rect 1142 2239 1143 2243
rect 1147 2239 1148 2243
rect 1142 2238 1148 2239
rect 1238 2240 1244 2241
rect 1070 2235 1076 2236
rect 1070 2231 1071 2235
rect 1075 2231 1076 2235
rect 1070 2230 1076 2231
rect 1046 2217 1052 2218
rect 966 2212 972 2213
rect 1006 2215 1012 2216
rect 550 2211 556 2212
rect 550 2207 551 2211
rect 555 2207 556 2211
rect 550 2206 556 2207
rect 560 2203 562 2212
rect 578 2211 584 2212
rect 578 2207 579 2211
rect 583 2207 584 2211
rect 578 2206 584 2207
rect 648 2203 650 2212
rect 686 2211 692 2212
rect 686 2207 687 2211
rect 691 2207 692 2211
rect 686 2206 692 2207
rect 728 2203 730 2212
rect 808 2203 810 2212
rect 854 2211 860 2212
rect 854 2207 855 2211
rect 859 2207 860 2211
rect 854 2206 860 2207
rect 559 2202 563 2203
rect 559 2197 563 2198
rect 599 2202 603 2203
rect 599 2197 603 2198
rect 647 2202 651 2203
rect 647 2197 651 2198
rect 679 2202 683 2203
rect 679 2197 683 2198
rect 727 2202 731 2203
rect 727 2197 731 2198
rect 759 2202 763 2203
rect 759 2197 763 2198
rect 807 2202 811 2203
rect 807 2197 811 2198
rect 831 2202 835 2203
rect 831 2197 835 2198
rect 542 2191 548 2192
rect 450 2186 456 2187
rect 518 2187 524 2188
rect 438 2182 444 2183
rect 452 2168 454 2186
rect 518 2183 519 2187
rect 523 2183 524 2187
rect 542 2187 543 2191
rect 547 2187 548 2191
rect 600 2188 602 2197
rect 680 2188 682 2197
rect 746 2191 752 2192
rect 542 2186 548 2187
rect 598 2187 604 2188
rect 518 2182 524 2183
rect 598 2183 599 2187
rect 603 2183 604 2187
rect 598 2182 604 2183
rect 678 2187 684 2188
rect 678 2183 679 2187
rect 683 2183 684 2187
rect 746 2187 747 2191
rect 751 2187 752 2191
rect 760 2188 762 2197
rect 770 2191 776 2192
rect 746 2186 752 2187
rect 758 2187 764 2188
rect 678 2182 684 2183
rect 450 2167 456 2168
rect 450 2163 451 2167
rect 455 2163 456 2167
rect 450 2162 456 2163
rect 110 2159 116 2160
rect 162 2159 168 2160
rect 162 2155 163 2159
rect 167 2155 168 2159
rect 162 2154 168 2155
rect 198 2159 204 2160
rect 198 2155 199 2159
rect 203 2155 204 2159
rect 198 2154 204 2155
rect 350 2159 356 2160
rect 350 2155 351 2159
rect 355 2155 356 2159
rect 350 2154 356 2155
rect 450 2159 456 2160
rect 450 2155 451 2159
rect 455 2155 456 2159
rect 450 2154 456 2155
rect 110 2147 116 2148
rect 110 2143 111 2147
rect 115 2143 116 2147
rect 110 2142 116 2143
rect 112 2127 114 2142
rect 134 2140 140 2141
rect 134 2136 135 2140
rect 139 2136 140 2140
rect 134 2135 140 2136
rect 206 2140 212 2141
rect 206 2136 207 2140
rect 211 2136 212 2140
rect 206 2135 212 2136
rect 278 2140 284 2141
rect 278 2136 279 2140
rect 283 2136 284 2140
rect 278 2135 284 2136
rect 358 2140 364 2141
rect 358 2136 359 2140
rect 363 2136 364 2140
rect 358 2135 364 2136
rect 438 2140 444 2141
rect 438 2136 439 2140
rect 443 2136 444 2140
rect 438 2135 444 2136
rect 136 2127 138 2135
rect 208 2127 210 2135
rect 280 2127 282 2135
rect 360 2127 362 2135
rect 440 2127 442 2135
rect 111 2126 115 2127
rect 111 2121 115 2122
rect 135 2126 139 2127
rect 135 2121 139 2122
rect 191 2126 195 2127
rect 191 2121 195 2122
rect 207 2126 211 2127
rect 207 2121 211 2122
rect 271 2126 275 2127
rect 271 2121 275 2122
rect 279 2126 283 2127
rect 279 2121 283 2122
rect 343 2126 347 2127
rect 343 2121 347 2122
rect 359 2126 363 2127
rect 359 2121 363 2122
rect 415 2126 419 2127
rect 415 2121 419 2122
rect 439 2126 443 2127
rect 439 2121 443 2122
rect 112 2114 114 2121
rect 134 2120 140 2121
rect 134 2116 135 2120
rect 139 2116 140 2120
rect 134 2115 140 2116
rect 190 2120 196 2121
rect 190 2116 191 2120
rect 195 2116 196 2120
rect 190 2115 196 2116
rect 270 2120 276 2121
rect 270 2116 271 2120
rect 275 2116 276 2120
rect 270 2115 276 2116
rect 342 2120 348 2121
rect 342 2116 343 2120
rect 347 2116 348 2120
rect 342 2115 348 2116
rect 414 2120 420 2121
rect 414 2116 415 2120
rect 419 2116 420 2120
rect 414 2115 420 2116
rect 110 2113 116 2114
rect 110 2109 111 2113
rect 115 2109 116 2113
rect 110 2108 116 2109
rect 206 2099 212 2100
rect 110 2096 116 2097
rect 110 2092 111 2096
rect 115 2092 116 2096
rect 206 2095 207 2099
rect 211 2095 212 2099
rect 206 2094 212 2095
rect 110 2091 116 2092
rect 112 2055 114 2091
rect 134 2073 140 2074
rect 134 2069 135 2073
rect 139 2069 140 2073
rect 134 2068 140 2069
rect 190 2073 196 2074
rect 190 2069 191 2073
rect 195 2069 196 2073
rect 190 2068 196 2069
rect 208 2068 210 2094
rect 270 2073 276 2074
rect 270 2069 271 2073
rect 275 2069 276 2073
rect 270 2068 276 2069
rect 342 2073 348 2074
rect 342 2069 343 2073
rect 347 2069 348 2073
rect 342 2068 348 2069
rect 414 2073 420 2074
rect 414 2069 415 2073
rect 419 2069 420 2073
rect 452 2072 454 2154
rect 518 2140 524 2141
rect 518 2136 519 2140
rect 523 2136 524 2140
rect 518 2135 524 2136
rect 598 2140 604 2141
rect 598 2136 599 2140
rect 603 2136 604 2140
rect 598 2135 604 2136
rect 678 2140 684 2141
rect 678 2136 679 2140
rect 683 2136 684 2140
rect 678 2135 684 2136
rect 520 2127 522 2135
rect 600 2127 602 2135
rect 680 2127 682 2135
rect 479 2126 483 2127
rect 479 2121 483 2122
rect 519 2126 523 2127
rect 519 2121 523 2122
rect 543 2126 547 2127
rect 543 2121 547 2122
rect 599 2126 603 2127
rect 599 2121 603 2122
rect 607 2126 611 2127
rect 607 2121 611 2122
rect 671 2126 675 2127
rect 671 2121 675 2122
rect 679 2126 683 2127
rect 679 2121 683 2122
rect 735 2126 739 2127
rect 735 2121 739 2122
rect 478 2120 484 2121
rect 478 2116 479 2120
rect 483 2116 484 2120
rect 478 2115 484 2116
rect 542 2120 548 2121
rect 542 2116 543 2120
rect 547 2116 548 2120
rect 542 2115 548 2116
rect 606 2120 612 2121
rect 606 2116 607 2120
rect 611 2116 612 2120
rect 606 2115 612 2116
rect 670 2120 676 2121
rect 670 2116 671 2120
rect 675 2116 676 2120
rect 670 2115 676 2116
rect 734 2120 740 2121
rect 734 2116 735 2120
rect 739 2116 740 2120
rect 734 2115 740 2116
rect 748 2100 750 2186
rect 758 2183 759 2187
rect 763 2183 764 2187
rect 770 2187 771 2191
rect 775 2187 776 2191
rect 832 2188 834 2197
rect 842 2191 848 2192
rect 770 2186 776 2187
rect 830 2187 836 2188
rect 758 2182 764 2183
rect 772 2160 774 2186
rect 830 2183 831 2187
rect 835 2183 836 2187
rect 842 2187 843 2191
rect 847 2187 848 2191
rect 842 2186 848 2187
rect 830 2182 836 2183
rect 844 2160 846 2186
rect 856 2160 858 2206
rect 888 2203 890 2212
rect 968 2203 970 2212
rect 1006 2211 1007 2215
rect 1011 2211 1012 2215
rect 1046 2213 1047 2217
rect 1051 2213 1052 2217
rect 1046 2212 1052 2213
rect 1072 2212 1074 2230
rect 1126 2217 1132 2218
rect 1126 2213 1127 2217
rect 1131 2213 1132 2217
rect 1126 2212 1132 2213
rect 1136 2212 1138 2238
rect 1006 2210 1012 2211
rect 1048 2203 1050 2212
rect 1070 2211 1076 2212
rect 1070 2207 1071 2211
rect 1075 2207 1076 2211
rect 1070 2206 1076 2207
rect 1128 2203 1130 2212
rect 1134 2211 1140 2212
rect 1134 2207 1135 2211
rect 1139 2207 1140 2211
rect 1134 2206 1140 2207
rect 887 2202 891 2203
rect 887 2197 891 2198
rect 903 2202 907 2203
rect 903 2197 907 2198
rect 967 2202 971 2203
rect 967 2197 971 2198
rect 975 2202 979 2203
rect 975 2197 979 2198
rect 1047 2202 1051 2203
rect 1047 2197 1051 2198
rect 1119 2202 1123 2203
rect 1119 2197 1123 2198
rect 1127 2202 1131 2203
rect 1127 2197 1131 2198
rect 904 2188 906 2197
rect 966 2191 972 2192
rect 902 2187 908 2188
rect 902 2183 903 2187
rect 907 2183 908 2187
rect 966 2187 967 2191
rect 971 2187 972 2191
rect 976 2188 978 2197
rect 1038 2191 1044 2192
rect 966 2186 972 2187
rect 974 2187 980 2188
rect 902 2182 908 2183
rect 968 2160 970 2186
rect 974 2183 975 2187
rect 979 2183 980 2187
rect 1038 2187 1039 2191
rect 1043 2187 1044 2191
rect 1048 2188 1050 2197
rect 1110 2191 1116 2192
rect 1038 2186 1044 2187
rect 1046 2187 1052 2188
rect 974 2182 980 2183
rect 1040 2160 1042 2186
rect 1046 2183 1047 2187
rect 1051 2183 1052 2187
rect 1110 2187 1111 2191
rect 1115 2187 1116 2191
rect 1120 2188 1122 2197
rect 1144 2192 1146 2238
rect 1238 2236 1239 2240
rect 1243 2236 1244 2240
rect 1238 2235 1244 2236
rect 1240 2203 1242 2235
rect 1280 2207 1282 2247
rect 1334 2229 1340 2230
rect 1334 2225 1335 2229
rect 1339 2225 1340 2229
rect 1334 2224 1340 2225
rect 1406 2229 1412 2230
rect 1406 2225 1407 2229
rect 1411 2225 1412 2229
rect 1406 2224 1412 2225
rect 1486 2229 1492 2230
rect 1486 2225 1487 2229
rect 1491 2225 1492 2229
rect 1486 2224 1492 2225
rect 1558 2229 1564 2230
rect 1558 2225 1559 2229
rect 1563 2225 1564 2229
rect 1558 2224 1564 2225
rect 1336 2207 1338 2224
rect 1408 2207 1410 2224
rect 1488 2207 1490 2224
rect 1534 2223 1540 2224
rect 1534 2219 1535 2223
rect 1539 2219 1540 2223
rect 1534 2218 1540 2219
rect 1279 2206 1283 2207
rect 1239 2202 1243 2203
rect 1279 2201 1283 2202
rect 1335 2206 1339 2207
rect 1335 2201 1339 2202
rect 1375 2206 1379 2207
rect 1375 2201 1379 2202
rect 1407 2206 1411 2207
rect 1407 2201 1411 2202
rect 1439 2206 1443 2207
rect 1439 2201 1443 2202
rect 1487 2206 1491 2207
rect 1487 2201 1491 2202
rect 1511 2206 1515 2207
rect 1511 2201 1515 2202
rect 1239 2197 1243 2198
rect 1142 2191 1148 2192
rect 1110 2186 1116 2187
rect 1118 2187 1124 2188
rect 1046 2182 1052 2183
rect 1112 2160 1114 2186
rect 1118 2183 1119 2187
rect 1123 2183 1124 2187
rect 1142 2187 1143 2191
rect 1147 2187 1148 2191
rect 1142 2186 1148 2187
rect 1118 2182 1124 2183
rect 1240 2165 1242 2197
rect 1280 2169 1282 2201
rect 1376 2192 1378 2201
rect 1422 2195 1428 2196
rect 1374 2191 1380 2192
rect 1374 2187 1375 2191
rect 1379 2187 1380 2191
rect 1422 2191 1423 2195
rect 1427 2191 1428 2195
rect 1440 2192 1442 2201
rect 1450 2195 1456 2196
rect 1422 2190 1428 2191
rect 1438 2191 1444 2192
rect 1374 2186 1380 2187
rect 1278 2168 1284 2169
rect 1238 2164 1244 2165
rect 1238 2160 1239 2164
rect 1243 2160 1244 2164
rect 1278 2164 1279 2168
rect 1283 2164 1284 2168
rect 1278 2163 1284 2164
rect 770 2159 776 2160
rect 770 2155 771 2159
rect 775 2155 776 2159
rect 770 2154 776 2155
rect 842 2159 848 2160
rect 842 2155 843 2159
rect 847 2155 848 2159
rect 842 2154 848 2155
rect 854 2159 860 2160
rect 854 2155 855 2159
rect 859 2155 860 2159
rect 854 2154 860 2155
rect 966 2159 972 2160
rect 966 2155 967 2159
rect 971 2155 972 2159
rect 966 2154 972 2155
rect 1038 2159 1044 2160
rect 1038 2155 1039 2159
rect 1043 2155 1044 2159
rect 1038 2154 1044 2155
rect 1110 2159 1116 2160
rect 1238 2159 1244 2160
rect 1110 2155 1111 2159
rect 1115 2155 1116 2159
rect 1110 2154 1116 2155
rect 1070 2151 1076 2152
rect 1070 2147 1071 2151
rect 1075 2147 1076 2151
rect 1278 2151 1284 2152
rect 1070 2146 1076 2147
rect 1238 2147 1244 2148
rect 758 2140 764 2141
rect 758 2136 759 2140
rect 763 2136 764 2140
rect 758 2135 764 2136
rect 830 2140 836 2141
rect 830 2136 831 2140
rect 835 2136 836 2140
rect 830 2135 836 2136
rect 902 2140 908 2141
rect 902 2136 903 2140
rect 907 2136 908 2140
rect 902 2135 908 2136
rect 974 2140 980 2141
rect 974 2136 975 2140
rect 979 2136 980 2140
rect 974 2135 980 2136
rect 1046 2140 1052 2141
rect 1046 2136 1047 2140
rect 1051 2136 1052 2140
rect 1046 2135 1052 2136
rect 760 2127 762 2135
rect 832 2127 834 2135
rect 904 2127 906 2135
rect 976 2127 978 2135
rect 1048 2127 1050 2135
rect 759 2126 763 2127
rect 759 2121 763 2122
rect 791 2126 795 2127
rect 791 2121 795 2122
rect 831 2126 835 2127
rect 831 2121 835 2122
rect 839 2126 843 2127
rect 839 2121 843 2122
rect 887 2126 891 2127
rect 887 2121 891 2122
rect 903 2126 907 2127
rect 903 2121 907 2122
rect 935 2126 939 2127
rect 935 2121 939 2122
rect 975 2126 979 2127
rect 975 2121 979 2122
rect 991 2126 995 2127
rect 991 2121 995 2122
rect 1047 2126 1051 2127
rect 1047 2121 1051 2122
rect 790 2120 796 2121
rect 790 2116 791 2120
rect 795 2116 796 2120
rect 790 2115 796 2116
rect 838 2120 844 2121
rect 838 2116 839 2120
rect 843 2116 844 2120
rect 838 2115 844 2116
rect 886 2120 892 2121
rect 886 2116 887 2120
rect 891 2116 892 2120
rect 886 2115 892 2116
rect 934 2120 940 2121
rect 934 2116 935 2120
rect 939 2116 940 2120
rect 934 2115 940 2116
rect 990 2120 996 2121
rect 990 2116 991 2120
rect 995 2116 996 2120
rect 990 2115 996 2116
rect 1046 2120 1052 2121
rect 1046 2116 1047 2120
rect 1051 2116 1052 2120
rect 1046 2115 1052 2116
rect 506 2099 512 2100
rect 506 2095 507 2099
rect 511 2095 512 2099
rect 506 2094 512 2095
rect 622 2099 628 2100
rect 622 2095 623 2099
rect 627 2095 628 2099
rect 622 2094 628 2095
rect 686 2099 692 2100
rect 686 2095 687 2099
rect 691 2095 692 2099
rect 686 2094 692 2095
rect 698 2099 704 2100
rect 698 2095 699 2099
rect 703 2095 704 2099
rect 698 2094 704 2095
rect 746 2099 752 2100
rect 746 2095 747 2099
rect 751 2095 752 2099
rect 746 2094 752 2095
rect 498 2091 504 2092
rect 498 2087 499 2091
rect 503 2087 504 2091
rect 498 2086 504 2087
rect 478 2073 484 2074
rect 414 2068 420 2069
rect 450 2071 456 2072
rect 136 2055 138 2068
rect 158 2067 164 2068
rect 158 2063 159 2067
rect 163 2063 164 2067
rect 158 2062 164 2063
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 135 2054 139 2055
rect 135 2049 139 2050
rect 112 2017 114 2049
rect 136 2040 138 2049
rect 134 2039 140 2040
rect 134 2035 135 2039
rect 139 2035 140 2039
rect 134 2034 140 2035
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 160 2012 162 2062
rect 192 2055 194 2068
rect 206 2067 212 2068
rect 206 2063 207 2067
rect 211 2063 212 2067
rect 206 2062 212 2063
rect 272 2055 274 2068
rect 344 2055 346 2068
rect 416 2055 418 2068
rect 450 2067 451 2071
rect 455 2067 456 2071
rect 478 2069 479 2073
rect 483 2069 484 2073
rect 478 2068 484 2069
rect 500 2068 502 2086
rect 450 2066 456 2067
rect 480 2055 482 2068
rect 498 2067 504 2068
rect 498 2063 499 2067
rect 503 2063 504 2067
rect 498 2062 504 2063
rect 175 2054 179 2055
rect 175 2049 179 2050
rect 191 2054 195 2055
rect 191 2049 195 2050
rect 215 2054 219 2055
rect 215 2049 219 2050
rect 271 2054 275 2055
rect 271 2049 275 2050
rect 279 2054 283 2055
rect 279 2049 283 2050
rect 343 2054 347 2055
rect 343 2049 347 2050
rect 351 2054 355 2055
rect 351 2049 355 2050
rect 415 2054 419 2055
rect 415 2049 419 2050
rect 423 2054 427 2055
rect 423 2049 427 2050
rect 479 2054 483 2055
rect 479 2049 483 2050
rect 487 2054 491 2055
rect 487 2049 491 2050
rect 176 2040 178 2049
rect 182 2047 188 2048
rect 182 2043 183 2047
rect 187 2043 188 2047
rect 182 2042 188 2043
rect 202 2043 208 2044
rect 174 2039 180 2040
rect 174 2035 175 2039
rect 179 2035 180 2039
rect 174 2034 180 2035
rect 184 2012 186 2042
rect 202 2039 203 2043
rect 207 2039 208 2043
rect 216 2040 218 2049
rect 270 2043 276 2044
rect 202 2038 208 2039
rect 214 2039 220 2040
rect 110 2011 116 2012
rect 158 2011 164 2012
rect 158 2007 159 2011
rect 163 2007 164 2011
rect 158 2006 164 2007
rect 182 2011 188 2012
rect 182 2007 183 2011
rect 187 2007 188 2011
rect 204 2010 206 2038
rect 214 2035 215 2039
rect 219 2035 220 2039
rect 270 2039 271 2043
rect 275 2039 276 2043
rect 280 2040 282 2049
rect 342 2043 348 2044
rect 270 2038 276 2039
rect 278 2039 284 2040
rect 214 2034 220 2035
rect 272 2012 274 2038
rect 278 2035 279 2039
rect 283 2035 284 2039
rect 342 2039 343 2043
rect 347 2039 348 2043
rect 352 2040 354 2049
rect 414 2043 420 2044
rect 342 2038 348 2039
rect 350 2039 356 2040
rect 278 2034 284 2035
rect 344 2012 346 2038
rect 350 2035 351 2039
rect 355 2035 356 2039
rect 414 2039 415 2043
rect 419 2039 420 2043
rect 424 2040 426 2049
rect 434 2043 440 2044
rect 414 2038 420 2039
rect 422 2039 428 2040
rect 350 2034 356 2035
rect 416 2012 418 2038
rect 422 2035 423 2039
rect 427 2035 428 2039
rect 434 2039 435 2043
rect 439 2039 440 2043
rect 488 2040 490 2049
rect 508 2044 510 2094
rect 542 2073 548 2074
rect 542 2069 543 2073
rect 547 2069 548 2073
rect 542 2068 548 2069
rect 606 2073 612 2074
rect 606 2069 607 2073
rect 611 2069 612 2073
rect 606 2068 612 2069
rect 624 2068 626 2094
rect 670 2073 676 2074
rect 670 2069 671 2073
rect 675 2069 676 2073
rect 670 2068 676 2069
rect 688 2068 690 2094
rect 544 2055 546 2068
rect 608 2055 610 2068
rect 622 2067 628 2068
rect 622 2063 623 2067
rect 627 2063 628 2067
rect 622 2062 628 2063
rect 672 2055 674 2068
rect 686 2067 692 2068
rect 686 2063 687 2067
rect 691 2063 692 2067
rect 686 2062 692 2063
rect 543 2054 547 2055
rect 543 2049 547 2050
rect 551 2054 555 2055
rect 551 2049 555 2050
rect 607 2054 611 2055
rect 607 2049 611 2050
rect 615 2054 619 2055
rect 615 2049 619 2050
rect 671 2054 675 2055
rect 671 2049 675 2050
rect 679 2054 683 2055
rect 679 2049 683 2050
rect 506 2043 512 2044
rect 434 2038 440 2039
rect 486 2039 492 2040
rect 422 2034 428 2035
rect 210 2011 216 2012
rect 210 2010 211 2011
rect 204 2008 211 2010
rect 182 2006 188 2007
rect 210 2007 211 2008
rect 215 2007 216 2011
rect 210 2006 216 2007
rect 270 2011 276 2012
rect 270 2007 271 2011
rect 275 2007 276 2011
rect 270 2006 276 2007
rect 342 2011 348 2012
rect 342 2007 343 2011
rect 347 2007 348 2011
rect 342 2006 348 2007
rect 414 2011 420 2012
rect 414 2007 415 2011
rect 419 2007 420 2011
rect 414 2006 420 2007
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 112 1987 114 1994
rect 134 1992 140 1993
rect 134 1988 135 1992
rect 139 1988 140 1992
rect 134 1987 140 1988
rect 174 1992 180 1993
rect 174 1988 175 1992
rect 179 1988 180 1992
rect 174 1987 180 1988
rect 214 1992 220 1993
rect 214 1988 215 1992
rect 219 1988 220 1992
rect 214 1987 220 1988
rect 278 1992 284 1993
rect 278 1988 279 1992
rect 283 1988 284 1992
rect 278 1987 284 1988
rect 350 1992 356 1993
rect 350 1988 351 1992
rect 355 1988 356 1992
rect 350 1987 356 1988
rect 422 1992 428 1993
rect 422 1988 423 1992
rect 427 1988 428 1992
rect 422 1987 428 1988
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 135 1986 139 1987
rect 135 1981 139 1982
rect 175 1986 179 1987
rect 175 1981 179 1982
rect 215 1986 219 1987
rect 215 1981 219 1982
rect 271 1986 275 1987
rect 271 1981 275 1982
rect 279 1986 283 1987
rect 279 1981 283 1982
rect 343 1986 347 1987
rect 343 1981 347 1982
rect 351 1986 355 1987
rect 351 1981 355 1982
rect 415 1986 419 1987
rect 415 1981 419 1982
rect 423 1986 427 1987
rect 423 1981 427 1982
rect 112 1974 114 1981
rect 134 1980 140 1981
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 174 1980 180 1981
rect 174 1976 175 1980
rect 179 1976 180 1980
rect 174 1975 180 1976
rect 214 1980 220 1981
rect 214 1976 215 1980
rect 219 1976 220 1980
rect 214 1975 220 1976
rect 270 1980 276 1981
rect 270 1976 271 1980
rect 275 1976 276 1980
rect 270 1975 276 1976
rect 342 1980 348 1981
rect 342 1976 343 1980
rect 347 1976 348 1980
rect 342 1975 348 1976
rect 414 1980 420 1981
rect 414 1976 415 1980
rect 419 1976 420 1980
rect 414 1975 420 1976
rect 110 1973 116 1974
rect 110 1969 111 1973
rect 115 1969 116 1973
rect 110 1968 116 1969
rect 436 1968 438 2038
rect 486 2035 487 2039
rect 491 2035 492 2039
rect 506 2039 507 2043
rect 511 2039 512 2043
rect 552 2040 554 2049
rect 562 2043 568 2044
rect 506 2038 512 2039
rect 550 2039 556 2040
rect 486 2034 492 2035
rect 550 2035 551 2039
rect 555 2035 556 2039
rect 562 2039 563 2043
rect 567 2039 568 2043
rect 616 2040 618 2049
rect 680 2040 682 2049
rect 700 2044 702 2094
rect 734 2073 740 2074
rect 734 2069 735 2073
rect 739 2069 740 2073
rect 734 2068 740 2069
rect 790 2073 796 2074
rect 790 2069 791 2073
rect 795 2069 796 2073
rect 790 2068 796 2069
rect 838 2073 844 2074
rect 838 2069 839 2073
rect 843 2069 844 2073
rect 838 2068 844 2069
rect 886 2073 892 2074
rect 886 2069 887 2073
rect 891 2069 892 2073
rect 886 2068 892 2069
rect 934 2073 940 2074
rect 934 2069 935 2073
rect 939 2069 940 2073
rect 934 2068 940 2069
rect 990 2073 996 2074
rect 990 2069 991 2073
rect 995 2069 996 2073
rect 990 2068 996 2069
rect 1046 2073 1052 2074
rect 1046 2069 1047 2073
rect 1051 2069 1052 2073
rect 1046 2068 1052 2069
rect 1072 2068 1074 2146
rect 1238 2143 1239 2147
rect 1243 2143 1244 2147
rect 1278 2147 1279 2151
rect 1283 2147 1284 2151
rect 1278 2146 1284 2147
rect 1238 2142 1244 2143
rect 1118 2140 1124 2141
rect 1118 2136 1119 2140
rect 1123 2136 1124 2140
rect 1118 2135 1124 2136
rect 1120 2127 1122 2135
rect 1240 2127 1242 2142
rect 1280 2139 1282 2146
rect 1374 2144 1380 2145
rect 1374 2140 1375 2144
rect 1379 2140 1380 2144
rect 1374 2139 1380 2140
rect 1279 2138 1283 2139
rect 1279 2133 1283 2134
rect 1375 2138 1379 2139
rect 1375 2133 1379 2134
rect 1399 2138 1403 2139
rect 1399 2133 1403 2134
rect 1119 2126 1123 2127
rect 1119 2121 1123 2122
rect 1239 2126 1243 2127
rect 1280 2126 1282 2133
rect 1398 2132 1404 2133
rect 1398 2128 1399 2132
rect 1403 2128 1404 2132
rect 1398 2127 1404 2128
rect 1239 2121 1243 2122
rect 1278 2125 1284 2126
rect 1278 2121 1279 2125
rect 1283 2121 1284 2125
rect 1240 2114 1242 2121
rect 1278 2120 1284 2121
rect 1238 2113 1244 2114
rect 1238 2109 1239 2113
rect 1243 2109 1244 2113
rect 1424 2112 1426 2190
rect 1438 2187 1439 2191
rect 1443 2187 1444 2191
rect 1450 2191 1451 2195
rect 1455 2191 1456 2195
rect 1512 2192 1514 2201
rect 1522 2195 1528 2196
rect 1450 2190 1456 2191
rect 1510 2191 1516 2192
rect 1438 2186 1444 2187
rect 1452 2164 1454 2190
rect 1510 2187 1511 2191
rect 1515 2187 1516 2191
rect 1522 2191 1523 2195
rect 1527 2191 1528 2195
rect 1522 2190 1528 2191
rect 1510 2186 1516 2187
rect 1524 2164 1526 2190
rect 1536 2164 1538 2218
rect 1560 2207 1562 2224
rect 1559 2206 1563 2207
rect 1559 2201 1563 2202
rect 1591 2206 1595 2207
rect 1591 2201 1595 2202
rect 1592 2192 1594 2201
rect 1616 2196 1618 2250
rect 1624 2224 1626 2250
rect 1630 2229 1636 2230
rect 1630 2225 1631 2229
rect 1635 2225 1636 2229
rect 1630 2224 1636 2225
rect 1702 2229 1708 2230
rect 1702 2225 1703 2229
rect 1707 2225 1708 2229
rect 1702 2224 1708 2225
rect 1774 2229 1780 2230
rect 1774 2225 1775 2229
rect 1779 2225 1780 2229
rect 1774 2224 1780 2225
rect 1792 2224 1794 2294
rect 1798 2288 1804 2289
rect 1798 2284 1799 2288
rect 1803 2284 1804 2288
rect 1798 2283 1804 2284
rect 1878 2288 1884 2289
rect 1878 2284 1879 2288
rect 1883 2284 1884 2288
rect 1878 2283 1884 2284
rect 1966 2288 1972 2289
rect 1966 2284 1967 2288
rect 1971 2284 1972 2288
rect 1966 2283 1972 2284
rect 1799 2282 1803 2283
rect 1799 2277 1803 2278
rect 1839 2282 1843 2283
rect 1839 2277 1843 2278
rect 1879 2282 1883 2283
rect 1879 2277 1883 2278
rect 1911 2282 1915 2283
rect 1911 2277 1915 2278
rect 1967 2282 1971 2283
rect 1967 2277 1971 2278
rect 1838 2276 1844 2277
rect 1838 2272 1839 2276
rect 1843 2272 1844 2276
rect 1838 2271 1844 2272
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1910 2271 1916 2272
rect 1980 2264 1982 2334
rect 2062 2331 2063 2335
rect 2067 2331 2068 2335
rect 2074 2335 2075 2339
rect 2079 2335 2080 2339
rect 2168 2336 2170 2345
rect 2178 2339 2184 2340
rect 2074 2334 2080 2335
rect 2166 2335 2172 2336
rect 2062 2330 2068 2331
rect 2076 2308 2078 2334
rect 2166 2331 2167 2335
rect 2171 2331 2172 2335
rect 2178 2335 2179 2339
rect 2183 2335 2184 2339
rect 2178 2334 2184 2335
rect 2166 2330 2172 2331
rect 2180 2308 2182 2334
rect 2188 2308 2190 2358
rect 2264 2351 2266 2364
rect 2286 2363 2292 2364
rect 2286 2359 2287 2363
rect 2291 2359 2292 2363
rect 2286 2358 2292 2359
rect 2360 2351 2362 2364
rect 2382 2363 2388 2364
rect 2382 2359 2383 2363
rect 2387 2359 2388 2363
rect 2382 2358 2388 2359
rect 2408 2351 2410 2387
rect 2263 2350 2267 2351
rect 2263 2345 2267 2346
rect 2271 2350 2275 2351
rect 2271 2345 2275 2346
rect 2359 2350 2363 2351
rect 2359 2345 2363 2346
rect 2407 2350 2411 2351
rect 2407 2345 2411 2346
rect 2272 2336 2274 2345
rect 2350 2339 2356 2340
rect 2270 2335 2276 2336
rect 2270 2331 2271 2335
rect 2275 2331 2276 2335
rect 2350 2335 2351 2339
rect 2355 2335 2356 2339
rect 2360 2336 2362 2345
rect 2350 2334 2356 2335
rect 2358 2335 2364 2336
rect 2270 2330 2276 2331
rect 2352 2308 2354 2334
rect 2358 2331 2359 2335
rect 2363 2331 2364 2335
rect 2358 2330 2364 2331
rect 2408 2313 2410 2345
rect 2406 2312 2412 2313
rect 2406 2308 2407 2312
rect 2411 2308 2412 2312
rect 2074 2307 2080 2308
rect 2074 2303 2075 2307
rect 2079 2303 2080 2307
rect 2074 2302 2080 2303
rect 2178 2307 2184 2308
rect 2178 2303 2179 2307
rect 2183 2303 2184 2307
rect 2178 2302 2184 2303
rect 2186 2307 2192 2308
rect 2186 2303 2187 2307
rect 2191 2303 2192 2307
rect 2186 2302 2192 2303
rect 2342 2307 2348 2308
rect 2342 2303 2343 2307
rect 2347 2303 2348 2307
rect 2342 2302 2348 2303
rect 2350 2307 2356 2308
rect 2406 2307 2412 2308
rect 2350 2303 2351 2307
rect 2355 2303 2356 2307
rect 2350 2302 2356 2303
rect 2062 2288 2068 2289
rect 2062 2284 2063 2288
rect 2067 2284 2068 2288
rect 2062 2283 2068 2284
rect 2166 2288 2172 2289
rect 2166 2284 2167 2288
rect 2171 2284 2172 2288
rect 2166 2283 2172 2284
rect 2270 2288 2276 2289
rect 2270 2284 2271 2288
rect 2275 2284 2276 2288
rect 2270 2283 2276 2284
rect 1991 2282 1995 2283
rect 1991 2277 1995 2278
rect 2063 2282 2067 2283
rect 2063 2277 2067 2278
rect 2079 2282 2083 2283
rect 2079 2277 2083 2278
rect 2167 2282 2171 2283
rect 2167 2277 2171 2278
rect 2175 2282 2179 2283
rect 2175 2277 2179 2278
rect 2271 2282 2275 2283
rect 2271 2277 2275 2278
rect 2279 2282 2283 2283
rect 2279 2277 2283 2278
rect 1990 2276 1996 2277
rect 1990 2272 1991 2276
rect 1995 2272 1996 2276
rect 1990 2271 1996 2272
rect 2078 2276 2084 2277
rect 2078 2272 2079 2276
rect 2083 2272 2084 2276
rect 2078 2271 2084 2272
rect 2174 2276 2180 2277
rect 2174 2272 2175 2276
rect 2179 2272 2180 2276
rect 2174 2271 2180 2272
rect 2278 2276 2284 2277
rect 2278 2272 2279 2276
rect 2283 2272 2284 2276
rect 2278 2271 2284 2272
rect 1978 2263 1984 2264
rect 1978 2259 1979 2263
rect 1983 2259 1984 2263
rect 1978 2258 1984 2259
rect 1838 2229 1844 2230
rect 1838 2225 1839 2229
rect 1843 2225 1844 2229
rect 1838 2224 1844 2225
rect 1910 2229 1916 2230
rect 1910 2225 1911 2229
rect 1915 2225 1916 2229
rect 1910 2224 1916 2225
rect 1990 2229 1996 2230
rect 1990 2225 1991 2229
rect 1995 2225 1996 2229
rect 1990 2224 1996 2225
rect 2078 2229 2084 2230
rect 2078 2225 2079 2229
rect 2083 2225 2084 2229
rect 2078 2224 2084 2225
rect 2174 2229 2180 2230
rect 2174 2225 2175 2229
rect 2179 2225 2180 2229
rect 2174 2224 2180 2225
rect 2278 2229 2284 2230
rect 2278 2225 2279 2229
rect 2283 2225 2284 2229
rect 2278 2224 2284 2225
rect 2344 2224 2346 2302
rect 2406 2295 2412 2296
rect 2406 2291 2407 2295
rect 2411 2291 2412 2295
rect 2406 2290 2412 2291
rect 2358 2288 2364 2289
rect 2358 2284 2359 2288
rect 2363 2284 2364 2288
rect 2358 2283 2364 2284
rect 2408 2283 2410 2290
rect 2359 2282 2363 2283
rect 2359 2277 2363 2278
rect 2407 2282 2411 2283
rect 2407 2277 2411 2278
rect 2358 2276 2364 2277
rect 2358 2272 2359 2276
rect 2363 2272 2364 2276
rect 2358 2271 2364 2272
rect 2408 2270 2410 2277
rect 2406 2269 2412 2270
rect 2406 2265 2407 2269
rect 2411 2265 2412 2269
rect 2406 2264 2412 2265
rect 2382 2255 2388 2256
rect 2382 2251 2383 2255
rect 2387 2251 2388 2255
rect 2382 2250 2388 2251
rect 2406 2252 2412 2253
rect 2358 2229 2364 2230
rect 2358 2225 2359 2229
rect 2363 2225 2364 2229
rect 2358 2224 2364 2225
rect 1622 2223 1628 2224
rect 1622 2219 1623 2223
rect 1627 2219 1628 2223
rect 1622 2218 1628 2219
rect 1632 2207 1634 2224
rect 1704 2207 1706 2224
rect 1776 2207 1778 2224
rect 1790 2223 1796 2224
rect 1790 2219 1791 2223
rect 1795 2219 1796 2223
rect 1790 2218 1796 2219
rect 1840 2207 1842 2224
rect 1858 2215 1864 2216
rect 1858 2211 1859 2215
rect 1863 2211 1864 2215
rect 1858 2210 1864 2211
rect 1631 2206 1635 2207
rect 1631 2201 1635 2202
rect 1671 2206 1675 2207
rect 1671 2201 1675 2202
rect 1703 2206 1707 2207
rect 1703 2201 1707 2202
rect 1751 2206 1755 2207
rect 1751 2201 1755 2202
rect 1775 2206 1779 2207
rect 1775 2201 1779 2202
rect 1831 2206 1835 2207
rect 1831 2201 1835 2202
rect 1839 2206 1843 2207
rect 1839 2201 1843 2202
rect 1614 2195 1620 2196
rect 1590 2191 1596 2192
rect 1590 2187 1591 2191
rect 1595 2187 1596 2191
rect 1614 2191 1615 2195
rect 1619 2191 1620 2195
rect 1672 2192 1674 2201
rect 1682 2195 1688 2196
rect 1614 2190 1620 2191
rect 1670 2191 1676 2192
rect 1590 2186 1596 2187
rect 1670 2187 1671 2191
rect 1675 2187 1676 2191
rect 1682 2191 1683 2195
rect 1687 2191 1688 2195
rect 1752 2192 1754 2201
rect 1762 2195 1768 2196
rect 1682 2190 1688 2191
rect 1750 2191 1756 2192
rect 1670 2186 1676 2187
rect 1684 2164 1686 2190
rect 1750 2187 1751 2191
rect 1755 2187 1756 2191
rect 1762 2191 1763 2195
rect 1767 2191 1768 2195
rect 1832 2192 1834 2201
rect 1762 2190 1768 2191
rect 1830 2191 1836 2192
rect 1750 2186 1756 2187
rect 1764 2164 1766 2190
rect 1830 2187 1831 2191
rect 1835 2187 1836 2191
rect 1830 2186 1836 2187
rect 1860 2164 1862 2210
rect 1912 2207 1914 2224
rect 1992 2207 1994 2224
rect 2080 2207 2082 2224
rect 2176 2207 2178 2224
rect 2280 2207 2282 2224
rect 2342 2223 2348 2224
rect 2342 2219 2343 2223
rect 2347 2219 2348 2223
rect 2342 2218 2348 2219
rect 2360 2207 2362 2224
rect 1903 2206 1907 2207
rect 1903 2201 1907 2202
rect 1911 2206 1915 2207
rect 1911 2201 1915 2202
rect 1967 2206 1971 2207
rect 1967 2201 1971 2202
rect 1991 2206 1995 2207
rect 1991 2201 1995 2202
rect 2031 2206 2035 2207
rect 2031 2201 2035 2202
rect 2079 2206 2083 2207
rect 2079 2201 2083 2202
rect 2095 2206 2099 2207
rect 2095 2201 2099 2202
rect 2167 2206 2171 2207
rect 2167 2201 2171 2202
rect 2175 2206 2179 2207
rect 2175 2201 2179 2202
rect 2239 2206 2243 2207
rect 2239 2201 2243 2202
rect 2279 2206 2283 2207
rect 2279 2201 2283 2202
rect 2311 2206 2315 2207
rect 2311 2201 2315 2202
rect 2359 2206 2363 2207
rect 2359 2201 2363 2202
rect 1894 2195 1900 2196
rect 1894 2191 1895 2195
rect 1899 2191 1900 2195
rect 1904 2192 1906 2201
rect 1958 2195 1964 2196
rect 1894 2190 1900 2191
rect 1902 2191 1908 2192
rect 1896 2164 1898 2190
rect 1902 2187 1903 2191
rect 1907 2187 1908 2191
rect 1958 2191 1959 2195
rect 1963 2191 1964 2195
rect 1968 2192 1970 2201
rect 2022 2195 2028 2196
rect 1958 2190 1964 2191
rect 1966 2191 1972 2192
rect 1902 2186 1908 2187
rect 1960 2164 1962 2190
rect 1966 2187 1967 2191
rect 1971 2187 1972 2191
rect 2022 2191 2023 2195
rect 2027 2191 2028 2195
rect 2032 2192 2034 2201
rect 2086 2195 2092 2196
rect 2022 2190 2028 2191
rect 2030 2191 2036 2192
rect 1966 2186 1972 2187
rect 2024 2164 2026 2190
rect 2030 2187 2031 2191
rect 2035 2187 2036 2191
rect 2086 2191 2087 2195
rect 2091 2191 2092 2195
rect 2096 2192 2098 2201
rect 2158 2195 2164 2196
rect 2086 2190 2092 2191
rect 2094 2191 2100 2192
rect 2030 2186 2036 2187
rect 2088 2164 2090 2190
rect 2094 2187 2095 2191
rect 2099 2187 2100 2191
rect 2158 2191 2159 2195
rect 2163 2191 2164 2195
rect 2168 2192 2170 2201
rect 2230 2195 2236 2196
rect 2158 2190 2164 2191
rect 2166 2191 2172 2192
rect 2094 2186 2100 2187
rect 2160 2164 2162 2190
rect 2166 2187 2167 2191
rect 2171 2187 2172 2191
rect 2230 2191 2231 2195
rect 2235 2191 2236 2195
rect 2240 2192 2242 2201
rect 2250 2195 2256 2196
rect 2230 2190 2236 2191
rect 2238 2191 2244 2192
rect 2166 2186 2172 2187
rect 2232 2164 2234 2190
rect 2238 2187 2239 2191
rect 2243 2187 2244 2191
rect 2250 2191 2251 2195
rect 2255 2191 2256 2195
rect 2312 2192 2314 2201
rect 2350 2195 2356 2196
rect 2250 2190 2256 2191
rect 2310 2191 2316 2192
rect 2238 2186 2244 2187
rect 1450 2163 1456 2164
rect 1450 2159 1451 2163
rect 1455 2159 1456 2163
rect 1450 2158 1456 2159
rect 1522 2163 1528 2164
rect 1522 2159 1523 2163
rect 1527 2159 1528 2163
rect 1522 2158 1528 2159
rect 1534 2163 1540 2164
rect 1534 2159 1535 2163
rect 1539 2159 1540 2163
rect 1534 2158 1540 2159
rect 1682 2163 1688 2164
rect 1682 2159 1683 2163
rect 1687 2159 1688 2163
rect 1682 2158 1688 2159
rect 1762 2163 1768 2164
rect 1762 2159 1763 2163
rect 1767 2159 1768 2163
rect 1762 2158 1768 2159
rect 1846 2163 1852 2164
rect 1846 2159 1847 2163
rect 1851 2159 1852 2163
rect 1846 2158 1852 2159
rect 1858 2163 1864 2164
rect 1858 2159 1859 2163
rect 1863 2159 1864 2163
rect 1858 2158 1864 2159
rect 1894 2163 1900 2164
rect 1894 2159 1895 2163
rect 1899 2159 1900 2163
rect 1894 2158 1900 2159
rect 1958 2163 1964 2164
rect 1958 2159 1959 2163
rect 1963 2159 1964 2163
rect 1958 2158 1964 2159
rect 2022 2163 2028 2164
rect 2022 2159 2023 2163
rect 2027 2159 2028 2163
rect 2022 2158 2028 2159
rect 2086 2163 2092 2164
rect 2086 2159 2087 2163
rect 2091 2159 2092 2163
rect 2086 2158 2092 2159
rect 2158 2163 2164 2164
rect 2158 2159 2159 2163
rect 2163 2159 2164 2163
rect 2158 2158 2164 2159
rect 2230 2163 2236 2164
rect 2230 2159 2231 2163
rect 2235 2159 2236 2163
rect 2230 2158 2236 2159
rect 1438 2144 1444 2145
rect 1438 2140 1439 2144
rect 1443 2140 1444 2144
rect 1438 2139 1444 2140
rect 1510 2144 1516 2145
rect 1510 2140 1511 2144
rect 1515 2140 1516 2144
rect 1510 2139 1516 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1670 2144 1676 2145
rect 1670 2140 1671 2144
rect 1675 2140 1676 2144
rect 1670 2139 1676 2140
rect 1750 2144 1756 2145
rect 1750 2140 1751 2144
rect 1755 2140 1756 2144
rect 1750 2139 1756 2140
rect 1830 2144 1836 2145
rect 1830 2140 1831 2144
rect 1835 2140 1836 2144
rect 1830 2139 1836 2140
rect 1439 2138 1443 2139
rect 1439 2133 1443 2134
rect 1495 2138 1499 2139
rect 1495 2133 1499 2134
rect 1511 2138 1515 2139
rect 1511 2133 1515 2134
rect 1567 2138 1571 2139
rect 1567 2133 1571 2134
rect 1591 2138 1595 2139
rect 1591 2133 1595 2134
rect 1647 2138 1651 2139
rect 1647 2133 1651 2134
rect 1671 2138 1675 2139
rect 1671 2133 1675 2134
rect 1735 2138 1739 2139
rect 1735 2133 1739 2134
rect 1751 2138 1755 2139
rect 1751 2133 1755 2134
rect 1823 2138 1827 2139
rect 1823 2133 1827 2134
rect 1831 2138 1835 2139
rect 1831 2133 1835 2134
rect 1438 2132 1444 2133
rect 1438 2128 1439 2132
rect 1443 2128 1444 2132
rect 1438 2127 1444 2128
rect 1494 2132 1500 2133
rect 1494 2128 1495 2132
rect 1499 2128 1500 2132
rect 1494 2127 1500 2128
rect 1566 2132 1572 2133
rect 1566 2128 1567 2132
rect 1571 2128 1572 2132
rect 1566 2127 1572 2128
rect 1646 2132 1652 2133
rect 1646 2128 1647 2132
rect 1651 2128 1652 2132
rect 1646 2127 1652 2128
rect 1734 2132 1740 2133
rect 1734 2128 1735 2132
rect 1739 2128 1740 2132
rect 1734 2127 1740 2128
rect 1822 2132 1828 2133
rect 1822 2128 1823 2132
rect 1827 2128 1828 2132
rect 1822 2127 1828 2128
rect 1422 2111 1428 2112
rect 1238 2108 1244 2109
rect 1278 2108 1284 2109
rect 1278 2104 1279 2108
rect 1283 2104 1284 2108
rect 1422 2107 1423 2111
rect 1427 2107 1428 2111
rect 1422 2106 1428 2107
rect 1446 2111 1452 2112
rect 1446 2107 1447 2111
rect 1451 2107 1452 2111
rect 1446 2106 1452 2107
rect 1278 2103 1284 2104
rect 1238 2096 1244 2097
rect 1238 2092 1239 2096
rect 1243 2092 1244 2096
rect 1238 2091 1244 2092
rect 736 2055 738 2068
rect 792 2055 794 2068
rect 840 2055 842 2068
rect 888 2055 890 2068
rect 936 2055 938 2068
rect 992 2055 994 2068
rect 1048 2055 1050 2068
rect 1070 2067 1076 2068
rect 1070 2063 1071 2067
rect 1075 2063 1076 2067
rect 1070 2062 1076 2063
rect 1240 2055 1242 2091
rect 1280 2071 1282 2103
rect 1398 2085 1404 2086
rect 1398 2081 1399 2085
rect 1403 2081 1404 2085
rect 1398 2080 1404 2081
rect 1438 2085 1444 2086
rect 1438 2081 1439 2085
rect 1443 2081 1444 2085
rect 1438 2080 1444 2081
rect 1448 2080 1450 2106
rect 1494 2085 1500 2086
rect 1494 2081 1495 2085
rect 1499 2081 1500 2085
rect 1494 2080 1500 2081
rect 1566 2085 1572 2086
rect 1566 2081 1567 2085
rect 1571 2081 1572 2085
rect 1566 2080 1572 2081
rect 1646 2085 1652 2086
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1646 2080 1652 2081
rect 1734 2085 1740 2086
rect 1734 2081 1735 2085
rect 1739 2081 1740 2085
rect 1734 2080 1740 2081
rect 1822 2085 1828 2086
rect 1822 2081 1823 2085
rect 1827 2081 1828 2085
rect 1822 2080 1828 2081
rect 1848 2080 1850 2158
rect 1902 2144 1908 2145
rect 1902 2140 1903 2144
rect 1907 2140 1908 2144
rect 1902 2139 1908 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2030 2144 2036 2145
rect 2030 2140 2031 2144
rect 2035 2140 2036 2144
rect 2030 2139 2036 2140
rect 2094 2144 2100 2145
rect 2094 2140 2095 2144
rect 2099 2140 2100 2144
rect 2094 2139 2100 2140
rect 2166 2144 2172 2145
rect 2166 2140 2167 2144
rect 2171 2140 2172 2144
rect 2166 2139 2172 2140
rect 2238 2144 2244 2145
rect 2238 2140 2239 2144
rect 2243 2140 2244 2144
rect 2238 2139 2244 2140
rect 1903 2138 1907 2139
rect 1903 2133 1907 2134
rect 1911 2138 1915 2139
rect 1911 2133 1915 2134
rect 1967 2138 1971 2139
rect 1967 2133 1971 2134
rect 1999 2138 2003 2139
rect 1999 2133 2003 2134
rect 2031 2138 2035 2139
rect 2031 2133 2035 2134
rect 2087 2138 2091 2139
rect 2087 2133 2091 2134
rect 2095 2138 2099 2139
rect 2095 2133 2099 2134
rect 2167 2138 2171 2139
rect 2167 2133 2171 2134
rect 2175 2138 2179 2139
rect 2175 2133 2179 2134
rect 2239 2138 2243 2139
rect 2239 2133 2243 2134
rect 1910 2132 1916 2133
rect 1910 2128 1911 2132
rect 1915 2128 1916 2132
rect 1910 2127 1916 2128
rect 1998 2132 2004 2133
rect 1998 2128 1999 2132
rect 2003 2128 2004 2132
rect 1998 2127 2004 2128
rect 2086 2132 2092 2133
rect 2086 2128 2087 2132
rect 2091 2128 2092 2132
rect 2086 2127 2092 2128
rect 2174 2132 2180 2133
rect 2174 2128 2175 2132
rect 2179 2128 2180 2132
rect 2174 2127 2180 2128
rect 2252 2117 2254 2190
rect 2310 2187 2311 2191
rect 2315 2187 2316 2191
rect 2350 2191 2351 2195
rect 2355 2191 2356 2195
rect 2360 2192 2362 2201
rect 2384 2196 2386 2250
rect 2406 2248 2407 2252
rect 2411 2248 2412 2252
rect 2406 2247 2412 2248
rect 2408 2207 2410 2247
rect 2407 2206 2411 2207
rect 2407 2201 2411 2202
rect 2382 2195 2388 2196
rect 2350 2190 2356 2191
rect 2358 2191 2364 2192
rect 2310 2186 2316 2187
rect 2352 2164 2354 2190
rect 2358 2187 2359 2191
rect 2363 2187 2364 2191
rect 2382 2191 2383 2195
rect 2387 2191 2388 2195
rect 2382 2190 2388 2191
rect 2358 2186 2364 2187
rect 2408 2169 2410 2201
rect 2406 2168 2412 2169
rect 2406 2164 2407 2168
rect 2411 2164 2412 2168
rect 2338 2163 2344 2164
rect 2338 2159 2339 2163
rect 2343 2159 2344 2163
rect 2338 2158 2344 2159
rect 2350 2163 2356 2164
rect 2406 2163 2412 2164
rect 2350 2159 2351 2163
rect 2355 2159 2356 2163
rect 2350 2158 2356 2159
rect 2310 2144 2316 2145
rect 2310 2140 2311 2144
rect 2315 2140 2316 2144
rect 2310 2139 2316 2140
rect 2271 2138 2275 2139
rect 2271 2133 2275 2134
rect 2311 2138 2315 2139
rect 2311 2133 2315 2134
rect 2270 2132 2276 2133
rect 2270 2128 2271 2132
rect 2275 2128 2276 2132
rect 2270 2127 2276 2128
rect 1939 2116 1943 2117
rect 2251 2116 2255 2117
rect 1938 2111 1944 2112
rect 1938 2107 1939 2111
rect 1943 2107 1944 2111
rect 1938 2106 1944 2107
rect 1946 2111 1952 2112
rect 2251 2111 2255 2112
rect 1946 2107 1947 2111
rect 1951 2107 1952 2111
rect 1946 2106 1952 2107
rect 1910 2085 1916 2086
rect 1910 2081 1911 2085
rect 1915 2081 1916 2085
rect 1910 2080 1916 2081
rect 1948 2080 1950 2106
rect 1998 2085 2004 2086
rect 1998 2081 1999 2085
rect 2003 2081 2004 2085
rect 1998 2080 2004 2081
rect 2086 2085 2092 2086
rect 2086 2081 2087 2085
rect 2091 2081 2092 2085
rect 2086 2080 2092 2081
rect 2174 2085 2180 2086
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2174 2080 2180 2081
rect 2270 2085 2276 2086
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2270 2080 2276 2081
rect 2340 2080 2342 2158
rect 2406 2151 2412 2152
rect 2406 2147 2407 2151
rect 2411 2147 2412 2151
rect 2406 2146 2412 2147
rect 2358 2144 2364 2145
rect 2358 2140 2359 2144
rect 2363 2140 2364 2144
rect 2358 2139 2364 2140
rect 2408 2139 2410 2146
rect 2359 2138 2363 2139
rect 2359 2133 2363 2134
rect 2407 2138 2411 2139
rect 2407 2133 2411 2134
rect 2358 2132 2364 2133
rect 2358 2128 2359 2132
rect 2363 2128 2364 2132
rect 2358 2127 2364 2128
rect 2408 2126 2410 2133
rect 2406 2125 2412 2126
rect 2406 2121 2407 2125
rect 2411 2121 2412 2125
rect 2406 2120 2412 2121
rect 2346 2111 2352 2112
rect 2346 2107 2347 2111
rect 2351 2107 2352 2111
rect 2346 2106 2352 2107
rect 2406 2108 2412 2109
rect 1400 2071 1402 2080
rect 1440 2071 1442 2080
rect 1446 2079 1452 2080
rect 1446 2075 1447 2079
rect 1451 2075 1452 2079
rect 1446 2074 1452 2075
rect 1496 2071 1498 2080
rect 1568 2071 1570 2080
rect 1648 2071 1650 2080
rect 1736 2071 1738 2080
rect 1824 2071 1826 2080
rect 1846 2079 1852 2080
rect 1846 2075 1847 2079
rect 1851 2075 1852 2079
rect 1846 2074 1852 2075
rect 1912 2071 1914 2080
rect 1946 2079 1952 2080
rect 1946 2075 1947 2079
rect 1951 2075 1952 2079
rect 1946 2074 1952 2075
rect 2000 2071 2002 2080
rect 2088 2071 2090 2080
rect 2106 2071 2112 2072
rect 2176 2071 2178 2080
rect 2272 2071 2274 2080
rect 2338 2079 2344 2080
rect 2338 2075 2339 2079
rect 2343 2075 2344 2079
rect 2338 2074 2344 2075
rect 1279 2070 1283 2071
rect 1279 2065 1283 2066
rect 1399 2070 1403 2071
rect 1399 2065 1403 2066
rect 1439 2070 1443 2071
rect 1439 2065 1443 2066
rect 1495 2070 1499 2071
rect 1495 2065 1499 2066
rect 1567 2070 1571 2071
rect 1567 2065 1571 2066
rect 1647 2070 1651 2071
rect 1647 2065 1651 2066
rect 1735 2070 1739 2071
rect 1735 2065 1739 2066
rect 1823 2070 1827 2071
rect 1823 2065 1827 2066
rect 1911 2070 1915 2071
rect 1911 2065 1915 2066
rect 1999 2070 2003 2071
rect 1999 2065 2003 2066
rect 2039 2070 2043 2071
rect 2039 2065 2043 2066
rect 2079 2070 2083 2071
rect 2079 2065 2083 2066
rect 2087 2070 2091 2071
rect 2106 2067 2107 2071
rect 2111 2067 2112 2071
rect 2106 2066 2112 2067
rect 2119 2070 2123 2071
rect 2087 2065 2091 2066
rect 735 2054 739 2055
rect 735 2049 739 2050
rect 743 2054 747 2055
rect 743 2049 747 2050
rect 791 2054 795 2055
rect 791 2049 795 2050
rect 815 2054 819 2055
rect 815 2049 819 2050
rect 839 2054 843 2055
rect 839 2049 843 2050
rect 887 2054 891 2055
rect 887 2049 891 2050
rect 935 2054 939 2055
rect 935 2049 939 2050
rect 991 2054 995 2055
rect 991 2049 995 2050
rect 1047 2054 1051 2055
rect 1047 2049 1051 2050
rect 1239 2054 1243 2055
rect 1239 2049 1243 2050
rect 698 2043 704 2044
rect 562 2038 568 2039
rect 614 2039 620 2040
rect 550 2034 556 2035
rect 564 2012 566 2038
rect 614 2035 615 2039
rect 619 2035 620 2039
rect 614 2034 620 2035
rect 678 2039 684 2040
rect 678 2035 679 2039
rect 683 2035 684 2039
rect 698 2039 699 2043
rect 703 2039 704 2043
rect 744 2040 746 2049
rect 754 2043 760 2044
rect 698 2038 704 2039
rect 742 2039 748 2040
rect 678 2034 684 2035
rect 742 2035 743 2039
rect 747 2035 748 2039
rect 754 2039 755 2043
rect 759 2039 760 2043
rect 816 2040 818 2049
rect 826 2043 832 2044
rect 754 2038 760 2039
rect 814 2039 820 2040
rect 742 2034 748 2035
rect 756 2020 758 2038
rect 814 2035 815 2039
rect 819 2035 820 2039
rect 826 2039 827 2043
rect 831 2039 832 2043
rect 826 2038 832 2039
rect 814 2034 820 2035
rect 754 2019 760 2020
rect 828 2019 830 2038
rect 754 2015 755 2019
rect 759 2015 760 2019
rect 754 2014 760 2015
rect 824 2017 830 2019
rect 1240 2017 1242 2049
rect 1280 2033 1282 2065
rect 1942 2063 1948 2064
rect 1942 2059 1943 2063
rect 1947 2059 1948 2063
rect 1942 2058 1948 2059
rect 1278 2032 1284 2033
rect 1278 2028 1279 2032
rect 1283 2028 1284 2032
rect 1278 2027 1284 2028
rect 824 2012 826 2017
rect 1238 2016 1244 2017
rect 1238 2012 1239 2016
rect 1243 2012 1244 2016
rect 562 2011 568 2012
rect 562 2007 563 2011
rect 567 2007 568 2011
rect 562 2006 568 2007
rect 602 2011 608 2012
rect 602 2007 603 2011
rect 607 2007 608 2011
rect 602 2006 608 2007
rect 822 2011 828 2012
rect 822 2007 823 2011
rect 827 2007 828 2011
rect 822 2006 828 2007
rect 830 2011 836 2012
rect 1238 2011 1244 2012
rect 1278 2015 1284 2016
rect 1278 2011 1279 2015
rect 1283 2011 1284 2015
rect 830 2007 831 2011
rect 835 2007 836 2011
rect 1278 2010 1284 2011
rect 830 2006 836 2007
rect 486 1992 492 1993
rect 486 1988 487 1992
rect 491 1988 492 1992
rect 486 1987 492 1988
rect 550 1992 556 1993
rect 550 1988 551 1992
rect 555 1988 556 1992
rect 550 1987 556 1988
rect 487 1986 491 1987
rect 487 1981 491 1982
rect 495 1986 499 1987
rect 495 1981 499 1982
rect 551 1986 555 1987
rect 551 1981 555 1982
rect 575 1986 579 1987
rect 575 1981 579 1982
rect 494 1980 500 1981
rect 494 1976 495 1980
rect 499 1976 500 1980
rect 494 1975 500 1976
rect 574 1980 580 1981
rect 574 1976 575 1980
rect 579 1976 580 1980
rect 574 1975 580 1976
rect 434 1967 440 1968
rect 434 1963 435 1967
rect 439 1963 440 1967
rect 434 1962 440 1963
rect 182 1959 188 1960
rect 110 1956 116 1957
rect 110 1952 111 1956
rect 115 1952 116 1956
rect 182 1955 183 1959
rect 187 1955 188 1959
rect 182 1954 188 1955
rect 222 1959 228 1960
rect 222 1955 223 1959
rect 227 1955 228 1959
rect 222 1954 228 1955
rect 110 1951 116 1952
rect 112 1915 114 1951
rect 134 1933 140 1934
rect 134 1929 135 1933
rect 139 1929 140 1933
rect 134 1928 140 1929
rect 174 1933 180 1934
rect 174 1929 175 1933
rect 179 1929 180 1933
rect 174 1928 180 1929
rect 184 1928 186 1954
rect 214 1933 220 1934
rect 214 1929 215 1933
rect 219 1929 220 1933
rect 214 1928 220 1929
rect 224 1928 226 1954
rect 438 1951 444 1952
rect 438 1947 439 1951
rect 443 1947 444 1951
rect 438 1946 444 1947
rect 270 1933 276 1934
rect 270 1929 271 1933
rect 275 1929 276 1933
rect 270 1928 276 1929
rect 342 1933 348 1934
rect 342 1929 343 1933
rect 347 1929 348 1933
rect 342 1928 348 1929
rect 414 1933 420 1934
rect 414 1929 415 1933
rect 419 1929 420 1933
rect 414 1928 420 1929
rect 440 1928 442 1946
rect 494 1933 500 1934
rect 494 1929 495 1933
rect 499 1929 500 1933
rect 494 1928 500 1929
rect 574 1933 580 1934
rect 574 1929 575 1933
rect 579 1929 580 1933
rect 574 1928 580 1929
rect 604 1928 606 2006
rect 614 1992 620 1993
rect 614 1988 615 1992
rect 619 1988 620 1992
rect 614 1987 620 1988
rect 678 1992 684 1993
rect 678 1988 679 1992
rect 683 1988 684 1992
rect 678 1987 684 1988
rect 742 1992 748 1993
rect 742 1988 743 1992
rect 747 1988 748 1992
rect 742 1987 748 1988
rect 814 1992 820 1993
rect 814 1988 815 1992
rect 819 1988 820 1992
rect 814 1987 820 1988
rect 615 1986 619 1987
rect 615 1981 619 1982
rect 647 1986 651 1987
rect 647 1981 651 1982
rect 679 1986 683 1987
rect 679 1981 683 1982
rect 719 1986 723 1987
rect 719 1981 723 1982
rect 743 1986 747 1987
rect 743 1981 747 1982
rect 791 1986 795 1987
rect 791 1981 795 1982
rect 815 1986 819 1987
rect 815 1981 819 1982
rect 646 1980 652 1981
rect 646 1976 647 1980
rect 651 1976 652 1980
rect 646 1975 652 1976
rect 718 1980 724 1981
rect 718 1976 719 1980
rect 723 1976 724 1980
rect 718 1975 724 1976
rect 790 1980 796 1981
rect 790 1976 791 1980
rect 795 1976 796 1980
rect 790 1975 796 1976
rect 662 1959 668 1960
rect 662 1955 663 1959
rect 667 1955 668 1959
rect 662 1954 668 1955
rect 682 1959 688 1960
rect 682 1955 683 1959
rect 687 1955 688 1959
rect 682 1954 688 1955
rect 690 1959 696 1960
rect 690 1955 691 1959
rect 695 1955 696 1959
rect 690 1954 696 1955
rect 646 1933 652 1934
rect 646 1929 647 1933
rect 651 1929 652 1933
rect 646 1928 652 1929
rect 664 1928 666 1954
rect 684 1928 686 1954
rect 136 1915 138 1928
rect 176 1915 178 1928
rect 182 1927 188 1928
rect 182 1923 183 1927
rect 187 1923 188 1927
rect 182 1922 188 1923
rect 216 1915 218 1928
rect 222 1927 228 1928
rect 222 1923 223 1927
rect 227 1923 228 1927
rect 222 1922 228 1923
rect 272 1915 274 1928
rect 294 1919 300 1920
rect 294 1915 295 1919
rect 299 1915 300 1919
rect 344 1915 346 1928
rect 416 1915 418 1928
rect 438 1927 444 1928
rect 438 1923 439 1927
rect 443 1923 444 1927
rect 438 1922 444 1923
rect 496 1915 498 1928
rect 576 1915 578 1928
rect 602 1927 608 1928
rect 602 1923 603 1927
rect 607 1923 608 1927
rect 602 1922 608 1923
rect 648 1915 650 1928
rect 662 1927 668 1928
rect 662 1923 663 1927
rect 667 1923 668 1927
rect 662 1922 668 1923
rect 682 1927 688 1928
rect 682 1923 683 1927
rect 687 1923 688 1927
rect 682 1922 688 1923
rect 111 1914 115 1915
rect 111 1909 115 1910
rect 135 1914 139 1915
rect 135 1909 139 1910
rect 175 1914 179 1915
rect 175 1909 179 1910
rect 215 1914 219 1915
rect 215 1909 219 1910
rect 247 1914 251 1915
rect 247 1909 251 1910
rect 271 1914 275 1915
rect 271 1909 275 1910
rect 287 1914 291 1915
rect 294 1914 300 1915
rect 327 1914 331 1915
rect 287 1909 291 1910
rect 112 1877 114 1909
rect 248 1900 250 1909
rect 288 1900 290 1909
rect 246 1899 252 1900
rect 246 1895 247 1899
rect 251 1895 252 1899
rect 246 1894 252 1895
rect 286 1899 292 1900
rect 286 1895 287 1899
rect 291 1895 292 1899
rect 286 1894 292 1895
rect 110 1876 116 1877
rect 296 1876 298 1914
rect 327 1909 331 1910
rect 343 1914 347 1915
rect 343 1909 347 1910
rect 367 1914 371 1915
rect 367 1909 371 1910
rect 415 1914 419 1915
rect 415 1909 419 1910
rect 471 1914 475 1915
rect 471 1909 475 1910
rect 495 1914 499 1915
rect 495 1909 499 1910
rect 535 1914 539 1915
rect 535 1909 539 1910
rect 575 1914 579 1915
rect 575 1909 579 1910
rect 599 1914 603 1915
rect 599 1909 603 1910
rect 647 1914 651 1915
rect 647 1909 651 1910
rect 663 1914 667 1915
rect 663 1909 667 1910
rect 302 1907 308 1908
rect 302 1903 303 1907
rect 307 1903 308 1907
rect 302 1902 308 1903
rect 314 1903 320 1904
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 294 1875 300 1876
rect 294 1871 295 1875
rect 299 1871 300 1875
rect 304 1872 306 1902
rect 314 1899 315 1903
rect 319 1899 320 1903
rect 328 1900 330 1909
rect 354 1903 360 1904
rect 314 1898 320 1899
rect 326 1899 332 1900
rect 316 1880 318 1898
rect 326 1895 327 1899
rect 331 1895 332 1899
rect 354 1899 355 1903
rect 359 1899 360 1903
rect 368 1900 370 1909
rect 406 1903 412 1904
rect 354 1898 360 1899
rect 366 1899 372 1900
rect 326 1894 332 1895
rect 314 1879 320 1880
rect 314 1875 315 1879
rect 319 1875 320 1879
rect 314 1874 320 1875
rect 294 1870 300 1871
rect 302 1871 308 1872
rect 302 1867 303 1871
rect 307 1867 308 1871
rect 356 1870 358 1898
rect 366 1895 367 1899
rect 371 1895 372 1899
rect 406 1899 407 1903
rect 411 1899 412 1903
rect 416 1900 418 1909
rect 462 1903 468 1904
rect 406 1898 412 1899
rect 414 1899 420 1900
rect 366 1894 372 1895
rect 408 1872 410 1898
rect 414 1895 415 1899
rect 419 1895 420 1899
rect 462 1899 463 1903
rect 467 1899 468 1903
rect 472 1900 474 1909
rect 526 1903 532 1904
rect 462 1898 468 1899
rect 470 1899 476 1900
rect 414 1894 420 1895
rect 464 1872 466 1898
rect 470 1895 471 1899
rect 475 1895 476 1899
rect 526 1899 527 1903
rect 531 1899 532 1903
rect 536 1900 538 1909
rect 590 1903 596 1904
rect 526 1898 532 1899
rect 534 1899 540 1900
rect 470 1894 476 1895
rect 528 1872 530 1898
rect 534 1895 535 1899
rect 539 1895 540 1899
rect 590 1899 591 1903
rect 595 1899 596 1903
rect 600 1900 602 1909
rect 610 1903 616 1904
rect 590 1898 596 1899
rect 598 1899 604 1900
rect 534 1894 540 1895
rect 592 1872 594 1898
rect 598 1895 599 1899
rect 603 1895 604 1899
rect 610 1899 611 1903
rect 615 1899 616 1903
rect 664 1900 666 1909
rect 692 1904 694 1954
rect 718 1933 724 1934
rect 718 1929 719 1933
rect 723 1929 724 1933
rect 718 1928 724 1929
rect 790 1933 796 1934
rect 790 1929 791 1933
rect 795 1929 796 1933
rect 790 1928 796 1929
rect 832 1928 834 2006
rect 1280 2003 1282 2010
rect 1279 2002 1283 2003
rect 1238 1999 1244 2000
rect 1238 1995 1239 1999
rect 1243 1995 1244 1999
rect 1279 1997 1283 1998
rect 1399 2002 1403 2003
rect 1399 1997 1403 1998
rect 1439 2002 1443 2003
rect 1439 1997 1443 1998
rect 1479 2002 1483 2003
rect 1479 1997 1483 1998
rect 1519 2002 1523 2003
rect 1519 1997 1523 1998
rect 1559 2002 1563 2003
rect 1559 1997 1563 1998
rect 1599 2002 1603 2003
rect 1599 1997 1603 1998
rect 1639 2002 1643 2003
rect 1639 1997 1643 1998
rect 1679 2002 1683 2003
rect 1679 1997 1683 1998
rect 1719 2002 1723 2003
rect 1719 1997 1723 1998
rect 1767 2002 1771 2003
rect 1767 1997 1771 1998
rect 1823 2002 1827 2003
rect 1823 1997 1827 1998
rect 1871 2002 1875 2003
rect 1871 1997 1875 1998
rect 1919 2002 1923 2003
rect 1919 1997 1923 1998
rect 1238 1994 1244 1995
rect 1240 1987 1242 1994
rect 1280 1990 1282 1997
rect 1398 1996 1404 1997
rect 1398 1992 1399 1996
rect 1403 1992 1404 1996
rect 1398 1991 1404 1992
rect 1438 1996 1444 1997
rect 1438 1992 1439 1996
rect 1443 1992 1444 1996
rect 1438 1991 1444 1992
rect 1478 1996 1484 1997
rect 1478 1992 1479 1996
rect 1483 1992 1484 1996
rect 1478 1991 1484 1992
rect 1518 1996 1524 1997
rect 1518 1992 1519 1996
rect 1523 1992 1524 1996
rect 1518 1991 1524 1992
rect 1558 1996 1564 1997
rect 1558 1992 1559 1996
rect 1563 1992 1564 1996
rect 1558 1991 1564 1992
rect 1598 1996 1604 1997
rect 1598 1992 1599 1996
rect 1603 1992 1604 1996
rect 1598 1991 1604 1992
rect 1638 1996 1644 1997
rect 1638 1992 1639 1996
rect 1643 1992 1644 1996
rect 1638 1991 1644 1992
rect 1678 1996 1684 1997
rect 1678 1992 1679 1996
rect 1683 1992 1684 1996
rect 1678 1991 1684 1992
rect 1718 1996 1724 1997
rect 1718 1992 1719 1996
rect 1723 1992 1724 1996
rect 1718 1991 1724 1992
rect 1766 1996 1772 1997
rect 1766 1992 1767 1996
rect 1771 1992 1772 1996
rect 1766 1991 1772 1992
rect 1822 1996 1828 1997
rect 1822 1992 1823 1996
rect 1827 1992 1828 1996
rect 1822 1991 1828 1992
rect 1870 1996 1876 1997
rect 1870 1992 1871 1996
rect 1875 1992 1876 1996
rect 1870 1991 1876 1992
rect 1918 1996 1924 1997
rect 1918 1992 1919 1996
rect 1923 1992 1924 1996
rect 1918 1991 1924 1992
rect 1278 1989 1284 1990
rect 863 1986 867 1987
rect 863 1981 867 1982
rect 935 1986 939 1987
rect 935 1981 939 1982
rect 1007 1986 1011 1987
rect 1007 1981 1011 1982
rect 1239 1986 1243 1987
rect 1278 1985 1279 1989
rect 1283 1985 1284 1989
rect 1278 1984 1284 1985
rect 1239 1981 1243 1982
rect 862 1980 868 1981
rect 862 1976 863 1980
rect 867 1976 868 1980
rect 862 1975 868 1976
rect 934 1980 940 1981
rect 934 1976 935 1980
rect 939 1976 940 1980
rect 934 1975 940 1976
rect 1006 1980 1012 1981
rect 1006 1976 1007 1980
rect 1011 1976 1012 1980
rect 1006 1975 1012 1976
rect 1240 1974 1242 1981
rect 1944 1976 1946 2058
rect 2040 2056 2042 2065
rect 2080 2056 2082 2065
rect 2090 2059 2096 2060
rect 2038 2055 2044 2056
rect 2038 2051 2039 2055
rect 2043 2051 2044 2055
rect 2038 2050 2044 2051
rect 2078 2055 2084 2056
rect 2078 2051 2079 2055
rect 2083 2051 2084 2055
rect 2090 2055 2091 2059
rect 2095 2055 2096 2059
rect 2090 2054 2096 2055
rect 2078 2050 2084 2051
rect 2092 2028 2094 2054
rect 2108 2028 2110 2066
rect 2119 2065 2123 2066
rect 2159 2070 2163 2071
rect 2159 2065 2163 2066
rect 2175 2070 2179 2071
rect 2175 2065 2179 2066
rect 2199 2070 2203 2071
rect 2199 2065 2203 2066
rect 2239 2070 2243 2071
rect 2239 2065 2243 2066
rect 2271 2070 2275 2071
rect 2271 2065 2275 2066
rect 2279 2070 2283 2071
rect 2279 2065 2283 2066
rect 2319 2070 2323 2071
rect 2319 2065 2323 2066
rect 2120 2056 2122 2065
rect 2146 2059 2152 2060
rect 2118 2055 2124 2056
rect 2118 2051 2119 2055
rect 2123 2051 2124 2055
rect 2146 2055 2147 2059
rect 2151 2055 2152 2059
rect 2160 2056 2162 2065
rect 2200 2056 2202 2065
rect 2206 2063 2212 2064
rect 2206 2059 2207 2063
rect 2211 2059 2212 2063
rect 2206 2058 2212 2059
rect 2146 2054 2152 2055
rect 2158 2055 2164 2056
rect 2118 2050 2124 2051
rect 2148 2036 2150 2054
rect 2158 2051 2159 2055
rect 2163 2051 2164 2055
rect 2158 2050 2164 2051
rect 2198 2055 2204 2056
rect 2198 2051 2199 2055
rect 2203 2051 2204 2055
rect 2198 2050 2204 2051
rect 2146 2035 2152 2036
rect 2146 2031 2147 2035
rect 2151 2031 2152 2035
rect 2146 2030 2152 2031
rect 2208 2028 2210 2058
rect 2240 2056 2242 2065
rect 2254 2063 2260 2064
rect 2254 2059 2255 2063
rect 2259 2059 2260 2063
rect 2254 2058 2260 2059
rect 2266 2059 2272 2060
rect 2238 2055 2244 2056
rect 2238 2051 2239 2055
rect 2243 2051 2244 2055
rect 2238 2050 2244 2051
rect 2256 2028 2258 2058
rect 2266 2055 2267 2059
rect 2271 2055 2272 2059
rect 2280 2056 2282 2065
rect 2294 2059 2300 2060
rect 2266 2054 2272 2055
rect 2278 2055 2284 2056
rect 2268 2036 2270 2054
rect 2278 2051 2279 2055
rect 2283 2051 2284 2055
rect 2294 2055 2295 2059
rect 2299 2055 2300 2059
rect 2320 2056 2322 2065
rect 2348 2060 2350 2106
rect 2406 2104 2407 2108
rect 2411 2104 2412 2108
rect 2406 2103 2412 2104
rect 2358 2085 2364 2086
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2358 2080 2364 2081
rect 2360 2071 2362 2080
rect 2408 2071 2410 2103
rect 2359 2070 2363 2071
rect 2359 2065 2363 2066
rect 2407 2070 2411 2071
rect 2407 2065 2411 2066
rect 2346 2059 2352 2060
rect 2294 2054 2300 2055
rect 2318 2055 2324 2056
rect 2278 2050 2284 2051
rect 2266 2035 2272 2036
rect 2266 2031 2267 2035
rect 2271 2031 2272 2035
rect 2266 2030 2272 2031
rect 2090 2027 2096 2028
rect 2090 2023 2091 2027
rect 2095 2023 2096 2027
rect 2090 2022 2096 2023
rect 2106 2027 2112 2028
rect 2106 2023 2107 2027
rect 2111 2023 2112 2027
rect 2106 2022 2112 2023
rect 2206 2027 2212 2028
rect 2206 2023 2207 2027
rect 2211 2023 2212 2027
rect 2206 2022 2212 2023
rect 2254 2027 2260 2028
rect 2254 2023 2255 2027
rect 2259 2023 2260 2027
rect 2254 2022 2260 2023
rect 2214 2019 2220 2020
rect 2214 2015 2215 2019
rect 2219 2015 2220 2019
rect 2214 2014 2220 2015
rect 2038 2008 2044 2009
rect 2038 2004 2039 2008
rect 2043 2004 2044 2008
rect 2038 2003 2044 2004
rect 2078 2008 2084 2009
rect 2078 2004 2079 2008
rect 2083 2004 2084 2008
rect 2078 2003 2084 2004
rect 2118 2008 2124 2009
rect 2118 2004 2119 2008
rect 2123 2004 2124 2008
rect 2118 2003 2124 2004
rect 2158 2008 2164 2009
rect 2158 2004 2159 2008
rect 2163 2004 2164 2008
rect 2158 2003 2164 2004
rect 2198 2008 2204 2009
rect 2198 2004 2199 2008
rect 2203 2004 2204 2008
rect 2198 2003 2204 2004
rect 1967 2002 1971 2003
rect 1967 1997 1971 1998
rect 2015 2002 2019 2003
rect 2015 1997 2019 1998
rect 2039 2002 2043 2003
rect 2039 1997 2043 1998
rect 2055 2002 2059 2003
rect 2055 1997 2059 1998
rect 2079 2002 2083 2003
rect 2079 1997 2083 1998
rect 2095 2002 2099 2003
rect 2095 1997 2099 1998
rect 2119 2002 2123 2003
rect 2119 1997 2123 1998
rect 2143 2002 2147 2003
rect 2143 1997 2147 1998
rect 2159 2002 2163 2003
rect 2159 1997 2163 1998
rect 2191 2002 2195 2003
rect 2191 1997 2195 1998
rect 2199 2002 2203 2003
rect 2199 1997 2203 1998
rect 1966 1996 1972 1997
rect 1966 1992 1967 1996
rect 1971 1992 1972 1996
rect 1966 1991 1972 1992
rect 2014 1996 2020 1997
rect 2014 1992 2015 1996
rect 2019 1992 2020 1996
rect 2014 1991 2020 1992
rect 2054 1996 2060 1997
rect 2054 1992 2055 1996
rect 2059 1992 2060 1996
rect 2054 1991 2060 1992
rect 2094 1996 2100 1997
rect 2094 1992 2095 1996
rect 2099 1992 2100 1996
rect 2094 1991 2100 1992
rect 2142 1996 2148 1997
rect 2142 1992 2143 1996
rect 2147 1992 2148 1996
rect 2142 1991 2148 1992
rect 2190 1996 2196 1997
rect 2190 1992 2191 1996
rect 2195 1992 2196 1996
rect 2190 1991 2196 1992
rect 1446 1975 1452 1976
rect 1238 1973 1244 1974
rect 1238 1969 1239 1973
rect 1243 1969 1244 1973
rect 1238 1968 1244 1969
rect 1278 1972 1284 1973
rect 1278 1968 1279 1972
rect 1283 1968 1284 1972
rect 1446 1971 1447 1975
rect 1451 1971 1452 1975
rect 1446 1970 1452 1971
rect 1486 1975 1492 1976
rect 1486 1971 1487 1975
rect 1491 1971 1492 1975
rect 1486 1970 1492 1971
rect 1574 1975 1580 1976
rect 1574 1971 1575 1975
rect 1579 1971 1580 1975
rect 1574 1970 1580 1971
rect 1614 1975 1620 1976
rect 1614 1971 1615 1975
rect 1619 1971 1620 1975
rect 1614 1970 1620 1971
rect 1654 1975 1660 1976
rect 1654 1971 1655 1975
rect 1659 1971 1660 1975
rect 1654 1970 1660 1971
rect 1694 1975 1700 1976
rect 1694 1971 1695 1975
rect 1699 1971 1700 1975
rect 1694 1970 1700 1971
rect 1734 1975 1740 1976
rect 1734 1971 1735 1975
rect 1739 1971 1740 1975
rect 1734 1970 1740 1971
rect 1782 1975 1788 1976
rect 1782 1971 1783 1975
rect 1787 1971 1788 1975
rect 1782 1970 1788 1971
rect 1838 1975 1844 1976
rect 1838 1971 1839 1975
rect 1843 1971 1844 1975
rect 1838 1970 1844 1971
rect 1878 1975 1884 1976
rect 1878 1971 1879 1975
rect 1883 1971 1884 1975
rect 1878 1970 1884 1971
rect 1942 1975 1948 1976
rect 1942 1971 1943 1975
rect 1947 1971 1948 1975
rect 1942 1970 1948 1971
rect 2022 1975 2028 1976
rect 2022 1971 2023 1975
rect 2027 1971 2028 1975
rect 2022 1970 2028 1971
rect 2082 1975 2088 1976
rect 2082 1971 2083 1975
rect 2087 1971 2088 1975
rect 2082 1970 2088 1971
rect 2102 1975 2108 1976
rect 2102 1971 2103 1975
rect 2107 1971 2108 1975
rect 2102 1970 2108 1971
rect 1278 1967 1284 1968
rect 878 1959 884 1960
rect 878 1955 879 1959
rect 883 1955 884 1959
rect 878 1954 884 1955
rect 950 1959 956 1960
rect 950 1955 951 1959
rect 955 1955 956 1959
rect 950 1954 956 1955
rect 1014 1959 1020 1960
rect 1014 1955 1015 1959
rect 1019 1955 1020 1959
rect 1014 1954 1020 1955
rect 1022 1959 1028 1960
rect 1022 1955 1023 1959
rect 1027 1955 1028 1959
rect 1022 1954 1028 1955
rect 1238 1956 1244 1957
rect 862 1933 868 1934
rect 862 1929 863 1933
rect 867 1929 868 1933
rect 862 1928 868 1929
rect 880 1928 882 1954
rect 934 1933 940 1934
rect 934 1929 935 1933
rect 939 1929 940 1933
rect 934 1928 940 1929
rect 952 1928 954 1954
rect 1006 1933 1012 1934
rect 1006 1929 1007 1933
rect 1011 1929 1012 1933
rect 1006 1928 1012 1929
rect 1016 1928 1018 1954
rect 720 1915 722 1928
rect 792 1915 794 1928
rect 830 1927 836 1928
rect 830 1923 831 1927
rect 835 1923 836 1927
rect 830 1922 836 1923
rect 864 1915 866 1928
rect 878 1927 884 1928
rect 878 1923 879 1927
rect 883 1923 884 1927
rect 878 1922 884 1923
rect 936 1915 938 1928
rect 950 1927 956 1928
rect 950 1923 951 1927
rect 955 1923 956 1927
rect 950 1922 956 1923
rect 1008 1915 1010 1928
rect 1014 1927 1020 1928
rect 1014 1923 1015 1927
rect 1019 1923 1020 1927
rect 1014 1922 1020 1923
rect 719 1914 723 1915
rect 719 1909 723 1910
rect 727 1914 731 1915
rect 727 1909 731 1910
rect 791 1914 795 1915
rect 791 1909 795 1910
rect 855 1914 859 1915
rect 855 1909 859 1910
rect 863 1914 867 1915
rect 863 1909 867 1910
rect 919 1914 923 1915
rect 919 1909 923 1910
rect 935 1914 939 1915
rect 935 1909 939 1910
rect 983 1914 987 1915
rect 983 1909 987 1910
rect 1007 1914 1011 1915
rect 1007 1909 1011 1910
rect 690 1903 696 1904
rect 610 1898 616 1899
rect 662 1899 668 1900
rect 598 1894 604 1895
rect 362 1871 368 1872
rect 362 1870 363 1871
rect 356 1868 363 1870
rect 302 1866 308 1867
rect 362 1867 363 1868
rect 367 1867 368 1871
rect 362 1866 368 1867
rect 406 1871 412 1872
rect 406 1867 407 1871
rect 411 1867 412 1871
rect 406 1866 412 1867
rect 462 1871 468 1872
rect 462 1867 463 1871
rect 467 1867 468 1871
rect 462 1866 468 1867
rect 526 1871 532 1872
rect 526 1867 527 1871
rect 531 1867 532 1871
rect 526 1866 532 1867
rect 590 1871 596 1872
rect 590 1867 591 1871
rect 595 1867 596 1871
rect 590 1866 596 1867
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 110 1854 116 1855
rect 112 1843 114 1854
rect 246 1852 252 1853
rect 246 1848 247 1852
rect 251 1848 252 1852
rect 246 1847 252 1848
rect 286 1852 292 1853
rect 286 1848 287 1852
rect 291 1848 292 1852
rect 286 1847 292 1848
rect 326 1852 332 1853
rect 326 1848 327 1852
rect 331 1848 332 1852
rect 326 1847 332 1848
rect 366 1852 372 1853
rect 366 1848 367 1852
rect 371 1848 372 1852
rect 366 1847 372 1848
rect 414 1852 420 1853
rect 414 1848 415 1852
rect 419 1848 420 1852
rect 414 1847 420 1848
rect 470 1852 476 1853
rect 470 1848 471 1852
rect 475 1848 476 1852
rect 470 1847 476 1848
rect 534 1852 540 1853
rect 534 1848 535 1852
rect 539 1848 540 1852
rect 534 1847 540 1848
rect 598 1852 604 1853
rect 598 1848 599 1852
rect 603 1848 604 1852
rect 598 1847 604 1848
rect 248 1843 250 1847
rect 288 1843 290 1847
rect 328 1843 330 1847
rect 368 1843 370 1847
rect 416 1843 418 1847
rect 472 1843 474 1847
rect 536 1843 538 1847
rect 600 1843 602 1847
rect 111 1842 115 1843
rect 111 1837 115 1838
rect 247 1842 251 1843
rect 247 1837 251 1838
rect 287 1842 291 1843
rect 287 1837 291 1838
rect 327 1842 331 1843
rect 327 1837 331 1838
rect 367 1842 371 1843
rect 367 1837 371 1838
rect 399 1842 403 1843
rect 399 1837 403 1838
rect 415 1842 419 1843
rect 415 1837 419 1838
rect 439 1842 443 1843
rect 439 1837 443 1838
rect 471 1842 475 1843
rect 471 1837 475 1838
rect 479 1842 483 1843
rect 479 1837 483 1838
rect 519 1842 523 1843
rect 519 1837 523 1838
rect 535 1842 539 1843
rect 535 1837 539 1838
rect 567 1842 571 1843
rect 567 1837 571 1838
rect 599 1842 603 1843
rect 599 1837 603 1838
rect 112 1830 114 1837
rect 398 1836 404 1837
rect 398 1832 399 1836
rect 403 1832 404 1836
rect 398 1831 404 1832
rect 438 1836 444 1837
rect 438 1832 439 1836
rect 443 1832 444 1836
rect 438 1831 444 1832
rect 478 1836 484 1837
rect 478 1832 479 1836
rect 483 1832 484 1836
rect 478 1831 484 1832
rect 518 1836 524 1837
rect 518 1832 519 1836
rect 523 1832 524 1836
rect 518 1831 524 1832
rect 566 1836 572 1837
rect 566 1832 567 1836
rect 571 1832 572 1836
rect 566 1831 572 1832
rect 110 1829 116 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 612 1824 614 1898
rect 662 1895 663 1899
rect 667 1895 668 1899
rect 690 1899 691 1903
rect 695 1899 696 1903
rect 728 1900 730 1909
rect 738 1903 744 1904
rect 690 1898 696 1899
rect 726 1899 732 1900
rect 662 1894 668 1895
rect 726 1895 727 1899
rect 731 1895 732 1899
rect 738 1899 739 1903
rect 743 1899 744 1903
rect 792 1900 794 1909
rect 802 1903 808 1904
rect 738 1898 744 1899
rect 790 1899 796 1900
rect 726 1894 732 1895
rect 740 1872 742 1898
rect 790 1895 791 1899
rect 795 1895 796 1899
rect 802 1899 803 1903
rect 807 1899 808 1903
rect 856 1900 858 1909
rect 866 1903 872 1904
rect 866 1902 867 1903
rect 802 1898 808 1899
rect 854 1899 860 1900
rect 790 1894 796 1895
rect 804 1872 806 1898
rect 854 1895 855 1899
rect 859 1895 860 1899
rect 854 1894 860 1895
rect 864 1899 867 1902
rect 871 1899 872 1903
rect 920 1900 922 1909
rect 974 1903 980 1904
rect 864 1898 872 1899
rect 918 1899 924 1900
rect 864 1872 866 1898
rect 918 1895 919 1899
rect 923 1895 924 1899
rect 974 1899 975 1903
rect 979 1899 980 1903
rect 984 1900 986 1909
rect 1024 1908 1026 1954
rect 1238 1952 1239 1956
rect 1243 1952 1244 1956
rect 1238 1951 1244 1952
rect 1240 1915 1242 1951
rect 1280 1931 1282 1967
rect 1398 1949 1404 1950
rect 1398 1945 1399 1949
rect 1403 1945 1404 1949
rect 1398 1944 1404 1945
rect 1438 1949 1444 1950
rect 1438 1945 1439 1949
rect 1443 1945 1444 1949
rect 1438 1944 1444 1945
rect 1448 1944 1450 1970
rect 1478 1949 1484 1950
rect 1478 1945 1479 1949
rect 1483 1945 1484 1949
rect 1478 1944 1484 1945
rect 1488 1944 1490 1970
rect 1542 1967 1548 1968
rect 1542 1963 1543 1967
rect 1547 1963 1548 1967
rect 1542 1962 1548 1963
rect 1518 1949 1524 1950
rect 1518 1945 1519 1949
rect 1523 1945 1524 1949
rect 1518 1944 1524 1945
rect 1544 1944 1546 1962
rect 1558 1949 1564 1950
rect 1558 1945 1559 1949
rect 1563 1945 1564 1949
rect 1558 1944 1564 1945
rect 1576 1944 1578 1970
rect 1598 1949 1604 1950
rect 1598 1945 1599 1949
rect 1603 1945 1604 1949
rect 1598 1944 1604 1945
rect 1616 1944 1618 1970
rect 1638 1949 1644 1950
rect 1638 1945 1639 1949
rect 1643 1945 1644 1949
rect 1638 1944 1644 1945
rect 1656 1944 1658 1970
rect 1678 1949 1684 1950
rect 1678 1945 1679 1949
rect 1683 1945 1684 1949
rect 1678 1944 1684 1945
rect 1696 1944 1698 1970
rect 1718 1949 1724 1950
rect 1718 1945 1719 1949
rect 1723 1945 1724 1949
rect 1718 1944 1724 1945
rect 1736 1944 1738 1970
rect 1766 1949 1772 1950
rect 1766 1945 1767 1949
rect 1771 1945 1772 1949
rect 1766 1944 1772 1945
rect 1784 1944 1786 1970
rect 1822 1949 1828 1950
rect 1822 1945 1823 1949
rect 1827 1945 1828 1949
rect 1822 1944 1828 1945
rect 1840 1944 1842 1970
rect 1870 1949 1876 1950
rect 1870 1945 1871 1949
rect 1875 1945 1876 1949
rect 1870 1944 1876 1945
rect 1880 1944 1882 1970
rect 1918 1949 1924 1950
rect 1918 1945 1919 1949
rect 1923 1945 1924 1949
rect 1918 1944 1924 1945
rect 1966 1949 1972 1950
rect 1966 1945 1967 1949
rect 1971 1945 1972 1949
rect 1966 1944 1972 1945
rect 2014 1949 2020 1950
rect 2014 1945 2015 1949
rect 2019 1945 2020 1949
rect 2014 1944 2020 1945
rect 2024 1944 2026 1970
rect 2046 1967 2052 1968
rect 2046 1963 2047 1967
rect 2051 1963 2052 1967
rect 2046 1962 2052 1963
rect 1400 1931 1402 1944
rect 1440 1931 1442 1944
rect 1446 1943 1452 1944
rect 1446 1939 1447 1943
rect 1451 1939 1452 1943
rect 1446 1938 1452 1939
rect 1480 1931 1482 1944
rect 1486 1943 1492 1944
rect 1486 1939 1487 1943
rect 1491 1939 1492 1943
rect 1486 1938 1492 1939
rect 1520 1931 1522 1944
rect 1534 1943 1540 1944
rect 1534 1939 1535 1943
rect 1539 1939 1540 1943
rect 1534 1938 1540 1939
rect 1542 1943 1548 1944
rect 1542 1939 1543 1943
rect 1547 1939 1548 1943
rect 1542 1938 1548 1939
rect 1279 1930 1283 1931
rect 1279 1925 1283 1926
rect 1343 1930 1347 1931
rect 1343 1925 1347 1926
rect 1383 1930 1387 1931
rect 1383 1925 1387 1926
rect 1399 1930 1403 1931
rect 1399 1925 1403 1926
rect 1423 1930 1427 1931
rect 1423 1925 1427 1926
rect 1439 1930 1443 1931
rect 1439 1925 1443 1926
rect 1463 1930 1467 1931
rect 1463 1925 1467 1926
rect 1479 1930 1483 1931
rect 1479 1925 1483 1926
rect 1511 1930 1515 1931
rect 1511 1925 1515 1926
rect 1519 1930 1523 1931
rect 1519 1925 1523 1926
rect 1055 1914 1059 1915
rect 1055 1909 1059 1910
rect 1127 1914 1131 1915
rect 1127 1909 1131 1910
rect 1239 1914 1243 1915
rect 1239 1909 1243 1910
rect 1022 1907 1028 1908
rect 1022 1903 1023 1907
rect 1027 1903 1028 1907
rect 1022 1902 1028 1903
rect 1056 1900 1058 1909
rect 1118 1903 1124 1904
rect 974 1898 980 1899
rect 982 1899 988 1900
rect 918 1894 924 1895
rect 976 1872 978 1898
rect 982 1895 983 1899
rect 987 1895 988 1899
rect 982 1894 988 1895
rect 1054 1899 1060 1900
rect 1054 1895 1055 1899
rect 1059 1895 1060 1899
rect 1118 1899 1119 1903
rect 1123 1899 1124 1903
rect 1128 1900 1130 1909
rect 1138 1903 1144 1904
rect 1118 1898 1124 1899
rect 1126 1899 1132 1900
rect 1054 1894 1060 1895
rect 1120 1872 1122 1898
rect 1126 1895 1127 1899
rect 1131 1895 1132 1899
rect 1138 1899 1139 1903
rect 1143 1899 1144 1903
rect 1138 1898 1144 1899
rect 1126 1894 1132 1895
rect 1140 1880 1142 1898
rect 1138 1879 1144 1880
rect 1138 1875 1139 1879
rect 1143 1875 1144 1879
rect 1240 1877 1242 1909
rect 1280 1893 1282 1925
rect 1344 1916 1346 1925
rect 1370 1919 1376 1920
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1370 1915 1371 1919
rect 1375 1915 1376 1919
rect 1384 1916 1386 1925
rect 1394 1919 1400 1920
rect 1370 1914 1376 1915
rect 1382 1915 1388 1916
rect 1342 1910 1348 1911
rect 1278 1892 1284 1893
rect 1278 1888 1279 1892
rect 1283 1888 1284 1892
rect 1278 1887 1284 1888
rect 1138 1874 1144 1875
rect 1238 1876 1244 1877
rect 1238 1872 1239 1876
rect 1243 1872 1244 1876
rect 738 1871 744 1872
rect 738 1867 739 1871
rect 743 1867 744 1871
rect 738 1866 744 1867
rect 802 1871 808 1872
rect 802 1867 803 1871
rect 807 1867 808 1871
rect 802 1866 808 1867
rect 862 1871 868 1872
rect 862 1867 863 1871
rect 867 1867 868 1871
rect 862 1866 868 1867
rect 870 1871 876 1872
rect 870 1867 871 1871
rect 875 1867 876 1871
rect 870 1866 876 1867
rect 974 1871 980 1872
rect 974 1867 975 1871
rect 979 1867 980 1871
rect 974 1866 980 1867
rect 1070 1871 1076 1872
rect 1070 1867 1071 1871
rect 1075 1867 1076 1871
rect 1070 1866 1076 1867
rect 1118 1871 1124 1872
rect 1238 1871 1244 1872
rect 1278 1875 1284 1876
rect 1278 1871 1279 1875
rect 1283 1871 1284 1875
rect 1118 1867 1119 1871
rect 1123 1867 1124 1871
rect 1278 1870 1284 1871
rect 1118 1866 1124 1867
rect 662 1852 668 1853
rect 662 1848 663 1852
rect 667 1848 668 1852
rect 662 1847 668 1848
rect 726 1852 732 1853
rect 726 1848 727 1852
rect 731 1848 732 1852
rect 726 1847 732 1848
rect 790 1852 796 1853
rect 790 1848 791 1852
rect 795 1848 796 1852
rect 790 1847 796 1848
rect 854 1852 860 1853
rect 854 1848 855 1852
rect 859 1848 860 1852
rect 854 1847 860 1848
rect 664 1843 666 1847
rect 728 1843 730 1847
rect 792 1843 794 1847
rect 856 1843 858 1847
rect 623 1842 627 1843
rect 623 1837 627 1838
rect 663 1842 667 1843
rect 663 1837 667 1838
rect 687 1842 691 1843
rect 687 1837 691 1838
rect 727 1842 731 1843
rect 727 1837 731 1838
rect 759 1842 763 1843
rect 759 1837 763 1838
rect 791 1842 795 1843
rect 791 1837 795 1838
rect 831 1842 835 1843
rect 831 1837 835 1838
rect 855 1842 859 1843
rect 855 1837 859 1838
rect 622 1836 628 1837
rect 622 1832 623 1836
rect 627 1832 628 1836
rect 622 1831 628 1832
rect 686 1836 692 1837
rect 686 1832 687 1836
rect 691 1832 692 1836
rect 686 1831 692 1832
rect 758 1836 764 1837
rect 758 1832 759 1836
rect 763 1832 764 1836
rect 758 1831 764 1832
rect 830 1836 836 1837
rect 830 1832 831 1836
rect 835 1832 836 1836
rect 830 1831 836 1832
rect 610 1823 616 1824
rect 610 1819 611 1823
rect 615 1819 616 1823
rect 610 1818 616 1819
rect 446 1815 452 1816
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 446 1811 447 1815
rect 451 1811 452 1815
rect 446 1810 452 1811
rect 486 1815 492 1816
rect 486 1811 487 1815
rect 491 1811 492 1815
rect 486 1810 492 1811
rect 526 1815 532 1816
rect 526 1811 527 1815
rect 531 1811 532 1815
rect 526 1810 532 1811
rect 110 1807 116 1808
rect 112 1775 114 1807
rect 398 1789 404 1790
rect 398 1785 399 1789
rect 403 1785 404 1789
rect 398 1784 404 1785
rect 438 1789 444 1790
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 438 1784 444 1785
rect 448 1784 450 1810
rect 478 1789 484 1790
rect 478 1785 479 1789
rect 483 1785 484 1789
rect 478 1784 484 1785
rect 488 1784 490 1810
rect 518 1789 524 1790
rect 518 1785 519 1789
rect 523 1785 524 1789
rect 518 1784 524 1785
rect 528 1784 530 1810
rect 566 1789 572 1790
rect 566 1785 567 1789
rect 571 1785 572 1789
rect 566 1784 572 1785
rect 622 1789 628 1790
rect 622 1785 623 1789
rect 627 1785 628 1789
rect 622 1784 628 1785
rect 686 1789 692 1790
rect 686 1785 687 1789
rect 691 1785 692 1789
rect 686 1784 692 1785
rect 758 1789 764 1790
rect 758 1785 759 1789
rect 763 1785 764 1789
rect 758 1784 764 1785
rect 830 1789 836 1790
rect 830 1785 831 1789
rect 835 1785 836 1789
rect 872 1788 874 1866
rect 918 1852 924 1853
rect 918 1848 919 1852
rect 923 1848 924 1852
rect 918 1847 924 1848
rect 982 1852 988 1853
rect 982 1848 983 1852
rect 987 1848 988 1852
rect 982 1847 988 1848
rect 1054 1852 1060 1853
rect 1054 1848 1055 1852
rect 1059 1848 1060 1852
rect 1054 1847 1060 1848
rect 920 1843 922 1847
rect 984 1843 986 1847
rect 1056 1843 1058 1847
rect 903 1842 907 1843
rect 903 1837 907 1838
rect 919 1842 923 1843
rect 919 1837 923 1838
rect 975 1842 979 1843
rect 975 1837 979 1838
rect 983 1842 987 1843
rect 983 1837 987 1838
rect 1047 1842 1051 1843
rect 1047 1837 1051 1838
rect 1055 1842 1059 1843
rect 1055 1837 1059 1838
rect 902 1836 908 1837
rect 902 1832 903 1836
rect 907 1832 908 1836
rect 902 1831 908 1832
rect 974 1836 980 1837
rect 974 1832 975 1836
rect 979 1832 980 1836
rect 974 1831 980 1832
rect 1046 1836 1052 1837
rect 1046 1832 1047 1836
rect 1051 1832 1052 1836
rect 1046 1831 1052 1832
rect 958 1815 964 1816
rect 958 1811 959 1815
rect 963 1811 964 1815
rect 958 1810 964 1811
rect 926 1807 932 1808
rect 926 1803 927 1807
rect 931 1803 932 1807
rect 926 1802 932 1803
rect 902 1789 908 1790
rect 830 1784 836 1785
rect 870 1787 876 1788
rect 400 1775 402 1784
rect 440 1775 442 1784
rect 446 1783 452 1784
rect 446 1779 447 1783
rect 451 1779 452 1783
rect 446 1778 452 1779
rect 480 1775 482 1784
rect 486 1783 492 1784
rect 486 1779 487 1783
rect 491 1779 492 1783
rect 486 1778 492 1779
rect 520 1775 522 1784
rect 526 1783 532 1784
rect 526 1779 527 1783
rect 531 1779 532 1783
rect 526 1778 532 1779
rect 568 1775 570 1784
rect 624 1775 626 1784
rect 674 1783 680 1784
rect 674 1779 675 1783
rect 679 1779 680 1783
rect 674 1778 680 1779
rect 111 1774 115 1775
rect 111 1769 115 1770
rect 399 1774 403 1775
rect 399 1769 403 1770
rect 407 1774 411 1775
rect 407 1769 411 1770
rect 439 1774 443 1775
rect 439 1769 443 1770
rect 447 1774 451 1775
rect 447 1769 451 1770
rect 479 1774 483 1775
rect 479 1769 483 1770
rect 487 1774 491 1775
rect 487 1769 491 1770
rect 519 1774 523 1775
rect 519 1769 523 1770
rect 527 1774 531 1775
rect 527 1769 531 1770
rect 567 1774 571 1775
rect 567 1769 571 1770
rect 607 1774 611 1775
rect 607 1769 611 1770
rect 623 1774 627 1775
rect 623 1769 627 1770
rect 647 1774 651 1775
rect 647 1769 651 1770
rect 112 1737 114 1769
rect 408 1760 410 1769
rect 434 1763 440 1764
rect 406 1759 412 1760
rect 406 1755 407 1759
rect 411 1755 412 1759
rect 434 1759 435 1763
rect 439 1759 440 1763
rect 448 1760 450 1769
rect 458 1763 464 1764
rect 434 1758 440 1759
rect 446 1759 452 1760
rect 406 1754 412 1755
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 110 1714 116 1715
rect 112 1703 114 1714
rect 406 1712 412 1713
rect 406 1708 407 1712
rect 411 1708 412 1712
rect 406 1707 412 1708
rect 408 1703 410 1707
rect 111 1702 115 1703
rect 111 1697 115 1698
rect 279 1702 283 1703
rect 279 1697 283 1698
rect 319 1702 323 1703
rect 319 1697 323 1698
rect 359 1702 363 1703
rect 359 1697 363 1698
rect 399 1702 403 1703
rect 399 1697 403 1698
rect 407 1702 411 1703
rect 407 1697 411 1698
rect 112 1690 114 1697
rect 278 1696 284 1697
rect 278 1692 279 1696
rect 283 1692 284 1696
rect 278 1691 284 1692
rect 318 1696 324 1697
rect 318 1692 319 1696
rect 323 1692 324 1696
rect 318 1691 324 1692
rect 358 1696 364 1697
rect 358 1692 359 1696
rect 363 1692 364 1696
rect 358 1691 364 1692
rect 398 1696 404 1697
rect 398 1692 399 1696
rect 403 1692 404 1696
rect 398 1691 404 1692
rect 110 1689 116 1690
rect 110 1685 111 1689
rect 115 1685 116 1689
rect 110 1684 116 1685
rect 436 1676 438 1758
rect 446 1755 447 1759
rect 451 1755 452 1759
rect 458 1759 459 1763
rect 463 1759 464 1763
rect 488 1760 490 1769
rect 498 1763 504 1764
rect 458 1758 464 1759
rect 486 1759 492 1760
rect 446 1754 452 1755
rect 460 1732 462 1758
rect 486 1755 487 1759
rect 491 1755 492 1759
rect 498 1759 499 1763
rect 503 1759 504 1763
rect 528 1760 530 1769
rect 538 1763 544 1764
rect 498 1758 504 1759
rect 526 1759 532 1760
rect 486 1754 492 1755
rect 500 1732 502 1758
rect 526 1755 527 1759
rect 531 1755 532 1759
rect 538 1759 539 1763
rect 543 1759 544 1763
rect 568 1760 570 1769
rect 578 1763 584 1764
rect 538 1758 544 1759
rect 566 1759 572 1760
rect 526 1754 532 1755
rect 540 1732 542 1758
rect 566 1755 567 1759
rect 571 1755 572 1759
rect 578 1759 579 1763
rect 583 1759 584 1763
rect 608 1760 610 1769
rect 618 1763 624 1764
rect 578 1758 584 1759
rect 606 1759 612 1760
rect 566 1754 572 1755
rect 580 1732 582 1758
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 618 1759 619 1763
rect 623 1759 624 1763
rect 648 1760 650 1769
rect 658 1763 664 1764
rect 618 1758 624 1759
rect 646 1759 652 1760
rect 606 1754 612 1755
rect 620 1732 622 1758
rect 646 1755 647 1759
rect 651 1755 652 1759
rect 658 1759 659 1763
rect 663 1759 664 1763
rect 658 1758 664 1759
rect 646 1754 652 1755
rect 660 1732 662 1758
rect 676 1732 678 1778
rect 688 1775 690 1784
rect 760 1775 762 1784
rect 832 1775 834 1784
rect 870 1783 871 1787
rect 875 1783 876 1787
rect 902 1785 903 1789
rect 907 1785 908 1789
rect 902 1784 908 1785
rect 928 1784 930 1802
rect 870 1782 876 1783
rect 904 1775 906 1784
rect 926 1783 932 1784
rect 926 1779 927 1783
rect 931 1779 932 1783
rect 926 1778 932 1779
rect 687 1774 691 1775
rect 687 1769 691 1770
rect 695 1774 699 1775
rect 695 1769 699 1770
rect 751 1774 755 1775
rect 751 1769 755 1770
rect 759 1774 763 1775
rect 759 1769 763 1770
rect 807 1774 811 1775
rect 807 1769 811 1770
rect 831 1774 835 1775
rect 831 1769 835 1770
rect 871 1774 875 1775
rect 871 1769 875 1770
rect 903 1774 907 1775
rect 903 1769 907 1770
rect 935 1774 939 1775
rect 935 1769 939 1770
rect 696 1760 698 1769
rect 742 1763 748 1764
rect 694 1759 700 1760
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 742 1759 743 1763
rect 747 1759 748 1763
rect 752 1760 754 1769
rect 798 1763 804 1764
rect 742 1758 748 1759
rect 750 1759 756 1760
rect 694 1754 700 1755
rect 744 1732 746 1758
rect 750 1755 751 1759
rect 755 1755 756 1759
rect 798 1759 799 1763
rect 803 1759 804 1763
rect 808 1760 810 1769
rect 862 1763 868 1764
rect 798 1758 804 1759
rect 806 1759 812 1760
rect 750 1754 756 1755
rect 800 1732 802 1758
rect 806 1755 807 1759
rect 811 1755 812 1759
rect 862 1759 863 1763
rect 867 1759 868 1763
rect 872 1760 874 1769
rect 926 1763 932 1764
rect 862 1758 868 1759
rect 870 1759 876 1760
rect 806 1754 812 1755
rect 864 1732 866 1758
rect 870 1755 871 1759
rect 875 1755 876 1759
rect 926 1759 927 1763
rect 931 1759 932 1763
rect 936 1760 938 1769
rect 960 1764 962 1810
rect 974 1789 980 1790
rect 974 1785 975 1789
rect 979 1785 980 1789
rect 974 1784 980 1785
rect 1046 1789 1052 1790
rect 1046 1785 1047 1789
rect 1051 1785 1052 1789
rect 1046 1784 1052 1785
rect 1072 1784 1074 1866
rect 1238 1859 1244 1860
rect 1238 1855 1239 1859
rect 1243 1855 1244 1859
rect 1280 1855 1282 1870
rect 1342 1868 1348 1869
rect 1342 1864 1343 1868
rect 1347 1864 1348 1868
rect 1342 1863 1348 1864
rect 1344 1855 1346 1863
rect 1238 1854 1244 1855
rect 1279 1854 1283 1855
rect 1126 1852 1132 1853
rect 1126 1848 1127 1852
rect 1131 1848 1132 1852
rect 1126 1847 1132 1848
rect 1128 1843 1130 1847
rect 1240 1843 1242 1854
rect 1279 1849 1283 1850
rect 1343 1854 1347 1855
rect 1343 1849 1347 1850
rect 1359 1854 1363 1855
rect 1359 1849 1363 1850
rect 1127 1842 1131 1843
rect 1127 1837 1131 1838
rect 1191 1842 1195 1843
rect 1191 1837 1195 1838
rect 1239 1842 1243 1843
rect 1280 1842 1282 1849
rect 1358 1848 1364 1849
rect 1358 1844 1359 1848
rect 1363 1844 1364 1848
rect 1358 1843 1364 1844
rect 1239 1837 1243 1838
rect 1278 1841 1284 1842
rect 1278 1837 1279 1841
rect 1283 1837 1284 1841
rect 1126 1836 1132 1837
rect 1126 1832 1127 1836
rect 1131 1832 1132 1836
rect 1126 1831 1132 1832
rect 1190 1836 1196 1837
rect 1190 1832 1191 1836
rect 1195 1832 1196 1836
rect 1190 1831 1196 1832
rect 1240 1830 1242 1837
rect 1278 1836 1284 1837
rect 1238 1829 1244 1830
rect 1238 1825 1239 1829
rect 1243 1825 1244 1829
rect 1372 1828 1374 1914
rect 1382 1911 1383 1915
rect 1387 1911 1388 1915
rect 1394 1915 1395 1919
rect 1399 1915 1400 1919
rect 1424 1916 1426 1925
rect 1434 1919 1440 1920
rect 1394 1914 1400 1915
rect 1422 1915 1428 1916
rect 1382 1910 1388 1911
rect 1396 1888 1398 1914
rect 1422 1911 1423 1915
rect 1427 1911 1428 1915
rect 1434 1915 1435 1919
rect 1439 1915 1440 1919
rect 1464 1916 1466 1925
rect 1474 1919 1480 1920
rect 1434 1914 1440 1915
rect 1462 1915 1468 1916
rect 1422 1910 1428 1911
rect 1436 1888 1438 1914
rect 1462 1911 1463 1915
rect 1467 1911 1468 1915
rect 1474 1915 1475 1919
rect 1479 1915 1480 1919
rect 1512 1916 1514 1925
rect 1474 1914 1480 1915
rect 1510 1915 1516 1916
rect 1462 1910 1468 1911
rect 1476 1888 1478 1914
rect 1510 1911 1511 1915
rect 1515 1911 1516 1915
rect 1510 1910 1516 1911
rect 1536 1888 1538 1938
rect 1560 1931 1562 1944
rect 1574 1943 1580 1944
rect 1574 1939 1575 1943
rect 1579 1939 1580 1943
rect 1574 1938 1580 1939
rect 1600 1931 1602 1944
rect 1614 1943 1620 1944
rect 1614 1939 1615 1943
rect 1619 1939 1620 1943
rect 1614 1938 1620 1939
rect 1640 1931 1642 1944
rect 1654 1943 1660 1944
rect 1654 1939 1655 1943
rect 1659 1939 1660 1943
rect 1654 1938 1660 1939
rect 1680 1931 1682 1944
rect 1694 1943 1700 1944
rect 1694 1939 1695 1943
rect 1699 1939 1700 1943
rect 1694 1938 1700 1939
rect 1720 1931 1722 1944
rect 1734 1943 1740 1944
rect 1734 1939 1735 1943
rect 1739 1939 1740 1943
rect 1734 1938 1740 1939
rect 1768 1931 1770 1944
rect 1782 1943 1788 1944
rect 1782 1939 1783 1943
rect 1787 1939 1788 1943
rect 1782 1938 1788 1939
rect 1824 1931 1826 1944
rect 1838 1943 1844 1944
rect 1838 1939 1839 1943
rect 1843 1939 1844 1943
rect 1838 1938 1844 1939
rect 1872 1931 1874 1944
rect 1878 1943 1884 1944
rect 1878 1939 1879 1943
rect 1883 1939 1884 1943
rect 1878 1938 1884 1939
rect 1920 1931 1922 1944
rect 1968 1931 1970 1944
rect 2016 1931 2018 1944
rect 2022 1943 2028 1944
rect 2022 1939 2023 1943
rect 2027 1939 2028 1943
rect 2022 1938 2028 1939
rect 1559 1930 1563 1931
rect 1559 1925 1563 1926
rect 1567 1930 1571 1931
rect 1567 1925 1571 1926
rect 1599 1930 1603 1931
rect 1599 1925 1603 1926
rect 1631 1930 1635 1931
rect 1631 1925 1635 1926
rect 1639 1930 1643 1931
rect 1639 1925 1643 1926
rect 1679 1930 1683 1931
rect 1679 1925 1683 1926
rect 1711 1930 1715 1931
rect 1711 1925 1715 1926
rect 1719 1930 1723 1931
rect 1719 1925 1723 1926
rect 1767 1930 1771 1931
rect 1767 1925 1771 1926
rect 1807 1930 1811 1931
rect 1807 1925 1811 1926
rect 1823 1930 1827 1931
rect 1823 1925 1827 1926
rect 1871 1930 1875 1931
rect 1871 1925 1875 1926
rect 1919 1930 1923 1931
rect 1919 1925 1923 1926
rect 1967 1930 1971 1931
rect 1967 1925 1971 1926
rect 2015 1930 2019 1931
rect 2015 1925 2019 1926
rect 2031 1930 2035 1931
rect 2031 1925 2035 1926
rect 1558 1919 1564 1920
rect 1558 1915 1559 1919
rect 1563 1915 1564 1919
rect 1568 1916 1570 1925
rect 1622 1919 1628 1920
rect 1558 1914 1564 1915
rect 1566 1915 1572 1916
rect 1560 1888 1562 1914
rect 1566 1911 1567 1915
rect 1571 1911 1572 1915
rect 1622 1915 1623 1919
rect 1627 1915 1628 1919
rect 1632 1916 1634 1925
rect 1642 1919 1648 1920
rect 1622 1914 1628 1915
rect 1630 1915 1636 1916
rect 1566 1910 1572 1911
rect 1624 1888 1626 1914
rect 1630 1911 1631 1915
rect 1635 1911 1636 1915
rect 1642 1915 1643 1919
rect 1647 1915 1648 1919
rect 1712 1916 1714 1925
rect 1798 1919 1804 1920
rect 1642 1914 1648 1915
rect 1710 1915 1716 1916
rect 1630 1910 1636 1911
rect 1644 1896 1646 1914
rect 1710 1911 1711 1915
rect 1715 1911 1716 1915
rect 1798 1915 1799 1919
rect 1803 1915 1804 1919
rect 1808 1916 1810 1925
rect 1910 1919 1916 1920
rect 1798 1914 1804 1915
rect 1806 1915 1812 1916
rect 1710 1910 1716 1911
rect 1642 1895 1648 1896
rect 1642 1891 1643 1895
rect 1647 1891 1648 1895
rect 1642 1890 1648 1891
rect 1800 1888 1802 1914
rect 1806 1911 1807 1915
rect 1811 1911 1812 1915
rect 1910 1915 1911 1919
rect 1915 1915 1916 1919
rect 1920 1916 1922 1925
rect 2022 1919 2028 1920
rect 1910 1914 1916 1915
rect 1918 1915 1924 1916
rect 1806 1910 1812 1911
rect 1912 1888 1914 1914
rect 1918 1911 1919 1915
rect 1923 1911 1924 1915
rect 2022 1915 2023 1919
rect 2027 1915 2028 1919
rect 2032 1916 2034 1925
rect 2048 1920 2050 1962
rect 2054 1949 2060 1950
rect 2054 1945 2055 1949
rect 2059 1945 2060 1949
rect 2054 1944 2060 1945
rect 2056 1931 2058 1944
rect 2070 1943 2076 1944
rect 2070 1939 2071 1943
rect 2075 1939 2076 1943
rect 2070 1938 2076 1939
rect 2055 1930 2059 1931
rect 2055 1925 2059 1926
rect 2046 1919 2052 1920
rect 2022 1914 2028 1915
rect 2030 1915 2036 1916
rect 1918 1910 1924 1911
rect 2024 1888 2026 1914
rect 2030 1911 2031 1915
rect 2035 1911 2036 1915
rect 2046 1915 2047 1919
rect 2051 1915 2052 1919
rect 2046 1914 2052 1915
rect 2030 1910 2036 1911
rect 2072 1888 2074 1938
rect 2084 1924 2086 1970
rect 2094 1949 2100 1950
rect 2094 1945 2095 1949
rect 2099 1945 2100 1949
rect 2094 1944 2100 1945
rect 2104 1944 2106 1970
rect 2142 1949 2148 1950
rect 2142 1945 2143 1949
rect 2147 1945 2148 1949
rect 2142 1944 2148 1945
rect 2190 1949 2196 1950
rect 2190 1945 2191 1949
rect 2195 1945 2196 1949
rect 2190 1944 2196 1945
rect 2216 1944 2218 2014
rect 2238 2008 2244 2009
rect 2238 2004 2239 2008
rect 2243 2004 2244 2008
rect 2238 2003 2244 2004
rect 2278 2008 2284 2009
rect 2278 2004 2279 2008
rect 2283 2004 2284 2008
rect 2278 2003 2284 2004
rect 2239 2002 2243 2003
rect 2239 1997 2243 1998
rect 2279 2002 2283 2003
rect 2279 1997 2283 1998
rect 2238 1996 2244 1997
rect 2238 1992 2239 1996
rect 2243 1992 2244 1996
rect 2238 1991 2244 1992
rect 2278 1996 2284 1997
rect 2278 1992 2279 1996
rect 2283 1992 2284 1996
rect 2278 1991 2284 1992
rect 2296 1976 2298 2054
rect 2318 2051 2319 2055
rect 2323 2051 2324 2055
rect 2346 2055 2347 2059
rect 2351 2055 2352 2059
rect 2360 2056 2362 2065
rect 2370 2059 2376 2060
rect 2346 2054 2352 2055
rect 2358 2055 2364 2056
rect 2318 2050 2324 2051
rect 2358 2051 2359 2055
rect 2363 2051 2364 2055
rect 2370 2055 2371 2059
rect 2375 2055 2376 2059
rect 2370 2054 2376 2055
rect 2358 2050 2364 2051
rect 2372 2028 2374 2054
rect 2408 2033 2410 2065
rect 2406 2032 2412 2033
rect 2406 2028 2407 2032
rect 2411 2028 2412 2032
rect 2370 2027 2376 2028
rect 2370 2023 2371 2027
rect 2375 2023 2376 2027
rect 2370 2022 2376 2023
rect 2382 2027 2388 2028
rect 2406 2027 2412 2028
rect 2382 2023 2383 2027
rect 2387 2023 2388 2027
rect 2382 2022 2388 2023
rect 2318 2008 2324 2009
rect 2318 2004 2319 2008
rect 2323 2004 2324 2008
rect 2318 2003 2324 2004
rect 2358 2008 2364 2009
rect 2358 2004 2359 2008
rect 2363 2004 2364 2008
rect 2358 2003 2364 2004
rect 2319 2002 2323 2003
rect 2319 1997 2323 1998
rect 2359 2002 2363 2003
rect 2359 1997 2363 1998
rect 2318 1996 2324 1997
rect 2318 1992 2319 1996
rect 2323 1992 2324 1996
rect 2318 1991 2324 1992
rect 2358 1996 2364 1997
rect 2358 1992 2359 1996
rect 2363 1992 2364 1996
rect 2358 1991 2364 1992
rect 2294 1975 2300 1976
rect 2294 1971 2295 1975
rect 2299 1971 2300 1975
rect 2294 1970 2300 1971
rect 2326 1975 2332 1976
rect 2326 1971 2327 1975
rect 2331 1971 2332 1975
rect 2326 1970 2332 1971
rect 2366 1975 2372 1976
rect 2366 1971 2367 1975
rect 2371 1971 2372 1975
rect 2366 1970 2372 1971
rect 2286 1967 2292 1968
rect 2286 1963 2287 1967
rect 2291 1963 2292 1967
rect 2286 1962 2292 1963
rect 2238 1949 2244 1950
rect 2238 1945 2239 1949
rect 2243 1945 2244 1949
rect 2238 1944 2244 1945
rect 2278 1949 2284 1950
rect 2278 1945 2279 1949
rect 2283 1945 2284 1949
rect 2278 1944 2284 1945
rect 2288 1944 2290 1962
rect 2318 1949 2324 1950
rect 2318 1945 2319 1949
rect 2323 1945 2324 1949
rect 2318 1944 2324 1945
rect 2328 1944 2330 1970
rect 2358 1949 2364 1950
rect 2358 1945 2359 1949
rect 2363 1945 2364 1949
rect 2358 1944 2364 1945
rect 2368 1944 2370 1970
rect 2384 1944 2386 2022
rect 2406 2015 2412 2016
rect 2406 2011 2407 2015
rect 2411 2011 2412 2015
rect 2406 2010 2412 2011
rect 2408 2003 2410 2010
rect 2407 2002 2411 2003
rect 2407 1997 2411 1998
rect 2408 1990 2410 1997
rect 2406 1989 2412 1990
rect 2406 1985 2407 1989
rect 2411 1985 2412 1989
rect 2406 1984 2412 1985
rect 2406 1972 2412 1973
rect 2406 1968 2407 1972
rect 2411 1968 2412 1972
rect 2406 1967 2412 1968
rect 2096 1931 2098 1944
rect 2102 1943 2108 1944
rect 2102 1939 2103 1943
rect 2107 1939 2108 1943
rect 2102 1938 2108 1939
rect 2144 1931 2146 1944
rect 2192 1931 2194 1944
rect 2214 1943 2220 1944
rect 2214 1939 2215 1943
rect 2219 1939 2220 1943
rect 2214 1938 2220 1939
rect 2240 1931 2242 1944
rect 2280 1931 2282 1944
rect 2286 1943 2292 1944
rect 2286 1939 2287 1943
rect 2291 1939 2292 1943
rect 2286 1938 2292 1939
rect 2320 1931 2322 1944
rect 2326 1943 2332 1944
rect 2326 1939 2327 1943
rect 2331 1939 2332 1943
rect 2326 1938 2332 1939
rect 2360 1931 2362 1944
rect 2366 1943 2372 1944
rect 2366 1939 2367 1943
rect 2371 1939 2372 1943
rect 2366 1938 2372 1939
rect 2382 1943 2388 1944
rect 2382 1939 2383 1943
rect 2387 1939 2388 1943
rect 2382 1938 2388 1939
rect 2408 1931 2410 1967
rect 2095 1930 2099 1931
rect 2095 1925 2099 1926
rect 2143 1930 2147 1931
rect 2143 1925 2147 1926
rect 2151 1930 2155 1931
rect 2151 1925 2155 1926
rect 2191 1930 2195 1931
rect 2191 1925 2195 1926
rect 2239 1930 2243 1931
rect 2239 1925 2243 1926
rect 2279 1930 2283 1931
rect 2279 1925 2283 1926
rect 2319 1930 2323 1931
rect 2319 1925 2323 1926
rect 2359 1930 2363 1931
rect 2359 1925 2363 1926
rect 2407 1930 2411 1931
rect 2407 1925 2411 1926
rect 2082 1923 2088 1924
rect 2082 1919 2083 1923
rect 2087 1919 2088 1923
rect 2082 1918 2088 1919
rect 2152 1916 2154 1925
rect 2150 1915 2156 1916
rect 2150 1911 2151 1915
rect 2155 1911 2156 1915
rect 2150 1910 2156 1911
rect 2408 1893 2410 1925
rect 2406 1892 2412 1893
rect 2406 1888 2407 1892
rect 2411 1888 2412 1892
rect 1394 1887 1400 1888
rect 1394 1883 1395 1887
rect 1399 1883 1400 1887
rect 1394 1882 1400 1883
rect 1434 1887 1440 1888
rect 1434 1883 1435 1887
rect 1439 1883 1440 1887
rect 1434 1882 1440 1883
rect 1474 1887 1480 1888
rect 1474 1883 1475 1887
rect 1479 1883 1480 1887
rect 1474 1882 1480 1883
rect 1534 1887 1540 1888
rect 1534 1883 1535 1887
rect 1539 1883 1540 1887
rect 1534 1882 1540 1883
rect 1558 1887 1564 1888
rect 1558 1883 1559 1887
rect 1563 1883 1564 1887
rect 1558 1882 1564 1883
rect 1622 1887 1628 1888
rect 1622 1883 1623 1887
rect 1627 1883 1628 1887
rect 1622 1882 1628 1883
rect 1798 1887 1804 1888
rect 1798 1883 1799 1887
rect 1803 1883 1804 1887
rect 1798 1882 1804 1883
rect 1910 1887 1916 1888
rect 1910 1883 1911 1887
rect 1915 1883 1916 1887
rect 1910 1882 1916 1883
rect 2022 1887 2028 1888
rect 2022 1883 2023 1887
rect 2027 1883 2028 1887
rect 2022 1882 2028 1883
rect 2070 1887 2076 1888
rect 2406 1887 2412 1888
rect 2070 1883 2071 1887
rect 2075 1883 2076 1887
rect 2070 1882 2076 1883
rect 2406 1875 2412 1876
rect 2406 1871 2407 1875
rect 2411 1871 2412 1875
rect 2406 1870 2412 1871
rect 1382 1868 1388 1869
rect 1382 1864 1383 1868
rect 1387 1864 1388 1868
rect 1382 1863 1388 1864
rect 1422 1868 1428 1869
rect 1422 1864 1423 1868
rect 1427 1864 1428 1868
rect 1422 1863 1428 1864
rect 1462 1868 1468 1869
rect 1462 1864 1463 1868
rect 1467 1864 1468 1868
rect 1462 1863 1468 1864
rect 1510 1868 1516 1869
rect 1510 1864 1511 1868
rect 1515 1864 1516 1868
rect 1510 1863 1516 1864
rect 1566 1868 1572 1869
rect 1566 1864 1567 1868
rect 1571 1864 1572 1868
rect 1566 1863 1572 1864
rect 1630 1868 1636 1869
rect 1630 1864 1631 1868
rect 1635 1864 1636 1868
rect 1630 1863 1636 1864
rect 1710 1868 1716 1869
rect 1710 1864 1711 1868
rect 1715 1864 1716 1868
rect 1710 1863 1716 1864
rect 1806 1868 1812 1869
rect 1806 1864 1807 1868
rect 1811 1864 1812 1868
rect 1806 1863 1812 1864
rect 1918 1868 1924 1869
rect 1918 1864 1919 1868
rect 1923 1864 1924 1868
rect 1918 1863 1924 1864
rect 2030 1868 2036 1869
rect 2030 1864 2031 1868
rect 2035 1864 2036 1868
rect 2030 1863 2036 1864
rect 2150 1868 2156 1869
rect 2150 1864 2151 1868
rect 2155 1864 2156 1868
rect 2150 1863 2156 1864
rect 1384 1855 1386 1863
rect 1424 1855 1426 1863
rect 1464 1855 1466 1863
rect 1512 1855 1514 1863
rect 1568 1855 1570 1863
rect 1632 1855 1634 1863
rect 1712 1855 1714 1863
rect 1808 1855 1810 1863
rect 1920 1855 1922 1863
rect 2032 1855 2034 1863
rect 2152 1855 2154 1863
rect 2408 1855 2410 1870
rect 1383 1854 1387 1855
rect 1383 1849 1387 1850
rect 1399 1854 1403 1855
rect 1399 1849 1403 1850
rect 1423 1854 1427 1855
rect 1423 1849 1427 1850
rect 1447 1854 1451 1855
rect 1447 1849 1451 1850
rect 1463 1854 1467 1855
rect 1463 1849 1467 1850
rect 1503 1854 1507 1855
rect 1503 1849 1507 1850
rect 1511 1854 1515 1855
rect 1511 1849 1515 1850
rect 1559 1854 1563 1855
rect 1559 1849 1563 1850
rect 1567 1854 1571 1855
rect 1567 1849 1571 1850
rect 1615 1854 1619 1855
rect 1615 1849 1619 1850
rect 1631 1854 1635 1855
rect 1631 1849 1635 1850
rect 1671 1854 1675 1855
rect 1671 1849 1675 1850
rect 1711 1854 1715 1855
rect 1711 1849 1715 1850
rect 1727 1854 1731 1855
rect 1727 1849 1731 1850
rect 1783 1854 1787 1855
rect 1783 1849 1787 1850
rect 1807 1854 1811 1855
rect 1807 1849 1811 1850
rect 1839 1854 1843 1855
rect 1839 1849 1843 1850
rect 1895 1854 1899 1855
rect 1895 1849 1899 1850
rect 1919 1854 1923 1855
rect 1919 1849 1923 1850
rect 1951 1854 1955 1855
rect 1951 1849 1955 1850
rect 2031 1854 2035 1855
rect 2031 1849 2035 1850
rect 2151 1854 2155 1855
rect 2151 1849 2155 1850
rect 2407 1854 2411 1855
rect 2407 1849 2411 1850
rect 1398 1848 1404 1849
rect 1398 1844 1399 1848
rect 1403 1844 1404 1848
rect 1398 1843 1404 1844
rect 1446 1848 1452 1849
rect 1446 1844 1447 1848
rect 1451 1844 1452 1848
rect 1446 1843 1452 1844
rect 1502 1848 1508 1849
rect 1502 1844 1503 1848
rect 1507 1844 1508 1848
rect 1502 1843 1508 1844
rect 1558 1848 1564 1849
rect 1558 1844 1559 1848
rect 1563 1844 1564 1848
rect 1558 1843 1564 1844
rect 1614 1848 1620 1849
rect 1614 1844 1615 1848
rect 1619 1844 1620 1848
rect 1614 1843 1620 1844
rect 1670 1848 1676 1849
rect 1670 1844 1671 1848
rect 1675 1844 1676 1848
rect 1670 1843 1676 1844
rect 1726 1848 1732 1849
rect 1726 1844 1727 1848
rect 1731 1844 1732 1848
rect 1726 1843 1732 1844
rect 1782 1848 1788 1849
rect 1782 1844 1783 1848
rect 1787 1844 1788 1848
rect 1782 1843 1788 1844
rect 1838 1848 1844 1849
rect 1838 1844 1839 1848
rect 1843 1844 1844 1848
rect 1838 1843 1844 1844
rect 1894 1848 1900 1849
rect 1894 1844 1895 1848
rect 1899 1844 1900 1848
rect 1894 1843 1900 1844
rect 1950 1848 1956 1849
rect 1950 1844 1951 1848
rect 1955 1844 1956 1848
rect 1950 1843 1956 1844
rect 2408 1842 2410 1849
rect 2406 1841 2412 1842
rect 2406 1837 2407 1841
rect 2411 1837 2412 1841
rect 2406 1836 2412 1837
rect 1370 1827 1376 1828
rect 1238 1824 1244 1825
rect 1278 1824 1284 1825
rect 1278 1820 1279 1824
rect 1283 1820 1284 1824
rect 1370 1823 1371 1827
rect 1375 1823 1376 1827
rect 1370 1822 1376 1823
rect 1406 1827 1412 1828
rect 1406 1823 1407 1827
rect 1411 1823 1412 1827
rect 1406 1822 1412 1823
rect 1742 1827 1748 1828
rect 1742 1823 1743 1827
rect 1747 1823 1748 1827
rect 1742 1822 1748 1823
rect 1798 1827 1804 1828
rect 1798 1823 1799 1827
rect 1803 1823 1804 1827
rect 1798 1822 1804 1823
rect 1854 1827 1860 1828
rect 1854 1823 1855 1827
rect 1859 1823 1860 1827
rect 1854 1822 1860 1823
rect 1902 1827 1908 1828
rect 1902 1823 1903 1827
rect 1907 1823 1908 1827
rect 1902 1822 1908 1823
rect 2406 1824 2412 1825
rect 1278 1819 1284 1820
rect 1206 1815 1212 1816
rect 1206 1811 1207 1815
rect 1211 1811 1212 1815
rect 1206 1810 1212 1811
rect 1238 1812 1244 1813
rect 1150 1807 1156 1808
rect 1150 1803 1151 1807
rect 1155 1803 1156 1807
rect 1150 1802 1156 1803
rect 1170 1807 1176 1808
rect 1170 1803 1171 1807
rect 1175 1803 1176 1807
rect 1170 1802 1176 1803
rect 1126 1789 1132 1790
rect 1126 1785 1127 1789
rect 1131 1785 1132 1789
rect 1126 1784 1132 1785
rect 1152 1784 1154 1802
rect 976 1775 978 1784
rect 1048 1775 1050 1784
rect 1070 1783 1076 1784
rect 1070 1779 1071 1783
rect 1075 1779 1076 1783
rect 1070 1778 1076 1779
rect 1128 1775 1130 1784
rect 1150 1783 1156 1784
rect 1150 1779 1151 1783
rect 1155 1779 1156 1783
rect 1150 1778 1156 1779
rect 975 1774 979 1775
rect 975 1769 979 1770
rect 999 1774 1003 1775
rect 999 1769 1003 1770
rect 1047 1774 1051 1775
rect 1047 1769 1051 1770
rect 1071 1774 1075 1775
rect 1071 1769 1075 1770
rect 1127 1774 1131 1775
rect 1127 1769 1131 1770
rect 1143 1774 1147 1775
rect 1143 1769 1147 1770
rect 958 1763 964 1764
rect 926 1758 932 1759
rect 934 1759 940 1760
rect 870 1754 876 1755
rect 928 1732 930 1758
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 958 1759 959 1763
rect 963 1759 964 1763
rect 1000 1760 1002 1769
rect 1072 1760 1074 1769
rect 1126 1763 1132 1764
rect 958 1758 964 1759
rect 998 1759 1004 1760
rect 934 1754 940 1755
rect 998 1755 999 1759
rect 1003 1755 1004 1759
rect 998 1754 1004 1755
rect 1070 1759 1076 1760
rect 1070 1755 1071 1759
rect 1075 1755 1076 1759
rect 1126 1759 1127 1763
rect 1131 1759 1132 1763
rect 1144 1760 1146 1769
rect 1172 1764 1174 1802
rect 1190 1789 1196 1790
rect 1190 1785 1191 1789
rect 1195 1785 1196 1789
rect 1190 1784 1196 1785
rect 1208 1784 1210 1810
rect 1238 1808 1239 1812
rect 1243 1808 1244 1812
rect 1238 1807 1244 1808
rect 1192 1775 1194 1784
rect 1206 1783 1212 1784
rect 1206 1779 1207 1783
rect 1211 1779 1212 1783
rect 1206 1778 1212 1779
rect 1240 1775 1242 1807
rect 1280 1775 1282 1819
rect 1358 1801 1364 1802
rect 1358 1797 1359 1801
rect 1363 1797 1364 1801
rect 1358 1796 1364 1797
rect 1398 1801 1404 1802
rect 1398 1797 1399 1801
rect 1403 1797 1404 1801
rect 1398 1796 1404 1797
rect 1408 1796 1410 1822
rect 1446 1801 1452 1802
rect 1446 1797 1447 1801
rect 1451 1797 1452 1801
rect 1446 1796 1452 1797
rect 1502 1801 1508 1802
rect 1502 1797 1503 1801
rect 1507 1797 1508 1801
rect 1502 1796 1508 1797
rect 1558 1801 1564 1802
rect 1558 1797 1559 1801
rect 1563 1797 1564 1801
rect 1558 1796 1564 1797
rect 1614 1801 1620 1802
rect 1614 1797 1615 1801
rect 1619 1797 1620 1801
rect 1614 1796 1620 1797
rect 1670 1801 1676 1802
rect 1670 1797 1671 1801
rect 1675 1797 1676 1801
rect 1670 1796 1676 1797
rect 1726 1801 1732 1802
rect 1726 1797 1727 1801
rect 1731 1797 1732 1801
rect 1726 1796 1732 1797
rect 1744 1796 1746 1822
rect 1782 1801 1788 1802
rect 1782 1797 1783 1801
rect 1787 1797 1788 1801
rect 1782 1796 1788 1797
rect 1800 1796 1802 1822
rect 1838 1801 1844 1802
rect 1838 1797 1839 1801
rect 1843 1797 1844 1801
rect 1838 1796 1844 1797
rect 1856 1796 1858 1822
rect 1894 1801 1900 1802
rect 1894 1797 1895 1801
rect 1899 1797 1900 1801
rect 1894 1796 1900 1797
rect 1360 1775 1362 1796
rect 1400 1775 1402 1796
rect 1406 1795 1412 1796
rect 1406 1791 1407 1795
rect 1411 1791 1412 1795
rect 1406 1790 1412 1791
rect 1448 1775 1450 1796
rect 1504 1775 1506 1796
rect 1560 1775 1562 1796
rect 1602 1795 1608 1796
rect 1602 1791 1603 1795
rect 1607 1791 1608 1795
rect 1602 1790 1608 1791
rect 1191 1774 1195 1775
rect 1191 1769 1195 1770
rect 1239 1774 1243 1775
rect 1239 1769 1243 1770
rect 1279 1774 1283 1775
rect 1279 1769 1283 1770
rect 1303 1774 1307 1775
rect 1303 1769 1307 1770
rect 1343 1774 1347 1775
rect 1343 1769 1347 1770
rect 1359 1774 1363 1775
rect 1359 1769 1363 1770
rect 1391 1774 1395 1775
rect 1391 1769 1395 1770
rect 1399 1774 1403 1775
rect 1399 1769 1403 1770
rect 1447 1774 1451 1775
rect 1447 1769 1451 1770
rect 1455 1774 1459 1775
rect 1455 1769 1459 1770
rect 1503 1774 1507 1775
rect 1503 1769 1507 1770
rect 1519 1774 1523 1775
rect 1519 1769 1523 1770
rect 1559 1774 1563 1775
rect 1559 1769 1563 1770
rect 1583 1774 1587 1775
rect 1583 1769 1587 1770
rect 1170 1763 1176 1764
rect 1126 1758 1132 1759
rect 1142 1759 1148 1760
rect 1070 1754 1076 1755
rect 1094 1751 1100 1752
rect 1094 1747 1095 1751
rect 1099 1747 1100 1751
rect 1094 1746 1100 1747
rect 1096 1732 1098 1746
rect 1128 1732 1130 1758
rect 1142 1755 1143 1759
rect 1147 1755 1148 1759
rect 1170 1759 1171 1763
rect 1175 1759 1176 1763
rect 1192 1760 1194 1769
rect 1202 1763 1208 1764
rect 1170 1758 1176 1759
rect 1190 1759 1196 1760
rect 1142 1754 1148 1755
rect 1190 1755 1191 1759
rect 1195 1755 1196 1759
rect 1202 1759 1203 1763
rect 1207 1759 1208 1763
rect 1202 1758 1208 1759
rect 1190 1754 1196 1755
rect 1204 1740 1206 1758
rect 1202 1739 1208 1740
rect 1202 1735 1203 1739
rect 1207 1735 1208 1739
rect 1240 1737 1242 1769
rect 1280 1737 1282 1769
rect 1304 1760 1306 1769
rect 1314 1763 1320 1764
rect 1302 1759 1308 1760
rect 1302 1755 1303 1759
rect 1307 1755 1308 1759
rect 1314 1759 1315 1763
rect 1319 1759 1320 1763
rect 1344 1760 1346 1769
rect 1354 1763 1360 1764
rect 1314 1758 1320 1759
rect 1342 1759 1348 1760
rect 1302 1754 1308 1755
rect 1202 1734 1208 1735
rect 1238 1736 1244 1737
rect 1238 1732 1239 1736
rect 1243 1732 1244 1736
rect 458 1731 464 1732
rect 458 1727 459 1731
rect 463 1727 464 1731
rect 458 1726 464 1727
rect 498 1731 504 1732
rect 498 1727 499 1731
rect 503 1727 504 1731
rect 498 1726 504 1727
rect 538 1731 544 1732
rect 538 1727 539 1731
rect 543 1727 544 1731
rect 538 1726 544 1727
rect 578 1731 584 1732
rect 578 1727 579 1731
rect 583 1727 584 1731
rect 578 1726 584 1727
rect 618 1731 624 1732
rect 618 1727 619 1731
rect 623 1727 624 1731
rect 618 1726 624 1727
rect 658 1731 664 1732
rect 658 1727 659 1731
rect 663 1727 664 1731
rect 658 1726 664 1727
rect 674 1731 680 1732
rect 674 1727 675 1731
rect 679 1727 680 1731
rect 674 1726 680 1727
rect 702 1731 708 1732
rect 702 1727 703 1731
rect 707 1727 708 1731
rect 702 1726 708 1727
rect 742 1731 748 1732
rect 742 1727 743 1731
rect 747 1727 748 1731
rect 742 1726 748 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 862 1731 868 1732
rect 862 1727 863 1731
rect 867 1727 868 1731
rect 862 1726 868 1727
rect 926 1731 932 1732
rect 926 1727 927 1731
rect 931 1727 932 1731
rect 926 1726 932 1727
rect 1094 1731 1100 1732
rect 1094 1727 1095 1731
rect 1099 1727 1100 1731
rect 1094 1726 1100 1727
rect 1126 1731 1132 1732
rect 1238 1731 1244 1732
rect 1278 1736 1284 1737
rect 1278 1732 1279 1736
rect 1283 1732 1284 1736
rect 1278 1731 1284 1732
rect 1126 1727 1127 1731
rect 1131 1727 1132 1731
rect 1316 1728 1318 1758
rect 1342 1755 1343 1759
rect 1347 1755 1348 1759
rect 1354 1759 1355 1763
rect 1359 1759 1360 1763
rect 1392 1760 1394 1769
rect 1446 1763 1452 1764
rect 1354 1758 1360 1759
rect 1390 1759 1396 1760
rect 1342 1754 1348 1755
rect 1356 1732 1358 1758
rect 1390 1755 1391 1759
rect 1395 1755 1396 1759
rect 1446 1759 1447 1763
rect 1451 1759 1452 1763
rect 1456 1760 1458 1769
rect 1510 1763 1516 1764
rect 1446 1758 1452 1759
rect 1454 1759 1460 1760
rect 1390 1754 1396 1755
rect 1448 1732 1450 1758
rect 1454 1755 1455 1759
rect 1459 1755 1460 1759
rect 1510 1759 1511 1763
rect 1515 1759 1516 1763
rect 1520 1760 1522 1769
rect 1574 1763 1580 1764
rect 1510 1758 1516 1759
rect 1518 1759 1524 1760
rect 1454 1754 1460 1755
rect 1512 1732 1514 1758
rect 1518 1755 1519 1759
rect 1523 1755 1524 1759
rect 1574 1759 1575 1763
rect 1579 1759 1580 1763
rect 1584 1760 1586 1769
rect 1594 1763 1600 1764
rect 1574 1758 1580 1759
rect 1582 1759 1588 1760
rect 1518 1754 1524 1755
rect 1576 1732 1578 1758
rect 1582 1755 1583 1759
rect 1587 1755 1588 1759
rect 1594 1759 1595 1763
rect 1599 1759 1600 1763
rect 1594 1758 1600 1759
rect 1582 1754 1588 1755
rect 1354 1731 1360 1732
rect 1126 1726 1132 1727
rect 1314 1727 1320 1728
rect 446 1712 452 1713
rect 446 1708 447 1712
rect 451 1708 452 1712
rect 446 1707 452 1708
rect 486 1712 492 1713
rect 486 1708 487 1712
rect 491 1708 492 1712
rect 486 1707 492 1708
rect 526 1712 532 1713
rect 526 1708 527 1712
rect 531 1708 532 1712
rect 526 1707 532 1708
rect 566 1712 572 1713
rect 566 1708 567 1712
rect 571 1708 572 1712
rect 566 1707 572 1708
rect 606 1712 612 1713
rect 606 1708 607 1712
rect 611 1708 612 1712
rect 606 1707 612 1708
rect 646 1712 652 1713
rect 646 1708 647 1712
rect 651 1708 652 1712
rect 646 1707 652 1708
rect 694 1712 700 1713
rect 694 1708 695 1712
rect 699 1708 700 1712
rect 694 1707 700 1708
rect 448 1703 450 1707
rect 488 1703 490 1707
rect 528 1703 530 1707
rect 568 1703 570 1707
rect 608 1703 610 1707
rect 648 1703 650 1707
rect 696 1703 698 1707
rect 447 1702 451 1703
rect 447 1697 451 1698
rect 487 1702 491 1703
rect 487 1697 491 1698
rect 495 1702 499 1703
rect 495 1697 499 1698
rect 527 1702 531 1703
rect 527 1697 531 1698
rect 543 1702 547 1703
rect 543 1697 547 1698
rect 567 1702 571 1703
rect 567 1697 571 1698
rect 591 1702 595 1703
rect 591 1697 595 1698
rect 607 1702 611 1703
rect 607 1697 611 1698
rect 639 1702 643 1703
rect 639 1697 643 1698
rect 647 1702 651 1703
rect 647 1697 651 1698
rect 687 1702 691 1703
rect 687 1697 691 1698
rect 695 1702 699 1703
rect 695 1697 699 1698
rect 446 1696 452 1697
rect 446 1692 447 1696
rect 451 1692 452 1696
rect 446 1691 452 1692
rect 494 1696 500 1697
rect 494 1692 495 1696
rect 499 1692 500 1696
rect 494 1691 500 1692
rect 542 1696 548 1697
rect 542 1692 543 1696
rect 547 1692 548 1696
rect 542 1691 548 1692
rect 590 1696 596 1697
rect 590 1692 591 1696
rect 595 1692 596 1696
rect 590 1691 596 1692
rect 638 1696 644 1697
rect 638 1692 639 1696
rect 643 1692 644 1696
rect 638 1691 644 1692
rect 686 1696 692 1697
rect 686 1692 687 1696
rect 691 1692 692 1696
rect 686 1691 692 1692
rect 566 1683 572 1684
rect 566 1679 567 1683
rect 571 1679 572 1683
rect 566 1678 572 1679
rect 330 1675 336 1676
rect 110 1672 116 1673
rect 110 1668 111 1672
rect 115 1668 116 1672
rect 330 1671 331 1675
rect 335 1671 336 1675
rect 330 1670 336 1671
rect 366 1675 372 1676
rect 366 1671 367 1675
rect 371 1671 372 1675
rect 366 1670 372 1671
rect 434 1675 440 1676
rect 434 1671 435 1675
rect 439 1671 440 1675
rect 434 1670 440 1671
rect 110 1667 116 1668
rect 112 1631 114 1667
rect 278 1649 284 1650
rect 278 1645 279 1649
rect 283 1645 284 1649
rect 278 1644 284 1645
rect 318 1649 324 1650
rect 318 1645 319 1649
rect 323 1645 324 1649
rect 318 1644 324 1645
rect 332 1644 334 1670
rect 358 1649 364 1650
rect 358 1645 359 1649
rect 363 1645 364 1649
rect 358 1644 364 1645
rect 368 1644 370 1670
rect 422 1667 428 1668
rect 422 1663 423 1667
rect 427 1663 428 1667
rect 422 1662 428 1663
rect 398 1649 404 1650
rect 398 1645 399 1649
rect 403 1645 404 1649
rect 398 1644 404 1645
rect 424 1644 426 1662
rect 446 1649 452 1650
rect 446 1645 447 1649
rect 451 1645 452 1649
rect 446 1644 452 1645
rect 494 1649 500 1650
rect 494 1645 495 1649
rect 499 1645 500 1649
rect 494 1644 500 1645
rect 542 1649 548 1650
rect 542 1645 543 1649
rect 547 1645 548 1649
rect 542 1644 548 1645
rect 568 1644 570 1678
rect 590 1649 596 1650
rect 590 1645 591 1649
rect 595 1645 596 1649
rect 590 1644 596 1645
rect 638 1649 644 1650
rect 638 1645 639 1649
rect 643 1645 644 1649
rect 638 1644 644 1645
rect 686 1649 692 1650
rect 686 1645 687 1649
rect 691 1645 692 1649
rect 686 1644 692 1645
rect 704 1644 706 1726
rect 1314 1723 1315 1727
rect 1319 1723 1320 1727
rect 1354 1727 1355 1731
rect 1359 1727 1360 1731
rect 1354 1726 1360 1727
rect 1366 1731 1372 1732
rect 1366 1727 1367 1731
rect 1371 1727 1372 1731
rect 1366 1726 1372 1727
rect 1446 1731 1452 1732
rect 1446 1727 1447 1731
rect 1451 1727 1452 1731
rect 1446 1726 1452 1727
rect 1510 1731 1516 1732
rect 1510 1727 1511 1731
rect 1515 1727 1516 1731
rect 1510 1726 1516 1727
rect 1574 1731 1580 1732
rect 1574 1727 1575 1731
rect 1579 1727 1580 1731
rect 1574 1726 1580 1727
rect 1314 1722 1320 1723
rect 1238 1719 1244 1720
rect 1238 1715 1239 1719
rect 1243 1715 1244 1719
rect 1238 1714 1244 1715
rect 1278 1719 1284 1720
rect 1278 1715 1279 1719
rect 1283 1715 1284 1719
rect 1278 1714 1284 1715
rect 750 1712 756 1713
rect 750 1708 751 1712
rect 755 1708 756 1712
rect 750 1707 756 1708
rect 806 1712 812 1713
rect 806 1708 807 1712
rect 811 1708 812 1712
rect 806 1707 812 1708
rect 870 1712 876 1713
rect 870 1708 871 1712
rect 875 1708 876 1712
rect 870 1707 876 1708
rect 934 1712 940 1713
rect 934 1708 935 1712
rect 939 1708 940 1712
rect 934 1707 940 1708
rect 998 1712 1004 1713
rect 998 1708 999 1712
rect 1003 1708 1004 1712
rect 998 1707 1004 1708
rect 1070 1712 1076 1713
rect 1070 1708 1071 1712
rect 1075 1708 1076 1712
rect 1070 1707 1076 1708
rect 1142 1712 1148 1713
rect 1142 1708 1143 1712
rect 1147 1708 1148 1712
rect 1142 1707 1148 1708
rect 1190 1712 1196 1713
rect 1190 1708 1191 1712
rect 1195 1708 1196 1712
rect 1190 1707 1196 1708
rect 752 1703 754 1707
rect 808 1703 810 1707
rect 872 1703 874 1707
rect 936 1703 938 1707
rect 1000 1703 1002 1707
rect 1072 1703 1074 1707
rect 1144 1703 1146 1707
rect 1192 1703 1194 1707
rect 1240 1703 1242 1714
rect 1280 1703 1282 1714
rect 1302 1712 1308 1713
rect 1302 1708 1303 1712
rect 1307 1708 1308 1712
rect 1302 1707 1308 1708
rect 1342 1712 1348 1713
rect 1342 1708 1343 1712
rect 1347 1708 1348 1712
rect 1342 1707 1348 1708
rect 1304 1703 1306 1707
rect 1344 1703 1346 1707
rect 735 1702 739 1703
rect 735 1697 739 1698
rect 751 1702 755 1703
rect 751 1697 755 1698
rect 783 1702 787 1703
rect 783 1697 787 1698
rect 807 1702 811 1703
rect 807 1697 811 1698
rect 839 1702 843 1703
rect 839 1697 843 1698
rect 871 1702 875 1703
rect 871 1697 875 1698
rect 895 1702 899 1703
rect 895 1697 899 1698
rect 935 1702 939 1703
rect 935 1697 939 1698
rect 999 1702 1003 1703
rect 999 1697 1003 1698
rect 1071 1702 1075 1703
rect 1071 1697 1075 1698
rect 1143 1702 1147 1703
rect 1143 1697 1147 1698
rect 1191 1702 1195 1703
rect 1191 1697 1195 1698
rect 1239 1702 1243 1703
rect 1239 1697 1243 1698
rect 1279 1702 1283 1703
rect 1279 1697 1283 1698
rect 1303 1702 1307 1703
rect 1303 1697 1307 1698
rect 1343 1702 1347 1703
rect 1343 1697 1347 1698
rect 734 1696 740 1697
rect 734 1692 735 1696
rect 739 1692 740 1696
rect 734 1691 740 1692
rect 782 1696 788 1697
rect 782 1692 783 1696
rect 787 1692 788 1696
rect 782 1691 788 1692
rect 838 1696 844 1697
rect 838 1692 839 1696
rect 843 1692 844 1696
rect 838 1691 844 1692
rect 894 1696 900 1697
rect 894 1692 895 1696
rect 899 1692 900 1696
rect 894 1691 900 1692
rect 1240 1690 1242 1697
rect 1280 1690 1282 1697
rect 1302 1696 1308 1697
rect 1302 1692 1303 1696
rect 1307 1692 1308 1696
rect 1302 1691 1308 1692
rect 1342 1696 1348 1697
rect 1342 1692 1343 1696
rect 1347 1692 1348 1696
rect 1342 1691 1348 1692
rect 1238 1689 1244 1690
rect 1238 1685 1239 1689
rect 1243 1685 1244 1689
rect 1238 1684 1244 1685
rect 1278 1689 1284 1690
rect 1278 1685 1279 1689
rect 1283 1685 1284 1689
rect 1278 1684 1284 1685
rect 750 1675 756 1676
rect 750 1671 751 1675
rect 755 1671 756 1675
rect 750 1670 756 1671
rect 798 1675 804 1676
rect 798 1671 799 1675
rect 803 1671 804 1675
rect 798 1670 804 1671
rect 818 1675 824 1676
rect 818 1671 819 1675
rect 823 1671 824 1675
rect 1350 1675 1356 1676
rect 818 1670 824 1671
rect 1238 1672 1244 1673
rect 710 1667 716 1668
rect 710 1663 711 1667
rect 715 1663 716 1667
rect 710 1662 716 1663
rect 712 1644 714 1662
rect 734 1649 740 1650
rect 734 1645 735 1649
rect 739 1645 740 1649
rect 734 1644 740 1645
rect 752 1644 754 1670
rect 782 1649 788 1650
rect 782 1645 783 1649
rect 787 1645 788 1649
rect 782 1644 788 1645
rect 800 1644 802 1670
rect 280 1631 282 1644
rect 320 1631 322 1644
rect 330 1643 336 1644
rect 330 1639 331 1643
rect 335 1639 336 1643
rect 330 1638 336 1639
rect 360 1631 362 1644
rect 366 1643 372 1644
rect 366 1639 367 1643
rect 371 1639 372 1643
rect 366 1638 372 1639
rect 400 1631 402 1644
rect 406 1643 412 1644
rect 406 1639 407 1643
rect 411 1639 412 1643
rect 406 1638 412 1639
rect 422 1643 428 1644
rect 422 1639 423 1643
rect 427 1639 428 1643
rect 422 1638 428 1639
rect 111 1630 115 1631
rect 111 1625 115 1626
rect 135 1630 139 1631
rect 135 1625 139 1626
rect 175 1630 179 1631
rect 175 1625 179 1626
rect 215 1630 219 1631
rect 215 1625 219 1626
rect 255 1630 259 1631
rect 255 1625 259 1626
rect 279 1630 283 1631
rect 279 1625 283 1626
rect 311 1630 315 1631
rect 311 1625 315 1626
rect 319 1630 323 1631
rect 319 1625 323 1626
rect 359 1630 363 1631
rect 359 1625 363 1626
rect 391 1630 395 1631
rect 391 1625 395 1626
rect 399 1630 403 1631
rect 399 1625 403 1626
rect 112 1593 114 1625
rect 136 1616 138 1625
rect 162 1619 168 1620
rect 134 1615 140 1616
rect 134 1611 135 1615
rect 139 1611 140 1615
rect 162 1615 163 1619
rect 167 1615 168 1619
rect 176 1616 178 1625
rect 186 1619 192 1620
rect 162 1614 168 1615
rect 174 1615 180 1616
rect 134 1610 140 1611
rect 164 1596 166 1614
rect 174 1611 175 1615
rect 179 1611 180 1615
rect 186 1615 187 1619
rect 191 1615 192 1619
rect 216 1616 218 1625
rect 256 1616 258 1625
rect 266 1619 272 1620
rect 186 1614 192 1615
rect 214 1615 220 1616
rect 174 1610 180 1611
rect 162 1595 168 1596
rect 110 1592 116 1593
rect 110 1588 111 1592
rect 115 1588 116 1592
rect 162 1591 163 1595
rect 167 1591 168 1595
rect 162 1590 168 1591
rect 110 1587 116 1588
rect 110 1575 116 1576
rect 110 1571 111 1575
rect 115 1571 116 1575
rect 110 1570 116 1571
rect 112 1559 114 1570
rect 134 1568 140 1569
rect 134 1564 135 1568
rect 139 1564 140 1568
rect 134 1563 140 1564
rect 174 1568 180 1569
rect 174 1564 175 1568
rect 179 1564 180 1568
rect 174 1563 180 1564
rect 136 1559 138 1563
rect 176 1559 178 1563
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 135 1558 139 1559
rect 135 1553 139 1554
rect 151 1558 155 1559
rect 151 1553 155 1554
rect 175 1558 179 1559
rect 175 1553 179 1554
rect 112 1546 114 1553
rect 150 1552 156 1553
rect 150 1548 151 1552
rect 155 1548 156 1552
rect 150 1547 156 1548
rect 110 1545 116 1546
rect 110 1541 111 1545
rect 115 1541 116 1545
rect 110 1540 116 1541
rect 188 1532 190 1614
rect 214 1611 215 1615
rect 219 1611 220 1615
rect 214 1610 220 1611
rect 254 1615 260 1616
rect 254 1611 255 1615
rect 259 1611 260 1615
rect 266 1615 267 1619
rect 271 1615 272 1619
rect 312 1616 314 1625
rect 326 1619 332 1620
rect 266 1614 272 1615
rect 310 1615 316 1616
rect 254 1610 260 1611
rect 268 1588 270 1614
rect 310 1611 311 1615
rect 315 1611 316 1615
rect 326 1615 327 1619
rect 331 1615 332 1619
rect 392 1616 394 1625
rect 326 1614 332 1615
rect 390 1615 396 1616
rect 310 1610 316 1611
rect 328 1588 330 1614
rect 390 1611 391 1615
rect 395 1611 396 1615
rect 390 1610 396 1611
rect 408 1588 410 1638
rect 448 1631 450 1644
rect 496 1631 498 1644
rect 544 1631 546 1644
rect 566 1643 572 1644
rect 566 1639 567 1643
rect 571 1639 572 1643
rect 566 1638 572 1639
rect 592 1631 594 1644
rect 640 1631 642 1644
rect 688 1631 690 1644
rect 702 1643 708 1644
rect 702 1639 703 1643
rect 707 1639 708 1643
rect 702 1638 708 1639
rect 710 1643 716 1644
rect 710 1639 711 1643
rect 715 1639 716 1643
rect 710 1638 716 1639
rect 736 1631 738 1644
rect 750 1643 756 1644
rect 750 1639 751 1643
rect 755 1639 756 1643
rect 750 1638 756 1639
rect 784 1631 786 1644
rect 798 1643 804 1644
rect 798 1639 799 1643
rect 803 1639 804 1643
rect 798 1638 804 1639
rect 447 1630 451 1631
rect 447 1625 451 1626
rect 471 1630 475 1631
rect 471 1625 475 1626
rect 495 1630 499 1631
rect 495 1625 499 1626
rect 543 1630 547 1631
rect 543 1625 547 1626
rect 559 1630 563 1631
rect 559 1625 563 1626
rect 591 1630 595 1631
rect 591 1625 595 1626
rect 639 1630 643 1631
rect 639 1625 643 1626
rect 687 1630 691 1631
rect 687 1625 691 1626
rect 719 1630 723 1631
rect 719 1625 723 1626
rect 735 1630 739 1631
rect 735 1625 739 1626
rect 783 1630 787 1631
rect 783 1625 787 1626
rect 791 1630 795 1631
rect 791 1625 795 1626
rect 462 1619 468 1620
rect 462 1615 463 1619
rect 467 1615 468 1619
rect 472 1616 474 1625
rect 550 1619 556 1620
rect 462 1614 468 1615
rect 470 1615 476 1616
rect 464 1588 466 1614
rect 470 1611 471 1615
rect 475 1611 476 1615
rect 550 1615 551 1619
rect 555 1615 556 1619
rect 560 1616 562 1625
rect 570 1619 576 1620
rect 550 1614 556 1615
rect 558 1615 564 1616
rect 470 1610 476 1611
rect 552 1588 554 1614
rect 558 1611 559 1615
rect 563 1611 564 1615
rect 570 1615 571 1619
rect 575 1615 576 1619
rect 640 1616 642 1625
rect 710 1619 716 1620
rect 570 1614 576 1615
rect 638 1615 644 1616
rect 558 1610 564 1611
rect 572 1596 574 1614
rect 638 1611 639 1615
rect 643 1611 644 1615
rect 710 1615 711 1619
rect 715 1615 716 1619
rect 720 1616 722 1625
rect 782 1619 788 1620
rect 710 1614 716 1615
rect 718 1615 724 1616
rect 638 1610 644 1611
rect 570 1595 576 1596
rect 570 1591 571 1595
rect 575 1591 576 1595
rect 570 1590 576 1591
rect 712 1588 714 1614
rect 718 1611 719 1615
rect 723 1611 724 1615
rect 782 1615 783 1619
rect 787 1615 788 1619
rect 792 1616 794 1625
rect 820 1620 822 1670
rect 1238 1668 1239 1672
rect 1243 1668 1244 1672
rect 918 1667 924 1668
rect 1238 1667 1244 1668
rect 1278 1672 1284 1673
rect 1278 1668 1279 1672
rect 1283 1668 1284 1672
rect 1350 1671 1351 1675
rect 1355 1671 1356 1675
rect 1350 1670 1356 1671
rect 1278 1667 1284 1668
rect 918 1663 919 1667
rect 923 1663 924 1667
rect 918 1662 924 1663
rect 838 1649 844 1650
rect 838 1645 839 1649
rect 843 1645 844 1649
rect 838 1644 844 1645
rect 894 1649 900 1650
rect 894 1645 895 1649
rect 899 1645 900 1649
rect 894 1644 900 1645
rect 920 1644 922 1662
rect 840 1631 842 1644
rect 896 1631 898 1644
rect 918 1643 924 1644
rect 918 1639 919 1643
rect 923 1639 924 1643
rect 918 1638 924 1639
rect 1240 1631 1242 1667
rect 1280 1631 1282 1667
rect 1302 1649 1308 1650
rect 1302 1645 1303 1649
rect 1307 1645 1308 1649
rect 1302 1644 1308 1645
rect 1342 1649 1348 1650
rect 1342 1645 1343 1649
rect 1347 1645 1348 1649
rect 1342 1644 1348 1645
rect 1352 1644 1354 1670
rect 1368 1644 1370 1726
rect 1390 1712 1396 1713
rect 1390 1708 1391 1712
rect 1395 1708 1396 1712
rect 1390 1707 1396 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1518 1712 1524 1713
rect 1518 1708 1519 1712
rect 1523 1708 1524 1712
rect 1518 1707 1524 1708
rect 1582 1712 1588 1713
rect 1582 1708 1583 1712
rect 1587 1708 1588 1712
rect 1582 1707 1588 1708
rect 1392 1703 1394 1707
rect 1456 1703 1458 1707
rect 1520 1703 1522 1707
rect 1584 1703 1586 1707
rect 1383 1702 1387 1703
rect 1383 1697 1387 1698
rect 1391 1702 1395 1703
rect 1391 1697 1395 1698
rect 1423 1702 1427 1703
rect 1423 1697 1427 1698
rect 1455 1702 1459 1703
rect 1455 1697 1459 1698
rect 1463 1702 1467 1703
rect 1463 1697 1467 1698
rect 1503 1702 1507 1703
rect 1503 1697 1507 1698
rect 1519 1702 1523 1703
rect 1519 1697 1523 1698
rect 1559 1702 1563 1703
rect 1559 1697 1563 1698
rect 1583 1702 1587 1703
rect 1583 1697 1587 1698
rect 1382 1696 1388 1697
rect 1382 1692 1383 1696
rect 1387 1692 1388 1696
rect 1382 1691 1388 1692
rect 1422 1696 1428 1697
rect 1422 1692 1423 1696
rect 1427 1692 1428 1696
rect 1422 1691 1428 1692
rect 1462 1696 1468 1697
rect 1462 1692 1463 1696
rect 1467 1692 1468 1696
rect 1462 1691 1468 1692
rect 1502 1696 1508 1697
rect 1502 1692 1503 1696
rect 1507 1692 1508 1696
rect 1502 1691 1508 1692
rect 1558 1696 1564 1697
rect 1558 1692 1559 1696
rect 1563 1692 1564 1696
rect 1558 1691 1564 1692
rect 1596 1684 1598 1758
rect 1604 1740 1606 1790
rect 1616 1775 1618 1796
rect 1672 1775 1674 1796
rect 1728 1775 1730 1796
rect 1742 1795 1748 1796
rect 1742 1791 1743 1795
rect 1747 1791 1748 1795
rect 1742 1790 1748 1791
rect 1784 1775 1786 1796
rect 1798 1795 1804 1796
rect 1798 1791 1799 1795
rect 1803 1791 1804 1795
rect 1798 1790 1804 1791
rect 1840 1775 1842 1796
rect 1854 1795 1860 1796
rect 1854 1791 1855 1795
rect 1859 1791 1860 1795
rect 1854 1790 1860 1791
rect 1896 1775 1898 1796
rect 1615 1774 1619 1775
rect 1615 1769 1619 1770
rect 1647 1774 1651 1775
rect 1647 1769 1651 1770
rect 1671 1774 1675 1775
rect 1671 1769 1675 1770
rect 1703 1774 1707 1775
rect 1703 1769 1707 1770
rect 1727 1774 1731 1775
rect 1727 1769 1731 1770
rect 1759 1774 1763 1775
rect 1759 1769 1763 1770
rect 1783 1774 1787 1775
rect 1783 1769 1787 1770
rect 1807 1774 1811 1775
rect 1807 1769 1811 1770
rect 1839 1774 1843 1775
rect 1839 1769 1843 1770
rect 1863 1774 1867 1775
rect 1863 1769 1867 1770
rect 1895 1774 1899 1775
rect 1895 1769 1899 1770
rect 1648 1760 1650 1769
rect 1694 1763 1700 1764
rect 1646 1759 1652 1760
rect 1646 1755 1647 1759
rect 1651 1755 1652 1759
rect 1694 1759 1695 1763
rect 1699 1759 1700 1763
rect 1704 1760 1706 1769
rect 1750 1763 1756 1764
rect 1694 1758 1700 1759
rect 1702 1759 1708 1760
rect 1646 1754 1652 1755
rect 1674 1751 1680 1752
rect 1674 1747 1675 1751
rect 1679 1747 1680 1751
rect 1674 1746 1680 1747
rect 1602 1739 1608 1740
rect 1602 1735 1603 1739
rect 1607 1735 1608 1739
rect 1602 1734 1608 1735
rect 1676 1732 1678 1746
rect 1696 1732 1698 1758
rect 1702 1755 1703 1759
rect 1707 1755 1708 1759
rect 1750 1759 1751 1763
rect 1755 1759 1756 1763
rect 1760 1760 1762 1769
rect 1798 1763 1804 1764
rect 1750 1758 1756 1759
rect 1758 1759 1764 1760
rect 1702 1754 1708 1755
rect 1752 1732 1754 1758
rect 1758 1755 1759 1759
rect 1763 1755 1764 1759
rect 1798 1759 1799 1763
rect 1803 1759 1804 1763
rect 1808 1760 1810 1769
rect 1864 1760 1866 1769
rect 1904 1764 1906 1822
rect 2406 1820 2407 1824
rect 2411 1820 2412 1824
rect 1974 1819 1980 1820
rect 2406 1819 2412 1820
rect 1974 1815 1975 1819
rect 1979 1815 1980 1819
rect 1974 1814 1980 1815
rect 1950 1801 1956 1802
rect 1950 1797 1951 1801
rect 1955 1797 1956 1801
rect 1950 1796 1956 1797
rect 1976 1796 1978 1814
rect 1952 1775 1954 1796
rect 1974 1795 1980 1796
rect 1974 1791 1975 1795
rect 1979 1791 1980 1795
rect 1974 1790 1980 1791
rect 2408 1775 2410 1819
rect 1919 1774 1923 1775
rect 1919 1769 1923 1770
rect 1951 1774 1955 1775
rect 1951 1769 1955 1770
rect 1975 1774 1979 1775
rect 1975 1769 1979 1770
rect 2407 1774 2411 1775
rect 2407 1769 2411 1770
rect 1902 1763 1908 1764
rect 1798 1758 1804 1759
rect 1806 1759 1812 1760
rect 1758 1754 1764 1755
rect 1800 1740 1802 1758
rect 1806 1755 1807 1759
rect 1811 1755 1812 1759
rect 1806 1754 1812 1755
rect 1862 1759 1868 1760
rect 1862 1755 1863 1759
rect 1867 1755 1868 1759
rect 1902 1759 1903 1763
rect 1907 1759 1908 1763
rect 1920 1760 1922 1769
rect 1966 1763 1972 1764
rect 1902 1758 1908 1759
rect 1918 1759 1924 1760
rect 1862 1754 1868 1755
rect 1918 1755 1919 1759
rect 1923 1755 1924 1759
rect 1966 1759 1967 1763
rect 1971 1759 1972 1763
rect 1976 1760 1978 1769
rect 1966 1758 1972 1759
rect 1974 1759 1980 1760
rect 1918 1754 1924 1755
rect 1830 1751 1836 1752
rect 1830 1747 1831 1751
rect 1835 1747 1836 1751
rect 1830 1746 1836 1747
rect 1798 1739 1804 1740
rect 1798 1735 1799 1739
rect 1803 1735 1804 1739
rect 1798 1734 1804 1735
rect 1832 1732 1834 1746
rect 1968 1732 1970 1758
rect 1974 1755 1975 1759
rect 1979 1755 1980 1759
rect 1974 1754 1980 1755
rect 2408 1737 2410 1769
rect 2406 1736 2412 1737
rect 2406 1732 2407 1736
rect 2411 1732 2412 1736
rect 1674 1731 1680 1732
rect 1674 1727 1675 1731
rect 1679 1727 1680 1731
rect 1674 1726 1680 1727
rect 1694 1731 1700 1732
rect 1694 1727 1695 1731
rect 1699 1727 1700 1731
rect 1694 1726 1700 1727
rect 1750 1731 1756 1732
rect 1750 1727 1751 1731
rect 1755 1727 1756 1731
rect 1750 1726 1756 1727
rect 1830 1731 1836 1732
rect 1830 1727 1831 1731
rect 1835 1727 1836 1731
rect 1830 1726 1836 1727
rect 1966 1731 1972 1732
rect 2406 1731 2412 1732
rect 1966 1727 1967 1731
rect 1971 1727 1972 1731
rect 1966 1726 1972 1727
rect 2406 1719 2412 1720
rect 2406 1715 2407 1719
rect 2411 1715 2412 1719
rect 2406 1714 2412 1715
rect 1646 1712 1652 1713
rect 1646 1708 1647 1712
rect 1651 1708 1652 1712
rect 1646 1707 1652 1708
rect 1702 1712 1708 1713
rect 1702 1708 1703 1712
rect 1707 1708 1708 1712
rect 1702 1707 1708 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1806 1712 1812 1713
rect 1806 1708 1807 1712
rect 1811 1708 1812 1712
rect 1806 1707 1812 1708
rect 1862 1712 1868 1713
rect 1862 1708 1863 1712
rect 1867 1708 1868 1712
rect 1862 1707 1868 1708
rect 1918 1712 1924 1713
rect 1918 1708 1919 1712
rect 1923 1708 1924 1712
rect 1918 1707 1924 1708
rect 1974 1712 1980 1713
rect 1974 1708 1975 1712
rect 1979 1708 1980 1712
rect 1974 1707 1980 1708
rect 1648 1703 1650 1707
rect 1704 1703 1706 1707
rect 1760 1703 1762 1707
rect 1808 1703 1810 1707
rect 1864 1703 1866 1707
rect 1920 1703 1922 1707
rect 1976 1703 1978 1707
rect 2408 1703 2410 1714
rect 1623 1702 1627 1703
rect 1623 1697 1627 1698
rect 1647 1702 1651 1703
rect 1647 1697 1651 1698
rect 1687 1702 1691 1703
rect 1687 1697 1691 1698
rect 1703 1702 1707 1703
rect 1703 1697 1707 1698
rect 1751 1702 1755 1703
rect 1751 1697 1755 1698
rect 1759 1702 1763 1703
rect 1759 1697 1763 1698
rect 1807 1702 1811 1703
rect 1807 1697 1811 1698
rect 1863 1702 1867 1703
rect 1863 1697 1867 1698
rect 1919 1702 1923 1703
rect 1919 1697 1923 1698
rect 1975 1702 1979 1703
rect 1975 1697 1979 1698
rect 2031 1702 2035 1703
rect 2031 1697 2035 1698
rect 2087 1702 2091 1703
rect 2087 1697 2091 1698
rect 2407 1702 2411 1703
rect 2407 1697 2411 1698
rect 1622 1696 1628 1697
rect 1622 1692 1623 1696
rect 1627 1692 1628 1696
rect 1622 1691 1628 1692
rect 1686 1696 1692 1697
rect 1686 1692 1687 1696
rect 1691 1692 1692 1696
rect 1686 1691 1692 1692
rect 1750 1696 1756 1697
rect 1750 1692 1751 1696
rect 1755 1692 1756 1696
rect 1750 1691 1756 1692
rect 1806 1696 1812 1697
rect 1806 1692 1807 1696
rect 1811 1692 1812 1696
rect 1806 1691 1812 1692
rect 1862 1696 1868 1697
rect 1862 1692 1863 1696
rect 1867 1692 1868 1696
rect 1862 1691 1868 1692
rect 1918 1696 1924 1697
rect 1918 1692 1919 1696
rect 1923 1692 1924 1696
rect 1918 1691 1924 1692
rect 1974 1696 1980 1697
rect 1974 1692 1975 1696
rect 1979 1692 1980 1696
rect 1974 1691 1980 1692
rect 2030 1696 2036 1697
rect 2030 1692 2031 1696
rect 2035 1692 2036 1696
rect 2030 1691 2036 1692
rect 2086 1696 2092 1697
rect 2086 1692 2087 1696
rect 2091 1692 2092 1696
rect 2086 1691 2092 1692
rect 2408 1690 2410 1697
rect 2406 1689 2412 1690
rect 2406 1685 2407 1689
rect 2411 1685 2412 1689
rect 2406 1684 2412 1685
rect 1594 1683 1600 1684
rect 1594 1679 1595 1683
rect 1599 1679 1600 1683
rect 1594 1678 1600 1679
rect 2110 1683 2116 1684
rect 2110 1679 2111 1683
rect 2115 1679 2116 1683
rect 2110 1678 2116 1679
rect 1430 1675 1436 1676
rect 1430 1671 1431 1675
rect 1435 1671 1436 1675
rect 1430 1670 1436 1671
rect 1470 1675 1476 1676
rect 1470 1671 1471 1675
rect 1475 1671 1476 1675
rect 1470 1670 1476 1671
rect 1786 1675 1792 1676
rect 1786 1671 1787 1675
rect 1791 1671 1792 1675
rect 1786 1670 1792 1671
rect 1954 1675 1960 1676
rect 1954 1671 1955 1675
rect 1959 1671 1960 1675
rect 1954 1670 1960 1671
rect 1406 1667 1412 1668
rect 1406 1663 1407 1667
rect 1411 1663 1412 1667
rect 1406 1662 1412 1663
rect 1382 1649 1388 1650
rect 1382 1645 1383 1649
rect 1387 1645 1388 1649
rect 1382 1644 1388 1645
rect 1408 1644 1410 1662
rect 1422 1649 1428 1650
rect 1422 1645 1423 1649
rect 1427 1645 1428 1649
rect 1422 1644 1428 1645
rect 1304 1631 1306 1644
rect 1344 1631 1346 1644
rect 1350 1643 1356 1644
rect 1350 1639 1351 1643
rect 1355 1639 1356 1643
rect 1350 1638 1356 1639
rect 1366 1643 1372 1644
rect 1366 1639 1367 1643
rect 1371 1639 1372 1643
rect 1366 1638 1372 1639
rect 1384 1631 1386 1644
rect 1406 1643 1412 1644
rect 1406 1639 1407 1643
rect 1411 1639 1412 1643
rect 1406 1638 1412 1639
rect 1424 1631 1426 1644
rect 839 1630 843 1631
rect 839 1625 843 1626
rect 855 1630 859 1631
rect 855 1625 859 1626
rect 895 1630 899 1631
rect 895 1625 899 1626
rect 919 1630 923 1631
rect 919 1625 923 1626
rect 983 1630 987 1631
rect 983 1625 987 1626
rect 1047 1630 1051 1631
rect 1047 1625 1051 1626
rect 1239 1630 1243 1631
rect 1239 1625 1243 1626
rect 1279 1630 1283 1631
rect 1279 1625 1283 1626
rect 1303 1630 1307 1631
rect 1303 1625 1307 1626
rect 1343 1630 1347 1631
rect 1343 1625 1347 1626
rect 1383 1630 1387 1631
rect 1383 1625 1387 1626
rect 1423 1630 1427 1631
rect 1423 1625 1427 1626
rect 818 1619 824 1620
rect 782 1614 788 1615
rect 790 1615 796 1616
rect 718 1610 724 1611
rect 784 1588 786 1614
rect 790 1611 791 1615
rect 795 1611 796 1615
rect 818 1615 819 1619
rect 823 1615 824 1619
rect 856 1616 858 1625
rect 866 1619 872 1620
rect 818 1614 824 1615
rect 854 1615 860 1616
rect 790 1610 796 1611
rect 854 1611 855 1615
rect 859 1611 860 1615
rect 866 1615 867 1619
rect 871 1615 872 1619
rect 920 1616 922 1625
rect 974 1619 980 1620
rect 866 1614 872 1615
rect 918 1615 924 1616
rect 854 1610 860 1611
rect 868 1596 870 1614
rect 918 1611 919 1615
rect 923 1611 924 1615
rect 974 1615 975 1619
rect 979 1615 980 1619
rect 984 1616 986 1625
rect 1038 1619 1044 1620
rect 974 1614 980 1615
rect 982 1615 988 1616
rect 918 1610 924 1611
rect 866 1595 872 1596
rect 866 1591 867 1595
rect 871 1591 872 1595
rect 866 1590 872 1591
rect 976 1588 978 1614
rect 982 1611 983 1615
rect 987 1611 988 1615
rect 1038 1615 1039 1619
rect 1043 1615 1044 1619
rect 1048 1616 1050 1625
rect 1058 1619 1064 1620
rect 1038 1614 1044 1615
rect 1046 1615 1052 1616
rect 982 1610 988 1611
rect 1040 1588 1042 1614
rect 1046 1611 1047 1615
rect 1051 1611 1052 1615
rect 1058 1615 1059 1619
rect 1063 1615 1064 1619
rect 1058 1614 1064 1615
rect 1046 1610 1052 1611
rect 1060 1596 1062 1614
rect 1058 1595 1064 1596
rect 1058 1591 1059 1595
rect 1063 1591 1064 1595
rect 1240 1593 1242 1625
rect 1280 1593 1282 1625
rect 1304 1616 1306 1625
rect 1344 1616 1346 1625
rect 1358 1623 1364 1624
rect 1358 1619 1359 1623
rect 1363 1619 1364 1623
rect 1358 1618 1364 1619
rect 1302 1615 1308 1616
rect 1302 1611 1303 1615
rect 1307 1611 1308 1615
rect 1302 1610 1308 1611
rect 1342 1615 1348 1616
rect 1342 1611 1343 1615
rect 1347 1611 1348 1615
rect 1342 1610 1348 1611
rect 1058 1590 1064 1591
rect 1238 1592 1244 1593
rect 1238 1588 1239 1592
rect 1243 1588 1244 1592
rect 266 1587 272 1588
rect 266 1583 267 1587
rect 271 1583 272 1587
rect 266 1582 272 1583
rect 326 1587 332 1588
rect 326 1583 327 1587
rect 331 1583 332 1587
rect 326 1582 332 1583
rect 406 1587 412 1588
rect 406 1583 407 1587
rect 411 1583 412 1587
rect 406 1582 412 1583
rect 462 1587 468 1588
rect 462 1583 463 1587
rect 467 1583 468 1587
rect 462 1582 468 1583
rect 550 1587 556 1588
rect 550 1583 551 1587
rect 555 1583 556 1587
rect 550 1582 556 1583
rect 710 1587 716 1588
rect 710 1583 711 1587
rect 715 1583 716 1587
rect 710 1582 716 1583
rect 782 1587 788 1588
rect 782 1583 783 1587
rect 787 1583 788 1587
rect 782 1582 788 1583
rect 930 1587 936 1588
rect 930 1583 931 1587
rect 935 1583 936 1587
rect 930 1582 936 1583
rect 974 1587 980 1588
rect 974 1583 975 1587
rect 979 1583 980 1587
rect 974 1582 980 1583
rect 1038 1587 1044 1588
rect 1238 1587 1244 1588
rect 1278 1592 1284 1593
rect 1278 1588 1279 1592
rect 1283 1588 1284 1592
rect 1360 1588 1362 1618
rect 1384 1616 1386 1625
rect 1398 1623 1404 1624
rect 1398 1619 1399 1623
rect 1403 1619 1404 1623
rect 1398 1618 1404 1619
rect 1382 1615 1388 1616
rect 1382 1611 1383 1615
rect 1387 1611 1388 1615
rect 1382 1610 1388 1611
rect 1400 1588 1402 1618
rect 1424 1616 1426 1625
rect 1432 1624 1434 1670
rect 1462 1649 1468 1650
rect 1462 1645 1463 1649
rect 1467 1645 1468 1649
rect 1462 1644 1468 1645
rect 1472 1644 1474 1670
rect 1486 1667 1492 1668
rect 1486 1663 1487 1667
rect 1491 1663 1492 1667
rect 1486 1662 1492 1663
rect 1488 1644 1490 1662
rect 1502 1649 1508 1650
rect 1502 1645 1503 1649
rect 1507 1645 1508 1649
rect 1502 1644 1508 1645
rect 1558 1649 1564 1650
rect 1558 1645 1559 1649
rect 1563 1645 1564 1649
rect 1558 1644 1564 1645
rect 1622 1649 1628 1650
rect 1622 1645 1623 1649
rect 1627 1645 1628 1649
rect 1622 1644 1628 1645
rect 1686 1649 1692 1650
rect 1686 1645 1687 1649
rect 1691 1645 1692 1649
rect 1686 1644 1692 1645
rect 1750 1649 1756 1650
rect 1750 1645 1751 1649
rect 1755 1645 1756 1649
rect 1750 1644 1756 1645
rect 1788 1644 1790 1670
rect 1942 1667 1948 1668
rect 1942 1663 1943 1667
rect 1947 1663 1948 1667
rect 1942 1662 1948 1663
rect 1806 1649 1812 1650
rect 1806 1645 1807 1649
rect 1811 1645 1812 1649
rect 1806 1644 1812 1645
rect 1862 1649 1868 1650
rect 1862 1645 1863 1649
rect 1867 1645 1868 1649
rect 1862 1644 1868 1645
rect 1918 1649 1924 1650
rect 1918 1645 1919 1649
rect 1923 1645 1924 1649
rect 1918 1644 1924 1645
rect 1944 1644 1946 1662
rect 1464 1631 1466 1644
rect 1470 1643 1476 1644
rect 1470 1639 1471 1643
rect 1475 1639 1476 1643
rect 1470 1638 1476 1639
rect 1486 1643 1492 1644
rect 1486 1639 1487 1643
rect 1491 1639 1492 1643
rect 1486 1638 1492 1639
rect 1504 1631 1506 1644
rect 1560 1631 1562 1644
rect 1624 1631 1626 1644
rect 1688 1631 1690 1644
rect 1752 1631 1754 1644
rect 1786 1643 1792 1644
rect 1786 1639 1787 1643
rect 1791 1639 1792 1643
rect 1786 1638 1792 1639
rect 1808 1631 1810 1644
rect 1864 1631 1866 1644
rect 1920 1631 1922 1644
rect 1942 1643 1948 1644
rect 1942 1639 1943 1643
rect 1947 1639 1948 1643
rect 1942 1638 1948 1639
rect 1463 1630 1467 1631
rect 1463 1625 1467 1626
rect 1503 1630 1507 1631
rect 1503 1625 1507 1626
rect 1559 1630 1563 1631
rect 1559 1625 1563 1626
rect 1623 1630 1627 1631
rect 1623 1625 1627 1626
rect 1631 1630 1635 1631
rect 1631 1625 1635 1626
rect 1687 1630 1691 1631
rect 1687 1625 1691 1626
rect 1703 1630 1707 1631
rect 1703 1625 1707 1626
rect 1751 1630 1755 1631
rect 1751 1625 1755 1626
rect 1783 1630 1787 1631
rect 1783 1625 1787 1626
rect 1807 1630 1811 1631
rect 1807 1625 1811 1626
rect 1855 1630 1859 1631
rect 1855 1625 1859 1626
rect 1863 1630 1867 1631
rect 1863 1625 1867 1626
rect 1919 1630 1923 1631
rect 1919 1625 1923 1626
rect 1927 1630 1931 1631
rect 1927 1625 1931 1626
rect 1430 1623 1436 1624
rect 1430 1619 1431 1623
rect 1435 1619 1436 1623
rect 1430 1618 1436 1619
rect 1438 1619 1444 1620
rect 1422 1615 1428 1616
rect 1422 1611 1423 1615
rect 1427 1611 1428 1615
rect 1438 1615 1439 1619
rect 1443 1615 1444 1619
rect 1464 1616 1466 1625
rect 1474 1619 1480 1620
rect 1438 1614 1444 1615
rect 1462 1615 1468 1616
rect 1422 1610 1428 1611
rect 1440 1596 1442 1614
rect 1462 1611 1463 1615
rect 1467 1611 1468 1615
rect 1474 1615 1475 1619
rect 1479 1615 1480 1619
rect 1504 1616 1506 1625
rect 1514 1619 1520 1620
rect 1474 1614 1480 1615
rect 1502 1615 1508 1616
rect 1462 1610 1468 1611
rect 1438 1595 1444 1596
rect 1438 1591 1439 1595
rect 1443 1591 1444 1595
rect 1438 1590 1444 1591
rect 1476 1588 1478 1614
rect 1502 1611 1503 1615
rect 1507 1611 1508 1615
rect 1514 1615 1515 1619
rect 1519 1615 1520 1619
rect 1560 1616 1562 1625
rect 1622 1619 1628 1620
rect 1514 1614 1520 1615
rect 1558 1615 1564 1616
rect 1502 1610 1508 1611
rect 1516 1596 1518 1614
rect 1558 1611 1559 1615
rect 1563 1611 1564 1615
rect 1622 1615 1623 1619
rect 1627 1615 1628 1619
rect 1632 1616 1634 1625
rect 1694 1619 1700 1620
rect 1622 1614 1628 1615
rect 1630 1615 1636 1616
rect 1558 1610 1564 1611
rect 1514 1595 1520 1596
rect 1514 1591 1515 1595
rect 1519 1591 1520 1595
rect 1514 1590 1520 1591
rect 1624 1588 1626 1614
rect 1630 1611 1631 1615
rect 1635 1611 1636 1615
rect 1694 1615 1695 1619
rect 1699 1615 1700 1619
rect 1704 1616 1706 1625
rect 1774 1619 1780 1620
rect 1694 1614 1700 1615
rect 1702 1615 1708 1616
rect 1630 1610 1636 1611
rect 1696 1588 1698 1614
rect 1702 1611 1703 1615
rect 1707 1611 1708 1615
rect 1774 1615 1775 1619
rect 1779 1615 1780 1619
rect 1784 1616 1786 1625
rect 1794 1619 1800 1620
rect 1774 1614 1780 1615
rect 1782 1615 1788 1616
rect 1702 1610 1708 1611
rect 1776 1588 1778 1614
rect 1782 1611 1783 1615
rect 1787 1611 1788 1615
rect 1794 1615 1795 1619
rect 1799 1615 1800 1619
rect 1856 1616 1858 1625
rect 1918 1619 1924 1620
rect 1794 1614 1800 1615
rect 1854 1615 1860 1616
rect 1782 1610 1788 1611
rect 1278 1587 1284 1588
rect 1358 1587 1364 1588
rect 1038 1583 1039 1587
rect 1043 1583 1044 1587
rect 1038 1582 1044 1583
rect 1358 1583 1359 1587
rect 1363 1583 1364 1587
rect 1358 1582 1364 1583
rect 1398 1587 1404 1588
rect 1398 1583 1399 1587
rect 1403 1583 1404 1587
rect 1398 1582 1404 1583
rect 1474 1587 1480 1588
rect 1474 1583 1475 1587
rect 1479 1583 1480 1587
rect 1474 1582 1480 1583
rect 1510 1587 1516 1588
rect 1510 1583 1511 1587
rect 1515 1583 1516 1587
rect 1510 1582 1516 1583
rect 1622 1587 1628 1588
rect 1622 1583 1623 1587
rect 1627 1583 1628 1587
rect 1622 1582 1628 1583
rect 1694 1587 1700 1588
rect 1694 1583 1695 1587
rect 1699 1583 1700 1587
rect 1694 1582 1700 1583
rect 1774 1587 1780 1588
rect 1774 1583 1775 1587
rect 1779 1583 1780 1587
rect 1774 1582 1780 1583
rect 214 1568 220 1569
rect 214 1564 215 1568
rect 219 1564 220 1568
rect 214 1563 220 1564
rect 254 1568 260 1569
rect 254 1564 255 1568
rect 259 1564 260 1568
rect 254 1563 260 1564
rect 310 1568 316 1569
rect 310 1564 311 1568
rect 315 1564 316 1568
rect 310 1563 316 1564
rect 390 1568 396 1569
rect 390 1564 391 1568
rect 395 1564 396 1568
rect 390 1563 396 1564
rect 470 1568 476 1569
rect 470 1564 471 1568
rect 475 1564 476 1568
rect 470 1563 476 1564
rect 558 1568 564 1569
rect 558 1564 559 1568
rect 563 1564 564 1568
rect 558 1563 564 1564
rect 638 1568 644 1569
rect 638 1564 639 1568
rect 643 1564 644 1568
rect 638 1563 644 1564
rect 718 1568 724 1569
rect 718 1564 719 1568
rect 723 1564 724 1568
rect 718 1563 724 1564
rect 790 1568 796 1569
rect 790 1564 791 1568
rect 795 1564 796 1568
rect 790 1563 796 1564
rect 854 1568 860 1569
rect 854 1564 855 1568
rect 859 1564 860 1568
rect 854 1563 860 1564
rect 918 1568 924 1569
rect 918 1564 919 1568
rect 923 1564 924 1568
rect 918 1563 924 1564
rect 216 1559 218 1563
rect 256 1559 258 1563
rect 312 1559 314 1563
rect 392 1559 394 1563
rect 472 1559 474 1563
rect 560 1559 562 1563
rect 640 1559 642 1563
rect 720 1559 722 1563
rect 792 1559 794 1563
rect 856 1559 858 1563
rect 920 1559 922 1563
rect 199 1558 203 1559
rect 199 1553 203 1554
rect 215 1558 219 1559
rect 215 1553 219 1554
rect 255 1558 259 1559
rect 255 1553 259 1554
rect 263 1558 267 1559
rect 263 1553 267 1554
rect 311 1558 315 1559
rect 311 1553 315 1554
rect 343 1558 347 1559
rect 343 1553 347 1554
rect 391 1558 395 1559
rect 391 1553 395 1554
rect 439 1558 443 1559
rect 439 1553 443 1554
rect 471 1558 475 1559
rect 471 1553 475 1554
rect 535 1558 539 1559
rect 535 1553 539 1554
rect 559 1558 563 1559
rect 559 1553 563 1554
rect 639 1558 643 1559
rect 639 1553 643 1554
rect 719 1558 723 1559
rect 719 1553 723 1554
rect 735 1558 739 1559
rect 735 1553 739 1554
rect 791 1558 795 1559
rect 791 1553 795 1554
rect 823 1558 827 1559
rect 823 1553 827 1554
rect 855 1558 859 1559
rect 855 1553 859 1554
rect 903 1558 907 1559
rect 903 1553 907 1554
rect 919 1558 923 1559
rect 919 1553 923 1554
rect 198 1552 204 1553
rect 198 1548 199 1552
rect 203 1548 204 1552
rect 198 1547 204 1548
rect 262 1552 268 1553
rect 262 1548 263 1552
rect 267 1548 268 1552
rect 262 1547 268 1548
rect 342 1552 348 1553
rect 342 1548 343 1552
rect 347 1548 348 1552
rect 342 1547 348 1548
rect 438 1552 444 1553
rect 438 1548 439 1552
rect 443 1548 444 1552
rect 438 1547 444 1548
rect 534 1552 540 1553
rect 534 1548 535 1552
rect 539 1548 540 1552
rect 534 1547 540 1548
rect 638 1552 644 1553
rect 638 1548 639 1552
rect 643 1548 644 1552
rect 638 1547 644 1548
rect 734 1552 740 1553
rect 734 1548 735 1552
rect 739 1548 740 1552
rect 734 1547 740 1548
rect 822 1552 828 1553
rect 822 1548 823 1552
rect 827 1548 828 1552
rect 822 1547 828 1548
rect 902 1552 908 1553
rect 902 1548 903 1552
rect 907 1548 908 1552
rect 902 1547 908 1548
rect 186 1531 192 1532
rect 110 1528 116 1529
rect 110 1524 111 1528
rect 115 1524 116 1528
rect 186 1527 187 1531
rect 191 1527 192 1531
rect 186 1526 192 1527
rect 206 1531 212 1532
rect 206 1527 207 1531
rect 211 1527 212 1531
rect 206 1526 212 1527
rect 110 1523 116 1524
rect 112 1487 114 1523
rect 150 1505 156 1506
rect 150 1501 151 1505
rect 155 1501 156 1505
rect 150 1500 156 1501
rect 198 1505 204 1506
rect 198 1501 199 1505
rect 203 1501 204 1505
rect 198 1500 204 1501
rect 208 1500 210 1526
rect 262 1505 268 1506
rect 262 1501 263 1505
rect 267 1501 268 1505
rect 262 1500 268 1501
rect 342 1505 348 1506
rect 342 1501 343 1505
rect 347 1501 348 1505
rect 342 1500 348 1501
rect 438 1505 444 1506
rect 438 1501 439 1505
rect 443 1501 444 1505
rect 438 1500 444 1501
rect 534 1505 540 1506
rect 534 1501 535 1505
rect 539 1501 540 1505
rect 534 1500 540 1501
rect 638 1505 644 1506
rect 638 1501 639 1505
rect 643 1501 644 1505
rect 638 1500 644 1501
rect 734 1505 740 1506
rect 734 1501 735 1505
rect 739 1501 740 1505
rect 734 1500 740 1501
rect 822 1505 828 1506
rect 822 1501 823 1505
rect 827 1501 828 1505
rect 822 1500 828 1501
rect 902 1505 908 1506
rect 902 1501 903 1505
rect 907 1501 908 1505
rect 902 1500 908 1501
rect 932 1500 934 1582
rect 1238 1575 1244 1576
rect 1238 1571 1239 1575
rect 1243 1571 1244 1575
rect 1238 1570 1244 1571
rect 1278 1575 1284 1576
rect 1278 1571 1279 1575
rect 1283 1571 1284 1575
rect 1278 1570 1284 1571
rect 982 1568 988 1569
rect 982 1564 983 1568
rect 987 1564 988 1568
rect 982 1563 988 1564
rect 1046 1568 1052 1569
rect 1046 1564 1047 1568
rect 1051 1564 1052 1568
rect 1046 1563 1052 1564
rect 984 1559 986 1563
rect 1048 1559 1050 1563
rect 1240 1559 1242 1570
rect 1280 1563 1282 1570
rect 1302 1568 1308 1569
rect 1302 1564 1303 1568
rect 1307 1564 1308 1568
rect 1302 1563 1308 1564
rect 1342 1568 1348 1569
rect 1342 1564 1343 1568
rect 1347 1564 1348 1568
rect 1342 1563 1348 1564
rect 1382 1568 1388 1569
rect 1382 1564 1383 1568
rect 1387 1564 1388 1568
rect 1382 1563 1388 1564
rect 1422 1568 1428 1569
rect 1422 1564 1423 1568
rect 1427 1564 1428 1568
rect 1422 1563 1428 1564
rect 1462 1568 1468 1569
rect 1462 1564 1463 1568
rect 1467 1564 1468 1568
rect 1462 1563 1468 1564
rect 1502 1568 1508 1569
rect 1502 1564 1503 1568
rect 1507 1564 1508 1568
rect 1502 1563 1508 1564
rect 1279 1562 1283 1563
rect 975 1558 979 1559
rect 975 1553 979 1554
rect 983 1558 987 1559
rect 983 1553 987 1554
rect 1047 1558 1051 1559
rect 1047 1553 1051 1554
rect 1119 1558 1123 1559
rect 1119 1553 1123 1554
rect 1191 1558 1195 1559
rect 1191 1553 1195 1554
rect 1239 1558 1243 1559
rect 1279 1557 1283 1558
rect 1303 1562 1307 1563
rect 1303 1557 1307 1558
rect 1343 1562 1347 1563
rect 1343 1557 1347 1558
rect 1383 1562 1387 1563
rect 1383 1557 1387 1558
rect 1423 1562 1427 1563
rect 1423 1557 1427 1558
rect 1463 1562 1467 1563
rect 1463 1557 1467 1558
rect 1471 1562 1475 1563
rect 1471 1557 1475 1558
rect 1503 1562 1507 1563
rect 1503 1557 1507 1558
rect 1239 1553 1243 1554
rect 974 1552 980 1553
rect 974 1548 975 1552
rect 979 1548 980 1552
rect 974 1547 980 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1118 1552 1124 1553
rect 1118 1548 1119 1552
rect 1123 1548 1124 1552
rect 1118 1547 1124 1548
rect 1190 1552 1196 1553
rect 1190 1548 1191 1552
rect 1195 1548 1196 1552
rect 1190 1547 1196 1548
rect 1240 1546 1242 1553
rect 1280 1550 1282 1557
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1278 1549 1284 1550
rect 1238 1545 1244 1546
rect 1238 1541 1239 1545
rect 1243 1541 1244 1545
rect 1278 1545 1279 1549
rect 1283 1545 1284 1549
rect 1278 1544 1284 1545
rect 1238 1540 1244 1541
rect 1278 1532 1284 1533
rect 1062 1531 1068 1532
rect 1062 1527 1063 1531
rect 1067 1527 1068 1531
rect 1062 1526 1068 1527
rect 1134 1531 1140 1532
rect 1134 1527 1135 1531
rect 1139 1527 1140 1531
rect 1134 1526 1140 1527
rect 1206 1531 1212 1532
rect 1206 1527 1207 1531
rect 1211 1527 1212 1531
rect 1206 1526 1212 1527
rect 1238 1528 1244 1529
rect 998 1523 1004 1524
rect 998 1519 999 1523
rect 1003 1519 1004 1523
rect 998 1518 1004 1519
rect 974 1505 980 1506
rect 974 1501 975 1505
rect 979 1501 980 1505
rect 974 1500 980 1501
rect 1000 1500 1002 1518
rect 1046 1505 1052 1506
rect 1046 1501 1047 1505
rect 1051 1501 1052 1505
rect 1046 1500 1052 1501
rect 1064 1500 1066 1526
rect 1118 1505 1124 1506
rect 1118 1501 1119 1505
rect 1123 1501 1124 1505
rect 1118 1500 1124 1501
rect 1136 1500 1138 1526
rect 1178 1523 1184 1524
rect 1178 1519 1179 1523
rect 1183 1519 1184 1523
rect 1178 1518 1184 1519
rect 152 1487 154 1500
rect 200 1487 202 1500
rect 206 1499 212 1500
rect 206 1495 207 1499
rect 211 1495 212 1499
rect 206 1494 212 1495
rect 264 1487 266 1500
rect 344 1487 346 1500
rect 440 1487 442 1500
rect 536 1487 538 1500
rect 578 1499 584 1500
rect 578 1495 579 1499
rect 583 1495 584 1499
rect 578 1494 584 1495
rect 111 1486 115 1487
rect 111 1481 115 1482
rect 151 1486 155 1487
rect 151 1481 155 1482
rect 199 1486 203 1487
rect 199 1481 203 1482
rect 263 1486 267 1487
rect 263 1481 267 1482
rect 319 1486 323 1487
rect 319 1481 323 1482
rect 343 1486 347 1487
rect 343 1481 347 1482
rect 359 1486 363 1487
rect 359 1481 363 1482
rect 399 1486 403 1487
rect 399 1481 403 1482
rect 439 1486 443 1487
rect 439 1481 443 1482
rect 447 1486 451 1487
rect 447 1481 451 1482
rect 503 1486 507 1487
rect 503 1481 507 1482
rect 535 1486 539 1487
rect 535 1481 539 1482
rect 559 1486 563 1487
rect 559 1481 563 1482
rect 112 1449 114 1481
rect 320 1472 322 1481
rect 346 1475 352 1476
rect 318 1471 324 1472
rect 318 1467 319 1471
rect 323 1467 324 1471
rect 346 1471 347 1475
rect 351 1471 352 1475
rect 360 1472 362 1481
rect 400 1472 402 1481
rect 414 1479 420 1480
rect 414 1475 415 1479
rect 419 1475 420 1479
rect 414 1474 420 1475
rect 438 1475 444 1476
rect 346 1470 352 1471
rect 358 1471 364 1472
rect 318 1466 324 1467
rect 348 1452 350 1470
rect 358 1467 359 1471
rect 363 1467 364 1471
rect 358 1466 364 1467
rect 398 1471 404 1472
rect 398 1467 399 1471
rect 403 1467 404 1471
rect 398 1466 404 1467
rect 346 1451 352 1452
rect 110 1448 116 1449
rect 110 1444 111 1448
rect 115 1444 116 1448
rect 346 1447 347 1451
rect 351 1447 352 1451
rect 346 1446 352 1447
rect 416 1444 418 1474
rect 438 1471 439 1475
rect 443 1471 444 1475
rect 448 1472 450 1481
rect 494 1475 500 1476
rect 438 1470 444 1471
rect 446 1471 452 1472
rect 440 1444 442 1470
rect 446 1467 447 1471
rect 451 1467 452 1471
rect 494 1471 495 1475
rect 499 1471 500 1475
rect 504 1472 506 1481
rect 550 1475 556 1476
rect 494 1470 500 1471
rect 502 1471 508 1472
rect 446 1466 452 1467
rect 496 1444 498 1470
rect 502 1467 503 1471
rect 507 1467 508 1471
rect 550 1471 551 1475
rect 555 1471 556 1475
rect 560 1472 562 1481
rect 550 1470 556 1471
rect 558 1471 564 1472
rect 502 1466 508 1467
rect 552 1444 554 1470
rect 558 1467 559 1471
rect 563 1467 564 1471
rect 558 1466 564 1467
rect 110 1443 116 1444
rect 414 1443 420 1444
rect 414 1439 415 1443
rect 419 1439 420 1443
rect 414 1438 420 1439
rect 438 1443 444 1444
rect 438 1439 439 1443
rect 443 1439 444 1443
rect 438 1438 444 1439
rect 494 1443 500 1444
rect 494 1439 495 1443
rect 499 1439 500 1443
rect 494 1438 500 1439
rect 550 1443 556 1444
rect 550 1439 551 1443
rect 555 1439 556 1443
rect 550 1438 556 1439
rect 580 1436 582 1494
rect 640 1487 642 1500
rect 736 1487 738 1500
rect 824 1487 826 1500
rect 904 1487 906 1500
rect 930 1499 936 1500
rect 930 1495 931 1499
rect 935 1495 936 1499
rect 930 1494 936 1495
rect 976 1487 978 1500
rect 998 1499 1004 1500
rect 998 1495 999 1499
rect 1003 1495 1004 1499
rect 998 1494 1004 1495
rect 1048 1487 1050 1500
rect 1062 1499 1068 1500
rect 1062 1495 1063 1499
rect 1067 1495 1068 1499
rect 1062 1494 1068 1495
rect 1120 1487 1122 1500
rect 1134 1499 1140 1500
rect 1134 1495 1135 1499
rect 1139 1495 1140 1499
rect 1134 1494 1140 1495
rect 615 1486 619 1487
rect 615 1481 619 1482
rect 639 1486 643 1487
rect 639 1481 643 1482
rect 671 1486 675 1487
rect 671 1481 675 1482
rect 735 1486 739 1487
rect 735 1481 739 1482
rect 799 1486 803 1487
rect 799 1481 803 1482
rect 823 1486 827 1487
rect 823 1481 827 1482
rect 855 1486 859 1487
rect 855 1481 859 1482
rect 903 1486 907 1487
rect 903 1481 907 1482
rect 911 1486 915 1487
rect 911 1481 915 1482
rect 967 1486 971 1487
rect 967 1481 971 1482
rect 975 1486 979 1487
rect 975 1481 979 1482
rect 1023 1486 1027 1487
rect 1023 1481 1027 1482
rect 1047 1486 1051 1487
rect 1047 1481 1051 1482
rect 1087 1486 1091 1487
rect 1087 1481 1091 1482
rect 1119 1486 1123 1487
rect 1119 1481 1123 1482
rect 1151 1486 1155 1487
rect 1151 1481 1155 1482
rect 606 1475 612 1476
rect 606 1471 607 1475
rect 611 1471 612 1475
rect 616 1472 618 1481
rect 630 1475 636 1476
rect 606 1470 612 1471
rect 614 1471 620 1472
rect 608 1444 610 1470
rect 614 1467 615 1471
rect 619 1467 620 1471
rect 630 1471 631 1475
rect 635 1471 636 1475
rect 672 1472 674 1481
rect 726 1475 732 1476
rect 630 1470 636 1471
rect 670 1471 676 1472
rect 614 1466 620 1467
rect 606 1443 612 1444
rect 606 1439 607 1443
rect 611 1439 612 1443
rect 606 1438 612 1439
rect 578 1435 584 1436
rect 110 1431 116 1432
rect 110 1427 111 1431
rect 115 1427 116 1431
rect 578 1431 579 1435
rect 583 1431 584 1435
rect 578 1430 584 1431
rect 110 1426 116 1427
rect 112 1415 114 1426
rect 318 1424 324 1425
rect 318 1420 319 1424
rect 323 1420 324 1424
rect 318 1419 324 1420
rect 358 1424 364 1425
rect 358 1420 359 1424
rect 363 1420 364 1424
rect 358 1419 364 1420
rect 398 1424 404 1425
rect 398 1420 399 1424
rect 403 1420 404 1424
rect 398 1419 404 1420
rect 446 1424 452 1425
rect 446 1420 447 1424
rect 451 1420 452 1424
rect 446 1419 452 1420
rect 502 1424 508 1425
rect 502 1420 503 1424
rect 507 1420 508 1424
rect 502 1419 508 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 614 1424 620 1425
rect 614 1420 615 1424
rect 619 1420 620 1424
rect 614 1419 620 1420
rect 320 1415 322 1419
rect 360 1415 362 1419
rect 400 1415 402 1419
rect 448 1415 450 1419
rect 504 1415 506 1419
rect 560 1415 562 1419
rect 616 1415 618 1419
rect 111 1414 115 1415
rect 111 1409 115 1410
rect 263 1414 267 1415
rect 263 1409 267 1410
rect 303 1414 307 1415
rect 303 1409 307 1410
rect 319 1414 323 1415
rect 319 1409 323 1410
rect 343 1414 347 1415
rect 343 1409 347 1410
rect 359 1414 363 1415
rect 359 1409 363 1410
rect 391 1414 395 1415
rect 391 1409 395 1410
rect 399 1414 403 1415
rect 399 1409 403 1410
rect 447 1414 451 1415
rect 447 1409 451 1410
rect 503 1414 507 1415
rect 503 1409 507 1410
rect 559 1414 563 1415
rect 559 1409 563 1410
rect 615 1414 619 1415
rect 615 1409 619 1410
rect 623 1414 627 1415
rect 623 1409 627 1410
rect 112 1402 114 1409
rect 262 1408 268 1409
rect 262 1404 263 1408
rect 267 1404 268 1408
rect 262 1403 268 1404
rect 302 1408 308 1409
rect 302 1404 303 1408
rect 307 1404 308 1408
rect 302 1403 308 1404
rect 342 1408 348 1409
rect 342 1404 343 1408
rect 347 1404 348 1408
rect 342 1403 348 1404
rect 390 1408 396 1409
rect 390 1404 391 1408
rect 395 1404 396 1408
rect 390 1403 396 1404
rect 446 1408 452 1409
rect 446 1404 447 1408
rect 451 1404 452 1408
rect 446 1403 452 1404
rect 502 1408 508 1409
rect 502 1404 503 1408
rect 507 1404 508 1408
rect 502 1403 508 1404
rect 558 1408 564 1409
rect 558 1404 559 1408
rect 563 1404 564 1408
rect 558 1403 564 1404
rect 622 1408 628 1409
rect 622 1404 623 1408
rect 627 1404 628 1408
rect 622 1403 628 1404
rect 110 1401 116 1402
rect 110 1397 111 1401
rect 115 1397 116 1401
rect 110 1396 116 1397
rect 632 1388 634 1470
rect 670 1467 671 1471
rect 675 1467 676 1471
rect 726 1471 727 1475
rect 731 1471 732 1475
rect 736 1472 738 1481
rect 790 1475 796 1476
rect 726 1470 732 1471
rect 734 1471 740 1472
rect 670 1466 676 1467
rect 728 1444 730 1470
rect 734 1467 735 1471
rect 739 1467 740 1471
rect 790 1471 791 1475
rect 795 1471 796 1475
rect 800 1472 802 1481
rect 846 1475 852 1476
rect 790 1470 796 1471
rect 798 1471 804 1472
rect 734 1466 740 1467
rect 792 1444 794 1470
rect 798 1467 799 1471
rect 803 1467 804 1471
rect 846 1471 847 1475
rect 851 1471 852 1475
rect 856 1472 858 1481
rect 902 1475 908 1476
rect 846 1470 852 1471
rect 854 1471 860 1472
rect 798 1466 804 1467
rect 848 1444 850 1470
rect 854 1467 855 1471
rect 859 1467 860 1471
rect 902 1471 903 1475
rect 907 1471 908 1475
rect 912 1472 914 1481
rect 958 1475 964 1476
rect 902 1470 908 1471
rect 910 1471 916 1472
rect 854 1466 860 1467
rect 904 1444 906 1470
rect 910 1467 911 1471
rect 915 1467 916 1471
rect 958 1471 959 1475
rect 963 1471 964 1475
rect 968 1472 970 1481
rect 1014 1475 1020 1476
rect 958 1470 964 1471
rect 966 1471 972 1472
rect 910 1466 916 1467
rect 960 1444 962 1470
rect 966 1467 967 1471
rect 971 1467 972 1471
rect 1014 1471 1015 1475
rect 1019 1471 1020 1475
rect 1024 1472 1026 1481
rect 1088 1472 1090 1481
rect 1152 1472 1154 1481
rect 1180 1476 1182 1518
rect 1190 1505 1196 1506
rect 1190 1501 1191 1505
rect 1195 1501 1196 1505
rect 1190 1500 1196 1501
rect 1208 1500 1210 1526
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1278 1528 1279 1532
rect 1283 1528 1284 1532
rect 1278 1527 1284 1528
rect 1238 1523 1244 1524
rect 1192 1487 1194 1500
rect 1206 1499 1212 1500
rect 1206 1495 1207 1499
rect 1211 1495 1212 1499
rect 1206 1494 1212 1495
rect 1240 1487 1242 1523
rect 1191 1486 1195 1487
rect 1191 1481 1195 1482
rect 1239 1486 1243 1487
rect 1239 1481 1243 1482
rect 1178 1475 1184 1476
rect 1014 1470 1020 1471
rect 1022 1471 1028 1472
rect 966 1466 972 1467
rect 726 1443 732 1444
rect 726 1439 727 1443
rect 731 1439 732 1443
rect 726 1438 732 1439
rect 790 1443 796 1444
rect 790 1439 791 1443
rect 795 1439 796 1443
rect 790 1438 796 1439
rect 846 1443 852 1444
rect 846 1439 847 1443
rect 851 1439 852 1443
rect 846 1438 852 1439
rect 902 1443 908 1444
rect 902 1439 903 1443
rect 907 1439 908 1443
rect 902 1438 908 1439
rect 958 1443 964 1444
rect 958 1439 959 1443
rect 963 1439 964 1443
rect 958 1438 964 1439
rect 838 1435 844 1436
rect 838 1431 839 1435
rect 843 1431 844 1435
rect 838 1430 844 1431
rect 670 1424 676 1425
rect 670 1420 671 1424
rect 675 1420 676 1424
rect 670 1419 676 1420
rect 734 1424 740 1425
rect 734 1420 735 1424
rect 739 1420 740 1424
rect 734 1419 740 1420
rect 798 1424 804 1425
rect 798 1420 799 1424
rect 803 1420 804 1424
rect 798 1419 804 1420
rect 672 1415 674 1419
rect 736 1415 738 1419
rect 800 1415 802 1419
rect 671 1414 675 1415
rect 671 1409 675 1410
rect 687 1414 691 1415
rect 687 1409 691 1410
rect 735 1414 739 1415
rect 735 1409 739 1410
rect 751 1414 755 1415
rect 751 1409 755 1410
rect 799 1414 803 1415
rect 799 1409 803 1410
rect 815 1414 819 1415
rect 815 1409 819 1410
rect 686 1408 692 1409
rect 686 1404 687 1408
rect 691 1404 692 1408
rect 686 1403 692 1404
rect 750 1408 756 1409
rect 750 1404 751 1408
rect 755 1404 756 1408
rect 750 1403 756 1404
rect 814 1408 820 1409
rect 814 1404 815 1408
rect 819 1404 820 1408
rect 814 1403 820 1404
rect 310 1387 316 1388
rect 110 1384 116 1385
rect 110 1380 111 1384
rect 115 1380 116 1384
rect 310 1383 311 1387
rect 315 1383 316 1387
rect 310 1382 316 1383
rect 406 1387 412 1388
rect 406 1383 407 1387
rect 411 1383 412 1387
rect 406 1382 412 1383
rect 462 1387 468 1388
rect 462 1383 463 1387
rect 467 1383 468 1387
rect 462 1382 468 1383
rect 518 1387 524 1388
rect 518 1383 519 1387
rect 523 1383 524 1387
rect 518 1382 524 1383
rect 574 1387 580 1388
rect 574 1383 575 1387
rect 579 1383 580 1387
rect 574 1382 580 1383
rect 630 1387 636 1388
rect 630 1383 631 1387
rect 635 1383 636 1387
rect 630 1382 636 1383
rect 110 1379 116 1380
rect 112 1343 114 1379
rect 262 1361 268 1362
rect 262 1357 263 1361
rect 267 1357 268 1361
rect 262 1356 268 1357
rect 302 1361 308 1362
rect 302 1357 303 1361
rect 307 1357 308 1361
rect 302 1356 308 1357
rect 312 1356 314 1382
rect 366 1379 372 1380
rect 366 1375 367 1379
rect 371 1375 372 1379
rect 366 1374 372 1375
rect 342 1361 348 1362
rect 342 1357 343 1361
rect 347 1357 348 1361
rect 342 1356 348 1357
rect 368 1356 370 1374
rect 390 1361 396 1362
rect 390 1357 391 1361
rect 395 1357 396 1361
rect 390 1356 396 1357
rect 408 1356 410 1382
rect 446 1361 452 1362
rect 446 1357 447 1361
rect 451 1357 452 1361
rect 446 1356 452 1357
rect 464 1356 466 1382
rect 502 1361 508 1362
rect 502 1357 503 1361
rect 507 1357 508 1361
rect 502 1356 508 1357
rect 520 1356 522 1382
rect 558 1361 564 1362
rect 558 1357 559 1361
rect 563 1357 564 1361
rect 558 1356 564 1357
rect 576 1356 578 1382
rect 782 1379 788 1380
rect 782 1375 783 1379
rect 787 1375 788 1379
rect 782 1374 788 1375
rect 622 1361 628 1362
rect 622 1357 623 1361
rect 627 1357 628 1361
rect 622 1356 628 1357
rect 686 1361 692 1362
rect 686 1357 687 1361
rect 691 1357 692 1361
rect 686 1356 692 1357
rect 750 1361 756 1362
rect 750 1357 751 1361
rect 755 1357 756 1361
rect 750 1356 756 1357
rect 264 1343 266 1356
rect 304 1343 306 1356
rect 310 1355 316 1356
rect 310 1351 311 1355
rect 315 1351 316 1355
rect 310 1350 316 1351
rect 344 1343 346 1356
rect 350 1355 356 1356
rect 350 1351 351 1355
rect 355 1351 356 1355
rect 350 1350 356 1351
rect 366 1355 372 1356
rect 366 1351 367 1355
rect 371 1351 372 1355
rect 366 1350 372 1351
rect 111 1342 115 1343
rect 111 1337 115 1338
rect 135 1342 139 1343
rect 135 1337 139 1338
rect 175 1342 179 1343
rect 175 1337 179 1338
rect 215 1342 219 1343
rect 215 1337 219 1338
rect 255 1342 259 1343
rect 255 1337 259 1338
rect 263 1342 267 1343
rect 263 1337 267 1338
rect 303 1342 307 1343
rect 303 1337 307 1338
rect 327 1342 331 1343
rect 327 1337 331 1338
rect 343 1342 347 1343
rect 343 1337 347 1338
rect 112 1305 114 1337
rect 136 1328 138 1337
rect 176 1328 178 1337
rect 190 1335 196 1336
rect 190 1331 191 1335
rect 195 1331 196 1335
rect 190 1330 196 1331
rect 202 1331 208 1332
rect 134 1327 140 1328
rect 134 1323 135 1327
rect 139 1323 140 1327
rect 134 1322 140 1323
rect 174 1327 180 1328
rect 174 1323 175 1327
rect 179 1323 180 1327
rect 174 1322 180 1323
rect 162 1319 168 1320
rect 162 1315 163 1319
rect 167 1315 168 1319
rect 162 1314 168 1315
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 164 1300 166 1314
rect 192 1300 194 1330
rect 202 1327 203 1331
rect 207 1327 208 1331
rect 216 1328 218 1337
rect 238 1331 244 1332
rect 202 1326 208 1327
rect 214 1327 220 1328
rect 204 1308 206 1326
rect 214 1323 215 1327
rect 219 1323 220 1327
rect 238 1327 239 1331
rect 243 1327 244 1331
rect 256 1328 258 1337
rect 328 1328 330 1337
rect 238 1326 244 1327
rect 254 1327 260 1328
rect 214 1322 220 1323
rect 202 1307 208 1308
rect 202 1303 203 1307
rect 207 1303 208 1307
rect 202 1302 208 1303
rect 110 1299 116 1300
rect 162 1299 168 1300
rect 162 1295 163 1299
rect 167 1295 168 1299
rect 162 1294 168 1295
rect 190 1299 196 1300
rect 190 1295 191 1299
rect 195 1295 196 1299
rect 190 1294 196 1295
rect 110 1287 116 1288
rect 110 1283 111 1287
rect 115 1283 116 1287
rect 110 1282 116 1283
rect 112 1271 114 1282
rect 134 1280 140 1281
rect 134 1276 135 1280
rect 139 1276 140 1280
rect 134 1275 140 1276
rect 174 1280 180 1281
rect 174 1276 175 1280
rect 179 1276 180 1280
rect 174 1275 180 1276
rect 214 1280 220 1281
rect 214 1276 215 1280
rect 219 1276 220 1280
rect 214 1275 220 1276
rect 136 1271 138 1275
rect 176 1271 178 1275
rect 216 1271 218 1275
rect 111 1270 115 1271
rect 111 1265 115 1266
rect 135 1270 139 1271
rect 135 1265 139 1266
rect 175 1270 179 1271
rect 175 1265 179 1266
rect 215 1270 219 1271
rect 215 1265 219 1266
rect 112 1258 114 1265
rect 134 1264 140 1265
rect 134 1260 135 1264
rect 139 1260 140 1264
rect 134 1259 140 1260
rect 174 1264 180 1265
rect 174 1260 175 1264
rect 179 1260 180 1264
rect 174 1259 180 1260
rect 110 1257 116 1258
rect 110 1253 111 1257
rect 115 1253 116 1257
rect 110 1252 116 1253
rect 240 1244 242 1326
rect 254 1323 255 1327
rect 259 1323 260 1327
rect 254 1322 260 1323
rect 326 1327 332 1328
rect 326 1323 327 1327
rect 331 1323 332 1327
rect 326 1322 332 1323
rect 352 1300 354 1350
rect 392 1343 394 1356
rect 406 1355 412 1356
rect 406 1351 407 1355
rect 411 1351 412 1355
rect 406 1350 412 1351
rect 448 1343 450 1356
rect 462 1355 468 1356
rect 462 1351 463 1355
rect 467 1351 468 1355
rect 462 1350 468 1351
rect 504 1343 506 1356
rect 518 1355 524 1356
rect 518 1351 519 1355
rect 523 1351 524 1355
rect 518 1350 524 1351
rect 560 1343 562 1356
rect 574 1355 580 1356
rect 574 1351 575 1355
rect 579 1351 580 1355
rect 574 1350 580 1351
rect 624 1343 626 1356
rect 688 1343 690 1356
rect 752 1343 754 1356
rect 391 1342 395 1343
rect 391 1337 395 1338
rect 407 1342 411 1343
rect 407 1337 411 1338
rect 447 1342 451 1343
rect 447 1337 451 1338
rect 495 1342 499 1343
rect 495 1337 499 1338
rect 503 1342 507 1343
rect 503 1337 507 1338
rect 559 1342 563 1343
rect 559 1337 563 1338
rect 583 1342 587 1343
rect 583 1337 587 1338
rect 623 1342 627 1343
rect 623 1337 627 1338
rect 671 1342 675 1343
rect 671 1337 675 1338
rect 687 1342 691 1343
rect 687 1337 691 1338
rect 751 1342 755 1343
rect 751 1337 755 1338
rect 759 1342 763 1343
rect 759 1337 763 1338
rect 398 1331 404 1332
rect 398 1327 399 1331
rect 403 1327 404 1331
rect 408 1328 410 1337
rect 486 1331 492 1332
rect 398 1326 404 1327
rect 406 1327 412 1328
rect 400 1300 402 1326
rect 406 1323 407 1327
rect 411 1323 412 1327
rect 486 1327 487 1331
rect 491 1327 492 1331
rect 496 1328 498 1337
rect 506 1331 512 1332
rect 486 1326 492 1327
rect 494 1327 500 1328
rect 406 1322 412 1323
rect 488 1300 490 1326
rect 494 1323 495 1327
rect 499 1323 500 1327
rect 506 1327 507 1331
rect 511 1327 512 1331
rect 584 1328 586 1337
rect 662 1331 668 1332
rect 506 1326 512 1327
rect 582 1327 588 1328
rect 494 1322 500 1323
rect 508 1308 510 1326
rect 582 1323 583 1327
rect 587 1323 588 1327
rect 662 1327 663 1331
rect 667 1327 668 1331
rect 672 1328 674 1337
rect 750 1331 756 1332
rect 662 1326 668 1327
rect 670 1327 676 1328
rect 582 1322 588 1323
rect 506 1307 512 1308
rect 506 1303 507 1307
rect 511 1303 512 1307
rect 506 1302 512 1303
rect 664 1300 666 1326
rect 670 1323 671 1327
rect 675 1323 676 1327
rect 750 1327 751 1331
rect 755 1327 756 1331
rect 760 1328 762 1337
rect 784 1332 786 1374
rect 814 1361 820 1362
rect 814 1357 815 1361
rect 819 1357 820 1361
rect 814 1356 820 1357
rect 840 1356 842 1430
rect 854 1424 860 1425
rect 854 1420 855 1424
rect 859 1420 860 1424
rect 854 1419 860 1420
rect 910 1424 916 1425
rect 910 1420 911 1424
rect 915 1420 916 1424
rect 910 1419 916 1420
rect 966 1424 972 1425
rect 966 1420 967 1424
rect 971 1420 972 1424
rect 966 1419 972 1420
rect 856 1415 858 1419
rect 912 1415 914 1419
rect 968 1415 970 1419
rect 855 1414 859 1415
rect 855 1409 859 1410
rect 879 1414 883 1415
rect 879 1409 883 1410
rect 911 1414 915 1415
rect 911 1409 915 1410
rect 951 1414 955 1415
rect 951 1409 955 1410
rect 967 1414 971 1415
rect 967 1409 971 1410
rect 878 1408 884 1409
rect 878 1404 879 1408
rect 883 1404 884 1408
rect 878 1403 884 1404
rect 950 1408 956 1409
rect 950 1404 951 1408
rect 955 1404 956 1408
rect 950 1403 956 1404
rect 1016 1396 1018 1470
rect 1022 1467 1023 1471
rect 1027 1467 1028 1471
rect 1022 1466 1028 1467
rect 1086 1471 1092 1472
rect 1086 1467 1087 1471
rect 1091 1467 1092 1471
rect 1086 1466 1092 1467
rect 1150 1471 1156 1472
rect 1150 1467 1151 1471
rect 1155 1467 1156 1471
rect 1178 1471 1179 1475
rect 1183 1471 1184 1475
rect 1192 1472 1194 1481
rect 1202 1475 1208 1476
rect 1178 1470 1184 1471
rect 1190 1471 1196 1472
rect 1150 1466 1156 1467
rect 1190 1467 1191 1471
rect 1195 1467 1196 1471
rect 1202 1471 1203 1475
rect 1207 1471 1208 1475
rect 1202 1470 1208 1471
rect 1190 1466 1196 1467
rect 1110 1463 1116 1464
rect 1110 1459 1111 1463
rect 1115 1459 1116 1463
rect 1110 1458 1116 1459
rect 1112 1444 1114 1458
rect 1204 1452 1206 1470
rect 1218 1467 1224 1468
rect 1218 1463 1219 1467
rect 1223 1463 1224 1467
rect 1218 1462 1224 1463
rect 1202 1451 1208 1452
rect 1202 1447 1203 1451
rect 1207 1447 1208 1451
rect 1202 1446 1208 1447
rect 1220 1444 1222 1462
rect 1240 1449 1242 1481
rect 1280 1475 1282 1527
rect 1470 1509 1476 1510
rect 1470 1505 1471 1509
rect 1475 1505 1476 1509
rect 1470 1504 1476 1505
rect 1512 1504 1514 1582
rect 1558 1568 1564 1569
rect 1558 1564 1559 1568
rect 1563 1564 1564 1568
rect 1558 1563 1564 1564
rect 1630 1568 1636 1569
rect 1630 1564 1631 1568
rect 1635 1564 1636 1568
rect 1630 1563 1636 1564
rect 1702 1568 1708 1569
rect 1702 1564 1703 1568
rect 1707 1564 1708 1568
rect 1702 1563 1708 1564
rect 1782 1568 1788 1569
rect 1782 1564 1783 1568
rect 1787 1564 1788 1568
rect 1782 1563 1788 1564
rect 1559 1562 1563 1563
rect 1559 1557 1563 1558
rect 1623 1562 1627 1563
rect 1623 1557 1627 1558
rect 1631 1562 1635 1563
rect 1631 1557 1635 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1759 1562 1763 1563
rect 1759 1557 1763 1558
rect 1783 1562 1787 1563
rect 1783 1557 1787 1558
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1758 1556 1764 1557
rect 1758 1552 1759 1556
rect 1763 1552 1764 1556
rect 1758 1551 1764 1552
rect 1796 1544 1798 1614
rect 1854 1611 1855 1615
rect 1859 1611 1860 1615
rect 1918 1615 1919 1619
rect 1923 1615 1924 1619
rect 1928 1616 1930 1625
rect 1956 1620 1958 1670
rect 1974 1649 1980 1650
rect 1974 1645 1975 1649
rect 1979 1645 1980 1649
rect 1974 1644 1980 1645
rect 2030 1649 2036 1650
rect 2030 1645 2031 1649
rect 2035 1645 2036 1649
rect 2030 1644 2036 1645
rect 2086 1649 2092 1650
rect 2086 1645 2087 1649
rect 2091 1645 2092 1649
rect 2086 1644 2092 1645
rect 2112 1644 2114 1678
rect 2406 1672 2412 1673
rect 2406 1668 2407 1672
rect 2411 1668 2412 1672
rect 2406 1667 2412 1668
rect 1976 1631 1978 1644
rect 2032 1631 2034 1644
rect 2088 1631 2090 1644
rect 2110 1643 2116 1644
rect 2110 1639 2111 1643
rect 2115 1639 2116 1643
rect 2110 1638 2116 1639
rect 2408 1631 2410 1667
rect 1975 1630 1979 1631
rect 1975 1625 1979 1626
rect 1999 1630 2003 1631
rect 1999 1625 2003 1626
rect 2031 1630 2035 1631
rect 2031 1625 2035 1626
rect 2063 1630 2067 1631
rect 2063 1625 2067 1626
rect 2087 1630 2091 1631
rect 2087 1625 2091 1626
rect 2127 1630 2131 1631
rect 2127 1625 2131 1626
rect 2191 1630 2195 1631
rect 2191 1625 2195 1626
rect 2255 1630 2259 1631
rect 2255 1625 2259 1626
rect 2319 1630 2323 1631
rect 2319 1625 2323 1626
rect 2359 1630 2363 1631
rect 2359 1625 2363 1626
rect 2407 1630 2411 1631
rect 2407 1625 2411 1626
rect 1954 1619 1960 1620
rect 1918 1614 1924 1615
rect 1926 1615 1932 1616
rect 1854 1610 1860 1611
rect 1920 1588 1922 1614
rect 1926 1611 1927 1615
rect 1931 1611 1932 1615
rect 1954 1615 1955 1619
rect 1959 1615 1960 1619
rect 2000 1616 2002 1625
rect 2010 1619 2016 1620
rect 1954 1614 1960 1615
rect 1998 1615 2004 1616
rect 1926 1610 1932 1611
rect 1998 1611 1999 1615
rect 2003 1611 2004 1615
rect 2010 1615 2011 1619
rect 2015 1615 2016 1619
rect 2064 1616 2066 1625
rect 2118 1619 2124 1620
rect 2010 1614 2016 1615
rect 2062 1615 2068 1616
rect 1998 1610 2004 1611
rect 2012 1596 2014 1614
rect 2062 1611 2063 1615
rect 2067 1611 2068 1615
rect 2118 1615 2119 1619
rect 2123 1615 2124 1619
rect 2128 1616 2130 1625
rect 2182 1619 2188 1620
rect 2118 1614 2124 1615
rect 2126 1615 2132 1616
rect 2062 1610 2068 1611
rect 2010 1595 2016 1596
rect 2010 1591 2011 1595
rect 2015 1591 2016 1595
rect 2010 1590 2016 1591
rect 2120 1588 2122 1614
rect 2126 1611 2127 1615
rect 2131 1611 2132 1615
rect 2182 1615 2183 1619
rect 2187 1615 2188 1619
rect 2192 1616 2194 1625
rect 2202 1619 2208 1620
rect 2182 1614 2188 1615
rect 2190 1615 2196 1616
rect 2126 1610 2132 1611
rect 2184 1588 2186 1614
rect 2190 1611 2191 1615
rect 2195 1611 2196 1615
rect 2202 1615 2203 1619
rect 2207 1615 2208 1619
rect 2256 1616 2258 1625
rect 2278 1619 2284 1620
rect 2202 1614 2208 1615
rect 2254 1615 2260 1616
rect 2190 1610 2196 1611
rect 2204 1596 2206 1614
rect 2254 1611 2255 1615
rect 2259 1611 2260 1615
rect 2278 1615 2279 1619
rect 2283 1615 2284 1619
rect 2320 1616 2322 1625
rect 2330 1619 2336 1620
rect 2278 1614 2284 1615
rect 2318 1615 2324 1616
rect 2254 1610 2260 1611
rect 2202 1595 2208 1596
rect 2202 1591 2203 1595
rect 2207 1591 2208 1595
rect 2202 1590 2208 1591
rect 1918 1587 1924 1588
rect 1918 1583 1919 1587
rect 1923 1583 1924 1587
rect 1918 1582 1924 1583
rect 2042 1587 2048 1588
rect 2042 1583 2043 1587
rect 2047 1583 2048 1587
rect 2042 1582 2048 1583
rect 2118 1587 2124 1588
rect 2118 1583 2119 1587
rect 2123 1583 2124 1587
rect 2118 1582 2124 1583
rect 2182 1587 2188 1588
rect 2182 1583 2183 1587
rect 2187 1583 2188 1587
rect 2182 1582 2188 1583
rect 1854 1568 1860 1569
rect 1854 1564 1855 1568
rect 1859 1564 1860 1568
rect 1854 1563 1860 1564
rect 1926 1568 1932 1569
rect 1926 1564 1927 1568
rect 1931 1564 1932 1568
rect 1926 1563 1932 1564
rect 1998 1568 2004 1569
rect 1998 1564 1999 1568
rect 2003 1564 2004 1568
rect 1998 1563 2004 1564
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1871 1562 1875 1563
rect 1871 1557 1875 1558
rect 1927 1562 1931 1563
rect 1927 1557 1931 1558
rect 1967 1562 1971 1563
rect 1967 1557 1971 1558
rect 1999 1562 2003 1563
rect 1999 1557 2003 1558
rect 1870 1556 1876 1557
rect 1870 1552 1871 1556
rect 1875 1552 1876 1556
rect 1870 1551 1876 1552
rect 1966 1556 1972 1557
rect 1966 1552 1967 1556
rect 1971 1552 1972 1556
rect 1966 1551 1972 1552
rect 1794 1543 1800 1544
rect 1794 1539 1795 1543
rect 1799 1539 1800 1543
rect 1794 1538 1800 1539
rect 1638 1535 1644 1536
rect 1638 1531 1639 1535
rect 1643 1531 1644 1535
rect 1638 1530 1644 1531
rect 1622 1509 1628 1510
rect 1622 1505 1623 1509
rect 1627 1505 1628 1509
rect 1622 1504 1628 1505
rect 1640 1504 1642 1530
rect 1758 1509 1764 1510
rect 1758 1505 1759 1509
rect 1763 1505 1764 1509
rect 1758 1504 1764 1505
rect 1870 1509 1876 1510
rect 1870 1505 1871 1509
rect 1875 1505 1876 1509
rect 1870 1504 1876 1505
rect 1966 1509 1972 1510
rect 1966 1505 1967 1509
rect 1971 1505 1972 1509
rect 1966 1504 1972 1505
rect 2044 1504 2046 1582
rect 2062 1568 2068 1569
rect 2062 1564 2063 1568
rect 2067 1564 2068 1568
rect 2062 1563 2068 1564
rect 2126 1568 2132 1569
rect 2126 1564 2127 1568
rect 2131 1564 2132 1568
rect 2126 1563 2132 1564
rect 2190 1568 2196 1569
rect 2190 1564 2191 1568
rect 2195 1564 2196 1568
rect 2190 1563 2196 1564
rect 2254 1568 2260 1569
rect 2254 1564 2255 1568
rect 2259 1564 2260 1568
rect 2254 1563 2260 1564
rect 2055 1562 2059 1563
rect 2055 1557 2059 1558
rect 2063 1562 2067 1563
rect 2063 1557 2067 1558
rect 2127 1562 2131 1563
rect 2127 1557 2131 1558
rect 2191 1562 2195 1563
rect 2191 1557 2195 1558
rect 2255 1562 2259 1563
rect 2255 1557 2259 1558
rect 2054 1556 2060 1557
rect 2054 1552 2055 1556
rect 2059 1552 2060 1556
rect 2054 1551 2060 1552
rect 2126 1556 2132 1557
rect 2126 1552 2127 1556
rect 2131 1552 2132 1556
rect 2126 1551 2132 1552
rect 2190 1556 2196 1557
rect 2190 1552 2191 1556
rect 2195 1552 2196 1556
rect 2190 1551 2196 1552
rect 2254 1556 2260 1557
rect 2254 1552 2255 1556
rect 2259 1552 2260 1556
rect 2254 1551 2260 1552
rect 2280 1536 2282 1614
rect 2318 1611 2319 1615
rect 2323 1611 2324 1615
rect 2330 1615 2331 1619
rect 2335 1615 2336 1619
rect 2360 1616 2362 1625
rect 2370 1619 2376 1620
rect 2330 1614 2336 1615
rect 2358 1615 2364 1616
rect 2318 1610 2324 1611
rect 2332 1588 2334 1614
rect 2358 1611 2359 1615
rect 2363 1611 2364 1615
rect 2370 1615 2371 1619
rect 2375 1615 2376 1619
rect 2370 1614 2376 1615
rect 2358 1610 2364 1611
rect 2372 1588 2374 1614
rect 2408 1593 2410 1625
rect 2406 1592 2412 1593
rect 2406 1588 2407 1592
rect 2411 1588 2412 1592
rect 2330 1587 2336 1588
rect 2330 1583 2331 1587
rect 2335 1583 2336 1587
rect 2330 1582 2336 1583
rect 2370 1587 2376 1588
rect 2406 1587 2412 1588
rect 2370 1583 2371 1587
rect 2375 1583 2376 1587
rect 2370 1582 2376 1583
rect 2346 1579 2352 1580
rect 2346 1575 2347 1579
rect 2351 1575 2352 1579
rect 2346 1574 2352 1575
rect 2406 1575 2412 1576
rect 2318 1568 2324 1569
rect 2318 1564 2319 1568
rect 2323 1564 2324 1568
rect 2318 1563 2324 1564
rect 2319 1562 2323 1563
rect 2319 1557 2323 1558
rect 2318 1556 2324 1557
rect 2318 1552 2319 1556
rect 2323 1552 2324 1556
rect 2318 1551 2324 1552
rect 2142 1535 2148 1536
rect 2142 1531 2143 1535
rect 2147 1531 2148 1535
rect 2142 1530 2148 1531
rect 2206 1535 2212 1536
rect 2206 1531 2207 1535
rect 2211 1531 2212 1535
rect 2206 1530 2212 1531
rect 2270 1535 2276 1536
rect 2270 1531 2271 1535
rect 2275 1531 2276 1535
rect 2270 1530 2276 1531
rect 2278 1535 2284 1536
rect 2278 1531 2279 1535
rect 2283 1531 2284 1535
rect 2278 1530 2284 1531
rect 2078 1527 2084 1528
rect 2078 1523 2079 1527
rect 2083 1523 2084 1527
rect 2078 1522 2084 1523
rect 2054 1509 2060 1510
rect 2054 1505 2055 1509
rect 2059 1505 2060 1509
rect 2054 1504 2060 1505
rect 2080 1504 2082 1522
rect 2126 1509 2132 1510
rect 2126 1505 2127 1509
rect 2131 1505 2132 1509
rect 2126 1504 2132 1505
rect 2144 1504 2146 1530
rect 2190 1509 2196 1510
rect 2190 1505 2191 1509
rect 2195 1505 2196 1509
rect 2190 1504 2196 1505
rect 2208 1504 2210 1530
rect 2254 1509 2260 1510
rect 2254 1505 2255 1509
rect 2259 1505 2260 1509
rect 2254 1504 2260 1505
rect 2272 1504 2274 1530
rect 2318 1509 2324 1510
rect 2318 1505 2319 1509
rect 2323 1505 2324 1509
rect 2318 1504 2324 1505
rect 2348 1504 2350 1574
rect 2406 1571 2407 1575
rect 2411 1571 2412 1575
rect 2406 1570 2412 1571
rect 2358 1568 2364 1569
rect 2358 1564 2359 1568
rect 2363 1564 2364 1568
rect 2358 1563 2364 1564
rect 2408 1563 2410 1570
rect 2359 1562 2363 1563
rect 2359 1557 2363 1558
rect 2407 1562 2411 1563
rect 2407 1557 2411 1558
rect 2358 1556 2364 1557
rect 2358 1552 2359 1556
rect 2363 1552 2364 1556
rect 2358 1551 2364 1552
rect 2408 1550 2410 1557
rect 2406 1549 2412 1550
rect 2406 1545 2407 1549
rect 2411 1545 2412 1549
rect 2406 1544 2412 1545
rect 2374 1535 2380 1536
rect 2374 1531 2375 1535
rect 2379 1531 2380 1535
rect 2374 1530 2380 1531
rect 2382 1535 2388 1536
rect 2382 1531 2383 1535
rect 2387 1531 2388 1535
rect 2382 1530 2388 1531
rect 2406 1532 2412 1533
rect 2358 1509 2364 1510
rect 2358 1505 2359 1509
rect 2363 1505 2364 1509
rect 2358 1504 2364 1505
rect 2376 1504 2378 1530
rect 1472 1475 1474 1504
rect 1510 1503 1516 1504
rect 1510 1499 1511 1503
rect 1515 1499 1516 1503
rect 1510 1498 1516 1499
rect 1624 1475 1626 1504
rect 1638 1503 1644 1504
rect 1638 1499 1639 1503
rect 1643 1499 1644 1503
rect 1638 1498 1644 1499
rect 1760 1475 1762 1504
rect 1872 1475 1874 1504
rect 1968 1475 1970 1504
rect 2042 1503 2048 1504
rect 2042 1499 2043 1503
rect 2047 1499 2048 1503
rect 2042 1498 2048 1499
rect 2056 1475 2058 1504
rect 2078 1503 2084 1504
rect 2078 1499 2079 1503
rect 2083 1499 2084 1503
rect 2078 1498 2084 1499
rect 2128 1475 2130 1504
rect 2142 1503 2148 1504
rect 2142 1499 2143 1503
rect 2147 1499 2148 1503
rect 2142 1498 2148 1499
rect 2192 1475 2194 1504
rect 2206 1503 2212 1504
rect 2206 1499 2207 1503
rect 2211 1499 2212 1503
rect 2206 1498 2212 1499
rect 2256 1475 2258 1504
rect 2270 1503 2276 1504
rect 2270 1499 2271 1503
rect 2275 1499 2276 1503
rect 2270 1498 2276 1499
rect 2320 1475 2322 1504
rect 2346 1503 2352 1504
rect 2346 1499 2347 1503
rect 2351 1499 2352 1503
rect 2346 1498 2352 1499
rect 2360 1475 2362 1504
rect 2374 1503 2380 1504
rect 2374 1499 2375 1503
rect 2379 1499 2380 1503
rect 2374 1498 2380 1499
rect 1279 1474 1283 1475
rect 1279 1469 1283 1470
rect 1303 1474 1307 1475
rect 1303 1469 1307 1470
rect 1375 1474 1379 1475
rect 1375 1469 1379 1470
rect 1471 1474 1475 1475
rect 1471 1469 1475 1470
rect 1479 1474 1483 1475
rect 1479 1469 1483 1470
rect 1583 1474 1587 1475
rect 1583 1469 1587 1470
rect 1623 1474 1627 1475
rect 1623 1469 1627 1470
rect 1687 1474 1691 1475
rect 1687 1469 1691 1470
rect 1759 1474 1763 1475
rect 1759 1469 1763 1470
rect 1783 1474 1787 1475
rect 1783 1469 1787 1470
rect 1871 1474 1875 1475
rect 1871 1469 1875 1470
rect 1951 1474 1955 1475
rect 1951 1469 1955 1470
rect 1967 1474 1971 1475
rect 1967 1469 1971 1470
rect 2031 1474 2035 1475
rect 2031 1469 2035 1470
rect 2055 1474 2059 1475
rect 2055 1469 2059 1470
rect 2103 1474 2107 1475
rect 2103 1469 2107 1470
rect 2127 1474 2131 1475
rect 2127 1469 2131 1470
rect 2167 1474 2171 1475
rect 2167 1469 2171 1470
rect 2191 1474 2195 1475
rect 2191 1469 2195 1470
rect 2239 1474 2243 1475
rect 2239 1469 2243 1470
rect 2255 1474 2259 1475
rect 2255 1469 2259 1470
rect 2311 1474 2315 1475
rect 2311 1469 2315 1470
rect 2319 1474 2323 1475
rect 2319 1469 2323 1470
rect 2359 1474 2363 1475
rect 2359 1469 2363 1470
rect 1238 1448 1244 1449
rect 1238 1444 1239 1448
rect 1243 1444 1244 1448
rect 1110 1443 1116 1444
rect 1110 1439 1111 1443
rect 1115 1439 1116 1443
rect 1110 1438 1116 1439
rect 1218 1443 1224 1444
rect 1238 1443 1244 1444
rect 1218 1439 1219 1443
rect 1223 1439 1224 1443
rect 1218 1438 1224 1439
rect 1280 1437 1282 1469
rect 1304 1460 1306 1469
rect 1376 1460 1378 1469
rect 1386 1463 1392 1464
rect 1302 1459 1308 1460
rect 1302 1455 1303 1459
rect 1307 1455 1308 1459
rect 1302 1454 1308 1455
rect 1374 1459 1380 1460
rect 1374 1455 1375 1459
rect 1379 1455 1380 1459
rect 1386 1459 1387 1463
rect 1391 1459 1392 1463
rect 1480 1460 1482 1469
rect 1574 1463 1580 1464
rect 1386 1458 1392 1459
rect 1478 1459 1484 1460
rect 1374 1454 1380 1455
rect 1278 1436 1284 1437
rect 1278 1432 1279 1436
rect 1283 1432 1284 1436
rect 1388 1432 1390 1458
rect 1478 1455 1479 1459
rect 1483 1455 1484 1459
rect 1574 1459 1575 1463
rect 1579 1459 1580 1463
rect 1584 1460 1586 1469
rect 1678 1463 1684 1464
rect 1574 1458 1580 1459
rect 1582 1459 1588 1460
rect 1478 1454 1484 1455
rect 1576 1432 1578 1458
rect 1582 1455 1583 1459
rect 1587 1455 1588 1459
rect 1678 1459 1679 1463
rect 1683 1459 1684 1463
rect 1688 1460 1690 1469
rect 1698 1463 1704 1464
rect 1678 1458 1684 1459
rect 1686 1459 1692 1460
rect 1582 1454 1588 1455
rect 1680 1432 1682 1458
rect 1686 1455 1687 1459
rect 1691 1455 1692 1459
rect 1698 1459 1699 1463
rect 1703 1459 1704 1463
rect 1784 1460 1786 1469
rect 1872 1460 1874 1469
rect 1942 1463 1948 1464
rect 1698 1458 1704 1459
rect 1782 1459 1788 1460
rect 1686 1454 1692 1455
rect 1700 1440 1702 1458
rect 1782 1455 1783 1459
rect 1787 1455 1788 1459
rect 1782 1454 1788 1455
rect 1870 1459 1876 1460
rect 1870 1455 1871 1459
rect 1875 1455 1876 1459
rect 1942 1459 1943 1463
rect 1947 1459 1948 1463
rect 1952 1460 1954 1469
rect 2022 1463 2028 1464
rect 1942 1458 1948 1459
rect 1950 1459 1956 1460
rect 1870 1454 1876 1455
rect 1698 1439 1704 1440
rect 1698 1435 1699 1439
rect 1703 1435 1704 1439
rect 1698 1434 1704 1435
rect 1944 1432 1946 1458
rect 1950 1455 1951 1459
rect 1955 1455 1956 1459
rect 2022 1459 2023 1463
rect 2027 1459 2028 1463
rect 2032 1460 2034 1469
rect 2094 1463 2100 1464
rect 2022 1458 2028 1459
rect 2030 1459 2036 1460
rect 1950 1454 1956 1455
rect 2024 1432 2026 1458
rect 2030 1455 2031 1459
rect 2035 1455 2036 1459
rect 2094 1459 2095 1463
rect 2099 1459 2100 1463
rect 2104 1460 2106 1469
rect 2158 1463 2164 1464
rect 2094 1458 2100 1459
rect 2102 1459 2108 1460
rect 2030 1454 2036 1455
rect 2096 1432 2098 1458
rect 2102 1455 2103 1459
rect 2107 1455 2108 1459
rect 2158 1459 2159 1463
rect 2163 1459 2164 1463
rect 2168 1460 2170 1469
rect 2230 1463 2236 1464
rect 2158 1458 2164 1459
rect 2166 1459 2172 1460
rect 2102 1454 2108 1455
rect 2160 1432 2162 1458
rect 2166 1455 2167 1459
rect 2171 1455 2172 1459
rect 2230 1459 2231 1463
rect 2235 1459 2236 1463
rect 2240 1460 2242 1469
rect 2302 1463 2308 1464
rect 2230 1458 2236 1459
rect 2238 1459 2244 1460
rect 2166 1454 2172 1455
rect 2232 1432 2234 1458
rect 2238 1455 2239 1459
rect 2243 1455 2244 1459
rect 2302 1459 2303 1463
rect 2307 1459 2308 1463
rect 2312 1460 2314 1469
rect 2322 1463 2328 1464
rect 2302 1458 2308 1459
rect 2310 1459 2316 1460
rect 2238 1454 2244 1455
rect 2304 1432 2306 1458
rect 2310 1455 2311 1459
rect 2315 1455 2316 1459
rect 2322 1459 2323 1463
rect 2327 1459 2328 1463
rect 2360 1460 2362 1469
rect 2384 1464 2386 1530
rect 2406 1528 2407 1532
rect 2411 1528 2412 1532
rect 2406 1527 2412 1528
rect 2408 1475 2410 1527
rect 2407 1474 2411 1475
rect 2407 1469 2411 1470
rect 2382 1463 2388 1464
rect 2322 1458 2328 1459
rect 2358 1459 2364 1460
rect 2310 1454 2316 1455
rect 1238 1431 1244 1432
rect 1278 1431 1284 1432
rect 1386 1431 1392 1432
rect 1238 1427 1239 1431
rect 1243 1427 1244 1431
rect 1238 1426 1244 1427
rect 1386 1427 1387 1431
rect 1391 1427 1392 1431
rect 1386 1426 1392 1427
rect 1458 1431 1464 1432
rect 1458 1427 1459 1431
rect 1463 1427 1464 1431
rect 1458 1426 1464 1427
rect 1574 1431 1580 1432
rect 1574 1427 1575 1431
rect 1579 1427 1580 1431
rect 1574 1426 1580 1427
rect 1678 1431 1684 1432
rect 1678 1427 1679 1431
rect 1683 1427 1684 1431
rect 1678 1426 1684 1427
rect 1942 1431 1948 1432
rect 1942 1427 1943 1431
rect 1947 1427 1948 1431
rect 1942 1426 1948 1427
rect 2022 1431 2028 1432
rect 2022 1427 2023 1431
rect 2027 1427 2028 1431
rect 2022 1426 2028 1427
rect 2094 1431 2100 1432
rect 2094 1427 2095 1431
rect 2099 1427 2100 1431
rect 2094 1426 2100 1427
rect 2158 1431 2164 1432
rect 2158 1427 2159 1431
rect 2163 1427 2164 1431
rect 2158 1426 2164 1427
rect 2230 1431 2236 1432
rect 2230 1427 2231 1431
rect 2235 1427 2236 1431
rect 2230 1426 2236 1427
rect 2302 1431 2308 1432
rect 2302 1427 2303 1431
rect 2307 1427 2308 1431
rect 2302 1426 2308 1427
rect 1022 1424 1028 1425
rect 1022 1420 1023 1424
rect 1027 1420 1028 1424
rect 1022 1419 1028 1420
rect 1086 1424 1092 1425
rect 1086 1420 1087 1424
rect 1091 1420 1092 1424
rect 1086 1419 1092 1420
rect 1150 1424 1156 1425
rect 1150 1420 1151 1424
rect 1155 1420 1156 1424
rect 1150 1419 1156 1420
rect 1190 1424 1196 1425
rect 1190 1420 1191 1424
rect 1195 1420 1196 1424
rect 1190 1419 1196 1420
rect 1024 1415 1026 1419
rect 1088 1415 1090 1419
rect 1152 1415 1154 1419
rect 1192 1415 1194 1419
rect 1240 1415 1242 1426
rect 1278 1419 1284 1420
rect 1278 1415 1279 1419
rect 1283 1415 1284 1419
rect 1023 1414 1027 1415
rect 1023 1409 1027 1410
rect 1087 1414 1091 1415
rect 1087 1409 1091 1410
rect 1151 1414 1155 1415
rect 1151 1409 1155 1410
rect 1191 1414 1195 1415
rect 1191 1409 1195 1410
rect 1239 1414 1243 1415
rect 1278 1414 1284 1415
rect 1239 1409 1243 1410
rect 1022 1408 1028 1409
rect 1022 1404 1023 1408
rect 1027 1404 1028 1408
rect 1022 1403 1028 1404
rect 1240 1402 1242 1409
rect 1280 1407 1282 1414
rect 1302 1412 1308 1413
rect 1302 1408 1303 1412
rect 1307 1408 1308 1412
rect 1302 1407 1308 1408
rect 1374 1412 1380 1413
rect 1374 1408 1375 1412
rect 1379 1408 1380 1412
rect 1374 1407 1380 1408
rect 1279 1406 1283 1407
rect 1238 1401 1244 1402
rect 1279 1401 1283 1402
rect 1303 1406 1307 1407
rect 1303 1401 1307 1402
rect 1343 1406 1347 1407
rect 1343 1401 1347 1402
rect 1375 1406 1379 1407
rect 1375 1401 1379 1402
rect 1399 1406 1403 1407
rect 1399 1401 1403 1402
rect 1238 1397 1239 1401
rect 1243 1397 1244 1401
rect 1238 1396 1244 1397
rect 1014 1395 1020 1396
rect 1014 1391 1015 1395
rect 1019 1391 1020 1395
rect 1280 1394 1282 1401
rect 1302 1400 1308 1401
rect 1302 1396 1303 1400
rect 1307 1396 1308 1400
rect 1302 1395 1308 1396
rect 1342 1400 1348 1401
rect 1342 1396 1343 1400
rect 1347 1396 1348 1400
rect 1342 1395 1348 1396
rect 1398 1400 1404 1401
rect 1398 1396 1399 1400
rect 1403 1396 1404 1400
rect 1398 1395 1404 1396
rect 1014 1390 1020 1391
rect 1278 1393 1284 1394
rect 1278 1389 1279 1393
rect 1283 1389 1284 1393
rect 1278 1388 1284 1389
rect 966 1387 972 1388
rect 966 1383 967 1387
rect 971 1383 972 1387
rect 966 1382 972 1383
rect 1038 1387 1044 1388
rect 1038 1383 1039 1387
rect 1043 1383 1044 1387
rect 1038 1382 1044 1383
rect 1238 1384 1244 1385
rect 878 1361 884 1362
rect 878 1357 879 1361
rect 883 1357 884 1361
rect 878 1356 884 1357
rect 950 1361 956 1362
rect 950 1357 951 1361
rect 955 1357 956 1361
rect 950 1356 956 1357
rect 968 1356 970 1382
rect 1022 1361 1028 1362
rect 1022 1357 1023 1361
rect 1027 1357 1028 1361
rect 1022 1356 1028 1357
rect 1040 1356 1042 1382
rect 1238 1380 1239 1384
rect 1243 1380 1244 1384
rect 1238 1379 1244 1380
rect 1350 1379 1356 1380
rect 816 1343 818 1356
rect 838 1355 844 1356
rect 838 1351 839 1355
rect 843 1351 844 1355
rect 838 1350 844 1351
rect 866 1355 872 1356
rect 866 1351 867 1355
rect 871 1351 872 1355
rect 866 1350 872 1351
rect 815 1342 819 1343
rect 815 1337 819 1338
rect 839 1342 843 1343
rect 839 1337 843 1338
rect 782 1331 788 1332
rect 750 1326 756 1327
rect 758 1327 764 1328
rect 670 1322 676 1323
rect 752 1300 754 1326
rect 758 1323 759 1327
rect 763 1323 764 1327
rect 782 1327 783 1331
rect 787 1327 788 1331
rect 840 1328 842 1337
rect 782 1326 788 1327
rect 838 1327 844 1328
rect 758 1322 764 1323
rect 838 1323 839 1327
rect 843 1323 844 1327
rect 838 1322 844 1323
rect 868 1300 870 1350
rect 880 1343 882 1356
rect 952 1343 954 1356
rect 966 1355 972 1356
rect 966 1351 967 1355
rect 971 1351 972 1355
rect 966 1350 972 1351
rect 1024 1343 1026 1356
rect 1038 1355 1044 1356
rect 1038 1351 1039 1355
rect 1043 1351 1044 1355
rect 1038 1350 1044 1351
rect 1240 1343 1242 1379
rect 1278 1376 1284 1377
rect 1278 1372 1279 1376
rect 1283 1372 1284 1376
rect 1350 1375 1351 1379
rect 1355 1375 1356 1379
rect 1350 1374 1356 1375
rect 1278 1371 1284 1372
rect 879 1342 883 1343
rect 879 1337 883 1338
rect 919 1342 923 1343
rect 919 1337 923 1338
rect 951 1342 955 1343
rect 951 1337 955 1338
rect 1007 1342 1011 1343
rect 1007 1337 1011 1338
rect 1023 1342 1027 1343
rect 1023 1337 1027 1338
rect 1095 1342 1099 1343
rect 1095 1337 1099 1338
rect 1239 1342 1243 1343
rect 1239 1337 1243 1338
rect 910 1331 916 1332
rect 910 1327 911 1331
rect 915 1327 916 1331
rect 920 1328 922 1337
rect 998 1331 1004 1332
rect 910 1326 916 1327
rect 918 1327 924 1328
rect 912 1300 914 1326
rect 918 1323 919 1327
rect 923 1323 924 1327
rect 998 1327 999 1331
rect 1003 1327 1004 1331
rect 1008 1328 1010 1337
rect 1086 1331 1092 1332
rect 998 1326 1004 1327
rect 1006 1327 1012 1328
rect 918 1322 924 1323
rect 1000 1300 1002 1326
rect 1006 1323 1007 1327
rect 1011 1323 1012 1327
rect 1086 1327 1087 1331
rect 1091 1327 1092 1331
rect 1096 1328 1098 1337
rect 1106 1331 1112 1332
rect 1086 1326 1092 1327
rect 1094 1327 1100 1328
rect 1006 1322 1012 1323
rect 1088 1300 1090 1326
rect 1094 1323 1095 1327
rect 1099 1323 1100 1327
rect 1106 1327 1107 1331
rect 1111 1327 1112 1331
rect 1106 1326 1112 1327
rect 1094 1322 1100 1323
rect 350 1299 356 1300
rect 350 1295 351 1299
rect 355 1295 356 1299
rect 350 1294 356 1295
rect 398 1299 404 1300
rect 398 1295 399 1299
rect 403 1295 404 1299
rect 398 1294 404 1295
rect 486 1299 492 1300
rect 486 1295 487 1299
rect 491 1295 492 1299
rect 486 1294 492 1295
rect 542 1299 548 1300
rect 542 1295 543 1299
rect 547 1295 548 1299
rect 542 1294 548 1295
rect 662 1299 668 1300
rect 662 1295 663 1299
rect 667 1295 668 1299
rect 662 1294 668 1295
rect 750 1299 756 1300
rect 750 1295 751 1299
rect 755 1295 756 1299
rect 750 1294 756 1295
rect 866 1299 872 1300
rect 866 1295 867 1299
rect 871 1295 872 1299
rect 866 1294 872 1295
rect 910 1299 916 1300
rect 910 1295 911 1299
rect 915 1295 916 1299
rect 910 1294 916 1295
rect 998 1299 1004 1300
rect 998 1295 999 1299
rect 1003 1295 1004 1299
rect 998 1294 1004 1295
rect 1086 1299 1092 1300
rect 1086 1295 1087 1299
rect 1091 1295 1092 1299
rect 1086 1294 1092 1295
rect 254 1280 260 1281
rect 254 1276 255 1280
rect 259 1276 260 1280
rect 254 1275 260 1276
rect 326 1280 332 1281
rect 326 1276 327 1280
rect 331 1276 332 1280
rect 326 1275 332 1276
rect 406 1280 412 1281
rect 406 1276 407 1280
rect 411 1276 412 1280
rect 406 1275 412 1276
rect 494 1280 500 1281
rect 494 1276 495 1280
rect 499 1276 500 1280
rect 494 1275 500 1276
rect 256 1271 258 1275
rect 328 1271 330 1275
rect 408 1271 410 1275
rect 496 1271 498 1275
rect 247 1270 251 1271
rect 247 1265 251 1266
rect 255 1270 259 1271
rect 255 1265 259 1266
rect 327 1270 331 1271
rect 327 1265 331 1266
rect 407 1270 411 1271
rect 407 1265 411 1266
rect 415 1270 419 1271
rect 415 1265 419 1266
rect 495 1270 499 1271
rect 495 1265 499 1266
rect 503 1270 507 1271
rect 503 1265 507 1266
rect 246 1264 252 1265
rect 246 1260 247 1264
rect 251 1260 252 1264
rect 246 1259 252 1260
rect 326 1264 332 1265
rect 326 1260 327 1264
rect 331 1260 332 1264
rect 326 1259 332 1260
rect 414 1264 420 1265
rect 414 1260 415 1264
rect 419 1260 420 1264
rect 414 1259 420 1260
rect 502 1264 508 1265
rect 502 1260 503 1264
rect 507 1260 508 1264
rect 502 1259 508 1260
rect 190 1243 196 1244
rect 110 1240 116 1241
rect 110 1236 111 1240
rect 115 1236 116 1240
rect 190 1239 191 1243
rect 195 1239 196 1243
rect 190 1238 196 1239
rect 238 1243 244 1244
rect 238 1239 239 1243
rect 243 1239 244 1243
rect 238 1238 244 1239
rect 110 1235 116 1236
rect 112 1195 114 1235
rect 134 1217 140 1218
rect 134 1213 135 1217
rect 139 1213 140 1217
rect 134 1212 140 1213
rect 174 1217 180 1218
rect 174 1213 175 1217
rect 179 1213 180 1217
rect 174 1212 180 1213
rect 192 1212 194 1238
rect 422 1235 428 1236
rect 422 1231 423 1235
rect 427 1231 428 1235
rect 422 1230 428 1231
rect 246 1217 252 1218
rect 246 1213 247 1217
rect 251 1213 252 1217
rect 246 1212 252 1213
rect 326 1217 332 1218
rect 326 1213 327 1217
rect 331 1213 332 1217
rect 326 1212 332 1213
rect 414 1217 420 1218
rect 414 1213 415 1217
rect 419 1213 420 1217
rect 414 1212 420 1213
rect 424 1212 426 1230
rect 502 1217 508 1218
rect 502 1213 503 1217
rect 507 1213 508 1217
rect 502 1212 508 1213
rect 544 1212 546 1294
rect 582 1280 588 1281
rect 582 1276 583 1280
rect 587 1276 588 1280
rect 582 1275 588 1276
rect 670 1280 676 1281
rect 670 1276 671 1280
rect 675 1276 676 1280
rect 670 1275 676 1276
rect 758 1280 764 1281
rect 758 1276 759 1280
rect 763 1276 764 1280
rect 758 1275 764 1276
rect 838 1280 844 1281
rect 838 1276 839 1280
rect 843 1276 844 1280
rect 838 1275 844 1276
rect 918 1280 924 1281
rect 918 1276 919 1280
rect 923 1276 924 1280
rect 918 1275 924 1276
rect 1006 1280 1012 1281
rect 1006 1276 1007 1280
rect 1011 1276 1012 1280
rect 1006 1275 1012 1276
rect 1094 1280 1100 1281
rect 1094 1276 1095 1280
rect 1099 1276 1100 1280
rect 1094 1275 1100 1276
rect 584 1271 586 1275
rect 672 1271 674 1275
rect 760 1271 762 1275
rect 840 1271 842 1275
rect 920 1271 922 1275
rect 1008 1271 1010 1275
rect 1096 1271 1098 1275
rect 583 1270 587 1271
rect 583 1265 587 1266
rect 591 1270 595 1271
rect 591 1265 595 1266
rect 671 1270 675 1271
rect 671 1265 675 1266
rect 743 1270 747 1271
rect 743 1265 747 1266
rect 759 1270 763 1271
rect 759 1265 763 1266
rect 815 1270 819 1271
rect 815 1265 819 1266
rect 839 1270 843 1271
rect 839 1265 843 1266
rect 879 1270 883 1271
rect 879 1265 883 1266
rect 919 1270 923 1271
rect 919 1265 923 1266
rect 943 1270 947 1271
rect 943 1265 947 1266
rect 1007 1270 1011 1271
rect 1007 1265 1011 1266
rect 1071 1270 1075 1271
rect 1071 1265 1075 1266
rect 1095 1270 1099 1271
rect 1095 1265 1099 1266
rect 590 1264 596 1265
rect 590 1260 591 1264
rect 595 1260 596 1264
rect 590 1259 596 1260
rect 670 1264 676 1265
rect 670 1260 671 1264
rect 675 1260 676 1264
rect 670 1259 676 1260
rect 742 1264 748 1265
rect 742 1260 743 1264
rect 747 1260 748 1264
rect 742 1259 748 1260
rect 814 1264 820 1265
rect 814 1260 815 1264
rect 819 1260 820 1264
rect 814 1259 820 1260
rect 878 1264 884 1265
rect 878 1260 879 1264
rect 883 1260 884 1264
rect 878 1259 884 1260
rect 942 1264 948 1265
rect 942 1260 943 1264
rect 947 1260 948 1264
rect 942 1259 948 1260
rect 1006 1264 1012 1265
rect 1006 1260 1007 1264
rect 1011 1260 1012 1264
rect 1006 1259 1012 1260
rect 1070 1264 1076 1265
rect 1070 1260 1071 1264
rect 1075 1260 1076 1264
rect 1070 1259 1076 1260
rect 1108 1244 1110 1326
rect 1240 1305 1242 1337
rect 1280 1335 1282 1371
rect 1302 1353 1308 1354
rect 1302 1349 1303 1353
rect 1307 1349 1308 1353
rect 1302 1348 1308 1349
rect 1342 1353 1348 1354
rect 1342 1349 1343 1353
rect 1347 1349 1348 1353
rect 1342 1348 1348 1349
rect 1352 1348 1354 1374
rect 1398 1353 1404 1354
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1398 1348 1404 1349
rect 1460 1348 1462 1426
rect 2094 1423 2100 1424
rect 2094 1419 2095 1423
rect 2099 1419 2100 1423
rect 2094 1418 2100 1419
rect 1478 1412 1484 1413
rect 1478 1408 1479 1412
rect 1483 1408 1484 1412
rect 1478 1407 1484 1408
rect 1582 1412 1588 1413
rect 1582 1408 1583 1412
rect 1587 1408 1588 1412
rect 1582 1407 1588 1408
rect 1686 1412 1692 1413
rect 1686 1408 1687 1412
rect 1691 1408 1692 1412
rect 1686 1407 1692 1408
rect 1782 1412 1788 1413
rect 1782 1408 1783 1412
rect 1787 1408 1788 1412
rect 1782 1407 1788 1408
rect 1870 1412 1876 1413
rect 1870 1408 1871 1412
rect 1875 1408 1876 1412
rect 1870 1407 1876 1408
rect 1950 1412 1956 1413
rect 1950 1408 1951 1412
rect 1955 1408 1956 1412
rect 1950 1407 1956 1408
rect 2030 1412 2036 1413
rect 2030 1408 2031 1412
rect 2035 1408 2036 1412
rect 2030 1407 2036 1408
rect 1471 1406 1475 1407
rect 1471 1401 1475 1402
rect 1479 1406 1483 1407
rect 1479 1401 1483 1402
rect 1551 1406 1555 1407
rect 1551 1401 1555 1402
rect 1583 1406 1587 1407
rect 1583 1401 1587 1402
rect 1639 1406 1643 1407
rect 1639 1401 1643 1402
rect 1687 1406 1691 1407
rect 1687 1401 1691 1402
rect 1727 1406 1731 1407
rect 1727 1401 1731 1402
rect 1783 1406 1787 1407
rect 1783 1401 1787 1402
rect 1815 1406 1819 1407
rect 1815 1401 1819 1402
rect 1871 1406 1875 1407
rect 1871 1401 1875 1402
rect 1903 1406 1907 1407
rect 1903 1401 1907 1402
rect 1951 1406 1955 1407
rect 1951 1401 1955 1402
rect 1991 1406 1995 1407
rect 1991 1401 1995 1402
rect 2031 1406 2035 1407
rect 2031 1401 2035 1402
rect 2071 1406 2075 1407
rect 2071 1401 2075 1402
rect 1470 1400 1476 1401
rect 1470 1396 1471 1400
rect 1475 1396 1476 1400
rect 1470 1395 1476 1396
rect 1550 1400 1556 1401
rect 1550 1396 1551 1400
rect 1555 1396 1556 1400
rect 1550 1395 1556 1396
rect 1638 1400 1644 1401
rect 1638 1396 1639 1400
rect 1643 1396 1644 1400
rect 1638 1395 1644 1396
rect 1726 1400 1732 1401
rect 1726 1396 1727 1400
rect 1731 1396 1732 1400
rect 1726 1395 1732 1396
rect 1814 1400 1820 1401
rect 1814 1396 1815 1400
rect 1819 1396 1820 1400
rect 1814 1395 1820 1396
rect 1902 1400 1908 1401
rect 1902 1396 1903 1400
rect 1907 1396 1908 1400
rect 1902 1395 1908 1396
rect 1990 1400 1996 1401
rect 1990 1396 1991 1400
rect 1995 1396 1996 1400
rect 1990 1395 1996 1396
rect 2070 1400 2076 1401
rect 2070 1396 2071 1400
rect 2075 1396 2076 1400
rect 2070 1395 2076 1396
rect 1574 1379 1580 1380
rect 1574 1375 1575 1379
rect 1579 1375 1580 1379
rect 1574 1374 1580 1375
rect 1926 1379 1932 1380
rect 1926 1375 1927 1379
rect 1931 1375 1932 1379
rect 1926 1374 1932 1375
rect 1494 1371 1500 1372
rect 1494 1367 1495 1371
rect 1499 1367 1500 1371
rect 1494 1366 1500 1367
rect 1470 1353 1476 1354
rect 1470 1349 1471 1353
rect 1475 1349 1476 1353
rect 1470 1348 1476 1349
rect 1496 1348 1498 1366
rect 1550 1353 1556 1354
rect 1550 1349 1551 1353
rect 1555 1349 1556 1353
rect 1550 1348 1556 1349
rect 1304 1335 1306 1348
rect 1344 1335 1346 1348
rect 1350 1347 1356 1348
rect 1350 1343 1351 1347
rect 1355 1343 1356 1347
rect 1350 1342 1356 1343
rect 1400 1335 1402 1348
rect 1458 1347 1464 1348
rect 1458 1343 1459 1347
rect 1463 1343 1464 1347
rect 1458 1342 1464 1343
rect 1472 1335 1474 1348
rect 1494 1347 1500 1348
rect 1494 1343 1495 1347
rect 1499 1343 1500 1347
rect 1494 1342 1500 1343
rect 1552 1335 1554 1348
rect 1279 1334 1283 1335
rect 1279 1329 1283 1330
rect 1303 1334 1307 1335
rect 1303 1329 1307 1330
rect 1343 1334 1347 1335
rect 1343 1329 1347 1330
rect 1399 1334 1403 1335
rect 1399 1329 1403 1330
rect 1447 1334 1451 1335
rect 1447 1329 1451 1330
rect 1471 1334 1475 1335
rect 1471 1329 1475 1330
rect 1487 1334 1491 1335
rect 1487 1329 1491 1330
rect 1527 1334 1531 1335
rect 1527 1329 1531 1330
rect 1551 1334 1555 1335
rect 1551 1329 1555 1330
rect 1567 1334 1571 1335
rect 1567 1329 1571 1330
rect 1238 1304 1244 1305
rect 1238 1300 1239 1304
rect 1243 1300 1244 1304
rect 1238 1299 1244 1300
rect 1280 1297 1282 1329
rect 1448 1320 1450 1329
rect 1488 1320 1490 1329
rect 1502 1327 1508 1328
rect 1502 1323 1503 1327
rect 1507 1323 1508 1327
rect 1502 1322 1508 1323
rect 1446 1319 1452 1320
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1486 1319 1492 1320
rect 1486 1315 1487 1319
rect 1491 1315 1492 1319
rect 1486 1314 1492 1315
rect 1278 1296 1284 1297
rect 1278 1292 1279 1296
rect 1283 1292 1284 1296
rect 1504 1292 1506 1322
rect 1528 1320 1530 1329
rect 1542 1327 1548 1328
rect 1542 1323 1543 1327
rect 1547 1323 1548 1327
rect 1542 1322 1548 1323
rect 1526 1319 1532 1320
rect 1526 1315 1527 1319
rect 1531 1315 1532 1319
rect 1526 1314 1532 1315
rect 1544 1292 1546 1322
rect 1568 1320 1570 1329
rect 1576 1328 1578 1374
rect 1746 1371 1752 1372
rect 1746 1367 1747 1371
rect 1751 1367 1752 1371
rect 1746 1366 1752 1367
rect 1638 1353 1644 1354
rect 1638 1349 1639 1353
rect 1643 1349 1644 1353
rect 1638 1348 1644 1349
rect 1726 1353 1732 1354
rect 1726 1349 1727 1353
rect 1731 1349 1732 1353
rect 1726 1348 1732 1349
rect 1748 1348 1750 1366
rect 1928 1356 1930 1374
rect 1926 1355 1932 1356
rect 1814 1353 1820 1354
rect 1814 1349 1815 1353
rect 1819 1349 1820 1353
rect 1814 1348 1820 1349
rect 1902 1353 1908 1354
rect 1902 1349 1903 1353
rect 1907 1349 1908 1353
rect 1926 1351 1927 1355
rect 1931 1351 1932 1355
rect 1926 1350 1932 1351
rect 1990 1353 1996 1354
rect 1902 1348 1908 1349
rect 1990 1349 1991 1353
rect 1995 1349 1996 1353
rect 1990 1348 1996 1349
rect 2070 1353 2076 1354
rect 2070 1349 2071 1353
rect 2075 1349 2076 1353
rect 2070 1348 2076 1349
rect 2096 1348 2098 1418
rect 2102 1412 2108 1413
rect 2102 1408 2103 1412
rect 2107 1408 2108 1412
rect 2102 1407 2108 1408
rect 2166 1412 2172 1413
rect 2166 1408 2167 1412
rect 2171 1408 2172 1412
rect 2166 1407 2172 1408
rect 2238 1412 2244 1413
rect 2238 1408 2239 1412
rect 2243 1408 2244 1412
rect 2238 1407 2244 1408
rect 2310 1412 2316 1413
rect 2310 1408 2311 1412
rect 2315 1408 2316 1412
rect 2310 1407 2316 1408
rect 2103 1406 2107 1407
rect 2103 1401 2107 1402
rect 2151 1406 2155 1407
rect 2151 1401 2155 1402
rect 2167 1406 2171 1407
rect 2167 1401 2171 1402
rect 2223 1406 2227 1407
rect 2223 1401 2227 1402
rect 2239 1406 2243 1407
rect 2239 1401 2243 1402
rect 2303 1406 2307 1407
rect 2303 1401 2307 1402
rect 2311 1406 2315 1407
rect 2311 1401 2315 1402
rect 2150 1400 2156 1401
rect 2150 1396 2151 1400
rect 2155 1396 2156 1400
rect 2150 1395 2156 1396
rect 2222 1400 2228 1401
rect 2222 1396 2223 1400
rect 2227 1396 2228 1400
rect 2222 1395 2228 1396
rect 2302 1400 2308 1401
rect 2302 1396 2303 1400
rect 2307 1396 2308 1400
rect 2302 1395 2308 1396
rect 2324 1388 2326 1458
rect 2358 1455 2359 1459
rect 2363 1455 2364 1459
rect 2382 1459 2383 1463
rect 2387 1459 2388 1463
rect 2382 1458 2388 1459
rect 2358 1454 2364 1455
rect 2408 1437 2410 1469
rect 2406 1436 2412 1437
rect 2406 1432 2407 1436
rect 2411 1432 2412 1436
rect 2406 1431 2412 1432
rect 2406 1419 2412 1420
rect 2406 1415 2407 1419
rect 2411 1415 2412 1419
rect 2406 1414 2412 1415
rect 2358 1412 2364 1413
rect 2358 1408 2359 1412
rect 2363 1408 2364 1412
rect 2358 1407 2364 1408
rect 2408 1407 2410 1414
rect 2359 1406 2363 1407
rect 2359 1401 2363 1402
rect 2407 1406 2411 1407
rect 2407 1401 2411 1402
rect 2358 1400 2364 1401
rect 2358 1396 2359 1400
rect 2363 1396 2364 1400
rect 2358 1395 2364 1396
rect 2408 1394 2410 1401
rect 2406 1393 2412 1394
rect 2406 1389 2407 1393
rect 2411 1389 2412 1393
rect 2406 1388 2412 1389
rect 2322 1387 2328 1388
rect 2322 1383 2323 1387
rect 2327 1383 2328 1387
rect 2322 1382 2328 1383
rect 2374 1379 2380 1380
rect 2374 1375 2375 1379
rect 2379 1375 2380 1379
rect 2374 1374 2380 1375
rect 2382 1379 2388 1380
rect 2382 1375 2383 1379
rect 2387 1375 2388 1379
rect 2382 1374 2388 1375
rect 2406 1376 2412 1377
rect 2190 1371 2196 1372
rect 2190 1367 2191 1371
rect 2195 1367 2196 1371
rect 2190 1366 2196 1367
rect 2150 1353 2156 1354
rect 2150 1349 2151 1353
rect 2155 1349 2156 1353
rect 2150 1348 2156 1349
rect 1640 1335 1642 1348
rect 1728 1335 1730 1348
rect 1746 1347 1752 1348
rect 1746 1343 1747 1347
rect 1751 1343 1752 1347
rect 1746 1342 1752 1343
rect 1816 1335 1818 1348
rect 1904 1335 1906 1348
rect 1992 1335 1994 1348
rect 2072 1335 2074 1348
rect 2094 1347 2100 1348
rect 2094 1343 2095 1347
rect 2099 1343 2100 1347
rect 2094 1342 2100 1343
rect 2152 1335 2154 1348
rect 1615 1334 1619 1335
rect 1615 1329 1619 1330
rect 1639 1334 1643 1335
rect 1639 1329 1643 1330
rect 1671 1334 1675 1335
rect 1671 1329 1675 1330
rect 1719 1334 1723 1335
rect 1719 1329 1723 1330
rect 1727 1334 1731 1335
rect 1727 1329 1731 1330
rect 1775 1334 1779 1335
rect 1775 1329 1779 1330
rect 1815 1334 1819 1335
rect 1815 1329 1819 1330
rect 1831 1334 1835 1335
rect 1831 1329 1835 1330
rect 1903 1334 1907 1335
rect 1903 1329 1907 1330
rect 1983 1334 1987 1335
rect 1983 1329 1987 1330
rect 1991 1334 1995 1335
rect 1991 1329 1995 1330
rect 2071 1334 2075 1335
rect 2071 1329 2075 1330
rect 2151 1334 2155 1335
rect 2151 1329 2155 1330
rect 2167 1334 2171 1335
rect 2167 1329 2171 1330
rect 1574 1327 1580 1328
rect 1574 1323 1575 1327
rect 1579 1323 1580 1327
rect 1574 1322 1580 1323
rect 1582 1323 1588 1324
rect 1566 1319 1572 1320
rect 1566 1315 1567 1319
rect 1571 1315 1572 1319
rect 1582 1319 1583 1323
rect 1587 1319 1588 1323
rect 1616 1320 1618 1329
rect 1662 1323 1668 1324
rect 1582 1318 1588 1319
rect 1614 1319 1620 1320
rect 1566 1314 1572 1315
rect 1584 1300 1586 1318
rect 1614 1315 1615 1319
rect 1619 1315 1620 1319
rect 1662 1319 1663 1323
rect 1667 1319 1668 1323
rect 1672 1320 1674 1329
rect 1710 1323 1716 1324
rect 1662 1318 1668 1319
rect 1670 1319 1676 1320
rect 1614 1314 1620 1315
rect 1582 1299 1588 1300
rect 1582 1295 1583 1299
rect 1587 1295 1588 1299
rect 1582 1294 1588 1295
rect 1664 1292 1666 1318
rect 1670 1315 1671 1319
rect 1675 1315 1676 1319
rect 1710 1319 1711 1323
rect 1715 1319 1716 1323
rect 1720 1320 1722 1329
rect 1730 1323 1736 1324
rect 1710 1318 1716 1319
rect 1718 1319 1724 1320
rect 1670 1314 1676 1315
rect 1712 1292 1714 1318
rect 1718 1315 1719 1319
rect 1723 1315 1724 1319
rect 1730 1319 1731 1323
rect 1735 1319 1736 1323
rect 1776 1320 1778 1329
rect 1822 1323 1828 1324
rect 1730 1318 1736 1319
rect 1774 1319 1780 1320
rect 1718 1314 1724 1315
rect 1732 1300 1734 1318
rect 1774 1315 1775 1319
rect 1779 1315 1780 1319
rect 1822 1319 1823 1323
rect 1827 1319 1828 1323
rect 1832 1320 1834 1329
rect 1894 1323 1900 1324
rect 1822 1318 1828 1319
rect 1830 1319 1836 1320
rect 1774 1314 1780 1315
rect 1730 1299 1736 1300
rect 1730 1295 1731 1299
rect 1735 1295 1736 1299
rect 1730 1294 1736 1295
rect 1824 1292 1826 1318
rect 1830 1315 1831 1319
rect 1835 1315 1836 1319
rect 1894 1319 1895 1323
rect 1899 1319 1900 1323
rect 1904 1320 1906 1329
rect 1962 1323 1968 1324
rect 1894 1318 1900 1319
rect 1902 1319 1908 1320
rect 1830 1314 1836 1315
rect 1896 1292 1898 1318
rect 1902 1315 1903 1319
rect 1907 1315 1908 1319
rect 1962 1319 1963 1323
rect 1967 1319 1968 1323
rect 1984 1320 1986 1329
rect 2062 1323 2068 1324
rect 1962 1318 1968 1319
rect 1982 1319 1988 1320
rect 1902 1314 1908 1315
rect 1964 1292 1966 1318
rect 1982 1315 1983 1319
rect 1987 1315 1988 1319
rect 2062 1319 2063 1323
rect 2067 1319 2068 1323
rect 2072 1320 2074 1329
rect 2158 1323 2164 1324
rect 2062 1318 2068 1319
rect 2070 1319 2076 1320
rect 1982 1314 1988 1315
rect 2064 1292 2066 1318
rect 2070 1315 2071 1319
rect 2075 1315 2076 1319
rect 2158 1319 2159 1323
rect 2163 1319 2164 1323
rect 2168 1320 2170 1329
rect 2192 1324 2194 1366
rect 2222 1353 2228 1354
rect 2222 1349 2223 1353
rect 2227 1349 2228 1353
rect 2222 1348 2228 1349
rect 2302 1353 2308 1354
rect 2302 1349 2303 1353
rect 2307 1349 2308 1353
rect 2302 1348 2308 1349
rect 2358 1353 2364 1354
rect 2358 1349 2359 1353
rect 2363 1349 2364 1353
rect 2358 1348 2364 1349
rect 2376 1348 2378 1374
rect 2224 1335 2226 1348
rect 2294 1347 2300 1348
rect 2294 1343 2295 1347
rect 2299 1343 2300 1347
rect 2294 1342 2300 1343
rect 2223 1334 2227 1335
rect 2223 1329 2227 1330
rect 2271 1334 2275 1335
rect 2271 1329 2275 1330
rect 2190 1323 2196 1324
rect 2158 1318 2164 1319
rect 2166 1319 2172 1320
rect 2070 1314 2076 1315
rect 2160 1292 2162 1318
rect 2166 1315 2167 1319
rect 2171 1315 2172 1319
rect 2190 1319 2191 1323
rect 2195 1319 2196 1323
rect 2272 1320 2274 1329
rect 2282 1323 2288 1324
rect 2190 1318 2196 1319
rect 2270 1319 2276 1320
rect 2166 1314 2172 1315
rect 2270 1315 2271 1319
rect 2275 1315 2276 1319
rect 2282 1319 2283 1323
rect 2287 1319 2288 1323
rect 2282 1318 2288 1319
rect 2270 1314 2276 1315
rect 1278 1291 1284 1292
rect 1502 1291 1508 1292
rect 1238 1287 1244 1288
rect 1238 1283 1239 1287
rect 1243 1283 1244 1287
rect 1502 1287 1503 1291
rect 1507 1287 1508 1291
rect 1502 1286 1508 1287
rect 1542 1291 1548 1292
rect 1542 1287 1543 1291
rect 1547 1287 1548 1291
rect 1542 1286 1548 1287
rect 1622 1291 1628 1292
rect 1622 1287 1623 1291
rect 1627 1287 1628 1291
rect 1622 1286 1628 1287
rect 1662 1291 1668 1292
rect 1662 1287 1663 1291
rect 1667 1287 1668 1291
rect 1662 1286 1668 1287
rect 1710 1291 1716 1292
rect 1710 1287 1711 1291
rect 1715 1287 1716 1291
rect 1710 1286 1716 1287
rect 1822 1291 1828 1292
rect 1822 1287 1823 1291
rect 1827 1287 1828 1291
rect 1822 1286 1828 1287
rect 1894 1291 1900 1292
rect 1894 1287 1895 1291
rect 1899 1287 1900 1291
rect 1894 1286 1900 1287
rect 1962 1291 1968 1292
rect 1962 1287 1963 1291
rect 1967 1287 1968 1291
rect 1962 1286 1968 1287
rect 2062 1291 2068 1292
rect 2062 1287 2063 1291
rect 2067 1287 2068 1291
rect 2062 1286 2068 1287
rect 2158 1291 2164 1292
rect 2158 1287 2159 1291
rect 2163 1287 2164 1291
rect 2158 1286 2164 1287
rect 1238 1282 1244 1283
rect 1240 1271 1242 1282
rect 1278 1279 1284 1280
rect 1278 1275 1279 1279
rect 1283 1275 1284 1279
rect 1278 1274 1284 1275
rect 1239 1270 1243 1271
rect 1239 1265 1243 1266
rect 1240 1258 1242 1265
rect 1280 1263 1282 1274
rect 1446 1272 1452 1273
rect 1446 1268 1447 1272
rect 1451 1268 1452 1272
rect 1446 1267 1452 1268
rect 1486 1272 1492 1273
rect 1486 1268 1487 1272
rect 1491 1268 1492 1272
rect 1486 1267 1492 1268
rect 1526 1272 1532 1273
rect 1526 1268 1527 1272
rect 1531 1268 1532 1272
rect 1526 1267 1532 1268
rect 1566 1272 1572 1273
rect 1566 1268 1567 1272
rect 1571 1268 1572 1272
rect 1566 1267 1572 1268
rect 1614 1272 1620 1273
rect 1614 1268 1615 1272
rect 1619 1268 1620 1272
rect 1614 1267 1620 1268
rect 1448 1263 1450 1267
rect 1488 1263 1490 1267
rect 1528 1263 1530 1267
rect 1568 1263 1570 1267
rect 1616 1263 1618 1267
rect 1279 1262 1283 1263
rect 1238 1257 1244 1258
rect 1279 1257 1283 1258
rect 1447 1262 1451 1263
rect 1447 1257 1451 1258
rect 1487 1262 1491 1263
rect 1487 1257 1491 1258
rect 1511 1262 1515 1263
rect 1511 1257 1515 1258
rect 1527 1262 1531 1263
rect 1527 1257 1531 1258
rect 1551 1262 1555 1263
rect 1551 1257 1555 1258
rect 1567 1262 1571 1263
rect 1567 1257 1571 1258
rect 1591 1262 1595 1263
rect 1591 1257 1595 1258
rect 1615 1262 1619 1263
rect 1615 1257 1619 1258
rect 1238 1253 1239 1257
rect 1243 1253 1244 1257
rect 1238 1252 1244 1253
rect 1280 1250 1282 1257
rect 1510 1256 1516 1257
rect 1510 1252 1511 1256
rect 1515 1252 1516 1256
rect 1510 1251 1516 1252
rect 1550 1256 1556 1257
rect 1550 1252 1551 1256
rect 1555 1252 1556 1256
rect 1550 1251 1556 1252
rect 1590 1256 1596 1257
rect 1590 1252 1591 1256
rect 1595 1252 1596 1256
rect 1590 1251 1596 1252
rect 1278 1249 1284 1250
rect 1278 1245 1279 1249
rect 1283 1245 1284 1249
rect 1278 1244 1284 1245
rect 606 1243 612 1244
rect 606 1239 607 1243
rect 611 1239 612 1243
rect 606 1238 612 1239
rect 662 1243 668 1244
rect 662 1239 663 1243
rect 667 1239 668 1243
rect 662 1238 668 1239
rect 678 1243 684 1244
rect 678 1239 679 1243
rect 683 1239 684 1243
rect 678 1238 684 1239
rect 958 1243 964 1244
rect 958 1239 959 1243
rect 963 1239 964 1243
rect 958 1238 964 1239
rect 1022 1243 1028 1244
rect 1022 1239 1023 1243
rect 1027 1239 1028 1243
rect 1022 1238 1028 1239
rect 1086 1243 1092 1244
rect 1086 1239 1087 1243
rect 1091 1239 1092 1243
rect 1086 1238 1092 1239
rect 1106 1243 1112 1244
rect 1106 1239 1107 1243
rect 1111 1239 1112 1243
rect 1106 1238 1112 1239
rect 1238 1240 1244 1241
rect 590 1217 596 1218
rect 590 1213 591 1217
rect 595 1213 596 1217
rect 590 1212 596 1213
rect 608 1212 610 1238
rect 664 1212 666 1238
rect 670 1217 676 1218
rect 670 1213 671 1217
rect 675 1213 676 1217
rect 670 1212 676 1213
rect 136 1195 138 1212
rect 158 1211 164 1212
rect 158 1207 159 1211
rect 163 1207 164 1211
rect 158 1206 164 1207
rect 111 1194 115 1195
rect 111 1189 115 1190
rect 135 1194 139 1195
rect 135 1189 139 1190
rect 112 1157 114 1189
rect 136 1180 138 1189
rect 134 1179 140 1180
rect 134 1175 135 1179
rect 139 1175 140 1179
rect 134 1174 140 1175
rect 110 1156 116 1157
rect 110 1152 111 1156
rect 115 1152 116 1156
rect 160 1152 162 1206
rect 176 1195 178 1212
rect 190 1211 196 1212
rect 190 1207 191 1211
rect 195 1207 196 1211
rect 190 1206 196 1207
rect 248 1195 250 1212
rect 328 1195 330 1212
rect 416 1195 418 1212
rect 422 1211 428 1212
rect 422 1207 423 1211
rect 427 1207 428 1211
rect 422 1206 428 1207
rect 504 1195 506 1212
rect 542 1211 548 1212
rect 542 1207 543 1211
rect 547 1207 548 1211
rect 542 1206 548 1207
rect 592 1195 594 1212
rect 606 1211 612 1212
rect 606 1207 607 1211
rect 611 1207 612 1211
rect 606 1206 612 1207
rect 662 1211 668 1212
rect 662 1207 663 1211
rect 667 1207 668 1211
rect 662 1206 668 1207
rect 672 1195 674 1212
rect 175 1194 179 1195
rect 175 1189 179 1190
rect 231 1194 235 1195
rect 231 1189 235 1190
rect 247 1194 251 1195
rect 247 1189 251 1190
rect 303 1194 307 1195
rect 303 1189 307 1190
rect 327 1194 331 1195
rect 327 1189 331 1190
rect 383 1194 387 1195
rect 383 1189 387 1190
rect 415 1194 419 1195
rect 415 1189 419 1190
rect 471 1194 475 1195
rect 471 1189 475 1190
rect 503 1194 507 1195
rect 503 1189 507 1190
rect 559 1194 563 1195
rect 559 1189 563 1190
rect 591 1194 595 1195
rect 591 1189 595 1190
rect 639 1194 643 1195
rect 639 1189 643 1190
rect 671 1194 675 1195
rect 671 1189 675 1190
rect 176 1180 178 1189
rect 190 1187 196 1188
rect 190 1183 191 1187
rect 195 1183 196 1187
rect 190 1182 196 1183
rect 222 1183 228 1184
rect 174 1179 180 1180
rect 174 1175 175 1179
rect 179 1175 180 1179
rect 174 1174 180 1175
rect 192 1152 194 1182
rect 222 1179 223 1183
rect 227 1179 228 1183
rect 232 1180 234 1189
rect 294 1183 300 1184
rect 222 1178 228 1179
rect 230 1179 236 1180
rect 224 1152 226 1178
rect 230 1175 231 1179
rect 235 1175 236 1179
rect 294 1179 295 1183
rect 299 1179 300 1183
rect 304 1180 306 1189
rect 374 1183 380 1184
rect 294 1178 300 1179
rect 302 1179 308 1180
rect 230 1174 236 1175
rect 296 1152 298 1178
rect 302 1175 303 1179
rect 307 1175 308 1179
rect 374 1179 375 1183
rect 379 1179 380 1183
rect 384 1180 386 1189
rect 398 1183 404 1184
rect 374 1178 380 1179
rect 382 1179 388 1180
rect 302 1174 308 1175
rect 376 1152 378 1178
rect 382 1175 383 1179
rect 387 1175 388 1179
rect 398 1179 399 1183
rect 403 1179 404 1183
rect 472 1180 474 1189
rect 550 1183 556 1184
rect 398 1178 404 1179
rect 470 1179 476 1180
rect 382 1174 388 1175
rect 110 1151 116 1152
rect 158 1151 164 1152
rect 158 1147 159 1151
rect 163 1147 164 1151
rect 158 1146 164 1147
rect 190 1151 196 1152
rect 190 1147 191 1151
rect 195 1147 196 1151
rect 190 1146 196 1147
rect 222 1151 228 1152
rect 222 1147 223 1151
rect 227 1147 228 1151
rect 222 1146 228 1147
rect 294 1151 300 1152
rect 294 1147 295 1151
rect 299 1147 300 1151
rect 294 1146 300 1147
rect 374 1151 380 1152
rect 374 1147 375 1151
rect 379 1147 380 1151
rect 374 1146 380 1147
rect 110 1139 116 1140
rect 110 1135 111 1139
rect 115 1135 116 1139
rect 110 1134 116 1135
rect 112 1127 114 1134
rect 134 1132 140 1133
rect 134 1128 135 1132
rect 139 1128 140 1132
rect 134 1127 140 1128
rect 174 1132 180 1133
rect 174 1128 175 1132
rect 179 1128 180 1132
rect 174 1127 180 1128
rect 230 1132 236 1133
rect 230 1128 231 1132
rect 235 1128 236 1132
rect 230 1127 236 1128
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 382 1132 388 1133
rect 382 1128 383 1132
rect 387 1128 388 1132
rect 382 1127 388 1128
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 135 1126 139 1127
rect 135 1121 139 1122
rect 175 1126 179 1127
rect 175 1121 179 1122
rect 215 1126 219 1127
rect 215 1121 219 1122
rect 231 1126 235 1127
rect 231 1121 235 1122
rect 303 1126 307 1127
rect 303 1121 307 1122
rect 383 1126 387 1127
rect 383 1121 387 1122
rect 391 1126 395 1127
rect 391 1121 395 1122
rect 112 1114 114 1121
rect 134 1120 140 1121
rect 134 1116 135 1120
rect 139 1116 140 1120
rect 134 1115 140 1116
rect 214 1120 220 1121
rect 214 1116 215 1120
rect 219 1116 220 1120
rect 214 1115 220 1116
rect 302 1120 308 1121
rect 302 1116 303 1120
rect 307 1116 308 1120
rect 302 1115 308 1116
rect 390 1120 396 1121
rect 390 1116 391 1120
rect 395 1116 396 1120
rect 390 1115 396 1116
rect 110 1113 116 1114
rect 110 1109 111 1113
rect 115 1109 116 1113
rect 110 1108 116 1109
rect 400 1108 402 1178
rect 470 1175 471 1179
rect 475 1175 476 1179
rect 550 1179 551 1183
rect 555 1179 556 1183
rect 560 1180 562 1189
rect 630 1183 636 1184
rect 550 1178 556 1179
rect 558 1179 564 1180
rect 470 1174 476 1175
rect 552 1152 554 1178
rect 558 1175 559 1179
rect 563 1175 564 1179
rect 630 1179 631 1183
rect 635 1179 636 1183
rect 640 1180 642 1189
rect 680 1184 682 1238
rect 902 1235 908 1236
rect 902 1231 903 1235
rect 907 1231 908 1235
rect 902 1230 908 1231
rect 742 1217 748 1218
rect 742 1213 743 1217
rect 747 1213 748 1217
rect 742 1212 748 1213
rect 814 1217 820 1218
rect 814 1213 815 1217
rect 819 1213 820 1217
rect 814 1212 820 1213
rect 878 1217 884 1218
rect 878 1213 879 1217
rect 883 1213 884 1217
rect 878 1212 884 1213
rect 904 1212 906 1230
rect 942 1217 948 1218
rect 942 1213 943 1217
rect 947 1213 948 1217
rect 942 1212 948 1213
rect 960 1212 962 1238
rect 1006 1217 1012 1218
rect 1006 1213 1007 1217
rect 1011 1213 1012 1217
rect 1006 1212 1012 1213
rect 1024 1212 1026 1238
rect 1070 1217 1076 1218
rect 1070 1213 1071 1217
rect 1075 1213 1076 1217
rect 1070 1212 1076 1213
rect 1088 1212 1090 1238
rect 1238 1236 1239 1240
rect 1243 1236 1244 1240
rect 1238 1235 1244 1236
rect 1558 1235 1564 1236
rect 744 1195 746 1212
rect 816 1195 818 1212
rect 880 1195 882 1212
rect 894 1211 900 1212
rect 894 1207 895 1211
rect 899 1207 900 1211
rect 894 1206 900 1207
rect 902 1211 908 1212
rect 902 1207 903 1211
rect 907 1207 908 1211
rect 902 1206 908 1207
rect 719 1194 723 1195
rect 719 1189 723 1190
rect 743 1194 747 1195
rect 743 1189 747 1190
rect 799 1194 803 1195
rect 799 1189 803 1190
rect 815 1194 819 1195
rect 815 1189 819 1190
rect 871 1194 875 1195
rect 871 1189 875 1190
rect 879 1194 883 1195
rect 879 1189 883 1190
rect 678 1183 684 1184
rect 630 1178 636 1179
rect 638 1179 644 1180
rect 558 1174 564 1175
rect 632 1152 634 1178
rect 638 1175 639 1179
rect 643 1175 644 1179
rect 678 1179 679 1183
rect 683 1179 684 1183
rect 720 1180 722 1189
rect 738 1183 744 1184
rect 678 1178 684 1179
rect 718 1179 724 1180
rect 638 1174 644 1175
rect 718 1175 719 1179
rect 723 1175 724 1179
rect 738 1179 739 1183
rect 743 1179 744 1183
rect 800 1180 802 1189
rect 810 1183 816 1184
rect 738 1178 744 1179
rect 798 1179 804 1180
rect 718 1174 724 1175
rect 498 1151 504 1152
rect 498 1147 499 1151
rect 503 1147 504 1151
rect 498 1146 504 1147
rect 550 1151 556 1152
rect 550 1147 551 1151
rect 555 1147 556 1151
rect 550 1146 556 1147
rect 630 1151 636 1152
rect 630 1147 631 1151
rect 635 1147 636 1151
rect 630 1146 636 1147
rect 470 1132 476 1133
rect 470 1128 471 1132
rect 475 1128 476 1132
rect 470 1127 476 1128
rect 471 1126 475 1127
rect 471 1121 475 1122
rect 479 1126 483 1127
rect 479 1121 483 1122
rect 478 1120 484 1121
rect 478 1116 479 1120
rect 483 1116 484 1120
rect 478 1115 484 1116
rect 398 1107 404 1108
rect 398 1103 399 1107
rect 403 1103 404 1107
rect 398 1102 404 1103
rect 110 1096 116 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 112 1055 114 1091
rect 134 1073 140 1074
rect 134 1069 135 1073
rect 139 1069 140 1073
rect 134 1068 140 1069
rect 214 1073 220 1074
rect 214 1069 215 1073
rect 219 1069 220 1073
rect 214 1068 220 1069
rect 302 1073 308 1074
rect 302 1069 303 1073
rect 307 1069 308 1073
rect 302 1068 308 1069
rect 390 1073 396 1074
rect 390 1069 391 1073
rect 395 1069 396 1073
rect 390 1068 396 1069
rect 478 1073 484 1074
rect 478 1069 479 1073
rect 483 1069 484 1073
rect 478 1068 484 1069
rect 500 1068 502 1146
rect 558 1132 564 1133
rect 558 1128 559 1132
rect 563 1128 564 1132
rect 558 1127 564 1128
rect 638 1132 644 1133
rect 638 1128 639 1132
rect 643 1128 644 1132
rect 638 1127 644 1128
rect 718 1132 724 1133
rect 718 1128 719 1132
rect 723 1128 724 1132
rect 718 1127 724 1128
rect 559 1126 563 1127
rect 559 1121 563 1122
rect 639 1126 643 1127
rect 639 1121 643 1122
rect 711 1126 715 1127
rect 711 1121 715 1122
rect 719 1126 723 1127
rect 719 1121 723 1122
rect 558 1120 564 1121
rect 558 1116 559 1120
rect 563 1116 564 1120
rect 558 1115 564 1116
rect 638 1120 644 1121
rect 638 1116 639 1120
rect 643 1116 644 1120
rect 638 1115 644 1116
rect 710 1120 716 1121
rect 710 1116 711 1120
rect 715 1116 716 1120
rect 710 1115 716 1116
rect 740 1100 742 1178
rect 798 1175 799 1179
rect 803 1175 804 1179
rect 810 1179 811 1183
rect 815 1179 816 1183
rect 872 1180 874 1189
rect 882 1183 888 1184
rect 810 1178 816 1179
rect 870 1179 876 1180
rect 798 1174 804 1175
rect 812 1152 814 1178
rect 870 1175 871 1179
rect 875 1175 876 1179
rect 882 1179 883 1183
rect 887 1179 888 1183
rect 882 1178 888 1179
rect 870 1174 876 1175
rect 884 1152 886 1178
rect 896 1152 898 1206
rect 944 1195 946 1212
rect 958 1211 964 1212
rect 958 1207 959 1211
rect 963 1207 964 1211
rect 958 1206 964 1207
rect 1008 1195 1010 1212
rect 1022 1211 1028 1212
rect 1022 1207 1023 1211
rect 1027 1207 1028 1211
rect 1022 1206 1028 1207
rect 1072 1195 1074 1212
rect 1086 1211 1092 1212
rect 1086 1207 1087 1211
rect 1091 1207 1092 1211
rect 1086 1206 1092 1207
rect 1240 1195 1242 1235
rect 1278 1232 1284 1233
rect 1278 1228 1279 1232
rect 1283 1228 1284 1232
rect 1558 1231 1559 1235
rect 1563 1231 1564 1235
rect 1558 1230 1564 1231
rect 1598 1235 1604 1236
rect 1598 1231 1599 1235
rect 1603 1231 1604 1235
rect 1598 1230 1604 1231
rect 1278 1227 1284 1228
rect 935 1194 939 1195
rect 935 1189 939 1190
rect 943 1194 947 1195
rect 943 1189 947 1190
rect 991 1194 995 1195
rect 991 1189 995 1190
rect 1007 1194 1011 1195
rect 1007 1189 1011 1190
rect 1047 1194 1051 1195
rect 1047 1189 1051 1190
rect 1071 1194 1075 1195
rect 1071 1189 1075 1190
rect 1103 1194 1107 1195
rect 1103 1189 1107 1190
rect 1151 1194 1155 1195
rect 1151 1189 1155 1190
rect 1191 1194 1195 1195
rect 1191 1189 1195 1190
rect 1239 1194 1243 1195
rect 1280 1191 1282 1227
rect 1510 1209 1516 1210
rect 1510 1205 1511 1209
rect 1515 1205 1516 1209
rect 1510 1204 1516 1205
rect 1550 1209 1556 1210
rect 1550 1205 1551 1209
rect 1555 1205 1556 1209
rect 1550 1204 1556 1205
rect 1560 1204 1562 1230
rect 1590 1209 1596 1210
rect 1590 1205 1591 1209
rect 1595 1205 1596 1209
rect 1590 1204 1596 1205
rect 1600 1204 1602 1230
rect 1512 1191 1514 1204
rect 1552 1191 1554 1204
rect 1558 1203 1564 1204
rect 1558 1199 1559 1203
rect 1563 1199 1564 1203
rect 1558 1198 1564 1199
rect 1592 1191 1594 1204
rect 1598 1203 1604 1204
rect 1598 1199 1599 1203
rect 1603 1199 1604 1203
rect 1598 1198 1604 1199
rect 1615 1203 1621 1204
rect 1615 1199 1616 1203
rect 1620 1202 1621 1203
rect 1624 1202 1626 1286
rect 2142 1283 2148 1284
rect 2142 1279 2143 1283
rect 2147 1279 2148 1283
rect 2142 1278 2148 1279
rect 1670 1272 1676 1273
rect 1670 1268 1671 1272
rect 1675 1268 1676 1272
rect 1670 1267 1676 1268
rect 1718 1272 1724 1273
rect 1718 1268 1719 1272
rect 1723 1268 1724 1272
rect 1718 1267 1724 1268
rect 1774 1272 1780 1273
rect 1774 1268 1775 1272
rect 1779 1268 1780 1272
rect 1774 1267 1780 1268
rect 1830 1272 1836 1273
rect 1830 1268 1831 1272
rect 1835 1268 1836 1272
rect 1830 1267 1836 1268
rect 1902 1272 1908 1273
rect 1902 1268 1903 1272
rect 1907 1268 1908 1272
rect 1902 1267 1908 1268
rect 1982 1272 1988 1273
rect 1982 1268 1983 1272
rect 1987 1268 1988 1272
rect 1982 1267 1988 1268
rect 2070 1272 2076 1273
rect 2070 1268 2071 1272
rect 2075 1268 2076 1272
rect 2070 1267 2076 1268
rect 1672 1263 1674 1267
rect 1720 1263 1722 1267
rect 1776 1263 1778 1267
rect 1832 1263 1834 1267
rect 1904 1263 1906 1267
rect 1984 1263 1986 1267
rect 2072 1263 2074 1267
rect 1631 1262 1635 1263
rect 1631 1257 1635 1258
rect 1671 1262 1675 1263
rect 1671 1257 1675 1258
rect 1711 1262 1715 1263
rect 1711 1257 1715 1258
rect 1719 1262 1723 1263
rect 1719 1257 1723 1258
rect 1751 1262 1755 1263
rect 1751 1257 1755 1258
rect 1775 1262 1779 1263
rect 1775 1257 1779 1258
rect 1791 1262 1795 1263
rect 1791 1257 1795 1258
rect 1831 1262 1835 1263
rect 1831 1257 1835 1258
rect 1839 1262 1843 1263
rect 1839 1257 1843 1258
rect 1903 1262 1907 1263
rect 1903 1257 1907 1258
rect 1967 1262 1971 1263
rect 1967 1257 1971 1258
rect 1983 1262 1987 1263
rect 1983 1257 1987 1258
rect 2039 1262 2043 1263
rect 2039 1257 2043 1258
rect 2071 1262 2075 1263
rect 2071 1257 2075 1258
rect 2119 1262 2123 1263
rect 2119 1257 2123 1258
rect 1630 1256 1636 1257
rect 1630 1252 1631 1256
rect 1635 1252 1636 1256
rect 1630 1251 1636 1252
rect 1670 1256 1676 1257
rect 1670 1252 1671 1256
rect 1675 1252 1676 1256
rect 1670 1251 1676 1252
rect 1710 1256 1716 1257
rect 1710 1252 1711 1256
rect 1715 1252 1716 1256
rect 1710 1251 1716 1252
rect 1750 1256 1756 1257
rect 1750 1252 1751 1256
rect 1755 1252 1756 1256
rect 1750 1251 1756 1252
rect 1790 1256 1796 1257
rect 1790 1252 1791 1256
rect 1795 1252 1796 1256
rect 1790 1251 1796 1252
rect 1838 1256 1844 1257
rect 1838 1252 1839 1256
rect 1843 1252 1844 1256
rect 1838 1251 1844 1252
rect 1902 1256 1908 1257
rect 1902 1252 1903 1256
rect 1907 1252 1908 1256
rect 1902 1251 1908 1252
rect 1966 1256 1972 1257
rect 1966 1252 1967 1256
rect 1971 1252 1972 1256
rect 1966 1251 1972 1252
rect 2038 1256 2044 1257
rect 2038 1252 2039 1256
rect 2043 1252 2044 1256
rect 2038 1251 2044 1252
rect 2118 1256 2124 1257
rect 2118 1252 2119 1256
rect 2123 1252 2124 1256
rect 2118 1251 2124 1252
rect 1686 1235 1692 1236
rect 1686 1231 1687 1235
rect 1691 1231 1692 1235
rect 1686 1230 1692 1231
rect 1726 1235 1732 1236
rect 1726 1231 1727 1235
rect 1731 1231 1732 1235
rect 1726 1230 1732 1231
rect 1758 1235 1764 1236
rect 1758 1231 1759 1235
rect 1763 1231 1764 1235
rect 1758 1230 1764 1231
rect 1766 1235 1772 1236
rect 1766 1231 1767 1235
rect 1771 1231 1772 1235
rect 1766 1230 1772 1231
rect 1806 1235 1812 1236
rect 1806 1231 1807 1235
rect 1811 1231 1812 1235
rect 1806 1230 1812 1231
rect 2030 1235 2036 1236
rect 2030 1231 2031 1235
rect 2035 1231 2036 1235
rect 2030 1230 2036 1231
rect 1654 1227 1660 1228
rect 1654 1223 1655 1227
rect 1659 1223 1660 1227
rect 1654 1222 1660 1223
rect 1630 1209 1636 1210
rect 1630 1205 1631 1209
rect 1635 1205 1636 1209
rect 1630 1204 1636 1205
rect 1656 1204 1658 1222
rect 1670 1209 1676 1210
rect 1670 1205 1671 1209
rect 1675 1205 1676 1209
rect 1670 1204 1676 1205
rect 1688 1204 1690 1230
rect 1710 1209 1716 1210
rect 1710 1205 1711 1209
rect 1715 1205 1716 1209
rect 1710 1204 1716 1205
rect 1728 1204 1730 1230
rect 1750 1209 1756 1210
rect 1750 1205 1751 1209
rect 1755 1205 1756 1209
rect 1750 1204 1756 1205
rect 1760 1204 1762 1230
rect 1620 1200 1626 1202
rect 1620 1199 1621 1200
rect 1615 1198 1621 1199
rect 1632 1191 1634 1204
rect 1654 1203 1660 1204
rect 1654 1199 1655 1203
rect 1659 1199 1660 1203
rect 1654 1198 1660 1199
rect 1672 1191 1674 1204
rect 1686 1203 1692 1204
rect 1686 1199 1687 1203
rect 1691 1199 1692 1203
rect 1686 1198 1692 1199
rect 1712 1191 1714 1204
rect 1726 1203 1732 1204
rect 1726 1199 1727 1203
rect 1731 1199 1732 1203
rect 1726 1198 1732 1199
rect 1752 1191 1754 1204
rect 1758 1203 1764 1204
rect 1758 1199 1759 1203
rect 1763 1199 1764 1203
rect 1758 1198 1764 1199
rect 1239 1189 1243 1190
rect 1279 1190 1283 1191
rect 936 1180 938 1189
rect 982 1183 988 1184
rect 934 1179 940 1180
rect 934 1175 935 1179
rect 939 1175 940 1179
rect 982 1179 983 1183
rect 987 1179 988 1183
rect 992 1180 994 1189
rect 1038 1183 1044 1184
rect 982 1178 988 1179
rect 990 1179 996 1180
rect 934 1174 940 1175
rect 984 1152 986 1178
rect 990 1175 991 1179
rect 995 1175 996 1179
rect 1038 1179 1039 1183
rect 1043 1179 1044 1183
rect 1048 1180 1050 1189
rect 1094 1183 1100 1184
rect 1038 1178 1044 1179
rect 1046 1179 1052 1180
rect 990 1174 996 1175
rect 1040 1152 1042 1178
rect 1046 1175 1047 1179
rect 1051 1175 1052 1179
rect 1094 1179 1095 1183
rect 1099 1179 1100 1183
rect 1104 1180 1106 1189
rect 1142 1183 1148 1184
rect 1094 1178 1100 1179
rect 1102 1179 1108 1180
rect 1046 1174 1052 1175
rect 1096 1152 1098 1178
rect 1102 1175 1103 1179
rect 1107 1175 1108 1179
rect 1142 1179 1143 1183
rect 1147 1179 1148 1183
rect 1152 1180 1154 1189
rect 1192 1180 1194 1189
rect 1206 1187 1212 1188
rect 1206 1183 1207 1187
rect 1211 1183 1212 1187
rect 1206 1182 1212 1183
rect 1214 1183 1220 1184
rect 1142 1178 1148 1179
rect 1150 1179 1156 1180
rect 1102 1174 1108 1175
rect 1144 1152 1146 1178
rect 1150 1175 1151 1179
rect 1155 1175 1156 1179
rect 1150 1174 1156 1175
rect 1190 1179 1196 1180
rect 1190 1175 1191 1179
rect 1195 1175 1196 1179
rect 1190 1174 1196 1175
rect 1208 1152 1210 1182
rect 1214 1179 1215 1183
rect 1219 1179 1220 1183
rect 1214 1178 1220 1179
rect 810 1151 816 1152
rect 810 1147 811 1151
rect 815 1147 816 1151
rect 810 1146 816 1147
rect 882 1151 888 1152
rect 882 1147 883 1151
rect 887 1147 888 1151
rect 882 1146 888 1147
rect 894 1151 900 1152
rect 894 1147 895 1151
rect 899 1147 900 1151
rect 894 1146 900 1147
rect 982 1151 988 1152
rect 982 1147 983 1151
rect 987 1147 988 1151
rect 982 1146 988 1147
rect 1038 1151 1044 1152
rect 1038 1147 1039 1151
rect 1043 1147 1044 1151
rect 1038 1146 1044 1147
rect 1094 1151 1100 1152
rect 1094 1147 1095 1151
rect 1099 1147 1100 1151
rect 1094 1146 1100 1147
rect 1142 1151 1148 1152
rect 1142 1147 1143 1151
rect 1147 1147 1148 1151
rect 1142 1146 1148 1147
rect 1206 1151 1212 1152
rect 1206 1147 1207 1151
rect 1211 1147 1212 1151
rect 1206 1146 1212 1147
rect 1014 1143 1020 1144
rect 1014 1139 1015 1143
rect 1019 1139 1020 1143
rect 1014 1138 1020 1139
rect 798 1132 804 1133
rect 798 1128 799 1132
rect 803 1128 804 1132
rect 798 1127 804 1128
rect 870 1132 876 1133
rect 870 1128 871 1132
rect 875 1128 876 1132
rect 870 1127 876 1128
rect 934 1132 940 1133
rect 934 1128 935 1132
rect 939 1128 940 1132
rect 934 1127 940 1128
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 775 1126 779 1127
rect 775 1121 779 1122
rect 799 1126 803 1127
rect 799 1121 803 1122
rect 839 1126 843 1127
rect 839 1121 843 1122
rect 871 1126 875 1127
rect 871 1121 875 1122
rect 903 1126 907 1127
rect 903 1121 907 1122
rect 935 1126 939 1127
rect 935 1121 939 1122
rect 959 1126 963 1127
rect 959 1121 963 1122
rect 991 1126 995 1127
rect 991 1121 995 1122
rect 774 1120 780 1121
rect 774 1116 775 1120
rect 779 1116 780 1120
rect 774 1115 780 1116
rect 838 1120 844 1121
rect 838 1116 839 1120
rect 843 1116 844 1120
rect 838 1115 844 1116
rect 902 1120 908 1121
rect 902 1116 903 1120
rect 907 1116 908 1120
rect 902 1115 908 1116
rect 958 1120 964 1121
rect 958 1116 959 1120
rect 963 1116 964 1120
rect 958 1115 964 1116
rect 566 1099 572 1100
rect 566 1095 567 1099
rect 571 1095 572 1099
rect 566 1094 572 1095
rect 574 1099 580 1100
rect 574 1095 575 1099
rect 579 1095 580 1099
rect 574 1094 580 1095
rect 726 1099 732 1100
rect 726 1095 727 1099
rect 731 1095 732 1099
rect 726 1094 732 1095
rect 738 1099 744 1100
rect 738 1095 739 1099
rect 743 1095 744 1099
rect 738 1094 744 1095
rect 558 1073 564 1074
rect 558 1069 559 1073
rect 563 1069 564 1073
rect 558 1068 564 1069
rect 568 1068 570 1094
rect 136 1055 138 1068
rect 216 1055 218 1068
rect 266 1059 272 1060
rect 266 1055 267 1059
rect 271 1055 272 1059
rect 304 1055 306 1068
rect 392 1055 394 1068
rect 480 1055 482 1068
rect 498 1067 504 1068
rect 498 1063 499 1067
rect 503 1063 504 1067
rect 498 1062 504 1063
rect 560 1055 562 1068
rect 566 1067 572 1068
rect 566 1063 567 1067
rect 571 1063 572 1067
rect 566 1062 572 1063
rect 111 1054 115 1055
rect 111 1049 115 1050
rect 135 1054 139 1055
rect 135 1049 139 1050
rect 199 1054 203 1055
rect 199 1049 203 1050
rect 215 1054 219 1055
rect 215 1049 219 1050
rect 239 1054 243 1055
rect 266 1054 272 1055
rect 287 1054 291 1055
rect 239 1049 243 1050
rect 112 1017 114 1049
rect 200 1040 202 1049
rect 226 1043 232 1044
rect 198 1039 204 1040
rect 198 1035 199 1039
rect 203 1035 204 1039
rect 226 1039 227 1043
rect 231 1039 232 1043
rect 240 1040 242 1049
rect 226 1038 232 1039
rect 238 1039 244 1040
rect 198 1034 204 1035
rect 110 1016 116 1017
rect 110 1012 111 1016
rect 115 1012 116 1016
rect 110 1011 116 1012
rect 228 1010 230 1038
rect 238 1035 239 1039
rect 243 1035 244 1039
rect 238 1034 244 1035
rect 268 1020 270 1054
rect 287 1049 291 1050
rect 303 1054 307 1055
rect 303 1049 307 1050
rect 343 1054 347 1055
rect 343 1049 347 1050
rect 391 1054 395 1055
rect 391 1049 395 1050
rect 439 1054 443 1055
rect 439 1049 443 1050
rect 479 1054 483 1055
rect 479 1049 483 1050
rect 487 1054 491 1055
rect 487 1049 491 1050
rect 535 1054 539 1055
rect 535 1049 539 1050
rect 559 1054 563 1055
rect 559 1049 563 1050
rect 278 1043 284 1044
rect 278 1039 279 1043
rect 283 1039 284 1043
rect 288 1040 290 1049
rect 334 1043 340 1044
rect 278 1038 284 1039
rect 286 1039 292 1040
rect 266 1019 272 1020
rect 266 1015 267 1019
rect 271 1015 272 1019
rect 266 1014 272 1015
rect 280 1012 282 1038
rect 286 1035 287 1039
rect 291 1035 292 1039
rect 334 1039 335 1043
rect 339 1039 340 1043
rect 344 1040 346 1049
rect 382 1043 388 1044
rect 334 1038 340 1039
rect 342 1039 348 1040
rect 286 1034 292 1035
rect 336 1012 338 1038
rect 342 1035 343 1039
rect 347 1035 348 1039
rect 382 1039 383 1043
rect 387 1039 388 1043
rect 392 1040 394 1049
rect 406 1043 412 1044
rect 382 1038 388 1039
rect 390 1039 396 1040
rect 342 1034 348 1035
rect 384 1012 386 1038
rect 390 1035 391 1039
rect 395 1035 396 1039
rect 406 1039 407 1043
rect 411 1039 412 1043
rect 440 1040 442 1049
rect 478 1043 484 1044
rect 406 1038 412 1039
rect 438 1039 444 1040
rect 390 1034 396 1035
rect 234 1011 240 1012
rect 234 1010 235 1011
rect 228 1008 235 1010
rect 234 1007 235 1008
rect 239 1007 240 1011
rect 234 1006 240 1007
rect 278 1011 284 1012
rect 278 1007 279 1011
rect 283 1007 284 1011
rect 278 1006 284 1007
rect 334 1011 340 1012
rect 334 1007 335 1011
rect 339 1007 340 1011
rect 334 1006 340 1007
rect 382 1011 388 1012
rect 382 1007 383 1011
rect 387 1007 388 1011
rect 382 1006 388 1007
rect 110 999 116 1000
rect 110 995 111 999
rect 115 995 116 999
rect 110 994 116 995
rect 112 975 114 994
rect 198 992 204 993
rect 198 988 199 992
rect 203 988 204 992
rect 198 987 204 988
rect 238 992 244 993
rect 238 988 239 992
rect 243 988 244 992
rect 238 987 244 988
rect 286 992 292 993
rect 286 988 287 992
rect 291 988 292 992
rect 286 987 292 988
rect 342 992 348 993
rect 342 988 343 992
rect 347 988 348 992
rect 342 987 348 988
rect 390 992 396 993
rect 390 988 391 992
rect 395 988 396 992
rect 390 987 396 988
rect 200 975 202 987
rect 240 975 242 987
rect 288 975 290 987
rect 344 975 346 987
rect 392 975 394 987
rect 111 974 115 975
rect 111 969 115 970
rect 199 974 203 975
rect 199 969 203 970
rect 239 974 243 975
rect 239 969 243 970
rect 287 974 291 975
rect 287 969 291 970
rect 295 974 299 975
rect 295 969 299 970
rect 343 974 347 975
rect 343 969 347 970
rect 391 974 395 975
rect 391 969 395 970
rect 399 974 403 975
rect 399 969 403 970
rect 112 962 114 969
rect 294 968 300 969
rect 294 964 295 968
rect 299 964 300 968
rect 294 963 300 964
rect 342 968 348 969
rect 342 964 343 968
rect 347 964 348 968
rect 342 963 348 964
rect 398 968 404 969
rect 398 964 399 968
rect 403 964 404 968
rect 398 963 404 964
rect 110 961 116 962
rect 110 957 111 961
rect 115 957 116 961
rect 110 956 116 957
rect 408 956 410 1038
rect 438 1035 439 1039
rect 443 1035 444 1039
rect 478 1039 479 1043
rect 483 1039 484 1043
rect 488 1040 490 1049
rect 526 1043 532 1044
rect 478 1038 484 1039
rect 486 1039 492 1040
rect 438 1034 444 1035
rect 480 1012 482 1038
rect 486 1035 487 1039
rect 491 1035 492 1039
rect 526 1039 527 1043
rect 531 1039 532 1043
rect 536 1040 538 1049
rect 576 1048 578 1094
rect 638 1073 644 1074
rect 638 1069 639 1073
rect 643 1069 644 1073
rect 638 1068 644 1069
rect 710 1073 716 1074
rect 710 1069 711 1073
rect 715 1069 716 1073
rect 710 1068 716 1069
rect 728 1068 730 1094
rect 982 1091 988 1092
rect 982 1087 983 1091
rect 987 1087 988 1091
rect 982 1086 988 1087
rect 774 1073 780 1074
rect 774 1069 775 1073
rect 779 1069 780 1073
rect 774 1068 780 1069
rect 838 1073 844 1074
rect 838 1069 839 1073
rect 843 1069 844 1073
rect 838 1068 844 1069
rect 902 1073 908 1074
rect 902 1069 903 1073
rect 907 1069 908 1073
rect 902 1068 908 1069
rect 958 1073 964 1074
rect 958 1069 959 1073
rect 963 1069 964 1073
rect 958 1068 964 1069
rect 610 1067 616 1068
rect 610 1063 611 1067
rect 615 1063 616 1067
rect 610 1062 616 1063
rect 583 1054 587 1055
rect 583 1049 587 1050
rect 574 1047 580 1048
rect 574 1043 575 1047
rect 579 1043 580 1047
rect 574 1042 580 1043
rect 584 1040 586 1049
rect 526 1038 532 1039
rect 534 1039 540 1040
rect 486 1034 492 1035
rect 528 1012 530 1038
rect 534 1035 535 1039
rect 539 1035 540 1039
rect 534 1034 540 1035
rect 582 1039 588 1040
rect 582 1035 583 1039
rect 587 1035 588 1039
rect 582 1034 588 1035
rect 612 1012 614 1062
rect 640 1055 642 1068
rect 712 1055 714 1068
rect 726 1067 732 1068
rect 726 1063 727 1067
rect 731 1063 732 1067
rect 726 1062 732 1063
rect 776 1055 778 1068
rect 840 1055 842 1068
rect 904 1055 906 1068
rect 960 1055 962 1068
rect 631 1054 635 1055
rect 631 1049 635 1050
rect 639 1054 643 1055
rect 639 1049 643 1050
rect 679 1054 683 1055
rect 679 1049 683 1050
rect 711 1054 715 1055
rect 711 1049 715 1050
rect 727 1054 731 1055
rect 727 1049 731 1050
rect 775 1054 779 1055
rect 775 1049 779 1050
rect 783 1054 787 1055
rect 783 1049 787 1050
rect 839 1054 843 1055
rect 839 1049 843 1050
rect 895 1054 899 1055
rect 895 1049 899 1050
rect 903 1054 907 1055
rect 903 1049 907 1050
rect 959 1054 963 1055
rect 959 1049 963 1050
rect 622 1043 628 1044
rect 622 1039 623 1043
rect 627 1039 628 1043
rect 632 1040 634 1049
rect 680 1040 682 1049
rect 718 1043 724 1044
rect 622 1038 628 1039
rect 630 1039 636 1040
rect 624 1012 626 1038
rect 630 1035 631 1039
rect 635 1035 636 1039
rect 630 1034 636 1035
rect 678 1039 684 1040
rect 678 1035 679 1039
rect 683 1035 684 1039
rect 718 1039 719 1043
rect 723 1039 724 1043
rect 728 1040 730 1049
rect 774 1043 780 1044
rect 718 1038 724 1039
rect 726 1039 732 1040
rect 678 1034 684 1035
rect 720 1012 722 1038
rect 726 1035 727 1039
rect 731 1035 732 1039
rect 774 1039 775 1043
rect 779 1039 780 1043
rect 784 1040 786 1049
rect 830 1043 836 1044
rect 774 1038 780 1039
rect 782 1039 788 1040
rect 726 1034 732 1035
rect 776 1012 778 1038
rect 782 1035 783 1039
rect 787 1035 788 1039
rect 830 1039 831 1043
rect 835 1039 836 1043
rect 840 1040 842 1049
rect 886 1043 892 1044
rect 830 1038 836 1039
rect 838 1039 844 1040
rect 782 1034 788 1035
rect 832 1012 834 1038
rect 838 1035 839 1039
rect 843 1035 844 1039
rect 886 1039 887 1043
rect 891 1039 892 1043
rect 896 1040 898 1049
rect 950 1043 956 1044
rect 886 1038 892 1039
rect 894 1039 900 1040
rect 838 1034 844 1035
rect 888 1012 890 1038
rect 894 1035 895 1039
rect 899 1035 900 1039
rect 950 1039 951 1043
rect 955 1039 956 1043
rect 960 1040 962 1049
rect 984 1044 986 1086
rect 1016 1068 1018 1138
rect 1046 1132 1052 1133
rect 1046 1128 1047 1132
rect 1051 1128 1052 1132
rect 1046 1127 1052 1128
rect 1102 1132 1108 1133
rect 1102 1128 1103 1132
rect 1107 1128 1108 1132
rect 1102 1127 1108 1128
rect 1150 1132 1156 1133
rect 1150 1128 1151 1132
rect 1155 1128 1156 1132
rect 1150 1127 1156 1128
rect 1190 1132 1196 1133
rect 1190 1128 1191 1132
rect 1195 1128 1196 1132
rect 1190 1127 1196 1128
rect 1023 1126 1027 1127
rect 1023 1121 1027 1122
rect 1047 1126 1051 1127
rect 1047 1121 1051 1122
rect 1087 1126 1091 1127
rect 1087 1121 1091 1122
rect 1103 1126 1107 1127
rect 1103 1121 1107 1122
rect 1151 1126 1155 1127
rect 1151 1121 1155 1122
rect 1191 1126 1195 1127
rect 1191 1121 1195 1122
rect 1022 1120 1028 1121
rect 1022 1116 1023 1120
rect 1027 1116 1028 1120
rect 1022 1115 1028 1116
rect 1086 1120 1092 1121
rect 1086 1116 1087 1120
rect 1091 1116 1092 1120
rect 1086 1115 1092 1116
rect 1150 1120 1156 1121
rect 1150 1116 1151 1120
rect 1155 1116 1156 1120
rect 1150 1115 1156 1116
rect 1190 1120 1196 1121
rect 1190 1116 1191 1120
rect 1195 1116 1196 1120
rect 1190 1115 1196 1116
rect 1216 1108 1218 1178
rect 1240 1157 1242 1189
rect 1279 1185 1283 1186
rect 1511 1190 1515 1191
rect 1511 1185 1515 1186
rect 1551 1190 1555 1191
rect 1551 1185 1555 1186
rect 1559 1190 1563 1191
rect 1559 1185 1563 1186
rect 1591 1190 1595 1191
rect 1591 1185 1595 1186
rect 1599 1190 1603 1191
rect 1599 1185 1603 1186
rect 1631 1190 1635 1191
rect 1631 1185 1635 1186
rect 1639 1190 1643 1191
rect 1639 1185 1643 1186
rect 1671 1190 1675 1191
rect 1671 1185 1675 1186
rect 1679 1190 1683 1191
rect 1679 1185 1683 1186
rect 1711 1190 1715 1191
rect 1711 1185 1715 1186
rect 1719 1190 1723 1191
rect 1719 1185 1723 1186
rect 1751 1190 1755 1191
rect 1751 1185 1755 1186
rect 1759 1190 1763 1191
rect 1759 1185 1763 1186
rect 1238 1156 1244 1157
rect 1238 1152 1239 1156
rect 1243 1152 1244 1156
rect 1280 1153 1282 1185
rect 1560 1176 1562 1185
rect 1600 1176 1602 1185
rect 1614 1183 1620 1184
rect 1614 1179 1615 1183
rect 1619 1179 1620 1183
rect 1614 1178 1620 1179
rect 1626 1179 1632 1180
rect 1558 1175 1564 1176
rect 1558 1171 1559 1175
rect 1563 1171 1564 1175
rect 1558 1170 1564 1171
rect 1598 1175 1604 1176
rect 1598 1171 1599 1175
rect 1603 1171 1604 1175
rect 1598 1170 1604 1171
rect 1238 1151 1244 1152
rect 1278 1152 1284 1153
rect 1278 1148 1279 1152
rect 1283 1148 1284 1152
rect 1616 1148 1618 1178
rect 1626 1175 1627 1179
rect 1631 1175 1632 1179
rect 1640 1176 1642 1185
rect 1680 1176 1682 1185
rect 1694 1183 1700 1184
rect 1694 1179 1695 1183
rect 1699 1179 1700 1183
rect 1694 1178 1700 1179
rect 1626 1174 1632 1175
rect 1638 1175 1644 1176
rect 1628 1156 1630 1174
rect 1638 1171 1639 1175
rect 1643 1171 1644 1175
rect 1638 1170 1644 1171
rect 1678 1175 1684 1176
rect 1678 1171 1679 1175
rect 1683 1171 1684 1175
rect 1678 1170 1684 1171
rect 1626 1155 1632 1156
rect 1626 1151 1627 1155
rect 1631 1151 1632 1155
rect 1626 1150 1632 1151
rect 1696 1148 1698 1178
rect 1720 1176 1722 1185
rect 1734 1183 1740 1184
rect 1734 1179 1735 1183
rect 1739 1179 1740 1183
rect 1734 1178 1740 1179
rect 1718 1175 1724 1176
rect 1718 1171 1719 1175
rect 1723 1171 1724 1175
rect 1718 1170 1724 1171
rect 1736 1148 1738 1178
rect 1760 1176 1762 1185
rect 1768 1184 1770 1230
rect 1790 1209 1796 1210
rect 1790 1205 1791 1209
rect 1795 1205 1796 1209
rect 1790 1204 1796 1205
rect 1792 1191 1794 1204
rect 1791 1190 1795 1191
rect 1791 1185 1795 1186
rect 1799 1190 1803 1191
rect 1799 1185 1803 1186
rect 1766 1183 1772 1184
rect 1766 1179 1767 1183
rect 1771 1179 1772 1183
rect 1766 1178 1772 1179
rect 1800 1176 1802 1185
rect 1808 1184 1810 1230
rect 1838 1209 1844 1210
rect 1838 1205 1839 1209
rect 1843 1205 1844 1209
rect 1838 1204 1844 1205
rect 1902 1209 1908 1210
rect 1902 1205 1903 1209
rect 1907 1205 1908 1209
rect 1902 1204 1908 1205
rect 1966 1209 1972 1210
rect 1966 1205 1967 1209
rect 1971 1205 1972 1209
rect 1966 1204 1972 1205
rect 2032 1204 2034 1230
rect 2038 1209 2044 1210
rect 2038 1205 2039 1209
rect 2043 1205 2044 1209
rect 2038 1204 2044 1205
rect 2118 1209 2124 1210
rect 2118 1205 2119 1209
rect 2123 1205 2124 1209
rect 2118 1204 2124 1205
rect 2144 1204 2146 1278
rect 2166 1272 2172 1273
rect 2166 1268 2167 1272
rect 2171 1268 2172 1272
rect 2166 1267 2172 1268
rect 2270 1272 2276 1273
rect 2270 1268 2271 1272
rect 2275 1268 2276 1272
rect 2270 1267 2276 1268
rect 2168 1263 2170 1267
rect 2272 1263 2274 1267
rect 2167 1262 2171 1263
rect 2167 1257 2171 1258
rect 2207 1262 2211 1263
rect 2207 1257 2211 1258
rect 2271 1262 2275 1263
rect 2271 1257 2275 1258
rect 2206 1256 2212 1257
rect 2206 1252 2207 1256
rect 2211 1252 2212 1256
rect 2206 1251 2212 1252
rect 2284 1236 2286 1318
rect 2296 1292 2298 1342
rect 2304 1335 2306 1348
rect 2360 1335 2362 1348
rect 2374 1347 2380 1348
rect 2374 1343 2375 1347
rect 2379 1343 2380 1347
rect 2374 1342 2380 1343
rect 2303 1334 2307 1335
rect 2303 1329 2307 1330
rect 2359 1334 2363 1335
rect 2359 1329 2363 1330
rect 2360 1320 2362 1329
rect 2384 1324 2386 1374
rect 2406 1372 2407 1376
rect 2411 1372 2412 1376
rect 2406 1371 2412 1372
rect 2408 1335 2410 1371
rect 2407 1334 2411 1335
rect 2407 1329 2411 1330
rect 2382 1323 2388 1324
rect 2358 1319 2364 1320
rect 2358 1315 2359 1319
rect 2363 1315 2364 1319
rect 2382 1319 2383 1323
rect 2387 1319 2388 1323
rect 2382 1318 2388 1319
rect 2358 1314 2364 1315
rect 2408 1297 2410 1329
rect 2406 1296 2412 1297
rect 2406 1292 2407 1296
rect 2411 1292 2412 1296
rect 2294 1291 2300 1292
rect 2294 1287 2295 1291
rect 2299 1287 2300 1291
rect 2294 1286 2300 1287
rect 2382 1291 2388 1292
rect 2406 1291 2412 1292
rect 2382 1287 2383 1291
rect 2387 1287 2388 1291
rect 2382 1286 2388 1287
rect 2358 1272 2364 1273
rect 2358 1268 2359 1272
rect 2363 1268 2364 1272
rect 2358 1267 2364 1268
rect 2360 1263 2362 1267
rect 2295 1262 2299 1263
rect 2295 1257 2299 1258
rect 2359 1262 2363 1263
rect 2359 1257 2363 1258
rect 2294 1256 2300 1257
rect 2294 1252 2295 1256
rect 2299 1252 2300 1256
rect 2294 1251 2300 1252
rect 2358 1256 2364 1257
rect 2358 1252 2359 1256
rect 2363 1252 2364 1256
rect 2358 1251 2364 1252
rect 2282 1235 2288 1236
rect 2282 1231 2283 1235
rect 2287 1231 2288 1235
rect 2282 1230 2288 1231
rect 2318 1235 2324 1236
rect 2318 1231 2319 1235
rect 2323 1231 2324 1235
rect 2318 1230 2324 1231
rect 2206 1209 2212 1210
rect 2206 1205 2207 1209
rect 2211 1205 2212 1209
rect 2206 1204 2212 1205
rect 2294 1209 2300 1210
rect 2294 1205 2295 1209
rect 2299 1205 2300 1209
rect 2294 1204 2300 1205
rect 1840 1191 1842 1204
rect 1904 1191 1906 1204
rect 1968 1191 1970 1204
rect 2030 1203 2036 1204
rect 2030 1199 2031 1203
rect 2035 1199 2036 1203
rect 2030 1198 2036 1199
rect 2040 1191 2042 1204
rect 2120 1191 2122 1204
rect 2142 1203 2148 1204
rect 2142 1199 2143 1203
rect 2147 1199 2148 1203
rect 2142 1198 2148 1199
rect 2208 1191 2210 1204
rect 2218 1203 2224 1204
rect 2218 1199 2219 1203
rect 2223 1199 2224 1203
rect 2218 1198 2224 1199
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1855 1190 1859 1191
rect 1855 1185 1859 1186
rect 1903 1190 1907 1191
rect 1903 1185 1907 1186
rect 1927 1190 1931 1191
rect 1927 1185 1931 1186
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 2023 1190 2027 1191
rect 2023 1185 2027 1186
rect 2039 1190 2043 1191
rect 2039 1185 2043 1186
rect 2119 1190 2123 1191
rect 2119 1185 2123 1186
rect 2135 1190 2139 1191
rect 2135 1185 2139 1186
rect 2207 1190 2211 1191
rect 2207 1185 2211 1186
rect 1806 1183 1812 1184
rect 1806 1179 1807 1183
rect 1811 1179 1812 1183
rect 1806 1178 1812 1179
rect 1814 1179 1820 1180
rect 1758 1175 1764 1176
rect 1758 1171 1759 1175
rect 1763 1171 1764 1175
rect 1758 1170 1764 1171
rect 1798 1175 1804 1176
rect 1798 1171 1799 1175
rect 1803 1171 1804 1175
rect 1814 1175 1815 1179
rect 1819 1175 1820 1179
rect 1856 1176 1858 1185
rect 1866 1179 1872 1180
rect 1814 1174 1820 1175
rect 1854 1175 1860 1176
rect 1798 1170 1804 1171
rect 1816 1148 1818 1174
rect 1854 1171 1855 1175
rect 1859 1171 1860 1175
rect 1866 1175 1867 1179
rect 1871 1175 1872 1179
rect 1928 1176 1930 1185
rect 1938 1179 1944 1180
rect 1866 1174 1872 1175
rect 1926 1175 1932 1176
rect 1854 1170 1860 1171
rect 1868 1148 1870 1174
rect 1926 1171 1927 1175
rect 1931 1171 1932 1175
rect 1938 1175 1939 1179
rect 1943 1175 1944 1179
rect 2024 1176 2026 1185
rect 2126 1179 2132 1180
rect 1938 1174 1944 1175
rect 2022 1175 2028 1176
rect 1926 1170 1932 1171
rect 1940 1148 1942 1174
rect 2022 1171 2023 1175
rect 2027 1171 2028 1175
rect 2126 1175 2127 1179
rect 2131 1175 2132 1179
rect 2136 1176 2138 1185
rect 2126 1174 2132 1175
rect 2134 1175 2140 1176
rect 2022 1170 2028 1171
rect 2128 1148 2130 1174
rect 2134 1171 2135 1175
rect 2139 1171 2140 1175
rect 2134 1170 2140 1171
rect 1278 1147 1284 1148
rect 1614 1147 1620 1148
rect 1614 1143 1615 1147
rect 1619 1143 1620 1147
rect 1614 1142 1620 1143
rect 1694 1147 1700 1148
rect 1694 1143 1695 1147
rect 1699 1143 1700 1147
rect 1694 1142 1700 1143
rect 1734 1147 1740 1148
rect 1734 1143 1735 1147
rect 1739 1143 1740 1147
rect 1734 1142 1740 1143
rect 1814 1147 1820 1148
rect 1814 1143 1815 1147
rect 1819 1143 1820 1147
rect 1814 1142 1820 1143
rect 1866 1147 1872 1148
rect 1866 1143 1867 1147
rect 1871 1143 1872 1147
rect 1866 1142 1872 1143
rect 1938 1147 1944 1148
rect 1938 1143 1939 1147
rect 1943 1143 1944 1147
rect 1938 1142 1944 1143
rect 1974 1147 1980 1148
rect 1974 1143 1975 1147
rect 1979 1143 1980 1147
rect 1974 1142 1980 1143
rect 2126 1147 2132 1148
rect 2126 1143 2127 1147
rect 2131 1143 2132 1147
rect 2126 1142 2132 1143
rect 1238 1139 1244 1140
rect 1238 1135 1239 1139
rect 1243 1135 1244 1139
rect 1750 1139 1756 1140
rect 1238 1134 1244 1135
rect 1278 1135 1284 1136
rect 1240 1127 1242 1134
rect 1278 1131 1279 1135
rect 1283 1131 1284 1135
rect 1750 1135 1751 1139
rect 1755 1135 1756 1139
rect 1750 1134 1756 1135
rect 1278 1130 1284 1131
rect 1239 1126 1243 1127
rect 1239 1121 1243 1122
rect 1240 1114 1242 1121
rect 1280 1115 1282 1130
rect 1558 1128 1564 1129
rect 1558 1124 1559 1128
rect 1563 1124 1564 1128
rect 1558 1123 1564 1124
rect 1598 1128 1604 1129
rect 1598 1124 1599 1128
rect 1603 1124 1604 1128
rect 1598 1123 1604 1124
rect 1638 1128 1644 1129
rect 1638 1124 1639 1128
rect 1643 1124 1644 1128
rect 1638 1123 1644 1124
rect 1678 1128 1684 1129
rect 1678 1124 1679 1128
rect 1683 1124 1684 1128
rect 1678 1123 1684 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1560 1115 1562 1123
rect 1600 1115 1602 1123
rect 1640 1115 1642 1123
rect 1680 1115 1682 1123
rect 1720 1115 1722 1123
rect 1279 1114 1283 1115
rect 1238 1113 1244 1114
rect 1238 1109 1239 1113
rect 1243 1109 1244 1113
rect 1279 1109 1283 1110
rect 1535 1114 1539 1115
rect 1535 1109 1539 1110
rect 1559 1114 1563 1115
rect 1559 1109 1563 1110
rect 1599 1114 1603 1115
rect 1599 1109 1603 1110
rect 1639 1114 1643 1115
rect 1639 1109 1643 1110
rect 1663 1114 1667 1115
rect 1663 1109 1667 1110
rect 1679 1114 1683 1115
rect 1679 1109 1683 1110
rect 1719 1114 1723 1115
rect 1719 1109 1723 1110
rect 1727 1114 1731 1115
rect 1727 1109 1731 1110
rect 1238 1108 1244 1109
rect 1214 1107 1220 1108
rect 1214 1103 1215 1107
rect 1219 1103 1220 1107
rect 1214 1102 1220 1103
rect 1280 1102 1282 1109
rect 1534 1108 1540 1109
rect 1534 1104 1535 1108
rect 1539 1104 1540 1108
rect 1534 1103 1540 1104
rect 1598 1108 1604 1109
rect 1598 1104 1599 1108
rect 1603 1104 1604 1108
rect 1598 1103 1604 1104
rect 1662 1108 1668 1109
rect 1662 1104 1663 1108
rect 1667 1104 1668 1108
rect 1662 1103 1668 1104
rect 1726 1108 1732 1109
rect 1726 1104 1727 1108
rect 1731 1104 1732 1108
rect 1726 1103 1732 1104
rect 1278 1101 1284 1102
rect 1198 1099 1204 1100
rect 1198 1095 1199 1099
rect 1203 1095 1204 1099
rect 1278 1097 1279 1101
rect 1283 1097 1284 1101
rect 1198 1094 1204 1095
rect 1238 1096 1244 1097
rect 1278 1096 1284 1097
rect 1022 1073 1028 1074
rect 1022 1069 1023 1073
rect 1027 1069 1028 1073
rect 1022 1068 1028 1069
rect 1086 1073 1092 1074
rect 1086 1069 1087 1073
rect 1091 1069 1092 1073
rect 1086 1068 1092 1069
rect 1150 1073 1156 1074
rect 1150 1069 1151 1073
rect 1155 1069 1156 1073
rect 1150 1068 1156 1069
rect 1190 1073 1196 1074
rect 1190 1069 1191 1073
rect 1195 1069 1196 1073
rect 1190 1068 1196 1069
rect 1200 1068 1202 1094
rect 1238 1092 1239 1096
rect 1243 1092 1244 1096
rect 1238 1091 1244 1092
rect 1014 1067 1020 1068
rect 1014 1063 1015 1067
rect 1019 1063 1020 1067
rect 1014 1062 1020 1063
rect 1024 1055 1026 1068
rect 1088 1055 1090 1068
rect 1152 1055 1154 1068
rect 1192 1055 1194 1068
rect 1198 1067 1204 1068
rect 1198 1063 1199 1067
rect 1203 1063 1204 1067
rect 1198 1062 1204 1063
rect 1214 1067 1220 1068
rect 1214 1063 1215 1067
rect 1219 1063 1220 1067
rect 1214 1062 1220 1063
rect 1023 1054 1027 1055
rect 1023 1049 1027 1050
rect 1087 1054 1091 1055
rect 1087 1049 1091 1050
rect 1151 1054 1155 1055
rect 1151 1049 1155 1050
rect 1191 1054 1195 1055
rect 1191 1049 1195 1050
rect 982 1043 988 1044
rect 950 1038 956 1039
rect 958 1039 964 1040
rect 894 1034 900 1035
rect 952 1012 954 1038
rect 958 1035 959 1039
rect 963 1035 964 1039
rect 982 1039 983 1043
rect 987 1039 988 1043
rect 1024 1040 1026 1049
rect 1078 1043 1084 1044
rect 982 1038 988 1039
rect 1022 1039 1028 1040
rect 958 1034 964 1035
rect 1022 1035 1023 1039
rect 1027 1035 1028 1039
rect 1078 1039 1079 1043
rect 1083 1039 1084 1043
rect 1088 1040 1090 1049
rect 1110 1043 1116 1044
rect 1078 1038 1084 1039
rect 1086 1039 1092 1040
rect 1022 1034 1028 1035
rect 1080 1012 1082 1038
rect 1086 1035 1087 1039
rect 1091 1035 1092 1039
rect 1110 1039 1111 1043
rect 1115 1039 1116 1043
rect 1152 1040 1154 1049
rect 1166 1043 1172 1044
rect 1110 1038 1116 1039
rect 1150 1039 1156 1040
rect 1086 1034 1092 1035
rect 478 1011 484 1012
rect 478 1007 479 1011
rect 483 1007 484 1011
rect 478 1006 484 1007
rect 526 1011 532 1012
rect 526 1007 527 1011
rect 531 1007 532 1011
rect 526 1006 532 1007
rect 610 1011 616 1012
rect 610 1007 611 1011
rect 615 1007 616 1011
rect 610 1006 616 1007
rect 622 1011 628 1012
rect 622 1007 623 1011
rect 627 1007 628 1011
rect 622 1006 628 1007
rect 718 1011 724 1012
rect 718 1007 719 1011
rect 723 1007 724 1011
rect 718 1006 724 1007
rect 774 1011 780 1012
rect 774 1007 775 1011
rect 779 1007 780 1011
rect 774 1006 780 1007
rect 830 1011 836 1012
rect 830 1007 831 1011
rect 835 1007 836 1011
rect 830 1006 836 1007
rect 886 1011 892 1012
rect 886 1007 887 1011
rect 891 1007 892 1011
rect 886 1006 892 1007
rect 950 1011 956 1012
rect 950 1007 951 1011
rect 955 1007 956 1011
rect 950 1006 956 1007
rect 1078 1011 1084 1012
rect 1078 1007 1079 1011
rect 1083 1007 1084 1011
rect 1078 1006 1084 1007
rect 574 1003 580 1004
rect 574 999 575 1003
rect 579 999 580 1003
rect 574 998 580 999
rect 438 992 444 993
rect 438 988 439 992
rect 443 988 444 992
rect 438 987 444 988
rect 486 992 492 993
rect 486 988 487 992
rect 491 988 492 992
rect 486 987 492 988
rect 534 992 540 993
rect 534 988 535 992
rect 539 988 540 992
rect 534 987 540 988
rect 440 975 442 987
rect 488 975 490 987
rect 536 975 538 987
rect 439 974 443 975
rect 439 969 443 970
rect 471 974 475 975
rect 471 969 475 970
rect 487 974 491 975
rect 487 969 491 970
rect 535 974 539 975
rect 535 969 539 970
rect 551 974 555 975
rect 551 969 555 970
rect 470 968 476 969
rect 470 964 471 968
rect 475 964 476 968
rect 470 963 476 964
rect 550 968 556 969
rect 550 964 551 968
rect 555 964 556 968
rect 550 963 556 964
rect 406 955 412 956
rect 406 951 407 955
rect 411 951 412 955
rect 406 950 412 951
rect 110 944 116 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 112 899 114 939
rect 294 921 300 922
rect 294 917 295 921
rect 299 917 300 921
rect 294 916 300 917
rect 342 921 348 922
rect 342 917 343 921
rect 347 917 348 921
rect 342 916 348 917
rect 398 921 404 922
rect 398 917 399 921
rect 403 917 404 921
rect 398 916 404 917
rect 470 921 476 922
rect 470 917 471 921
rect 475 917 476 921
rect 470 916 476 917
rect 550 921 556 922
rect 550 917 551 921
rect 555 917 556 921
rect 550 916 556 917
rect 576 916 578 998
rect 582 992 588 993
rect 582 988 583 992
rect 587 988 588 992
rect 582 987 588 988
rect 630 992 636 993
rect 630 988 631 992
rect 635 988 636 992
rect 630 987 636 988
rect 678 992 684 993
rect 678 988 679 992
rect 683 988 684 992
rect 678 987 684 988
rect 726 992 732 993
rect 726 988 727 992
rect 731 988 732 992
rect 726 987 732 988
rect 782 992 788 993
rect 782 988 783 992
rect 787 988 788 992
rect 782 987 788 988
rect 838 992 844 993
rect 838 988 839 992
rect 843 988 844 992
rect 838 987 844 988
rect 894 992 900 993
rect 894 988 895 992
rect 899 988 900 992
rect 894 987 900 988
rect 958 992 964 993
rect 958 988 959 992
rect 963 988 964 992
rect 958 987 964 988
rect 1022 992 1028 993
rect 1022 988 1023 992
rect 1027 988 1028 992
rect 1022 987 1028 988
rect 1086 992 1092 993
rect 1086 988 1087 992
rect 1091 988 1092 992
rect 1086 987 1092 988
rect 584 975 586 987
rect 632 975 634 987
rect 680 975 682 987
rect 728 975 730 987
rect 784 975 786 987
rect 840 975 842 987
rect 896 975 898 987
rect 960 975 962 987
rect 1024 975 1026 987
rect 1088 975 1090 987
rect 583 974 587 975
rect 583 969 587 970
rect 631 974 635 975
rect 631 969 635 970
rect 639 974 643 975
rect 639 969 643 970
rect 679 974 683 975
rect 679 969 683 970
rect 727 974 731 975
rect 727 969 731 970
rect 783 974 787 975
rect 783 969 787 970
rect 807 974 811 975
rect 807 969 811 970
rect 839 974 843 975
rect 839 969 843 970
rect 887 974 891 975
rect 887 969 891 970
rect 895 974 899 975
rect 895 969 899 970
rect 959 974 963 975
rect 959 969 963 970
rect 1023 974 1027 975
rect 1023 969 1027 970
rect 1087 974 1091 975
rect 1087 969 1091 970
rect 638 968 644 969
rect 638 964 639 968
rect 643 964 644 968
rect 638 963 644 964
rect 726 968 732 969
rect 726 964 727 968
rect 731 964 732 968
rect 726 963 732 964
rect 806 968 812 969
rect 806 964 807 968
rect 811 964 812 968
rect 806 963 812 964
rect 886 968 892 969
rect 886 964 887 968
rect 891 964 892 968
rect 886 963 892 964
rect 958 968 964 969
rect 958 964 959 968
rect 963 964 964 968
rect 958 963 964 964
rect 1022 968 1028 969
rect 1022 964 1023 968
rect 1027 964 1028 968
rect 1022 963 1028 964
rect 1086 968 1092 969
rect 1086 964 1087 968
rect 1091 964 1092 968
rect 1086 963 1092 964
rect 1112 948 1114 1038
rect 1150 1035 1151 1039
rect 1155 1035 1156 1039
rect 1166 1039 1167 1043
rect 1171 1039 1172 1043
rect 1192 1040 1194 1049
rect 1202 1043 1208 1044
rect 1166 1038 1172 1039
rect 1190 1039 1196 1040
rect 1150 1034 1156 1035
rect 1168 1020 1170 1038
rect 1190 1035 1191 1039
rect 1195 1035 1196 1039
rect 1202 1039 1203 1043
rect 1207 1039 1208 1043
rect 1202 1038 1208 1039
rect 1190 1034 1196 1035
rect 1166 1019 1172 1020
rect 1166 1015 1167 1019
rect 1171 1015 1172 1019
rect 1166 1014 1172 1015
rect 1204 1012 1206 1038
rect 1216 1012 1218 1062
rect 1240 1055 1242 1091
rect 1278 1084 1284 1085
rect 1278 1080 1279 1084
rect 1283 1080 1284 1084
rect 1278 1079 1284 1080
rect 1239 1054 1243 1055
rect 1239 1049 1243 1050
rect 1240 1017 1242 1049
rect 1280 1035 1282 1079
rect 1534 1061 1540 1062
rect 1534 1057 1535 1061
rect 1539 1057 1540 1061
rect 1534 1056 1540 1057
rect 1598 1061 1604 1062
rect 1598 1057 1599 1061
rect 1603 1057 1604 1061
rect 1598 1056 1604 1057
rect 1662 1061 1668 1062
rect 1662 1057 1663 1061
rect 1667 1057 1668 1061
rect 1662 1056 1668 1057
rect 1726 1061 1732 1062
rect 1726 1057 1727 1061
rect 1731 1057 1732 1061
rect 1726 1056 1732 1057
rect 1752 1056 1754 1134
rect 1758 1128 1764 1129
rect 1758 1124 1759 1128
rect 1763 1124 1764 1128
rect 1758 1123 1764 1124
rect 1798 1128 1804 1129
rect 1798 1124 1799 1128
rect 1803 1124 1804 1128
rect 1798 1123 1804 1124
rect 1854 1128 1860 1129
rect 1854 1124 1855 1128
rect 1859 1124 1860 1128
rect 1854 1123 1860 1124
rect 1926 1128 1932 1129
rect 1926 1124 1927 1128
rect 1931 1124 1932 1128
rect 1926 1123 1932 1124
rect 1760 1115 1762 1123
rect 1800 1115 1802 1123
rect 1856 1115 1858 1123
rect 1928 1115 1930 1123
rect 1759 1114 1763 1115
rect 1759 1109 1763 1110
rect 1791 1114 1795 1115
rect 1791 1109 1795 1110
rect 1799 1114 1803 1115
rect 1799 1109 1803 1110
rect 1855 1114 1859 1115
rect 1855 1109 1859 1110
rect 1911 1114 1915 1115
rect 1911 1109 1915 1110
rect 1927 1114 1931 1115
rect 1927 1109 1931 1110
rect 1967 1114 1971 1115
rect 1967 1109 1971 1110
rect 1790 1108 1796 1109
rect 1790 1104 1791 1108
rect 1795 1104 1796 1108
rect 1790 1103 1796 1104
rect 1854 1108 1860 1109
rect 1854 1104 1855 1108
rect 1859 1104 1860 1108
rect 1854 1103 1860 1104
rect 1910 1108 1916 1109
rect 1910 1104 1911 1108
rect 1915 1104 1916 1108
rect 1910 1103 1916 1104
rect 1966 1108 1972 1109
rect 1966 1104 1967 1108
rect 1971 1104 1972 1108
rect 1966 1103 1972 1104
rect 1758 1079 1764 1080
rect 1758 1075 1759 1079
rect 1763 1075 1764 1079
rect 1758 1074 1764 1075
rect 1536 1035 1538 1056
rect 1600 1035 1602 1056
rect 1664 1035 1666 1056
rect 1728 1035 1730 1056
rect 1750 1055 1756 1056
rect 1750 1051 1751 1055
rect 1755 1051 1756 1055
rect 1750 1050 1756 1051
rect 1279 1034 1283 1035
rect 1279 1029 1283 1030
rect 1503 1034 1507 1035
rect 1503 1029 1507 1030
rect 1535 1034 1539 1035
rect 1535 1029 1539 1030
rect 1599 1034 1603 1035
rect 1599 1029 1603 1030
rect 1623 1034 1627 1035
rect 1623 1029 1627 1030
rect 1663 1034 1667 1035
rect 1663 1029 1667 1030
rect 1727 1034 1731 1035
rect 1727 1029 1731 1030
rect 1735 1034 1739 1035
rect 1735 1029 1739 1030
rect 1238 1016 1244 1017
rect 1238 1012 1239 1016
rect 1243 1012 1244 1016
rect 1202 1011 1208 1012
rect 1202 1007 1203 1011
rect 1207 1007 1208 1011
rect 1202 1006 1208 1007
rect 1214 1011 1220 1012
rect 1238 1011 1244 1012
rect 1214 1007 1215 1011
rect 1219 1007 1220 1011
rect 1214 1006 1220 1007
rect 1238 999 1244 1000
rect 1238 995 1239 999
rect 1243 995 1244 999
rect 1280 997 1282 1029
rect 1504 1020 1506 1029
rect 1614 1023 1620 1024
rect 1502 1019 1508 1020
rect 1502 1015 1503 1019
rect 1507 1015 1508 1019
rect 1614 1019 1615 1023
rect 1619 1019 1620 1023
rect 1624 1020 1626 1029
rect 1726 1023 1732 1024
rect 1614 1018 1620 1019
rect 1622 1019 1628 1020
rect 1502 1014 1508 1015
rect 1238 994 1244 995
rect 1278 996 1284 997
rect 1150 992 1156 993
rect 1150 988 1151 992
rect 1155 988 1156 992
rect 1150 987 1156 988
rect 1190 992 1196 993
rect 1190 988 1191 992
rect 1195 988 1196 992
rect 1190 987 1196 988
rect 1152 975 1154 987
rect 1192 975 1194 987
rect 1240 975 1242 994
rect 1278 992 1279 996
rect 1283 992 1284 996
rect 1616 992 1618 1018
rect 1622 1015 1623 1019
rect 1627 1015 1628 1019
rect 1726 1019 1727 1023
rect 1731 1019 1732 1023
rect 1736 1020 1738 1029
rect 1760 1024 1762 1074
rect 1790 1061 1796 1062
rect 1790 1057 1791 1061
rect 1795 1057 1796 1061
rect 1790 1056 1796 1057
rect 1854 1061 1860 1062
rect 1854 1057 1855 1061
rect 1859 1057 1860 1061
rect 1854 1056 1860 1057
rect 1910 1061 1916 1062
rect 1910 1057 1911 1061
rect 1915 1057 1916 1061
rect 1910 1056 1916 1057
rect 1966 1061 1972 1062
rect 1966 1057 1967 1061
rect 1971 1057 1972 1061
rect 1966 1056 1972 1057
rect 1976 1056 1978 1142
rect 2022 1128 2028 1129
rect 2022 1124 2023 1128
rect 2027 1124 2028 1128
rect 2022 1123 2028 1124
rect 2134 1128 2140 1129
rect 2134 1124 2135 1128
rect 2139 1124 2140 1128
rect 2134 1123 2140 1124
rect 2024 1115 2026 1123
rect 2136 1115 2138 1123
rect 2023 1114 2027 1115
rect 2023 1109 2027 1110
rect 2079 1114 2083 1115
rect 2079 1109 2083 1110
rect 2135 1114 2139 1115
rect 2135 1109 2139 1110
rect 2191 1114 2195 1115
rect 2191 1109 2195 1110
rect 2022 1108 2028 1109
rect 2022 1104 2023 1108
rect 2027 1104 2028 1108
rect 2022 1103 2028 1104
rect 2078 1108 2084 1109
rect 2078 1104 2079 1108
rect 2083 1104 2084 1108
rect 2078 1103 2084 1104
rect 2134 1108 2140 1109
rect 2134 1104 2135 1108
rect 2139 1104 2140 1108
rect 2134 1103 2140 1104
rect 2190 1108 2196 1109
rect 2190 1104 2191 1108
rect 2195 1104 2196 1108
rect 2190 1103 2196 1104
rect 2220 1088 2222 1198
rect 2296 1191 2298 1204
rect 2255 1190 2259 1191
rect 2255 1185 2259 1186
rect 2295 1190 2299 1191
rect 2295 1185 2299 1186
rect 2246 1179 2252 1180
rect 2246 1175 2247 1179
rect 2251 1175 2252 1179
rect 2256 1176 2258 1185
rect 2320 1184 2322 1230
rect 2358 1209 2364 1210
rect 2358 1205 2359 1209
rect 2363 1205 2364 1209
rect 2358 1204 2364 1205
rect 2384 1204 2386 1286
rect 2406 1279 2412 1280
rect 2406 1275 2407 1279
rect 2411 1275 2412 1279
rect 2406 1274 2412 1275
rect 2408 1263 2410 1274
rect 2407 1262 2411 1263
rect 2407 1257 2411 1258
rect 2408 1250 2410 1257
rect 2406 1249 2412 1250
rect 2406 1245 2407 1249
rect 2411 1245 2412 1249
rect 2406 1244 2412 1245
rect 2406 1232 2412 1233
rect 2406 1228 2407 1232
rect 2411 1228 2412 1232
rect 2406 1227 2412 1228
rect 2360 1191 2362 1204
rect 2382 1203 2388 1204
rect 2382 1199 2383 1203
rect 2387 1199 2388 1203
rect 2382 1198 2388 1199
rect 2408 1191 2410 1227
rect 2359 1190 2363 1191
rect 2359 1185 2363 1186
rect 2407 1190 2411 1191
rect 2407 1185 2411 1186
rect 2318 1183 2324 1184
rect 2266 1179 2272 1180
rect 2246 1174 2252 1175
rect 2254 1175 2260 1176
rect 2248 1148 2250 1174
rect 2254 1171 2255 1175
rect 2259 1171 2260 1175
rect 2266 1175 2267 1179
rect 2271 1175 2272 1179
rect 2318 1179 2319 1183
rect 2323 1179 2324 1183
rect 2318 1178 2324 1179
rect 2360 1176 2362 1185
rect 2266 1174 2272 1175
rect 2358 1175 2364 1176
rect 2254 1170 2260 1171
rect 2268 1156 2270 1174
rect 2358 1171 2359 1175
rect 2363 1171 2364 1175
rect 2358 1170 2364 1171
rect 2266 1155 2272 1156
rect 2266 1151 2267 1155
rect 2271 1151 2272 1155
rect 2408 1153 2410 1185
rect 2266 1150 2272 1151
rect 2406 1152 2412 1153
rect 2406 1148 2407 1152
rect 2411 1148 2412 1152
rect 2246 1147 2252 1148
rect 2246 1143 2247 1147
rect 2251 1143 2252 1147
rect 2246 1142 2252 1143
rect 2382 1147 2388 1148
rect 2406 1147 2412 1148
rect 2382 1143 2383 1147
rect 2387 1143 2388 1147
rect 2382 1142 2388 1143
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 2256 1115 2258 1123
rect 2360 1115 2362 1123
rect 2255 1114 2259 1115
rect 2255 1109 2259 1110
rect 2319 1114 2323 1115
rect 2319 1109 2323 1110
rect 2359 1114 2363 1115
rect 2359 1109 2363 1110
rect 2254 1108 2260 1109
rect 2254 1104 2255 1108
rect 2259 1104 2260 1108
rect 2254 1103 2260 1104
rect 2318 1108 2324 1109
rect 2318 1104 2319 1108
rect 2323 1104 2324 1108
rect 2318 1103 2324 1104
rect 2358 1108 2364 1109
rect 2358 1104 2359 1108
rect 2363 1104 2364 1108
rect 2358 1103 2364 1104
rect 2038 1087 2044 1088
rect 2038 1083 2039 1087
rect 2043 1083 2044 1087
rect 2038 1082 2044 1083
rect 2218 1087 2224 1088
rect 2218 1083 2219 1087
rect 2223 1083 2224 1087
rect 2218 1082 2224 1083
rect 2226 1087 2232 1088
rect 2226 1083 2227 1087
rect 2231 1083 2232 1087
rect 2226 1082 2232 1083
rect 2366 1087 2372 1088
rect 2366 1083 2367 1087
rect 2371 1083 2372 1087
rect 2366 1082 2372 1083
rect 1990 1079 1996 1080
rect 1990 1075 1991 1079
rect 1995 1075 1996 1079
rect 1990 1074 1996 1075
rect 1992 1056 1994 1074
rect 2022 1061 2028 1062
rect 2022 1057 2023 1061
rect 2027 1057 2028 1061
rect 2022 1056 2028 1057
rect 1792 1035 1794 1056
rect 1856 1035 1858 1056
rect 1912 1035 1914 1056
rect 1968 1035 1970 1056
rect 1974 1055 1980 1056
rect 1974 1051 1975 1055
rect 1979 1051 1980 1055
rect 1974 1050 1980 1051
rect 1990 1055 1996 1056
rect 1990 1051 1991 1055
rect 1995 1051 1996 1055
rect 1990 1050 1996 1051
rect 2024 1035 2026 1056
rect 1791 1034 1795 1035
rect 1791 1029 1795 1030
rect 1831 1034 1835 1035
rect 1831 1029 1835 1030
rect 1855 1034 1859 1035
rect 1855 1029 1859 1030
rect 1911 1034 1915 1035
rect 1911 1029 1915 1030
rect 1919 1034 1923 1035
rect 1919 1029 1923 1030
rect 1967 1034 1971 1035
rect 1967 1029 1971 1030
rect 1999 1034 2003 1035
rect 1999 1029 2003 1030
rect 2023 1034 2027 1035
rect 2023 1029 2027 1030
rect 1758 1023 1764 1024
rect 1726 1018 1732 1019
rect 1734 1019 1740 1020
rect 1622 1014 1628 1015
rect 1728 992 1730 1018
rect 1734 1015 1735 1019
rect 1739 1015 1740 1019
rect 1758 1019 1759 1023
rect 1763 1019 1764 1023
rect 1832 1020 1834 1029
rect 1920 1020 1922 1029
rect 1934 1027 1940 1028
rect 1934 1023 1935 1027
rect 1939 1023 1940 1027
rect 1934 1022 1940 1023
rect 1758 1018 1764 1019
rect 1830 1019 1836 1020
rect 1734 1014 1740 1015
rect 1830 1015 1831 1019
rect 1835 1015 1836 1019
rect 1830 1014 1836 1015
rect 1918 1019 1924 1020
rect 1918 1015 1919 1019
rect 1923 1015 1924 1019
rect 1918 1014 1924 1015
rect 1936 992 1938 1022
rect 2000 1020 2002 1029
rect 2040 1028 2042 1082
rect 2146 1079 2152 1080
rect 2146 1075 2147 1079
rect 2151 1075 2152 1079
rect 2146 1074 2152 1075
rect 2078 1061 2084 1062
rect 2078 1057 2079 1061
rect 2083 1057 2084 1061
rect 2078 1056 2084 1057
rect 2134 1061 2140 1062
rect 2134 1057 2135 1061
rect 2139 1057 2140 1061
rect 2134 1056 2140 1057
rect 2148 1056 2150 1074
rect 2190 1061 2196 1062
rect 2190 1057 2191 1061
rect 2195 1057 2196 1061
rect 2190 1056 2196 1057
rect 2228 1056 2230 1082
rect 2254 1061 2260 1062
rect 2254 1057 2255 1061
rect 2259 1057 2260 1061
rect 2254 1056 2260 1057
rect 2318 1061 2324 1062
rect 2318 1057 2319 1061
rect 2323 1057 2324 1061
rect 2318 1056 2324 1057
rect 2358 1061 2364 1062
rect 2358 1057 2359 1061
rect 2363 1057 2364 1061
rect 2358 1056 2364 1057
rect 2368 1056 2370 1082
rect 2384 1056 2386 1142
rect 2406 1135 2412 1136
rect 2406 1131 2407 1135
rect 2411 1131 2412 1135
rect 2406 1130 2412 1131
rect 2408 1115 2410 1130
rect 2407 1114 2411 1115
rect 2407 1109 2411 1110
rect 2408 1102 2410 1109
rect 2406 1101 2412 1102
rect 2406 1097 2407 1101
rect 2411 1097 2412 1101
rect 2406 1096 2412 1097
rect 2406 1084 2412 1085
rect 2406 1080 2407 1084
rect 2411 1080 2412 1084
rect 2406 1079 2412 1080
rect 2080 1035 2082 1056
rect 2136 1035 2138 1056
rect 2146 1055 2152 1056
rect 2146 1051 2147 1055
rect 2151 1051 2152 1055
rect 2146 1050 2152 1051
rect 2192 1035 2194 1056
rect 2226 1055 2232 1056
rect 2226 1051 2227 1055
rect 2231 1051 2232 1055
rect 2226 1050 2232 1051
rect 2256 1035 2258 1056
rect 2320 1035 2322 1056
rect 2360 1035 2362 1056
rect 2366 1055 2372 1056
rect 2366 1051 2367 1055
rect 2371 1051 2372 1055
rect 2366 1050 2372 1051
rect 2382 1055 2388 1056
rect 2382 1051 2383 1055
rect 2387 1051 2388 1055
rect 2382 1050 2388 1051
rect 2408 1035 2410 1079
rect 2071 1034 2075 1035
rect 2071 1029 2075 1030
rect 2079 1034 2083 1035
rect 2079 1029 2083 1030
rect 2135 1034 2139 1035
rect 2135 1029 2139 1030
rect 2143 1034 2147 1035
rect 2143 1029 2147 1030
rect 2191 1034 2195 1035
rect 2191 1029 2195 1030
rect 2207 1034 2211 1035
rect 2207 1029 2211 1030
rect 2255 1034 2259 1035
rect 2255 1029 2259 1030
rect 2279 1034 2283 1035
rect 2279 1029 2283 1030
rect 2319 1034 2323 1035
rect 2319 1029 2323 1030
rect 2359 1034 2363 1035
rect 2359 1029 2363 1030
rect 2407 1034 2411 1035
rect 2407 1029 2411 1030
rect 2038 1027 2044 1028
rect 2038 1023 2039 1027
rect 2043 1023 2044 1027
rect 2038 1022 2044 1023
rect 2072 1020 2074 1029
rect 2082 1023 2088 1024
rect 1998 1019 2004 1020
rect 1998 1015 1999 1019
rect 2003 1015 2004 1019
rect 1998 1014 2004 1015
rect 2070 1019 2076 1020
rect 2070 1015 2071 1019
rect 2075 1015 2076 1019
rect 2082 1019 2083 1023
rect 2087 1019 2088 1023
rect 2144 1020 2146 1029
rect 2198 1023 2204 1024
rect 2082 1018 2088 1019
rect 2142 1019 2148 1020
rect 2070 1014 2076 1015
rect 2084 1000 2086 1018
rect 2142 1015 2143 1019
rect 2147 1015 2148 1019
rect 2198 1019 2199 1023
rect 2203 1019 2204 1023
rect 2208 1020 2210 1029
rect 2270 1023 2276 1024
rect 2198 1018 2204 1019
rect 2206 1019 2212 1020
rect 2142 1014 2148 1015
rect 2082 999 2088 1000
rect 2082 995 2083 999
rect 2087 995 2088 999
rect 2082 994 2088 995
rect 2200 992 2202 1018
rect 2206 1015 2207 1019
rect 2211 1015 2212 1019
rect 2270 1019 2271 1023
rect 2275 1019 2276 1023
rect 2280 1020 2282 1029
rect 2290 1023 2296 1024
rect 2270 1018 2276 1019
rect 2278 1019 2284 1020
rect 2206 1014 2212 1015
rect 2272 992 2274 1018
rect 2278 1015 2279 1019
rect 2283 1015 2284 1019
rect 2290 1019 2291 1023
rect 2295 1019 2296 1023
rect 2290 1018 2296 1019
rect 2278 1014 2284 1015
rect 2292 1000 2294 1018
rect 2290 999 2296 1000
rect 2290 995 2291 999
rect 2295 995 2296 999
rect 2408 997 2410 1029
rect 2290 994 2296 995
rect 2406 996 2412 997
rect 2406 992 2407 996
rect 2411 992 2412 996
rect 1278 991 1284 992
rect 1614 991 1620 992
rect 1614 987 1615 991
rect 1619 987 1620 991
rect 1614 986 1620 987
rect 1726 991 1732 992
rect 1726 987 1727 991
rect 1731 987 1732 991
rect 1726 986 1732 987
rect 1934 991 1940 992
rect 1934 987 1935 991
rect 1939 987 1940 991
rect 1934 986 1940 987
rect 2130 991 2136 992
rect 2130 987 2131 991
rect 2135 987 2136 991
rect 2130 986 2136 987
rect 2198 991 2204 992
rect 2198 987 2199 991
rect 2203 987 2204 991
rect 2198 986 2204 987
rect 2270 991 2276 992
rect 2406 991 2412 992
rect 2270 987 2271 991
rect 2275 987 2276 991
rect 2270 986 2276 987
rect 1278 979 1284 980
rect 1278 975 1279 979
rect 1283 975 1284 979
rect 1151 974 1155 975
rect 1151 969 1155 970
rect 1191 974 1195 975
rect 1191 969 1195 970
rect 1239 974 1243 975
rect 1278 974 1284 975
rect 1239 969 1243 970
rect 1150 968 1156 969
rect 1150 964 1151 968
rect 1155 964 1156 968
rect 1150 963 1156 964
rect 1190 968 1196 969
rect 1190 964 1191 968
rect 1195 964 1196 968
rect 1190 963 1196 964
rect 1240 962 1242 969
rect 1238 961 1244 962
rect 1238 957 1239 961
rect 1243 957 1244 961
rect 1280 959 1282 974
rect 1502 972 1508 973
rect 1502 968 1503 972
rect 1507 968 1508 972
rect 1502 967 1508 968
rect 1622 972 1628 973
rect 1622 968 1623 972
rect 1627 968 1628 972
rect 1622 967 1628 968
rect 1734 972 1740 973
rect 1734 968 1735 972
rect 1739 968 1740 972
rect 1734 967 1740 968
rect 1830 972 1836 973
rect 1830 968 1831 972
rect 1835 968 1836 972
rect 1830 967 1836 968
rect 1918 972 1924 973
rect 1918 968 1919 972
rect 1923 968 1924 972
rect 1918 967 1924 968
rect 1998 972 2004 973
rect 1998 968 1999 972
rect 2003 968 2004 972
rect 1998 967 2004 968
rect 2070 972 2076 973
rect 2070 968 2071 972
rect 2075 968 2076 972
rect 2070 967 2076 968
rect 1504 959 1506 967
rect 1624 959 1626 967
rect 1736 959 1738 967
rect 1832 959 1834 967
rect 1920 959 1922 967
rect 2000 959 2002 967
rect 2072 959 2074 967
rect 1238 956 1244 957
rect 1279 958 1283 959
rect 1279 953 1283 954
rect 1319 958 1323 959
rect 1319 953 1323 954
rect 1359 958 1363 959
rect 1359 953 1363 954
rect 1399 958 1403 959
rect 1399 953 1403 954
rect 1463 958 1467 959
rect 1463 953 1467 954
rect 1503 958 1507 959
rect 1503 953 1507 954
rect 1543 958 1547 959
rect 1543 953 1547 954
rect 1623 958 1627 959
rect 1623 953 1627 954
rect 1639 958 1643 959
rect 1639 953 1643 954
rect 1735 958 1739 959
rect 1735 953 1739 954
rect 1831 958 1835 959
rect 1831 953 1835 954
rect 1839 958 1843 959
rect 1839 953 1843 954
rect 1919 958 1923 959
rect 1919 953 1923 954
rect 1935 958 1939 959
rect 1935 953 1939 954
rect 1999 958 2003 959
rect 1999 953 2003 954
rect 2023 958 2027 959
rect 2023 953 2027 954
rect 2071 958 2075 959
rect 2071 953 2075 954
rect 2103 958 2107 959
rect 2103 953 2107 954
rect 654 947 660 948
rect 654 943 655 947
rect 659 943 660 947
rect 654 942 660 943
rect 718 947 724 948
rect 718 943 719 947
rect 723 943 724 947
rect 718 942 724 943
rect 738 947 744 948
rect 738 943 739 947
rect 743 943 744 947
rect 738 942 744 943
rect 1110 947 1116 948
rect 1110 943 1111 947
rect 1115 943 1116 947
rect 1110 942 1116 943
rect 1198 947 1204 948
rect 1198 943 1199 947
rect 1203 943 1204 947
rect 1280 946 1282 953
rect 1318 952 1324 953
rect 1318 948 1319 952
rect 1323 948 1324 952
rect 1318 947 1324 948
rect 1358 952 1364 953
rect 1358 948 1359 952
rect 1363 948 1364 952
rect 1358 947 1364 948
rect 1398 952 1404 953
rect 1398 948 1399 952
rect 1403 948 1404 952
rect 1398 947 1404 948
rect 1462 952 1468 953
rect 1462 948 1463 952
rect 1467 948 1468 952
rect 1462 947 1468 948
rect 1542 952 1548 953
rect 1542 948 1543 952
rect 1547 948 1548 952
rect 1542 947 1548 948
rect 1638 952 1644 953
rect 1638 948 1639 952
rect 1643 948 1644 952
rect 1638 947 1644 948
rect 1734 952 1740 953
rect 1734 948 1735 952
rect 1739 948 1740 952
rect 1734 947 1740 948
rect 1838 952 1844 953
rect 1838 948 1839 952
rect 1843 948 1844 952
rect 1838 947 1844 948
rect 1934 952 1940 953
rect 1934 948 1935 952
rect 1939 948 1940 952
rect 1934 947 1940 948
rect 2022 952 2028 953
rect 2022 948 2023 952
rect 2027 948 2028 952
rect 2022 947 2028 948
rect 2102 952 2108 953
rect 2102 948 2103 952
rect 2107 948 2108 952
rect 2102 947 2108 948
rect 1278 945 1284 946
rect 1198 942 1204 943
rect 1238 944 1244 945
rect 638 921 644 922
rect 638 917 639 921
rect 643 917 644 921
rect 638 916 644 917
rect 656 916 658 942
rect 720 916 722 942
rect 726 921 732 922
rect 726 917 727 921
rect 731 917 732 921
rect 726 916 732 917
rect 296 899 298 916
rect 344 899 346 916
rect 400 899 402 916
rect 472 899 474 916
rect 552 899 554 916
rect 558 915 564 916
rect 558 911 559 915
rect 563 911 564 915
rect 558 910 564 911
rect 574 915 580 916
rect 574 911 575 915
rect 579 911 580 915
rect 574 910 580 911
rect 111 898 115 899
rect 111 893 115 894
rect 255 898 259 899
rect 255 893 259 894
rect 295 898 299 899
rect 295 893 299 894
rect 311 898 315 899
rect 311 893 315 894
rect 343 898 347 899
rect 343 893 347 894
rect 375 898 379 899
rect 375 893 379 894
rect 399 898 403 899
rect 399 893 403 894
rect 455 898 459 899
rect 455 893 459 894
rect 471 898 475 899
rect 471 893 475 894
rect 535 898 539 899
rect 535 893 539 894
rect 551 898 555 899
rect 551 893 555 894
rect 112 861 114 893
rect 256 884 258 893
rect 312 884 314 893
rect 334 887 340 888
rect 254 883 260 884
rect 254 879 255 883
rect 259 879 260 883
rect 254 878 260 879
rect 310 883 316 884
rect 310 879 311 883
rect 315 879 316 883
rect 334 883 335 887
rect 339 883 340 887
rect 376 884 378 893
rect 386 887 392 888
rect 334 882 340 883
rect 374 883 380 884
rect 310 878 316 879
rect 110 860 116 861
rect 110 856 111 860
rect 115 856 116 860
rect 110 855 116 856
rect 110 843 116 844
rect 110 839 111 843
rect 115 839 116 843
rect 110 838 116 839
rect 112 831 114 838
rect 254 836 260 837
rect 254 832 255 836
rect 259 832 260 836
rect 254 831 260 832
rect 310 836 316 837
rect 310 832 311 836
rect 315 832 316 836
rect 310 831 316 832
rect 111 830 115 831
rect 111 825 115 826
rect 191 830 195 831
rect 191 825 195 826
rect 247 830 251 831
rect 247 825 251 826
rect 255 830 259 831
rect 255 825 259 826
rect 311 830 315 831
rect 311 825 315 826
rect 112 818 114 825
rect 190 824 196 825
rect 190 820 191 824
rect 195 820 196 824
rect 190 819 196 820
rect 246 824 252 825
rect 246 820 247 824
rect 251 820 252 824
rect 246 819 252 820
rect 310 824 316 825
rect 310 820 311 824
rect 315 820 316 824
rect 310 819 316 820
rect 110 817 116 818
rect 110 813 111 817
rect 115 813 116 817
rect 110 812 116 813
rect 336 804 338 882
rect 374 879 375 883
rect 379 879 380 883
rect 386 883 387 887
rect 391 883 392 887
rect 456 884 458 893
rect 466 887 472 888
rect 386 882 392 883
rect 454 883 460 884
rect 374 878 380 879
rect 388 864 390 882
rect 454 879 455 883
rect 459 879 460 883
rect 466 883 467 887
rect 471 883 472 887
rect 536 884 538 893
rect 546 887 552 888
rect 466 882 472 883
rect 534 883 540 884
rect 454 878 460 879
rect 386 863 392 864
rect 386 859 387 863
rect 391 859 392 863
rect 386 858 392 859
rect 468 856 470 882
rect 534 879 535 883
rect 539 879 540 883
rect 546 883 547 887
rect 551 883 552 887
rect 546 882 552 883
rect 534 878 540 879
rect 548 856 550 882
rect 560 856 562 910
rect 640 899 642 916
rect 654 915 660 916
rect 654 911 655 915
rect 659 911 660 915
rect 654 910 660 911
rect 718 915 724 916
rect 718 911 719 915
rect 723 911 724 915
rect 718 910 724 911
rect 728 899 730 916
rect 623 898 627 899
rect 623 893 627 894
rect 639 898 643 899
rect 639 893 643 894
rect 711 898 715 899
rect 711 893 715 894
rect 727 898 731 899
rect 727 893 731 894
rect 624 884 626 893
rect 702 887 708 888
rect 622 883 628 884
rect 622 879 623 883
rect 627 879 628 883
rect 702 883 703 887
rect 707 883 708 887
rect 712 884 714 893
rect 740 888 742 942
rect 806 921 812 922
rect 806 917 807 921
rect 811 917 812 921
rect 806 916 812 917
rect 886 921 892 922
rect 886 917 887 921
rect 891 917 892 921
rect 886 916 892 917
rect 958 921 964 922
rect 958 917 959 921
rect 963 917 964 921
rect 958 916 964 917
rect 1022 921 1028 922
rect 1022 917 1023 921
rect 1027 917 1028 921
rect 1022 916 1028 917
rect 1086 921 1092 922
rect 1086 917 1087 921
rect 1091 917 1092 921
rect 1086 916 1092 917
rect 1150 921 1156 922
rect 1150 917 1151 921
rect 1155 917 1156 921
rect 1150 916 1156 917
rect 1190 921 1196 922
rect 1190 917 1191 921
rect 1195 917 1196 921
rect 1190 916 1196 917
rect 1200 916 1202 942
rect 1238 940 1239 944
rect 1243 940 1244 944
rect 1278 941 1279 945
rect 1283 941 1284 945
rect 1278 940 1284 941
rect 1214 939 1220 940
rect 1238 939 1244 940
rect 1214 935 1215 939
rect 1219 935 1220 939
rect 1214 934 1220 935
rect 1216 916 1218 934
rect 808 899 810 916
rect 888 899 890 916
rect 960 899 962 916
rect 1024 899 1026 916
rect 1078 915 1084 916
rect 1078 911 1079 915
rect 1083 911 1084 915
rect 1078 910 1084 911
rect 791 898 795 899
rect 791 893 795 894
rect 807 898 811 899
rect 807 893 811 894
rect 863 898 867 899
rect 863 893 867 894
rect 887 898 891 899
rect 887 893 891 894
rect 935 898 939 899
rect 935 893 939 894
rect 959 898 963 899
rect 959 893 963 894
rect 999 898 1003 899
rect 999 893 1003 894
rect 1023 898 1027 899
rect 1023 893 1027 894
rect 1055 898 1059 899
rect 1055 893 1059 894
rect 738 887 744 888
rect 702 882 708 883
rect 710 883 716 884
rect 622 878 628 879
rect 704 856 706 882
rect 710 879 711 883
rect 715 879 716 883
rect 738 883 739 887
rect 743 883 744 887
rect 792 884 794 893
rect 854 887 860 888
rect 738 882 744 883
rect 790 883 796 884
rect 710 878 716 879
rect 790 879 791 883
rect 795 879 796 883
rect 854 883 855 887
rect 859 883 860 887
rect 864 884 866 893
rect 918 887 924 888
rect 854 882 860 883
rect 862 883 868 884
rect 790 878 796 879
rect 856 856 858 882
rect 862 879 863 883
rect 867 879 868 883
rect 918 883 919 887
rect 923 883 924 887
rect 936 884 938 893
rect 946 887 952 888
rect 918 882 924 883
rect 934 883 940 884
rect 862 878 868 879
rect 466 855 472 856
rect 466 851 467 855
rect 471 851 472 855
rect 466 850 472 851
rect 546 855 552 856
rect 546 851 547 855
rect 551 851 552 855
rect 546 850 552 851
rect 558 855 564 856
rect 558 851 559 855
rect 563 851 564 855
rect 558 850 564 851
rect 638 855 644 856
rect 638 851 639 855
rect 643 851 644 855
rect 638 850 644 851
rect 702 855 708 856
rect 702 851 703 855
rect 707 851 708 855
rect 702 850 708 851
rect 854 855 860 856
rect 854 851 855 855
rect 859 851 860 855
rect 854 850 860 851
rect 374 836 380 837
rect 374 832 375 836
rect 379 832 380 836
rect 374 831 380 832
rect 454 836 460 837
rect 454 832 455 836
rect 459 832 460 836
rect 454 831 460 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 622 836 628 837
rect 622 832 623 836
rect 627 832 628 836
rect 622 831 628 832
rect 375 830 379 831
rect 375 825 379 826
rect 383 830 387 831
rect 383 825 387 826
rect 455 830 459 831
rect 455 825 459 826
rect 463 830 467 831
rect 463 825 467 826
rect 535 830 539 831
rect 535 825 539 826
rect 543 830 547 831
rect 543 825 547 826
rect 615 830 619 831
rect 615 825 619 826
rect 623 830 627 831
rect 623 825 627 826
rect 382 824 388 825
rect 382 820 383 824
rect 387 820 388 824
rect 382 819 388 820
rect 462 824 468 825
rect 462 820 463 824
rect 467 820 468 824
rect 462 819 468 820
rect 542 824 548 825
rect 542 820 543 824
rect 547 820 548 824
rect 542 819 548 820
rect 614 824 620 825
rect 614 820 615 824
rect 619 820 620 824
rect 614 819 620 820
rect 270 803 276 804
rect 270 802 271 803
rect 110 800 116 801
rect 110 796 111 800
rect 115 796 116 800
rect 110 795 116 796
rect 264 800 271 802
rect 112 763 114 795
rect 190 777 196 778
rect 190 773 191 777
rect 195 773 196 777
rect 190 772 196 773
rect 246 777 252 778
rect 246 773 247 777
rect 251 773 252 777
rect 246 772 252 773
rect 264 772 266 800
rect 270 799 271 800
rect 275 799 276 803
rect 270 798 276 799
rect 334 803 340 804
rect 334 799 335 803
rect 339 799 340 803
rect 334 798 340 799
rect 346 803 352 804
rect 346 799 347 803
rect 351 799 352 803
rect 346 798 352 799
rect 518 803 524 804
rect 518 799 519 803
rect 523 799 524 803
rect 518 798 524 799
rect 526 803 532 804
rect 526 799 527 803
rect 531 799 532 803
rect 526 798 532 799
rect 310 777 316 778
rect 310 773 311 777
rect 315 773 316 777
rect 310 772 316 773
rect 348 772 350 798
rect 406 795 412 796
rect 406 791 407 795
rect 411 791 412 795
rect 406 790 412 791
rect 382 777 388 778
rect 382 773 383 777
rect 387 773 388 777
rect 382 772 388 773
rect 408 772 410 790
rect 462 777 468 778
rect 462 773 463 777
rect 467 773 468 777
rect 462 772 468 773
rect 192 763 194 772
rect 248 763 250 772
rect 262 771 268 772
rect 262 767 263 771
rect 267 767 268 771
rect 262 766 268 767
rect 302 771 308 772
rect 302 767 303 771
rect 307 767 308 771
rect 302 766 308 767
rect 111 762 115 763
rect 111 757 115 758
rect 135 762 139 763
rect 135 757 139 758
rect 175 762 179 763
rect 175 757 179 758
rect 191 762 195 763
rect 191 757 195 758
rect 215 762 219 763
rect 215 757 219 758
rect 247 762 251 763
rect 247 757 251 758
rect 279 762 283 763
rect 279 757 283 758
rect 112 725 114 757
rect 136 748 138 757
rect 162 751 168 752
rect 134 747 140 748
rect 134 743 135 747
rect 139 743 140 747
rect 162 747 163 751
rect 167 747 168 751
rect 176 748 178 757
rect 198 751 204 752
rect 162 746 168 747
rect 174 747 180 748
rect 134 742 140 743
rect 164 728 166 746
rect 174 743 175 747
rect 179 743 180 747
rect 198 747 199 751
rect 203 747 204 751
rect 216 748 218 757
rect 280 748 282 757
rect 198 746 204 747
rect 214 747 220 748
rect 174 742 180 743
rect 162 727 168 728
rect 110 724 116 725
rect 110 720 111 724
rect 115 720 116 724
rect 162 723 163 727
rect 167 723 168 727
rect 162 722 168 723
rect 110 719 116 720
rect 110 707 116 708
rect 110 703 111 707
rect 115 703 116 707
rect 110 702 116 703
rect 112 687 114 702
rect 134 700 140 701
rect 134 696 135 700
rect 139 696 140 700
rect 134 695 140 696
rect 174 700 180 701
rect 174 696 175 700
rect 179 696 180 700
rect 174 695 180 696
rect 136 687 138 695
rect 176 687 178 695
rect 111 686 115 687
rect 111 681 115 682
rect 135 686 139 687
rect 135 681 139 682
rect 175 686 179 687
rect 175 681 179 682
rect 112 674 114 681
rect 134 680 140 681
rect 134 676 135 680
rect 139 676 140 680
rect 134 675 140 676
rect 174 680 180 681
rect 174 676 175 680
rect 179 676 180 680
rect 174 675 180 676
rect 110 673 116 674
rect 110 669 111 673
rect 115 669 116 673
rect 110 668 116 669
rect 200 660 202 746
rect 214 743 215 747
rect 219 743 220 747
rect 214 742 220 743
rect 278 747 284 748
rect 278 743 279 747
rect 283 743 284 747
rect 278 742 284 743
rect 304 720 306 766
rect 312 763 314 772
rect 346 771 352 772
rect 346 767 347 771
rect 351 767 352 771
rect 346 766 352 767
rect 384 763 386 772
rect 406 771 412 772
rect 406 767 407 771
rect 411 767 412 771
rect 406 766 412 767
rect 464 763 466 772
rect 311 762 315 763
rect 311 757 315 758
rect 351 762 355 763
rect 351 757 355 758
rect 383 762 387 763
rect 383 757 387 758
rect 423 762 427 763
rect 423 757 427 758
rect 463 762 467 763
rect 463 757 467 758
rect 495 762 499 763
rect 495 757 499 758
rect 342 751 348 752
rect 342 747 343 751
rect 347 747 348 751
rect 352 748 354 757
rect 362 751 368 752
rect 342 746 348 747
rect 350 747 356 748
rect 344 720 346 746
rect 350 743 351 747
rect 355 743 356 747
rect 362 747 363 751
rect 367 747 368 751
rect 424 748 426 757
rect 486 751 492 752
rect 362 746 368 747
rect 422 747 428 748
rect 350 742 356 743
rect 364 728 366 746
rect 422 743 423 747
rect 427 743 428 747
rect 486 747 487 751
rect 491 747 492 751
rect 496 748 498 757
rect 520 752 522 798
rect 528 772 530 798
rect 542 777 548 778
rect 542 773 543 777
rect 547 773 548 777
rect 542 772 548 773
rect 614 777 620 778
rect 614 773 615 777
rect 619 773 620 777
rect 614 772 620 773
rect 640 772 642 850
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 790 836 796 837
rect 790 832 791 836
rect 795 832 796 836
rect 790 831 796 832
rect 862 836 868 837
rect 862 832 863 836
rect 867 832 868 836
rect 862 831 868 832
rect 687 830 691 831
rect 687 825 691 826
rect 711 830 715 831
rect 711 825 715 826
rect 751 830 755 831
rect 751 825 755 826
rect 791 830 795 831
rect 791 825 795 826
rect 815 830 819 831
rect 815 825 819 826
rect 863 830 867 831
rect 863 825 867 826
rect 871 830 875 831
rect 871 825 875 826
rect 686 824 692 825
rect 686 820 687 824
rect 691 820 692 824
rect 686 819 692 820
rect 750 824 756 825
rect 750 820 751 824
rect 755 820 756 824
rect 750 819 756 820
rect 814 824 820 825
rect 814 820 815 824
rect 819 820 820 824
rect 814 819 820 820
rect 870 824 876 825
rect 870 820 871 824
rect 875 820 876 824
rect 870 819 876 820
rect 920 804 922 882
rect 934 879 935 883
rect 939 879 940 883
rect 946 883 947 887
rect 951 883 952 887
rect 1000 884 1002 893
rect 1010 887 1016 888
rect 946 882 952 883
rect 998 883 1004 884
rect 934 878 940 879
rect 948 864 950 882
rect 998 879 999 883
rect 1003 879 1004 883
rect 1010 883 1011 887
rect 1015 883 1016 887
rect 1056 884 1058 893
rect 1010 882 1016 883
rect 1054 883 1060 884
rect 998 878 1004 879
rect 946 863 952 864
rect 946 859 947 863
rect 951 859 952 863
rect 946 858 952 859
rect 1012 856 1014 882
rect 1054 879 1055 883
rect 1059 879 1060 883
rect 1054 878 1060 879
rect 1080 856 1082 910
rect 1088 899 1090 916
rect 1152 899 1154 916
rect 1192 899 1194 916
rect 1198 915 1204 916
rect 1198 911 1199 915
rect 1203 911 1204 915
rect 1198 910 1204 911
rect 1214 915 1220 916
rect 1214 911 1215 915
rect 1219 911 1220 915
rect 1214 910 1220 911
rect 1240 899 1242 939
rect 1346 931 1352 932
rect 1278 928 1284 929
rect 1278 924 1279 928
rect 1283 924 1284 928
rect 1346 927 1347 931
rect 1351 927 1352 931
rect 1346 926 1352 927
rect 1366 931 1372 932
rect 1366 927 1367 931
rect 1371 927 1372 931
rect 1366 926 1372 927
rect 1406 931 1412 932
rect 1406 927 1407 931
rect 1411 927 1412 931
rect 1406 926 1412 927
rect 1490 931 1496 932
rect 1490 927 1491 931
rect 1495 927 1496 931
rect 1490 926 1496 927
rect 1986 931 1992 932
rect 1986 927 1987 931
rect 1991 927 1992 931
rect 1986 926 1992 927
rect 1278 923 1284 924
rect 1087 898 1091 899
rect 1087 893 1091 894
rect 1119 898 1123 899
rect 1119 893 1123 894
rect 1151 898 1155 899
rect 1151 893 1155 894
rect 1183 898 1187 899
rect 1183 893 1187 894
rect 1191 898 1195 899
rect 1191 893 1195 894
rect 1239 898 1243 899
rect 1239 893 1243 894
rect 1110 887 1116 888
rect 1110 883 1111 887
rect 1115 883 1116 887
rect 1120 884 1122 893
rect 1174 887 1180 888
rect 1110 882 1116 883
rect 1118 883 1124 884
rect 1112 856 1114 882
rect 1118 879 1119 883
rect 1123 879 1124 883
rect 1174 883 1175 887
rect 1179 883 1180 887
rect 1184 884 1186 893
rect 1194 887 1200 888
rect 1174 882 1180 883
rect 1182 883 1188 884
rect 1118 878 1124 879
rect 1176 856 1178 882
rect 1182 879 1183 883
rect 1187 879 1188 883
rect 1194 883 1195 887
rect 1199 883 1200 887
rect 1194 882 1200 883
rect 1182 878 1188 879
rect 1196 864 1198 882
rect 1194 863 1200 864
rect 1194 859 1195 863
rect 1199 859 1200 863
rect 1240 861 1242 893
rect 1280 883 1282 923
rect 1318 905 1324 906
rect 1318 901 1319 905
rect 1323 901 1324 905
rect 1318 900 1324 901
rect 1320 883 1322 900
rect 1279 882 1283 883
rect 1279 877 1283 878
rect 1319 882 1323 883
rect 1319 877 1323 878
rect 1335 882 1339 883
rect 1348 880 1350 926
rect 1358 905 1364 906
rect 1358 901 1359 905
rect 1363 901 1364 905
rect 1358 900 1364 901
rect 1368 900 1370 926
rect 1398 905 1404 906
rect 1398 901 1399 905
rect 1403 901 1404 905
rect 1398 900 1404 901
rect 1408 900 1410 926
rect 1426 923 1432 924
rect 1426 919 1427 923
rect 1431 919 1432 923
rect 1426 918 1432 919
rect 1428 900 1430 918
rect 1462 905 1468 906
rect 1462 901 1463 905
rect 1467 901 1468 905
rect 1462 900 1468 901
rect 1360 883 1362 900
rect 1366 899 1372 900
rect 1366 895 1367 899
rect 1371 895 1372 899
rect 1366 894 1372 895
rect 1400 883 1402 900
rect 1406 899 1412 900
rect 1406 895 1407 899
rect 1411 895 1412 899
rect 1406 894 1412 895
rect 1426 899 1432 900
rect 1426 895 1427 899
rect 1431 895 1432 899
rect 1426 894 1432 895
rect 1464 883 1466 900
rect 1359 882 1363 883
rect 1335 877 1339 878
rect 1346 879 1352 880
rect 1194 858 1200 859
rect 1238 860 1244 861
rect 1238 856 1239 860
rect 1243 856 1244 860
rect 1010 855 1016 856
rect 1010 851 1011 855
rect 1015 851 1016 855
rect 1010 850 1016 851
rect 1078 855 1084 856
rect 1078 851 1079 855
rect 1083 851 1084 855
rect 1078 850 1084 851
rect 1110 855 1116 856
rect 1110 851 1111 855
rect 1115 851 1116 855
rect 1110 850 1116 851
rect 1174 855 1180 856
rect 1238 855 1244 856
rect 1174 851 1175 855
rect 1179 851 1180 855
rect 1174 850 1180 851
rect 1280 845 1282 877
rect 1336 868 1338 877
rect 1346 875 1347 879
rect 1351 875 1352 879
rect 1359 877 1363 878
rect 1375 882 1379 883
rect 1375 877 1379 878
rect 1399 882 1403 883
rect 1399 877 1403 878
rect 1415 882 1419 883
rect 1415 877 1419 878
rect 1463 882 1467 883
rect 1463 877 1467 878
rect 1471 882 1475 883
rect 1471 877 1475 878
rect 1346 874 1352 875
rect 1362 871 1368 872
rect 1334 867 1340 868
rect 1334 863 1335 867
rect 1339 863 1340 867
rect 1362 867 1363 871
rect 1367 867 1368 871
rect 1376 868 1378 877
rect 1402 871 1408 872
rect 1362 866 1368 867
rect 1374 867 1380 868
rect 1334 862 1340 863
rect 1278 844 1284 845
rect 1238 843 1244 844
rect 1238 839 1239 843
rect 1243 839 1244 843
rect 1278 840 1279 844
rect 1283 840 1284 844
rect 1278 839 1284 840
rect 1350 839 1356 840
rect 1238 838 1244 839
rect 934 836 940 837
rect 934 832 935 836
rect 939 832 940 836
rect 934 831 940 832
rect 998 836 1004 837
rect 998 832 999 836
rect 1003 832 1004 836
rect 998 831 1004 832
rect 1054 836 1060 837
rect 1054 832 1055 836
rect 1059 832 1060 836
rect 1054 831 1060 832
rect 1118 836 1124 837
rect 1118 832 1119 836
rect 1123 832 1124 836
rect 1118 831 1124 832
rect 1182 836 1188 837
rect 1182 832 1183 836
rect 1187 832 1188 836
rect 1182 831 1188 832
rect 1240 831 1242 838
rect 1350 835 1351 839
rect 1355 835 1356 839
rect 1364 838 1366 866
rect 1374 863 1375 867
rect 1379 863 1380 867
rect 1402 867 1403 871
rect 1407 867 1408 871
rect 1416 868 1418 877
rect 1472 868 1474 877
rect 1492 872 1494 926
rect 1542 905 1548 906
rect 1542 901 1543 905
rect 1547 901 1548 905
rect 1542 900 1548 901
rect 1638 905 1644 906
rect 1638 901 1639 905
rect 1643 901 1644 905
rect 1638 900 1644 901
rect 1734 905 1740 906
rect 1734 901 1735 905
rect 1739 901 1740 905
rect 1734 900 1740 901
rect 1838 905 1844 906
rect 1838 901 1839 905
rect 1843 901 1844 905
rect 1838 900 1844 901
rect 1934 905 1940 906
rect 1934 901 1935 905
rect 1939 901 1940 905
rect 1934 900 1940 901
rect 1988 900 1990 926
rect 2022 905 2028 906
rect 2022 901 2023 905
rect 2027 901 2028 905
rect 2022 900 2028 901
rect 2102 905 2108 906
rect 2102 901 2103 905
rect 2107 901 2108 905
rect 2102 900 2108 901
rect 2132 900 2134 986
rect 2406 979 2412 980
rect 2406 975 2407 979
rect 2411 975 2412 979
rect 2406 974 2412 975
rect 2142 972 2148 973
rect 2142 968 2143 972
rect 2147 968 2148 972
rect 2142 967 2148 968
rect 2206 972 2212 973
rect 2206 968 2207 972
rect 2211 968 2212 972
rect 2206 967 2212 968
rect 2278 972 2284 973
rect 2278 968 2279 972
rect 2283 968 2284 972
rect 2278 967 2284 968
rect 2144 959 2146 967
rect 2208 959 2210 967
rect 2280 959 2282 967
rect 2408 959 2410 974
rect 2143 958 2147 959
rect 2143 953 2147 954
rect 2175 958 2179 959
rect 2175 953 2179 954
rect 2207 958 2211 959
rect 2207 953 2211 954
rect 2239 958 2243 959
rect 2239 953 2243 954
rect 2279 958 2283 959
rect 2279 953 2283 954
rect 2311 958 2315 959
rect 2311 953 2315 954
rect 2359 958 2363 959
rect 2359 953 2363 954
rect 2407 958 2411 959
rect 2407 953 2411 954
rect 2174 952 2180 953
rect 2174 948 2175 952
rect 2179 948 2180 952
rect 2174 947 2180 948
rect 2238 952 2244 953
rect 2238 948 2239 952
rect 2243 948 2244 952
rect 2238 947 2244 948
rect 2310 952 2316 953
rect 2310 948 2311 952
rect 2315 948 2316 952
rect 2310 947 2316 948
rect 2358 952 2364 953
rect 2358 948 2359 952
rect 2363 948 2364 952
rect 2358 947 2364 948
rect 2408 946 2410 953
rect 2406 945 2412 946
rect 2406 941 2407 945
rect 2411 941 2412 945
rect 2406 940 2412 941
rect 2254 931 2260 932
rect 2254 927 2255 931
rect 2259 927 2260 931
rect 2254 926 2260 927
rect 2326 931 2332 932
rect 2326 927 2327 931
rect 2331 927 2332 931
rect 2326 926 2332 927
rect 2374 931 2380 932
rect 2374 927 2375 931
rect 2379 927 2380 931
rect 2374 926 2380 927
rect 2382 931 2388 932
rect 2382 927 2383 931
rect 2387 927 2388 931
rect 2382 926 2388 927
rect 2406 928 2412 929
rect 2198 923 2204 924
rect 2198 919 2199 923
rect 2203 919 2204 923
rect 2198 918 2204 919
rect 2174 905 2180 906
rect 2174 901 2175 905
rect 2179 901 2180 905
rect 2174 900 2180 901
rect 2200 900 2202 918
rect 2238 905 2244 906
rect 2238 901 2239 905
rect 2243 901 2244 905
rect 2238 900 2244 901
rect 2256 900 2258 926
rect 2310 905 2316 906
rect 2310 901 2311 905
rect 2315 901 2316 905
rect 2310 900 2316 901
rect 2328 900 2330 926
rect 2358 905 2364 906
rect 2358 901 2359 905
rect 2363 901 2364 905
rect 2358 900 2364 901
rect 2376 900 2378 926
rect 1544 883 1546 900
rect 1640 883 1642 900
rect 1736 883 1738 900
rect 1778 899 1784 900
rect 1778 895 1779 899
rect 1783 895 1784 899
rect 1778 894 1784 895
rect 1535 882 1539 883
rect 1535 877 1539 878
rect 1543 882 1547 883
rect 1543 877 1547 878
rect 1607 882 1611 883
rect 1607 877 1611 878
rect 1639 882 1643 883
rect 1639 877 1643 878
rect 1679 882 1683 883
rect 1679 877 1683 878
rect 1735 882 1739 883
rect 1735 877 1739 878
rect 1751 882 1755 883
rect 1751 877 1755 878
rect 1490 871 1496 872
rect 1402 866 1408 867
rect 1414 867 1420 868
rect 1374 862 1380 863
rect 1370 839 1376 840
rect 1370 838 1371 839
rect 1364 836 1371 838
rect 1350 834 1356 835
rect 1370 835 1371 836
rect 1375 835 1376 839
rect 1404 838 1406 866
rect 1414 863 1415 867
rect 1419 863 1420 867
rect 1414 862 1420 863
rect 1470 867 1476 868
rect 1470 863 1471 867
rect 1475 863 1476 867
rect 1490 867 1491 871
rect 1495 867 1496 871
rect 1536 868 1538 877
rect 1546 871 1552 872
rect 1490 866 1496 867
rect 1534 867 1540 868
rect 1470 862 1476 863
rect 1534 863 1535 867
rect 1539 863 1540 867
rect 1546 867 1547 871
rect 1551 867 1552 871
rect 1608 868 1610 877
rect 1646 871 1652 872
rect 1546 866 1552 867
rect 1606 867 1612 868
rect 1534 862 1540 863
rect 1548 840 1550 866
rect 1606 863 1607 867
rect 1611 863 1612 867
rect 1646 867 1647 871
rect 1651 867 1652 871
rect 1680 868 1682 877
rect 1690 871 1696 872
rect 1646 866 1652 867
rect 1678 867 1684 868
rect 1606 862 1612 863
rect 1410 839 1416 840
rect 1410 838 1411 839
rect 1404 836 1411 838
rect 1370 834 1376 835
rect 1410 835 1411 836
rect 1415 835 1416 839
rect 1410 834 1416 835
rect 1546 839 1552 840
rect 1546 835 1547 839
rect 1551 835 1552 839
rect 1546 834 1552 835
rect 1574 839 1580 840
rect 1574 835 1575 839
rect 1579 835 1580 839
rect 1574 834 1580 835
rect 927 830 931 831
rect 927 825 931 826
rect 935 830 939 831
rect 935 825 939 826
rect 983 830 987 831
rect 983 825 987 826
rect 999 830 1003 831
rect 999 825 1003 826
rect 1047 830 1051 831
rect 1047 825 1051 826
rect 1055 830 1059 831
rect 1055 825 1059 826
rect 1119 830 1123 831
rect 1119 825 1123 826
rect 1183 830 1187 831
rect 1183 825 1187 826
rect 1239 830 1243 831
rect 1239 825 1243 826
rect 1278 827 1284 828
rect 926 824 932 825
rect 926 820 927 824
rect 931 820 932 824
rect 926 819 932 820
rect 982 824 988 825
rect 982 820 983 824
rect 987 820 988 824
rect 982 819 988 820
rect 1046 824 1052 825
rect 1046 820 1047 824
rect 1051 820 1052 824
rect 1046 819 1052 820
rect 1240 818 1242 825
rect 1278 823 1279 827
rect 1283 823 1284 827
rect 1278 822 1284 823
rect 1238 817 1244 818
rect 1238 813 1239 817
rect 1243 813 1244 817
rect 1238 812 1244 813
rect 1280 811 1282 822
rect 1334 820 1340 821
rect 1334 816 1335 820
rect 1339 816 1340 820
rect 1334 815 1340 816
rect 1336 811 1338 815
rect 1279 810 1283 811
rect 1279 805 1283 806
rect 1303 810 1307 811
rect 1303 805 1307 806
rect 1335 810 1339 811
rect 1335 805 1339 806
rect 1343 810 1347 811
rect 1343 805 1347 806
rect 918 803 924 804
rect 918 799 919 803
rect 923 799 924 803
rect 918 798 924 799
rect 1238 800 1244 801
rect 1238 796 1239 800
rect 1243 796 1244 800
rect 1280 798 1282 805
rect 1302 804 1308 805
rect 1302 800 1303 804
rect 1307 800 1308 804
rect 1302 799 1308 800
rect 1342 804 1348 805
rect 1342 800 1343 804
rect 1347 800 1348 804
rect 1342 799 1348 800
rect 894 795 900 796
rect 894 791 895 795
rect 899 791 900 795
rect 894 790 900 791
rect 1070 795 1076 796
rect 1238 795 1244 796
rect 1278 797 1284 798
rect 1070 791 1071 795
rect 1075 791 1076 795
rect 1070 790 1076 791
rect 686 777 692 778
rect 686 773 687 777
rect 691 773 692 777
rect 686 772 692 773
rect 750 777 756 778
rect 750 773 751 777
rect 755 773 756 777
rect 750 772 756 773
rect 814 777 820 778
rect 814 773 815 777
rect 819 773 820 777
rect 814 772 820 773
rect 870 777 876 778
rect 870 773 871 777
rect 875 773 876 777
rect 870 772 876 773
rect 896 772 898 790
rect 926 777 932 778
rect 926 773 927 777
rect 931 773 932 777
rect 926 772 932 773
rect 982 777 988 778
rect 982 773 983 777
rect 987 773 988 777
rect 982 772 988 773
rect 1046 777 1052 778
rect 1046 773 1047 777
rect 1051 773 1052 777
rect 1046 772 1052 773
rect 1072 772 1074 790
rect 526 771 532 772
rect 526 767 527 771
rect 531 767 532 771
rect 526 766 532 767
rect 544 763 546 772
rect 616 763 618 772
rect 638 771 644 772
rect 638 767 639 771
rect 643 767 644 771
rect 638 766 644 767
rect 688 763 690 772
rect 752 763 754 772
rect 816 763 818 772
rect 872 763 874 772
rect 886 771 892 772
rect 886 767 887 771
rect 891 767 892 771
rect 886 766 892 767
rect 894 771 900 772
rect 894 767 895 771
rect 899 767 900 771
rect 894 766 900 767
rect 543 762 547 763
rect 543 757 547 758
rect 559 762 563 763
rect 559 757 563 758
rect 615 762 619 763
rect 615 757 619 758
rect 623 762 627 763
rect 623 757 627 758
rect 687 762 691 763
rect 687 757 691 758
rect 695 762 699 763
rect 695 757 699 758
rect 751 762 755 763
rect 751 757 755 758
rect 783 762 787 763
rect 783 757 787 758
rect 815 762 819 763
rect 815 757 819 758
rect 871 762 875 763
rect 871 757 875 758
rect 879 762 883 763
rect 879 757 883 758
rect 518 751 524 752
rect 486 746 492 747
rect 494 747 500 748
rect 422 742 428 743
rect 362 727 368 728
rect 362 723 363 727
rect 367 723 368 727
rect 362 722 368 723
rect 488 720 490 746
rect 494 743 495 747
rect 499 743 500 747
rect 518 747 519 751
rect 523 747 524 751
rect 560 748 562 757
rect 614 751 620 752
rect 518 746 524 747
rect 558 747 564 748
rect 494 742 500 743
rect 558 743 559 747
rect 563 743 564 747
rect 614 747 615 751
rect 619 747 620 751
rect 624 748 626 757
rect 686 751 692 752
rect 614 746 620 747
rect 622 747 628 748
rect 558 742 564 743
rect 616 720 618 746
rect 622 743 623 747
rect 627 743 628 747
rect 686 747 687 751
rect 691 747 692 751
rect 696 748 698 757
rect 758 751 764 752
rect 686 746 692 747
rect 694 747 700 748
rect 622 742 628 743
rect 688 720 690 746
rect 694 743 695 747
rect 699 743 700 747
rect 758 747 759 751
rect 763 747 764 751
rect 784 748 786 757
rect 794 751 800 752
rect 758 746 764 747
rect 782 747 788 748
rect 694 742 700 743
rect 302 719 308 720
rect 302 715 303 719
rect 307 715 308 719
rect 302 714 308 715
rect 342 719 348 720
rect 342 715 343 719
rect 347 715 348 719
rect 342 714 348 715
rect 438 719 444 720
rect 438 715 439 719
rect 443 715 444 719
rect 438 714 444 715
rect 486 719 492 720
rect 486 715 487 719
rect 491 715 492 719
rect 486 714 492 715
rect 614 719 620 720
rect 614 715 615 719
rect 619 715 620 719
rect 614 714 620 715
rect 686 719 692 720
rect 686 715 687 719
rect 691 715 692 719
rect 686 714 692 715
rect 214 700 220 701
rect 214 696 215 700
rect 219 696 220 700
rect 214 695 220 696
rect 278 700 284 701
rect 278 696 279 700
rect 283 696 284 700
rect 278 695 284 696
rect 350 700 356 701
rect 350 696 351 700
rect 355 696 356 700
rect 350 695 356 696
rect 422 700 428 701
rect 422 696 423 700
rect 427 696 428 700
rect 422 695 428 696
rect 216 687 218 695
rect 280 687 282 695
rect 352 687 354 695
rect 424 687 426 695
rect 215 686 219 687
rect 215 681 219 682
rect 231 686 235 687
rect 231 681 235 682
rect 279 686 283 687
rect 279 681 283 682
rect 287 686 291 687
rect 287 681 291 682
rect 343 686 347 687
rect 343 681 347 682
rect 351 686 355 687
rect 351 681 355 682
rect 399 686 403 687
rect 399 681 403 682
rect 423 686 427 687
rect 423 681 427 682
rect 230 680 236 681
rect 230 676 231 680
rect 235 676 236 680
rect 230 675 236 676
rect 286 680 292 681
rect 286 676 287 680
rect 291 676 292 680
rect 286 675 292 676
rect 342 680 348 681
rect 342 676 343 680
rect 347 676 348 680
rect 342 675 348 676
rect 398 680 404 681
rect 398 676 399 680
rect 403 676 404 680
rect 398 675 404 676
rect 198 659 204 660
rect 110 656 116 657
rect 110 652 111 656
rect 115 652 116 656
rect 198 655 199 659
rect 203 655 204 659
rect 198 654 204 655
rect 210 659 216 660
rect 210 655 211 659
rect 215 655 216 659
rect 210 654 216 655
rect 110 651 116 652
rect 112 619 114 651
rect 134 633 140 634
rect 134 629 135 633
rect 139 629 140 633
rect 134 628 140 629
rect 174 633 180 634
rect 174 629 175 633
rect 179 629 180 633
rect 174 628 180 629
rect 212 628 214 654
rect 310 651 316 652
rect 310 647 311 651
rect 315 647 316 651
rect 310 646 316 647
rect 230 633 236 634
rect 230 629 231 633
rect 235 629 236 633
rect 230 628 236 629
rect 286 633 292 634
rect 286 629 287 633
rect 291 629 292 633
rect 286 628 292 629
rect 312 628 314 646
rect 342 633 348 634
rect 342 629 343 633
rect 347 629 348 633
rect 342 628 348 629
rect 398 633 404 634
rect 398 629 399 633
rect 403 629 404 633
rect 398 628 404 629
rect 440 628 442 714
rect 494 700 500 701
rect 494 696 495 700
rect 499 696 500 700
rect 494 695 500 696
rect 558 700 564 701
rect 558 696 559 700
rect 563 696 564 700
rect 558 695 564 696
rect 622 700 628 701
rect 622 696 623 700
rect 627 696 628 700
rect 622 695 628 696
rect 694 700 700 701
rect 694 696 695 700
rect 699 696 700 700
rect 694 695 700 696
rect 496 687 498 695
rect 560 687 562 695
rect 624 687 626 695
rect 696 687 698 695
rect 455 686 459 687
rect 455 681 459 682
rect 495 686 499 687
rect 495 681 499 682
rect 503 686 507 687
rect 503 681 507 682
rect 559 686 563 687
rect 559 681 563 682
rect 623 686 627 687
rect 623 681 627 682
rect 695 686 699 687
rect 695 681 699 682
rect 454 680 460 681
rect 454 676 455 680
rect 459 676 460 680
rect 454 675 460 676
rect 502 680 508 681
rect 502 676 503 680
rect 507 676 508 680
rect 502 675 508 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 694 680 700 681
rect 694 676 695 680
rect 699 676 700 680
rect 694 675 700 676
rect 760 660 762 746
rect 782 743 783 747
rect 787 743 788 747
rect 794 747 795 751
rect 799 747 800 751
rect 880 748 882 757
rect 794 746 800 747
rect 878 747 884 748
rect 782 742 788 743
rect 796 728 798 746
rect 878 743 879 747
rect 883 743 884 747
rect 878 742 884 743
rect 794 727 800 728
rect 794 723 795 727
rect 799 723 800 727
rect 794 722 800 723
rect 888 720 890 766
rect 928 763 930 772
rect 984 763 986 772
rect 1048 763 1050 772
rect 1070 771 1076 772
rect 1070 767 1071 771
rect 1075 767 1076 771
rect 1070 766 1076 767
rect 1240 763 1242 795
rect 1278 793 1279 797
rect 1283 793 1284 797
rect 1278 792 1284 793
rect 1278 780 1284 781
rect 1278 776 1279 780
rect 1283 776 1284 780
rect 1278 775 1284 776
rect 927 762 931 763
rect 927 757 931 758
rect 983 762 987 763
rect 983 757 987 758
rect 1047 762 1051 763
rect 1047 757 1051 758
rect 1095 762 1099 763
rect 1095 757 1099 758
rect 1191 762 1195 763
rect 1191 757 1195 758
rect 1239 762 1243 763
rect 1239 757 1243 758
rect 974 751 980 752
rect 974 747 975 751
rect 979 747 980 751
rect 984 748 986 757
rect 1086 751 1092 752
rect 974 746 980 747
rect 982 747 988 748
rect 976 720 978 746
rect 982 743 983 747
rect 987 743 988 747
rect 1086 747 1087 751
rect 1091 747 1092 751
rect 1096 748 1098 757
rect 1106 751 1112 752
rect 1086 746 1092 747
rect 1094 747 1100 748
rect 982 742 988 743
rect 1088 720 1090 746
rect 1094 743 1095 747
rect 1099 743 1100 747
rect 1106 747 1107 751
rect 1111 747 1112 751
rect 1192 748 1194 757
rect 1106 746 1112 747
rect 1190 747 1196 748
rect 1094 742 1100 743
rect 1108 728 1110 746
rect 1190 743 1191 747
rect 1195 743 1196 747
rect 1190 742 1196 743
rect 1106 727 1112 728
rect 1106 723 1107 727
rect 1111 723 1112 727
rect 1240 725 1242 757
rect 1280 743 1282 775
rect 1302 757 1308 758
rect 1302 753 1303 757
rect 1307 753 1308 757
rect 1302 752 1308 753
rect 1342 757 1348 758
rect 1342 753 1343 757
rect 1347 753 1348 757
rect 1342 752 1348 753
rect 1352 752 1354 834
rect 1374 820 1380 821
rect 1374 816 1375 820
rect 1379 816 1380 820
rect 1374 815 1380 816
rect 1414 820 1420 821
rect 1414 816 1415 820
rect 1419 816 1420 820
rect 1414 815 1420 816
rect 1470 820 1476 821
rect 1470 816 1471 820
rect 1475 816 1476 820
rect 1470 815 1476 816
rect 1534 820 1540 821
rect 1534 816 1535 820
rect 1539 816 1540 820
rect 1534 815 1540 816
rect 1376 811 1378 815
rect 1416 811 1418 815
rect 1472 811 1474 815
rect 1536 811 1538 815
rect 1375 810 1379 811
rect 1375 805 1379 806
rect 1407 810 1411 811
rect 1407 805 1411 806
rect 1415 810 1419 811
rect 1415 805 1419 806
rect 1471 810 1475 811
rect 1471 805 1475 806
rect 1479 810 1483 811
rect 1479 805 1483 806
rect 1535 810 1539 811
rect 1535 805 1539 806
rect 1551 810 1555 811
rect 1551 805 1555 806
rect 1406 804 1412 805
rect 1406 800 1407 804
rect 1411 800 1412 804
rect 1406 799 1412 800
rect 1478 804 1484 805
rect 1478 800 1479 804
rect 1483 800 1484 804
rect 1478 799 1484 800
rect 1550 804 1556 805
rect 1550 800 1551 804
rect 1555 800 1556 804
rect 1550 799 1556 800
rect 1358 783 1364 784
rect 1358 779 1359 783
rect 1363 779 1364 783
rect 1358 778 1364 779
rect 1386 783 1392 784
rect 1386 779 1387 783
rect 1391 779 1392 783
rect 1386 778 1392 779
rect 1394 783 1400 784
rect 1394 779 1395 783
rect 1399 779 1400 783
rect 1394 778 1400 779
rect 1490 783 1496 784
rect 1490 779 1491 783
rect 1495 779 1496 783
rect 1490 778 1496 779
rect 1360 752 1362 778
rect 1388 752 1390 778
rect 1304 743 1306 752
rect 1318 751 1324 752
rect 1318 747 1319 751
rect 1323 747 1324 751
rect 1318 746 1324 747
rect 1279 742 1283 743
rect 1279 737 1283 738
rect 1303 742 1307 743
rect 1303 737 1307 738
rect 1106 722 1112 723
rect 1238 724 1244 725
rect 1238 720 1239 724
rect 1243 720 1244 724
rect 886 719 892 720
rect 886 715 887 719
rect 891 715 892 719
rect 886 714 892 715
rect 974 719 980 720
rect 974 715 975 719
rect 979 715 980 719
rect 974 714 980 715
rect 1086 719 1092 720
rect 1086 715 1087 719
rect 1091 715 1092 719
rect 1086 714 1092 715
rect 1174 719 1180 720
rect 1238 719 1244 720
rect 1174 715 1175 719
rect 1179 715 1180 719
rect 1174 714 1180 715
rect 782 700 788 701
rect 782 696 783 700
rect 787 696 788 700
rect 782 695 788 696
rect 878 700 884 701
rect 878 696 879 700
rect 883 696 884 700
rect 878 695 884 696
rect 982 700 988 701
rect 982 696 983 700
rect 987 696 988 700
rect 982 695 988 696
rect 1094 700 1100 701
rect 1094 696 1095 700
rect 1099 696 1100 700
rect 1094 695 1100 696
rect 784 687 786 695
rect 880 687 882 695
rect 984 687 986 695
rect 1096 687 1098 695
rect 767 686 771 687
rect 767 681 771 682
rect 783 686 787 687
rect 783 681 787 682
rect 839 686 843 687
rect 839 681 843 682
rect 879 686 883 687
rect 879 681 883 682
rect 903 686 907 687
rect 903 681 907 682
rect 967 686 971 687
rect 967 681 971 682
rect 983 686 987 687
rect 983 681 987 682
rect 1023 686 1027 687
rect 1023 681 1027 682
rect 1087 686 1091 687
rect 1087 681 1091 682
rect 1095 686 1099 687
rect 1095 681 1099 682
rect 1151 686 1155 687
rect 1151 681 1155 682
rect 766 680 772 681
rect 766 676 767 680
rect 771 676 772 680
rect 766 675 772 676
rect 838 680 844 681
rect 838 676 839 680
rect 843 676 844 680
rect 838 675 844 676
rect 902 680 908 681
rect 902 676 903 680
rect 907 676 908 680
rect 902 675 908 676
rect 966 680 972 681
rect 966 676 967 680
rect 971 676 972 680
rect 966 675 972 676
rect 1022 680 1028 681
rect 1022 676 1023 680
rect 1027 676 1028 680
rect 1022 675 1028 676
rect 1086 680 1092 681
rect 1086 676 1087 680
rect 1091 676 1092 680
rect 1086 675 1092 676
rect 1150 680 1156 681
rect 1150 676 1151 680
rect 1155 676 1156 680
rect 1150 675 1156 676
rect 494 659 500 660
rect 494 655 495 659
rect 499 655 500 659
rect 494 654 500 655
rect 514 659 520 660
rect 514 655 515 659
rect 519 655 520 659
rect 514 654 520 655
rect 638 659 644 660
rect 638 655 639 659
rect 643 655 644 659
rect 638 654 644 655
rect 758 659 764 660
rect 758 655 759 659
rect 763 655 764 659
rect 758 654 764 655
rect 914 659 920 660
rect 914 655 915 659
rect 919 655 920 659
rect 914 654 920 655
rect 478 651 484 652
rect 478 647 479 651
rect 483 647 484 651
rect 478 646 484 647
rect 454 633 460 634
rect 454 629 455 633
rect 459 629 460 633
rect 454 628 460 629
rect 480 628 482 646
rect 496 628 498 654
rect 502 633 508 634
rect 502 629 503 633
rect 507 629 508 633
rect 502 628 508 629
rect 136 619 138 628
rect 158 627 164 628
rect 158 623 159 627
rect 163 623 164 627
rect 158 622 164 623
rect 111 618 115 619
rect 111 613 115 614
rect 135 618 139 619
rect 135 613 139 614
rect 112 581 114 613
rect 136 604 138 613
rect 134 603 140 604
rect 134 599 135 603
rect 139 599 140 603
rect 134 598 140 599
rect 110 580 116 581
rect 110 576 111 580
rect 115 576 116 580
rect 160 576 162 622
rect 176 619 178 628
rect 210 627 216 628
rect 210 623 211 627
rect 215 623 216 627
rect 210 622 216 623
rect 232 619 234 628
rect 288 619 290 628
rect 310 627 316 628
rect 310 623 311 627
rect 315 623 316 627
rect 310 622 316 623
rect 344 619 346 628
rect 400 619 402 628
rect 438 627 444 628
rect 438 623 439 627
rect 443 623 444 627
rect 438 622 444 623
rect 456 619 458 628
rect 478 627 484 628
rect 478 623 479 627
rect 483 623 484 627
rect 478 622 484 623
rect 494 627 500 628
rect 494 623 495 627
rect 499 623 500 627
rect 494 622 500 623
rect 504 619 506 628
rect 175 618 179 619
rect 175 613 179 614
rect 183 618 187 619
rect 183 613 187 614
rect 231 618 235 619
rect 231 613 235 614
rect 255 618 259 619
rect 255 613 259 614
rect 287 618 291 619
rect 287 613 291 614
rect 327 618 331 619
rect 327 613 331 614
rect 343 618 347 619
rect 343 613 347 614
rect 399 618 403 619
rect 399 613 403 614
rect 455 618 459 619
rect 455 613 459 614
rect 479 618 483 619
rect 479 613 483 614
rect 503 618 507 619
rect 503 613 507 614
rect 174 607 180 608
rect 174 603 175 607
rect 179 603 180 607
rect 184 604 186 613
rect 246 607 252 608
rect 174 602 180 603
rect 182 603 188 604
rect 176 576 178 602
rect 182 599 183 603
rect 187 599 188 603
rect 246 603 247 607
rect 251 603 252 607
rect 256 604 258 613
rect 318 607 324 608
rect 246 602 252 603
rect 254 603 260 604
rect 182 598 188 599
rect 248 576 250 602
rect 254 599 255 603
rect 259 599 260 603
rect 318 603 319 607
rect 323 603 324 607
rect 328 604 330 613
rect 338 607 344 608
rect 318 602 324 603
rect 326 603 332 604
rect 254 598 260 599
rect 320 576 322 602
rect 326 599 327 603
rect 331 599 332 603
rect 338 603 339 607
rect 343 603 344 607
rect 400 604 402 613
rect 470 607 476 608
rect 338 602 344 603
rect 398 603 404 604
rect 326 598 332 599
rect 110 575 116 576
rect 158 575 164 576
rect 158 571 159 575
rect 163 571 164 575
rect 158 570 164 571
rect 174 575 180 576
rect 174 571 175 575
rect 179 571 180 575
rect 174 570 180 571
rect 246 575 252 576
rect 246 571 247 575
rect 251 571 252 575
rect 246 570 252 571
rect 318 575 324 576
rect 318 571 319 575
rect 323 571 324 575
rect 318 570 324 571
rect 110 563 116 564
rect 110 559 111 563
rect 115 559 116 563
rect 110 558 116 559
rect 112 547 114 558
rect 134 556 140 557
rect 134 552 135 556
rect 139 552 140 556
rect 134 551 140 552
rect 182 556 188 557
rect 182 552 183 556
rect 187 552 188 556
rect 182 551 188 552
rect 254 556 260 557
rect 254 552 255 556
rect 259 552 260 556
rect 254 551 260 552
rect 326 556 332 557
rect 326 552 327 556
rect 331 552 332 556
rect 326 551 332 552
rect 136 547 138 551
rect 184 547 186 551
rect 256 547 258 551
rect 328 547 330 551
rect 111 546 115 547
rect 111 541 115 542
rect 135 546 139 547
rect 135 541 139 542
rect 151 546 155 547
rect 151 541 155 542
rect 183 546 187 547
rect 183 541 187 542
rect 223 546 227 547
rect 223 541 227 542
rect 255 546 259 547
rect 255 541 259 542
rect 287 546 291 547
rect 287 541 291 542
rect 327 546 331 547
rect 327 541 331 542
rect 112 534 114 541
rect 150 540 156 541
rect 150 536 151 540
rect 155 536 156 540
rect 150 535 156 536
rect 222 540 228 541
rect 222 536 223 540
rect 227 536 228 540
rect 222 535 228 536
rect 286 540 292 541
rect 286 536 287 540
rect 291 536 292 540
rect 286 535 292 536
rect 110 533 116 534
rect 110 529 111 533
rect 115 529 116 533
rect 110 528 116 529
rect 340 520 342 602
rect 398 599 399 603
rect 403 599 404 603
rect 470 603 471 607
rect 475 603 476 607
rect 480 604 482 613
rect 516 608 518 654
rect 558 633 564 634
rect 558 629 559 633
rect 563 629 564 633
rect 558 628 564 629
rect 622 633 628 634
rect 622 629 623 633
rect 627 629 628 633
rect 622 628 628 629
rect 640 628 642 654
rect 718 651 724 652
rect 718 647 719 651
rect 723 647 724 651
rect 718 646 724 647
rect 862 651 868 652
rect 862 647 863 651
rect 867 647 868 651
rect 862 646 868 647
rect 694 633 700 634
rect 694 629 695 633
rect 699 629 700 633
rect 694 628 700 629
rect 720 628 722 646
rect 766 633 772 634
rect 766 629 767 633
rect 771 629 772 633
rect 766 628 772 629
rect 838 633 844 634
rect 838 629 839 633
rect 843 629 844 633
rect 838 628 844 629
rect 864 628 866 646
rect 902 633 908 634
rect 902 629 903 633
rect 907 629 908 633
rect 902 628 908 629
rect 560 619 562 628
rect 624 619 626 628
rect 638 627 644 628
rect 638 623 639 627
rect 643 623 644 627
rect 638 622 644 623
rect 662 627 668 628
rect 662 623 663 627
rect 667 623 668 627
rect 662 622 668 623
rect 559 618 563 619
rect 559 613 563 614
rect 623 618 627 619
rect 623 613 627 614
rect 639 618 643 619
rect 639 613 643 614
rect 514 607 520 608
rect 470 602 476 603
rect 478 603 484 604
rect 398 598 404 599
rect 472 576 474 602
rect 478 599 479 603
rect 483 599 484 603
rect 514 603 515 607
rect 519 603 520 607
rect 560 604 562 613
rect 570 607 576 608
rect 514 602 520 603
rect 558 603 564 604
rect 478 598 484 599
rect 558 599 559 603
rect 563 599 564 603
rect 570 603 571 607
rect 575 603 576 607
rect 640 604 642 613
rect 570 602 576 603
rect 638 603 644 604
rect 558 598 564 599
rect 572 584 574 602
rect 638 599 639 603
rect 643 599 644 603
rect 638 598 644 599
rect 570 583 576 584
rect 570 579 571 583
rect 575 579 576 583
rect 570 578 576 579
rect 664 576 666 622
rect 696 619 698 628
rect 718 627 724 628
rect 718 623 719 627
rect 723 623 724 627
rect 718 622 724 623
rect 768 619 770 628
rect 840 619 842 628
rect 862 627 868 628
rect 862 623 863 627
rect 867 623 868 627
rect 862 622 868 623
rect 904 619 906 628
rect 695 618 699 619
rect 695 613 699 614
rect 719 618 723 619
rect 719 613 723 614
rect 767 618 771 619
rect 767 613 771 614
rect 799 618 803 619
rect 799 613 803 614
rect 839 618 843 619
rect 839 613 843 614
rect 879 618 883 619
rect 879 613 883 614
rect 903 618 907 619
rect 903 613 907 614
rect 710 607 716 608
rect 710 603 711 607
rect 715 603 716 607
rect 720 604 722 613
rect 790 607 796 608
rect 710 602 716 603
rect 718 603 724 604
rect 712 576 714 602
rect 718 599 719 603
rect 723 599 724 603
rect 790 603 791 607
rect 795 603 796 607
rect 800 604 802 613
rect 810 607 816 608
rect 790 602 796 603
rect 798 603 804 604
rect 718 598 724 599
rect 792 576 794 602
rect 798 599 799 603
rect 803 599 804 603
rect 810 603 811 607
rect 815 603 816 607
rect 880 604 882 613
rect 916 608 918 654
rect 966 633 972 634
rect 966 629 967 633
rect 971 629 972 633
rect 966 628 972 629
rect 1022 633 1028 634
rect 1022 629 1023 633
rect 1027 629 1028 633
rect 1022 628 1028 629
rect 1086 633 1092 634
rect 1086 629 1087 633
rect 1091 629 1092 633
rect 1086 628 1092 629
rect 1150 633 1156 634
rect 1150 629 1151 633
rect 1155 629 1156 633
rect 1150 628 1156 629
rect 1176 628 1178 714
rect 1238 707 1244 708
rect 1238 703 1239 707
rect 1243 703 1244 707
rect 1280 705 1282 737
rect 1304 728 1306 737
rect 1302 727 1308 728
rect 1302 723 1303 727
rect 1307 723 1308 727
rect 1302 722 1308 723
rect 1238 702 1244 703
rect 1278 704 1284 705
rect 1190 700 1196 701
rect 1190 696 1191 700
rect 1195 696 1196 700
rect 1190 695 1196 696
rect 1192 687 1194 695
rect 1240 687 1242 702
rect 1278 700 1279 704
rect 1283 700 1284 704
rect 1320 700 1322 746
rect 1344 743 1346 752
rect 1350 751 1356 752
rect 1350 747 1351 751
rect 1355 747 1356 751
rect 1350 746 1356 747
rect 1358 751 1364 752
rect 1358 747 1359 751
rect 1363 747 1364 751
rect 1358 746 1364 747
rect 1386 751 1392 752
rect 1386 747 1387 751
rect 1391 747 1392 751
rect 1386 746 1392 747
rect 1343 742 1347 743
rect 1343 737 1347 738
rect 1367 742 1371 743
rect 1367 737 1371 738
rect 1358 731 1364 732
rect 1358 727 1359 731
rect 1363 727 1364 731
rect 1368 728 1370 737
rect 1396 732 1398 778
rect 1406 757 1412 758
rect 1406 753 1407 757
rect 1411 753 1412 757
rect 1406 752 1412 753
rect 1478 757 1484 758
rect 1478 753 1479 757
rect 1483 753 1484 757
rect 1478 752 1484 753
rect 1408 743 1410 752
rect 1480 743 1482 752
rect 1407 742 1411 743
rect 1407 737 1411 738
rect 1455 742 1459 743
rect 1455 737 1459 738
rect 1479 742 1483 743
rect 1479 737 1483 738
rect 1394 731 1400 732
rect 1358 726 1364 727
rect 1366 727 1372 728
rect 1360 700 1362 726
rect 1366 723 1367 727
rect 1371 723 1372 727
rect 1394 727 1395 731
rect 1399 727 1400 731
rect 1456 728 1458 737
rect 1492 732 1494 778
rect 1550 757 1556 758
rect 1550 753 1551 757
rect 1555 753 1556 757
rect 1550 752 1556 753
rect 1576 752 1578 834
rect 1606 820 1612 821
rect 1606 816 1607 820
rect 1611 816 1612 820
rect 1606 815 1612 816
rect 1608 811 1610 815
rect 1607 810 1611 811
rect 1607 805 1611 806
rect 1623 810 1627 811
rect 1623 805 1627 806
rect 1622 804 1628 805
rect 1622 800 1623 804
rect 1627 800 1628 804
rect 1622 799 1628 800
rect 1648 784 1650 866
rect 1678 863 1679 867
rect 1683 863 1684 867
rect 1690 867 1691 871
rect 1695 867 1696 871
rect 1752 868 1754 877
rect 1762 871 1768 872
rect 1690 866 1696 867
rect 1750 867 1756 868
rect 1678 862 1684 863
rect 1692 840 1694 866
rect 1750 863 1751 867
rect 1755 863 1756 867
rect 1762 867 1763 871
rect 1767 867 1768 871
rect 1762 866 1768 867
rect 1750 862 1756 863
rect 1764 840 1766 866
rect 1780 840 1782 894
rect 1840 883 1842 900
rect 1936 883 1938 900
rect 1986 899 1992 900
rect 1986 895 1987 899
rect 1991 895 1992 899
rect 1986 894 1992 895
rect 2024 883 2026 900
rect 2104 883 2106 900
rect 2130 899 2136 900
rect 2130 895 2131 899
rect 2135 895 2136 899
rect 2130 894 2136 895
rect 2176 883 2178 900
rect 2198 899 2204 900
rect 2198 895 2199 899
rect 2203 895 2204 899
rect 2198 894 2204 895
rect 2240 883 2242 900
rect 2254 899 2260 900
rect 2254 895 2255 899
rect 2259 895 2260 899
rect 2254 894 2260 895
rect 2312 883 2314 900
rect 2326 899 2332 900
rect 2326 895 2327 899
rect 2331 895 2332 899
rect 2326 894 2332 895
rect 2360 883 2362 900
rect 2374 899 2380 900
rect 2374 895 2375 899
rect 2379 895 2380 899
rect 2374 894 2380 895
rect 1823 882 1827 883
rect 1823 877 1827 878
rect 1839 882 1843 883
rect 1839 877 1843 878
rect 1895 882 1899 883
rect 1895 877 1899 878
rect 1935 882 1939 883
rect 1935 877 1939 878
rect 1959 882 1963 883
rect 1959 877 1963 878
rect 2023 882 2027 883
rect 2023 877 2027 878
rect 2087 882 2091 883
rect 2087 877 2091 878
rect 2103 882 2107 883
rect 2103 877 2107 878
rect 2143 882 2147 883
rect 2143 877 2147 878
rect 2175 882 2179 883
rect 2175 877 2179 878
rect 2199 882 2203 883
rect 2199 877 2203 878
rect 2239 882 2243 883
rect 2239 877 2243 878
rect 2255 882 2259 883
rect 2255 877 2259 878
rect 2311 882 2315 883
rect 2311 877 2315 878
rect 2319 882 2323 883
rect 2319 877 2323 878
rect 2359 882 2363 883
rect 2359 877 2363 878
rect 1824 868 1826 877
rect 1886 871 1892 872
rect 1822 867 1828 868
rect 1822 863 1823 867
rect 1827 863 1828 867
rect 1886 867 1887 871
rect 1891 867 1892 871
rect 1896 868 1898 877
rect 1950 871 1956 872
rect 1886 866 1892 867
rect 1894 867 1900 868
rect 1822 862 1828 863
rect 1888 848 1890 866
rect 1894 863 1895 867
rect 1899 863 1900 867
rect 1950 867 1951 871
rect 1955 867 1956 871
rect 1960 868 1962 877
rect 2014 871 2020 872
rect 1950 866 1956 867
rect 1958 867 1964 868
rect 1894 862 1900 863
rect 1886 847 1892 848
rect 1886 843 1887 847
rect 1891 843 1892 847
rect 1886 842 1892 843
rect 1952 840 1954 866
rect 1958 863 1959 867
rect 1963 863 1964 867
rect 2014 867 2015 871
rect 2019 867 2020 871
rect 2024 868 2026 877
rect 2078 871 2084 872
rect 2014 866 2020 867
rect 2022 867 2028 868
rect 1958 862 1964 863
rect 2016 840 2018 866
rect 2022 863 2023 867
rect 2027 863 2028 867
rect 2078 867 2079 871
rect 2083 867 2084 871
rect 2088 868 2090 877
rect 2134 871 2140 872
rect 2078 866 2084 867
rect 2086 867 2092 868
rect 2022 862 2028 863
rect 2080 840 2082 866
rect 2086 863 2087 867
rect 2091 863 2092 867
rect 2134 867 2135 871
rect 2139 867 2140 871
rect 2144 868 2146 877
rect 2200 868 2202 877
rect 2246 871 2252 872
rect 2134 866 2140 867
rect 2142 867 2148 868
rect 2086 862 2092 863
rect 2136 840 2138 866
rect 2142 863 2143 867
rect 2147 863 2148 867
rect 2142 862 2148 863
rect 2198 867 2204 868
rect 2198 863 2199 867
rect 2203 863 2204 867
rect 2246 867 2247 871
rect 2251 867 2252 871
rect 2256 868 2258 877
rect 2310 871 2316 872
rect 2246 866 2252 867
rect 2254 867 2260 868
rect 2198 862 2204 863
rect 2248 840 2250 866
rect 2254 863 2255 867
rect 2259 863 2260 867
rect 2310 867 2311 871
rect 2315 867 2316 871
rect 2320 868 2322 877
rect 2346 871 2352 872
rect 2310 866 2316 867
rect 2318 867 2324 868
rect 2254 862 2260 863
rect 2312 840 2314 866
rect 2318 863 2319 867
rect 2323 863 2324 867
rect 2346 867 2347 871
rect 2351 867 2352 871
rect 2360 868 2362 877
rect 2384 872 2386 926
rect 2406 924 2407 928
rect 2411 924 2412 928
rect 2406 923 2412 924
rect 2408 883 2410 923
rect 2407 882 2411 883
rect 2407 877 2411 878
rect 2382 871 2388 872
rect 2346 866 2352 867
rect 2358 867 2364 868
rect 2318 862 2324 863
rect 2348 848 2350 866
rect 2358 863 2359 867
rect 2363 863 2364 867
rect 2382 867 2383 871
rect 2387 867 2388 871
rect 2382 866 2388 867
rect 2358 862 2364 863
rect 2346 847 2352 848
rect 2346 843 2347 847
rect 2351 843 2352 847
rect 2408 845 2410 877
rect 2346 842 2352 843
rect 2406 844 2412 845
rect 2406 840 2407 844
rect 2411 840 2412 844
rect 1690 839 1696 840
rect 1690 835 1691 839
rect 1695 835 1696 839
rect 1690 834 1696 835
rect 1762 839 1768 840
rect 1762 835 1763 839
rect 1767 835 1768 839
rect 1762 834 1768 835
rect 1778 839 1784 840
rect 1778 835 1779 839
rect 1783 835 1784 839
rect 1778 834 1784 835
rect 1950 839 1956 840
rect 1950 835 1951 839
rect 1955 835 1956 839
rect 1950 834 1956 835
rect 2014 839 2020 840
rect 2014 835 2015 839
rect 2019 835 2020 839
rect 2014 834 2020 835
rect 2078 839 2084 840
rect 2078 835 2079 839
rect 2083 835 2084 839
rect 2078 834 2084 835
rect 2134 839 2140 840
rect 2134 835 2135 839
rect 2139 835 2140 839
rect 2134 834 2140 835
rect 2246 839 2252 840
rect 2246 835 2247 839
rect 2251 835 2252 839
rect 2246 834 2252 835
rect 2310 839 2316 840
rect 2406 839 2412 840
rect 2310 835 2311 839
rect 2315 835 2316 839
rect 2310 834 2316 835
rect 2046 831 2052 832
rect 2046 827 2047 831
rect 2051 827 2052 831
rect 2046 826 2052 827
rect 2382 831 2388 832
rect 2382 827 2383 831
rect 2387 827 2388 831
rect 2382 826 2388 827
rect 2406 827 2412 828
rect 1678 820 1684 821
rect 1678 816 1679 820
rect 1683 816 1684 820
rect 1678 815 1684 816
rect 1750 820 1756 821
rect 1750 816 1751 820
rect 1755 816 1756 820
rect 1750 815 1756 816
rect 1822 820 1828 821
rect 1822 816 1823 820
rect 1827 816 1828 820
rect 1822 815 1828 816
rect 1894 820 1900 821
rect 1894 816 1895 820
rect 1899 816 1900 820
rect 1894 815 1900 816
rect 1958 820 1964 821
rect 1958 816 1959 820
rect 1963 816 1964 820
rect 1958 815 1964 816
rect 2022 820 2028 821
rect 2022 816 2023 820
rect 2027 816 2028 820
rect 2022 815 2028 816
rect 1680 811 1682 815
rect 1752 811 1754 815
rect 1824 811 1826 815
rect 1896 811 1898 815
rect 1960 811 1962 815
rect 2024 811 2026 815
rect 1679 810 1683 811
rect 1679 805 1683 806
rect 1695 810 1699 811
rect 1695 805 1699 806
rect 1751 810 1755 811
rect 1751 805 1755 806
rect 1759 810 1763 811
rect 1759 805 1763 806
rect 1823 810 1827 811
rect 1823 805 1827 806
rect 1887 810 1891 811
rect 1887 805 1891 806
rect 1895 810 1899 811
rect 1895 805 1899 806
rect 1951 810 1955 811
rect 1951 805 1955 806
rect 1959 810 1963 811
rect 1959 805 1963 806
rect 2023 810 2027 811
rect 2023 805 2027 806
rect 1694 804 1700 805
rect 1694 800 1695 804
rect 1699 800 1700 804
rect 1694 799 1700 800
rect 1758 804 1764 805
rect 1758 800 1759 804
rect 1763 800 1764 804
rect 1758 799 1764 800
rect 1822 804 1828 805
rect 1822 800 1823 804
rect 1827 800 1828 804
rect 1822 799 1828 800
rect 1886 804 1892 805
rect 1886 800 1887 804
rect 1891 800 1892 804
rect 1886 799 1892 800
rect 1950 804 1956 805
rect 1950 800 1951 804
rect 1955 800 1956 804
rect 1950 799 1956 800
rect 2022 804 2028 805
rect 2022 800 2023 804
rect 2027 800 2028 804
rect 2022 799 2028 800
rect 1646 783 1652 784
rect 1646 779 1647 783
rect 1651 779 1652 783
rect 1646 778 1652 779
rect 1798 783 1804 784
rect 1798 779 1799 783
rect 1803 779 1804 783
rect 1798 778 1804 779
rect 1622 757 1628 758
rect 1622 753 1623 757
rect 1627 753 1628 757
rect 1622 752 1628 753
rect 1694 757 1700 758
rect 1694 753 1695 757
rect 1699 753 1700 757
rect 1694 752 1700 753
rect 1758 757 1764 758
rect 1758 753 1759 757
rect 1763 753 1764 757
rect 1758 752 1764 753
rect 1552 743 1554 752
rect 1574 751 1580 752
rect 1574 747 1575 751
rect 1579 747 1580 751
rect 1574 746 1580 747
rect 1624 743 1626 752
rect 1696 743 1698 752
rect 1718 751 1724 752
rect 1718 747 1719 751
rect 1723 747 1724 751
rect 1718 746 1724 747
rect 1535 742 1539 743
rect 1535 737 1539 738
rect 1551 742 1555 743
rect 1551 737 1555 738
rect 1615 742 1619 743
rect 1615 737 1619 738
rect 1623 742 1627 743
rect 1623 737 1627 738
rect 1695 742 1699 743
rect 1695 737 1699 738
rect 1490 731 1496 732
rect 1394 726 1400 727
rect 1454 727 1460 728
rect 1366 722 1372 723
rect 1454 723 1455 727
rect 1459 723 1460 727
rect 1490 727 1491 731
rect 1495 727 1496 731
rect 1536 728 1538 737
rect 1546 731 1552 732
rect 1490 726 1496 727
rect 1534 727 1540 728
rect 1454 722 1460 723
rect 1534 723 1535 727
rect 1539 723 1540 727
rect 1546 727 1547 731
rect 1551 727 1552 731
rect 1616 728 1618 737
rect 1662 731 1668 732
rect 1546 726 1552 727
rect 1614 727 1620 728
rect 1534 722 1540 723
rect 1548 700 1550 726
rect 1614 723 1615 727
rect 1619 723 1620 727
rect 1662 727 1663 731
rect 1667 727 1668 731
rect 1696 728 1698 737
rect 1706 731 1712 732
rect 1662 726 1668 727
rect 1694 727 1700 728
rect 1614 722 1620 723
rect 1278 699 1284 700
rect 1318 699 1324 700
rect 1318 695 1319 699
rect 1323 695 1324 699
rect 1318 694 1324 695
rect 1358 699 1364 700
rect 1358 695 1359 699
rect 1363 695 1364 699
rect 1358 694 1364 695
rect 1546 699 1552 700
rect 1546 695 1547 699
rect 1551 695 1552 699
rect 1546 694 1552 695
rect 1606 699 1612 700
rect 1606 695 1607 699
rect 1611 695 1612 699
rect 1606 694 1612 695
rect 1278 687 1284 688
rect 1191 686 1195 687
rect 1191 681 1195 682
rect 1239 686 1243 687
rect 1278 683 1279 687
rect 1283 683 1284 687
rect 1278 682 1284 683
rect 1239 681 1243 682
rect 1190 680 1196 681
rect 1190 676 1191 680
rect 1195 676 1196 680
rect 1190 675 1196 676
rect 1240 674 1242 681
rect 1280 675 1282 682
rect 1302 680 1308 681
rect 1302 676 1303 680
rect 1307 676 1308 680
rect 1302 675 1308 676
rect 1366 680 1372 681
rect 1366 676 1367 680
rect 1371 676 1372 680
rect 1366 675 1372 676
rect 1454 680 1460 681
rect 1454 676 1455 680
rect 1459 676 1460 680
rect 1454 675 1460 676
rect 1534 680 1540 681
rect 1534 676 1535 680
rect 1539 676 1540 680
rect 1534 675 1540 676
rect 1279 674 1283 675
rect 1238 673 1244 674
rect 1238 669 1239 673
rect 1243 669 1244 673
rect 1279 669 1283 670
rect 1303 674 1307 675
rect 1303 669 1307 670
rect 1367 674 1371 675
rect 1367 669 1371 670
rect 1455 674 1459 675
rect 1455 669 1459 670
rect 1535 674 1539 675
rect 1535 669 1539 670
rect 1591 674 1595 675
rect 1591 669 1595 670
rect 1238 668 1244 669
rect 1280 662 1282 669
rect 1590 668 1596 669
rect 1590 664 1591 668
rect 1595 664 1596 668
rect 1590 663 1596 664
rect 1278 661 1284 662
rect 1214 659 1220 660
rect 1214 655 1215 659
rect 1219 655 1220 659
rect 1278 657 1279 661
rect 1283 657 1284 661
rect 1214 654 1220 655
rect 1238 656 1244 657
rect 1278 656 1284 657
rect 1198 651 1204 652
rect 1198 647 1199 651
rect 1203 647 1204 651
rect 1198 646 1204 647
rect 1190 633 1196 634
rect 1190 629 1191 633
rect 1195 629 1196 633
rect 1190 628 1196 629
rect 1200 628 1202 646
rect 968 619 970 628
rect 1024 619 1026 628
rect 1088 619 1090 628
rect 1102 627 1108 628
rect 1102 623 1103 627
rect 1107 623 1108 627
rect 1102 622 1108 623
rect 951 618 955 619
rect 951 613 955 614
rect 967 618 971 619
rect 967 613 971 614
rect 1015 618 1019 619
rect 1015 613 1019 614
rect 1023 618 1027 619
rect 1023 613 1027 614
rect 1079 618 1083 619
rect 1079 613 1083 614
rect 1087 618 1091 619
rect 1087 613 1091 614
rect 914 607 920 608
rect 810 602 816 603
rect 878 603 884 604
rect 798 598 804 599
rect 470 575 476 576
rect 470 571 471 575
rect 475 571 476 575
rect 470 570 476 571
rect 578 575 584 576
rect 578 571 579 575
rect 583 571 584 575
rect 578 570 584 571
rect 662 575 668 576
rect 662 571 663 575
rect 667 571 668 575
rect 662 570 668 571
rect 710 575 716 576
rect 710 571 711 575
rect 715 571 716 575
rect 710 570 716 571
rect 790 575 796 576
rect 790 571 791 575
rect 795 571 796 575
rect 790 570 796 571
rect 398 556 404 557
rect 398 552 399 556
rect 403 552 404 556
rect 398 551 404 552
rect 478 556 484 557
rect 478 552 479 556
rect 483 552 484 556
rect 478 551 484 552
rect 558 556 564 557
rect 558 552 559 556
rect 563 552 564 556
rect 558 551 564 552
rect 400 547 402 551
rect 480 547 482 551
rect 560 547 562 551
rect 351 546 355 547
rect 351 541 355 542
rect 399 546 403 547
rect 399 541 403 542
rect 415 546 419 547
rect 415 541 419 542
rect 479 546 483 547
rect 479 541 483 542
rect 551 546 555 547
rect 551 541 555 542
rect 559 546 563 547
rect 559 541 563 542
rect 350 540 356 541
rect 350 536 351 540
rect 355 536 356 540
rect 350 535 356 536
rect 414 540 420 541
rect 414 536 415 540
rect 419 536 420 540
rect 414 535 420 536
rect 478 540 484 541
rect 478 536 479 540
rect 483 536 484 540
rect 478 535 484 536
rect 550 540 556 541
rect 550 536 551 540
rect 555 536 556 540
rect 550 535 556 536
rect 338 519 344 520
rect 110 516 116 517
rect 110 512 111 516
rect 115 512 116 516
rect 338 515 339 519
rect 343 515 344 519
rect 338 514 344 515
rect 110 511 116 512
rect 310 511 316 512
rect 112 479 114 511
rect 310 507 311 511
rect 315 507 316 511
rect 310 506 316 507
rect 462 511 468 512
rect 462 507 463 511
rect 467 507 468 511
rect 462 506 468 507
rect 150 493 156 494
rect 150 489 151 493
rect 155 489 156 493
rect 150 488 156 489
rect 222 493 228 494
rect 222 489 223 493
rect 227 489 228 493
rect 222 488 228 489
rect 286 493 292 494
rect 286 489 287 493
rect 291 489 292 493
rect 286 488 292 489
rect 312 488 314 506
rect 350 493 356 494
rect 350 489 351 493
rect 355 489 356 493
rect 350 488 356 489
rect 414 493 420 494
rect 414 489 415 493
rect 419 489 420 493
rect 414 488 420 489
rect 152 479 154 488
rect 224 479 226 488
rect 262 487 268 488
rect 262 483 263 487
rect 267 483 268 487
rect 262 482 268 483
rect 111 478 115 479
rect 111 473 115 474
rect 151 478 155 479
rect 151 473 155 474
rect 223 478 227 479
rect 223 473 227 474
rect 239 478 243 479
rect 239 473 243 474
rect 112 441 114 473
rect 240 464 242 473
rect 238 463 244 464
rect 238 459 239 463
rect 243 459 244 463
rect 238 458 244 459
rect 110 440 116 441
rect 110 436 111 440
rect 115 436 116 440
rect 264 436 266 482
rect 288 479 290 488
rect 310 487 316 488
rect 310 483 311 487
rect 315 483 316 487
rect 310 482 316 483
rect 352 479 354 488
rect 416 479 418 488
rect 279 478 283 479
rect 279 473 283 474
rect 287 478 291 479
rect 287 473 291 474
rect 327 478 331 479
rect 327 473 331 474
rect 351 478 355 479
rect 351 473 355 474
rect 383 478 387 479
rect 383 473 387 474
rect 415 478 419 479
rect 415 473 419 474
rect 439 478 443 479
rect 439 473 443 474
rect 280 464 282 473
rect 294 471 300 472
rect 294 467 295 471
rect 299 467 300 471
rect 294 466 300 467
rect 318 467 324 468
rect 278 463 284 464
rect 278 459 279 463
rect 283 459 284 463
rect 278 458 284 459
rect 296 436 298 466
rect 318 463 319 467
rect 323 463 324 467
rect 328 464 330 473
rect 374 467 380 468
rect 318 462 324 463
rect 326 463 332 464
rect 320 436 322 462
rect 326 459 327 463
rect 331 459 332 463
rect 374 463 375 467
rect 379 463 380 467
rect 384 464 386 473
rect 406 467 412 468
rect 374 462 380 463
rect 382 463 388 464
rect 326 458 332 459
rect 376 436 378 462
rect 382 459 383 463
rect 387 459 388 463
rect 406 463 407 467
rect 411 463 412 467
rect 440 464 442 473
rect 464 468 466 506
rect 478 493 484 494
rect 478 489 479 493
rect 483 489 484 493
rect 478 488 484 489
rect 550 493 556 494
rect 550 489 551 493
rect 555 489 556 493
rect 550 488 556 489
rect 580 488 582 570
rect 638 556 644 557
rect 638 552 639 556
rect 643 552 644 556
rect 638 551 644 552
rect 718 556 724 557
rect 718 552 719 556
rect 723 552 724 556
rect 718 551 724 552
rect 798 556 804 557
rect 798 552 799 556
rect 803 552 804 556
rect 798 551 804 552
rect 640 547 642 551
rect 720 547 722 551
rect 800 547 802 551
rect 623 546 627 547
rect 623 541 627 542
rect 639 546 643 547
rect 639 541 643 542
rect 695 546 699 547
rect 695 541 699 542
rect 719 546 723 547
rect 719 541 723 542
rect 767 546 771 547
rect 767 541 771 542
rect 799 546 803 547
rect 799 541 803 542
rect 622 540 628 541
rect 622 536 623 540
rect 627 536 628 540
rect 622 535 628 536
rect 694 540 700 541
rect 694 536 695 540
rect 699 536 700 540
rect 694 535 700 536
rect 766 540 772 541
rect 766 536 767 540
rect 771 536 772 540
rect 766 535 772 536
rect 812 528 814 602
rect 878 599 879 603
rect 883 599 884 603
rect 914 603 915 607
rect 919 603 920 607
rect 952 604 954 613
rect 962 607 968 608
rect 914 602 920 603
rect 950 603 956 604
rect 878 598 884 599
rect 950 599 951 603
rect 955 599 956 603
rect 962 603 963 607
rect 967 603 968 607
rect 1016 604 1018 613
rect 1026 607 1032 608
rect 962 602 968 603
rect 1014 603 1020 604
rect 950 598 956 599
rect 964 576 966 602
rect 1014 599 1015 603
rect 1019 599 1020 603
rect 1026 603 1027 607
rect 1031 603 1032 607
rect 1080 604 1082 613
rect 1026 602 1032 603
rect 1078 603 1084 604
rect 1014 598 1020 599
rect 1028 576 1030 602
rect 1078 599 1079 603
rect 1083 599 1084 603
rect 1078 598 1084 599
rect 1104 576 1106 622
rect 1152 619 1154 628
rect 1174 627 1180 628
rect 1174 623 1175 627
rect 1179 623 1180 627
rect 1174 622 1180 623
rect 1192 619 1194 628
rect 1198 627 1204 628
rect 1198 623 1199 627
rect 1203 623 1204 627
rect 1198 622 1204 623
rect 1143 618 1147 619
rect 1143 613 1147 614
rect 1151 618 1155 619
rect 1151 613 1155 614
rect 1191 618 1195 619
rect 1191 613 1195 614
rect 1134 607 1140 608
rect 1134 603 1135 607
rect 1139 603 1140 607
rect 1144 604 1146 613
rect 1182 607 1188 608
rect 1134 602 1140 603
rect 1142 603 1148 604
rect 1136 576 1138 602
rect 1142 599 1143 603
rect 1147 599 1148 603
rect 1182 603 1183 607
rect 1187 603 1188 607
rect 1192 604 1194 613
rect 1216 608 1218 654
rect 1238 652 1239 656
rect 1243 652 1244 656
rect 1238 651 1244 652
rect 1240 619 1242 651
rect 1582 647 1588 648
rect 1278 644 1284 645
rect 1278 640 1279 644
rect 1283 640 1284 644
rect 1582 643 1583 647
rect 1587 643 1588 647
rect 1582 642 1588 643
rect 1278 639 1284 640
rect 1239 618 1243 619
rect 1239 613 1243 614
rect 1214 607 1220 608
rect 1182 602 1188 603
rect 1190 603 1196 604
rect 1142 598 1148 599
rect 1184 576 1186 602
rect 1190 599 1191 603
rect 1195 599 1196 603
rect 1214 603 1215 607
rect 1219 603 1220 607
rect 1214 602 1220 603
rect 1190 598 1196 599
rect 1240 581 1242 613
rect 1280 599 1282 639
rect 1279 598 1283 599
rect 1279 593 1283 594
rect 1559 598 1563 599
rect 1559 593 1563 594
rect 1238 580 1244 581
rect 1238 576 1239 580
rect 1243 576 1244 580
rect 962 575 968 576
rect 962 571 963 575
rect 967 571 968 575
rect 962 570 968 571
rect 1026 575 1032 576
rect 1026 571 1027 575
rect 1031 571 1032 575
rect 1026 570 1032 571
rect 1094 575 1100 576
rect 1094 571 1095 575
rect 1099 571 1100 575
rect 1094 570 1100 571
rect 1102 575 1108 576
rect 1102 571 1103 575
rect 1107 571 1108 575
rect 1102 570 1108 571
rect 1134 575 1140 576
rect 1134 571 1135 575
rect 1139 571 1140 575
rect 1134 570 1140 571
rect 1182 575 1188 576
rect 1238 575 1244 576
rect 1182 571 1183 575
rect 1187 571 1188 575
rect 1182 570 1188 571
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 950 556 956 557
rect 950 552 951 556
rect 955 552 956 556
rect 950 551 956 552
rect 1014 556 1020 557
rect 1014 552 1015 556
rect 1019 552 1020 556
rect 1014 551 1020 552
rect 1078 556 1084 557
rect 1078 552 1079 556
rect 1083 552 1084 556
rect 1078 551 1084 552
rect 880 547 882 551
rect 952 547 954 551
rect 1016 547 1018 551
rect 1080 547 1082 551
rect 839 546 843 547
rect 839 541 843 542
rect 879 546 883 547
rect 879 541 883 542
rect 919 546 923 547
rect 919 541 923 542
rect 951 546 955 547
rect 951 541 955 542
rect 999 546 1003 547
rect 999 541 1003 542
rect 1015 546 1019 547
rect 1015 541 1019 542
rect 1079 546 1083 547
rect 1079 541 1083 542
rect 838 540 844 541
rect 838 536 839 540
rect 843 536 844 540
rect 838 535 844 536
rect 918 540 924 541
rect 918 536 919 540
rect 923 536 924 540
rect 918 535 924 536
rect 998 540 1004 541
rect 998 536 999 540
rect 1003 536 1004 540
rect 998 535 1004 536
rect 1078 540 1084 541
rect 1078 536 1079 540
rect 1083 536 1084 540
rect 1078 535 1084 536
rect 810 527 816 528
rect 810 523 811 527
rect 815 523 816 527
rect 810 522 816 523
rect 830 519 836 520
rect 670 515 676 516
rect 670 511 671 515
rect 675 511 676 515
rect 830 515 831 519
rect 835 515 836 519
rect 830 514 836 515
rect 974 519 980 520
rect 974 515 975 519
rect 979 515 980 519
rect 974 514 980 515
rect 982 519 988 520
rect 982 515 983 519
rect 987 515 988 519
rect 982 514 988 515
rect 670 510 676 511
rect 622 493 628 494
rect 622 489 623 493
rect 627 489 628 493
rect 622 488 628 489
rect 672 488 674 510
rect 832 496 834 514
rect 830 495 836 496
rect 694 493 700 494
rect 694 489 695 493
rect 699 489 700 493
rect 694 488 700 489
rect 766 493 772 494
rect 766 489 767 493
rect 771 489 772 493
rect 830 491 831 495
rect 835 491 836 495
rect 830 490 836 491
rect 838 493 844 494
rect 766 488 772 489
rect 838 489 839 493
rect 843 489 844 493
rect 838 488 844 489
rect 918 493 924 494
rect 918 489 919 493
rect 923 489 924 493
rect 918 488 924 489
rect 480 479 482 488
rect 552 479 554 488
rect 578 487 584 488
rect 578 483 579 487
rect 583 483 584 487
rect 578 482 584 483
rect 624 479 626 488
rect 670 487 676 488
rect 670 483 671 487
rect 675 483 676 487
rect 670 482 676 483
rect 658 479 664 480
rect 696 479 698 488
rect 768 479 770 488
rect 840 479 842 488
rect 920 479 922 488
rect 479 478 483 479
rect 479 473 483 474
rect 503 478 507 479
rect 503 473 507 474
rect 551 478 555 479
rect 551 473 555 474
rect 567 478 571 479
rect 567 473 571 474
rect 623 478 627 479
rect 623 473 627 474
rect 631 478 635 479
rect 658 475 659 479
rect 663 475 664 479
rect 658 474 664 475
rect 695 478 699 479
rect 631 473 635 474
rect 462 467 468 468
rect 406 462 412 463
rect 438 463 444 464
rect 382 458 388 459
rect 110 435 116 436
rect 262 435 268 436
rect 262 431 263 435
rect 267 431 268 435
rect 262 430 268 431
rect 294 435 300 436
rect 294 431 295 435
rect 299 431 300 435
rect 294 430 300 431
rect 318 435 324 436
rect 318 431 319 435
rect 323 431 324 435
rect 318 430 324 431
rect 374 435 380 436
rect 374 431 375 435
rect 379 431 380 435
rect 374 430 380 431
rect 110 423 116 424
rect 110 419 111 423
rect 115 419 116 423
rect 110 418 116 419
rect 112 407 114 418
rect 238 416 244 417
rect 238 412 239 416
rect 243 412 244 416
rect 238 411 244 412
rect 278 416 284 417
rect 278 412 279 416
rect 283 412 284 416
rect 278 411 284 412
rect 326 416 332 417
rect 326 412 327 416
rect 331 412 332 416
rect 326 411 332 412
rect 382 416 388 417
rect 382 412 383 416
rect 387 412 388 416
rect 382 411 388 412
rect 240 407 242 411
rect 280 407 282 411
rect 328 407 330 411
rect 384 407 386 411
rect 111 406 115 407
rect 111 401 115 402
rect 143 406 147 407
rect 143 401 147 402
rect 183 406 187 407
rect 183 401 187 402
rect 223 406 227 407
rect 223 401 227 402
rect 239 406 243 407
rect 239 401 243 402
rect 271 406 275 407
rect 271 401 275 402
rect 279 406 283 407
rect 279 401 283 402
rect 327 406 331 407
rect 327 401 331 402
rect 335 406 339 407
rect 335 401 339 402
rect 383 406 387 407
rect 383 401 387 402
rect 399 406 403 407
rect 399 401 403 402
rect 112 394 114 401
rect 142 400 148 401
rect 142 396 143 400
rect 147 396 148 400
rect 142 395 148 396
rect 182 400 188 401
rect 182 396 183 400
rect 187 396 188 400
rect 182 395 188 396
rect 222 400 228 401
rect 222 396 223 400
rect 227 396 228 400
rect 222 395 228 396
rect 270 400 276 401
rect 270 396 271 400
rect 275 396 276 400
rect 270 395 276 396
rect 334 400 340 401
rect 334 396 335 400
rect 339 396 340 400
rect 334 395 340 396
rect 398 400 404 401
rect 398 396 399 400
rect 403 396 404 400
rect 398 395 404 396
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 110 388 116 389
rect 408 388 410 462
rect 438 459 439 463
rect 443 459 444 463
rect 462 463 463 467
rect 467 463 468 467
rect 504 464 506 473
rect 514 467 520 468
rect 462 462 468 463
rect 502 463 508 464
rect 438 458 444 459
rect 502 459 503 463
rect 507 459 508 463
rect 514 463 515 467
rect 519 463 520 467
rect 568 464 570 473
rect 578 467 584 468
rect 578 466 579 467
rect 514 462 520 463
rect 566 463 572 464
rect 502 458 508 459
rect 516 436 518 462
rect 566 459 567 463
rect 571 459 572 463
rect 566 458 572 459
rect 576 463 579 466
rect 583 463 584 467
rect 632 464 634 473
rect 576 462 584 463
rect 630 463 636 464
rect 576 436 578 462
rect 630 459 631 463
rect 635 459 636 463
rect 630 458 636 459
rect 660 436 662 474
rect 695 473 699 474
rect 759 478 763 479
rect 759 473 763 474
rect 767 478 771 479
rect 767 473 771 474
rect 823 478 827 479
rect 823 473 827 474
rect 839 478 843 479
rect 839 473 843 474
rect 887 478 891 479
rect 887 473 891 474
rect 919 478 923 479
rect 919 473 923 474
rect 951 478 955 479
rect 951 473 955 474
rect 686 467 692 468
rect 686 463 687 467
rect 691 463 692 467
rect 696 464 698 473
rect 750 467 756 468
rect 686 462 692 463
rect 694 463 700 464
rect 688 436 690 462
rect 694 459 695 463
rect 699 459 700 463
rect 750 463 751 467
rect 755 463 756 467
rect 760 464 762 473
rect 814 467 820 468
rect 750 462 756 463
rect 758 463 764 464
rect 694 458 700 459
rect 752 436 754 462
rect 758 459 759 463
rect 763 459 764 463
rect 814 463 815 467
rect 819 463 820 467
rect 824 464 826 473
rect 878 467 884 468
rect 814 462 820 463
rect 822 463 828 464
rect 758 458 764 459
rect 816 436 818 462
rect 822 459 823 463
rect 827 459 828 463
rect 878 463 879 467
rect 883 463 884 467
rect 888 464 890 473
rect 898 467 904 468
rect 878 462 884 463
rect 886 463 892 464
rect 822 458 828 459
rect 880 436 882 462
rect 886 459 887 463
rect 891 459 892 463
rect 898 463 899 467
rect 903 463 904 467
rect 952 464 954 473
rect 976 468 978 514
rect 984 488 986 514
rect 998 493 1004 494
rect 998 489 999 493
rect 1003 489 1004 493
rect 998 488 1004 489
rect 1078 493 1084 494
rect 1078 489 1079 493
rect 1083 489 1084 493
rect 1078 488 1084 489
rect 1096 488 1098 570
rect 1238 563 1244 564
rect 1238 559 1239 563
rect 1243 559 1244 563
rect 1280 561 1282 593
rect 1560 584 1562 593
rect 1584 588 1586 642
rect 1590 621 1596 622
rect 1590 617 1591 621
rect 1595 617 1596 621
rect 1590 616 1596 617
rect 1608 616 1610 694
rect 1614 680 1620 681
rect 1614 676 1615 680
rect 1619 676 1620 680
rect 1614 675 1620 676
rect 1615 674 1619 675
rect 1615 669 1619 670
rect 1639 674 1643 675
rect 1639 669 1643 670
rect 1638 668 1644 669
rect 1638 664 1639 668
rect 1643 664 1644 668
rect 1638 663 1644 664
rect 1664 648 1666 726
rect 1694 723 1695 727
rect 1699 723 1700 727
rect 1706 727 1707 731
rect 1711 727 1712 731
rect 1706 726 1712 727
rect 1694 722 1700 723
rect 1708 700 1710 726
rect 1720 700 1722 746
rect 1760 743 1762 752
rect 1759 742 1763 743
rect 1759 737 1763 738
rect 1775 742 1779 743
rect 1775 737 1779 738
rect 1776 728 1778 737
rect 1800 732 1802 778
rect 1822 757 1828 758
rect 1822 753 1823 757
rect 1827 753 1828 757
rect 1822 752 1828 753
rect 1886 757 1892 758
rect 1886 753 1887 757
rect 1891 753 1892 757
rect 1886 752 1892 753
rect 1950 757 1956 758
rect 1950 753 1951 757
rect 1955 753 1956 757
rect 1950 752 1956 753
rect 2022 757 2028 758
rect 2022 753 2023 757
rect 2027 753 2028 757
rect 2022 752 2028 753
rect 2048 752 2050 826
rect 2086 820 2092 821
rect 2086 816 2087 820
rect 2091 816 2092 820
rect 2086 815 2092 816
rect 2142 820 2148 821
rect 2142 816 2143 820
rect 2147 816 2148 820
rect 2142 815 2148 816
rect 2198 820 2204 821
rect 2198 816 2199 820
rect 2203 816 2204 820
rect 2198 815 2204 816
rect 2254 820 2260 821
rect 2254 816 2255 820
rect 2259 816 2260 820
rect 2254 815 2260 816
rect 2318 820 2324 821
rect 2318 816 2319 820
rect 2323 816 2324 820
rect 2318 815 2324 816
rect 2358 820 2364 821
rect 2358 816 2359 820
rect 2363 816 2364 820
rect 2358 815 2364 816
rect 2088 811 2090 815
rect 2144 811 2146 815
rect 2200 811 2202 815
rect 2256 811 2258 815
rect 2320 811 2322 815
rect 2360 811 2362 815
rect 2087 810 2091 811
rect 2087 805 2091 806
rect 2103 810 2107 811
rect 2103 805 2107 806
rect 2143 810 2147 811
rect 2143 805 2147 806
rect 2191 810 2195 811
rect 2191 805 2195 806
rect 2199 810 2203 811
rect 2199 805 2203 806
rect 2255 810 2259 811
rect 2255 805 2259 806
rect 2279 810 2283 811
rect 2279 805 2283 806
rect 2319 810 2323 811
rect 2319 805 2323 806
rect 2359 810 2363 811
rect 2359 805 2363 806
rect 2102 804 2108 805
rect 2102 800 2103 804
rect 2107 800 2108 804
rect 2102 799 2108 800
rect 2190 804 2196 805
rect 2190 800 2191 804
rect 2195 800 2196 804
rect 2190 799 2196 800
rect 2278 804 2284 805
rect 2278 800 2279 804
rect 2283 800 2284 804
rect 2278 799 2284 800
rect 2358 804 2364 805
rect 2358 800 2359 804
rect 2363 800 2364 804
rect 2358 799 2364 800
rect 2322 783 2328 784
rect 2322 779 2323 783
rect 2327 779 2328 783
rect 2322 778 2328 779
rect 2302 775 2308 776
rect 2302 771 2303 775
rect 2307 771 2308 775
rect 2302 770 2308 771
rect 2102 757 2108 758
rect 2102 753 2103 757
rect 2107 753 2108 757
rect 2102 752 2108 753
rect 2190 757 2196 758
rect 2190 753 2191 757
rect 2195 753 2196 757
rect 2190 752 2196 753
rect 2278 757 2284 758
rect 2278 753 2279 757
rect 2283 753 2284 757
rect 2278 752 2284 753
rect 2304 752 2306 770
rect 1824 743 1826 752
rect 1888 743 1890 752
rect 1952 743 1954 752
rect 2024 743 2026 752
rect 2046 751 2052 752
rect 2046 747 2047 751
rect 2051 747 2052 751
rect 2046 746 2052 747
rect 2104 743 2106 752
rect 2142 751 2148 752
rect 2142 747 2143 751
rect 2147 747 2148 751
rect 2142 746 2148 747
rect 1823 742 1827 743
rect 1823 737 1827 738
rect 1855 742 1859 743
rect 1855 737 1859 738
rect 1887 742 1891 743
rect 1887 737 1891 738
rect 1943 742 1947 743
rect 1943 737 1947 738
rect 1951 742 1955 743
rect 1951 737 1955 738
rect 2023 742 2027 743
rect 2023 737 2027 738
rect 2031 742 2035 743
rect 2031 737 2035 738
rect 2103 742 2107 743
rect 2103 737 2107 738
rect 2119 742 2123 743
rect 2119 737 2123 738
rect 1798 731 1804 732
rect 1774 727 1780 728
rect 1774 723 1775 727
rect 1779 723 1780 727
rect 1798 727 1799 731
rect 1803 727 1804 731
rect 1856 728 1858 737
rect 1866 731 1872 732
rect 1798 726 1804 727
rect 1854 727 1860 728
rect 1774 722 1780 723
rect 1854 723 1855 727
rect 1859 723 1860 727
rect 1866 727 1867 731
rect 1871 727 1872 731
rect 1944 728 1946 737
rect 1954 731 1960 732
rect 1866 726 1872 727
rect 1942 727 1948 728
rect 1854 722 1860 723
rect 1868 700 1870 726
rect 1942 723 1943 727
rect 1947 723 1948 727
rect 1954 727 1955 731
rect 1959 727 1960 731
rect 2032 728 2034 737
rect 2042 731 2048 732
rect 1954 726 1960 727
rect 2030 727 2036 728
rect 1942 722 1948 723
rect 1956 700 1958 726
rect 2030 723 2031 727
rect 2035 723 2036 727
rect 2042 727 2043 731
rect 2047 727 2048 731
rect 2120 728 2122 737
rect 2042 726 2048 727
rect 2118 727 2124 728
rect 2030 722 2036 723
rect 2044 700 2046 726
rect 2118 723 2119 727
rect 2123 723 2124 727
rect 2118 722 2124 723
rect 2144 700 2146 746
rect 2192 743 2194 752
rect 2280 743 2282 752
rect 2302 751 2308 752
rect 2302 747 2303 751
rect 2307 747 2308 751
rect 2302 746 2308 747
rect 2191 742 2195 743
rect 2191 737 2195 738
rect 2207 742 2211 743
rect 2207 737 2211 738
rect 2279 742 2283 743
rect 2279 737 2283 738
rect 2295 742 2299 743
rect 2295 737 2299 738
rect 2198 731 2204 732
rect 2198 727 2199 731
rect 2203 727 2204 731
rect 2208 728 2210 737
rect 2286 731 2292 732
rect 2198 726 2204 727
rect 2206 727 2212 728
rect 2200 700 2202 726
rect 2206 723 2207 727
rect 2211 723 2212 727
rect 2286 727 2287 731
rect 2291 727 2292 731
rect 2296 728 2298 737
rect 2324 732 2326 778
rect 2358 757 2364 758
rect 2358 753 2359 757
rect 2363 753 2364 757
rect 2358 752 2364 753
rect 2384 752 2386 826
rect 2406 823 2407 827
rect 2411 823 2412 827
rect 2406 822 2412 823
rect 2408 811 2410 822
rect 2407 810 2411 811
rect 2407 805 2411 806
rect 2408 798 2410 805
rect 2406 797 2412 798
rect 2406 793 2407 797
rect 2411 793 2412 797
rect 2406 792 2412 793
rect 2406 780 2412 781
rect 2406 776 2407 780
rect 2411 776 2412 780
rect 2406 775 2412 776
rect 2360 743 2362 752
rect 2382 751 2388 752
rect 2382 747 2383 751
rect 2387 747 2388 751
rect 2382 746 2388 747
rect 2408 743 2410 775
rect 2359 742 2363 743
rect 2359 737 2363 738
rect 2407 742 2411 743
rect 2407 737 2411 738
rect 2322 731 2328 732
rect 2286 726 2292 727
rect 2294 727 2300 728
rect 2206 722 2212 723
rect 1706 699 1712 700
rect 1706 695 1707 699
rect 1711 695 1712 699
rect 1706 694 1712 695
rect 1718 699 1724 700
rect 1718 695 1719 699
rect 1723 695 1724 699
rect 1718 694 1724 695
rect 1866 699 1872 700
rect 1866 695 1867 699
rect 1871 695 1872 699
rect 1866 694 1872 695
rect 1954 699 1960 700
rect 1954 695 1955 699
rect 1959 695 1960 699
rect 1954 694 1960 695
rect 2042 699 2048 700
rect 2042 695 2043 699
rect 2047 695 2048 699
rect 2042 694 2048 695
rect 2134 699 2140 700
rect 2134 695 2135 699
rect 2139 695 2140 699
rect 2134 694 2140 695
rect 2142 699 2148 700
rect 2142 695 2143 699
rect 2147 695 2148 699
rect 2142 694 2148 695
rect 2198 699 2204 700
rect 2198 695 2199 699
rect 2203 695 2204 699
rect 2198 694 2204 695
rect 1694 680 1700 681
rect 1694 676 1695 680
rect 1699 676 1700 680
rect 1694 675 1700 676
rect 1774 680 1780 681
rect 1774 676 1775 680
rect 1779 676 1780 680
rect 1774 675 1780 676
rect 1854 680 1860 681
rect 1854 676 1855 680
rect 1859 676 1860 680
rect 1854 675 1860 676
rect 1942 680 1948 681
rect 1942 676 1943 680
rect 1947 676 1948 680
rect 1942 675 1948 676
rect 2030 680 2036 681
rect 2030 676 2031 680
rect 2035 676 2036 680
rect 2030 675 2036 676
rect 2118 680 2124 681
rect 2118 676 2119 680
rect 2123 676 2124 680
rect 2118 675 2124 676
rect 1687 674 1691 675
rect 1687 669 1691 670
rect 1695 674 1699 675
rect 1695 669 1699 670
rect 1743 674 1747 675
rect 1743 669 1747 670
rect 1775 674 1779 675
rect 1775 669 1779 670
rect 1799 674 1803 675
rect 1799 669 1803 670
rect 1855 674 1859 675
rect 1855 669 1859 670
rect 1871 674 1875 675
rect 1871 669 1875 670
rect 1943 674 1947 675
rect 1943 669 1947 670
rect 1951 674 1955 675
rect 1951 669 1955 670
rect 2031 674 2035 675
rect 2031 669 2035 670
rect 2047 674 2051 675
rect 2047 669 2051 670
rect 2119 674 2123 675
rect 2119 669 2123 670
rect 1686 668 1692 669
rect 1686 664 1687 668
rect 1691 664 1692 668
rect 1686 663 1692 664
rect 1742 668 1748 669
rect 1742 664 1743 668
rect 1747 664 1748 668
rect 1742 663 1748 664
rect 1798 668 1804 669
rect 1798 664 1799 668
rect 1803 664 1804 668
rect 1798 663 1804 664
rect 1870 668 1876 669
rect 1870 664 1871 668
rect 1875 664 1876 668
rect 1870 663 1876 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 1662 647 1668 648
rect 1662 643 1663 647
rect 1667 643 1668 647
rect 1662 642 1668 643
rect 1974 647 1980 648
rect 1974 643 1975 647
rect 1979 643 1980 647
rect 1974 642 1980 643
rect 2082 647 2088 648
rect 2082 643 2083 647
rect 2087 643 2088 647
rect 2082 642 2088 643
rect 1638 621 1644 622
rect 1638 617 1639 621
rect 1643 617 1644 621
rect 1638 616 1644 617
rect 1686 621 1692 622
rect 1686 617 1687 621
rect 1691 617 1692 621
rect 1686 616 1692 617
rect 1742 621 1748 622
rect 1742 617 1743 621
rect 1747 617 1748 621
rect 1742 616 1748 617
rect 1798 621 1804 622
rect 1798 617 1799 621
rect 1803 617 1804 621
rect 1798 616 1804 617
rect 1870 621 1876 622
rect 1870 617 1871 621
rect 1875 617 1876 621
rect 1870 616 1876 617
rect 1950 621 1956 622
rect 1950 617 1951 621
rect 1955 617 1956 621
rect 1950 616 1956 617
rect 1592 599 1594 616
rect 1606 615 1612 616
rect 1606 611 1607 615
rect 1611 611 1612 615
rect 1606 610 1612 611
rect 1640 599 1642 616
rect 1688 599 1690 616
rect 1744 599 1746 616
rect 1800 599 1802 616
rect 1872 599 1874 616
rect 1890 615 1896 616
rect 1890 611 1891 615
rect 1895 611 1896 615
rect 1890 610 1896 611
rect 1591 598 1595 599
rect 1591 593 1595 594
rect 1599 598 1603 599
rect 1599 593 1603 594
rect 1639 598 1643 599
rect 1639 593 1643 594
rect 1679 598 1683 599
rect 1679 593 1683 594
rect 1687 598 1691 599
rect 1687 593 1691 594
rect 1719 598 1723 599
rect 1719 593 1723 594
rect 1743 598 1747 599
rect 1743 593 1747 594
rect 1759 598 1763 599
rect 1759 593 1763 594
rect 1799 598 1803 599
rect 1799 593 1803 594
rect 1807 598 1811 599
rect 1807 593 1811 594
rect 1855 598 1859 599
rect 1855 593 1859 594
rect 1871 598 1875 599
rect 1871 593 1875 594
rect 1582 587 1588 588
rect 1558 583 1564 584
rect 1558 579 1559 583
rect 1563 579 1564 583
rect 1582 583 1583 587
rect 1587 583 1588 587
rect 1600 584 1602 593
rect 1610 587 1616 588
rect 1582 582 1588 583
rect 1598 583 1604 584
rect 1558 578 1564 579
rect 1598 579 1599 583
rect 1603 579 1604 583
rect 1610 583 1611 587
rect 1615 583 1616 587
rect 1640 584 1642 593
rect 1650 587 1656 588
rect 1610 582 1616 583
rect 1638 583 1644 584
rect 1598 578 1604 579
rect 1238 558 1244 559
rect 1278 560 1284 561
rect 1142 556 1148 557
rect 1142 552 1143 556
rect 1147 552 1148 556
rect 1142 551 1148 552
rect 1190 556 1196 557
rect 1190 552 1191 556
rect 1195 552 1196 556
rect 1190 551 1196 552
rect 1144 547 1146 551
rect 1192 547 1194 551
rect 1240 547 1242 558
rect 1278 556 1279 560
rect 1283 556 1284 560
rect 1612 556 1614 582
rect 1638 579 1639 583
rect 1643 579 1644 583
rect 1650 583 1651 587
rect 1655 583 1656 587
rect 1680 584 1682 593
rect 1706 587 1712 588
rect 1650 582 1656 583
rect 1678 583 1684 584
rect 1638 578 1644 579
rect 1652 556 1654 582
rect 1678 579 1679 583
rect 1683 579 1684 583
rect 1706 583 1707 587
rect 1711 583 1712 587
rect 1720 584 1722 593
rect 1746 587 1752 588
rect 1706 582 1712 583
rect 1718 583 1724 584
rect 1678 578 1684 579
rect 1666 575 1672 576
rect 1666 571 1667 575
rect 1671 571 1672 575
rect 1666 570 1672 571
rect 1668 556 1670 570
rect 1278 555 1284 556
rect 1610 555 1616 556
rect 1610 551 1611 555
rect 1615 551 1616 555
rect 1610 550 1616 551
rect 1650 555 1656 556
rect 1650 551 1651 555
rect 1655 551 1656 555
rect 1650 550 1656 551
rect 1666 555 1672 556
rect 1666 551 1667 555
rect 1671 551 1672 555
rect 1666 550 1672 551
rect 1708 548 1710 582
rect 1718 579 1719 583
rect 1723 579 1724 583
rect 1746 583 1747 587
rect 1751 583 1752 587
rect 1760 584 1762 593
rect 1798 587 1804 588
rect 1746 582 1752 583
rect 1758 583 1764 584
rect 1718 578 1724 579
rect 1748 564 1750 582
rect 1758 579 1759 583
rect 1763 579 1764 583
rect 1798 583 1799 587
rect 1803 583 1804 587
rect 1808 584 1810 593
rect 1856 584 1858 593
rect 1798 582 1804 583
rect 1806 583 1812 584
rect 1758 578 1764 579
rect 1746 563 1752 564
rect 1746 559 1747 563
rect 1751 559 1752 563
rect 1746 558 1752 559
rect 1800 556 1802 582
rect 1806 579 1807 583
rect 1811 579 1812 583
rect 1806 578 1812 579
rect 1854 583 1860 584
rect 1854 579 1855 583
rect 1859 579 1860 583
rect 1854 578 1860 579
rect 1892 556 1894 610
rect 1952 599 1954 616
rect 1911 598 1915 599
rect 1911 593 1915 594
rect 1951 598 1955 599
rect 1951 593 1955 594
rect 1967 598 1971 599
rect 1967 593 1971 594
rect 1902 587 1908 588
rect 1902 583 1903 587
rect 1907 583 1908 587
rect 1912 584 1914 593
rect 1958 587 1964 588
rect 1902 582 1908 583
rect 1910 583 1916 584
rect 1904 556 1906 582
rect 1910 579 1911 583
rect 1915 579 1916 583
rect 1958 583 1959 587
rect 1963 583 1964 587
rect 1968 584 1970 593
rect 1976 592 1978 642
rect 2046 621 2052 622
rect 2046 617 2047 621
rect 2051 617 2052 621
rect 2046 616 2052 617
rect 2084 616 2086 642
rect 2136 616 2138 694
rect 2206 680 2212 681
rect 2206 676 2207 680
rect 2211 676 2212 680
rect 2206 675 2212 676
rect 2151 674 2155 675
rect 2151 669 2155 670
rect 2207 674 2211 675
rect 2207 669 2211 670
rect 2263 674 2267 675
rect 2263 669 2267 670
rect 2150 668 2156 669
rect 2150 664 2151 668
rect 2155 664 2156 668
rect 2150 663 2156 664
rect 2262 668 2268 669
rect 2262 664 2263 668
rect 2267 664 2268 668
rect 2262 663 2268 664
rect 2288 648 2290 726
rect 2294 723 2295 727
rect 2299 723 2300 727
rect 2322 727 2323 731
rect 2327 727 2328 731
rect 2360 728 2362 737
rect 2370 731 2376 732
rect 2322 726 2328 727
rect 2358 727 2364 728
rect 2294 722 2300 723
rect 2358 723 2359 727
rect 2363 723 2364 727
rect 2370 727 2371 731
rect 2375 727 2376 731
rect 2370 726 2376 727
rect 2358 722 2364 723
rect 2372 700 2374 726
rect 2408 705 2410 737
rect 2406 704 2412 705
rect 2406 700 2407 704
rect 2411 700 2412 704
rect 2370 699 2376 700
rect 2370 695 2371 699
rect 2375 695 2376 699
rect 2370 694 2376 695
rect 2382 699 2388 700
rect 2406 699 2412 700
rect 2382 695 2383 699
rect 2387 695 2388 699
rect 2382 694 2388 695
rect 2294 680 2300 681
rect 2294 676 2295 680
rect 2299 676 2300 680
rect 2294 675 2300 676
rect 2358 680 2364 681
rect 2358 676 2359 680
rect 2363 676 2364 680
rect 2358 675 2364 676
rect 2295 674 2299 675
rect 2295 669 2299 670
rect 2359 674 2363 675
rect 2359 669 2363 670
rect 2358 668 2364 669
rect 2358 664 2359 668
rect 2363 664 2364 668
rect 2358 663 2364 664
rect 2286 647 2292 648
rect 2286 643 2287 647
rect 2291 643 2292 647
rect 2286 642 2292 643
rect 2150 621 2156 622
rect 2150 617 2151 621
rect 2155 617 2156 621
rect 2150 616 2156 617
rect 2262 621 2268 622
rect 2262 617 2263 621
rect 2267 617 2268 621
rect 2262 616 2268 617
rect 2358 621 2364 622
rect 2358 617 2359 621
rect 2363 617 2364 621
rect 2358 616 2364 617
rect 2384 616 2386 694
rect 2406 687 2412 688
rect 2406 683 2407 687
rect 2411 683 2412 687
rect 2406 682 2412 683
rect 2408 675 2410 682
rect 2407 674 2411 675
rect 2407 669 2411 670
rect 2408 662 2410 669
rect 2406 661 2412 662
rect 2406 657 2407 661
rect 2411 657 2412 661
rect 2406 656 2412 657
rect 2406 644 2412 645
rect 2406 640 2407 644
rect 2411 640 2412 644
rect 2406 639 2412 640
rect 2048 599 2050 616
rect 2082 615 2088 616
rect 2082 611 2083 615
rect 2087 611 2088 615
rect 2082 610 2088 611
rect 2134 615 2140 616
rect 2134 611 2135 615
rect 2139 611 2140 615
rect 2134 610 2140 611
rect 2152 599 2154 616
rect 2264 599 2266 616
rect 2360 599 2362 616
rect 2382 615 2388 616
rect 2382 611 2383 615
rect 2387 611 2388 615
rect 2382 610 2388 611
rect 2408 599 2410 639
rect 2031 598 2035 599
rect 2031 593 2035 594
rect 2047 598 2051 599
rect 2047 593 2051 594
rect 2095 598 2099 599
rect 2095 593 2099 594
rect 2151 598 2155 599
rect 2151 593 2155 594
rect 2167 598 2171 599
rect 2167 593 2171 594
rect 2239 598 2243 599
rect 2239 593 2243 594
rect 2263 598 2267 599
rect 2263 593 2267 594
rect 2311 598 2315 599
rect 2311 593 2315 594
rect 2359 598 2363 599
rect 2359 593 2363 594
rect 2407 598 2411 599
rect 2407 593 2411 594
rect 1974 591 1980 592
rect 1974 587 1975 591
rect 1979 587 1980 591
rect 1974 586 1980 587
rect 2032 584 2034 593
rect 2042 587 2048 588
rect 1958 582 1964 583
rect 1966 583 1972 584
rect 1910 578 1916 579
rect 1734 555 1740 556
rect 1734 551 1735 555
rect 1739 551 1740 555
rect 1734 550 1740 551
rect 1798 555 1804 556
rect 1798 551 1799 555
rect 1803 551 1804 555
rect 1798 550 1804 551
rect 1890 555 1896 556
rect 1890 551 1891 555
rect 1895 551 1896 555
rect 1890 550 1896 551
rect 1902 555 1908 556
rect 1902 551 1903 555
rect 1907 551 1908 555
rect 1902 550 1908 551
rect 1706 547 1712 548
rect 1143 546 1147 547
rect 1143 541 1147 542
rect 1191 546 1195 547
rect 1191 541 1195 542
rect 1239 546 1243 547
rect 1239 541 1243 542
rect 1278 543 1284 544
rect 1240 534 1242 541
rect 1278 539 1279 543
rect 1283 539 1284 543
rect 1706 543 1707 547
rect 1711 543 1712 547
rect 1706 542 1712 543
rect 1278 538 1284 539
rect 1238 533 1244 534
rect 1238 529 1239 533
rect 1243 529 1244 533
rect 1280 531 1282 538
rect 1558 536 1564 537
rect 1558 532 1559 536
rect 1563 532 1564 536
rect 1558 531 1564 532
rect 1598 536 1604 537
rect 1598 532 1599 536
rect 1603 532 1604 536
rect 1598 531 1604 532
rect 1638 536 1644 537
rect 1638 532 1639 536
rect 1643 532 1644 536
rect 1638 531 1644 532
rect 1678 536 1684 537
rect 1678 532 1679 536
rect 1683 532 1684 536
rect 1678 531 1684 532
rect 1718 536 1724 537
rect 1718 532 1719 536
rect 1723 532 1724 536
rect 1718 531 1724 532
rect 1238 528 1244 529
rect 1279 530 1283 531
rect 1279 525 1283 526
rect 1407 530 1411 531
rect 1407 525 1411 526
rect 1447 530 1451 531
rect 1447 525 1451 526
rect 1487 530 1491 531
rect 1487 525 1491 526
rect 1535 530 1539 531
rect 1535 525 1539 526
rect 1559 530 1563 531
rect 1559 525 1563 526
rect 1591 530 1595 531
rect 1591 525 1595 526
rect 1599 530 1603 531
rect 1599 525 1603 526
rect 1639 530 1643 531
rect 1639 525 1643 526
rect 1647 530 1651 531
rect 1647 525 1651 526
rect 1679 530 1683 531
rect 1679 525 1683 526
rect 1711 530 1715 531
rect 1711 525 1715 526
rect 1719 530 1723 531
rect 1719 525 1723 526
rect 1280 518 1282 525
rect 1406 524 1412 525
rect 1406 520 1407 524
rect 1411 520 1412 524
rect 1406 519 1412 520
rect 1446 524 1452 525
rect 1446 520 1447 524
rect 1451 520 1452 524
rect 1446 519 1452 520
rect 1486 524 1492 525
rect 1486 520 1487 524
rect 1491 520 1492 524
rect 1486 519 1492 520
rect 1534 524 1540 525
rect 1534 520 1535 524
rect 1539 520 1540 524
rect 1534 519 1540 520
rect 1590 524 1596 525
rect 1590 520 1591 524
rect 1595 520 1596 524
rect 1590 519 1596 520
rect 1646 524 1652 525
rect 1646 520 1647 524
rect 1651 520 1652 524
rect 1646 519 1652 520
rect 1710 524 1716 525
rect 1710 520 1711 524
rect 1715 520 1716 524
rect 1710 519 1716 520
rect 1278 517 1284 518
rect 1238 516 1244 517
rect 1238 512 1239 516
rect 1243 512 1244 516
rect 1278 513 1279 517
rect 1283 513 1284 517
rect 1278 512 1284 513
rect 1238 511 1244 512
rect 982 487 988 488
rect 982 483 983 487
rect 987 483 988 487
rect 982 482 988 483
rect 1000 479 1002 488
rect 1080 479 1082 488
rect 1094 487 1100 488
rect 1094 483 1095 487
rect 1099 483 1100 487
rect 1094 482 1100 483
rect 1240 479 1242 511
rect 1454 503 1460 504
rect 1278 500 1284 501
rect 1278 496 1279 500
rect 1283 496 1284 500
rect 1454 499 1455 503
rect 1459 499 1460 503
rect 1454 498 1460 499
rect 1494 503 1500 504
rect 1494 499 1495 503
rect 1499 499 1500 503
rect 1494 498 1500 499
rect 1278 495 1284 496
rect 999 478 1003 479
rect 999 473 1003 474
rect 1015 478 1019 479
rect 1015 473 1019 474
rect 1079 478 1083 479
rect 1079 473 1083 474
rect 1239 478 1243 479
rect 1239 473 1243 474
rect 974 467 980 468
rect 898 462 904 463
rect 950 463 956 464
rect 886 458 892 459
rect 514 435 520 436
rect 514 431 515 435
rect 519 431 520 435
rect 514 430 520 431
rect 574 435 580 436
rect 574 431 575 435
rect 579 431 580 435
rect 574 430 580 431
rect 582 435 588 436
rect 582 431 583 435
rect 587 431 588 435
rect 582 430 588 431
rect 658 435 664 436
rect 658 431 659 435
rect 663 431 664 435
rect 658 430 664 431
rect 686 435 692 436
rect 686 431 687 435
rect 691 431 692 435
rect 686 430 692 431
rect 750 435 756 436
rect 750 431 751 435
rect 755 431 756 435
rect 750 430 756 431
rect 814 435 820 436
rect 814 431 815 435
rect 819 431 820 435
rect 814 430 820 431
rect 878 435 884 436
rect 878 431 879 435
rect 883 431 884 435
rect 878 430 884 431
rect 438 416 444 417
rect 438 412 439 416
rect 443 412 444 416
rect 438 411 444 412
rect 502 416 508 417
rect 502 412 503 416
rect 507 412 508 416
rect 502 411 508 412
rect 566 416 572 417
rect 566 412 567 416
rect 571 412 572 416
rect 566 411 572 412
rect 440 407 442 411
rect 504 407 506 411
rect 568 407 570 411
rect 439 406 443 407
rect 439 401 443 402
rect 471 406 475 407
rect 471 401 475 402
rect 503 406 507 407
rect 503 401 507 402
rect 543 406 547 407
rect 543 401 547 402
rect 567 406 571 407
rect 567 401 571 402
rect 470 400 476 401
rect 470 396 471 400
rect 475 396 476 400
rect 470 395 476 396
rect 542 400 548 401
rect 542 396 543 400
rect 547 396 548 400
rect 542 395 548 396
rect 406 387 412 388
rect 406 383 407 387
rect 411 383 412 387
rect 406 382 412 383
rect 198 379 204 380
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 198 375 199 379
rect 203 375 204 379
rect 198 374 204 375
rect 238 379 244 380
rect 238 375 239 379
rect 243 375 244 379
rect 238 374 244 375
rect 286 379 292 380
rect 286 375 287 379
rect 291 375 292 379
rect 286 374 292 375
rect 506 379 512 380
rect 506 375 507 379
rect 511 375 512 379
rect 506 374 512 375
rect 110 371 116 372
rect 112 331 114 371
rect 200 363 202 374
rect 200 361 210 363
rect 142 353 148 354
rect 142 349 143 353
rect 147 349 148 353
rect 142 348 148 349
rect 182 353 188 354
rect 182 349 183 353
rect 187 349 188 353
rect 182 348 188 349
rect 208 348 210 361
rect 222 353 228 354
rect 222 349 223 353
rect 227 349 228 353
rect 222 348 228 349
rect 240 348 242 374
rect 270 353 276 354
rect 270 349 271 353
rect 275 349 276 353
rect 270 348 276 349
rect 288 348 290 374
rect 462 371 468 372
rect 462 367 463 371
rect 467 367 468 371
rect 462 366 468 367
rect 334 353 340 354
rect 334 349 335 353
rect 339 349 340 353
rect 334 348 340 349
rect 398 353 404 354
rect 398 349 399 353
rect 403 349 404 353
rect 398 348 404 349
rect 144 331 146 348
rect 184 331 186 348
rect 198 347 204 348
rect 198 343 199 347
rect 203 343 204 347
rect 198 342 204 343
rect 206 347 212 348
rect 206 343 207 347
rect 211 343 212 347
rect 206 342 212 343
rect 111 330 115 331
rect 111 325 115 326
rect 135 330 139 331
rect 135 325 139 326
rect 143 330 147 331
rect 143 325 147 326
rect 175 330 179 331
rect 175 325 179 326
rect 183 330 187 331
rect 183 325 187 326
rect 112 293 114 325
rect 136 316 138 325
rect 158 319 164 320
rect 134 315 140 316
rect 134 311 135 315
rect 139 311 140 315
rect 158 315 159 319
rect 163 315 164 319
rect 176 316 178 325
rect 158 314 164 315
rect 174 315 180 316
rect 134 310 140 311
rect 110 292 116 293
rect 110 288 111 292
rect 115 288 116 292
rect 110 287 116 288
rect 150 279 156 280
rect 110 275 116 276
rect 110 271 111 275
rect 115 271 116 275
rect 150 275 151 279
rect 155 275 156 279
rect 150 274 156 275
rect 110 270 116 271
rect 112 255 114 270
rect 134 268 140 269
rect 134 264 135 268
rect 139 264 140 268
rect 134 263 140 264
rect 136 255 138 263
rect 111 254 115 255
rect 111 249 115 250
rect 135 254 139 255
rect 135 249 139 250
rect 112 242 114 249
rect 134 248 140 249
rect 134 244 135 248
rect 139 244 140 248
rect 134 243 140 244
rect 110 241 116 242
rect 110 237 111 241
rect 115 237 116 241
rect 110 236 116 237
rect 110 224 116 225
rect 110 220 111 224
rect 115 220 116 224
rect 110 219 116 220
rect 112 155 114 219
rect 134 201 140 202
rect 134 197 135 201
rect 139 197 140 201
rect 134 196 140 197
rect 152 196 154 274
rect 160 228 162 314
rect 174 311 175 315
rect 179 311 180 315
rect 174 310 180 311
rect 200 288 202 342
rect 224 331 226 348
rect 238 347 244 348
rect 238 343 239 347
rect 243 343 244 347
rect 238 342 244 343
rect 272 331 274 348
rect 286 347 292 348
rect 286 343 287 347
rect 291 343 292 347
rect 286 342 292 343
rect 336 331 338 348
rect 400 331 402 348
rect 215 330 219 331
rect 215 325 219 326
rect 223 330 227 331
rect 223 325 227 326
rect 255 330 259 331
rect 255 325 259 326
rect 271 330 275 331
rect 271 325 275 326
rect 295 330 299 331
rect 295 325 299 326
rect 335 330 339 331
rect 335 325 339 326
rect 391 330 395 331
rect 391 325 395 326
rect 399 330 403 331
rect 399 325 403 326
rect 447 330 451 331
rect 447 325 451 326
rect 216 316 218 325
rect 230 323 236 324
rect 230 319 231 323
rect 235 319 236 323
rect 230 318 236 319
rect 242 319 248 320
rect 214 315 220 316
rect 214 311 215 315
rect 219 311 220 315
rect 214 310 220 311
rect 232 288 234 318
rect 242 315 243 319
rect 247 315 248 319
rect 256 316 258 325
rect 266 319 272 320
rect 242 314 248 315
rect 254 315 260 316
rect 198 287 204 288
rect 198 283 199 287
rect 203 283 204 287
rect 198 282 204 283
rect 230 287 236 288
rect 230 283 231 287
rect 235 283 236 287
rect 244 286 246 314
rect 254 311 255 315
rect 259 311 260 315
rect 266 315 267 319
rect 271 315 272 319
rect 296 316 298 325
rect 322 319 328 320
rect 266 314 272 315
rect 294 315 300 316
rect 254 310 260 311
rect 268 296 270 314
rect 294 311 295 315
rect 299 311 300 315
rect 322 315 323 319
rect 327 315 328 319
rect 336 316 338 325
rect 382 319 388 320
rect 322 314 328 315
rect 334 315 340 316
rect 294 310 300 311
rect 324 296 326 314
rect 334 311 335 315
rect 339 311 340 315
rect 382 315 383 319
rect 387 315 388 319
rect 392 316 394 325
rect 438 319 444 320
rect 382 314 388 315
rect 390 315 396 316
rect 334 310 340 311
rect 266 295 272 296
rect 266 291 267 295
rect 271 291 272 295
rect 266 290 272 291
rect 322 295 328 296
rect 322 291 323 295
rect 327 291 328 295
rect 322 290 328 291
rect 384 288 386 314
rect 390 311 391 315
rect 395 311 396 315
rect 438 315 439 319
rect 443 315 444 319
rect 448 316 450 325
rect 464 320 466 366
rect 470 353 476 354
rect 470 349 471 353
rect 475 349 476 353
rect 470 348 476 349
rect 508 348 510 374
rect 542 353 548 354
rect 542 349 543 353
rect 547 349 548 353
rect 584 352 586 430
rect 630 416 636 417
rect 630 412 631 416
rect 635 412 636 416
rect 630 411 636 412
rect 694 416 700 417
rect 694 412 695 416
rect 699 412 700 416
rect 694 411 700 412
rect 758 416 764 417
rect 758 412 759 416
rect 763 412 764 416
rect 758 411 764 412
rect 822 416 828 417
rect 822 412 823 416
rect 827 412 828 416
rect 822 411 828 412
rect 886 416 892 417
rect 886 412 887 416
rect 891 412 892 416
rect 886 411 892 412
rect 632 407 634 411
rect 696 407 698 411
rect 760 407 762 411
rect 824 407 826 411
rect 888 407 890 411
rect 615 406 619 407
rect 615 401 619 402
rect 631 406 635 407
rect 631 401 635 402
rect 687 406 691 407
rect 687 401 691 402
rect 695 406 699 407
rect 695 401 699 402
rect 751 406 755 407
rect 751 401 755 402
rect 759 406 763 407
rect 759 401 763 402
rect 807 406 811 407
rect 807 401 811 402
rect 823 406 827 407
rect 823 401 827 402
rect 863 406 867 407
rect 863 401 867 402
rect 887 406 891 407
rect 887 401 891 402
rect 614 400 620 401
rect 614 396 615 400
rect 619 396 620 400
rect 614 395 620 396
rect 686 400 692 401
rect 686 396 687 400
rect 691 396 692 400
rect 686 395 692 396
rect 750 400 756 401
rect 750 396 751 400
rect 755 396 756 400
rect 750 395 756 396
rect 806 400 812 401
rect 806 396 807 400
rect 811 396 812 400
rect 806 395 812 396
rect 862 400 868 401
rect 862 396 863 400
rect 867 396 868 400
rect 862 395 868 396
rect 900 380 902 462
rect 950 459 951 463
rect 955 459 956 463
rect 974 463 975 467
rect 979 463 980 467
rect 1016 464 1018 473
rect 1026 467 1032 468
rect 974 462 980 463
rect 1014 463 1020 464
rect 950 458 956 459
rect 1014 459 1015 463
rect 1019 459 1020 463
rect 1026 463 1027 467
rect 1031 463 1032 467
rect 1026 462 1032 463
rect 1014 458 1020 459
rect 1028 436 1030 462
rect 1240 441 1242 473
rect 1280 463 1282 495
rect 1406 477 1412 478
rect 1406 473 1407 477
rect 1411 473 1412 477
rect 1406 472 1412 473
rect 1446 477 1452 478
rect 1446 473 1447 477
rect 1451 473 1452 477
rect 1446 472 1452 473
rect 1456 472 1458 498
rect 1486 477 1492 478
rect 1486 473 1487 477
rect 1491 473 1492 477
rect 1486 472 1492 473
rect 1496 472 1498 498
rect 1534 477 1540 478
rect 1534 473 1535 477
rect 1539 473 1540 477
rect 1534 472 1540 473
rect 1590 477 1596 478
rect 1590 473 1591 477
rect 1595 473 1596 477
rect 1590 472 1596 473
rect 1646 477 1652 478
rect 1646 473 1647 477
rect 1651 473 1652 477
rect 1646 472 1652 473
rect 1710 477 1716 478
rect 1710 473 1711 477
rect 1715 473 1716 477
rect 1710 472 1716 473
rect 1736 472 1738 550
rect 1758 536 1764 537
rect 1758 532 1759 536
rect 1763 532 1764 536
rect 1758 531 1764 532
rect 1806 536 1812 537
rect 1806 532 1807 536
rect 1811 532 1812 536
rect 1806 531 1812 532
rect 1854 536 1860 537
rect 1854 532 1855 536
rect 1859 532 1860 536
rect 1854 531 1860 532
rect 1910 536 1916 537
rect 1910 532 1911 536
rect 1915 532 1916 536
rect 1910 531 1916 532
rect 1759 530 1763 531
rect 1759 525 1763 526
rect 1783 530 1787 531
rect 1783 525 1787 526
rect 1807 530 1811 531
rect 1807 525 1811 526
rect 1855 530 1859 531
rect 1855 525 1859 526
rect 1863 530 1867 531
rect 1863 525 1867 526
rect 1911 530 1915 531
rect 1911 525 1915 526
rect 1943 530 1947 531
rect 1943 525 1947 526
rect 1782 524 1788 525
rect 1782 520 1783 524
rect 1787 520 1788 524
rect 1782 519 1788 520
rect 1862 524 1868 525
rect 1862 520 1863 524
rect 1867 520 1868 524
rect 1862 519 1868 520
rect 1942 524 1948 525
rect 1942 520 1943 524
rect 1947 520 1948 524
rect 1942 519 1948 520
rect 1960 504 1962 582
rect 1966 579 1967 583
rect 1971 579 1972 583
rect 1966 578 1972 579
rect 2030 583 2036 584
rect 2030 579 2031 583
rect 2035 579 2036 583
rect 2042 583 2043 587
rect 2047 583 2048 587
rect 2096 584 2098 593
rect 2106 587 2112 588
rect 2042 582 2048 583
rect 2094 583 2100 584
rect 2030 578 2036 579
rect 2044 556 2046 582
rect 2094 579 2095 583
rect 2099 579 2100 583
rect 2106 583 2107 587
rect 2111 583 2112 587
rect 2168 584 2170 593
rect 2230 587 2236 588
rect 2106 582 2112 583
rect 2166 583 2172 584
rect 2094 578 2100 579
rect 2108 556 2110 582
rect 2166 579 2167 583
rect 2171 579 2172 583
rect 2230 583 2231 587
rect 2235 583 2236 587
rect 2240 584 2242 593
rect 2302 587 2308 588
rect 2230 582 2236 583
rect 2238 583 2244 584
rect 2166 578 2172 579
rect 2232 556 2234 582
rect 2238 579 2239 583
rect 2243 579 2244 583
rect 2302 583 2303 587
rect 2307 583 2308 587
rect 2312 584 2314 593
rect 2350 587 2356 588
rect 2302 582 2308 583
rect 2310 583 2316 584
rect 2238 578 2244 579
rect 2042 555 2048 556
rect 2042 551 2043 555
rect 2047 551 2048 555
rect 2042 550 2048 551
rect 2106 555 2112 556
rect 2106 551 2107 555
rect 2111 551 2112 555
rect 2106 550 2112 551
rect 2122 555 2128 556
rect 2122 551 2123 555
rect 2127 551 2128 555
rect 2122 550 2128 551
rect 2230 555 2236 556
rect 2230 551 2231 555
rect 2235 551 2236 555
rect 2230 550 2236 551
rect 1966 536 1972 537
rect 1966 532 1967 536
rect 1971 532 1972 536
rect 1966 531 1972 532
rect 2030 536 2036 537
rect 2030 532 2031 536
rect 2035 532 2036 536
rect 2030 531 2036 532
rect 2094 536 2100 537
rect 2094 532 2095 536
rect 2099 532 2100 536
rect 2094 531 2100 532
rect 1967 530 1971 531
rect 1967 525 1971 526
rect 2023 530 2027 531
rect 2023 525 2027 526
rect 2031 530 2035 531
rect 2031 525 2035 526
rect 2095 530 2099 531
rect 2095 525 2099 526
rect 2103 530 2107 531
rect 2103 525 2107 526
rect 2022 524 2028 525
rect 2022 520 2023 524
rect 2027 520 2028 524
rect 2022 519 2028 520
rect 2102 524 2108 525
rect 2102 520 2103 524
rect 2107 520 2108 524
rect 2102 519 2108 520
rect 1878 503 1884 504
rect 1878 499 1879 503
rect 1883 499 1884 503
rect 1878 498 1884 499
rect 1950 503 1956 504
rect 1950 499 1951 503
rect 1955 499 1956 503
rect 1950 498 1956 499
rect 1958 503 1964 504
rect 1958 499 1959 503
rect 1963 499 1964 503
rect 1958 498 1964 499
rect 2038 503 2044 504
rect 2038 499 2039 503
rect 2043 499 2044 503
rect 2038 498 2044 499
rect 1758 495 1764 496
rect 1758 491 1759 495
rect 1763 491 1764 495
rect 1758 490 1764 491
rect 1408 463 1410 472
rect 1448 463 1450 472
rect 1454 471 1460 472
rect 1454 467 1455 471
rect 1459 467 1460 471
rect 1454 466 1460 467
rect 1488 463 1490 472
rect 1494 471 1500 472
rect 1494 467 1495 471
rect 1499 467 1500 471
rect 1494 466 1500 467
rect 1536 463 1538 472
rect 1592 463 1594 472
rect 1648 463 1650 472
rect 1712 463 1714 472
rect 1734 471 1740 472
rect 1734 467 1735 471
rect 1739 467 1740 471
rect 1734 466 1740 467
rect 1279 462 1283 463
rect 1279 457 1283 458
rect 1303 462 1307 463
rect 1303 457 1307 458
rect 1343 462 1347 463
rect 1343 457 1347 458
rect 1383 462 1387 463
rect 1383 457 1387 458
rect 1407 462 1411 463
rect 1407 457 1411 458
rect 1447 462 1451 463
rect 1447 457 1451 458
rect 1487 462 1491 463
rect 1487 457 1491 458
rect 1535 462 1539 463
rect 1535 457 1539 458
rect 1591 462 1595 463
rect 1591 457 1595 458
rect 1631 462 1635 463
rect 1631 457 1635 458
rect 1647 462 1651 463
rect 1647 457 1651 458
rect 1711 462 1715 463
rect 1711 457 1715 458
rect 1735 462 1739 463
rect 1735 457 1739 458
rect 1238 440 1244 441
rect 1238 436 1239 440
rect 1243 436 1244 440
rect 1026 435 1032 436
rect 1026 431 1027 435
rect 1031 431 1032 435
rect 1026 430 1032 431
rect 1054 435 1060 436
rect 1238 435 1244 436
rect 1054 431 1055 435
rect 1059 431 1060 435
rect 1054 430 1060 431
rect 950 416 956 417
rect 950 412 951 416
rect 955 412 956 416
rect 950 411 956 412
rect 1014 416 1020 417
rect 1014 412 1015 416
rect 1019 412 1020 416
rect 1014 411 1020 412
rect 952 407 954 411
rect 1016 407 1018 411
rect 919 406 923 407
rect 919 401 923 402
rect 951 406 955 407
rect 951 401 955 402
rect 975 406 979 407
rect 975 401 979 402
rect 1015 406 1019 407
rect 1015 401 1019 402
rect 1031 406 1035 407
rect 1031 401 1035 402
rect 918 400 924 401
rect 918 396 919 400
rect 923 396 924 400
rect 918 395 924 396
rect 974 400 980 401
rect 974 396 975 400
rect 979 396 980 400
rect 974 395 980 396
rect 1030 400 1036 401
rect 1030 396 1031 400
rect 1035 396 1036 400
rect 1030 395 1036 396
rect 702 379 708 380
rect 702 375 703 379
rect 707 375 708 379
rect 702 374 708 375
rect 766 379 772 380
rect 766 375 767 379
rect 771 375 772 379
rect 766 374 772 375
rect 822 379 828 380
rect 822 375 823 379
rect 827 375 828 379
rect 822 374 828 375
rect 878 379 884 380
rect 878 375 879 379
rect 883 375 884 379
rect 878 374 884 375
rect 898 379 904 380
rect 898 375 899 379
rect 903 375 904 379
rect 898 374 904 375
rect 906 379 912 380
rect 906 375 907 379
rect 911 375 912 379
rect 906 374 912 375
rect 614 353 620 354
rect 542 348 548 349
rect 582 351 588 352
rect 472 331 474 348
rect 506 347 512 348
rect 506 343 507 347
rect 511 343 512 347
rect 506 342 512 343
rect 544 331 546 348
rect 582 347 583 351
rect 587 347 588 351
rect 614 349 615 353
rect 619 349 620 353
rect 614 348 620 349
rect 686 353 692 354
rect 686 349 687 353
rect 691 349 692 353
rect 686 348 692 349
rect 704 348 706 374
rect 750 353 756 354
rect 750 349 751 353
rect 755 349 756 353
rect 750 348 756 349
rect 768 348 770 374
rect 806 353 812 354
rect 806 349 807 353
rect 811 349 812 353
rect 806 348 812 349
rect 824 348 826 374
rect 862 353 868 354
rect 862 349 863 353
rect 867 349 868 353
rect 862 348 868 349
rect 880 348 882 374
rect 582 346 588 347
rect 616 331 618 348
rect 630 347 636 348
rect 630 343 631 347
rect 635 343 636 347
rect 630 342 636 343
rect 471 330 475 331
rect 471 325 475 326
rect 495 330 499 331
rect 495 325 499 326
rect 543 330 547 331
rect 543 325 547 326
rect 591 330 595 331
rect 591 325 595 326
rect 615 330 619 331
rect 615 325 619 326
rect 462 319 468 320
rect 438 314 444 315
rect 446 315 452 316
rect 390 310 396 311
rect 440 288 442 314
rect 446 311 447 315
rect 451 311 452 315
rect 462 315 463 319
rect 467 315 468 319
rect 496 316 498 325
rect 534 319 540 320
rect 462 314 468 315
rect 494 315 500 316
rect 446 310 452 311
rect 494 311 495 315
rect 499 311 500 315
rect 534 315 535 319
rect 539 315 540 319
rect 544 316 546 325
rect 592 316 594 325
rect 534 314 540 315
rect 542 315 548 316
rect 494 310 500 311
rect 536 288 538 314
rect 542 311 543 315
rect 547 311 548 315
rect 542 310 548 311
rect 590 315 596 316
rect 590 311 591 315
rect 595 311 596 315
rect 590 310 596 311
rect 632 288 634 342
rect 688 331 690 348
rect 702 347 708 348
rect 702 343 703 347
rect 707 343 708 347
rect 702 342 708 343
rect 752 331 754 348
rect 766 347 772 348
rect 766 343 767 347
rect 771 343 772 347
rect 766 342 772 343
rect 808 331 810 348
rect 822 347 828 348
rect 822 343 823 347
rect 827 343 828 347
rect 822 342 828 343
rect 864 331 866 348
rect 878 347 884 348
rect 878 343 879 347
rect 883 343 884 347
rect 878 342 884 343
rect 639 330 643 331
rect 639 325 643 326
rect 687 330 691 331
rect 687 325 691 326
rect 735 330 739 331
rect 735 325 739 326
rect 751 330 755 331
rect 751 325 755 326
rect 783 330 787 331
rect 783 325 787 326
rect 807 330 811 331
rect 807 325 811 326
rect 839 330 843 331
rect 839 325 843 326
rect 863 330 867 331
rect 863 325 867 326
rect 640 316 642 325
rect 654 323 660 324
rect 654 319 655 323
rect 659 319 660 323
rect 654 318 660 319
rect 678 319 684 320
rect 638 315 644 316
rect 638 311 639 315
rect 643 311 644 315
rect 638 310 644 311
rect 656 288 658 318
rect 678 315 679 319
rect 683 315 684 319
rect 688 316 690 325
rect 726 319 732 320
rect 678 314 684 315
rect 686 315 692 316
rect 680 288 682 314
rect 686 311 687 315
rect 691 311 692 315
rect 726 315 727 319
rect 731 315 732 319
rect 736 316 738 325
rect 774 319 780 320
rect 726 314 732 315
rect 734 315 740 316
rect 686 310 692 311
rect 728 288 730 314
rect 734 311 735 315
rect 739 311 740 315
rect 774 315 775 319
rect 779 315 780 319
rect 784 316 786 325
rect 794 319 800 320
rect 774 314 780 315
rect 782 315 788 316
rect 734 310 740 311
rect 776 288 778 314
rect 782 311 783 315
rect 787 311 788 315
rect 794 315 795 319
rect 799 315 800 319
rect 840 316 842 325
rect 908 320 910 374
rect 918 353 924 354
rect 918 349 919 353
rect 923 349 924 353
rect 918 348 924 349
rect 974 353 980 354
rect 974 349 975 353
rect 979 349 980 353
rect 974 348 980 349
rect 1030 353 1036 354
rect 1030 349 1031 353
rect 1035 349 1036 353
rect 1030 348 1036 349
rect 1056 348 1058 430
rect 1280 425 1282 457
rect 1304 448 1306 457
rect 1344 448 1346 457
rect 1358 455 1364 456
rect 1358 451 1359 455
rect 1363 451 1364 455
rect 1358 450 1364 451
rect 1302 447 1308 448
rect 1302 443 1303 447
rect 1307 443 1308 447
rect 1302 442 1308 443
rect 1342 447 1348 448
rect 1342 443 1343 447
rect 1347 443 1348 447
rect 1342 442 1348 443
rect 1278 424 1284 425
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1278 420 1279 424
rect 1283 420 1284 424
rect 1360 420 1362 450
rect 1384 448 1386 457
rect 1398 455 1404 456
rect 1398 451 1399 455
rect 1403 451 1404 455
rect 1398 450 1404 451
rect 1438 451 1444 452
rect 1382 447 1388 448
rect 1382 443 1383 447
rect 1387 443 1388 447
rect 1382 442 1388 443
rect 1400 420 1402 450
rect 1438 447 1439 451
rect 1443 447 1444 451
rect 1448 448 1450 457
rect 1526 451 1532 452
rect 1438 446 1444 447
rect 1446 447 1452 448
rect 1440 420 1442 446
rect 1446 443 1447 447
rect 1451 443 1452 447
rect 1526 447 1527 451
rect 1531 447 1532 451
rect 1536 448 1538 457
rect 1606 451 1612 452
rect 1526 446 1532 447
rect 1534 447 1540 448
rect 1446 442 1452 443
rect 1528 420 1530 446
rect 1534 443 1535 447
rect 1539 443 1540 447
rect 1606 447 1607 451
rect 1611 447 1612 451
rect 1632 448 1634 457
rect 1726 451 1732 452
rect 1606 446 1612 447
rect 1630 447 1636 448
rect 1534 442 1540 443
rect 1608 420 1610 446
rect 1630 443 1631 447
rect 1635 443 1636 447
rect 1726 447 1727 451
rect 1731 447 1732 451
rect 1736 448 1738 457
rect 1760 452 1762 490
rect 1782 477 1788 478
rect 1782 473 1783 477
rect 1787 473 1788 477
rect 1782 472 1788 473
rect 1862 477 1868 478
rect 1862 473 1863 477
rect 1867 473 1868 477
rect 1862 472 1868 473
rect 1880 472 1882 498
rect 1942 477 1948 478
rect 1942 473 1943 477
rect 1947 473 1948 477
rect 1942 472 1948 473
rect 1952 472 1954 498
rect 2022 477 2028 478
rect 2022 473 2023 477
rect 2027 473 2028 477
rect 2022 472 2028 473
rect 1784 463 1786 472
rect 1854 471 1860 472
rect 1854 467 1855 471
rect 1859 467 1860 471
rect 1854 466 1860 467
rect 1783 462 1787 463
rect 1783 457 1787 458
rect 1831 462 1835 463
rect 1831 457 1835 458
rect 1758 451 1764 452
rect 1726 446 1732 447
rect 1734 447 1740 448
rect 1630 442 1636 443
rect 1728 420 1730 446
rect 1734 443 1735 447
rect 1739 443 1740 447
rect 1758 447 1759 451
rect 1763 447 1764 451
rect 1832 448 1834 457
rect 1758 446 1764 447
rect 1830 447 1836 448
rect 1734 442 1740 443
rect 1830 443 1831 447
rect 1835 443 1836 447
rect 1830 442 1836 443
rect 1856 420 1858 466
rect 1864 463 1866 472
rect 1878 471 1884 472
rect 1878 467 1879 471
rect 1883 467 1884 471
rect 1878 466 1884 467
rect 1944 463 1946 472
rect 1950 471 1956 472
rect 1950 467 1951 471
rect 1955 467 1956 471
rect 1950 466 1956 467
rect 2024 463 2026 472
rect 1863 462 1867 463
rect 1863 457 1867 458
rect 1919 462 1923 463
rect 1919 457 1923 458
rect 1943 462 1947 463
rect 1943 457 1947 458
rect 1999 462 2003 463
rect 1999 457 2003 458
rect 2023 462 2027 463
rect 2023 457 2027 458
rect 1910 451 1916 452
rect 1910 447 1911 451
rect 1915 447 1916 451
rect 1920 448 1922 457
rect 1978 451 1984 452
rect 1910 446 1916 447
rect 1918 447 1924 448
rect 1278 419 1284 420
rect 1350 419 1356 420
rect 1238 418 1244 419
rect 1240 407 1242 418
rect 1350 415 1351 419
rect 1355 415 1356 419
rect 1350 414 1356 415
rect 1358 419 1364 420
rect 1358 415 1359 419
rect 1363 415 1364 419
rect 1358 414 1364 415
rect 1398 419 1404 420
rect 1398 415 1399 419
rect 1403 415 1404 419
rect 1398 414 1404 415
rect 1438 419 1444 420
rect 1438 415 1439 419
rect 1443 415 1444 419
rect 1438 414 1444 415
rect 1526 419 1532 420
rect 1526 415 1527 419
rect 1531 415 1532 419
rect 1526 414 1532 415
rect 1606 419 1612 420
rect 1606 415 1607 419
rect 1611 415 1612 419
rect 1606 414 1612 415
rect 1726 419 1732 420
rect 1726 415 1727 419
rect 1731 415 1732 419
rect 1726 414 1732 415
rect 1854 419 1860 420
rect 1854 415 1855 419
rect 1859 415 1860 419
rect 1854 414 1860 415
rect 1278 407 1284 408
rect 1239 406 1243 407
rect 1278 403 1279 407
rect 1283 403 1284 407
rect 1278 402 1284 403
rect 1239 401 1243 402
rect 1240 394 1242 401
rect 1280 395 1282 402
rect 1302 400 1308 401
rect 1302 396 1303 400
rect 1307 396 1308 400
rect 1302 395 1308 396
rect 1342 400 1348 401
rect 1342 396 1343 400
rect 1347 396 1348 400
rect 1342 395 1348 396
rect 1279 394 1283 395
rect 1238 393 1244 394
rect 1238 389 1239 393
rect 1243 389 1244 393
rect 1279 389 1283 390
rect 1303 394 1307 395
rect 1303 389 1307 390
rect 1343 394 1347 395
rect 1343 389 1347 390
rect 1238 388 1244 389
rect 1280 382 1282 389
rect 1278 381 1284 382
rect 1278 377 1279 381
rect 1283 377 1284 381
rect 1238 376 1244 377
rect 1278 376 1284 377
rect 1238 372 1239 376
rect 1243 372 1244 376
rect 1238 371 1244 372
rect 920 331 922 348
rect 976 331 978 348
rect 1032 331 1034 348
rect 1054 347 1060 348
rect 1054 343 1055 347
rect 1059 343 1060 347
rect 1054 342 1060 343
rect 1240 331 1242 371
rect 1278 364 1284 365
rect 1278 360 1279 364
rect 1283 360 1284 364
rect 1278 359 1284 360
rect 919 330 923 331
rect 919 325 923 326
rect 975 330 979 331
rect 975 325 979 326
rect 1031 330 1035 331
rect 1031 325 1035 326
rect 1239 330 1243 331
rect 1239 325 1243 326
rect 906 319 912 320
rect 794 314 800 315
rect 838 315 844 316
rect 782 310 788 311
rect 250 287 256 288
rect 250 286 251 287
rect 244 284 251 286
rect 230 282 236 283
rect 250 283 251 284
rect 255 283 256 287
rect 250 282 256 283
rect 382 287 388 288
rect 382 283 383 287
rect 387 283 388 287
rect 382 282 388 283
rect 438 287 444 288
rect 438 283 439 287
rect 443 283 444 287
rect 438 282 444 283
rect 534 287 540 288
rect 534 283 535 287
rect 539 283 540 287
rect 534 282 540 283
rect 630 287 636 288
rect 630 283 631 287
rect 635 283 636 287
rect 630 282 636 283
rect 654 287 660 288
rect 654 283 655 287
rect 659 283 660 287
rect 654 282 660 283
rect 678 287 684 288
rect 678 283 679 287
rect 683 283 684 287
rect 678 282 684 283
rect 726 287 732 288
rect 726 283 727 287
rect 731 283 732 287
rect 726 282 732 283
rect 774 287 780 288
rect 774 283 775 287
rect 779 283 780 287
rect 774 282 780 283
rect 670 279 676 280
rect 670 275 671 279
rect 675 275 676 279
rect 670 274 676 275
rect 174 268 180 269
rect 174 264 175 268
rect 179 264 180 268
rect 174 263 180 264
rect 214 268 220 269
rect 214 264 215 268
rect 219 264 220 268
rect 214 263 220 264
rect 254 268 260 269
rect 254 264 255 268
rect 259 264 260 268
rect 254 263 260 264
rect 294 268 300 269
rect 294 264 295 268
rect 299 264 300 268
rect 294 263 300 264
rect 334 268 340 269
rect 334 264 335 268
rect 339 264 340 268
rect 334 263 340 264
rect 390 268 396 269
rect 390 264 391 268
rect 395 264 396 268
rect 390 263 396 264
rect 446 268 452 269
rect 446 264 447 268
rect 451 264 452 268
rect 446 263 452 264
rect 494 268 500 269
rect 494 264 495 268
rect 499 264 500 268
rect 494 263 500 264
rect 542 268 548 269
rect 542 264 543 268
rect 547 264 548 268
rect 542 263 548 264
rect 590 268 596 269
rect 590 264 591 268
rect 595 264 596 268
rect 590 263 596 264
rect 638 268 644 269
rect 638 264 639 268
rect 643 264 644 268
rect 638 263 644 264
rect 176 255 178 263
rect 216 255 218 263
rect 256 255 258 263
rect 296 255 298 263
rect 336 255 338 263
rect 392 255 394 263
rect 448 255 450 263
rect 496 255 498 263
rect 544 255 546 263
rect 592 255 594 263
rect 640 255 642 263
rect 175 254 179 255
rect 175 249 179 250
rect 215 254 219 255
rect 215 249 219 250
rect 223 254 227 255
rect 223 249 227 250
rect 255 254 259 255
rect 255 249 259 250
rect 295 254 299 255
rect 295 249 299 250
rect 311 254 315 255
rect 311 249 315 250
rect 335 254 339 255
rect 335 249 339 250
rect 391 254 395 255
rect 391 249 395 250
rect 447 254 451 255
rect 447 249 451 250
rect 463 254 467 255
rect 463 249 467 250
rect 495 254 499 255
rect 495 249 499 250
rect 527 254 531 255
rect 527 249 531 250
rect 543 254 547 255
rect 543 249 547 250
rect 591 254 595 255
rect 591 249 595 250
rect 639 254 643 255
rect 639 249 643 250
rect 647 254 651 255
rect 647 249 651 250
rect 222 248 228 249
rect 222 244 223 248
rect 227 244 228 248
rect 222 243 228 244
rect 310 248 316 249
rect 310 244 311 248
rect 315 244 316 248
rect 310 243 316 244
rect 390 248 396 249
rect 390 244 391 248
rect 395 244 396 248
rect 390 243 396 244
rect 462 248 468 249
rect 462 244 463 248
rect 467 244 468 248
rect 462 243 468 244
rect 526 248 532 249
rect 526 244 527 248
rect 531 244 532 248
rect 526 243 532 244
rect 590 248 596 249
rect 590 244 591 248
rect 595 244 596 248
rect 590 243 596 244
rect 646 248 652 249
rect 646 244 647 248
rect 651 244 652 248
rect 646 243 652 244
rect 158 227 164 228
rect 158 223 159 227
rect 163 223 164 227
rect 158 222 164 223
rect 286 227 292 228
rect 286 223 287 227
rect 291 223 292 227
rect 286 222 292 223
rect 222 201 228 202
rect 222 197 223 201
rect 227 197 228 201
rect 222 196 228 197
rect 288 196 290 222
rect 614 219 620 220
rect 614 215 615 219
rect 619 215 620 219
rect 614 214 620 215
rect 310 201 316 202
rect 310 197 311 201
rect 315 197 316 201
rect 310 196 316 197
rect 390 201 396 202
rect 390 197 391 201
rect 395 197 396 201
rect 390 196 396 197
rect 462 201 468 202
rect 462 197 463 201
rect 467 197 468 201
rect 462 196 468 197
rect 526 201 532 202
rect 526 197 527 201
rect 531 197 532 201
rect 526 196 532 197
rect 590 201 596 202
rect 590 197 591 201
rect 595 197 596 201
rect 590 196 596 197
rect 136 155 138 196
rect 150 195 156 196
rect 150 191 151 195
rect 155 191 156 195
rect 150 190 156 191
rect 224 155 226 196
rect 286 195 292 196
rect 286 191 287 195
rect 291 191 292 195
rect 286 190 292 191
rect 312 155 314 196
rect 392 155 394 196
rect 464 155 466 196
rect 528 155 530 196
rect 592 155 594 196
rect 111 154 115 155
rect 111 149 115 150
rect 135 154 139 155
rect 135 149 139 150
rect 151 154 155 155
rect 151 149 155 150
rect 191 154 195 155
rect 191 149 195 150
rect 223 154 227 155
rect 223 149 227 150
rect 231 154 235 155
rect 231 149 235 150
rect 271 154 275 155
rect 271 149 275 150
rect 311 154 315 155
rect 311 149 315 150
rect 351 154 355 155
rect 351 149 355 150
rect 391 154 395 155
rect 391 149 395 150
rect 431 154 435 155
rect 431 149 435 150
rect 463 154 467 155
rect 463 149 467 150
rect 471 154 475 155
rect 471 149 475 150
rect 511 154 515 155
rect 511 149 515 150
rect 527 154 531 155
rect 527 149 531 150
rect 551 154 555 155
rect 551 149 555 150
rect 591 154 595 155
rect 591 149 595 150
rect 112 117 114 149
rect 152 140 154 149
rect 178 143 184 144
rect 150 139 156 140
rect 150 135 151 139
rect 155 135 156 139
rect 178 139 179 143
rect 183 139 184 143
rect 192 140 194 149
rect 218 143 224 144
rect 178 138 184 139
rect 190 139 196 140
rect 150 134 156 135
rect 110 116 116 117
rect 110 112 111 116
rect 115 112 116 116
rect 180 112 182 138
rect 190 135 191 139
rect 195 135 196 139
rect 218 139 219 143
rect 223 139 224 143
rect 232 140 234 149
rect 258 143 264 144
rect 218 138 224 139
rect 230 139 236 140
rect 190 134 196 135
rect 110 111 116 112
rect 178 111 184 112
rect 178 107 179 111
rect 183 107 184 111
rect 220 110 222 138
rect 230 135 231 139
rect 235 135 236 139
rect 258 139 259 143
rect 263 139 264 143
rect 272 140 274 149
rect 298 143 304 144
rect 258 138 264 139
rect 270 139 276 140
rect 230 134 236 135
rect 226 111 232 112
rect 226 110 227 111
rect 220 108 227 110
rect 178 106 184 107
rect 226 107 227 108
rect 231 107 232 111
rect 260 110 262 138
rect 270 135 271 139
rect 275 135 276 139
rect 298 139 299 143
rect 303 139 304 143
rect 312 140 314 149
rect 338 143 344 144
rect 298 138 304 139
rect 310 139 316 140
rect 270 134 276 135
rect 300 120 302 138
rect 310 135 311 139
rect 315 135 316 139
rect 338 139 339 143
rect 343 139 344 143
rect 352 140 354 149
rect 378 143 384 144
rect 338 138 344 139
rect 350 139 356 140
rect 310 134 316 135
rect 298 119 304 120
rect 298 115 299 119
rect 303 115 304 119
rect 298 114 304 115
rect 266 111 272 112
rect 266 110 267 111
rect 260 108 267 110
rect 226 106 232 107
rect 266 107 267 108
rect 271 107 272 111
rect 340 110 342 138
rect 350 135 351 139
rect 355 135 356 139
rect 378 139 379 143
rect 383 139 384 143
rect 392 140 394 149
rect 432 140 434 149
rect 446 147 452 148
rect 446 143 447 147
rect 451 143 452 147
rect 446 142 452 143
rect 458 143 464 144
rect 378 138 384 139
rect 390 139 396 140
rect 350 134 356 135
rect 346 111 352 112
rect 346 110 347 111
rect 340 108 347 110
rect 266 106 272 107
rect 346 107 347 108
rect 351 107 352 111
rect 380 110 382 138
rect 390 135 391 139
rect 395 135 396 139
rect 390 134 396 135
rect 430 139 436 140
rect 430 135 431 139
rect 435 135 436 139
rect 430 134 436 135
rect 448 112 450 142
rect 458 139 459 143
rect 463 139 464 143
rect 472 140 474 149
rect 498 143 504 144
rect 458 138 464 139
rect 470 139 476 140
rect 386 111 392 112
rect 386 110 387 111
rect 380 108 387 110
rect 346 106 352 107
rect 386 107 387 108
rect 391 107 392 111
rect 386 106 392 107
rect 446 111 452 112
rect 446 107 447 111
rect 451 107 452 111
rect 460 110 462 138
rect 470 135 471 139
rect 475 135 476 139
rect 498 139 499 143
rect 503 139 504 143
rect 512 140 514 149
rect 538 143 544 144
rect 498 138 504 139
rect 510 139 516 140
rect 470 134 476 135
rect 466 111 472 112
rect 466 110 467 111
rect 460 108 467 110
rect 446 106 452 107
rect 466 107 467 108
rect 471 107 472 111
rect 500 110 502 138
rect 510 135 511 139
rect 515 135 516 139
rect 538 139 539 143
rect 543 139 544 143
rect 552 140 554 149
rect 578 143 584 144
rect 538 138 544 139
rect 550 139 556 140
rect 510 134 516 135
rect 506 111 512 112
rect 506 110 507 111
rect 500 108 507 110
rect 466 106 472 107
rect 506 107 507 108
rect 511 107 512 111
rect 540 110 542 138
rect 550 135 551 139
rect 555 135 556 139
rect 578 139 579 143
rect 583 139 584 143
rect 592 140 594 149
rect 616 144 618 214
rect 646 201 652 202
rect 646 197 647 201
rect 651 197 652 201
rect 646 196 652 197
rect 672 196 674 274
rect 686 268 692 269
rect 686 264 687 268
rect 691 264 692 268
rect 686 263 692 264
rect 734 268 740 269
rect 734 264 735 268
rect 739 264 740 268
rect 734 263 740 264
rect 782 268 788 269
rect 782 264 783 268
rect 787 264 788 268
rect 782 263 788 264
rect 688 255 690 263
rect 736 255 738 263
rect 784 255 786 263
rect 687 254 691 255
rect 687 249 691 250
rect 695 254 699 255
rect 695 249 699 250
rect 735 254 739 255
rect 735 249 739 250
rect 783 254 787 255
rect 783 249 787 250
rect 694 248 700 249
rect 694 244 695 248
rect 699 244 700 248
rect 694 243 700 244
rect 734 248 740 249
rect 734 244 735 248
rect 739 244 740 248
rect 734 243 740 244
rect 782 248 788 249
rect 782 244 783 248
rect 787 244 788 248
rect 782 243 788 244
rect 796 236 798 314
rect 838 311 839 315
rect 843 311 844 315
rect 906 315 907 319
rect 911 315 912 319
rect 906 314 912 315
rect 838 310 844 311
rect 862 307 868 308
rect 862 303 863 307
rect 867 303 868 307
rect 862 302 868 303
rect 864 288 866 302
rect 1240 293 1242 325
rect 1280 319 1282 359
rect 1352 336 1354 414
rect 1382 400 1388 401
rect 1382 396 1383 400
rect 1387 396 1388 400
rect 1382 395 1388 396
rect 1446 400 1452 401
rect 1446 396 1447 400
rect 1451 396 1452 400
rect 1446 395 1452 396
rect 1534 400 1540 401
rect 1534 396 1535 400
rect 1539 396 1540 400
rect 1534 395 1540 396
rect 1630 400 1636 401
rect 1630 396 1631 400
rect 1635 396 1636 400
rect 1630 395 1636 396
rect 1734 400 1740 401
rect 1734 396 1735 400
rect 1739 396 1740 400
rect 1734 395 1740 396
rect 1830 400 1836 401
rect 1830 396 1831 400
rect 1835 396 1836 400
rect 1830 395 1836 396
rect 1359 394 1363 395
rect 1359 389 1363 390
rect 1383 394 1387 395
rect 1383 389 1387 390
rect 1399 394 1403 395
rect 1399 389 1403 390
rect 1439 394 1443 395
rect 1439 389 1443 390
rect 1447 394 1451 395
rect 1447 389 1451 390
rect 1487 394 1491 395
rect 1487 389 1491 390
rect 1535 394 1539 395
rect 1535 389 1539 390
rect 1543 394 1547 395
rect 1543 389 1547 390
rect 1607 394 1611 395
rect 1607 389 1611 390
rect 1631 394 1635 395
rect 1631 389 1635 390
rect 1679 394 1683 395
rect 1679 389 1683 390
rect 1735 394 1739 395
rect 1735 389 1739 390
rect 1759 394 1763 395
rect 1759 389 1763 390
rect 1831 394 1835 395
rect 1831 389 1835 390
rect 1839 394 1843 395
rect 1839 389 1843 390
rect 1358 388 1364 389
rect 1358 384 1359 388
rect 1363 384 1364 388
rect 1358 383 1364 384
rect 1398 388 1404 389
rect 1398 384 1399 388
rect 1403 384 1404 388
rect 1398 383 1404 384
rect 1438 388 1444 389
rect 1438 384 1439 388
rect 1443 384 1444 388
rect 1438 383 1444 384
rect 1486 388 1492 389
rect 1486 384 1487 388
rect 1491 384 1492 388
rect 1486 383 1492 384
rect 1542 388 1548 389
rect 1542 384 1543 388
rect 1547 384 1548 388
rect 1542 383 1548 384
rect 1606 388 1612 389
rect 1606 384 1607 388
rect 1611 384 1612 388
rect 1606 383 1612 384
rect 1678 388 1684 389
rect 1678 384 1679 388
rect 1683 384 1684 388
rect 1678 383 1684 384
rect 1758 388 1764 389
rect 1758 384 1759 388
rect 1763 384 1764 388
rect 1758 383 1764 384
rect 1838 388 1844 389
rect 1838 384 1839 388
rect 1843 384 1844 388
rect 1838 383 1844 384
rect 1912 368 1914 446
rect 1918 443 1919 447
rect 1923 443 1924 447
rect 1978 447 1979 451
rect 1983 447 1984 451
rect 2000 448 2002 457
rect 2040 456 2042 498
rect 2102 477 2108 478
rect 2102 473 2103 477
rect 2107 473 2108 477
rect 2102 472 2108 473
rect 2124 472 2126 550
rect 2166 536 2172 537
rect 2166 532 2167 536
rect 2171 532 2172 536
rect 2166 531 2172 532
rect 2238 536 2244 537
rect 2238 532 2239 536
rect 2243 532 2244 536
rect 2238 531 2244 532
rect 2167 530 2171 531
rect 2167 525 2171 526
rect 2191 530 2195 531
rect 2191 525 2195 526
rect 2239 530 2243 531
rect 2239 525 2243 526
rect 2287 530 2291 531
rect 2287 525 2291 526
rect 2190 524 2196 525
rect 2190 520 2191 524
rect 2195 520 2196 524
rect 2190 519 2196 520
rect 2286 524 2292 525
rect 2286 520 2287 524
rect 2291 520 2292 524
rect 2286 519 2292 520
rect 2304 504 2306 582
rect 2310 579 2311 583
rect 2315 579 2316 583
rect 2350 583 2351 587
rect 2355 583 2356 587
rect 2360 584 2362 593
rect 2350 582 2356 583
rect 2358 583 2364 584
rect 2310 578 2316 579
rect 2352 556 2354 582
rect 2358 579 2359 583
rect 2363 579 2364 583
rect 2358 578 2364 579
rect 2408 561 2410 593
rect 2406 560 2412 561
rect 2406 556 2407 560
rect 2411 556 2412 560
rect 2338 555 2344 556
rect 2338 551 2339 555
rect 2343 551 2344 555
rect 2338 550 2344 551
rect 2350 555 2356 556
rect 2406 555 2412 556
rect 2350 551 2351 555
rect 2355 551 2356 555
rect 2350 550 2356 551
rect 2310 536 2316 537
rect 2310 532 2311 536
rect 2315 532 2316 536
rect 2310 531 2316 532
rect 2311 530 2315 531
rect 2311 525 2315 526
rect 2294 503 2300 504
rect 2294 499 2295 503
rect 2299 499 2300 503
rect 2294 498 2300 499
rect 2302 503 2308 504
rect 2302 499 2303 503
rect 2307 499 2308 503
rect 2302 498 2308 499
rect 2190 477 2196 478
rect 2190 473 2191 477
rect 2195 473 2196 477
rect 2190 472 2196 473
rect 2286 477 2292 478
rect 2286 473 2287 477
rect 2291 473 2292 477
rect 2286 472 2292 473
rect 2296 472 2298 498
rect 2340 472 2342 550
rect 2406 543 2412 544
rect 2406 539 2407 543
rect 2411 539 2412 543
rect 2406 538 2412 539
rect 2358 536 2364 537
rect 2358 532 2359 536
rect 2363 532 2364 536
rect 2358 531 2364 532
rect 2408 531 2410 538
rect 2359 530 2363 531
rect 2359 525 2363 526
rect 2407 530 2411 531
rect 2407 525 2411 526
rect 2358 524 2364 525
rect 2358 520 2359 524
rect 2363 520 2364 524
rect 2358 519 2364 520
rect 2408 518 2410 525
rect 2406 517 2412 518
rect 2406 513 2407 517
rect 2411 513 2412 517
rect 2406 512 2412 513
rect 2382 503 2388 504
rect 2382 499 2383 503
rect 2387 499 2388 503
rect 2382 498 2388 499
rect 2406 500 2412 501
rect 2358 477 2364 478
rect 2358 473 2359 477
rect 2363 473 2364 477
rect 2358 472 2364 473
rect 2104 463 2106 472
rect 2122 471 2128 472
rect 2122 467 2123 471
rect 2127 467 2128 471
rect 2122 466 2128 467
rect 2110 463 2116 464
rect 2192 463 2194 472
rect 2288 463 2290 472
rect 2294 471 2300 472
rect 2294 467 2295 471
rect 2299 467 2300 471
rect 2294 466 2300 467
rect 2338 471 2344 472
rect 2338 467 2339 471
rect 2343 467 2344 471
rect 2338 466 2344 467
rect 2360 463 2362 472
rect 2071 462 2075 463
rect 2071 457 2075 458
rect 2103 462 2107 463
rect 2110 459 2111 463
rect 2115 459 2116 463
rect 2110 458 2116 459
rect 2135 462 2139 463
rect 2103 457 2107 458
rect 2038 455 2044 456
rect 2038 451 2039 455
rect 2043 451 2044 455
rect 2038 450 2044 451
rect 2072 448 2074 457
rect 1978 446 1984 447
rect 1998 447 2004 448
rect 1918 442 1924 443
rect 1980 420 1982 446
rect 1998 443 1999 447
rect 2003 443 2004 447
rect 1998 442 2004 443
rect 2070 447 2076 448
rect 2070 443 2071 447
rect 2075 443 2076 447
rect 2070 442 2076 443
rect 2112 420 2114 458
rect 2135 457 2139 458
rect 2191 462 2195 463
rect 2191 457 2195 458
rect 2199 462 2203 463
rect 2199 457 2203 458
rect 2255 462 2259 463
rect 2255 457 2259 458
rect 2287 462 2291 463
rect 2287 457 2291 458
rect 2319 462 2323 463
rect 2319 457 2323 458
rect 2359 462 2363 463
rect 2359 457 2363 458
rect 2126 451 2132 452
rect 2126 447 2127 451
rect 2131 447 2132 451
rect 2136 448 2138 457
rect 2190 451 2196 452
rect 2126 446 2132 447
rect 2134 447 2140 448
rect 2128 420 2130 446
rect 2134 443 2135 447
rect 2139 443 2140 447
rect 2190 447 2191 451
rect 2195 447 2196 451
rect 2200 448 2202 457
rect 2246 451 2252 452
rect 2190 446 2196 447
rect 2198 447 2204 448
rect 2134 442 2140 443
rect 2192 420 2194 446
rect 2198 443 2199 447
rect 2203 443 2204 447
rect 2246 447 2247 451
rect 2251 447 2252 451
rect 2256 448 2258 457
rect 2310 451 2316 452
rect 2246 446 2252 447
rect 2254 447 2260 448
rect 2198 442 2204 443
rect 2248 420 2250 446
rect 2254 443 2255 447
rect 2259 443 2260 447
rect 2310 447 2311 451
rect 2315 447 2316 451
rect 2320 448 2322 457
rect 2346 451 2352 452
rect 2310 446 2316 447
rect 2318 447 2324 448
rect 2254 442 2260 443
rect 1978 419 1984 420
rect 1978 415 1979 419
rect 1983 415 1984 419
rect 1978 414 1984 415
rect 2110 419 2116 420
rect 2110 415 2111 419
rect 2115 415 2116 419
rect 2110 414 2116 415
rect 2126 419 2132 420
rect 2126 415 2127 419
rect 2131 415 2132 419
rect 2126 414 2132 415
rect 2190 419 2196 420
rect 2190 415 2191 419
rect 2195 415 2196 419
rect 2190 414 2196 415
rect 2246 419 2252 420
rect 2246 415 2247 419
rect 2251 415 2252 419
rect 2246 414 2252 415
rect 2098 411 2104 412
rect 2098 407 2099 411
rect 2103 407 2104 411
rect 2098 406 2104 407
rect 1918 400 1924 401
rect 1918 396 1919 400
rect 1923 396 1924 400
rect 1918 395 1924 396
rect 1998 400 2004 401
rect 1998 396 1999 400
rect 2003 396 2004 400
rect 1998 395 2004 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 1919 394 1923 395
rect 1919 389 1923 390
rect 1999 394 2003 395
rect 1999 389 2003 390
rect 2071 394 2075 395
rect 2071 389 2075 390
rect 2079 394 2083 395
rect 2079 389 2083 390
rect 1918 388 1924 389
rect 1918 384 1919 388
rect 1923 384 1924 388
rect 1918 383 1924 384
rect 1998 388 2004 389
rect 1998 384 1999 388
rect 2003 384 2004 388
rect 1998 383 2004 384
rect 2078 388 2084 389
rect 2078 384 2079 388
rect 2083 384 2084 388
rect 2078 383 2084 384
rect 1414 367 1420 368
rect 1414 363 1415 367
rect 1419 363 1420 367
rect 1414 362 1420 363
rect 1454 367 1460 368
rect 1454 363 1455 367
rect 1459 363 1460 367
rect 1454 362 1460 363
rect 1502 367 1508 368
rect 1502 363 1503 367
rect 1507 363 1508 367
rect 1502 362 1508 363
rect 1558 367 1564 368
rect 1558 363 1559 367
rect 1563 363 1564 367
rect 1558 362 1564 363
rect 1614 367 1620 368
rect 1614 363 1615 367
rect 1619 363 1620 367
rect 1614 362 1620 363
rect 1854 367 1860 368
rect 1854 363 1855 367
rect 1859 363 1860 367
rect 1854 362 1860 363
rect 1910 367 1916 368
rect 1910 363 1911 367
rect 1915 363 1916 367
rect 1910 362 1916 363
rect 1358 341 1364 342
rect 1358 337 1359 341
rect 1363 337 1364 341
rect 1358 336 1364 337
rect 1398 341 1404 342
rect 1398 337 1399 341
rect 1403 337 1404 341
rect 1398 336 1404 337
rect 1416 336 1418 362
rect 1438 341 1444 342
rect 1438 337 1439 341
rect 1443 337 1444 341
rect 1438 336 1444 337
rect 1456 336 1458 362
rect 1486 341 1492 342
rect 1486 337 1487 341
rect 1491 337 1492 341
rect 1486 336 1492 337
rect 1504 336 1506 362
rect 1542 341 1548 342
rect 1542 337 1543 341
rect 1547 337 1548 341
rect 1542 336 1548 337
rect 1560 336 1562 362
rect 1606 341 1612 342
rect 1606 337 1607 341
rect 1611 337 1612 341
rect 1606 336 1612 337
rect 1350 335 1356 336
rect 1350 331 1351 335
rect 1355 331 1356 335
rect 1350 330 1356 331
rect 1360 319 1362 336
rect 1400 319 1402 336
rect 1414 335 1420 336
rect 1414 331 1415 335
rect 1419 331 1420 335
rect 1414 330 1420 331
rect 1440 319 1442 336
rect 1454 335 1460 336
rect 1454 331 1455 335
rect 1459 331 1460 335
rect 1454 330 1460 331
rect 1488 319 1490 336
rect 1502 335 1508 336
rect 1502 331 1503 335
rect 1507 331 1508 335
rect 1502 330 1508 331
rect 1544 319 1546 336
rect 1558 335 1564 336
rect 1558 331 1559 335
rect 1563 331 1564 335
rect 1558 330 1564 331
rect 1608 319 1610 336
rect 1279 318 1283 319
rect 1279 313 1283 314
rect 1359 318 1363 319
rect 1359 313 1363 314
rect 1399 318 1403 319
rect 1399 313 1403 314
rect 1439 318 1443 319
rect 1439 313 1443 314
rect 1487 318 1491 319
rect 1487 313 1491 314
rect 1511 318 1515 319
rect 1511 313 1515 314
rect 1543 318 1547 319
rect 1543 313 1547 314
rect 1551 318 1555 319
rect 1551 313 1555 314
rect 1591 318 1595 319
rect 1591 313 1595 314
rect 1607 318 1611 319
rect 1607 313 1611 314
rect 1238 292 1244 293
rect 1238 288 1239 292
rect 1243 288 1244 292
rect 862 287 868 288
rect 1238 287 1244 288
rect 862 283 863 287
rect 867 283 868 287
rect 862 282 868 283
rect 1280 281 1282 313
rect 1512 304 1514 313
rect 1538 307 1544 308
rect 1510 303 1516 304
rect 1510 299 1511 303
rect 1515 299 1516 303
rect 1538 303 1539 307
rect 1543 303 1544 307
rect 1552 304 1554 313
rect 1592 304 1594 313
rect 1598 311 1604 312
rect 1598 307 1599 311
rect 1603 307 1604 311
rect 1616 308 1618 362
rect 1702 359 1708 360
rect 1702 355 1703 359
rect 1707 355 1708 359
rect 1702 354 1708 355
rect 1678 341 1684 342
rect 1678 337 1679 341
rect 1683 337 1684 341
rect 1678 336 1684 337
rect 1704 336 1706 354
rect 1758 341 1764 342
rect 1758 337 1759 341
rect 1763 337 1764 341
rect 1758 336 1764 337
rect 1838 341 1844 342
rect 1838 337 1839 341
rect 1843 337 1844 341
rect 1838 336 1844 337
rect 1856 336 1858 362
rect 2022 359 2028 360
rect 2022 355 2023 359
rect 2027 355 2028 359
rect 2022 354 2028 355
rect 1918 341 1924 342
rect 1918 337 1919 341
rect 1923 337 1924 341
rect 1918 336 1924 337
rect 1998 341 2004 342
rect 1998 337 1999 341
rect 2003 337 2004 341
rect 1998 336 2004 337
rect 2024 336 2026 354
rect 2078 341 2084 342
rect 2078 337 2079 341
rect 2083 337 2084 341
rect 2078 336 2084 337
rect 2100 336 2102 406
rect 2134 400 2140 401
rect 2134 396 2135 400
rect 2139 396 2140 400
rect 2134 395 2140 396
rect 2198 400 2204 401
rect 2198 396 2199 400
rect 2203 396 2204 400
rect 2198 395 2204 396
rect 2254 400 2260 401
rect 2254 396 2255 400
rect 2259 396 2260 400
rect 2254 395 2260 396
rect 2135 394 2139 395
rect 2135 389 2139 390
rect 2159 394 2163 395
rect 2159 389 2163 390
rect 2199 394 2203 395
rect 2199 389 2203 390
rect 2247 394 2251 395
rect 2247 389 2251 390
rect 2255 394 2259 395
rect 2255 389 2259 390
rect 2158 388 2164 389
rect 2158 384 2159 388
rect 2163 384 2164 388
rect 2158 383 2164 384
rect 2246 388 2252 389
rect 2246 384 2247 388
rect 2251 384 2252 388
rect 2246 383 2252 384
rect 2312 368 2314 446
rect 2318 443 2319 447
rect 2323 443 2324 447
rect 2346 447 2347 451
rect 2351 447 2352 451
rect 2360 448 2362 457
rect 2384 452 2386 498
rect 2406 496 2407 500
rect 2411 496 2412 500
rect 2406 495 2412 496
rect 2408 463 2410 495
rect 2407 462 2411 463
rect 2407 457 2411 458
rect 2382 451 2388 452
rect 2346 446 2352 447
rect 2358 447 2364 448
rect 2318 442 2324 443
rect 2348 428 2350 446
rect 2358 443 2359 447
rect 2363 443 2364 447
rect 2382 447 2383 451
rect 2387 447 2388 451
rect 2382 446 2388 447
rect 2358 442 2364 443
rect 2346 427 2352 428
rect 2346 423 2347 427
rect 2351 423 2352 427
rect 2408 425 2410 457
rect 2346 422 2352 423
rect 2406 424 2412 425
rect 2406 420 2407 424
rect 2411 420 2412 424
rect 2346 419 2352 420
rect 2406 419 2412 420
rect 2346 415 2347 419
rect 2351 415 2352 419
rect 2346 414 2352 415
rect 2318 400 2324 401
rect 2318 396 2319 400
rect 2323 396 2324 400
rect 2318 395 2324 396
rect 2319 394 2323 395
rect 2319 389 2323 390
rect 2335 394 2339 395
rect 2335 389 2339 390
rect 2334 388 2340 389
rect 2334 384 2335 388
rect 2339 384 2340 388
rect 2334 383 2340 384
rect 2174 367 2180 368
rect 2174 363 2175 367
rect 2179 363 2180 367
rect 2174 362 2180 363
rect 2218 367 2224 368
rect 2218 363 2219 367
rect 2223 363 2224 367
rect 2218 362 2224 363
rect 2226 367 2232 368
rect 2226 363 2227 367
rect 2231 363 2232 367
rect 2226 362 2232 363
rect 2310 367 2316 368
rect 2310 363 2311 367
rect 2315 363 2316 367
rect 2310 362 2316 363
rect 2158 341 2164 342
rect 2158 337 2159 341
rect 2163 337 2164 341
rect 2158 336 2164 337
rect 2176 336 2178 362
rect 2220 336 2222 362
rect 1680 319 1682 336
rect 1702 335 1708 336
rect 1702 331 1703 335
rect 1707 331 1708 335
rect 1702 330 1708 331
rect 1760 319 1762 336
rect 1840 319 1842 336
rect 1846 335 1852 336
rect 1846 331 1847 335
rect 1851 331 1852 335
rect 1846 330 1852 331
rect 1854 335 1860 336
rect 1854 331 1855 335
rect 1859 331 1860 335
rect 1854 330 1860 331
rect 1631 318 1635 319
rect 1631 313 1635 314
rect 1671 318 1675 319
rect 1671 313 1675 314
rect 1679 318 1683 319
rect 1679 313 1683 314
rect 1711 318 1715 319
rect 1711 313 1715 314
rect 1751 318 1755 319
rect 1751 313 1755 314
rect 1759 318 1763 319
rect 1759 313 1763 314
rect 1791 318 1795 319
rect 1791 313 1795 314
rect 1839 318 1843 319
rect 1839 313 1843 314
rect 1598 306 1604 307
rect 1614 307 1620 308
rect 1538 302 1544 303
rect 1550 303 1556 304
rect 1510 298 1516 299
rect 1540 284 1542 302
rect 1550 299 1551 303
rect 1555 299 1556 303
rect 1550 298 1556 299
rect 1590 303 1596 304
rect 1590 299 1591 303
rect 1595 299 1596 303
rect 1590 298 1596 299
rect 1538 283 1544 284
rect 1278 280 1284 281
rect 1278 276 1279 280
rect 1283 276 1284 280
rect 1538 279 1539 283
rect 1543 279 1544 283
rect 1538 278 1544 279
rect 1600 276 1602 306
rect 1614 303 1615 307
rect 1619 303 1620 307
rect 1632 304 1634 313
rect 1672 304 1674 313
rect 1686 311 1692 312
rect 1686 307 1687 311
rect 1691 307 1692 311
rect 1686 306 1692 307
rect 1698 307 1704 308
rect 1614 302 1620 303
rect 1630 303 1636 304
rect 1630 299 1631 303
rect 1635 299 1636 303
rect 1630 298 1636 299
rect 1670 303 1676 304
rect 1670 299 1671 303
rect 1675 299 1676 303
rect 1670 298 1676 299
rect 1688 276 1690 306
rect 1698 303 1699 307
rect 1703 303 1704 307
rect 1712 304 1714 313
rect 1752 304 1754 313
rect 1766 311 1772 312
rect 1766 307 1767 311
rect 1771 307 1772 311
rect 1766 306 1772 307
rect 1778 307 1784 308
rect 1698 302 1704 303
rect 1710 303 1716 304
rect 1700 284 1702 302
rect 1710 299 1711 303
rect 1715 299 1716 303
rect 1710 298 1716 299
rect 1750 303 1756 304
rect 1750 299 1751 303
rect 1755 299 1756 303
rect 1750 298 1756 299
rect 1698 283 1704 284
rect 1698 279 1699 283
rect 1703 279 1704 283
rect 1698 278 1704 279
rect 1768 276 1770 306
rect 1778 303 1779 307
rect 1783 303 1784 307
rect 1792 304 1794 313
rect 1840 304 1842 313
rect 1778 302 1784 303
rect 1790 303 1796 304
rect 1780 284 1782 302
rect 1790 299 1791 303
rect 1795 299 1796 303
rect 1790 298 1796 299
rect 1838 303 1844 304
rect 1838 299 1839 303
rect 1843 299 1844 303
rect 1838 298 1844 299
rect 1778 283 1784 284
rect 1778 279 1779 283
rect 1783 279 1784 283
rect 1778 278 1784 279
rect 1848 276 1850 330
rect 1920 319 1922 336
rect 2000 319 2002 336
rect 2022 335 2028 336
rect 2022 331 2023 335
rect 2027 331 2028 335
rect 2022 330 2028 331
rect 2080 319 2082 336
rect 2098 335 2104 336
rect 2098 331 2099 335
rect 2103 331 2104 335
rect 2098 330 2104 331
rect 2160 319 2162 336
rect 2174 335 2180 336
rect 2174 331 2175 335
rect 2179 331 2180 335
rect 2174 330 2180 331
rect 2218 335 2224 336
rect 2218 331 2219 335
rect 2223 331 2224 335
rect 2218 330 2224 331
rect 1903 318 1907 319
rect 1903 313 1907 314
rect 1919 318 1923 319
rect 1919 313 1923 314
rect 1967 318 1971 319
rect 1967 313 1971 314
rect 1999 318 2003 319
rect 1999 313 2003 314
rect 2039 318 2043 319
rect 2039 313 2043 314
rect 2079 318 2083 319
rect 2079 313 2083 314
rect 2119 318 2123 319
rect 2119 313 2123 314
rect 2159 318 2163 319
rect 2159 313 2163 314
rect 2199 318 2203 319
rect 2199 313 2203 314
rect 1894 307 1900 308
rect 1894 303 1895 307
rect 1899 303 1900 307
rect 1904 304 1906 313
rect 1958 307 1964 308
rect 1894 302 1900 303
rect 1902 303 1908 304
rect 1896 276 1898 302
rect 1902 299 1903 303
rect 1907 299 1908 303
rect 1958 303 1959 307
rect 1963 303 1964 307
rect 1968 304 1970 313
rect 2026 307 2032 308
rect 1958 302 1964 303
rect 1966 303 1972 304
rect 1902 298 1908 299
rect 1960 276 1962 302
rect 1966 299 1967 303
rect 1971 299 1972 303
rect 2026 303 2027 307
rect 2031 303 2032 307
rect 2040 304 2042 313
rect 2110 307 2116 308
rect 2026 302 2032 303
rect 2038 303 2044 304
rect 1966 298 1972 299
rect 2028 276 2030 302
rect 2038 299 2039 303
rect 2043 299 2044 303
rect 2110 303 2111 307
rect 2115 303 2116 307
rect 2120 304 2122 313
rect 2130 307 2136 308
rect 2110 302 2116 303
rect 2118 303 2124 304
rect 2038 298 2044 299
rect 2112 276 2114 302
rect 2118 299 2119 303
rect 2123 299 2124 303
rect 2130 303 2131 307
rect 2135 303 2136 307
rect 2200 304 2202 313
rect 2228 308 2230 362
rect 2246 341 2252 342
rect 2246 337 2247 341
rect 2251 337 2252 341
rect 2246 336 2252 337
rect 2334 341 2340 342
rect 2334 337 2335 341
rect 2339 337 2340 341
rect 2334 336 2340 337
rect 2348 336 2350 414
rect 2406 407 2412 408
rect 2406 403 2407 407
rect 2411 403 2412 407
rect 2406 402 2412 403
rect 2358 400 2364 401
rect 2358 396 2359 400
rect 2363 396 2364 400
rect 2358 395 2364 396
rect 2408 395 2410 402
rect 2359 394 2363 395
rect 2359 389 2363 390
rect 2407 394 2411 395
rect 2407 389 2411 390
rect 2408 382 2410 389
rect 2406 381 2412 382
rect 2406 377 2407 381
rect 2411 377 2412 381
rect 2406 376 2412 377
rect 2406 364 2412 365
rect 2406 360 2407 364
rect 2411 360 2412 364
rect 2406 359 2412 360
rect 2248 319 2250 336
rect 2336 319 2338 336
rect 2346 335 2352 336
rect 2346 331 2347 335
rect 2351 331 2352 335
rect 2346 330 2352 331
rect 2408 319 2410 359
rect 2247 318 2251 319
rect 2247 313 2251 314
rect 2279 318 2283 319
rect 2279 313 2283 314
rect 2335 318 2339 319
rect 2335 313 2339 314
rect 2359 318 2363 319
rect 2359 313 2363 314
rect 2407 318 2411 319
rect 2407 313 2411 314
rect 2226 307 2232 308
rect 2130 302 2136 303
rect 2198 303 2204 304
rect 2118 298 2124 299
rect 1238 275 1244 276
rect 1278 275 1284 276
rect 1598 275 1604 276
rect 1238 271 1239 275
rect 1243 271 1244 275
rect 1238 270 1244 271
rect 1598 271 1599 275
rect 1603 271 1604 275
rect 1598 270 1604 271
rect 1678 275 1684 276
rect 1678 271 1679 275
rect 1683 271 1684 275
rect 1678 270 1684 271
rect 1686 275 1692 276
rect 1686 271 1687 275
rect 1691 271 1692 275
rect 1686 270 1692 271
rect 1766 275 1772 276
rect 1766 271 1767 275
rect 1771 271 1772 275
rect 1766 270 1772 271
rect 1846 275 1852 276
rect 1846 271 1847 275
rect 1851 271 1852 275
rect 1846 270 1852 271
rect 1894 275 1900 276
rect 1894 271 1895 275
rect 1899 271 1900 275
rect 1894 270 1900 271
rect 1958 275 1964 276
rect 1958 271 1959 275
rect 1963 271 1964 275
rect 1958 270 1964 271
rect 2026 275 2032 276
rect 2026 271 2027 275
rect 2031 271 2032 275
rect 2026 270 2032 271
rect 2110 275 2116 276
rect 2110 271 2111 275
rect 2115 271 2116 275
rect 2110 270 2116 271
rect 838 268 844 269
rect 838 264 839 268
rect 843 264 844 268
rect 838 263 844 264
rect 840 255 842 263
rect 1240 255 1242 270
rect 1278 263 1284 264
rect 1278 259 1279 263
rect 1283 259 1284 263
rect 1278 258 1284 259
rect 831 254 835 255
rect 831 249 835 250
rect 839 254 843 255
rect 839 249 843 250
rect 879 254 883 255
rect 879 249 883 250
rect 927 254 931 255
rect 927 249 931 250
rect 975 254 979 255
rect 975 249 979 250
rect 1023 254 1027 255
rect 1023 249 1027 250
rect 1239 254 1243 255
rect 1239 249 1243 250
rect 830 248 836 249
rect 830 244 831 248
rect 835 244 836 248
rect 830 243 836 244
rect 878 248 884 249
rect 878 244 879 248
rect 883 244 884 248
rect 878 243 884 244
rect 926 248 932 249
rect 926 244 927 248
rect 931 244 932 248
rect 926 243 932 244
rect 974 248 980 249
rect 974 244 975 248
rect 979 244 980 248
rect 974 243 980 244
rect 1022 248 1028 249
rect 1022 244 1023 248
rect 1027 244 1028 248
rect 1022 243 1028 244
rect 1240 242 1242 249
rect 1280 247 1282 258
rect 1510 256 1516 257
rect 1510 252 1511 256
rect 1515 252 1516 256
rect 1510 251 1516 252
rect 1550 256 1556 257
rect 1550 252 1551 256
rect 1555 252 1556 256
rect 1550 251 1556 252
rect 1590 256 1596 257
rect 1590 252 1591 256
rect 1595 252 1596 256
rect 1590 251 1596 252
rect 1630 256 1636 257
rect 1630 252 1631 256
rect 1635 252 1636 256
rect 1630 251 1636 252
rect 1670 256 1676 257
rect 1670 252 1671 256
rect 1675 252 1676 256
rect 1670 251 1676 252
rect 1512 247 1514 251
rect 1552 247 1554 251
rect 1592 247 1594 251
rect 1632 247 1634 251
rect 1672 247 1674 251
rect 1279 246 1283 247
rect 1238 241 1244 242
rect 1279 241 1283 242
rect 1367 246 1371 247
rect 1367 241 1371 242
rect 1407 246 1411 247
rect 1407 241 1411 242
rect 1455 246 1459 247
rect 1455 241 1459 242
rect 1511 246 1515 247
rect 1511 241 1515 242
rect 1551 246 1555 247
rect 1551 241 1555 242
rect 1567 246 1571 247
rect 1567 241 1571 242
rect 1591 246 1595 247
rect 1591 241 1595 242
rect 1631 246 1635 247
rect 1631 241 1635 242
rect 1671 246 1675 247
rect 1671 241 1675 242
rect 1238 237 1239 241
rect 1243 237 1244 241
rect 1238 236 1244 237
rect 794 235 800 236
rect 794 231 795 235
rect 799 231 800 235
rect 1280 234 1282 241
rect 1366 240 1372 241
rect 1366 236 1367 240
rect 1371 236 1372 240
rect 1366 235 1372 236
rect 1406 240 1412 241
rect 1406 236 1407 240
rect 1411 236 1412 240
rect 1406 235 1412 236
rect 1454 240 1460 241
rect 1454 236 1455 240
rect 1459 236 1460 240
rect 1454 235 1460 236
rect 1510 240 1516 241
rect 1510 236 1511 240
rect 1515 236 1516 240
rect 1510 235 1516 236
rect 1566 240 1572 241
rect 1566 236 1567 240
rect 1571 236 1572 240
rect 1566 235 1572 236
rect 1630 240 1636 241
rect 1630 236 1631 240
rect 1635 236 1636 240
rect 1630 235 1636 236
rect 794 230 800 231
rect 1278 233 1284 234
rect 1278 229 1279 233
rect 1283 229 1284 233
rect 1278 228 1284 229
rect 742 227 748 228
rect 742 223 743 227
rect 747 223 748 227
rect 742 222 748 223
rect 1238 224 1244 225
rect 694 201 700 202
rect 694 197 695 201
rect 699 197 700 201
rect 694 196 700 197
rect 734 201 740 202
rect 734 197 735 201
rect 739 197 740 201
rect 734 196 740 197
rect 744 196 746 222
rect 1238 220 1239 224
rect 1243 220 1244 224
rect 1238 219 1244 220
rect 1414 219 1420 220
rect 782 201 788 202
rect 782 197 783 201
rect 787 197 788 201
rect 782 196 788 197
rect 830 201 836 202
rect 830 197 831 201
rect 835 197 836 201
rect 830 196 836 197
rect 878 201 884 202
rect 878 197 879 201
rect 883 197 884 201
rect 878 196 884 197
rect 926 201 932 202
rect 926 197 927 201
rect 931 197 932 201
rect 926 196 932 197
rect 974 201 980 202
rect 974 197 975 201
rect 979 197 980 201
rect 974 196 980 197
rect 1022 201 1028 202
rect 1022 197 1023 201
rect 1027 197 1028 201
rect 1022 196 1028 197
rect 648 155 650 196
rect 670 195 676 196
rect 670 191 671 195
rect 675 191 676 195
rect 670 190 676 191
rect 696 155 698 196
rect 736 155 738 196
rect 742 195 748 196
rect 742 191 743 195
rect 747 191 748 195
rect 742 190 748 191
rect 784 155 786 196
rect 832 155 834 196
rect 880 155 882 196
rect 928 155 930 196
rect 976 155 978 196
rect 1024 155 1026 196
rect 1038 195 1044 196
rect 1038 191 1039 195
rect 1043 191 1044 195
rect 1038 190 1044 191
rect 631 154 635 155
rect 631 149 635 150
rect 647 154 651 155
rect 647 149 651 150
rect 671 154 675 155
rect 671 149 675 150
rect 695 154 699 155
rect 695 149 699 150
rect 711 154 715 155
rect 711 149 715 150
rect 735 154 739 155
rect 735 149 739 150
rect 751 154 755 155
rect 751 149 755 150
rect 783 154 787 155
rect 783 149 787 150
rect 791 154 795 155
rect 791 149 795 150
rect 831 154 835 155
rect 831 149 835 150
rect 871 154 875 155
rect 871 149 875 150
rect 879 154 883 155
rect 879 149 883 150
rect 911 154 915 155
rect 911 149 915 150
rect 927 154 931 155
rect 927 149 931 150
rect 951 154 955 155
rect 951 149 955 150
rect 975 154 979 155
rect 975 149 979 150
rect 991 154 995 155
rect 991 149 995 150
rect 1023 154 1027 155
rect 1023 149 1027 150
rect 1031 154 1035 155
rect 1031 149 1035 150
rect 614 143 620 144
rect 578 138 584 139
rect 590 139 596 140
rect 550 134 556 135
rect 546 111 552 112
rect 546 110 547 111
rect 540 108 547 110
rect 506 106 512 107
rect 546 107 547 108
rect 551 107 552 111
rect 580 110 582 138
rect 590 135 591 139
rect 595 135 596 139
rect 614 139 615 143
rect 619 139 620 143
rect 632 140 634 149
rect 658 143 664 144
rect 614 138 620 139
rect 630 139 636 140
rect 590 134 596 135
rect 630 135 631 139
rect 635 135 636 139
rect 658 139 659 143
rect 663 139 664 143
rect 672 140 674 149
rect 698 143 704 144
rect 658 138 664 139
rect 670 139 676 140
rect 630 134 636 135
rect 651 116 655 117
rect 586 111 592 112
rect 586 110 587 111
rect 580 108 587 110
rect 546 106 552 107
rect 586 107 587 108
rect 591 107 592 111
rect 586 106 592 107
rect 650 111 656 112
rect 650 107 651 111
rect 655 107 656 111
rect 660 110 662 138
rect 670 135 671 139
rect 675 135 676 139
rect 698 139 699 143
rect 703 139 704 143
rect 712 140 714 149
rect 738 143 744 144
rect 698 138 704 139
rect 710 139 716 140
rect 670 134 676 135
rect 666 111 672 112
rect 666 110 667 111
rect 660 108 667 110
rect 650 106 656 107
rect 666 107 667 108
rect 671 107 672 111
rect 700 110 702 138
rect 710 135 711 139
rect 715 135 716 139
rect 738 139 739 143
rect 743 139 744 143
rect 752 140 754 149
rect 778 143 784 144
rect 738 138 744 139
rect 750 139 756 140
rect 710 134 716 135
rect 706 111 712 112
rect 706 110 707 111
rect 700 108 707 110
rect 666 106 672 107
rect 706 107 707 108
rect 711 107 712 111
rect 740 110 742 138
rect 750 135 751 139
rect 755 135 756 139
rect 778 139 779 143
rect 783 139 784 143
rect 792 140 794 149
rect 818 143 824 144
rect 778 138 784 139
rect 790 139 796 140
rect 750 134 756 135
rect 746 111 752 112
rect 746 110 747 111
rect 740 108 747 110
rect 706 106 712 107
rect 746 107 747 108
rect 751 107 752 111
rect 780 110 782 138
rect 790 135 791 139
rect 795 135 796 139
rect 818 139 819 143
rect 823 139 824 143
rect 832 140 834 149
rect 858 143 864 144
rect 818 138 824 139
rect 830 139 836 140
rect 790 134 796 135
rect 786 111 792 112
rect 786 110 787 111
rect 780 108 787 110
rect 746 106 752 107
rect 786 107 787 108
rect 791 107 792 111
rect 820 110 822 138
rect 830 135 831 139
rect 835 135 836 139
rect 858 139 859 143
rect 863 139 864 143
rect 872 140 874 149
rect 898 143 904 144
rect 858 138 864 139
rect 870 139 876 140
rect 830 134 836 135
rect 826 111 832 112
rect 826 110 827 111
rect 820 108 827 110
rect 786 106 792 107
rect 826 107 827 108
rect 831 107 832 111
rect 860 110 862 138
rect 870 135 871 139
rect 875 135 876 139
rect 898 139 899 143
rect 903 139 904 143
rect 912 140 914 149
rect 938 143 944 144
rect 898 138 904 139
rect 910 139 916 140
rect 870 134 876 135
rect 866 111 872 112
rect 866 110 867 111
rect 860 108 867 110
rect 826 106 832 107
rect 866 107 867 108
rect 871 107 872 111
rect 900 110 902 138
rect 910 135 911 139
rect 915 135 916 139
rect 938 139 939 143
rect 943 139 944 143
rect 952 140 954 149
rect 978 143 984 144
rect 938 138 944 139
rect 950 139 956 140
rect 910 134 916 135
rect 906 111 912 112
rect 906 110 907 111
rect 900 108 907 110
rect 866 106 872 107
rect 906 107 907 108
rect 911 107 912 111
rect 940 110 942 138
rect 950 135 951 139
rect 955 135 956 139
rect 978 139 979 143
rect 983 139 984 143
rect 992 140 994 149
rect 1018 143 1024 144
rect 978 138 984 139
rect 990 139 996 140
rect 950 134 956 135
rect 946 111 952 112
rect 946 110 947 111
rect 940 108 947 110
rect 906 106 912 107
rect 946 107 947 108
rect 951 107 952 111
rect 980 110 982 138
rect 990 135 991 139
rect 995 135 996 139
rect 1018 139 1019 143
rect 1023 139 1024 143
rect 1032 140 1034 149
rect 1018 138 1024 139
rect 1030 139 1036 140
rect 990 134 996 135
rect 986 111 992 112
rect 986 110 987 111
rect 980 108 987 110
rect 946 106 952 107
rect 986 107 987 108
rect 991 107 992 111
rect 1020 110 1022 138
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1040 117 1042 190
rect 1240 155 1242 219
rect 1278 216 1284 217
rect 1278 212 1279 216
rect 1283 212 1284 216
rect 1414 215 1415 219
rect 1419 215 1420 219
rect 1414 214 1420 215
rect 1278 211 1284 212
rect 1280 171 1282 211
rect 1366 193 1372 194
rect 1366 189 1367 193
rect 1371 189 1372 193
rect 1366 188 1372 189
rect 1406 193 1412 194
rect 1406 189 1407 193
rect 1411 189 1412 193
rect 1406 188 1412 189
rect 1416 188 1418 214
rect 1670 211 1676 212
rect 1670 207 1671 211
rect 1675 207 1676 211
rect 1670 206 1676 207
rect 1454 193 1460 194
rect 1454 189 1455 193
rect 1459 189 1460 193
rect 1454 188 1460 189
rect 1510 193 1516 194
rect 1510 189 1511 193
rect 1515 189 1516 193
rect 1510 188 1516 189
rect 1566 193 1572 194
rect 1566 189 1567 193
rect 1571 189 1572 193
rect 1566 188 1572 189
rect 1630 193 1636 194
rect 1630 189 1631 193
rect 1635 189 1636 193
rect 1630 188 1636 189
rect 1368 171 1370 188
rect 1408 171 1410 188
rect 1414 187 1420 188
rect 1414 183 1415 187
rect 1419 183 1420 187
rect 1414 182 1420 183
rect 1456 171 1458 188
rect 1512 171 1514 188
rect 1568 171 1570 188
rect 1632 171 1634 188
rect 1279 170 1283 171
rect 1279 165 1283 166
rect 1303 170 1307 171
rect 1303 165 1307 166
rect 1343 170 1347 171
rect 1343 165 1347 166
rect 1367 170 1371 171
rect 1367 165 1371 166
rect 1383 170 1387 171
rect 1383 165 1387 166
rect 1407 170 1411 171
rect 1407 165 1411 166
rect 1423 170 1427 171
rect 1423 165 1427 166
rect 1455 170 1459 171
rect 1455 165 1459 166
rect 1463 170 1467 171
rect 1463 165 1467 166
rect 1511 170 1515 171
rect 1511 165 1515 166
rect 1519 170 1523 171
rect 1519 165 1523 166
rect 1567 170 1571 171
rect 1567 165 1571 166
rect 1583 170 1587 171
rect 1583 165 1587 166
rect 1631 170 1635 171
rect 1631 165 1635 166
rect 1647 170 1651 171
rect 1647 165 1651 166
rect 1071 154 1075 155
rect 1071 149 1075 150
rect 1111 154 1115 155
rect 1111 149 1115 150
rect 1151 154 1155 155
rect 1151 149 1155 150
rect 1191 154 1195 155
rect 1191 149 1195 150
rect 1239 154 1243 155
rect 1239 149 1243 150
rect 1058 143 1064 144
rect 1058 139 1059 143
rect 1063 139 1064 143
rect 1072 140 1074 149
rect 1098 143 1104 144
rect 1058 138 1064 139
rect 1070 139 1076 140
rect 1039 116 1043 117
rect 1026 111 1032 112
rect 1039 111 1043 112
rect 1026 110 1027 111
rect 1020 108 1027 110
rect 986 106 992 107
rect 1026 107 1027 108
rect 1031 107 1032 111
rect 1060 110 1062 138
rect 1070 135 1071 139
rect 1075 135 1076 139
rect 1098 139 1099 143
rect 1103 139 1104 143
rect 1112 140 1114 149
rect 1152 140 1154 149
rect 1166 147 1172 148
rect 1166 143 1167 147
rect 1171 143 1172 147
rect 1166 142 1172 143
rect 1098 138 1104 139
rect 1110 139 1116 140
rect 1070 134 1076 135
rect 1066 111 1072 112
rect 1066 110 1067 111
rect 1060 108 1067 110
rect 1026 106 1032 107
rect 1066 107 1067 108
rect 1071 107 1072 111
rect 1100 110 1102 138
rect 1110 135 1111 139
rect 1115 135 1116 139
rect 1110 134 1116 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1168 112 1170 142
rect 1192 140 1194 149
rect 1198 147 1204 148
rect 1198 143 1199 147
rect 1203 143 1204 147
rect 1198 142 1204 143
rect 1190 139 1196 140
rect 1190 135 1191 139
rect 1195 135 1196 139
rect 1190 134 1196 135
rect 1200 112 1202 142
rect 1240 117 1242 149
rect 1280 133 1282 165
rect 1304 156 1306 165
rect 1330 159 1336 160
rect 1302 155 1308 156
rect 1302 151 1303 155
rect 1307 151 1308 155
rect 1330 155 1331 159
rect 1335 155 1336 159
rect 1344 156 1346 165
rect 1370 159 1376 160
rect 1330 154 1336 155
rect 1342 155 1348 156
rect 1302 150 1308 151
rect 1278 132 1284 133
rect 1278 128 1279 132
rect 1283 128 1284 132
rect 1278 127 1284 128
rect 1332 126 1334 154
rect 1342 151 1343 155
rect 1347 151 1348 155
rect 1370 155 1371 159
rect 1375 155 1376 159
rect 1384 156 1386 165
rect 1410 159 1416 160
rect 1370 154 1376 155
rect 1382 155 1388 156
rect 1342 150 1348 151
rect 1338 127 1344 128
rect 1338 126 1339 127
rect 1332 124 1339 126
rect 1338 123 1339 124
rect 1343 123 1344 127
rect 1372 126 1374 154
rect 1382 151 1383 155
rect 1387 151 1388 155
rect 1410 155 1411 159
rect 1415 155 1416 159
rect 1424 156 1426 165
rect 1450 159 1456 160
rect 1410 154 1416 155
rect 1422 155 1428 156
rect 1382 150 1388 151
rect 1378 127 1384 128
rect 1378 126 1379 127
rect 1372 124 1379 126
rect 1338 122 1344 123
rect 1378 123 1379 124
rect 1383 123 1384 127
rect 1412 126 1414 154
rect 1422 151 1423 155
rect 1427 151 1428 155
rect 1450 155 1451 159
rect 1455 155 1456 159
rect 1464 156 1466 165
rect 1510 159 1516 160
rect 1450 154 1456 155
rect 1462 155 1468 156
rect 1422 150 1428 151
rect 1418 127 1424 128
rect 1418 126 1419 127
rect 1412 124 1419 126
rect 1378 122 1384 123
rect 1418 123 1419 124
rect 1423 123 1424 127
rect 1452 126 1454 154
rect 1462 151 1463 155
rect 1467 151 1468 155
rect 1510 155 1511 159
rect 1515 155 1516 159
rect 1520 156 1522 165
rect 1574 159 1580 160
rect 1510 154 1516 155
rect 1518 155 1524 156
rect 1462 150 1468 151
rect 1512 128 1514 154
rect 1518 151 1519 155
rect 1523 151 1524 155
rect 1574 155 1575 159
rect 1579 155 1580 159
rect 1584 156 1586 165
rect 1638 159 1644 160
rect 1574 154 1580 155
rect 1582 155 1588 156
rect 1518 150 1524 151
rect 1576 128 1578 154
rect 1582 151 1583 155
rect 1587 151 1588 155
rect 1638 155 1639 159
rect 1643 155 1644 159
rect 1648 156 1650 165
rect 1672 160 1674 206
rect 1680 188 1682 270
rect 1710 256 1716 257
rect 1710 252 1711 256
rect 1715 252 1716 256
rect 1710 251 1716 252
rect 1750 256 1756 257
rect 1750 252 1751 256
rect 1755 252 1756 256
rect 1750 251 1756 252
rect 1790 256 1796 257
rect 1790 252 1791 256
rect 1795 252 1796 256
rect 1790 251 1796 252
rect 1838 256 1844 257
rect 1838 252 1839 256
rect 1843 252 1844 256
rect 1838 251 1844 252
rect 1902 256 1908 257
rect 1902 252 1903 256
rect 1907 252 1908 256
rect 1902 251 1908 252
rect 1966 256 1972 257
rect 1966 252 1967 256
rect 1971 252 1972 256
rect 1966 251 1972 252
rect 2038 256 2044 257
rect 2038 252 2039 256
rect 2043 252 2044 256
rect 2038 251 2044 252
rect 2118 256 2124 257
rect 2118 252 2119 256
rect 2123 252 2124 256
rect 2118 251 2124 252
rect 1712 247 1714 251
rect 1752 247 1754 251
rect 1792 247 1794 251
rect 1840 247 1842 251
rect 1904 247 1906 251
rect 1968 247 1970 251
rect 2040 247 2042 251
rect 2120 247 2122 251
rect 1703 246 1707 247
rect 1703 241 1707 242
rect 1711 246 1715 247
rect 1711 241 1715 242
rect 1751 246 1755 247
rect 1751 241 1755 242
rect 1775 246 1779 247
rect 1775 241 1779 242
rect 1791 246 1795 247
rect 1791 241 1795 242
rect 1839 246 1843 247
rect 1839 241 1843 242
rect 1855 246 1859 247
rect 1855 241 1859 242
rect 1903 246 1907 247
rect 1903 241 1907 242
rect 1943 246 1947 247
rect 1943 241 1947 242
rect 1967 246 1971 247
rect 1967 241 1971 242
rect 2031 246 2035 247
rect 2031 241 2035 242
rect 2039 246 2043 247
rect 2039 241 2043 242
rect 2119 246 2123 247
rect 2119 241 2123 242
rect 1702 240 1708 241
rect 1702 236 1703 240
rect 1707 236 1708 240
rect 1702 235 1708 236
rect 1774 240 1780 241
rect 1774 236 1775 240
rect 1779 236 1780 240
rect 1774 235 1780 236
rect 1854 240 1860 241
rect 1854 236 1855 240
rect 1859 236 1860 240
rect 1854 235 1860 236
rect 1942 240 1948 241
rect 1942 236 1943 240
rect 1947 236 1948 240
rect 1942 235 1948 236
rect 2030 240 2036 241
rect 2030 236 2031 240
rect 2035 236 2036 240
rect 2030 235 2036 236
rect 2118 240 2124 241
rect 2118 236 2119 240
rect 2123 236 2124 240
rect 2118 235 2124 236
rect 2132 228 2134 302
rect 2198 299 2199 303
rect 2203 299 2204 303
rect 2226 303 2227 307
rect 2231 303 2232 307
rect 2280 304 2282 313
rect 2290 307 2296 308
rect 2226 302 2232 303
rect 2278 303 2284 304
rect 2198 298 2204 299
rect 2278 299 2279 303
rect 2283 299 2284 303
rect 2290 303 2291 307
rect 2295 303 2296 307
rect 2360 304 2362 313
rect 2370 307 2376 308
rect 2290 302 2296 303
rect 2358 303 2364 304
rect 2278 298 2284 299
rect 2292 276 2294 302
rect 2358 299 2359 303
rect 2363 299 2364 303
rect 2370 303 2371 307
rect 2375 303 2376 307
rect 2370 302 2376 303
rect 2358 298 2364 299
rect 2372 276 2374 302
rect 2408 281 2410 313
rect 2406 280 2412 281
rect 2406 276 2407 280
rect 2411 276 2412 280
rect 2290 275 2296 276
rect 2290 271 2291 275
rect 2295 271 2296 275
rect 2290 270 2296 271
rect 2370 275 2376 276
rect 2406 275 2412 276
rect 2370 271 2371 275
rect 2375 271 2376 275
rect 2370 270 2376 271
rect 2322 267 2328 268
rect 2322 263 2323 267
rect 2327 263 2328 267
rect 2322 262 2328 263
rect 2406 263 2412 264
rect 2198 256 2204 257
rect 2198 252 2199 256
rect 2203 252 2204 256
rect 2198 251 2204 252
rect 2278 256 2284 257
rect 2278 252 2279 256
rect 2283 252 2284 256
rect 2278 251 2284 252
rect 2200 247 2202 251
rect 2280 247 2282 251
rect 2199 246 2203 247
rect 2199 241 2203 242
rect 2207 246 2211 247
rect 2207 241 2211 242
rect 2279 246 2283 247
rect 2279 241 2283 242
rect 2295 246 2299 247
rect 2295 241 2299 242
rect 2206 240 2212 241
rect 2206 236 2207 240
rect 2211 236 2212 240
rect 2206 235 2212 236
rect 2294 240 2300 241
rect 2294 236 2295 240
rect 2299 236 2300 240
rect 2294 235 2300 236
rect 2130 227 2136 228
rect 2130 223 2131 227
rect 2135 223 2136 227
rect 2130 222 2136 223
rect 2226 219 2232 220
rect 2226 215 2227 219
rect 2231 215 2232 219
rect 2226 214 2232 215
rect 1702 193 1708 194
rect 1702 189 1703 193
rect 1707 189 1708 193
rect 1702 188 1708 189
rect 1774 193 1780 194
rect 1774 189 1775 193
rect 1779 189 1780 193
rect 1774 188 1780 189
rect 1854 193 1860 194
rect 1854 189 1855 193
rect 1859 189 1860 193
rect 1854 188 1860 189
rect 1942 193 1948 194
rect 1942 189 1943 193
rect 1947 189 1948 193
rect 1942 188 1948 189
rect 2030 193 2036 194
rect 2030 189 2031 193
rect 2035 189 2036 193
rect 2030 188 2036 189
rect 2118 193 2124 194
rect 2118 189 2119 193
rect 2123 189 2124 193
rect 2118 188 2124 189
rect 2206 193 2212 194
rect 2206 189 2207 193
rect 2211 189 2212 193
rect 2206 188 2212 189
rect 1678 187 1684 188
rect 1678 183 1679 187
rect 1683 183 1684 187
rect 1678 182 1684 183
rect 1704 171 1706 188
rect 1738 179 1744 180
rect 1738 175 1739 179
rect 1743 175 1744 179
rect 1738 174 1744 175
rect 1703 170 1707 171
rect 1703 165 1707 166
rect 1711 170 1715 171
rect 1711 165 1715 166
rect 1670 159 1676 160
rect 1638 154 1644 155
rect 1646 155 1652 156
rect 1582 150 1588 151
rect 1640 128 1642 154
rect 1646 151 1647 155
rect 1651 151 1652 155
rect 1670 155 1671 159
rect 1675 155 1676 159
rect 1712 156 1714 165
rect 1670 154 1676 155
rect 1710 155 1716 156
rect 1646 150 1652 151
rect 1710 151 1711 155
rect 1715 151 1716 155
rect 1710 150 1716 151
rect 1740 128 1742 174
rect 1776 171 1778 188
rect 1856 171 1858 188
rect 1944 171 1946 188
rect 2032 171 2034 188
rect 2120 171 2122 188
rect 2208 171 2210 188
rect 1775 170 1779 171
rect 1775 165 1779 166
rect 1831 170 1835 171
rect 1831 165 1835 166
rect 1855 170 1859 171
rect 1855 165 1859 166
rect 1887 170 1891 171
rect 1887 165 1891 166
rect 1935 170 1939 171
rect 1935 165 1939 166
rect 1943 170 1947 171
rect 1943 165 1947 166
rect 1975 170 1979 171
rect 1975 165 1979 166
rect 2015 170 2019 171
rect 2015 165 2019 166
rect 2031 170 2035 171
rect 2031 165 2035 166
rect 2055 170 2059 171
rect 2055 165 2059 166
rect 2095 170 2099 171
rect 2095 165 2099 166
rect 2119 170 2123 171
rect 2119 165 2123 166
rect 2143 170 2147 171
rect 2143 165 2147 166
rect 2191 170 2195 171
rect 2191 165 2195 166
rect 2207 170 2211 171
rect 2207 165 2211 166
rect 1766 159 1772 160
rect 1766 155 1767 159
rect 1771 155 1772 159
rect 1776 156 1778 165
rect 1822 159 1828 160
rect 1766 154 1772 155
rect 1774 155 1780 156
rect 1768 128 1770 154
rect 1774 151 1775 155
rect 1779 151 1780 155
rect 1822 155 1823 159
rect 1827 155 1828 159
rect 1832 156 1834 165
rect 1878 159 1884 160
rect 1822 154 1828 155
rect 1830 155 1836 156
rect 1774 150 1780 151
rect 1824 128 1826 154
rect 1830 151 1831 155
rect 1835 151 1836 155
rect 1878 155 1879 159
rect 1883 155 1884 159
rect 1888 156 1890 165
rect 1926 159 1932 160
rect 1878 154 1884 155
rect 1886 155 1892 156
rect 1830 150 1836 151
rect 1880 128 1882 154
rect 1886 151 1887 155
rect 1891 151 1892 155
rect 1926 155 1927 159
rect 1931 155 1932 159
rect 1936 156 1938 165
rect 1962 159 1968 160
rect 1926 154 1932 155
rect 1934 155 1940 156
rect 1886 150 1892 151
rect 1928 128 1930 154
rect 1934 151 1935 155
rect 1939 151 1940 155
rect 1962 155 1963 159
rect 1967 155 1968 159
rect 1976 156 1978 165
rect 2016 156 2018 165
rect 2022 163 2028 164
rect 2022 159 2023 163
rect 2027 159 2028 163
rect 2022 158 2028 159
rect 1962 154 1968 155
rect 1974 155 1980 156
rect 1934 150 1940 151
rect 1964 136 1966 154
rect 1974 151 1975 155
rect 1979 151 1980 155
rect 1974 150 1980 151
rect 2014 155 2020 156
rect 2014 151 2015 155
rect 2019 151 2020 155
rect 2014 150 2020 151
rect 1962 135 1968 136
rect 1962 131 1963 135
rect 1967 131 1968 135
rect 1962 130 1968 131
rect 2024 128 2026 158
rect 2056 156 2058 165
rect 2070 163 2076 164
rect 2070 159 2071 163
rect 2075 159 2076 163
rect 2070 158 2076 159
rect 2054 155 2060 156
rect 2054 151 2055 155
rect 2059 151 2060 155
rect 2054 150 2060 151
rect 2072 128 2074 158
rect 2096 156 2098 165
rect 2102 163 2108 164
rect 2102 159 2103 163
rect 2107 159 2108 163
rect 2102 158 2108 159
rect 2134 159 2140 160
rect 2094 155 2100 156
rect 2094 151 2095 155
rect 2099 151 2100 155
rect 2094 150 2100 151
rect 2104 128 2106 158
rect 2134 155 2135 159
rect 2139 155 2140 159
rect 2144 156 2146 165
rect 2182 159 2188 160
rect 2134 154 2140 155
rect 2142 155 2148 156
rect 2136 128 2138 154
rect 2142 151 2143 155
rect 2147 151 2148 155
rect 2182 155 2183 159
rect 2187 155 2188 159
rect 2192 156 2194 165
rect 2228 160 2230 214
rect 2294 193 2300 194
rect 2294 189 2295 193
rect 2299 189 2300 193
rect 2294 188 2300 189
rect 2324 188 2326 262
rect 2406 259 2407 263
rect 2411 259 2412 263
rect 2406 258 2412 259
rect 2358 256 2364 257
rect 2358 252 2359 256
rect 2363 252 2364 256
rect 2358 251 2364 252
rect 2360 247 2362 251
rect 2408 247 2410 258
rect 2359 246 2363 247
rect 2359 241 2363 242
rect 2407 246 2411 247
rect 2407 241 2411 242
rect 2358 240 2364 241
rect 2358 236 2359 240
rect 2363 236 2364 240
rect 2358 235 2364 236
rect 2408 234 2410 241
rect 2406 233 2412 234
rect 2406 229 2407 233
rect 2411 229 2412 233
rect 2406 228 2412 229
rect 2374 219 2380 220
rect 2374 215 2375 219
rect 2379 215 2380 219
rect 2374 214 2380 215
rect 2382 219 2388 220
rect 2382 215 2383 219
rect 2387 215 2388 219
rect 2382 214 2388 215
rect 2406 216 2412 217
rect 2358 193 2364 194
rect 2358 189 2359 193
rect 2363 189 2364 193
rect 2358 188 2364 189
rect 2376 188 2378 214
rect 2262 187 2268 188
rect 2262 183 2263 187
rect 2267 183 2268 187
rect 2262 182 2268 183
rect 2239 170 2243 171
rect 2239 165 2243 166
rect 2226 159 2232 160
rect 2182 154 2188 155
rect 2190 155 2196 156
rect 2142 150 2148 151
rect 2184 128 2186 154
rect 2190 151 2191 155
rect 2195 151 2196 155
rect 2226 155 2227 159
rect 2231 155 2232 159
rect 2240 156 2242 165
rect 2226 154 2232 155
rect 2238 155 2244 156
rect 2190 150 2196 151
rect 2238 151 2239 155
rect 2243 151 2244 155
rect 2238 150 2244 151
rect 2264 128 2266 182
rect 2296 171 2298 188
rect 2322 187 2328 188
rect 2322 183 2323 187
rect 2327 183 2328 187
rect 2322 182 2328 183
rect 2360 171 2362 188
rect 2374 187 2380 188
rect 2374 183 2375 187
rect 2379 183 2380 187
rect 2374 182 2380 183
rect 2279 170 2283 171
rect 2279 165 2283 166
rect 2295 170 2299 171
rect 2295 165 2299 166
rect 2319 170 2323 171
rect 2319 165 2323 166
rect 2359 170 2363 171
rect 2359 165 2363 166
rect 2280 156 2282 165
rect 2286 163 2292 164
rect 2286 159 2287 163
rect 2291 159 2292 163
rect 2286 158 2292 159
rect 2278 155 2284 156
rect 2278 151 2279 155
rect 2283 151 2284 155
rect 2278 150 2284 151
rect 2288 128 2290 158
rect 2320 156 2322 165
rect 2334 163 2340 164
rect 2334 159 2335 163
rect 2339 159 2340 163
rect 2334 158 2340 159
rect 2318 155 2324 156
rect 2318 151 2319 155
rect 2323 151 2324 155
rect 2318 150 2324 151
rect 2336 128 2338 158
rect 2360 156 2362 165
rect 2366 163 2372 164
rect 2366 159 2367 163
rect 2371 159 2372 163
rect 2384 160 2386 214
rect 2406 212 2407 216
rect 2411 212 2412 216
rect 2406 211 2412 212
rect 2408 171 2410 211
rect 2407 170 2411 171
rect 2407 165 2411 166
rect 2366 158 2372 159
rect 2382 159 2388 160
rect 2358 155 2364 156
rect 2358 151 2359 155
rect 2363 151 2364 155
rect 2358 150 2364 151
rect 2368 128 2370 158
rect 2382 155 2383 159
rect 2387 155 2388 159
rect 2382 154 2388 155
rect 2408 133 2410 165
rect 2406 132 2412 133
rect 2406 128 2407 132
rect 2411 128 2412 132
rect 1458 127 1464 128
rect 1458 126 1459 127
rect 1452 124 1459 126
rect 1418 122 1424 123
rect 1458 123 1459 124
rect 1463 123 1464 127
rect 1458 122 1464 123
rect 1510 127 1516 128
rect 1510 123 1511 127
rect 1515 123 1516 127
rect 1510 122 1516 123
rect 1574 127 1580 128
rect 1574 123 1575 127
rect 1579 123 1580 127
rect 1574 122 1580 123
rect 1638 127 1644 128
rect 1638 123 1639 127
rect 1643 123 1644 127
rect 1638 122 1644 123
rect 1738 127 1744 128
rect 1738 123 1739 127
rect 1743 123 1744 127
rect 1738 122 1744 123
rect 1766 127 1772 128
rect 1766 123 1767 127
rect 1771 123 1772 127
rect 1766 122 1772 123
rect 1822 127 1828 128
rect 1822 123 1823 127
rect 1827 123 1828 127
rect 1822 122 1828 123
rect 1878 127 1884 128
rect 1878 123 1879 127
rect 1883 123 1884 127
rect 1878 122 1884 123
rect 1926 127 1932 128
rect 1926 123 1927 127
rect 1931 123 1932 127
rect 1926 122 1932 123
rect 2022 127 2028 128
rect 2022 123 2023 127
rect 2027 123 2028 127
rect 2022 122 2028 123
rect 2070 127 2076 128
rect 2070 123 2071 127
rect 2075 123 2076 127
rect 2070 122 2076 123
rect 2102 127 2108 128
rect 2102 123 2103 127
rect 2107 123 2108 127
rect 2102 122 2108 123
rect 2134 127 2140 128
rect 2134 123 2135 127
rect 2139 123 2140 127
rect 2134 122 2140 123
rect 2182 127 2188 128
rect 2182 123 2183 127
rect 2187 123 2188 127
rect 2182 122 2188 123
rect 2262 127 2268 128
rect 2262 123 2263 127
rect 2267 123 2268 127
rect 2262 122 2268 123
rect 2286 127 2292 128
rect 2286 123 2287 127
rect 2291 123 2292 127
rect 2286 122 2292 123
rect 2334 127 2340 128
rect 2334 123 2335 127
rect 2339 123 2340 127
rect 2334 122 2340 123
rect 2366 127 2372 128
rect 2406 127 2412 128
rect 2366 123 2367 127
rect 2371 123 2372 127
rect 2366 122 2372 123
rect 1238 116 1244 117
rect 1238 112 1239 116
rect 1243 112 1244 116
rect 1106 111 1112 112
rect 1106 110 1107 111
rect 1100 108 1107 110
rect 1066 106 1072 107
rect 1106 107 1107 108
rect 1111 107 1112 111
rect 1106 106 1112 107
rect 1166 111 1172 112
rect 1166 107 1167 111
rect 1171 107 1172 111
rect 1166 106 1172 107
rect 1198 111 1204 112
rect 1238 111 1244 112
rect 1278 115 1284 116
rect 1278 111 1279 115
rect 1283 111 1284 115
rect 1198 107 1199 111
rect 1203 107 1204 111
rect 1278 110 1284 111
rect 2406 115 2412 116
rect 2406 111 2407 115
rect 2411 111 2412 115
rect 2406 110 2412 111
rect 1198 106 1204 107
rect 1280 103 1282 110
rect 1302 108 1308 109
rect 1302 104 1303 108
rect 1307 104 1308 108
rect 1302 103 1308 104
rect 1342 108 1348 109
rect 1342 104 1343 108
rect 1347 104 1348 108
rect 1342 103 1348 104
rect 1382 108 1388 109
rect 1382 104 1383 108
rect 1387 104 1388 108
rect 1382 103 1388 104
rect 1422 108 1428 109
rect 1422 104 1423 108
rect 1427 104 1428 108
rect 1422 103 1428 104
rect 1462 108 1468 109
rect 1462 104 1463 108
rect 1467 104 1468 108
rect 1462 103 1468 104
rect 1518 108 1524 109
rect 1518 104 1519 108
rect 1523 104 1524 108
rect 1518 103 1524 104
rect 1582 108 1588 109
rect 1582 104 1583 108
rect 1587 104 1588 108
rect 1582 103 1588 104
rect 1646 108 1652 109
rect 1646 104 1647 108
rect 1651 104 1652 108
rect 1646 103 1652 104
rect 1710 108 1716 109
rect 1710 104 1711 108
rect 1715 104 1716 108
rect 1710 103 1716 104
rect 1774 108 1780 109
rect 1774 104 1775 108
rect 1779 104 1780 108
rect 1774 103 1780 104
rect 1830 108 1836 109
rect 1830 104 1831 108
rect 1835 104 1836 108
rect 1830 103 1836 104
rect 1886 108 1892 109
rect 1886 104 1887 108
rect 1891 104 1892 108
rect 1886 103 1892 104
rect 1934 108 1940 109
rect 1934 104 1935 108
rect 1939 104 1940 108
rect 1934 103 1940 104
rect 1974 108 1980 109
rect 1974 104 1975 108
rect 1979 104 1980 108
rect 1974 103 1980 104
rect 2014 108 2020 109
rect 2014 104 2015 108
rect 2019 104 2020 108
rect 2014 103 2020 104
rect 2054 108 2060 109
rect 2054 104 2055 108
rect 2059 104 2060 108
rect 2054 103 2060 104
rect 2094 108 2100 109
rect 2094 104 2095 108
rect 2099 104 2100 108
rect 2094 103 2100 104
rect 2142 108 2148 109
rect 2142 104 2143 108
rect 2147 104 2148 108
rect 2142 103 2148 104
rect 2190 108 2196 109
rect 2190 104 2191 108
rect 2195 104 2196 108
rect 2190 103 2196 104
rect 2238 108 2244 109
rect 2238 104 2239 108
rect 2243 104 2244 108
rect 2238 103 2244 104
rect 2278 108 2284 109
rect 2278 104 2279 108
rect 2283 104 2284 108
rect 2278 103 2284 104
rect 2318 108 2324 109
rect 2318 104 2319 108
rect 2323 104 2324 108
rect 2318 103 2324 104
rect 2358 108 2364 109
rect 2358 104 2359 108
rect 2363 104 2364 108
rect 2358 103 2364 104
rect 2408 103 2410 110
rect 1279 102 1283 103
rect 110 99 116 100
rect 110 95 111 99
rect 115 95 116 99
rect 110 94 116 95
rect 1238 99 1244 100
rect 1238 95 1239 99
rect 1243 95 1244 99
rect 1279 97 1283 98
rect 1303 102 1307 103
rect 1303 97 1307 98
rect 1343 102 1347 103
rect 1343 97 1347 98
rect 1383 102 1387 103
rect 1383 97 1387 98
rect 1423 102 1427 103
rect 1423 97 1427 98
rect 1463 102 1467 103
rect 1463 97 1467 98
rect 1519 102 1523 103
rect 1519 97 1523 98
rect 1583 102 1587 103
rect 1583 97 1587 98
rect 1647 102 1651 103
rect 1647 97 1651 98
rect 1711 102 1715 103
rect 1711 97 1715 98
rect 1775 102 1779 103
rect 1775 97 1779 98
rect 1831 102 1835 103
rect 1831 97 1835 98
rect 1887 102 1891 103
rect 1887 97 1891 98
rect 1935 102 1939 103
rect 1935 97 1939 98
rect 1975 102 1979 103
rect 1975 97 1979 98
rect 2015 102 2019 103
rect 2015 97 2019 98
rect 2055 102 2059 103
rect 2055 97 2059 98
rect 2095 102 2099 103
rect 2095 97 2099 98
rect 2143 102 2147 103
rect 2143 97 2147 98
rect 2191 102 2195 103
rect 2191 97 2195 98
rect 2239 102 2243 103
rect 2239 97 2243 98
rect 2279 102 2283 103
rect 2279 97 2283 98
rect 2319 102 2323 103
rect 2319 97 2323 98
rect 2359 102 2363 103
rect 2359 97 2363 98
rect 2407 102 2411 103
rect 2407 97 2411 98
rect 1238 94 1244 95
rect 112 87 114 94
rect 150 92 156 93
rect 150 88 151 92
rect 155 88 156 92
rect 150 87 156 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 230 92 236 93
rect 230 88 231 92
rect 235 88 236 92
rect 230 87 236 88
rect 270 92 276 93
rect 270 88 271 92
rect 275 88 276 92
rect 270 87 276 88
rect 310 92 316 93
rect 310 88 311 92
rect 315 88 316 92
rect 310 87 316 88
rect 350 92 356 93
rect 350 88 351 92
rect 355 88 356 92
rect 350 87 356 88
rect 390 92 396 93
rect 390 88 391 92
rect 395 88 396 92
rect 390 87 396 88
rect 430 92 436 93
rect 430 88 431 92
rect 435 88 436 92
rect 430 87 436 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 510 92 516 93
rect 510 88 511 92
rect 515 88 516 92
rect 510 87 516 88
rect 550 92 556 93
rect 550 88 551 92
rect 555 88 556 92
rect 550 87 556 88
rect 590 92 596 93
rect 590 88 591 92
rect 595 88 596 92
rect 590 87 596 88
rect 630 92 636 93
rect 630 88 631 92
rect 635 88 636 92
rect 630 87 636 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 710 92 716 93
rect 710 88 711 92
rect 715 88 716 92
rect 710 87 716 88
rect 750 92 756 93
rect 750 88 751 92
rect 755 88 756 92
rect 750 87 756 88
rect 790 92 796 93
rect 790 88 791 92
rect 795 88 796 92
rect 790 87 796 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 870 92 876 93
rect 870 88 871 92
rect 875 88 876 92
rect 870 87 876 88
rect 910 92 916 93
rect 910 88 911 92
rect 915 88 916 92
rect 910 87 916 88
rect 950 92 956 93
rect 950 88 951 92
rect 955 88 956 92
rect 950 87 956 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1030 92 1036 93
rect 1030 88 1031 92
rect 1035 88 1036 92
rect 1030 87 1036 88
rect 1070 92 1076 93
rect 1070 88 1071 92
rect 1075 88 1076 92
rect 1070 87 1076 88
rect 1110 92 1116 93
rect 1110 88 1111 92
rect 1115 88 1116 92
rect 1110 87 1116 88
rect 1150 92 1156 93
rect 1150 88 1151 92
rect 1155 88 1156 92
rect 1150 87 1156 88
rect 1190 92 1196 93
rect 1190 88 1191 92
rect 1195 88 1196 92
rect 1190 87 1196 88
rect 1240 87 1242 94
rect 111 86 115 87
rect 111 81 115 82
rect 151 86 155 87
rect 151 81 155 82
rect 191 86 195 87
rect 191 81 195 82
rect 231 86 235 87
rect 231 81 235 82
rect 271 86 275 87
rect 271 81 275 82
rect 311 86 315 87
rect 311 81 315 82
rect 351 86 355 87
rect 351 81 355 82
rect 391 86 395 87
rect 391 81 395 82
rect 431 86 435 87
rect 431 81 435 82
rect 471 86 475 87
rect 471 81 475 82
rect 511 86 515 87
rect 511 81 515 82
rect 551 86 555 87
rect 551 81 555 82
rect 591 86 595 87
rect 591 81 595 82
rect 631 86 635 87
rect 631 81 635 82
rect 671 86 675 87
rect 671 81 675 82
rect 711 86 715 87
rect 711 81 715 82
rect 751 86 755 87
rect 751 81 755 82
rect 791 86 795 87
rect 791 81 795 82
rect 831 86 835 87
rect 831 81 835 82
rect 871 86 875 87
rect 871 81 875 82
rect 911 86 915 87
rect 911 81 915 82
rect 951 86 955 87
rect 951 81 955 82
rect 991 86 995 87
rect 991 81 995 82
rect 1031 86 1035 87
rect 1031 81 1035 82
rect 1071 86 1075 87
rect 1071 81 1075 82
rect 1111 86 1115 87
rect 1111 81 1115 82
rect 1151 86 1155 87
rect 1151 81 1155 82
rect 1191 86 1195 87
rect 1191 81 1195 82
rect 1239 86 1243 87
rect 1239 81 1243 82
<< m4c >>
rect 111 2490 115 2494
rect 231 2490 235 2494
rect 271 2490 275 2494
rect 311 2490 315 2494
rect 351 2490 355 2494
rect 399 2490 403 2494
rect 455 2490 459 2494
rect 511 2490 515 2494
rect 575 2490 579 2494
rect 639 2490 643 2494
rect 703 2490 707 2494
rect 767 2490 771 2494
rect 823 2490 827 2494
rect 879 2490 883 2494
rect 927 2490 931 2494
rect 975 2490 979 2494
rect 1023 2490 1027 2494
rect 1071 2490 1075 2494
rect 1111 2490 1115 2494
rect 1151 2490 1155 2494
rect 1191 2490 1195 2494
rect 1239 2490 1243 2494
rect 111 2414 115 2418
rect 199 2414 203 2418
rect 231 2414 235 2418
rect 263 2414 267 2418
rect 271 2414 275 2418
rect 311 2414 315 2418
rect 327 2414 331 2418
rect 351 2414 355 2418
rect 399 2414 403 2418
rect 455 2414 459 2418
rect 471 2414 475 2418
rect 511 2414 515 2418
rect 543 2414 547 2418
rect 575 2414 579 2418
rect 615 2414 619 2418
rect 639 2414 643 2418
rect 1279 2486 1283 2490
rect 1303 2486 1307 2490
rect 1343 2486 1347 2490
rect 1383 2486 1387 2490
rect 1439 2486 1443 2490
rect 1511 2486 1515 2490
rect 1583 2486 1587 2490
rect 1663 2486 1667 2490
rect 1735 2486 1739 2490
rect 1807 2486 1811 2490
rect 1887 2486 1891 2490
rect 1967 2486 1971 2490
rect 2063 2486 2067 2490
rect 2167 2486 2171 2490
rect 2271 2486 2275 2490
rect 2359 2486 2363 2490
rect 2407 2486 2411 2490
rect 687 2414 691 2418
rect 703 2414 707 2418
rect 751 2414 755 2418
rect 767 2414 771 2418
rect 111 2342 115 2346
rect 199 2342 203 2346
rect 263 2342 267 2346
rect 271 2342 275 2346
rect 327 2342 331 2346
rect 399 2342 403 2346
rect 823 2414 827 2418
rect 879 2414 883 2418
rect 895 2414 899 2418
rect 927 2414 931 2418
rect 967 2414 971 2418
rect 975 2414 979 2418
rect 1023 2414 1027 2418
rect 1071 2414 1075 2418
rect 1111 2414 1115 2418
rect 1151 2414 1155 2418
rect 1191 2414 1195 2418
rect 1239 2414 1243 2418
rect 1279 2418 1283 2422
rect 1303 2418 1307 2422
rect 1343 2418 1347 2422
rect 1375 2418 1379 2422
rect 1383 2418 1387 2422
rect 1415 2418 1419 2422
rect 1439 2418 1443 2422
rect 1455 2418 1459 2422
rect 1503 2418 1507 2422
rect 1511 2418 1515 2422
rect 1559 2418 1563 2422
rect 1583 2418 1587 2422
rect 1615 2418 1619 2422
rect 1663 2418 1667 2422
rect 1679 2418 1683 2422
rect 1735 2418 1739 2422
rect 1799 2418 1803 2422
rect 1807 2418 1811 2422
rect 1871 2418 1875 2422
rect 1887 2418 1891 2422
rect 1951 2418 1955 2422
rect 1967 2418 1971 2422
rect 471 2342 475 2346
rect 543 2342 547 2346
rect 551 2342 555 2346
rect 615 2342 619 2346
rect 631 2342 635 2346
rect 687 2342 691 2346
rect 711 2342 715 2346
rect 111 2266 115 2270
rect 143 2266 147 2270
rect 183 2266 187 2270
rect 223 2266 227 2270
rect 271 2266 275 2270
rect 279 2266 283 2270
rect 327 2266 331 2270
rect 335 2266 339 2270
rect 399 2266 403 2270
rect 407 2266 411 2270
rect 471 2266 475 2270
rect 479 2266 483 2270
rect 551 2266 555 2270
rect 559 2266 563 2270
rect 111 2198 115 2202
rect 135 2198 139 2202
rect 143 2198 147 2202
rect 183 2198 187 2202
rect 207 2198 211 2202
rect 223 2198 227 2202
rect 279 2198 283 2202
rect 335 2198 339 2202
rect 359 2198 363 2202
rect 407 2198 411 2202
rect 439 2198 443 2202
rect 479 2198 483 2202
rect 519 2198 523 2202
rect 631 2266 635 2270
rect 647 2266 651 2270
rect 751 2342 755 2346
rect 783 2342 787 2346
rect 823 2342 827 2346
rect 855 2342 859 2346
rect 895 2342 899 2346
rect 919 2342 923 2346
rect 967 2342 971 2346
rect 991 2342 995 2346
rect 1063 2342 1067 2346
rect 1239 2342 1243 2346
rect 1279 2346 1283 2350
rect 1327 2346 1331 2350
rect 1375 2346 1379 2350
rect 1383 2346 1387 2350
rect 1415 2346 1419 2350
rect 1439 2346 1443 2350
rect 1455 2346 1459 2350
rect 1503 2346 1507 2350
rect 1559 2346 1563 2350
rect 1575 2346 1579 2350
rect 1615 2346 1619 2350
rect 1647 2346 1651 2350
rect 711 2266 715 2270
rect 727 2266 731 2270
rect 783 2266 787 2270
rect 807 2266 811 2270
rect 855 2266 859 2270
rect 887 2266 891 2270
rect 919 2266 923 2270
rect 967 2266 971 2270
rect 991 2266 995 2270
rect 1279 2278 1283 2282
rect 1327 2278 1331 2282
rect 1335 2278 1339 2282
rect 1047 2266 1051 2270
rect 1063 2266 1067 2270
rect 1127 2266 1131 2270
rect 1239 2266 1243 2270
rect 1679 2346 1683 2350
rect 1719 2346 1723 2350
rect 1735 2346 1739 2350
rect 1799 2346 1803 2350
rect 1871 2346 1875 2350
rect 1879 2346 1883 2350
rect 2047 2418 2051 2422
rect 2063 2418 2067 2422
rect 2151 2418 2155 2422
rect 2167 2418 2171 2422
rect 2263 2418 2267 2422
rect 2271 2418 2275 2422
rect 2359 2418 2363 2422
rect 2407 2418 2411 2422
rect 1951 2346 1955 2350
rect 1967 2346 1971 2350
rect 2047 2346 2051 2350
rect 2063 2346 2067 2350
rect 2151 2346 2155 2350
rect 2167 2346 2171 2350
rect 1383 2278 1387 2282
rect 1407 2278 1411 2282
rect 1439 2278 1443 2282
rect 1487 2278 1491 2282
rect 1503 2278 1507 2282
rect 1559 2278 1563 2282
rect 1575 2278 1579 2282
rect 1631 2278 1635 2282
rect 1647 2278 1651 2282
rect 1703 2278 1707 2282
rect 1719 2278 1723 2282
rect 1775 2278 1779 2282
rect 559 2198 563 2202
rect 599 2198 603 2202
rect 647 2198 651 2202
rect 679 2198 683 2202
rect 727 2198 731 2202
rect 759 2198 763 2202
rect 807 2198 811 2202
rect 831 2198 835 2202
rect 111 2122 115 2126
rect 135 2122 139 2126
rect 191 2122 195 2126
rect 207 2122 211 2126
rect 271 2122 275 2126
rect 279 2122 283 2126
rect 343 2122 347 2126
rect 359 2122 363 2126
rect 415 2122 419 2126
rect 439 2122 443 2126
rect 479 2122 483 2126
rect 519 2122 523 2126
rect 543 2122 547 2126
rect 599 2122 603 2126
rect 607 2122 611 2126
rect 671 2122 675 2126
rect 679 2122 683 2126
rect 735 2122 739 2126
rect 887 2198 891 2202
rect 903 2198 907 2202
rect 967 2198 971 2202
rect 975 2198 979 2202
rect 1047 2198 1051 2202
rect 1119 2198 1123 2202
rect 1127 2198 1131 2202
rect 1239 2198 1243 2202
rect 1279 2202 1283 2206
rect 1335 2202 1339 2206
rect 1375 2202 1379 2206
rect 1407 2202 1411 2206
rect 1439 2202 1443 2206
rect 1487 2202 1491 2206
rect 1511 2202 1515 2206
rect 759 2122 763 2126
rect 791 2122 795 2126
rect 831 2122 835 2126
rect 839 2122 843 2126
rect 887 2122 891 2126
rect 903 2122 907 2126
rect 935 2122 939 2126
rect 975 2122 979 2126
rect 991 2122 995 2126
rect 1047 2122 1051 2126
rect 111 2050 115 2054
rect 135 2050 139 2054
rect 175 2050 179 2054
rect 191 2050 195 2054
rect 215 2050 219 2054
rect 271 2050 275 2054
rect 279 2050 283 2054
rect 343 2050 347 2054
rect 351 2050 355 2054
rect 415 2050 419 2054
rect 423 2050 427 2054
rect 479 2050 483 2054
rect 487 2050 491 2054
rect 543 2050 547 2054
rect 551 2050 555 2054
rect 607 2050 611 2054
rect 615 2050 619 2054
rect 671 2050 675 2054
rect 679 2050 683 2054
rect 111 1982 115 1986
rect 135 1982 139 1986
rect 175 1982 179 1986
rect 215 1982 219 1986
rect 271 1982 275 1986
rect 279 1982 283 1986
rect 343 1982 347 1986
rect 351 1982 355 1986
rect 415 1982 419 1986
rect 423 1982 427 1986
rect 1279 2134 1283 2138
rect 1375 2134 1379 2138
rect 1399 2134 1403 2138
rect 1119 2122 1123 2126
rect 1239 2122 1243 2126
rect 1559 2202 1563 2206
rect 1591 2202 1595 2206
rect 1799 2278 1803 2282
rect 1839 2278 1843 2282
rect 1879 2278 1883 2282
rect 1911 2278 1915 2282
rect 1967 2278 1971 2282
rect 2263 2346 2267 2350
rect 2271 2346 2275 2350
rect 2359 2346 2363 2350
rect 2407 2346 2411 2350
rect 1991 2278 1995 2282
rect 2063 2278 2067 2282
rect 2079 2278 2083 2282
rect 2167 2278 2171 2282
rect 2175 2278 2179 2282
rect 2271 2278 2275 2282
rect 2279 2278 2283 2282
rect 2359 2278 2363 2282
rect 2407 2278 2411 2282
rect 1631 2202 1635 2206
rect 1671 2202 1675 2206
rect 1703 2202 1707 2206
rect 1751 2202 1755 2206
rect 1775 2202 1779 2206
rect 1831 2202 1835 2206
rect 1839 2202 1843 2206
rect 1903 2202 1907 2206
rect 1911 2202 1915 2206
rect 1967 2202 1971 2206
rect 1991 2202 1995 2206
rect 2031 2202 2035 2206
rect 2079 2202 2083 2206
rect 2095 2202 2099 2206
rect 2167 2202 2171 2206
rect 2175 2202 2179 2206
rect 2239 2202 2243 2206
rect 2279 2202 2283 2206
rect 2311 2202 2315 2206
rect 2359 2202 2363 2206
rect 1439 2134 1443 2138
rect 1495 2134 1499 2138
rect 1511 2134 1515 2138
rect 1567 2134 1571 2138
rect 1591 2134 1595 2138
rect 1647 2134 1651 2138
rect 1671 2134 1675 2138
rect 1735 2134 1739 2138
rect 1751 2134 1755 2138
rect 1823 2134 1827 2138
rect 1831 2134 1835 2138
rect 1903 2134 1907 2138
rect 1911 2134 1915 2138
rect 1967 2134 1971 2138
rect 1999 2134 2003 2138
rect 2031 2134 2035 2138
rect 2087 2134 2091 2138
rect 2095 2134 2099 2138
rect 2167 2134 2171 2138
rect 2175 2134 2179 2138
rect 2239 2134 2243 2138
rect 2407 2202 2411 2206
rect 2271 2134 2275 2138
rect 2311 2134 2315 2138
rect 1939 2112 1943 2116
rect 2251 2112 2255 2116
rect 2359 2134 2363 2138
rect 2407 2134 2411 2138
rect 1279 2066 1283 2070
rect 1399 2066 1403 2070
rect 1439 2066 1443 2070
rect 1495 2066 1499 2070
rect 1567 2066 1571 2070
rect 1647 2066 1651 2070
rect 1735 2066 1739 2070
rect 1823 2066 1827 2070
rect 1911 2066 1915 2070
rect 1999 2066 2003 2070
rect 2039 2066 2043 2070
rect 2079 2066 2083 2070
rect 2087 2066 2091 2070
rect 2119 2066 2123 2070
rect 735 2050 739 2054
rect 743 2050 747 2054
rect 791 2050 795 2054
rect 815 2050 819 2054
rect 839 2050 843 2054
rect 887 2050 891 2054
rect 935 2050 939 2054
rect 991 2050 995 2054
rect 1047 2050 1051 2054
rect 1239 2050 1243 2054
rect 487 1982 491 1986
rect 495 1982 499 1986
rect 551 1982 555 1986
rect 575 1982 579 1986
rect 615 1982 619 1986
rect 647 1982 651 1986
rect 679 1982 683 1986
rect 719 1982 723 1986
rect 743 1982 747 1986
rect 791 1982 795 1986
rect 815 1982 819 1986
rect 111 1910 115 1914
rect 135 1910 139 1914
rect 175 1910 179 1914
rect 215 1910 219 1914
rect 247 1910 251 1914
rect 271 1910 275 1914
rect 287 1910 291 1914
rect 327 1910 331 1914
rect 343 1910 347 1914
rect 367 1910 371 1914
rect 415 1910 419 1914
rect 471 1910 475 1914
rect 495 1910 499 1914
rect 535 1910 539 1914
rect 575 1910 579 1914
rect 599 1910 603 1914
rect 647 1910 651 1914
rect 663 1910 667 1914
rect 1279 1998 1283 2002
rect 1399 1998 1403 2002
rect 1439 1998 1443 2002
rect 1479 1998 1483 2002
rect 1519 1998 1523 2002
rect 1559 1998 1563 2002
rect 1599 1998 1603 2002
rect 1639 1998 1643 2002
rect 1679 1998 1683 2002
rect 1719 1998 1723 2002
rect 1767 1998 1771 2002
rect 1823 1998 1827 2002
rect 1871 1998 1875 2002
rect 1919 1998 1923 2002
rect 863 1982 867 1986
rect 935 1982 939 1986
rect 1007 1982 1011 1986
rect 1239 1982 1243 1986
rect 2159 2066 2163 2070
rect 2175 2066 2179 2070
rect 2199 2066 2203 2070
rect 2239 2066 2243 2070
rect 2271 2066 2275 2070
rect 2279 2066 2283 2070
rect 2319 2066 2323 2070
rect 2359 2066 2363 2070
rect 2407 2066 2411 2070
rect 1967 1998 1971 2002
rect 2015 1998 2019 2002
rect 2039 1998 2043 2002
rect 2055 1998 2059 2002
rect 2079 1998 2083 2002
rect 2095 1998 2099 2002
rect 2119 1998 2123 2002
rect 2143 1998 2147 2002
rect 2159 1998 2163 2002
rect 2191 1998 2195 2002
rect 2199 1998 2203 2002
rect 719 1910 723 1914
rect 727 1910 731 1914
rect 791 1910 795 1914
rect 855 1910 859 1914
rect 863 1910 867 1914
rect 919 1910 923 1914
rect 935 1910 939 1914
rect 983 1910 987 1914
rect 1007 1910 1011 1914
rect 111 1838 115 1842
rect 247 1838 251 1842
rect 287 1838 291 1842
rect 327 1838 331 1842
rect 367 1838 371 1842
rect 399 1838 403 1842
rect 415 1838 419 1842
rect 439 1838 443 1842
rect 471 1838 475 1842
rect 479 1838 483 1842
rect 519 1838 523 1842
rect 535 1838 539 1842
rect 567 1838 571 1842
rect 599 1838 603 1842
rect 1279 1926 1283 1930
rect 1343 1926 1347 1930
rect 1383 1926 1387 1930
rect 1399 1926 1403 1930
rect 1423 1926 1427 1930
rect 1439 1926 1443 1930
rect 1463 1926 1467 1930
rect 1479 1926 1483 1930
rect 1511 1926 1515 1930
rect 1519 1926 1523 1930
rect 1055 1910 1059 1914
rect 1127 1910 1131 1914
rect 1239 1910 1243 1914
rect 623 1838 627 1842
rect 663 1838 667 1842
rect 687 1838 691 1842
rect 727 1838 731 1842
rect 759 1838 763 1842
rect 791 1838 795 1842
rect 831 1838 835 1842
rect 855 1838 859 1842
rect 903 1838 907 1842
rect 919 1838 923 1842
rect 975 1838 979 1842
rect 983 1838 987 1842
rect 1047 1838 1051 1842
rect 1055 1838 1059 1842
rect 111 1770 115 1774
rect 399 1770 403 1774
rect 407 1770 411 1774
rect 439 1770 443 1774
rect 447 1770 451 1774
rect 479 1770 483 1774
rect 487 1770 491 1774
rect 519 1770 523 1774
rect 527 1770 531 1774
rect 567 1770 571 1774
rect 607 1770 611 1774
rect 623 1770 627 1774
rect 647 1770 651 1774
rect 111 1698 115 1702
rect 279 1698 283 1702
rect 319 1698 323 1702
rect 359 1698 363 1702
rect 399 1698 403 1702
rect 407 1698 411 1702
rect 687 1770 691 1774
rect 695 1770 699 1774
rect 751 1770 755 1774
rect 759 1770 763 1774
rect 807 1770 811 1774
rect 831 1770 835 1774
rect 871 1770 875 1774
rect 903 1770 907 1774
rect 935 1770 939 1774
rect 1279 1850 1283 1854
rect 1343 1850 1347 1854
rect 1359 1850 1363 1854
rect 1127 1838 1131 1842
rect 1191 1838 1195 1842
rect 1239 1838 1243 1842
rect 1559 1926 1563 1930
rect 1567 1926 1571 1930
rect 1599 1926 1603 1930
rect 1631 1926 1635 1930
rect 1639 1926 1643 1930
rect 1679 1926 1683 1930
rect 1711 1926 1715 1930
rect 1719 1926 1723 1930
rect 1767 1926 1771 1930
rect 1807 1926 1811 1930
rect 1823 1926 1827 1930
rect 1871 1926 1875 1930
rect 1919 1926 1923 1930
rect 1967 1926 1971 1930
rect 2015 1926 2019 1930
rect 2031 1926 2035 1930
rect 2055 1926 2059 1930
rect 2239 1998 2243 2002
rect 2279 1998 2283 2002
rect 2319 1998 2323 2002
rect 2359 1998 2363 2002
rect 2407 1998 2411 2002
rect 2095 1926 2099 1930
rect 2143 1926 2147 1930
rect 2151 1926 2155 1930
rect 2191 1926 2195 1930
rect 2239 1926 2243 1930
rect 2279 1926 2283 1930
rect 2319 1926 2323 1930
rect 2359 1926 2363 1930
rect 2407 1926 2411 1930
rect 1383 1850 1387 1854
rect 1399 1850 1403 1854
rect 1423 1850 1427 1854
rect 1447 1850 1451 1854
rect 1463 1850 1467 1854
rect 1503 1850 1507 1854
rect 1511 1850 1515 1854
rect 1559 1850 1563 1854
rect 1567 1850 1571 1854
rect 1615 1850 1619 1854
rect 1631 1850 1635 1854
rect 1671 1850 1675 1854
rect 1711 1850 1715 1854
rect 1727 1850 1731 1854
rect 1783 1850 1787 1854
rect 1807 1850 1811 1854
rect 1839 1850 1843 1854
rect 1895 1850 1899 1854
rect 1919 1850 1923 1854
rect 1951 1850 1955 1854
rect 2031 1850 2035 1854
rect 2151 1850 2155 1854
rect 2407 1850 2411 1854
rect 975 1770 979 1774
rect 999 1770 1003 1774
rect 1047 1770 1051 1774
rect 1071 1770 1075 1774
rect 1127 1770 1131 1774
rect 1143 1770 1147 1774
rect 1191 1770 1195 1774
rect 1239 1770 1243 1774
rect 1279 1770 1283 1774
rect 1303 1770 1307 1774
rect 1343 1770 1347 1774
rect 1359 1770 1363 1774
rect 1391 1770 1395 1774
rect 1399 1770 1403 1774
rect 1447 1770 1451 1774
rect 1455 1770 1459 1774
rect 1503 1770 1507 1774
rect 1519 1770 1523 1774
rect 1559 1770 1563 1774
rect 1583 1770 1587 1774
rect 447 1698 451 1702
rect 487 1698 491 1702
rect 495 1698 499 1702
rect 527 1698 531 1702
rect 543 1698 547 1702
rect 567 1698 571 1702
rect 591 1698 595 1702
rect 607 1698 611 1702
rect 639 1698 643 1702
rect 647 1698 651 1702
rect 687 1698 691 1702
rect 695 1698 699 1702
rect 735 1698 739 1702
rect 751 1698 755 1702
rect 783 1698 787 1702
rect 807 1698 811 1702
rect 839 1698 843 1702
rect 871 1698 875 1702
rect 895 1698 899 1702
rect 935 1698 939 1702
rect 999 1698 1003 1702
rect 1071 1698 1075 1702
rect 1143 1698 1147 1702
rect 1191 1698 1195 1702
rect 1239 1698 1243 1702
rect 1279 1698 1283 1702
rect 1303 1698 1307 1702
rect 1343 1698 1347 1702
rect 111 1626 115 1630
rect 135 1626 139 1630
rect 175 1626 179 1630
rect 215 1626 219 1630
rect 255 1626 259 1630
rect 279 1626 283 1630
rect 311 1626 315 1630
rect 319 1626 323 1630
rect 359 1626 363 1630
rect 391 1626 395 1630
rect 399 1626 403 1630
rect 111 1554 115 1558
rect 135 1554 139 1558
rect 151 1554 155 1558
rect 175 1554 179 1558
rect 447 1626 451 1630
rect 471 1626 475 1630
rect 495 1626 499 1630
rect 543 1626 547 1630
rect 559 1626 563 1630
rect 591 1626 595 1630
rect 639 1626 643 1630
rect 687 1626 691 1630
rect 719 1626 723 1630
rect 735 1626 739 1630
rect 783 1626 787 1630
rect 791 1626 795 1630
rect 1383 1698 1387 1702
rect 1391 1698 1395 1702
rect 1423 1698 1427 1702
rect 1455 1698 1459 1702
rect 1463 1698 1467 1702
rect 1503 1698 1507 1702
rect 1519 1698 1523 1702
rect 1559 1698 1563 1702
rect 1583 1698 1587 1702
rect 1615 1770 1619 1774
rect 1647 1770 1651 1774
rect 1671 1770 1675 1774
rect 1703 1770 1707 1774
rect 1727 1770 1731 1774
rect 1759 1770 1763 1774
rect 1783 1770 1787 1774
rect 1807 1770 1811 1774
rect 1839 1770 1843 1774
rect 1863 1770 1867 1774
rect 1895 1770 1899 1774
rect 1919 1770 1923 1774
rect 1951 1770 1955 1774
rect 1975 1770 1979 1774
rect 2407 1770 2411 1774
rect 1623 1698 1627 1702
rect 1647 1698 1651 1702
rect 1687 1698 1691 1702
rect 1703 1698 1707 1702
rect 1751 1698 1755 1702
rect 1759 1698 1763 1702
rect 1807 1698 1811 1702
rect 1863 1698 1867 1702
rect 1919 1698 1923 1702
rect 1975 1698 1979 1702
rect 2031 1698 2035 1702
rect 2087 1698 2091 1702
rect 2407 1698 2411 1702
rect 839 1626 843 1630
rect 855 1626 859 1630
rect 895 1626 899 1630
rect 919 1626 923 1630
rect 983 1626 987 1630
rect 1047 1626 1051 1630
rect 1239 1626 1243 1630
rect 1279 1626 1283 1630
rect 1303 1626 1307 1630
rect 1343 1626 1347 1630
rect 1383 1626 1387 1630
rect 1423 1626 1427 1630
rect 1463 1626 1467 1630
rect 1503 1626 1507 1630
rect 1559 1626 1563 1630
rect 1623 1626 1627 1630
rect 1631 1626 1635 1630
rect 1687 1626 1691 1630
rect 1703 1626 1707 1630
rect 1751 1626 1755 1630
rect 1783 1626 1787 1630
rect 1807 1626 1811 1630
rect 1855 1626 1859 1630
rect 1863 1626 1867 1630
rect 1919 1626 1923 1630
rect 1927 1626 1931 1630
rect 199 1554 203 1558
rect 215 1554 219 1558
rect 255 1554 259 1558
rect 263 1554 267 1558
rect 311 1554 315 1558
rect 343 1554 347 1558
rect 391 1554 395 1558
rect 439 1554 443 1558
rect 471 1554 475 1558
rect 535 1554 539 1558
rect 559 1554 563 1558
rect 639 1554 643 1558
rect 719 1554 723 1558
rect 735 1554 739 1558
rect 791 1554 795 1558
rect 823 1554 827 1558
rect 855 1554 859 1558
rect 903 1554 907 1558
rect 919 1554 923 1558
rect 975 1554 979 1558
rect 983 1554 987 1558
rect 1047 1554 1051 1558
rect 1119 1554 1123 1558
rect 1191 1554 1195 1558
rect 1239 1554 1243 1558
rect 1279 1558 1283 1562
rect 1303 1558 1307 1562
rect 1343 1558 1347 1562
rect 1383 1558 1387 1562
rect 1423 1558 1427 1562
rect 1463 1558 1467 1562
rect 1471 1558 1475 1562
rect 1503 1558 1507 1562
rect 111 1482 115 1486
rect 151 1482 155 1486
rect 199 1482 203 1486
rect 263 1482 267 1486
rect 319 1482 323 1486
rect 343 1482 347 1486
rect 359 1482 363 1486
rect 399 1482 403 1486
rect 439 1482 443 1486
rect 447 1482 451 1486
rect 503 1482 507 1486
rect 535 1482 539 1486
rect 559 1482 563 1486
rect 615 1482 619 1486
rect 639 1482 643 1486
rect 671 1482 675 1486
rect 735 1482 739 1486
rect 799 1482 803 1486
rect 823 1482 827 1486
rect 855 1482 859 1486
rect 903 1482 907 1486
rect 911 1482 915 1486
rect 967 1482 971 1486
rect 975 1482 979 1486
rect 1023 1482 1027 1486
rect 1047 1482 1051 1486
rect 1087 1482 1091 1486
rect 1119 1482 1123 1486
rect 1151 1482 1155 1486
rect 111 1410 115 1414
rect 263 1410 267 1414
rect 303 1410 307 1414
rect 319 1410 323 1414
rect 343 1410 347 1414
rect 359 1410 363 1414
rect 391 1410 395 1414
rect 399 1410 403 1414
rect 447 1410 451 1414
rect 503 1410 507 1414
rect 559 1410 563 1414
rect 615 1410 619 1414
rect 623 1410 627 1414
rect 1191 1482 1195 1486
rect 1239 1482 1243 1486
rect 671 1410 675 1414
rect 687 1410 691 1414
rect 735 1410 739 1414
rect 751 1410 755 1414
rect 799 1410 803 1414
rect 815 1410 819 1414
rect 111 1338 115 1342
rect 135 1338 139 1342
rect 175 1338 179 1342
rect 215 1338 219 1342
rect 255 1338 259 1342
rect 263 1338 267 1342
rect 303 1338 307 1342
rect 327 1338 331 1342
rect 343 1338 347 1342
rect 111 1266 115 1270
rect 135 1266 139 1270
rect 175 1266 179 1270
rect 215 1266 219 1270
rect 391 1338 395 1342
rect 407 1338 411 1342
rect 447 1338 451 1342
rect 495 1338 499 1342
rect 503 1338 507 1342
rect 559 1338 563 1342
rect 583 1338 587 1342
rect 623 1338 627 1342
rect 671 1338 675 1342
rect 687 1338 691 1342
rect 751 1338 755 1342
rect 759 1338 763 1342
rect 855 1410 859 1414
rect 879 1410 883 1414
rect 911 1410 915 1414
rect 951 1410 955 1414
rect 967 1410 971 1414
rect 1559 1558 1563 1562
rect 1623 1558 1627 1562
rect 1631 1558 1635 1562
rect 1703 1558 1707 1562
rect 1759 1558 1763 1562
rect 1783 1558 1787 1562
rect 1975 1626 1979 1630
rect 1999 1626 2003 1630
rect 2031 1626 2035 1630
rect 2063 1626 2067 1630
rect 2087 1626 2091 1630
rect 2127 1626 2131 1630
rect 2191 1626 2195 1630
rect 2255 1626 2259 1630
rect 2319 1626 2323 1630
rect 2359 1626 2363 1630
rect 2407 1626 2411 1630
rect 1855 1558 1859 1562
rect 1871 1558 1875 1562
rect 1927 1558 1931 1562
rect 1967 1558 1971 1562
rect 1999 1558 2003 1562
rect 2055 1558 2059 1562
rect 2063 1558 2067 1562
rect 2127 1558 2131 1562
rect 2191 1558 2195 1562
rect 2255 1558 2259 1562
rect 2319 1558 2323 1562
rect 2359 1558 2363 1562
rect 2407 1558 2411 1562
rect 1279 1470 1283 1474
rect 1303 1470 1307 1474
rect 1375 1470 1379 1474
rect 1471 1470 1475 1474
rect 1479 1470 1483 1474
rect 1583 1470 1587 1474
rect 1623 1470 1627 1474
rect 1687 1470 1691 1474
rect 1759 1470 1763 1474
rect 1783 1470 1787 1474
rect 1871 1470 1875 1474
rect 1951 1470 1955 1474
rect 1967 1470 1971 1474
rect 2031 1470 2035 1474
rect 2055 1470 2059 1474
rect 2103 1470 2107 1474
rect 2127 1470 2131 1474
rect 2167 1470 2171 1474
rect 2191 1470 2195 1474
rect 2239 1470 2243 1474
rect 2255 1470 2259 1474
rect 2311 1470 2315 1474
rect 2319 1470 2323 1474
rect 2359 1470 2363 1474
rect 2407 1470 2411 1474
rect 1023 1410 1027 1414
rect 1087 1410 1091 1414
rect 1151 1410 1155 1414
rect 1191 1410 1195 1414
rect 1239 1410 1243 1414
rect 1279 1402 1283 1406
rect 1303 1402 1307 1406
rect 1343 1402 1347 1406
rect 1375 1402 1379 1406
rect 1399 1402 1403 1406
rect 815 1338 819 1342
rect 839 1338 843 1342
rect 879 1338 883 1342
rect 919 1338 923 1342
rect 951 1338 955 1342
rect 1007 1338 1011 1342
rect 1023 1338 1027 1342
rect 1095 1338 1099 1342
rect 1239 1338 1243 1342
rect 247 1266 251 1270
rect 255 1266 259 1270
rect 327 1266 331 1270
rect 407 1266 411 1270
rect 415 1266 419 1270
rect 495 1266 499 1270
rect 503 1266 507 1270
rect 583 1266 587 1270
rect 591 1266 595 1270
rect 671 1266 675 1270
rect 743 1266 747 1270
rect 759 1266 763 1270
rect 815 1266 819 1270
rect 839 1266 843 1270
rect 879 1266 883 1270
rect 919 1266 923 1270
rect 943 1266 947 1270
rect 1007 1266 1011 1270
rect 1071 1266 1075 1270
rect 1095 1266 1099 1270
rect 1471 1402 1475 1406
rect 1479 1402 1483 1406
rect 1551 1402 1555 1406
rect 1583 1402 1587 1406
rect 1639 1402 1643 1406
rect 1687 1402 1691 1406
rect 1727 1402 1731 1406
rect 1783 1402 1787 1406
rect 1815 1402 1819 1406
rect 1871 1402 1875 1406
rect 1903 1402 1907 1406
rect 1951 1402 1955 1406
rect 1991 1402 1995 1406
rect 2031 1402 2035 1406
rect 2071 1402 2075 1406
rect 1279 1330 1283 1334
rect 1303 1330 1307 1334
rect 1343 1330 1347 1334
rect 1399 1330 1403 1334
rect 1447 1330 1451 1334
rect 1471 1330 1475 1334
rect 1487 1330 1491 1334
rect 1527 1330 1531 1334
rect 1551 1330 1555 1334
rect 1567 1330 1571 1334
rect 2103 1402 2107 1406
rect 2151 1402 2155 1406
rect 2167 1402 2171 1406
rect 2223 1402 2227 1406
rect 2239 1402 2243 1406
rect 2303 1402 2307 1406
rect 2311 1402 2315 1406
rect 2359 1402 2363 1406
rect 2407 1402 2411 1406
rect 1615 1330 1619 1334
rect 1639 1330 1643 1334
rect 1671 1330 1675 1334
rect 1719 1330 1723 1334
rect 1727 1330 1731 1334
rect 1775 1330 1779 1334
rect 1815 1330 1819 1334
rect 1831 1330 1835 1334
rect 1903 1330 1907 1334
rect 1983 1330 1987 1334
rect 1991 1330 1995 1334
rect 2071 1330 2075 1334
rect 2151 1330 2155 1334
rect 2167 1330 2171 1334
rect 2223 1330 2227 1334
rect 2271 1330 2275 1334
rect 1239 1266 1243 1270
rect 1279 1258 1283 1262
rect 1447 1258 1451 1262
rect 1487 1258 1491 1262
rect 1511 1258 1515 1262
rect 1527 1258 1531 1262
rect 1551 1258 1555 1262
rect 1567 1258 1571 1262
rect 1591 1258 1595 1262
rect 1615 1258 1619 1262
rect 111 1190 115 1194
rect 135 1190 139 1194
rect 175 1190 179 1194
rect 231 1190 235 1194
rect 247 1190 251 1194
rect 303 1190 307 1194
rect 327 1190 331 1194
rect 383 1190 387 1194
rect 415 1190 419 1194
rect 471 1190 475 1194
rect 503 1190 507 1194
rect 559 1190 563 1194
rect 591 1190 595 1194
rect 639 1190 643 1194
rect 671 1190 675 1194
rect 111 1122 115 1126
rect 135 1122 139 1126
rect 175 1122 179 1126
rect 215 1122 219 1126
rect 231 1122 235 1126
rect 303 1122 307 1126
rect 383 1122 387 1126
rect 391 1122 395 1126
rect 719 1190 723 1194
rect 743 1190 747 1194
rect 799 1190 803 1194
rect 815 1190 819 1194
rect 871 1190 875 1194
rect 879 1190 883 1194
rect 471 1122 475 1126
rect 479 1122 483 1126
rect 559 1122 563 1126
rect 639 1122 643 1126
rect 711 1122 715 1126
rect 719 1122 723 1126
rect 935 1190 939 1194
rect 943 1190 947 1194
rect 991 1190 995 1194
rect 1007 1190 1011 1194
rect 1047 1190 1051 1194
rect 1071 1190 1075 1194
rect 1103 1190 1107 1194
rect 1151 1190 1155 1194
rect 1191 1190 1195 1194
rect 1239 1190 1243 1194
rect 1631 1258 1635 1262
rect 1671 1258 1675 1262
rect 1711 1258 1715 1262
rect 1719 1258 1723 1262
rect 1751 1258 1755 1262
rect 1775 1258 1779 1262
rect 1791 1258 1795 1262
rect 1831 1258 1835 1262
rect 1839 1258 1843 1262
rect 1903 1258 1907 1262
rect 1967 1258 1971 1262
rect 1983 1258 1987 1262
rect 2039 1258 2043 1262
rect 2071 1258 2075 1262
rect 2119 1258 2123 1262
rect 775 1122 779 1126
rect 799 1122 803 1126
rect 839 1122 843 1126
rect 871 1122 875 1126
rect 903 1122 907 1126
rect 935 1122 939 1126
rect 959 1122 963 1126
rect 991 1122 995 1126
rect 111 1050 115 1054
rect 135 1050 139 1054
rect 199 1050 203 1054
rect 215 1050 219 1054
rect 239 1050 243 1054
rect 287 1050 291 1054
rect 303 1050 307 1054
rect 343 1050 347 1054
rect 391 1050 395 1054
rect 439 1050 443 1054
rect 479 1050 483 1054
rect 487 1050 491 1054
rect 535 1050 539 1054
rect 559 1050 563 1054
rect 111 970 115 974
rect 199 970 203 974
rect 239 970 243 974
rect 287 970 291 974
rect 295 970 299 974
rect 343 970 347 974
rect 391 970 395 974
rect 399 970 403 974
rect 583 1050 587 1054
rect 631 1050 635 1054
rect 639 1050 643 1054
rect 679 1050 683 1054
rect 711 1050 715 1054
rect 727 1050 731 1054
rect 775 1050 779 1054
rect 783 1050 787 1054
rect 839 1050 843 1054
rect 895 1050 899 1054
rect 903 1050 907 1054
rect 959 1050 963 1054
rect 1023 1122 1027 1126
rect 1047 1122 1051 1126
rect 1087 1122 1091 1126
rect 1103 1122 1107 1126
rect 1151 1122 1155 1126
rect 1191 1122 1195 1126
rect 1279 1186 1283 1190
rect 1511 1186 1515 1190
rect 1551 1186 1555 1190
rect 1559 1186 1563 1190
rect 1591 1186 1595 1190
rect 1599 1186 1603 1190
rect 1631 1186 1635 1190
rect 1639 1186 1643 1190
rect 1671 1186 1675 1190
rect 1679 1186 1683 1190
rect 1711 1186 1715 1190
rect 1719 1186 1723 1190
rect 1751 1186 1755 1190
rect 1759 1186 1763 1190
rect 1791 1186 1795 1190
rect 1799 1186 1803 1190
rect 2167 1258 2171 1262
rect 2207 1258 2211 1262
rect 2271 1258 2275 1262
rect 2303 1330 2307 1334
rect 2359 1330 2363 1334
rect 2407 1330 2411 1334
rect 2295 1258 2299 1262
rect 2359 1258 2363 1262
rect 1839 1186 1843 1190
rect 1855 1186 1859 1190
rect 1903 1186 1907 1190
rect 1927 1186 1931 1190
rect 1967 1186 1971 1190
rect 2023 1186 2027 1190
rect 2039 1186 2043 1190
rect 2119 1186 2123 1190
rect 2135 1186 2139 1190
rect 2207 1186 2211 1190
rect 1239 1122 1243 1126
rect 1279 1110 1283 1114
rect 1535 1110 1539 1114
rect 1559 1110 1563 1114
rect 1599 1110 1603 1114
rect 1639 1110 1643 1114
rect 1663 1110 1667 1114
rect 1679 1110 1683 1114
rect 1719 1110 1723 1114
rect 1727 1110 1731 1114
rect 1023 1050 1027 1054
rect 1087 1050 1091 1054
rect 1151 1050 1155 1054
rect 1191 1050 1195 1054
rect 439 970 443 974
rect 471 970 475 974
rect 487 970 491 974
rect 535 970 539 974
rect 551 970 555 974
rect 583 970 587 974
rect 631 970 635 974
rect 639 970 643 974
rect 679 970 683 974
rect 727 970 731 974
rect 783 970 787 974
rect 807 970 811 974
rect 839 970 843 974
rect 887 970 891 974
rect 895 970 899 974
rect 959 970 963 974
rect 1023 970 1027 974
rect 1087 970 1091 974
rect 1239 1050 1243 1054
rect 1759 1110 1763 1114
rect 1791 1110 1795 1114
rect 1799 1110 1803 1114
rect 1855 1110 1859 1114
rect 1911 1110 1915 1114
rect 1927 1110 1931 1114
rect 1967 1110 1971 1114
rect 1279 1030 1283 1034
rect 1503 1030 1507 1034
rect 1535 1030 1539 1034
rect 1599 1030 1603 1034
rect 1623 1030 1627 1034
rect 1663 1030 1667 1034
rect 1727 1030 1731 1034
rect 1735 1030 1739 1034
rect 2023 1110 2027 1114
rect 2079 1110 2083 1114
rect 2135 1110 2139 1114
rect 2191 1110 2195 1114
rect 2255 1186 2259 1190
rect 2295 1186 2299 1190
rect 2407 1258 2411 1262
rect 2359 1186 2363 1190
rect 2407 1186 2411 1190
rect 2255 1110 2259 1114
rect 2319 1110 2323 1114
rect 2359 1110 2363 1114
rect 1791 1030 1795 1034
rect 1831 1030 1835 1034
rect 1855 1030 1859 1034
rect 1911 1030 1915 1034
rect 1919 1030 1923 1034
rect 1967 1030 1971 1034
rect 1999 1030 2003 1034
rect 2023 1030 2027 1034
rect 2407 1110 2411 1114
rect 2071 1030 2075 1034
rect 2079 1030 2083 1034
rect 2135 1030 2139 1034
rect 2143 1030 2147 1034
rect 2191 1030 2195 1034
rect 2207 1030 2211 1034
rect 2255 1030 2259 1034
rect 2279 1030 2283 1034
rect 2319 1030 2323 1034
rect 2359 1030 2363 1034
rect 2407 1030 2411 1034
rect 1151 970 1155 974
rect 1191 970 1195 974
rect 1239 970 1243 974
rect 1279 954 1283 958
rect 1319 954 1323 958
rect 1359 954 1363 958
rect 1399 954 1403 958
rect 1463 954 1467 958
rect 1503 954 1507 958
rect 1543 954 1547 958
rect 1623 954 1627 958
rect 1639 954 1643 958
rect 1735 954 1739 958
rect 1831 954 1835 958
rect 1839 954 1843 958
rect 1919 954 1923 958
rect 1935 954 1939 958
rect 1999 954 2003 958
rect 2023 954 2027 958
rect 2071 954 2075 958
rect 2103 954 2107 958
rect 111 894 115 898
rect 255 894 259 898
rect 295 894 299 898
rect 311 894 315 898
rect 343 894 347 898
rect 375 894 379 898
rect 399 894 403 898
rect 455 894 459 898
rect 471 894 475 898
rect 535 894 539 898
rect 551 894 555 898
rect 111 826 115 830
rect 191 826 195 830
rect 247 826 251 830
rect 255 826 259 830
rect 311 826 315 830
rect 623 894 627 898
rect 639 894 643 898
rect 711 894 715 898
rect 727 894 731 898
rect 791 894 795 898
rect 807 894 811 898
rect 863 894 867 898
rect 887 894 891 898
rect 935 894 939 898
rect 959 894 963 898
rect 999 894 1003 898
rect 1023 894 1027 898
rect 1055 894 1059 898
rect 375 826 379 830
rect 383 826 387 830
rect 455 826 459 830
rect 463 826 467 830
rect 535 826 539 830
rect 543 826 547 830
rect 615 826 619 830
rect 623 826 627 830
rect 111 758 115 762
rect 135 758 139 762
rect 175 758 179 762
rect 191 758 195 762
rect 215 758 219 762
rect 247 758 251 762
rect 279 758 283 762
rect 111 682 115 686
rect 135 682 139 686
rect 175 682 179 686
rect 311 758 315 762
rect 351 758 355 762
rect 383 758 387 762
rect 423 758 427 762
rect 463 758 467 762
rect 495 758 499 762
rect 687 826 691 830
rect 711 826 715 830
rect 751 826 755 830
rect 791 826 795 830
rect 815 826 819 830
rect 863 826 867 830
rect 871 826 875 830
rect 1087 894 1091 898
rect 1119 894 1123 898
rect 1151 894 1155 898
rect 1183 894 1187 898
rect 1191 894 1195 898
rect 1239 894 1243 898
rect 1279 878 1283 882
rect 1319 878 1323 882
rect 1335 878 1339 882
rect 1359 878 1363 882
rect 1375 878 1379 882
rect 1399 878 1403 882
rect 1415 878 1419 882
rect 1463 878 1467 882
rect 1471 878 1475 882
rect 2143 954 2147 958
rect 2175 954 2179 958
rect 2207 954 2211 958
rect 2239 954 2243 958
rect 2279 954 2283 958
rect 2311 954 2315 958
rect 2359 954 2363 958
rect 2407 954 2411 958
rect 1535 878 1539 882
rect 1543 878 1547 882
rect 1607 878 1611 882
rect 1639 878 1643 882
rect 1679 878 1683 882
rect 1735 878 1739 882
rect 1751 878 1755 882
rect 927 826 931 830
rect 935 826 939 830
rect 983 826 987 830
rect 999 826 1003 830
rect 1047 826 1051 830
rect 1055 826 1059 830
rect 1119 826 1123 830
rect 1183 826 1187 830
rect 1239 826 1243 830
rect 1279 806 1283 810
rect 1303 806 1307 810
rect 1335 806 1339 810
rect 1343 806 1347 810
rect 543 758 547 762
rect 559 758 563 762
rect 615 758 619 762
rect 623 758 627 762
rect 687 758 691 762
rect 695 758 699 762
rect 751 758 755 762
rect 783 758 787 762
rect 815 758 819 762
rect 871 758 875 762
rect 879 758 883 762
rect 215 682 219 686
rect 231 682 235 686
rect 279 682 283 686
rect 287 682 291 686
rect 343 682 347 686
rect 351 682 355 686
rect 399 682 403 686
rect 423 682 427 686
rect 455 682 459 686
rect 495 682 499 686
rect 503 682 507 686
rect 559 682 563 686
rect 623 682 627 686
rect 695 682 699 686
rect 927 758 931 762
rect 983 758 987 762
rect 1047 758 1051 762
rect 1095 758 1099 762
rect 1191 758 1195 762
rect 1239 758 1243 762
rect 1375 806 1379 810
rect 1407 806 1411 810
rect 1415 806 1419 810
rect 1471 806 1475 810
rect 1479 806 1483 810
rect 1535 806 1539 810
rect 1551 806 1555 810
rect 1279 738 1283 742
rect 1303 738 1307 742
rect 767 682 771 686
rect 783 682 787 686
rect 839 682 843 686
rect 879 682 883 686
rect 903 682 907 686
rect 967 682 971 686
rect 983 682 987 686
rect 1023 682 1027 686
rect 1087 682 1091 686
rect 1095 682 1099 686
rect 1151 682 1155 686
rect 111 614 115 618
rect 135 614 139 618
rect 175 614 179 618
rect 183 614 187 618
rect 231 614 235 618
rect 255 614 259 618
rect 287 614 291 618
rect 327 614 331 618
rect 343 614 347 618
rect 399 614 403 618
rect 455 614 459 618
rect 479 614 483 618
rect 503 614 507 618
rect 111 542 115 546
rect 135 542 139 546
rect 151 542 155 546
rect 183 542 187 546
rect 223 542 227 546
rect 255 542 259 546
rect 287 542 291 546
rect 327 542 331 546
rect 559 614 563 618
rect 623 614 627 618
rect 639 614 643 618
rect 695 614 699 618
rect 719 614 723 618
rect 767 614 771 618
rect 799 614 803 618
rect 839 614 843 618
rect 879 614 883 618
rect 903 614 907 618
rect 1343 738 1347 742
rect 1367 738 1371 742
rect 1407 738 1411 742
rect 1455 738 1459 742
rect 1479 738 1483 742
rect 1607 806 1611 810
rect 1623 806 1627 810
rect 1823 878 1827 882
rect 1839 878 1843 882
rect 1895 878 1899 882
rect 1935 878 1939 882
rect 1959 878 1963 882
rect 2023 878 2027 882
rect 2087 878 2091 882
rect 2103 878 2107 882
rect 2143 878 2147 882
rect 2175 878 2179 882
rect 2199 878 2203 882
rect 2239 878 2243 882
rect 2255 878 2259 882
rect 2311 878 2315 882
rect 2319 878 2323 882
rect 2359 878 2363 882
rect 2407 878 2411 882
rect 1679 806 1683 810
rect 1695 806 1699 810
rect 1751 806 1755 810
rect 1759 806 1763 810
rect 1823 806 1827 810
rect 1887 806 1891 810
rect 1895 806 1899 810
rect 1951 806 1955 810
rect 1959 806 1963 810
rect 2023 806 2027 810
rect 1535 738 1539 742
rect 1551 738 1555 742
rect 1615 738 1619 742
rect 1623 738 1627 742
rect 1695 738 1699 742
rect 1191 682 1195 686
rect 1239 682 1243 686
rect 1279 670 1283 674
rect 1303 670 1307 674
rect 1367 670 1371 674
rect 1455 670 1459 674
rect 1535 670 1539 674
rect 1591 670 1595 674
rect 951 614 955 618
rect 967 614 971 618
rect 1015 614 1019 618
rect 1023 614 1027 618
rect 1079 614 1083 618
rect 1087 614 1091 618
rect 351 542 355 546
rect 399 542 403 546
rect 415 542 419 546
rect 479 542 483 546
rect 551 542 555 546
rect 559 542 563 546
rect 111 474 115 478
rect 151 474 155 478
rect 223 474 227 478
rect 239 474 243 478
rect 279 474 283 478
rect 287 474 291 478
rect 327 474 331 478
rect 351 474 355 478
rect 383 474 387 478
rect 415 474 419 478
rect 439 474 443 478
rect 623 542 627 546
rect 639 542 643 546
rect 695 542 699 546
rect 719 542 723 546
rect 767 542 771 546
rect 799 542 803 546
rect 1143 614 1147 618
rect 1151 614 1155 618
rect 1191 614 1195 618
rect 1239 614 1243 618
rect 1279 594 1283 598
rect 1559 594 1563 598
rect 839 542 843 546
rect 879 542 883 546
rect 919 542 923 546
rect 951 542 955 546
rect 999 542 1003 546
rect 1015 542 1019 546
rect 1079 542 1083 546
rect 479 474 483 478
rect 503 474 507 478
rect 551 474 555 478
rect 567 474 571 478
rect 623 474 627 478
rect 631 474 635 478
rect 695 474 699 478
rect 111 402 115 406
rect 143 402 147 406
rect 183 402 187 406
rect 223 402 227 406
rect 239 402 243 406
rect 271 402 275 406
rect 279 402 283 406
rect 327 402 331 406
rect 335 402 339 406
rect 383 402 387 406
rect 399 402 403 406
rect 759 474 763 478
rect 767 474 771 478
rect 823 474 827 478
rect 839 474 843 478
rect 887 474 891 478
rect 919 474 923 478
rect 951 474 955 478
rect 1615 670 1619 674
rect 1639 670 1643 674
rect 1759 738 1763 742
rect 1775 738 1779 742
rect 2087 806 2091 810
rect 2103 806 2107 810
rect 2143 806 2147 810
rect 2191 806 2195 810
rect 2199 806 2203 810
rect 2255 806 2259 810
rect 2279 806 2283 810
rect 2319 806 2323 810
rect 2359 806 2363 810
rect 1823 738 1827 742
rect 1855 738 1859 742
rect 1887 738 1891 742
rect 1943 738 1947 742
rect 1951 738 1955 742
rect 2023 738 2027 742
rect 2031 738 2035 742
rect 2103 738 2107 742
rect 2119 738 2123 742
rect 2191 738 2195 742
rect 2207 738 2211 742
rect 2279 738 2283 742
rect 2295 738 2299 742
rect 2407 806 2411 810
rect 2359 738 2363 742
rect 2407 738 2411 742
rect 1687 670 1691 674
rect 1695 670 1699 674
rect 1743 670 1747 674
rect 1775 670 1779 674
rect 1799 670 1803 674
rect 1855 670 1859 674
rect 1871 670 1875 674
rect 1943 670 1947 674
rect 1951 670 1955 674
rect 2031 670 2035 674
rect 2047 670 2051 674
rect 2119 670 2123 674
rect 1591 594 1595 598
rect 1599 594 1603 598
rect 1639 594 1643 598
rect 1679 594 1683 598
rect 1687 594 1691 598
rect 1719 594 1723 598
rect 1743 594 1747 598
rect 1759 594 1763 598
rect 1799 594 1803 598
rect 1807 594 1811 598
rect 1855 594 1859 598
rect 1871 594 1875 598
rect 1911 594 1915 598
rect 1951 594 1955 598
rect 1967 594 1971 598
rect 2151 670 2155 674
rect 2207 670 2211 674
rect 2263 670 2267 674
rect 2295 670 2299 674
rect 2359 670 2363 674
rect 2407 670 2411 674
rect 2031 594 2035 598
rect 2047 594 2051 598
rect 2095 594 2099 598
rect 2151 594 2155 598
rect 2167 594 2171 598
rect 2239 594 2243 598
rect 2263 594 2267 598
rect 2311 594 2315 598
rect 2359 594 2363 598
rect 2407 594 2411 598
rect 1143 542 1147 546
rect 1191 542 1195 546
rect 1239 542 1243 546
rect 1279 526 1283 530
rect 1407 526 1411 530
rect 1447 526 1451 530
rect 1487 526 1491 530
rect 1535 526 1539 530
rect 1559 526 1563 530
rect 1591 526 1595 530
rect 1599 526 1603 530
rect 1639 526 1643 530
rect 1647 526 1651 530
rect 1679 526 1683 530
rect 1711 526 1715 530
rect 1719 526 1723 530
rect 999 474 1003 478
rect 1015 474 1019 478
rect 1079 474 1083 478
rect 1239 474 1243 478
rect 439 402 443 406
rect 471 402 475 406
rect 503 402 507 406
rect 543 402 547 406
rect 567 402 571 406
rect 111 326 115 330
rect 135 326 139 330
rect 143 326 147 330
rect 175 326 179 330
rect 183 326 187 330
rect 111 250 115 254
rect 135 250 139 254
rect 215 326 219 330
rect 223 326 227 330
rect 255 326 259 330
rect 271 326 275 330
rect 295 326 299 330
rect 335 326 339 330
rect 391 326 395 330
rect 399 326 403 330
rect 447 326 451 330
rect 615 402 619 406
rect 631 402 635 406
rect 687 402 691 406
rect 695 402 699 406
rect 751 402 755 406
rect 759 402 763 406
rect 807 402 811 406
rect 823 402 827 406
rect 863 402 867 406
rect 887 402 891 406
rect 1759 526 1763 530
rect 1783 526 1787 530
rect 1807 526 1811 530
rect 1855 526 1859 530
rect 1863 526 1867 530
rect 1911 526 1915 530
rect 1943 526 1947 530
rect 1967 526 1971 530
rect 2023 526 2027 530
rect 2031 526 2035 530
rect 2095 526 2099 530
rect 2103 526 2107 530
rect 1279 458 1283 462
rect 1303 458 1307 462
rect 1343 458 1347 462
rect 1383 458 1387 462
rect 1407 458 1411 462
rect 1447 458 1451 462
rect 1487 458 1491 462
rect 1535 458 1539 462
rect 1591 458 1595 462
rect 1631 458 1635 462
rect 1647 458 1651 462
rect 1711 458 1715 462
rect 1735 458 1739 462
rect 919 402 923 406
rect 951 402 955 406
rect 975 402 979 406
rect 1015 402 1019 406
rect 1031 402 1035 406
rect 471 326 475 330
rect 495 326 499 330
rect 543 326 547 330
rect 591 326 595 330
rect 615 326 619 330
rect 639 326 643 330
rect 687 326 691 330
rect 735 326 739 330
rect 751 326 755 330
rect 783 326 787 330
rect 807 326 811 330
rect 839 326 843 330
rect 863 326 867 330
rect 1783 458 1787 462
rect 1831 458 1835 462
rect 1863 458 1867 462
rect 1919 458 1923 462
rect 1943 458 1947 462
rect 1999 458 2003 462
rect 2023 458 2027 462
rect 1239 402 1243 406
rect 1279 390 1283 394
rect 1303 390 1307 394
rect 1343 390 1347 394
rect 919 326 923 330
rect 975 326 979 330
rect 1031 326 1035 330
rect 1239 326 1243 330
rect 175 250 179 254
rect 215 250 219 254
rect 223 250 227 254
rect 255 250 259 254
rect 295 250 299 254
rect 311 250 315 254
rect 335 250 339 254
rect 391 250 395 254
rect 447 250 451 254
rect 463 250 467 254
rect 495 250 499 254
rect 527 250 531 254
rect 543 250 547 254
rect 591 250 595 254
rect 639 250 643 254
rect 647 250 651 254
rect 111 150 115 154
rect 135 150 139 154
rect 151 150 155 154
rect 191 150 195 154
rect 223 150 227 154
rect 231 150 235 154
rect 271 150 275 154
rect 311 150 315 154
rect 351 150 355 154
rect 391 150 395 154
rect 431 150 435 154
rect 463 150 467 154
rect 471 150 475 154
rect 511 150 515 154
rect 527 150 531 154
rect 551 150 555 154
rect 591 150 595 154
rect 687 250 691 254
rect 695 250 699 254
rect 735 250 739 254
rect 783 250 787 254
rect 1359 390 1363 394
rect 1383 390 1387 394
rect 1399 390 1403 394
rect 1439 390 1443 394
rect 1447 390 1451 394
rect 1487 390 1491 394
rect 1535 390 1539 394
rect 1543 390 1547 394
rect 1607 390 1611 394
rect 1631 390 1635 394
rect 1679 390 1683 394
rect 1735 390 1739 394
rect 1759 390 1763 394
rect 1831 390 1835 394
rect 1839 390 1843 394
rect 2167 526 2171 530
rect 2191 526 2195 530
rect 2239 526 2243 530
rect 2287 526 2291 530
rect 2311 526 2315 530
rect 2359 526 2363 530
rect 2407 526 2411 530
rect 2071 458 2075 462
rect 2103 458 2107 462
rect 2135 458 2139 462
rect 2191 458 2195 462
rect 2199 458 2203 462
rect 2255 458 2259 462
rect 2287 458 2291 462
rect 2319 458 2323 462
rect 2359 458 2363 462
rect 1919 390 1923 394
rect 1999 390 2003 394
rect 2071 390 2075 394
rect 2079 390 2083 394
rect 1279 314 1283 318
rect 1359 314 1363 318
rect 1399 314 1403 318
rect 1439 314 1443 318
rect 1487 314 1491 318
rect 1511 314 1515 318
rect 1543 314 1547 318
rect 1551 314 1555 318
rect 1591 314 1595 318
rect 1607 314 1611 318
rect 2135 390 2139 394
rect 2159 390 2163 394
rect 2199 390 2203 394
rect 2247 390 2251 394
rect 2255 390 2259 394
rect 2407 458 2411 462
rect 2319 390 2323 394
rect 2335 390 2339 394
rect 1631 314 1635 318
rect 1671 314 1675 318
rect 1679 314 1683 318
rect 1711 314 1715 318
rect 1751 314 1755 318
rect 1759 314 1763 318
rect 1791 314 1795 318
rect 1839 314 1843 318
rect 1903 314 1907 318
rect 1919 314 1923 318
rect 1967 314 1971 318
rect 1999 314 2003 318
rect 2039 314 2043 318
rect 2079 314 2083 318
rect 2119 314 2123 318
rect 2159 314 2163 318
rect 2199 314 2203 318
rect 2359 390 2363 394
rect 2407 390 2411 394
rect 2247 314 2251 318
rect 2279 314 2283 318
rect 2335 314 2339 318
rect 2359 314 2363 318
rect 2407 314 2411 318
rect 831 250 835 254
rect 839 250 843 254
rect 879 250 883 254
rect 927 250 931 254
rect 975 250 979 254
rect 1023 250 1027 254
rect 1239 250 1243 254
rect 1279 242 1283 246
rect 1367 242 1371 246
rect 1407 242 1411 246
rect 1455 242 1459 246
rect 1511 242 1515 246
rect 1551 242 1555 246
rect 1567 242 1571 246
rect 1591 242 1595 246
rect 1631 242 1635 246
rect 1671 242 1675 246
rect 631 150 635 154
rect 647 150 651 154
rect 671 150 675 154
rect 695 150 699 154
rect 711 150 715 154
rect 735 150 739 154
rect 751 150 755 154
rect 783 150 787 154
rect 791 150 795 154
rect 831 150 835 154
rect 871 150 875 154
rect 879 150 883 154
rect 911 150 915 154
rect 927 150 931 154
rect 951 150 955 154
rect 975 150 979 154
rect 991 150 995 154
rect 1023 150 1027 154
rect 1031 150 1035 154
rect 651 112 655 116
rect 1279 166 1283 170
rect 1303 166 1307 170
rect 1343 166 1347 170
rect 1367 166 1371 170
rect 1383 166 1387 170
rect 1407 166 1411 170
rect 1423 166 1427 170
rect 1455 166 1459 170
rect 1463 166 1467 170
rect 1511 166 1515 170
rect 1519 166 1523 170
rect 1567 166 1571 170
rect 1583 166 1587 170
rect 1631 166 1635 170
rect 1647 166 1651 170
rect 1071 150 1075 154
rect 1111 150 1115 154
rect 1151 150 1155 154
rect 1191 150 1195 154
rect 1239 150 1243 154
rect 1039 112 1043 116
rect 1703 242 1707 246
rect 1711 242 1715 246
rect 1751 242 1755 246
rect 1775 242 1779 246
rect 1791 242 1795 246
rect 1839 242 1843 246
rect 1855 242 1859 246
rect 1903 242 1907 246
rect 1943 242 1947 246
rect 1967 242 1971 246
rect 2031 242 2035 246
rect 2039 242 2043 246
rect 2119 242 2123 246
rect 2199 242 2203 246
rect 2207 242 2211 246
rect 2279 242 2283 246
rect 2295 242 2299 246
rect 1703 166 1707 170
rect 1711 166 1715 170
rect 1775 166 1779 170
rect 1831 166 1835 170
rect 1855 166 1859 170
rect 1887 166 1891 170
rect 1935 166 1939 170
rect 1943 166 1947 170
rect 1975 166 1979 170
rect 2015 166 2019 170
rect 2031 166 2035 170
rect 2055 166 2059 170
rect 2095 166 2099 170
rect 2119 166 2123 170
rect 2143 166 2147 170
rect 2191 166 2195 170
rect 2207 166 2211 170
rect 2359 242 2363 246
rect 2407 242 2411 246
rect 2239 166 2243 170
rect 2279 166 2283 170
rect 2295 166 2299 170
rect 2319 166 2323 170
rect 2359 166 2363 170
rect 2407 166 2411 170
rect 1279 98 1283 102
rect 1303 98 1307 102
rect 1343 98 1347 102
rect 1383 98 1387 102
rect 1423 98 1427 102
rect 1463 98 1467 102
rect 1519 98 1523 102
rect 1583 98 1587 102
rect 1647 98 1651 102
rect 1711 98 1715 102
rect 1775 98 1779 102
rect 1831 98 1835 102
rect 1887 98 1891 102
rect 1935 98 1939 102
rect 1975 98 1979 102
rect 2015 98 2019 102
rect 2055 98 2059 102
rect 2095 98 2099 102
rect 2143 98 2147 102
rect 2191 98 2195 102
rect 2239 98 2243 102
rect 2279 98 2283 102
rect 2319 98 2323 102
rect 2359 98 2363 102
rect 2407 98 2411 102
rect 111 82 115 86
rect 151 82 155 86
rect 191 82 195 86
rect 231 82 235 86
rect 271 82 275 86
rect 311 82 315 86
rect 351 82 355 86
rect 391 82 395 86
rect 431 82 435 86
rect 471 82 475 86
rect 511 82 515 86
rect 551 82 555 86
rect 591 82 595 86
rect 631 82 635 86
rect 671 82 675 86
rect 711 82 715 86
rect 751 82 755 86
rect 791 82 795 86
rect 831 82 835 86
rect 871 82 875 86
rect 911 82 915 86
rect 951 82 955 86
rect 991 82 995 86
rect 1031 82 1035 86
rect 1071 82 1075 86
rect 1111 82 1115 86
rect 1151 82 1155 86
rect 1191 82 1195 86
rect 1239 82 1243 86
<< m4 >>
rect 96 2489 97 2495
rect 103 2494 1263 2495
rect 103 2490 111 2494
rect 115 2490 231 2494
rect 235 2490 271 2494
rect 275 2490 311 2494
rect 315 2490 351 2494
rect 355 2490 399 2494
rect 403 2490 455 2494
rect 459 2490 511 2494
rect 515 2490 575 2494
rect 579 2490 639 2494
rect 643 2490 703 2494
rect 707 2490 767 2494
rect 771 2490 823 2494
rect 827 2490 879 2494
rect 883 2490 927 2494
rect 931 2490 975 2494
rect 979 2490 1023 2494
rect 1027 2490 1071 2494
rect 1075 2490 1111 2494
rect 1115 2490 1151 2494
rect 1155 2490 1191 2494
rect 1195 2490 1239 2494
rect 1243 2490 1263 2494
rect 103 2489 1263 2490
rect 1269 2491 1270 2495
rect 1269 2490 2454 2491
rect 1269 2489 1279 2490
rect 1262 2486 1279 2489
rect 1283 2486 1303 2490
rect 1307 2486 1343 2490
rect 1347 2486 1383 2490
rect 1387 2486 1439 2490
rect 1443 2486 1511 2490
rect 1515 2486 1583 2490
rect 1587 2486 1663 2490
rect 1667 2486 1735 2490
rect 1739 2486 1807 2490
rect 1811 2486 1887 2490
rect 1891 2486 1967 2490
rect 1971 2486 2063 2490
rect 2067 2486 2167 2490
rect 2171 2486 2271 2490
rect 2275 2486 2359 2490
rect 2363 2486 2407 2490
rect 2411 2486 2454 2490
rect 1262 2485 2454 2486
rect 1250 2422 2442 2423
rect 1250 2419 1279 2422
rect 84 2413 85 2419
rect 91 2418 1251 2419
rect 91 2414 111 2418
rect 115 2414 199 2418
rect 203 2414 231 2418
rect 235 2414 263 2418
rect 267 2414 271 2418
rect 275 2414 311 2418
rect 315 2414 327 2418
rect 331 2414 351 2418
rect 355 2414 399 2418
rect 403 2414 455 2418
rect 459 2414 471 2418
rect 475 2414 511 2418
rect 515 2414 543 2418
rect 547 2414 575 2418
rect 579 2414 615 2418
rect 619 2414 639 2418
rect 643 2414 687 2418
rect 691 2414 703 2418
rect 707 2414 751 2418
rect 755 2414 767 2418
rect 771 2414 823 2418
rect 827 2414 879 2418
rect 883 2414 895 2418
rect 899 2414 927 2418
rect 931 2414 967 2418
rect 971 2414 975 2418
rect 979 2414 1023 2418
rect 1027 2414 1071 2418
rect 1075 2414 1111 2418
rect 1115 2414 1151 2418
rect 1155 2414 1191 2418
rect 1195 2414 1239 2418
rect 1243 2414 1251 2418
rect 91 2413 1251 2414
rect 1257 2418 1279 2419
rect 1283 2418 1303 2422
rect 1307 2418 1343 2422
rect 1347 2418 1375 2422
rect 1379 2418 1383 2422
rect 1387 2418 1415 2422
rect 1419 2418 1439 2422
rect 1443 2418 1455 2422
rect 1459 2418 1503 2422
rect 1507 2418 1511 2422
rect 1515 2418 1559 2422
rect 1563 2418 1583 2422
rect 1587 2418 1615 2422
rect 1619 2418 1663 2422
rect 1667 2418 1679 2422
rect 1683 2418 1735 2422
rect 1739 2418 1799 2422
rect 1803 2418 1807 2422
rect 1811 2418 1871 2422
rect 1875 2418 1887 2422
rect 1891 2418 1951 2422
rect 1955 2418 1967 2422
rect 1971 2418 2047 2422
rect 2051 2418 2063 2422
rect 2067 2418 2151 2422
rect 2155 2418 2167 2422
rect 2171 2418 2263 2422
rect 2267 2418 2271 2422
rect 2275 2418 2359 2422
rect 2363 2418 2407 2422
rect 2411 2418 2442 2422
rect 1257 2417 2442 2418
rect 1257 2413 1258 2417
rect 1262 2350 2454 2351
rect 1262 2347 1279 2350
rect 96 2341 97 2347
rect 103 2346 1263 2347
rect 103 2342 111 2346
rect 115 2342 199 2346
rect 203 2342 263 2346
rect 267 2342 271 2346
rect 275 2342 327 2346
rect 331 2342 399 2346
rect 403 2342 471 2346
rect 475 2342 543 2346
rect 547 2342 551 2346
rect 555 2342 615 2346
rect 619 2342 631 2346
rect 635 2342 687 2346
rect 691 2342 711 2346
rect 715 2342 751 2346
rect 755 2342 783 2346
rect 787 2342 823 2346
rect 827 2342 855 2346
rect 859 2342 895 2346
rect 899 2342 919 2346
rect 923 2342 967 2346
rect 971 2342 991 2346
rect 995 2342 1063 2346
rect 1067 2342 1239 2346
rect 1243 2342 1263 2346
rect 103 2341 1263 2342
rect 1269 2346 1279 2347
rect 1283 2346 1327 2350
rect 1331 2346 1375 2350
rect 1379 2346 1383 2350
rect 1387 2346 1415 2350
rect 1419 2346 1439 2350
rect 1443 2346 1455 2350
rect 1459 2346 1503 2350
rect 1507 2346 1559 2350
rect 1563 2346 1575 2350
rect 1579 2346 1615 2350
rect 1619 2346 1647 2350
rect 1651 2346 1679 2350
rect 1683 2346 1719 2350
rect 1723 2346 1735 2350
rect 1739 2346 1799 2350
rect 1803 2346 1871 2350
rect 1875 2346 1879 2350
rect 1883 2346 1951 2350
rect 1955 2346 1967 2350
rect 1971 2346 2047 2350
rect 2051 2346 2063 2350
rect 2067 2346 2151 2350
rect 2155 2346 2167 2350
rect 2171 2346 2263 2350
rect 2267 2346 2271 2350
rect 2275 2346 2359 2350
rect 2363 2346 2407 2350
rect 2411 2346 2454 2350
rect 1269 2345 2454 2346
rect 1269 2341 1270 2345
rect 1250 2277 1251 2283
rect 1257 2282 2435 2283
rect 1257 2278 1279 2282
rect 1283 2278 1327 2282
rect 1331 2278 1335 2282
rect 1339 2278 1383 2282
rect 1387 2278 1407 2282
rect 1411 2278 1439 2282
rect 1443 2278 1487 2282
rect 1491 2278 1503 2282
rect 1507 2278 1559 2282
rect 1563 2278 1575 2282
rect 1579 2278 1631 2282
rect 1635 2278 1647 2282
rect 1651 2278 1703 2282
rect 1707 2278 1719 2282
rect 1723 2278 1775 2282
rect 1779 2278 1799 2282
rect 1803 2278 1839 2282
rect 1843 2278 1879 2282
rect 1883 2278 1911 2282
rect 1915 2278 1967 2282
rect 1971 2278 1991 2282
rect 1995 2278 2063 2282
rect 2067 2278 2079 2282
rect 2083 2278 2167 2282
rect 2171 2278 2175 2282
rect 2179 2278 2271 2282
rect 2275 2278 2279 2282
rect 2283 2278 2359 2282
rect 2363 2278 2407 2282
rect 2411 2278 2435 2282
rect 1257 2277 2435 2278
rect 2441 2277 2442 2283
rect 84 2265 85 2271
rect 91 2270 1251 2271
rect 91 2266 111 2270
rect 115 2266 143 2270
rect 147 2266 183 2270
rect 187 2266 223 2270
rect 227 2266 271 2270
rect 275 2266 279 2270
rect 283 2266 327 2270
rect 331 2266 335 2270
rect 339 2266 399 2270
rect 403 2266 407 2270
rect 411 2266 471 2270
rect 475 2266 479 2270
rect 483 2266 551 2270
rect 555 2266 559 2270
rect 563 2266 631 2270
rect 635 2266 647 2270
rect 651 2266 711 2270
rect 715 2266 727 2270
rect 731 2266 783 2270
rect 787 2266 807 2270
rect 811 2266 855 2270
rect 859 2266 887 2270
rect 891 2266 919 2270
rect 923 2266 967 2270
rect 971 2266 991 2270
rect 995 2266 1047 2270
rect 1051 2266 1063 2270
rect 1067 2266 1127 2270
rect 1131 2266 1239 2270
rect 1243 2266 1251 2270
rect 91 2265 1251 2266
rect 1257 2265 1258 2271
rect 1262 2206 2454 2207
rect 1262 2203 1279 2206
rect 96 2197 97 2203
rect 103 2202 1263 2203
rect 103 2198 111 2202
rect 115 2198 135 2202
rect 139 2198 143 2202
rect 147 2198 183 2202
rect 187 2198 207 2202
rect 211 2198 223 2202
rect 227 2198 279 2202
rect 283 2198 335 2202
rect 339 2198 359 2202
rect 363 2198 407 2202
rect 411 2198 439 2202
rect 443 2198 479 2202
rect 483 2198 519 2202
rect 523 2198 559 2202
rect 563 2198 599 2202
rect 603 2198 647 2202
rect 651 2198 679 2202
rect 683 2198 727 2202
rect 731 2198 759 2202
rect 763 2198 807 2202
rect 811 2198 831 2202
rect 835 2198 887 2202
rect 891 2198 903 2202
rect 907 2198 967 2202
rect 971 2198 975 2202
rect 979 2198 1047 2202
rect 1051 2198 1119 2202
rect 1123 2198 1127 2202
rect 1131 2198 1239 2202
rect 1243 2198 1263 2202
rect 103 2197 1263 2198
rect 1269 2202 1279 2203
rect 1283 2202 1335 2206
rect 1339 2202 1375 2206
rect 1379 2202 1407 2206
rect 1411 2202 1439 2206
rect 1443 2202 1487 2206
rect 1491 2202 1511 2206
rect 1515 2202 1559 2206
rect 1563 2202 1591 2206
rect 1595 2202 1631 2206
rect 1635 2202 1671 2206
rect 1675 2202 1703 2206
rect 1707 2202 1751 2206
rect 1755 2202 1775 2206
rect 1779 2202 1831 2206
rect 1835 2202 1839 2206
rect 1843 2202 1903 2206
rect 1907 2202 1911 2206
rect 1915 2202 1967 2206
rect 1971 2202 1991 2206
rect 1995 2202 2031 2206
rect 2035 2202 2079 2206
rect 2083 2202 2095 2206
rect 2099 2202 2167 2206
rect 2171 2202 2175 2206
rect 2179 2202 2239 2206
rect 2243 2202 2279 2206
rect 2283 2202 2311 2206
rect 2315 2202 2359 2206
rect 2363 2202 2407 2206
rect 2411 2202 2454 2206
rect 1269 2201 2454 2202
rect 1269 2197 1270 2201
rect 1250 2133 1251 2139
rect 1257 2138 2435 2139
rect 1257 2134 1279 2138
rect 1283 2134 1375 2138
rect 1379 2134 1399 2138
rect 1403 2134 1439 2138
rect 1443 2134 1495 2138
rect 1499 2134 1511 2138
rect 1515 2134 1567 2138
rect 1571 2134 1591 2138
rect 1595 2134 1647 2138
rect 1651 2134 1671 2138
rect 1675 2134 1735 2138
rect 1739 2134 1751 2138
rect 1755 2134 1823 2138
rect 1827 2134 1831 2138
rect 1835 2134 1903 2138
rect 1907 2134 1911 2138
rect 1915 2134 1967 2138
rect 1971 2134 1999 2138
rect 2003 2134 2031 2138
rect 2035 2134 2087 2138
rect 2091 2134 2095 2138
rect 2099 2134 2167 2138
rect 2171 2134 2175 2138
rect 2179 2134 2239 2138
rect 2243 2134 2271 2138
rect 2275 2134 2311 2138
rect 2315 2134 2359 2138
rect 2363 2134 2407 2138
rect 2411 2134 2435 2138
rect 1257 2133 2435 2134
rect 2441 2133 2442 2139
rect 84 2121 85 2127
rect 91 2126 1251 2127
rect 91 2122 111 2126
rect 115 2122 135 2126
rect 139 2122 191 2126
rect 195 2122 207 2126
rect 211 2122 271 2126
rect 275 2122 279 2126
rect 283 2122 343 2126
rect 347 2122 359 2126
rect 363 2122 415 2126
rect 419 2122 439 2126
rect 443 2122 479 2126
rect 483 2122 519 2126
rect 523 2122 543 2126
rect 547 2122 599 2126
rect 603 2122 607 2126
rect 611 2122 671 2126
rect 675 2122 679 2126
rect 683 2122 735 2126
rect 739 2122 759 2126
rect 763 2122 791 2126
rect 795 2122 831 2126
rect 835 2122 839 2126
rect 843 2122 887 2126
rect 891 2122 903 2126
rect 907 2122 935 2126
rect 939 2122 975 2126
rect 979 2122 991 2126
rect 995 2122 1047 2126
rect 1051 2122 1119 2126
rect 1123 2122 1239 2126
rect 1243 2122 1251 2126
rect 91 2121 1251 2122
rect 1257 2121 1258 2127
rect 1938 2116 1944 2117
rect 2250 2116 2256 2117
rect 1938 2112 1939 2116
rect 1943 2112 2251 2116
rect 2255 2112 2256 2116
rect 1938 2111 1944 2112
rect 2250 2111 2256 2112
rect 1262 2065 1263 2071
rect 1269 2070 2447 2071
rect 1269 2066 1279 2070
rect 1283 2066 1399 2070
rect 1403 2066 1439 2070
rect 1443 2066 1495 2070
rect 1499 2066 1567 2070
rect 1571 2066 1647 2070
rect 1651 2066 1735 2070
rect 1739 2066 1823 2070
rect 1827 2066 1911 2070
rect 1915 2066 1999 2070
rect 2003 2066 2039 2070
rect 2043 2066 2079 2070
rect 2083 2066 2087 2070
rect 2091 2066 2119 2070
rect 2123 2066 2159 2070
rect 2163 2066 2175 2070
rect 2179 2066 2199 2070
rect 2203 2066 2239 2070
rect 2243 2066 2271 2070
rect 2275 2066 2279 2070
rect 2283 2066 2319 2070
rect 2323 2066 2359 2070
rect 2363 2066 2407 2070
rect 2411 2066 2447 2070
rect 1269 2065 2447 2066
rect 2453 2065 2454 2071
rect 96 2049 97 2055
rect 103 2054 1263 2055
rect 103 2050 111 2054
rect 115 2050 135 2054
rect 139 2050 175 2054
rect 179 2050 191 2054
rect 195 2050 215 2054
rect 219 2050 271 2054
rect 275 2050 279 2054
rect 283 2050 343 2054
rect 347 2050 351 2054
rect 355 2050 415 2054
rect 419 2050 423 2054
rect 427 2050 479 2054
rect 483 2050 487 2054
rect 491 2050 543 2054
rect 547 2050 551 2054
rect 555 2050 607 2054
rect 611 2050 615 2054
rect 619 2050 671 2054
rect 675 2050 679 2054
rect 683 2050 735 2054
rect 739 2050 743 2054
rect 747 2050 791 2054
rect 795 2050 815 2054
rect 819 2050 839 2054
rect 843 2050 887 2054
rect 891 2050 935 2054
rect 939 2050 991 2054
rect 995 2050 1047 2054
rect 1051 2050 1239 2054
rect 1243 2050 1263 2054
rect 103 2049 1263 2050
rect 1269 2049 1270 2055
rect 1250 1997 1251 2003
rect 1257 2002 2435 2003
rect 1257 1998 1279 2002
rect 1283 1998 1399 2002
rect 1403 1998 1439 2002
rect 1443 1998 1479 2002
rect 1483 1998 1519 2002
rect 1523 1998 1559 2002
rect 1563 1998 1599 2002
rect 1603 1998 1639 2002
rect 1643 1998 1679 2002
rect 1683 1998 1719 2002
rect 1723 1998 1767 2002
rect 1771 1998 1823 2002
rect 1827 1998 1871 2002
rect 1875 1998 1919 2002
rect 1923 1998 1967 2002
rect 1971 1998 2015 2002
rect 2019 1998 2039 2002
rect 2043 1998 2055 2002
rect 2059 1998 2079 2002
rect 2083 1998 2095 2002
rect 2099 1998 2119 2002
rect 2123 1998 2143 2002
rect 2147 1998 2159 2002
rect 2163 1998 2191 2002
rect 2195 1998 2199 2002
rect 2203 1998 2239 2002
rect 2243 1998 2279 2002
rect 2283 1998 2319 2002
rect 2323 1998 2359 2002
rect 2363 1998 2407 2002
rect 2411 1998 2435 2002
rect 1257 1997 2435 1998
rect 2441 1997 2442 2003
rect 84 1981 85 1987
rect 91 1986 1251 1987
rect 91 1982 111 1986
rect 115 1982 135 1986
rect 139 1982 175 1986
rect 179 1982 215 1986
rect 219 1982 271 1986
rect 275 1982 279 1986
rect 283 1982 343 1986
rect 347 1982 351 1986
rect 355 1982 415 1986
rect 419 1982 423 1986
rect 427 1982 487 1986
rect 491 1982 495 1986
rect 499 1982 551 1986
rect 555 1982 575 1986
rect 579 1982 615 1986
rect 619 1982 647 1986
rect 651 1982 679 1986
rect 683 1982 719 1986
rect 723 1982 743 1986
rect 747 1982 791 1986
rect 795 1982 815 1986
rect 819 1982 863 1986
rect 867 1982 935 1986
rect 939 1982 1007 1986
rect 1011 1982 1239 1986
rect 1243 1982 1251 1986
rect 91 1981 1251 1982
rect 1257 1981 1258 1987
rect 1262 1925 1263 1931
rect 1269 1930 2447 1931
rect 1269 1926 1279 1930
rect 1283 1926 1343 1930
rect 1347 1926 1383 1930
rect 1387 1926 1399 1930
rect 1403 1926 1423 1930
rect 1427 1926 1439 1930
rect 1443 1926 1463 1930
rect 1467 1926 1479 1930
rect 1483 1926 1511 1930
rect 1515 1926 1519 1930
rect 1523 1926 1559 1930
rect 1563 1926 1567 1930
rect 1571 1926 1599 1930
rect 1603 1926 1631 1930
rect 1635 1926 1639 1930
rect 1643 1926 1679 1930
rect 1683 1926 1711 1930
rect 1715 1926 1719 1930
rect 1723 1926 1767 1930
rect 1771 1926 1807 1930
rect 1811 1926 1823 1930
rect 1827 1926 1871 1930
rect 1875 1926 1919 1930
rect 1923 1926 1967 1930
rect 1971 1926 2015 1930
rect 2019 1926 2031 1930
rect 2035 1926 2055 1930
rect 2059 1926 2095 1930
rect 2099 1926 2143 1930
rect 2147 1926 2151 1930
rect 2155 1926 2191 1930
rect 2195 1926 2239 1930
rect 2243 1926 2279 1930
rect 2283 1926 2319 1930
rect 2323 1926 2359 1930
rect 2363 1926 2407 1930
rect 2411 1926 2447 1930
rect 1269 1925 2447 1926
rect 2453 1925 2454 1931
rect 96 1909 97 1915
rect 103 1914 1263 1915
rect 103 1910 111 1914
rect 115 1910 135 1914
rect 139 1910 175 1914
rect 179 1910 215 1914
rect 219 1910 247 1914
rect 251 1910 271 1914
rect 275 1910 287 1914
rect 291 1910 327 1914
rect 331 1910 343 1914
rect 347 1910 367 1914
rect 371 1910 415 1914
rect 419 1910 471 1914
rect 475 1910 495 1914
rect 499 1910 535 1914
rect 539 1910 575 1914
rect 579 1910 599 1914
rect 603 1910 647 1914
rect 651 1910 663 1914
rect 667 1910 719 1914
rect 723 1910 727 1914
rect 731 1910 791 1914
rect 795 1910 855 1914
rect 859 1910 863 1914
rect 867 1910 919 1914
rect 923 1910 935 1914
rect 939 1910 983 1914
rect 987 1910 1007 1914
rect 1011 1910 1055 1914
rect 1059 1910 1127 1914
rect 1131 1910 1239 1914
rect 1243 1910 1263 1914
rect 103 1909 1263 1910
rect 1269 1909 1270 1915
rect 1250 1849 1251 1855
rect 1257 1854 2435 1855
rect 1257 1850 1279 1854
rect 1283 1850 1343 1854
rect 1347 1850 1359 1854
rect 1363 1850 1383 1854
rect 1387 1850 1399 1854
rect 1403 1850 1423 1854
rect 1427 1850 1447 1854
rect 1451 1850 1463 1854
rect 1467 1850 1503 1854
rect 1507 1850 1511 1854
rect 1515 1850 1559 1854
rect 1563 1850 1567 1854
rect 1571 1850 1615 1854
rect 1619 1850 1631 1854
rect 1635 1850 1671 1854
rect 1675 1850 1711 1854
rect 1715 1850 1727 1854
rect 1731 1850 1783 1854
rect 1787 1850 1807 1854
rect 1811 1850 1839 1854
rect 1843 1850 1895 1854
rect 1899 1850 1919 1854
rect 1923 1850 1951 1854
rect 1955 1850 2031 1854
rect 2035 1850 2151 1854
rect 2155 1850 2407 1854
rect 2411 1850 2435 1854
rect 1257 1849 2435 1850
rect 2441 1849 2442 1855
rect 84 1837 85 1843
rect 91 1842 1251 1843
rect 91 1838 111 1842
rect 115 1838 247 1842
rect 251 1838 287 1842
rect 291 1838 327 1842
rect 331 1838 367 1842
rect 371 1838 399 1842
rect 403 1838 415 1842
rect 419 1838 439 1842
rect 443 1838 471 1842
rect 475 1838 479 1842
rect 483 1838 519 1842
rect 523 1838 535 1842
rect 539 1838 567 1842
rect 571 1838 599 1842
rect 603 1838 623 1842
rect 627 1838 663 1842
rect 667 1838 687 1842
rect 691 1838 727 1842
rect 731 1838 759 1842
rect 763 1838 791 1842
rect 795 1838 831 1842
rect 835 1838 855 1842
rect 859 1838 903 1842
rect 907 1838 919 1842
rect 923 1838 975 1842
rect 979 1838 983 1842
rect 987 1838 1047 1842
rect 1051 1838 1055 1842
rect 1059 1838 1127 1842
rect 1131 1838 1191 1842
rect 1195 1838 1239 1842
rect 1243 1838 1251 1842
rect 91 1837 1251 1838
rect 1257 1837 1258 1843
rect 96 1769 97 1775
rect 103 1774 1263 1775
rect 103 1770 111 1774
rect 115 1770 399 1774
rect 403 1770 407 1774
rect 411 1770 439 1774
rect 443 1770 447 1774
rect 451 1770 479 1774
rect 483 1770 487 1774
rect 491 1770 519 1774
rect 523 1770 527 1774
rect 531 1770 567 1774
rect 571 1770 607 1774
rect 611 1770 623 1774
rect 627 1770 647 1774
rect 651 1770 687 1774
rect 691 1770 695 1774
rect 699 1770 751 1774
rect 755 1770 759 1774
rect 763 1770 807 1774
rect 811 1770 831 1774
rect 835 1770 871 1774
rect 875 1770 903 1774
rect 907 1770 935 1774
rect 939 1770 975 1774
rect 979 1770 999 1774
rect 1003 1770 1047 1774
rect 1051 1770 1071 1774
rect 1075 1770 1127 1774
rect 1131 1770 1143 1774
rect 1147 1770 1191 1774
rect 1195 1770 1239 1774
rect 1243 1770 1263 1774
rect 103 1769 1263 1770
rect 1269 1774 2454 1775
rect 1269 1770 1279 1774
rect 1283 1770 1303 1774
rect 1307 1770 1343 1774
rect 1347 1770 1359 1774
rect 1363 1770 1391 1774
rect 1395 1770 1399 1774
rect 1403 1770 1447 1774
rect 1451 1770 1455 1774
rect 1459 1770 1503 1774
rect 1507 1770 1519 1774
rect 1523 1770 1559 1774
rect 1563 1770 1583 1774
rect 1587 1770 1615 1774
rect 1619 1770 1647 1774
rect 1651 1770 1671 1774
rect 1675 1770 1703 1774
rect 1707 1770 1727 1774
rect 1731 1770 1759 1774
rect 1763 1770 1783 1774
rect 1787 1770 1807 1774
rect 1811 1770 1839 1774
rect 1843 1770 1863 1774
rect 1867 1770 1895 1774
rect 1899 1770 1919 1774
rect 1923 1770 1951 1774
rect 1955 1770 1975 1774
rect 1979 1770 2407 1774
rect 2411 1770 2454 1774
rect 1269 1769 2454 1770
rect 84 1697 85 1703
rect 91 1702 1251 1703
rect 91 1698 111 1702
rect 115 1698 279 1702
rect 283 1698 319 1702
rect 323 1698 359 1702
rect 363 1698 399 1702
rect 403 1698 407 1702
rect 411 1698 447 1702
rect 451 1698 487 1702
rect 491 1698 495 1702
rect 499 1698 527 1702
rect 531 1698 543 1702
rect 547 1698 567 1702
rect 571 1698 591 1702
rect 595 1698 607 1702
rect 611 1698 639 1702
rect 643 1698 647 1702
rect 651 1698 687 1702
rect 691 1698 695 1702
rect 699 1698 735 1702
rect 739 1698 751 1702
rect 755 1698 783 1702
rect 787 1698 807 1702
rect 811 1698 839 1702
rect 843 1698 871 1702
rect 875 1698 895 1702
rect 899 1698 935 1702
rect 939 1698 999 1702
rect 1003 1698 1071 1702
rect 1075 1698 1143 1702
rect 1147 1698 1191 1702
rect 1195 1698 1239 1702
rect 1243 1698 1251 1702
rect 91 1697 1251 1698
rect 1257 1702 2442 1703
rect 1257 1698 1279 1702
rect 1283 1698 1303 1702
rect 1307 1698 1343 1702
rect 1347 1698 1383 1702
rect 1387 1698 1391 1702
rect 1395 1698 1423 1702
rect 1427 1698 1455 1702
rect 1459 1698 1463 1702
rect 1467 1698 1503 1702
rect 1507 1698 1519 1702
rect 1523 1698 1559 1702
rect 1563 1698 1583 1702
rect 1587 1698 1623 1702
rect 1627 1698 1647 1702
rect 1651 1698 1687 1702
rect 1691 1698 1703 1702
rect 1707 1698 1751 1702
rect 1755 1698 1759 1702
rect 1763 1698 1807 1702
rect 1811 1698 1863 1702
rect 1867 1698 1919 1702
rect 1923 1698 1975 1702
rect 1979 1698 2031 1702
rect 2035 1698 2087 1702
rect 2091 1698 2407 1702
rect 2411 1698 2442 1702
rect 1257 1697 2442 1698
rect 96 1625 97 1631
rect 103 1630 1263 1631
rect 103 1626 111 1630
rect 115 1626 135 1630
rect 139 1626 175 1630
rect 179 1626 215 1630
rect 219 1626 255 1630
rect 259 1626 279 1630
rect 283 1626 311 1630
rect 315 1626 319 1630
rect 323 1626 359 1630
rect 363 1626 391 1630
rect 395 1626 399 1630
rect 403 1626 447 1630
rect 451 1626 471 1630
rect 475 1626 495 1630
rect 499 1626 543 1630
rect 547 1626 559 1630
rect 563 1626 591 1630
rect 595 1626 639 1630
rect 643 1626 687 1630
rect 691 1626 719 1630
rect 723 1626 735 1630
rect 739 1626 783 1630
rect 787 1626 791 1630
rect 795 1626 839 1630
rect 843 1626 855 1630
rect 859 1626 895 1630
rect 899 1626 919 1630
rect 923 1626 983 1630
rect 987 1626 1047 1630
rect 1051 1626 1239 1630
rect 1243 1626 1263 1630
rect 103 1625 1263 1626
rect 1269 1630 2454 1631
rect 1269 1626 1279 1630
rect 1283 1626 1303 1630
rect 1307 1626 1343 1630
rect 1347 1626 1383 1630
rect 1387 1626 1423 1630
rect 1427 1626 1463 1630
rect 1467 1626 1503 1630
rect 1507 1626 1559 1630
rect 1563 1626 1623 1630
rect 1627 1626 1631 1630
rect 1635 1626 1687 1630
rect 1691 1626 1703 1630
rect 1707 1626 1751 1630
rect 1755 1626 1783 1630
rect 1787 1626 1807 1630
rect 1811 1626 1855 1630
rect 1859 1626 1863 1630
rect 1867 1626 1919 1630
rect 1923 1626 1927 1630
rect 1931 1626 1975 1630
rect 1979 1626 1999 1630
rect 2003 1626 2031 1630
rect 2035 1626 2063 1630
rect 2067 1626 2087 1630
rect 2091 1626 2127 1630
rect 2131 1626 2191 1630
rect 2195 1626 2255 1630
rect 2259 1626 2319 1630
rect 2323 1626 2359 1630
rect 2363 1626 2407 1630
rect 2411 1626 2454 1630
rect 1269 1625 2454 1626
rect 1250 1562 2442 1563
rect 1250 1559 1279 1562
rect 84 1553 85 1559
rect 91 1558 1251 1559
rect 91 1554 111 1558
rect 115 1554 135 1558
rect 139 1554 151 1558
rect 155 1554 175 1558
rect 179 1554 199 1558
rect 203 1554 215 1558
rect 219 1554 255 1558
rect 259 1554 263 1558
rect 267 1554 311 1558
rect 315 1554 343 1558
rect 347 1554 391 1558
rect 395 1554 439 1558
rect 443 1554 471 1558
rect 475 1554 535 1558
rect 539 1554 559 1558
rect 563 1554 639 1558
rect 643 1554 719 1558
rect 723 1554 735 1558
rect 739 1554 791 1558
rect 795 1554 823 1558
rect 827 1554 855 1558
rect 859 1554 903 1558
rect 907 1554 919 1558
rect 923 1554 975 1558
rect 979 1554 983 1558
rect 987 1554 1047 1558
rect 1051 1554 1119 1558
rect 1123 1554 1191 1558
rect 1195 1554 1239 1558
rect 1243 1554 1251 1558
rect 91 1553 1251 1554
rect 1257 1558 1279 1559
rect 1283 1558 1303 1562
rect 1307 1558 1343 1562
rect 1347 1558 1383 1562
rect 1387 1558 1423 1562
rect 1427 1558 1463 1562
rect 1467 1558 1471 1562
rect 1475 1558 1503 1562
rect 1507 1558 1559 1562
rect 1563 1558 1623 1562
rect 1627 1558 1631 1562
rect 1635 1558 1703 1562
rect 1707 1558 1759 1562
rect 1763 1558 1783 1562
rect 1787 1558 1855 1562
rect 1859 1558 1871 1562
rect 1875 1558 1927 1562
rect 1931 1558 1967 1562
rect 1971 1558 1999 1562
rect 2003 1558 2055 1562
rect 2059 1558 2063 1562
rect 2067 1558 2127 1562
rect 2131 1558 2191 1562
rect 2195 1558 2255 1562
rect 2259 1558 2319 1562
rect 2323 1558 2359 1562
rect 2363 1558 2407 1562
rect 2411 1558 2442 1562
rect 1257 1557 2442 1558
rect 1257 1553 1258 1557
rect 96 1481 97 1487
rect 103 1486 1263 1487
rect 103 1482 111 1486
rect 115 1482 151 1486
rect 155 1482 199 1486
rect 203 1482 263 1486
rect 267 1482 319 1486
rect 323 1482 343 1486
rect 347 1482 359 1486
rect 363 1482 399 1486
rect 403 1482 439 1486
rect 443 1482 447 1486
rect 451 1482 503 1486
rect 507 1482 535 1486
rect 539 1482 559 1486
rect 563 1482 615 1486
rect 619 1482 639 1486
rect 643 1482 671 1486
rect 675 1482 735 1486
rect 739 1482 799 1486
rect 803 1482 823 1486
rect 827 1482 855 1486
rect 859 1482 903 1486
rect 907 1482 911 1486
rect 915 1482 967 1486
rect 971 1482 975 1486
rect 979 1482 1023 1486
rect 1027 1482 1047 1486
rect 1051 1482 1087 1486
rect 1091 1482 1119 1486
rect 1123 1482 1151 1486
rect 1155 1482 1191 1486
rect 1195 1482 1239 1486
rect 1243 1482 1263 1486
rect 103 1481 1263 1482
rect 1269 1481 1270 1487
rect 1262 1469 1263 1475
rect 1269 1474 2447 1475
rect 1269 1470 1279 1474
rect 1283 1470 1303 1474
rect 1307 1470 1375 1474
rect 1379 1470 1471 1474
rect 1475 1470 1479 1474
rect 1483 1470 1583 1474
rect 1587 1470 1623 1474
rect 1627 1470 1687 1474
rect 1691 1470 1759 1474
rect 1763 1470 1783 1474
rect 1787 1470 1871 1474
rect 1875 1470 1951 1474
rect 1955 1470 1967 1474
rect 1971 1470 2031 1474
rect 2035 1470 2055 1474
rect 2059 1470 2103 1474
rect 2107 1470 2127 1474
rect 2131 1470 2167 1474
rect 2171 1470 2191 1474
rect 2195 1470 2239 1474
rect 2243 1470 2255 1474
rect 2259 1470 2311 1474
rect 2315 1470 2319 1474
rect 2323 1470 2359 1474
rect 2363 1470 2407 1474
rect 2411 1470 2447 1474
rect 1269 1469 2447 1470
rect 2453 1469 2454 1475
rect 84 1409 85 1415
rect 91 1414 1251 1415
rect 91 1410 111 1414
rect 115 1410 263 1414
rect 267 1410 303 1414
rect 307 1410 319 1414
rect 323 1410 343 1414
rect 347 1410 359 1414
rect 363 1410 391 1414
rect 395 1410 399 1414
rect 403 1410 447 1414
rect 451 1410 503 1414
rect 507 1410 559 1414
rect 563 1410 615 1414
rect 619 1410 623 1414
rect 627 1410 671 1414
rect 675 1410 687 1414
rect 691 1410 735 1414
rect 739 1410 751 1414
rect 755 1410 799 1414
rect 803 1410 815 1414
rect 819 1410 855 1414
rect 859 1410 879 1414
rect 883 1410 911 1414
rect 915 1410 951 1414
rect 955 1410 967 1414
rect 971 1410 1023 1414
rect 1027 1410 1087 1414
rect 1091 1410 1151 1414
rect 1155 1410 1191 1414
rect 1195 1410 1239 1414
rect 1243 1410 1251 1414
rect 91 1409 1251 1410
rect 1257 1409 1258 1415
rect 1250 1407 1258 1409
rect 1250 1401 1251 1407
rect 1257 1406 2435 1407
rect 1257 1402 1279 1406
rect 1283 1402 1303 1406
rect 1307 1402 1343 1406
rect 1347 1402 1375 1406
rect 1379 1402 1399 1406
rect 1403 1402 1471 1406
rect 1475 1402 1479 1406
rect 1483 1402 1551 1406
rect 1555 1402 1583 1406
rect 1587 1402 1639 1406
rect 1643 1402 1687 1406
rect 1691 1402 1727 1406
rect 1731 1402 1783 1406
rect 1787 1402 1815 1406
rect 1819 1402 1871 1406
rect 1875 1402 1903 1406
rect 1907 1402 1951 1406
rect 1955 1402 1991 1406
rect 1995 1402 2031 1406
rect 2035 1402 2071 1406
rect 2075 1402 2103 1406
rect 2107 1402 2151 1406
rect 2155 1402 2167 1406
rect 2171 1402 2223 1406
rect 2227 1402 2239 1406
rect 2243 1402 2303 1406
rect 2307 1402 2311 1406
rect 2315 1402 2359 1406
rect 2363 1402 2407 1406
rect 2411 1402 2435 1406
rect 1257 1401 2435 1402
rect 2441 1401 2442 1407
rect 96 1337 97 1343
rect 103 1342 1263 1343
rect 103 1338 111 1342
rect 115 1338 135 1342
rect 139 1338 175 1342
rect 179 1338 215 1342
rect 219 1338 255 1342
rect 259 1338 263 1342
rect 267 1338 303 1342
rect 307 1338 327 1342
rect 331 1338 343 1342
rect 347 1338 391 1342
rect 395 1338 407 1342
rect 411 1338 447 1342
rect 451 1338 495 1342
rect 499 1338 503 1342
rect 507 1338 559 1342
rect 563 1338 583 1342
rect 587 1338 623 1342
rect 627 1338 671 1342
rect 675 1338 687 1342
rect 691 1338 751 1342
rect 755 1338 759 1342
rect 763 1338 815 1342
rect 819 1338 839 1342
rect 843 1338 879 1342
rect 883 1338 919 1342
rect 923 1338 951 1342
rect 955 1338 1007 1342
rect 1011 1338 1023 1342
rect 1027 1338 1095 1342
rect 1099 1338 1239 1342
rect 1243 1338 1263 1342
rect 103 1337 1263 1338
rect 1269 1337 1270 1343
rect 1262 1335 1270 1337
rect 1262 1329 1263 1335
rect 1269 1334 2447 1335
rect 1269 1330 1279 1334
rect 1283 1330 1303 1334
rect 1307 1330 1343 1334
rect 1347 1330 1399 1334
rect 1403 1330 1447 1334
rect 1451 1330 1471 1334
rect 1475 1330 1487 1334
rect 1491 1330 1527 1334
rect 1531 1330 1551 1334
rect 1555 1330 1567 1334
rect 1571 1330 1615 1334
rect 1619 1330 1639 1334
rect 1643 1330 1671 1334
rect 1675 1330 1719 1334
rect 1723 1330 1727 1334
rect 1731 1330 1775 1334
rect 1779 1330 1815 1334
rect 1819 1330 1831 1334
rect 1835 1330 1903 1334
rect 1907 1330 1983 1334
rect 1987 1330 1991 1334
rect 1995 1330 2071 1334
rect 2075 1330 2151 1334
rect 2155 1330 2167 1334
rect 2171 1330 2223 1334
rect 2227 1330 2271 1334
rect 2275 1330 2303 1334
rect 2307 1330 2359 1334
rect 2363 1330 2407 1334
rect 2411 1330 2447 1334
rect 1269 1329 2447 1330
rect 2453 1329 2454 1335
rect 84 1265 85 1271
rect 91 1270 1251 1271
rect 91 1266 111 1270
rect 115 1266 135 1270
rect 139 1266 175 1270
rect 179 1266 215 1270
rect 219 1266 247 1270
rect 251 1266 255 1270
rect 259 1266 327 1270
rect 331 1266 407 1270
rect 411 1266 415 1270
rect 419 1266 495 1270
rect 499 1266 503 1270
rect 507 1266 583 1270
rect 587 1266 591 1270
rect 595 1266 671 1270
rect 675 1266 743 1270
rect 747 1266 759 1270
rect 763 1266 815 1270
rect 819 1266 839 1270
rect 843 1266 879 1270
rect 883 1266 919 1270
rect 923 1266 943 1270
rect 947 1266 1007 1270
rect 1011 1266 1071 1270
rect 1075 1266 1095 1270
rect 1099 1266 1239 1270
rect 1243 1266 1251 1270
rect 91 1265 1251 1266
rect 1257 1265 1258 1271
rect 1250 1263 1258 1265
rect 1250 1257 1251 1263
rect 1257 1262 2435 1263
rect 1257 1258 1279 1262
rect 1283 1258 1447 1262
rect 1451 1258 1487 1262
rect 1491 1258 1511 1262
rect 1515 1258 1527 1262
rect 1531 1258 1551 1262
rect 1555 1258 1567 1262
rect 1571 1258 1591 1262
rect 1595 1258 1615 1262
rect 1619 1258 1631 1262
rect 1635 1258 1671 1262
rect 1675 1258 1711 1262
rect 1715 1258 1719 1262
rect 1723 1258 1751 1262
rect 1755 1258 1775 1262
rect 1779 1258 1791 1262
rect 1795 1258 1831 1262
rect 1835 1258 1839 1262
rect 1843 1258 1903 1262
rect 1907 1258 1967 1262
rect 1971 1258 1983 1262
rect 1987 1258 2039 1262
rect 2043 1258 2071 1262
rect 2075 1258 2119 1262
rect 2123 1258 2167 1262
rect 2171 1258 2207 1262
rect 2211 1258 2271 1262
rect 2275 1258 2295 1262
rect 2299 1258 2359 1262
rect 2363 1258 2407 1262
rect 2411 1258 2435 1262
rect 1257 1257 2435 1258
rect 2441 1257 2442 1263
rect 96 1189 97 1195
rect 103 1194 1263 1195
rect 103 1190 111 1194
rect 115 1190 135 1194
rect 139 1190 175 1194
rect 179 1190 231 1194
rect 235 1190 247 1194
rect 251 1190 303 1194
rect 307 1190 327 1194
rect 331 1190 383 1194
rect 387 1190 415 1194
rect 419 1190 471 1194
rect 475 1190 503 1194
rect 507 1190 559 1194
rect 563 1190 591 1194
rect 595 1190 639 1194
rect 643 1190 671 1194
rect 675 1190 719 1194
rect 723 1190 743 1194
rect 747 1190 799 1194
rect 803 1190 815 1194
rect 819 1190 871 1194
rect 875 1190 879 1194
rect 883 1190 935 1194
rect 939 1190 943 1194
rect 947 1190 991 1194
rect 995 1190 1007 1194
rect 1011 1190 1047 1194
rect 1051 1190 1071 1194
rect 1075 1190 1103 1194
rect 1107 1190 1151 1194
rect 1155 1190 1191 1194
rect 1195 1190 1239 1194
rect 1243 1190 1263 1194
rect 103 1189 1263 1190
rect 1269 1191 1270 1195
rect 1269 1190 2454 1191
rect 1269 1189 1279 1190
rect 1262 1186 1279 1189
rect 1283 1186 1511 1190
rect 1515 1186 1551 1190
rect 1555 1186 1559 1190
rect 1563 1186 1591 1190
rect 1595 1186 1599 1190
rect 1603 1186 1631 1190
rect 1635 1186 1639 1190
rect 1643 1186 1671 1190
rect 1675 1186 1679 1190
rect 1683 1186 1711 1190
rect 1715 1186 1719 1190
rect 1723 1186 1751 1190
rect 1755 1186 1759 1190
rect 1763 1186 1791 1190
rect 1795 1186 1799 1190
rect 1803 1186 1839 1190
rect 1843 1186 1855 1190
rect 1859 1186 1903 1190
rect 1907 1186 1927 1190
rect 1931 1186 1967 1190
rect 1971 1186 2023 1190
rect 2027 1186 2039 1190
rect 2043 1186 2119 1190
rect 2123 1186 2135 1190
rect 2139 1186 2207 1190
rect 2211 1186 2255 1190
rect 2259 1186 2295 1190
rect 2299 1186 2359 1190
rect 2363 1186 2407 1190
rect 2411 1186 2454 1190
rect 1262 1185 2454 1186
rect 84 1121 85 1127
rect 91 1126 1251 1127
rect 91 1122 111 1126
rect 115 1122 135 1126
rect 139 1122 175 1126
rect 179 1122 215 1126
rect 219 1122 231 1126
rect 235 1122 303 1126
rect 307 1122 383 1126
rect 387 1122 391 1126
rect 395 1122 471 1126
rect 475 1122 479 1126
rect 483 1122 559 1126
rect 563 1122 639 1126
rect 643 1122 711 1126
rect 715 1122 719 1126
rect 723 1122 775 1126
rect 779 1122 799 1126
rect 803 1122 839 1126
rect 843 1122 871 1126
rect 875 1122 903 1126
rect 907 1122 935 1126
rect 939 1122 959 1126
rect 963 1122 991 1126
rect 995 1122 1023 1126
rect 1027 1122 1047 1126
rect 1051 1122 1087 1126
rect 1091 1122 1103 1126
rect 1107 1122 1151 1126
rect 1155 1122 1191 1126
rect 1195 1122 1239 1126
rect 1243 1122 1251 1126
rect 91 1121 1251 1122
rect 1257 1121 1258 1127
rect 1250 1109 1251 1115
rect 1257 1114 2435 1115
rect 1257 1110 1279 1114
rect 1283 1110 1535 1114
rect 1539 1110 1559 1114
rect 1563 1110 1599 1114
rect 1603 1110 1639 1114
rect 1643 1110 1663 1114
rect 1667 1110 1679 1114
rect 1683 1110 1719 1114
rect 1723 1110 1727 1114
rect 1731 1110 1759 1114
rect 1763 1110 1791 1114
rect 1795 1110 1799 1114
rect 1803 1110 1855 1114
rect 1859 1110 1911 1114
rect 1915 1110 1927 1114
rect 1931 1110 1967 1114
rect 1971 1110 2023 1114
rect 2027 1110 2079 1114
rect 2083 1110 2135 1114
rect 2139 1110 2191 1114
rect 2195 1110 2255 1114
rect 2259 1110 2319 1114
rect 2323 1110 2359 1114
rect 2363 1110 2407 1114
rect 2411 1110 2435 1114
rect 1257 1109 2435 1110
rect 2441 1109 2442 1115
rect 96 1049 97 1055
rect 103 1054 1263 1055
rect 103 1050 111 1054
rect 115 1050 135 1054
rect 139 1050 199 1054
rect 203 1050 215 1054
rect 219 1050 239 1054
rect 243 1050 287 1054
rect 291 1050 303 1054
rect 307 1050 343 1054
rect 347 1050 391 1054
rect 395 1050 439 1054
rect 443 1050 479 1054
rect 483 1050 487 1054
rect 491 1050 535 1054
rect 539 1050 559 1054
rect 563 1050 583 1054
rect 587 1050 631 1054
rect 635 1050 639 1054
rect 643 1050 679 1054
rect 683 1050 711 1054
rect 715 1050 727 1054
rect 731 1050 775 1054
rect 779 1050 783 1054
rect 787 1050 839 1054
rect 843 1050 895 1054
rect 899 1050 903 1054
rect 907 1050 959 1054
rect 963 1050 1023 1054
rect 1027 1050 1087 1054
rect 1091 1050 1151 1054
rect 1155 1050 1191 1054
rect 1195 1050 1239 1054
rect 1243 1050 1263 1054
rect 103 1049 1263 1050
rect 1269 1049 1270 1055
rect 1262 1029 1263 1035
rect 1269 1034 2447 1035
rect 1269 1030 1279 1034
rect 1283 1030 1503 1034
rect 1507 1030 1535 1034
rect 1539 1030 1599 1034
rect 1603 1030 1623 1034
rect 1627 1030 1663 1034
rect 1667 1030 1727 1034
rect 1731 1030 1735 1034
rect 1739 1030 1791 1034
rect 1795 1030 1831 1034
rect 1835 1030 1855 1034
rect 1859 1030 1911 1034
rect 1915 1030 1919 1034
rect 1923 1030 1967 1034
rect 1971 1030 1999 1034
rect 2003 1030 2023 1034
rect 2027 1030 2071 1034
rect 2075 1030 2079 1034
rect 2083 1030 2135 1034
rect 2139 1030 2143 1034
rect 2147 1030 2191 1034
rect 2195 1030 2207 1034
rect 2211 1030 2255 1034
rect 2259 1030 2279 1034
rect 2283 1030 2319 1034
rect 2323 1030 2359 1034
rect 2363 1030 2407 1034
rect 2411 1030 2447 1034
rect 1269 1029 2447 1030
rect 2453 1029 2454 1035
rect 84 969 85 975
rect 91 974 1251 975
rect 91 970 111 974
rect 115 970 199 974
rect 203 970 239 974
rect 243 970 287 974
rect 291 970 295 974
rect 299 970 343 974
rect 347 970 391 974
rect 395 970 399 974
rect 403 970 439 974
rect 443 970 471 974
rect 475 970 487 974
rect 491 970 535 974
rect 539 970 551 974
rect 555 970 583 974
rect 587 970 631 974
rect 635 970 639 974
rect 643 970 679 974
rect 683 970 727 974
rect 731 970 783 974
rect 787 970 807 974
rect 811 970 839 974
rect 843 970 887 974
rect 891 970 895 974
rect 899 970 959 974
rect 963 970 1023 974
rect 1027 970 1087 974
rect 1091 970 1151 974
rect 1155 970 1191 974
rect 1195 970 1239 974
rect 1243 970 1251 974
rect 91 969 1251 970
rect 1257 969 1258 975
rect 1250 953 1251 959
rect 1257 958 2435 959
rect 1257 954 1279 958
rect 1283 954 1319 958
rect 1323 954 1359 958
rect 1363 954 1399 958
rect 1403 954 1463 958
rect 1467 954 1503 958
rect 1507 954 1543 958
rect 1547 954 1623 958
rect 1627 954 1639 958
rect 1643 954 1735 958
rect 1739 954 1831 958
rect 1835 954 1839 958
rect 1843 954 1919 958
rect 1923 954 1935 958
rect 1939 954 1999 958
rect 2003 954 2023 958
rect 2027 954 2071 958
rect 2075 954 2103 958
rect 2107 954 2143 958
rect 2147 954 2175 958
rect 2179 954 2207 958
rect 2211 954 2239 958
rect 2243 954 2279 958
rect 2283 954 2311 958
rect 2315 954 2359 958
rect 2363 954 2407 958
rect 2411 954 2435 958
rect 1257 953 2435 954
rect 2441 953 2442 959
rect 96 893 97 899
rect 103 898 1263 899
rect 103 894 111 898
rect 115 894 255 898
rect 259 894 295 898
rect 299 894 311 898
rect 315 894 343 898
rect 347 894 375 898
rect 379 894 399 898
rect 403 894 455 898
rect 459 894 471 898
rect 475 894 535 898
rect 539 894 551 898
rect 555 894 623 898
rect 627 894 639 898
rect 643 894 711 898
rect 715 894 727 898
rect 731 894 791 898
rect 795 894 807 898
rect 811 894 863 898
rect 867 894 887 898
rect 891 894 935 898
rect 939 894 959 898
rect 963 894 999 898
rect 1003 894 1023 898
rect 1027 894 1055 898
rect 1059 894 1087 898
rect 1091 894 1119 898
rect 1123 894 1151 898
rect 1155 894 1183 898
rect 1187 894 1191 898
rect 1195 894 1239 898
rect 1243 894 1263 898
rect 103 893 1263 894
rect 1269 893 1270 899
rect 1262 877 1263 883
rect 1269 882 2447 883
rect 1269 878 1279 882
rect 1283 878 1319 882
rect 1323 878 1335 882
rect 1339 878 1359 882
rect 1363 878 1375 882
rect 1379 878 1399 882
rect 1403 878 1415 882
rect 1419 878 1463 882
rect 1467 878 1471 882
rect 1475 878 1535 882
rect 1539 878 1543 882
rect 1547 878 1607 882
rect 1611 878 1639 882
rect 1643 878 1679 882
rect 1683 878 1735 882
rect 1739 878 1751 882
rect 1755 878 1823 882
rect 1827 878 1839 882
rect 1843 878 1895 882
rect 1899 878 1935 882
rect 1939 878 1959 882
rect 1963 878 2023 882
rect 2027 878 2087 882
rect 2091 878 2103 882
rect 2107 878 2143 882
rect 2147 878 2175 882
rect 2179 878 2199 882
rect 2203 878 2239 882
rect 2243 878 2255 882
rect 2259 878 2311 882
rect 2315 878 2319 882
rect 2323 878 2359 882
rect 2363 878 2407 882
rect 2411 878 2447 882
rect 1269 877 2447 878
rect 2453 877 2454 883
rect 84 825 85 831
rect 91 830 1251 831
rect 91 826 111 830
rect 115 826 191 830
rect 195 826 247 830
rect 251 826 255 830
rect 259 826 311 830
rect 315 826 375 830
rect 379 826 383 830
rect 387 826 455 830
rect 459 826 463 830
rect 467 826 535 830
rect 539 826 543 830
rect 547 826 615 830
rect 619 826 623 830
rect 627 826 687 830
rect 691 826 711 830
rect 715 826 751 830
rect 755 826 791 830
rect 795 826 815 830
rect 819 826 863 830
rect 867 826 871 830
rect 875 826 927 830
rect 931 826 935 830
rect 939 826 983 830
rect 987 826 999 830
rect 1003 826 1047 830
rect 1051 826 1055 830
rect 1059 826 1119 830
rect 1123 826 1183 830
rect 1187 826 1239 830
rect 1243 826 1251 830
rect 91 825 1251 826
rect 1257 825 1258 831
rect 1250 805 1251 811
rect 1257 810 2435 811
rect 1257 806 1279 810
rect 1283 806 1303 810
rect 1307 806 1335 810
rect 1339 806 1343 810
rect 1347 806 1375 810
rect 1379 806 1407 810
rect 1411 806 1415 810
rect 1419 806 1471 810
rect 1475 806 1479 810
rect 1483 806 1535 810
rect 1539 806 1551 810
rect 1555 806 1607 810
rect 1611 806 1623 810
rect 1627 806 1679 810
rect 1683 806 1695 810
rect 1699 806 1751 810
rect 1755 806 1759 810
rect 1763 806 1823 810
rect 1827 806 1887 810
rect 1891 806 1895 810
rect 1899 806 1951 810
rect 1955 806 1959 810
rect 1963 806 2023 810
rect 2027 806 2087 810
rect 2091 806 2103 810
rect 2107 806 2143 810
rect 2147 806 2191 810
rect 2195 806 2199 810
rect 2203 806 2255 810
rect 2259 806 2279 810
rect 2283 806 2319 810
rect 2323 806 2359 810
rect 2363 806 2407 810
rect 2411 806 2435 810
rect 1257 805 2435 806
rect 2441 805 2442 811
rect 96 757 97 763
rect 103 762 1263 763
rect 103 758 111 762
rect 115 758 135 762
rect 139 758 175 762
rect 179 758 191 762
rect 195 758 215 762
rect 219 758 247 762
rect 251 758 279 762
rect 283 758 311 762
rect 315 758 351 762
rect 355 758 383 762
rect 387 758 423 762
rect 427 758 463 762
rect 467 758 495 762
rect 499 758 543 762
rect 547 758 559 762
rect 563 758 615 762
rect 619 758 623 762
rect 627 758 687 762
rect 691 758 695 762
rect 699 758 751 762
rect 755 758 783 762
rect 787 758 815 762
rect 819 758 871 762
rect 875 758 879 762
rect 883 758 927 762
rect 931 758 983 762
rect 987 758 1047 762
rect 1051 758 1095 762
rect 1099 758 1191 762
rect 1195 758 1239 762
rect 1243 758 1263 762
rect 103 757 1263 758
rect 1269 757 1270 763
rect 1262 737 1263 743
rect 1269 742 2447 743
rect 1269 738 1279 742
rect 1283 738 1303 742
rect 1307 738 1343 742
rect 1347 738 1367 742
rect 1371 738 1407 742
rect 1411 738 1455 742
rect 1459 738 1479 742
rect 1483 738 1535 742
rect 1539 738 1551 742
rect 1555 738 1615 742
rect 1619 738 1623 742
rect 1627 738 1695 742
rect 1699 738 1759 742
rect 1763 738 1775 742
rect 1779 738 1823 742
rect 1827 738 1855 742
rect 1859 738 1887 742
rect 1891 738 1943 742
rect 1947 738 1951 742
rect 1955 738 2023 742
rect 2027 738 2031 742
rect 2035 738 2103 742
rect 2107 738 2119 742
rect 2123 738 2191 742
rect 2195 738 2207 742
rect 2211 738 2279 742
rect 2283 738 2295 742
rect 2299 738 2359 742
rect 2363 738 2407 742
rect 2411 738 2447 742
rect 1269 737 2447 738
rect 2453 737 2454 743
rect 84 681 85 687
rect 91 686 1251 687
rect 91 682 111 686
rect 115 682 135 686
rect 139 682 175 686
rect 179 682 215 686
rect 219 682 231 686
rect 235 682 279 686
rect 283 682 287 686
rect 291 682 343 686
rect 347 682 351 686
rect 355 682 399 686
rect 403 682 423 686
rect 427 682 455 686
rect 459 682 495 686
rect 499 682 503 686
rect 507 682 559 686
rect 563 682 623 686
rect 627 682 695 686
rect 699 682 767 686
rect 771 682 783 686
rect 787 682 839 686
rect 843 682 879 686
rect 883 682 903 686
rect 907 682 967 686
rect 971 682 983 686
rect 987 682 1023 686
rect 1027 682 1087 686
rect 1091 682 1095 686
rect 1099 682 1151 686
rect 1155 682 1191 686
rect 1195 682 1239 686
rect 1243 682 1251 686
rect 91 681 1251 682
rect 1257 681 1258 687
rect 1250 669 1251 675
rect 1257 674 2435 675
rect 1257 670 1279 674
rect 1283 670 1303 674
rect 1307 670 1367 674
rect 1371 670 1455 674
rect 1459 670 1535 674
rect 1539 670 1591 674
rect 1595 670 1615 674
rect 1619 670 1639 674
rect 1643 670 1687 674
rect 1691 670 1695 674
rect 1699 670 1743 674
rect 1747 670 1775 674
rect 1779 670 1799 674
rect 1803 670 1855 674
rect 1859 670 1871 674
rect 1875 670 1943 674
rect 1947 670 1951 674
rect 1955 670 2031 674
rect 2035 670 2047 674
rect 2051 670 2119 674
rect 2123 670 2151 674
rect 2155 670 2207 674
rect 2211 670 2263 674
rect 2267 670 2295 674
rect 2299 670 2359 674
rect 2363 670 2407 674
rect 2411 670 2435 674
rect 1257 669 2435 670
rect 2441 669 2442 675
rect 96 613 97 619
rect 103 618 1263 619
rect 103 614 111 618
rect 115 614 135 618
rect 139 614 175 618
rect 179 614 183 618
rect 187 614 231 618
rect 235 614 255 618
rect 259 614 287 618
rect 291 614 327 618
rect 331 614 343 618
rect 347 614 399 618
rect 403 614 455 618
rect 459 614 479 618
rect 483 614 503 618
rect 507 614 559 618
rect 563 614 623 618
rect 627 614 639 618
rect 643 614 695 618
rect 699 614 719 618
rect 723 614 767 618
rect 771 614 799 618
rect 803 614 839 618
rect 843 614 879 618
rect 883 614 903 618
rect 907 614 951 618
rect 955 614 967 618
rect 971 614 1015 618
rect 1019 614 1023 618
rect 1027 614 1079 618
rect 1083 614 1087 618
rect 1091 614 1143 618
rect 1147 614 1151 618
rect 1155 614 1191 618
rect 1195 614 1239 618
rect 1243 614 1263 618
rect 103 613 1263 614
rect 1269 613 1270 619
rect 1262 593 1263 599
rect 1269 598 2447 599
rect 1269 594 1279 598
rect 1283 594 1559 598
rect 1563 594 1591 598
rect 1595 594 1599 598
rect 1603 594 1639 598
rect 1643 594 1679 598
rect 1683 594 1687 598
rect 1691 594 1719 598
rect 1723 594 1743 598
rect 1747 594 1759 598
rect 1763 594 1799 598
rect 1803 594 1807 598
rect 1811 594 1855 598
rect 1859 594 1871 598
rect 1875 594 1911 598
rect 1915 594 1951 598
rect 1955 594 1967 598
rect 1971 594 2031 598
rect 2035 594 2047 598
rect 2051 594 2095 598
rect 2099 594 2151 598
rect 2155 594 2167 598
rect 2171 594 2239 598
rect 2243 594 2263 598
rect 2267 594 2311 598
rect 2315 594 2359 598
rect 2363 594 2407 598
rect 2411 594 2447 598
rect 1269 593 2447 594
rect 2453 593 2454 599
rect 84 541 85 547
rect 91 546 1251 547
rect 91 542 111 546
rect 115 542 135 546
rect 139 542 151 546
rect 155 542 183 546
rect 187 542 223 546
rect 227 542 255 546
rect 259 542 287 546
rect 291 542 327 546
rect 331 542 351 546
rect 355 542 399 546
rect 403 542 415 546
rect 419 542 479 546
rect 483 542 551 546
rect 555 542 559 546
rect 563 542 623 546
rect 627 542 639 546
rect 643 542 695 546
rect 699 542 719 546
rect 723 542 767 546
rect 771 542 799 546
rect 803 542 839 546
rect 843 542 879 546
rect 883 542 919 546
rect 923 542 951 546
rect 955 542 999 546
rect 1003 542 1015 546
rect 1019 542 1079 546
rect 1083 542 1143 546
rect 1147 542 1191 546
rect 1195 542 1239 546
rect 1243 542 1251 546
rect 91 541 1251 542
rect 1257 541 1258 547
rect 1250 525 1251 531
rect 1257 530 2435 531
rect 1257 526 1279 530
rect 1283 526 1407 530
rect 1411 526 1447 530
rect 1451 526 1487 530
rect 1491 526 1535 530
rect 1539 526 1559 530
rect 1563 526 1591 530
rect 1595 526 1599 530
rect 1603 526 1639 530
rect 1643 526 1647 530
rect 1651 526 1679 530
rect 1683 526 1711 530
rect 1715 526 1719 530
rect 1723 526 1759 530
rect 1763 526 1783 530
rect 1787 526 1807 530
rect 1811 526 1855 530
rect 1859 526 1863 530
rect 1867 526 1911 530
rect 1915 526 1943 530
rect 1947 526 1967 530
rect 1971 526 2023 530
rect 2027 526 2031 530
rect 2035 526 2095 530
rect 2099 526 2103 530
rect 2107 526 2167 530
rect 2171 526 2191 530
rect 2195 526 2239 530
rect 2243 526 2287 530
rect 2291 526 2311 530
rect 2315 526 2359 530
rect 2363 526 2407 530
rect 2411 526 2435 530
rect 1257 525 2435 526
rect 2441 525 2442 531
rect 96 473 97 479
rect 103 478 1263 479
rect 103 474 111 478
rect 115 474 151 478
rect 155 474 223 478
rect 227 474 239 478
rect 243 474 279 478
rect 283 474 287 478
rect 291 474 327 478
rect 331 474 351 478
rect 355 474 383 478
rect 387 474 415 478
rect 419 474 439 478
rect 443 474 479 478
rect 483 474 503 478
rect 507 474 551 478
rect 555 474 567 478
rect 571 474 623 478
rect 627 474 631 478
rect 635 474 695 478
rect 699 474 759 478
rect 763 474 767 478
rect 771 474 823 478
rect 827 474 839 478
rect 843 474 887 478
rect 891 474 919 478
rect 923 474 951 478
rect 955 474 999 478
rect 1003 474 1015 478
rect 1019 474 1079 478
rect 1083 474 1239 478
rect 1243 474 1263 478
rect 103 473 1263 474
rect 1269 473 1270 479
rect 1262 457 1263 463
rect 1269 462 2447 463
rect 1269 458 1279 462
rect 1283 458 1303 462
rect 1307 458 1343 462
rect 1347 458 1383 462
rect 1387 458 1407 462
rect 1411 458 1447 462
rect 1451 458 1487 462
rect 1491 458 1535 462
rect 1539 458 1591 462
rect 1595 458 1631 462
rect 1635 458 1647 462
rect 1651 458 1711 462
rect 1715 458 1735 462
rect 1739 458 1783 462
rect 1787 458 1831 462
rect 1835 458 1863 462
rect 1867 458 1919 462
rect 1923 458 1943 462
rect 1947 458 1999 462
rect 2003 458 2023 462
rect 2027 458 2071 462
rect 2075 458 2103 462
rect 2107 458 2135 462
rect 2139 458 2191 462
rect 2195 458 2199 462
rect 2203 458 2255 462
rect 2259 458 2287 462
rect 2291 458 2319 462
rect 2323 458 2359 462
rect 2363 458 2407 462
rect 2411 458 2447 462
rect 1269 457 2447 458
rect 2453 457 2454 463
rect 84 401 85 407
rect 91 406 1251 407
rect 91 402 111 406
rect 115 402 143 406
rect 147 402 183 406
rect 187 402 223 406
rect 227 402 239 406
rect 243 402 271 406
rect 275 402 279 406
rect 283 402 327 406
rect 331 402 335 406
rect 339 402 383 406
rect 387 402 399 406
rect 403 402 439 406
rect 443 402 471 406
rect 475 402 503 406
rect 507 402 543 406
rect 547 402 567 406
rect 571 402 615 406
rect 619 402 631 406
rect 635 402 687 406
rect 691 402 695 406
rect 699 402 751 406
rect 755 402 759 406
rect 763 402 807 406
rect 811 402 823 406
rect 827 402 863 406
rect 867 402 887 406
rect 891 402 919 406
rect 923 402 951 406
rect 955 402 975 406
rect 979 402 1015 406
rect 1019 402 1031 406
rect 1035 402 1239 406
rect 1243 402 1251 406
rect 91 401 1251 402
rect 1257 401 1258 407
rect 1250 389 1251 395
rect 1257 394 2435 395
rect 1257 390 1279 394
rect 1283 390 1303 394
rect 1307 390 1343 394
rect 1347 390 1359 394
rect 1363 390 1383 394
rect 1387 390 1399 394
rect 1403 390 1439 394
rect 1443 390 1447 394
rect 1451 390 1487 394
rect 1491 390 1535 394
rect 1539 390 1543 394
rect 1547 390 1607 394
rect 1611 390 1631 394
rect 1635 390 1679 394
rect 1683 390 1735 394
rect 1739 390 1759 394
rect 1763 390 1831 394
rect 1835 390 1839 394
rect 1843 390 1919 394
rect 1923 390 1999 394
rect 2003 390 2071 394
rect 2075 390 2079 394
rect 2083 390 2135 394
rect 2139 390 2159 394
rect 2163 390 2199 394
rect 2203 390 2247 394
rect 2251 390 2255 394
rect 2259 390 2319 394
rect 2323 390 2335 394
rect 2339 390 2359 394
rect 2363 390 2407 394
rect 2411 390 2435 394
rect 1257 389 2435 390
rect 2441 389 2442 395
rect 96 325 97 331
rect 103 330 1263 331
rect 103 326 111 330
rect 115 326 135 330
rect 139 326 143 330
rect 147 326 175 330
rect 179 326 183 330
rect 187 326 215 330
rect 219 326 223 330
rect 227 326 255 330
rect 259 326 271 330
rect 275 326 295 330
rect 299 326 335 330
rect 339 326 391 330
rect 395 326 399 330
rect 403 326 447 330
rect 451 326 471 330
rect 475 326 495 330
rect 499 326 543 330
rect 547 326 591 330
rect 595 326 615 330
rect 619 326 639 330
rect 643 326 687 330
rect 691 326 735 330
rect 739 326 751 330
rect 755 326 783 330
rect 787 326 807 330
rect 811 326 839 330
rect 843 326 863 330
rect 867 326 919 330
rect 923 326 975 330
rect 979 326 1031 330
rect 1035 326 1239 330
rect 1243 326 1263 330
rect 103 325 1263 326
rect 1269 325 1270 331
rect 1262 313 1263 319
rect 1269 318 2447 319
rect 1269 314 1279 318
rect 1283 314 1359 318
rect 1363 314 1399 318
rect 1403 314 1439 318
rect 1443 314 1487 318
rect 1491 314 1511 318
rect 1515 314 1543 318
rect 1547 314 1551 318
rect 1555 314 1591 318
rect 1595 314 1607 318
rect 1611 314 1631 318
rect 1635 314 1671 318
rect 1675 314 1679 318
rect 1683 314 1711 318
rect 1715 314 1751 318
rect 1755 314 1759 318
rect 1763 314 1791 318
rect 1795 314 1839 318
rect 1843 314 1903 318
rect 1907 314 1919 318
rect 1923 314 1967 318
rect 1971 314 1999 318
rect 2003 314 2039 318
rect 2043 314 2079 318
rect 2083 314 2119 318
rect 2123 314 2159 318
rect 2163 314 2199 318
rect 2203 314 2247 318
rect 2251 314 2279 318
rect 2283 314 2335 318
rect 2339 314 2359 318
rect 2363 314 2407 318
rect 2411 314 2447 318
rect 1269 313 2447 314
rect 2453 313 2454 319
rect 84 249 85 255
rect 91 254 1251 255
rect 91 250 111 254
rect 115 250 135 254
rect 139 250 175 254
rect 179 250 215 254
rect 219 250 223 254
rect 227 250 255 254
rect 259 250 295 254
rect 299 250 311 254
rect 315 250 335 254
rect 339 250 391 254
rect 395 250 447 254
rect 451 250 463 254
rect 467 250 495 254
rect 499 250 527 254
rect 531 250 543 254
rect 547 250 591 254
rect 595 250 639 254
rect 643 250 647 254
rect 651 250 687 254
rect 691 250 695 254
rect 699 250 735 254
rect 739 250 783 254
rect 787 250 831 254
rect 835 250 839 254
rect 843 250 879 254
rect 883 250 927 254
rect 931 250 975 254
rect 979 250 1023 254
rect 1027 250 1239 254
rect 1243 250 1251 254
rect 91 249 1251 250
rect 1257 249 1258 255
rect 1250 247 1258 249
rect 1250 241 1251 247
rect 1257 246 2435 247
rect 1257 242 1279 246
rect 1283 242 1367 246
rect 1371 242 1407 246
rect 1411 242 1455 246
rect 1459 242 1511 246
rect 1515 242 1551 246
rect 1555 242 1567 246
rect 1571 242 1591 246
rect 1595 242 1631 246
rect 1635 242 1671 246
rect 1675 242 1703 246
rect 1707 242 1711 246
rect 1715 242 1751 246
rect 1755 242 1775 246
rect 1779 242 1791 246
rect 1795 242 1839 246
rect 1843 242 1855 246
rect 1859 242 1903 246
rect 1907 242 1943 246
rect 1947 242 1967 246
rect 1971 242 2031 246
rect 2035 242 2039 246
rect 2043 242 2119 246
rect 2123 242 2199 246
rect 2203 242 2207 246
rect 2211 242 2279 246
rect 2283 242 2295 246
rect 2299 242 2359 246
rect 2363 242 2407 246
rect 2411 242 2435 246
rect 1257 241 2435 242
rect 2441 241 2442 247
rect 1262 165 1263 171
rect 1269 170 2447 171
rect 1269 166 1279 170
rect 1283 166 1303 170
rect 1307 166 1343 170
rect 1347 166 1367 170
rect 1371 166 1383 170
rect 1387 166 1407 170
rect 1411 166 1423 170
rect 1427 166 1455 170
rect 1459 166 1463 170
rect 1467 166 1511 170
rect 1515 166 1519 170
rect 1523 166 1567 170
rect 1571 166 1583 170
rect 1587 166 1631 170
rect 1635 166 1647 170
rect 1651 166 1703 170
rect 1707 166 1711 170
rect 1715 166 1775 170
rect 1779 166 1831 170
rect 1835 166 1855 170
rect 1859 166 1887 170
rect 1891 166 1935 170
rect 1939 166 1943 170
rect 1947 166 1975 170
rect 1979 166 2015 170
rect 2019 166 2031 170
rect 2035 166 2055 170
rect 2059 166 2095 170
rect 2099 166 2119 170
rect 2123 166 2143 170
rect 2147 166 2191 170
rect 2195 166 2207 170
rect 2211 166 2239 170
rect 2243 166 2279 170
rect 2283 166 2295 170
rect 2299 166 2319 170
rect 2323 166 2359 170
rect 2363 166 2407 170
rect 2411 166 2447 170
rect 1269 165 2447 166
rect 2453 165 2454 171
rect 96 149 97 155
rect 103 154 1263 155
rect 103 150 111 154
rect 115 150 135 154
rect 139 150 151 154
rect 155 150 191 154
rect 195 150 223 154
rect 227 150 231 154
rect 235 150 271 154
rect 275 150 311 154
rect 315 150 351 154
rect 355 150 391 154
rect 395 150 431 154
rect 435 150 463 154
rect 467 150 471 154
rect 475 150 511 154
rect 515 150 527 154
rect 531 150 551 154
rect 555 150 591 154
rect 595 150 631 154
rect 635 150 647 154
rect 651 150 671 154
rect 675 150 695 154
rect 699 150 711 154
rect 715 150 735 154
rect 739 150 751 154
rect 755 150 783 154
rect 787 150 791 154
rect 795 150 831 154
rect 835 150 871 154
rect 875 150 879 154
rect 883 150 911 154
rect 915 150 927 154
rect 931 150 951 154
rect 955 150 975 154
rect 979 150 991 154
rect 995 150 1023 154
rect 1027 150 1031 154
rect 1035 150 1071 154
rect 1075 150 1111 154
rect 1115 150 1151 154
rect 1155 150 1191 154
rect 1195 150 1239 154
rect 1243 150 1263 154
rect 103 149 1263 150
rect 1269 149 1270 155
rect 650 116 656 117
rect 1038 116 1044 117
rect 650 112 651 116
rect 655 112 1039 116
rect 1043 112 1044 116
rect 650 111 656 112
rect 1038 111 1044 112
rect 1250 97 1251 103
rect 1257 102 2435 103
rect 1257 98 1279 102
rect 1283 98 1303 102
rect 1307 98 1343 102
rect 1347 98 1383 102
rect 1387 98 1423 102
rect 1427 98 1463 102
rect 1467 98 1519 102
rect 1523 98 1583 102
rect 1587 98 1647 102
rect 1651 98 1711 102
rect 1715 98 1775 102
rect 1779 98 1831 102
rect 1835 98 1887 102
rect 1891 98 1935 102
rect 1939 98 1975 102
rect 1979 98 2015 102
rect 2019 98 2055 102
rect 2059 98 2095 102
rect 2099 98 2143 102
rect 2147 98 2191 102
rect 2195 98 2239 102
rect 2243 98 2279 102
rect 2283 98 2319 102
rect 2323 98 2359 102
rect 2363 98 2407 102
rect 2411 98 2435 102
rect 1257 97 2435 98
rect 2441 97 2442 103
rect 84 81 85 87
rect 91 86 1251 87
rect 91 82 111 86
rect 115 82 151 86
rect 155 82 191 86
rect 195 82 231 86
rect 235 82 271 86
rect 275 82 311 86
rect 315 82 351 86
rect 355 82 391 86
rect 395 82 431 86
rect 435 82 471 86
rect 475 82 511 86
rect 515 82 551 86
rect 555 82 591 86
rect 595 82 631 86
rect 635 82 671 86
rect 675 82 711 86
rect 715 82 751 86
rect 755 82 791 86
rect 795 82 831 86
rect 835 82 871 86
rect 875 82 911 86
rect 915 82 951 86
rect 955 82 991 86
rect 995 82 1031 86
rect 1035 82 1071 86
rect 1075 82 1111 86
rect 1115 82 1151 86
rect 1155 82 1191 86
rect 1195 82 1239 86
rect 1243 82 1251 86
rect 91 81 1251 82
rect 1257 81 1258 87
<< m5c >>
rect 97 2489 103 2495
rect 1263 2489 1269 2495
rect 85 2413 91 2419
rect 1251 2413 1257 2419
rect 97 2341 103 2347
rect 1263 2341 1269 2347
rect 1251 2277 1257 2283
rect 2435 2277 2441 2283
rect 85 2265 91 2271
rect 1251 2265 1257 2271
rect 97 2197 103 2203
rect 1263 2197 1269 2203
rect 1251 2133 1257 2139
rect 2435 2133 2441 2139
rect 85 2121 91 2127
rect 1251 2121 1257 2127
rect 1263 2065 1269 2071
rect 2447 2065 2453 2071
rect 97 2049 103 2055
rect 1263 2049 1269 2055
rect 1251 1997 1257 2003
rect 2435 1997 2441 2003
rect 85 1981 91 1987
rect 1251 1981 1257 1987
rect 1263 1925 1269 1931
rect 2447 1925 2453 1931
rect 97 1909 103 1915
rect 1263 1909 1269 1915
rect 1251 1849 1257 1855
rect 2435 1849 2441 1855
rect 85 1837 91 1843
rect 1251 1837 1257 1843
rect 97 1769 103 1775
rect 1263 1769 1269 1775
rect 85 1697 91 1703
rect 1251 1697 1257 1703
rect 97 1625 103 1631
rect 1263 1625 1269 1631
rect 85 1553 91 1559
rect 1251 1553 1257 1559
rect 97 1481 103 1487
rect 1263 1481 1269 1487
rect 1263 1469 1269 1475
rect 2447 1469 2453 1475
rect 85 1409 91 1415
rect 1251 1409 1257 1415
rect 1251 1401 1257 1407
rect 2435 1401 2441 1407
rect 97 1337 103 1343
rect 1263 1337 1269 1343
rect 1263 1329 1269 1335
rect 2447 1329 2453 1335
rect 85 1265 91 1271
rect 1251 1265 1257 1271
rect 1251 1257 1257 1263
rect 2435 1257 2441 1263
rect 97 1189 103 1195
rect 1263 1189 1269 1195
rect 85 1121 91 1127
rect 1251 1121 1257 1127
rect 1251 1109 1257 1115
rect 2435 1109 2441 1115
rect 97 1049 103 1055
rect 1263 1049 1269 1055
rect 1263 1029 1269 1035
rect 2447 1029 2453 1035
rect 85 969 91 975
rect 1251 969 1257 975
rect 1251 953 1257 959
rect 2435 953 2441 959
rect 97 893 103 899
rect 1263 893 1269 899
rect 1263 877 1269 883
rect 2447 877 2453 883
rect 85 825 91 831
rect 1251 825 1257 831
rect 1251 805 1257 811
rect 2435 805 2441 811
rect 97 757 103 763
rect 1263 757 1269 763
rect 1263 737 1269 743
rect 2447 737 2453 743
rect 85 681 91 687
rect 1251 681 1257 687
rect 1251 669 1257 675
rect 2435 669 2441 675
rect 97 613 103 619
rect 1263 613 1269 619
rect 1263 593 1269 599
rect 2447 593 2453 599
rect 85 541 91 547
rect 1251 541 1257 547
rect 1251 525 1257 531
rect 2435 525 2441 531
rect 97 473 103 479
rect 1263 473 1269 479
rect 1263 457 1269 463
rect 2447 457 2453 463
rect 85 401 91 407
rect 1251 401 1257 407
rect 1251 389 1257 395
rect 2435 389 2441 395
rect 97 325 103 331
rect 1263 325 1269 331
rect 1263 313 1269 319
rect 2447 313 2453 319
rect 85 249 91 255
rect 1251 249 1257 255
rect 1251 241 1257 247
rect 2435 241 2441 247
rect 1263 165 1269 171
rect 2447 165 2453 171
rect 97 149 103 155
rect 1263 149 1269 155
rect 1251 97 1257 103
rect 2435 97 2441 103
rect 85 81 91 87
rect 1251 81 1257 87
<< m5 >>
rect 84 2419 92 2520
rect 84 2413 85 2419
rect 91 2413 92 2419
rect 84 2271 92 2413
rect 84 2265 85 2271
rect 91 2265 92 2271
rect 84 2127 92 2265
rect 84 2121 85 2127
rect 91 2121 92 2127
rect 84 1987 92 2121
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1843 92 1981
rect 84 1837 85 1843
rect 91 1837 92 1843
rect 84 1703 92 1837
rect 84 1697 85 1703
rect 91 1697 92 1703
rect 84 1559 92 1697
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1415 92 1553
rect 84 1409 85 1415
rect 91 1409 92 1415
rect 84 1271 92 1409
rect 84 1265 85 1271
rect 91 1265 92 1271
rect 84 1127 92 1265
rect 84 1121 85 1127
rect 91 1121 92 1127
rect 84 975 92 1121
rect 84 969 85 975
rect 91 969 92 975
rect 84 831 92 969
rect 84 825 85 831
rect 91 825 92 831
rect 84 687 92 825
rect 84 681 85 687
rect 91 681 92 687
rect 84 547 92 681
rect 84 541 85 547
rect 91 541 92 547
rect 84 407 92 541
rect 84 401 85 407
rect 91 401 92 407
rect 84 255 92 401
rect 84 249 85 255
rect 91 249 92 255
rect 84 87 92 249
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2495 104 2520
rect 96 2489 97 2495
rect 103 2489 104 2495
rect 96 2347 104 2489
rect 96 2341 97 2347
rect 103 2341 104 2347
rect 96 2203 104 2341
rect 96 2197 97 2203
rect 103 2197 104 2203
rect 96 2055 104 2197
rect 96 2049 97 2055
rect 103 2049 104 2055
rect 96 1915 104 2049
rect 96 1909 97 1915
rect 103 1909 104 1915
rect 96 1775 104 1909
rect 96 1769 97 1775
rect 103 1769 104 1775
rect 96 1631 104 1769
rect 96 1625 97 1631
rect 103 1625 104 1631
rect 96 1487 104 1625
rect 96 1481 97 1487
rect 103 1481 104 1487
rect 96 1343 104 1481
rect 96 1337 97 1343
rect 103 1337 104 1343
rect 96 1195 104 1337
rect 96 1189 97 1195
rect 103 1189 104 1195
rect 96 1055 104 1189
rect 96 1049 97 1055
rect 103 1049 104 1055
rect 96 899 104 1049
rect 96 893 97 899
rect 103 893 104 899
rect 96 763 104 893
rect 96 757 97 763
rect 103 757 104 763
rect 96 619 104 757
rect 96 613 97 619
rect 103 613 104 619
rect 96 479 104 613
rect 96 473 97 479
rect 103 473 104 479
rect 96 331 104 473
rect 96 325 97 331
rect 103 325 104 331
rect 96 155 104 325
rect 96 149 97 155
rect 103 149 104 155
rect 96 72 104 149
rect 1250 2419 1258 2520
rect 1250 2413 1251 2419
rect 1257 2413 1258 2419
rect 1250 2283 1258 2413
rect 1250 2277 1251 2283
rect 1257 2277 1258 2283
rect 1250 2271 1258 2277
rect 1250 2265 1251 2271
rect 1257 2265 1258 2271
rect 1250 2139 1258 2265
rect 1250 2133 1251 2139
rect 1257 2133 1258 2139
rect 1250 2127 1258 2133
rect 1250 2121 1251 2127
rect 1257 2121 1258 2127
rect 1250 2003 1258 2121
rect 1250 1997 1251 2003
rect 1257 1997 1258 2003
rect 1250 1987 1258 1997
rect 1250 1981 1251 1987
rect 1257 1981 1258 1987
rect 1250 1855 1258 1981
rect 1250 1849 1251 1855
rect 1257 1849 1258 1855
rect 1250 1843 1258 1849
rect 1250 1837 1251 1843
rect 1257 1837 1258 1843
rect 1250 1703 1258 1837
rect 1250 1697 1251 1703
rect 1257 1697 1258 1703
rect 1250 1559 1258 1697
rect 1250 1553 1251 1559
rect 1257 1553 1258 1559
rect 1250 1415 1258 1553
rect 1250 1409 1251 1415
rect 1257 1409 1258 1415
rect 1250 1407 1258 1409
rect 1250 1401 1251 1407
rect 1257 1401 1258 1407
rect 1250 1271 1258 1401
rect 1250 1265 1251 1271
rect 1257 1265 1258 1271
rect 1250 1263 1258 1265
rect 1250 1257 1251 1263
rect 1257 1257 1258 1263
rect 1250 1127 1258 1257
rect 1250 1121 1251 1127
rect 1257 1121 1258 1127
rect 1250 1115 1258 1121
rect 1250 1109 1251 1115
rect 1257 1109 1258 1115
rect 1250 975 1258 1109
rect 1250 969 1251 975
rect 1257 969 1258 975
rect 1250 959 1258 969
rect 1250 953 1251 959
rect 1257 953 1258 959
rect 1250 831 1258 953
rect 1250 825 1251 831
rect 1257 825 1258 831
rect 1250 811 1258 825
rect 1250 805 1251 811
rect 1257 805 1258 811
rect 1250 687 1258 805
rect 1250 681 1251 687
rect 1257 681 1258 687
rect 1250 675 1258 681
rect 1250 669 1251 675
rect 1257 669 1258 675
rect 1250 547 1258 669
rect 1250 541 1251 547
rect 1257 541 1258 547
rect 1250 531 1258 541
rect 1250 525 1251 531
rect 1257 525 1258 531
rect 1250 407 1258 525
rect 1250 401 1251 407
rect 1257 401 1258 407
rect 1250 395 1258 401
rect 1250 389 1251 395
rect 1257 389 1258 395
rect 1250 255 1258 389
rect 1250 249 1251 255
rect 1257 249 1258 255
rect 1250 247 1258 249
rect 1250 241 1251 247
rect 1257 241 1258 247
rect 1250 103 1258 241
rect 1250 97 1251 103
rect 1257 97 1258 103
rect 1250 87 1258 97
rect 1250 81 1251 87
rect 1257 81 1258 87
rect 1250 72 1258 81
rect 1262 2495 1270 2520
rect 1262 2489 1263 2495
rect 1269 2489 1270 2495
rect 1262 2347 1270 2489
rect 1262 2341 1263 2347
rect 1269 2341 1270 2347
rect 1262 2203 1270 2341
rect 1262 2197 1263 2203
rect 1269 2197 1270 2203
rect 1262 2071 1270 2197
rect 1262 2065 1263 2071
rect 1269 2065 1270 2071
rect 1262 2055 1270 2065
rect 1262 2049 1263 2055
rect 1269 2049 1270 2055
rect 1262 1931 1270 2049
rect 1262 1925 1263 1931
rect 1269 1925 1270 1931
rect 1262 1915 1270 1925
rect 1262 1909 1263 1915
rect 1269 1909 1270 1915
rect 1262 1775 1270 1909
rect 1262 1769 1263 1775
rect 1269 1769 1270 1775
rect 1262 1631 1270 1769
rect 1262 1625 1263 1631
rect 1269 1625 1270 1631
rect 1262 1487 1270 1625
rect 1262 1481 1263 1487
rect 1269 1481 1270 1487
rect 1262 1475 1270 1481
rect 1262 1469 1263 1475
rect 1269 1469 1270 1475
rect 1262 1343 1270 1469
rect 1262 1337 1263 1343
rect 1269 1337 1270 1343
rect 1262 1335 1270 1337
rect 1262 1329 1263 1335
rect 1269 1329 1270 1335
rect 1262 1195 1270 1329
rect 1262 1189 1263 1195
rect 1269 1189 1270 1195
rect 1262 1055 1270 1189
rect 1262 1049 1263 1055
rect 1269 1049 1270 1055
rect 1262 1035 1270 1049
rect 1262 1029 1263 1035
rect 1269 1029 1270 1035
rect 1262 899 1270 1029
rect 1262 893 1263 899
rect 1269 893 1270 899
rect 1262 883 1270 893
rect 1262 877 1263 883
rect 1269 877 1270 883
rect 1262 763 1270 877
rect 1262 757 1263 763
rect 1269 757 1270 763
rect 1262 743 1270 757
rect 1262 737 1263 743
rect 1269 737 1270 743
rect 1262 619 1270 737
rect 1262 613 1263 619
rect 1269 613 1270 619
rect 1262 599 1270 613
rect 1262 593 1263 599
rect 1269 593 1270 599
rect 1262 479 1270 593
rect 1262 473 1263 479
rect 1269 473 1270 479
rect 1262 463 1270 473
rect 1262 457 1263 463
rect 1269 457 1270 463
rect 1262 331 1270 457
rect 1262 325 1263 331
rect 1269 325 1270 331
rect 1262 319 1270 325
rect 1262 313 1263 319
rect 1269 313 1270 319
rect 1262 171 1270 313
rect 1262 165 1263 171
rect 1269 165 1270 171
rect 1262 155 1270 165
rect 1262 149 1263 155
rect 1269 149 1270 155
rect 1262 72 1270 149
rect 2434 2283 2442 2520
rect 2434 2277 2435 2283
rect 2441 2277 2442 2283
rect 2434 2139 2442 2277
rect 2434 2133 2435 2139
rect 2441 2133 2442 2139
rect 2434 2003 2442 2133
rect 2434 1997 2435 2003
rect 2441 1997 2442 2003
rect 2434 1855 2442 1997
rect 2434 1849 2435 1855
rect 2441 1849 2442 1855
rect 2434 1407 2442 1849
rect 2434 1401 2435 1407
rect 2441 1401 2442 1407
rect 2434 1263 2442 1401
rect 2434 1257 2435 1263
rect 2441 1257 2442 1263
rect 2434 1115 2442 1257
rect 2434 1109 2435 1115
rect 2441 1109 2442 1115
rect 2434 959 2442 1109
rect 2434 953 2435 959
rect 2441 953 2442 959
rect 2434 811 2442 953
rect 2434 805 2435 811
rect 2441 805 2442 811
rect 2434 675 2442 805
rect 2434 669 2435 675
rect 2441 669 2442 675
rect 2434 531 2442 669
rect 2434 525 2435 531
rect 2441 525 2442 531
rect 2434 395 2442 525
rect 2434 389 2435 395
rect 2441 389 2442 395
rect 2434 247 2442 389
rect 2434 241 2435 247
rect 2441 241 2442 247
rect 2434 103 2442 241
rect 2434 97 2435 103
rect 2441 97 2442 103
rect 2434 72 2442 97
rect 2446 2071 2454 2520
rect 2446 2065 2447 2071
rect 2453 2065 2454 2071
rect 2446 1931 2454 2065
rect 2446 1925 2447 1931
rect 2453 1925 2454 1931
rect 2446 1475 2454 1925
rect 2446 1469 2447 1475
rect 2453 1469 2454 1475
rect 2446 1335 2454 1469
rect 2446 1329 2447 1335
rect 2453 1329 2454 1335
rect 2446 1035 2454 1329
rect 2446 1029 2447 1035
rect 2453 1029 2454 1035
rect 2446 883 2454 1029
rect 2446 877 2447 883
rect 2453 877 2454 883
rect 2446 743 2454 877
rect 2446 737 2447 743
rect 2453 737 2454 743
rect 2446 599 2454 737
rect 2446 593 2447 599
rect 2453 593 2454 599
rect 2446 463 2454 593
rect 2446 457 2447 463
rect 2453 457 2454 463
rect 2446 319 2454 457
rect 2446 313 2447 319
rect 2453 313 2454 319
rect 2446 171 2454 313
rect 2446 165 2447 171
rect 2453 165 2454 171
rect 2446 72 2454 165
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__131
timestamp 1731220651
transform 1 0 2400 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220651
transform 1 0 1272 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220651
transform 1 0 2400 0 -1 2412
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220651
transform 1 0 1272 0 -1 2412
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220651
transform 1 0 2400 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220651
transform 1 0 1272 0 1 2288
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220651
transform 1 0 2400 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220651
transform 1 0 1272 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220651
transform 1 0 2400 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220651
transform 1 0 1272 0 1 2144
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220651
transform 1 0 2400 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220651
transform 1 0 1272 0 -1 2128
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220651
transform 1 0 2400 0 1 2008
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220651
transform 1 0 1272 0 1 2008
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220651
transform 1 0 2400 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220651
transform 1 0 1272 0 -1 1992
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220651
transform 1 0 2400 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220651
transform 1 0 1272 0 1 1868
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220651
transform 1 0 2400 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220651
transform 1 0 1272 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220651
transform 1 0 2400 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220651
transform 1 0 1272 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220651
transform 1 0 2400 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220651
transform 1 0 1272 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220651
transform 1 0 2400 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220651
transform 1 0 1272 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220651
transform 1 0 2400 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220651
transform 1 0 1272 0 -1 1552
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220651
transform 1 0 2400 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220651
transform 1 0 1272 0 1 1412
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220651
transform 1 0 2400 0 -1 1396
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220651
transform 1 0 1272 0 -1 1396
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220651
transform 1 0 2400 0 1 1272
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220651
transform 1 0 1272 0 1 1272
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220651
transform 1 0 2400 0 -1 1252
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220651
transform 1 0 1272 0 -1 1252
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220651
transform 1 0 2400 0 1 1128
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220651
transform 1 0 1272 0 1 1128
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220651
transform 1 0 2400 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220651
transform 1 0 1272 0 -1 1104
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220651
transform 1 0 2400 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220651
transform 1 0 1272 0 1 972
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220651
transform 1 0 2400 0 -1 948
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220651
transform 1 0 1272 0 -1 948
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220651
transform 1 0 2400 0 1 820
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220651
transform 1 0 1272 0 1 820
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220651
transform 1 0 2400 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220651
transform 1 0 1272 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220651
transform 1 0 2400 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220651
transform 1 0 1272 0 1 680
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220651
transform 1 0 2400 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220651
transform 1 0 1272 0 -1 664
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220651
transform 1 0 2400 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220651
transform 1 0 1272 0 1 536
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220651
transform 1 0 2400 0 -1 520
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220651
transform 1 0 1272 0 -1 520
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220651
transform 1 0 2400 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220651
transform 1 0 1272 0 1 400
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220651
transform 1 0 2400 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220651
transform 1 0 1272 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220651
transform 1 0 2400 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220651
transform 1 0 1272 0 1 256
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220651
transform 1 0 2400 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220651
transform 1 0 1272 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220651
transform 1 0 2400 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220651
transform 1 0 1272 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220651
transform 1 0 1232 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220651
transform 1 0 104 0 1 2432
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220651
transform 1 0 1232 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220651
transform 1 0 104 0 -1 2408
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220651
transform 1 0 1232 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220651
transform 1 0 104 0 1 2284
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220651
transform 1 0 1232 0 -1 2260
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220651
transform 1 0 104 0 -1 2260
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220651
transform 1 0 1232 0 1 2140
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220651
transform 1 0 104 0 1 2140
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220651
transform 1 0 1232 0 -1 2116
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220651
transform 1 0 104 0 -1 2116
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220651
transform 1 0 1232 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220651
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220651
transform 1 0 1232 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220651
transform 1 0 104 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220651
transform 1 0 1232 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220651
transform 1 0 104 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220651
transform 1 0 1232 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220651
transform 1 0 104 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220651
transform 1 0 1232 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220651
transform 1 0 104 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220651
transform 1 0 1232 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220651
transform 1 0 104 0 -1 1692
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220651
transform 1 0 1232 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220651
transform 1 0 104 0 1 1568
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220651
transform 1 0 1232 0 -1 1548
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220651
transform 1 0 104 0 -1 1548
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220651
transform 1 0 1232 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220651
transform 1 0 104 0 1 1424
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220651
transform 1 0 1232 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220651
transform 1 0 104 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220651
transform 1 0 1232 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220651
transform 1 0 104 0 1 1280
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220651
transform 1 0 1232 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220651
transform 1 0 104 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220651
transform 1 0 1232 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220651
transform 1 0 104 0 1 1132
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220651
transform 1 0 1232 0 -1 1116
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220651
transform 1 0 104 0 -1 1116
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220651
transform 1 0 1232 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220651
transform 1 0 104 0 1 992
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220651
transform 1 0 1232 0 -1 964
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220651
transform 1 0 104 0 -1 964
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220651
transform 1 0 1232 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220651
transform 1 0 104 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220651
transform 1 0 1232 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220651
transform 1 0 104 0 -1 820
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220651
transform 1 0 1232 0 1 700
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220651
transform 1 0 104 0 1 700
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220651
transform 1 0 1232 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220651
transform 1 0 104 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220651
transform 1 0 1232 0 1 556
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220651
transform 1 0 104 0 1 556
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220651
transform 1 0 1232 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220651
transform 1 0 104 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220651
transform 1 0 1232 0 1 416
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220651
transform 1 0 104 0 1 416
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220651
transform 1 0 1232 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220651
transform 1 0 104 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220651
transform 1 0 1232 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220651
transform 1 0 104 0 1 268
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220651
transform 1 0 1232 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220651
transform 1 0 104 0 -1 244
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220651
transform 1 0 1232 0 1 92
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220651
transform 1 0 104 0 1 92
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X2  tst_5999_6
timestamp 1731220651
transform 1 0 144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5998_6
timestamp 1731220651
transform 1 0 184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5997_6
timestamp 1731220651
transform 1 0 224 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5996_6
timestamp 1731220651
transform 1 0 264 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5995_6
timestamp 1731220651
transform 1 0 304 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5994_6
timestamp 1731220651
transform 1 0 344 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5993_6
timestamp 1731220651
transform 1 0 384 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5992_6
timestamp 1731220651
transform 1 0 424 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5991_6
timestamp 1731220651
transform 1 0 464 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5990_6
timestamp 1731220651
transform 1 0 504 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5989_6
timestamp 1731220651
transform 1 0 544 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5988_6
timestamp 1731220651
transform 1 0 584 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5987_6
timestamp 1731220651
transform 1 0 216 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5986_6
timestamp 1731220651
transform 1 0 304 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5985_6
timestamp 1731220651
transform 1 0 384 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5984_6
timestamp 1731220651
transform 1 0 456 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5983_6
timestamp 1731220651
transform 1 0 520 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5982_6
timestamp 1731220651
transform 1 0 584 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5981_6
timestamp 1731220651
transform 1 0 640 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5980_6
timestamp 1731220651
transform 1 0 488 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5979_6
timestamp 1731220651
transform 1 0 536 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5978_6
timestamp 1731220651
transform 1 0 832 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5977_6
timestamp 1731220651
transform 1 0 912 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5976_6
timestamp 1731220651
transform 1 0 968 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5975_6
timestamp 1731220651
transform 1 0 1024 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5974_6
timestamp 1731220651
transform 1 0 1008 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5973_6
timestamp 1731220651
transform 1 0 944 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5972_6
timestamp 1731220651
transform 1 0 912 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5971_6
timestamp 1731220651
transform 1 0 992 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5970_6
timestamp 1731220651
transform 1 0 1072 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5969_6
timestamp 1731220651
transform 1 0 1008 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5968_6
timestamp 1731220651
transform 1 0 944 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5967_6
timestamp 1731220651
transform 1 0 872 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5966_6
timestamp 1731220651
transform 1 0 896 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5965_6
timestamp 1731220651
transform 1 0 960 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5964_6
timestamp 1731220651
transform 1 0 1016 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5963_6
timestamp 1731220651
transform 1 0 1072 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5962_6
timestamp 1731220651
transform 1 0 1136 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5961_6
timestamp 1731220651
transform 1 0 1184 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5960_6
timestamp 1731220651
transform 1 0 1184 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5959_6
timestamp 1731220651
transform 1 0 1080 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5958_6
timestamp 1731220651
transform 1 0 1144 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5957_6
timestamp 1731220651
transform 1 0 1184 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5956_6
timestamp 1731220651
transform 1 0 1296 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5955_6
timestamp 1731220651
transform 1 0 1360 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5954_6
timestamp 1731220651
transform 1 0 1400 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5953_6
timestamp 1731220651
transform 1 0 1336 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5952_6
timestamp 1731220651
transform 1 0 1296 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5951_6
timestamp 1731220651
transform 1 0 1328 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5950_6
timestamp 1731220651
transform 1 0 1368 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5949_6
timestamp 1731220651
transform 1 0 1408 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5948_6
timestamp 1731220651
transform 1 0 1312 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5947_6
timestamp 1731220651
transform 1 0 1352 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5946_6
timestamp 1731220651
transform 1 0 1392 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5945_6
timestamp 1731220651
transform 1 0 1536 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5944_6
timestamp 1731220651
transform 1 0 1632 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5943_6
timestamp 1731220651
transform 1 0 1728 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5942_6
timestamp 1731220651
transform 1 0 1832 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5941_6
timestamp 1731220651
transform 1 0 1744 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5940_6
timestamp 1731220651
transform 1 0 1672 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5939_6
timestamp 1731220651
transform 1 0 1600 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5938_6
timestamp 1731220651
transform 1 0 1616 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5937_6
timestamp 1731220651
transform 1 0 1688 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5936_6
timestamp 1731220651
transform 1 0 1688 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5935_6
timestamp 1731220651
transform 1 0 1608 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5934_6
timestamp 1731220651
transform 1 0 1632 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5933_6
timestamp 1731220651
transform 1 0 1680 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5932_6
timestamp 1731220651
transform 1 0 1736 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5931_6
timestamp 1731220651
transform 1 0 1792 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5930_6
timestamp 1731220651
transform 1 0 1864 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5929_6
timestamp 1731220651
transform 1 0 1848 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5928_6
timestamp 1731220651
transform 1 0 1904 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5927_6
timestamp 1731220651
transform 1 0 1936 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5926_6
timestamp 1731220651
transform 1 0 1856 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5925_6
timestamp 1731220651
transform 1 0 1776 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5924_6
timestamp 1731220651
transform 1 0 1824 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5923_6
timestamp 1731220651
transform 1 0 1912 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5922_6
timestamp 1731220651
transform 1 0 1992 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5921_6
timestamp 1731220651
transform 1 0 1832 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5920_6
timestamp 1731220651
transform 1 0 1752 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5919_6
timestamp 1731220651
transform 1 0 1832 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5918_6
timestamp 1731220651
transform 1 0 1896 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5917_6
timestamp 1731220651
transform 1 0 1960 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5916_6
timestamp 1731220651
transform 1 0 2032 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5915_6
timestamp 1731220651
transform 1 0 2112 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5914_6
timestamp 1731220651
transform 1 0 1768 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5913_6
timestamp 1731220651
transform 1 0 1848 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5912_6
timestamp 1731220651
transform 1 0 1936 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5911_6
timestamp 1731220651
transform 1 0 2024 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5910_6
timestamp 1731220651
transform 1 0 2112 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5909_6
timestamp 1731220651
transform 1 0 1704 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5908_6
timestamp 1731220651
transform 1 0 1768 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5907_6
timestamp 1731220651
transform 1 0 1824 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5906_6
timestamp 1731220651
transform 1 0 1880 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5905_6
timestamp 1731220651
transform 1 0 1928 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5904_6
timestamp 1731220651
transform 1 0 1968 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5903_6
timestamp 1731220651
transform 1 0 2008 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5902_6
timestamp 1731220651
transform 1 0 2048 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5901_6
timestamp 1731220651
transform 1 0 2088 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5900_6
timestamp 1731220651
transform 1 0 2136 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5899_6
timestamp 1731220651
transform 1 0 2184 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5898_6
timestamp 1731220651
transform 1 0 2200 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5897_6
timestamp 1731220651
transform 1 0 2232 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5896_6
timestamp 1731220651
transform 1 0 2272 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5895_6
timestamp 1731220651
transform 1 0 2312 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5894_6
timestamp 1731220651
transform 1 0 2352 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5893_6
timestamp 1731220651
transform 1 0 2352 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5892_6
timestamp 1731220651
transform 1 0 2288 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5891_6
timestamp 1731220651
transform 1 0 2352 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5890_6
timestamp 1731220651
transform 1 0 2272 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5889_6
timestamp 1731220651
transform 1 0 2192 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5888_6
timestamp 1731220651
transform 1 0 2240 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5887_6
timestamp 1731220651
transform 1 0 2152 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5886_6
timestamp 1731220651
transform 1 0 2072 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5885_6
timestamp 1731220651
transform 1 0 1912 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5884_6
timestamp 1731220651
transform 1 0 1992 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5883_6
timestamp 1731220651
transform 1 0 2016 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5882_6
timestamp 1731220651
transform 1 0 2096 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5881_6
timestamp 1731220651
transform 1 0 2088 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5880_6
timestamp 1731220651
transform 1 0 2024 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5879_6
timestamp 1731220651
transform 1 0 1960 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5878_6
timestamp 1731220651
transform 1 0 1944 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5877_6
timestamp 1731220651
transform 1 0 2040 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5876_6
timestamp 1731220651
transform 1 0 2144 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5875_6
timestamp 1731220651
transform 1 0 2024 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5874_6
timestamp 1731220651
transform 1 0 1936 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5873_6
timestamp 1731220651
transform 1 0 1848 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5872_6
timestamp 1731220651
transform 1 0 1768 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5871_6
timestamp 1731220651
transform 1 0 1752 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5870_6
timestamp 1731220651
transform 1 0 1816 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5869_6
timestamp 1731220651
transform 1 0 1880 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5868_6
timestamp 1731220651
transform 1 0 1944 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5867_6
timestamp 1731220651
transform 1 0 2016 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5866_6
timestamp 1731220651
transform 1 0 1816 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5865_6
timestamp 1731220651
transform 1 0 1888 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5864_6
timestamp 1731220651
transform 1 0 1952 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5863_6
timestamp 1731220651
transform 1 0 2016 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5862_6
timestamp 1731220651
transform 1 0 2080 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5861_6
timestamp 1731220651
transform 1 0 2136 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5860_6
timestamp 1731220651
transform 1 0 2184 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5859_6
timestamp 1731220651
transform 1 0 2272 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5858_6
timestamp 1731220651
transform 1 0 2096 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5857_6
timestamp 1731220651
transform 1 0 2112 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5856_6
timestamp 1731220651
transform 1 0 2200 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5855_6
timestamp 1731220651
transform 1 0 2256 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5854_6
timestamp 1731220651
transform 1 0 2160 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5853_6
timestamp 1731220651
transform 1 0 2232 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5852_6
timestamp 1731220651
transform 1 0 2280 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5851_6
timestamp 1731220651
transform 1 0 2184 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5850_6
timestamp 1731220651
transform 1 0 2064 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5849_6
timestamp 1731220651
transform 1 0 2128 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5848_6
timestamp 1731220651
transform 1 0 2192 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5847_6
timestamp 1731220651
transform 1 0 2248 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5846_6
timestamp 1731220651
transform 1 0 2328 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5845_6
timestamp 1731220651
transform 1 0 2312 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5844_6
timestamp 1731220651
transform 1 0 2352 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5843_6
timestamp 1731220651
transform 1 0 2352 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5842_6
timestamp 1731220651
transform 1 0 2304 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5841_6
timestamp 1731220651
transform 1 0 2352 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5840_6
timestamp 1731220651
transform 1 0 2352 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5839_6
timestamp 1731220651
transform 1 0 2352 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5838_6
timestamp 1731220651
transform 1 0 2288 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5837_6
timestamp 1731220651
transform 1 0 2352 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5836_6
timestamp 1731220651
transform 1 0 2192 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5835_6
timestamp 1731220651
transform 1 0 2248 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5834_6
timestamp 1731220651
transform 1 0 2312 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5833_6
timestamp 1731220651
transform 1 0 2352 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5832_6
timestamp 1731220651
transform 1 0 2352 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5831_6
timestamp 1731220651
transform 1 0 2304 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5830_6
timestamp 1731220651
transform 1 0 2232 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5829_6
timestamp 1731220651
transform 1 0 2168 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5828_6
timestamp 1731220651
transform 1 0 1928 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5827_6
timestamp 1731220651
transform 1 0 2016 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5826_6
timestamp 1731220651
transform 1 0 2096 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5825_6
timestamp 1731220651
transform 1 0 2136 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5824_6
timestamp 1731220651
transform 1 0 2200 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5823_6
timestamp 1731220651
transform 1 0 2272 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5822_6
timestamp 1731220651
transform 1 0 2064 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5821_6
timestamp 1731220651
transform 1 0 1824 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5820_6
timestamp 1731220651
transform 1 0 1912 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5819_6
timestamp 1731220651
transform 1 0 1992 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5818_6
timestamp 1731220651
transform 1 0 2016 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5817_6
timestamp 1731220651
transform 1 0 2072 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5816_6
timestamp 1731220651
transform 1 0 2128 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5815_6
timestamp 1731220651
transform 1 0 1960 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5814_6
timestamp 1731220651
transform 1 0 1784 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5813_6
timestamp 1731220651
transform 1 0 1848 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5812_6
timestamp 1731220651
transform 1 0 1904 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5811_6
timestamp 1731220651
transform 1 0 2016 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5810_6
timestamp 1731220651
transform 1 0 2128 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5809_6
timestamp 1731220651
transform 1 0 2248 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5808_6
timestamp 1731220651
transform 1 0 1920 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5807_6
timestamp 1731220651
transform 1 0 1848 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5806_6
timestamp 1731220651
transform 1 0 1792 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5805_6
timestamp 1731220651
transform 1 0 1752 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5804_6
timestamp 1731220651
transform 1 0 1784 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5803_6
timestamp 1731220651
transform 1 0 1832 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5802_6
timestamp 1731220651
transform 1 0 1896 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5801_6
timestamp 1731220651
transform 1 0 1960 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5800_6
timestamp 1731220651
transform 1 0 2032 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5799_6
timestamp 1731220651
transform 1 0 2112 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5798_6
timestamp 1731220651
transform 1 0 1768 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5797_6
timestamp 1731220651
transform 1 0 1824 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5796_6
timestamp 1731220651
transform 1 0 1896 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5795_6
timestamp 1731220651
transform 1 0 1976 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5794_6
timestamp 1731220651
transform 1 0 2064 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5793_6
timestamp 1731220651
transform 1 0 2160 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5792_6
timestamp 1731220651
transform 1 0 1808 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5791_6
timestamp 1731220651
transform 1 0 1896 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5790_6
timestamp 1731220651
transform 1 0 1984 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5789_6
timestamp 1731220651
transform 1 0 2064 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5788_6
timestamp 1731220651
transform 1 0 1776 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5787_6
timestamp 1731220651
transform 1 0 1864 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5786_6
timestamp 1731220651
transform 1 0 1944 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5785_6
timestamp 1731220651
transform 1 0 2024 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5784_6
timestamp 1731220651
transform 1 0 2096 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5783_6
timestamp 1731220651
transform 1 0 2160 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5782_6
timestamp 1731220651
transform 1 0 2232 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5781_6
timestamp 1731220651
transform 1 0 2304 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5780_6
timestamp 1731220651
transform 1 0 2144 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5779_6
timestamp 1731220651
transform 1 0 2216 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5778_6
timestamp 1731220651
transform 1 0 2264 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5777_6
timestamp 1731220651
transform 1 0 2200 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5776_6
timestamp 1731220651
transform 1 0 2184 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5775_6
timestamp 1731220651
transform 1 0 2248 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5774_6
timestamp 1731220651
transform 1 0 2312 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5773_6
timestamp 1731220651
transform 1 0 2352 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5772_6
timestamp 1731220651
transform 1 0 2352 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5771_6
timestamp 1731220651
transform 1 0 2288 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5770_6
timestamp 1731220651
transform 1 0 2352 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5769_6
timestamp 1731220651
transform 1 0 2352 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5768_6
timestamp 1731220651
transform 1 0 2352 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5767_6
timestamp 1731220651
transform 1 0 2296 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5766_6
timestamp 1731220651
transform 1 0 2352 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5765_6
timestamp 1731220651
transform 1 0 2352 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5764_6
timestamp 1731220651
transform 1 0 2312 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5763_6
timestamp 1731220651
transform 1 0 2352 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5762_6
timestamp 1731220651
transform 1 0 2312 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5761_6
timestamp 1731220651
transform 1 0 2248 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5760_6
timestamp 1731220651
transform 1 0 2248 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5759_6
timestamp 1731220651
transform 1 0 2184 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5758_6
timestamp 1731220651
transform 1 0 2120 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5757_6
timestamp 1731220651
transform 1 0 2048 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5756_6
timestamp 1731220651
transform 1 0 1752 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5755_6
timestamp 1731220651
transform 1 0 1864 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5754_6
timestamp 1731220651
transform 1 0 1960 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5753_6
timestamp 1731220651
transform 1 0 2056 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5752_6
timestamp 1731220651
transform 1 0 2120 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5751_6
timestamp 1731220651
transform 1 0 2184 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5750_6
timestamp 1731220651
transform 1 0 1992 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5749_6
timestamp 1731220651
transform 1 0 1848 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5748_6
timestamp 1731220651
transform 1 0 1920 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5747_6
timestamp 1731220651
transform 1 0 1968 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5746_6
timestamp 1731220651
transform 1 0 2024 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5745_6
timestamp 1731220651
transform 1 0 2080 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5744_6
timestamp 1731220651
transform 1 0 1912 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5743_6
timestamp 1731220651
transform 1 0 1744 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5742_6
timestamp 1731220651
transform 1 0 1800 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5741_6
timestamp 1731220651
transform 1 0 1856 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5740_6
timestamp 1731220651
transform 1 0 1912 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5739_6
timestamp 1731220651
transform 1 0 1968 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5738_6
timestamp 1731220651
transform 1 0 1800 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5737_6
timestamp 1731220651
transform 1 0 1640 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5736_6
timestamp 1731220651
transform 1 0 1696 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5735_6
timestamp 1731220651
transform 1 0 1752 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5734_6
timestamp 1731220651
transform 1 0 1856 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5733_6
timestamp 1731220651
transform 1 0 1888 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5732_6
timestamp 1731220651
transform 1 0 1944 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5731_6
timestamp 1731220651
transform 1 0 1832 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5730_6
timestamp 1731220651
transform 1 0 1776 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5729_6
timestamp 1731220651
transform 1 0 1720 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5728_6
timestamp 1731220651
transform 1 0 1664 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5727_6
timestamp 1731220651
transform 1 0 1704 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5726_6
timestamp 1731220651
transform 1 0 1800 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5725_6
timestamp 1731220651
transform 1 0 1912 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5724_6
timestamp 1731220651
transform 1 0 2024 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5723_6
timestamp 1731220651
transform 1 0 1864 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5722_6
timestamp 1731220651
transform 1 0 1816 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5721_6
timestamp 1731220651
transform 1 0 1760 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5720_6
timestamp 1731220651
transform 1 0 1712 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5719_6
timestamp 1731220651
transform 1 0 1672 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5718_6
timestamp 1731220651
transform 1 0 1632 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5717_6
timestamp 1731220651
transform 1 0 1592 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5716_6
timestamp 1731220651
transform 1 0 1552 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5715_6
timestamp 1731220651
transform 1 0 1512 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5714_6
timestamp 1731220651
transform 1 0 1392 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5713_6
timestamp 1731220651
transform 1 0 1432 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5712_6
timestamp 1731220651
transform 1 0 1472 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5711_6
timestamp 1731220651
transform 1 0 1504 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5710_6
timestamp 1731220651
transform 1 0 1560 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5709_6
timestamp 1731220651
transform 1 0 1624 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5708_6
timestamp 1731220651
transform 1 0 1456 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5707_6
timestamp 1731220651
transform 1 0 1416 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5706_6
timestamp 1731220651
transform 1 0 1376 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5705_6
timestamp 1731220651
transform 1 0 1336 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5704_6
timestamp 1731220651
transform 1 0 1352 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5703_6
timestamp 1731220651
transform 1 0 1392 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5702_6
timestamp 1731220651
transform 1 0 1440 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5701_6
timestamp 1731220651
transform 1 0 1496 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5700_6
timestamp 1731220651
transform 1 0 1552 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5699_6
timestamp 1731220651
transform 1 0 1608 0 -1 1852
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5698_6
timestamp 1731220651
transform 1 0 1384 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5697_6
timestamp 1731220651
transform 1 0 1448 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5696_6
timestamp 1731220651
transform 1 0 1512 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5695_6
timestamp 1731220651
transform 1 0 1576 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5694_6
timestamp 1731220651
transform 1 0 1496 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5693_6
timestamp 1731220651
transform 1 0 1552 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5692_6
timestamp 1731220651
transform 1 0 1616 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5691_6
timestamp 1731220651
transform 1 0 1680 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5690_6
timestamp 1731220651
transform 1 0 1552 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5689_6
timestamp 1731220651
transform 1 0 1624 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5688_6
timestamp 1731220651
transform 1 0 1696 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5687_6
timestamp 1731220651
transform 1 0 1776 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5686_6
timestamp 1731220651
transform 1 0 1616 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5685_6
timestamp 1731220651
transform 1 0 1464 0 -1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5684_6
timestamp 1731220651
transform 1 0 1496 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5683_6
timestamp 1731220651
transform 1 0 1456 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5682_6
timestamp 1731220651
transform 1 0 1416 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5681_6
timestamp 1731220651
transform 1 0 1296 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5680_6
timestamp 1731220651
transform 1 0 1336 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5679_6
timestamp 1731220651
transform 1 0 1376 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5678_6
timestamp 1731220651
transform 1 0 1416 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5677_6
timestamp 1731220651
transform 1 0 1456 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5676_6
timestamp 1731220651
transform 1 0 1376 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5675_6
timestamp 1731220651
transform 1 0 1296 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5674_6
timestamp 1731220651
transform 1 0 1336 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5673_6
timestamp 1731220651
transform 1 0 1336 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5672_6
timestamp 1731220651
transform 1 0 1296 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5671_6
timestamp 1731220651
transform 1 0 1184 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5670_6
timestamp 1731220651
transform 1 0 992 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5669_6
timestamp 1731220651
transform 1 0 1064 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5668_6
timestamp 1731220651
transform 1 0 1136 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5667_6
timestamp 1731220651
transform 1 0 1184 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5666_6
timestamp 1731220651
transform 1 0 1120 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5665_6
timestamp 1731220651
transform 1 0 968 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5664_6
timestamp 1731220651
transform 1 0 1040 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5663_6
timestamp 1731220651
transform 1 0 1048 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5662_6
timestamp 1731220651
transform 1 0 1120 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5661_6
timestamp 1731220651
transform 1 0 912 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5660_6
timestamp 1731220651
transform 1 0 976 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5659_6
timestamp 1731220651
transform 1 0 1000 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5658_6
timestamp 1731220651
transform 1 0 928 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5657_6
timestamp 1731220651
transform 1 0 856 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5656_6
timestamp 1731220651
transform 1 0 784 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5655_6
timestamp 1731220651
transform 1 0 808 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5654_6
timestamp 1731220651
transform 1 0 736 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5653_6
timestamp 1731220651
transform 1 0 544 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5652_6
timestamp 1731220651
transform 1 0 480 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5651_6
timestamp 1731220651
transform 1 0 472 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5650_6
timestamp 1731220651
transform 1 0 336 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5649_6
timestamp 1731220651
transform 1 0 408 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5648_6
timestamp 1731220651
transform 1 0 432 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5647_6
timestamp 1731220651
transform 1 0 272 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5646_6
timestamp 1731220651
transform 1 0 352 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5645_6
timestamp 1731220651
transform 1 0 400 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5644_6
timestamp 1731220651
transform 1 0 328 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5643_6
timestamp 1731220651
transform 1 0 272 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5642_6
timestamp 1731220651
transform 1 0 216 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5641_6
timestamp 1731220651
transform 1 0 176 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5640_6
timestamp 1731220651
transform 1 0 136 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5639_6
timestamp 1731220651
transform 1 0 128 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5638_6
timestamp 1731220651
transform 1 0 200 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5637_6
timestamp 1731220651
transform 1 0 264 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5636_6
timestamp 1731220651
transform 1 0 184 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5635_6
timestamp 1731220651
transform 1 0 128 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5634_6
timestamp 1731220651
transform 1 0 128 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5633_6
timestamp 1731220651
transform 1 0 168 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5632_6
timestamp 1731220651
transform 1 0 208 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5631_6
timestamp 1731220651
transform 1 0 272 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5630_6
timestamp 1731220651
transform 1 0 344 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5629_6
timestamp 1731220651
transform 1 0 416 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5628_6
timestamp 1731220651
transform 1 0 128 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5627_6
timestamp 1731220651
transform 1 0 168 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5626_6
timestamp 1731220651
transform 1 0 208 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5625_6
timestamp 1731220651
transform 1 0 264 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5624_6
timestamp 1731220651
transform 1 0 336 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5623_6
timestamp 1731220651
transform 1 0 408 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5622_6
timestamp 1731220651
transform 1 0 488 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5621_6
timestamp 1731220651
transform 1 0 240 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5620_6
timestamp 1731220651
transform 1 0 280 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5619_6
timestamp 1731220651
transform 1 0 320 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5618_6
timestamp 1731220651
transform 1 0 360 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5617_6
timestamp 1731220651
transform 1 0 408 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5616_6
timestamp 1731220651
transform 1 0 464 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5615_6
timestamp 1731220651
transform 1 0 528 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5614_6
timestamp 1731220651
transform 1 0 592 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5613_6
timestamp 1731220651
transform 1 0 392 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5612_6
timestamp 1731220651
transform 1 0 432 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5611_6
timestamp 1731220651
transform 1 0 472 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5610_6
timestamp 1731220651
transform 1 0 512 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5609_6
timestamp 1731220651
transform 1 0 560 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5608_6
timestamp 1731220651
transform 1 0 616 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5607_6
timestamp 1731220651
transform 1 0 680 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5606_6
timestamp 1731220651
transform 1 0 640 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5605_6
timestamp 1731220651
transform 1 0 600 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5604_6
timestamp 1731220651
transform 1 0 560 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5603_6
timestamp 1731220651
transform 1 0 520 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5602_6
timestamp 1731220651
transform 1 0 480 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5601_6
timestamp 1731220651
transform 1 0 440 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5600_6
timestamp 1731220651
transform 1 0 400 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5599_6
timestamp 1731220651
transform 1 0 440 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5598_6
timestamp 1731220651
transform 1 0 488 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5597_6
timestamp 1731220651
transform 1 0 536 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5596_6
timestamp 1731220651
transform 1 0 392 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5595_6
timestamp 1731220651
transform 1 0 272 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5594_6
timestamp 1731220651
transform 1 0 312 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5593_6
timestamp 1731220651
transform 1 0 352 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5592_6
timestamp 1731220651
transform 1 0 384 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5591_6
timestamp 1731220651
transform 1 0 464 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5590_6
timestamp 1731220651
transform 1 0 552 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5589_6
timestamp 1731220651
transform 1 0 304 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5588_6
timestamp 1731220651
transform 1 0 248 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5587_6
timestamp 1731220651
transform 1 0 208 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5586_6
timestamp 1731220651
transform 1 0 128 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5585_6
timestamp 1731220651
transform 1 0 168 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5584_6
timestamp 1731220651
transform 1 0 144 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5583_6
timestamp 1731220651
transform 1 0 192 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5582_6
timestamp 1731220651
transform 1 0 256 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5581_6
timestamp 1731220651
transform 1 0 336 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5580_6
timestamp 1731220651
transform 1 0 432 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5579_6
timestamp 1731220651
transform 1 0 528 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5578_6
timestamp 1731220651
transform 1 0 632 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5577_6
timestamp 1731220651
transform 1 0 312 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5576_6
timestamp 1731220651
transform 1 0 352 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5575_6
timestamp 1731220651
transform 1 0 392 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5574_6
timestamp 1731220651
transform 1 0 440 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5573_6
timestamp 1731220651
transform 1 0 496 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5572_6
timestamp 1731220651
transform 1 0 552 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5571_6
timestamp 1731220651
transform 1 0 608 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5570_6
timestamp 1731220651
transform 1 0 552 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5569_6
timestamp 1731220651
transform 1 0 496 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5568_6
timestamp 1731220651
transform 1 0 440 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5567_6
timestamp 1731220651
transform 1 0 384 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5566_6
timestamp 1731220651
transform 1 0 336 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5565_6
timestamp 1731220651
transform 1 0 256 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5564_6
timestamp 1731220651
transform 1 0 296 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5563_6
timestamp 1731220651
transform 1 0 320 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5562_6
timestamp 1731220651
transform 1 0 400 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5561_6
timestamp 1731220651
transform 1 0 488 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5560_6
timestamp 1731220651
transform 1 0 248 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5559_6
timestamp 1731220651
transform 1 0 128 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5558_6
timestamp 1731220651
transform 1 0 168 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5557_6
timestamp 1731220651
transform 1 0 208 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5556_6
timestamp 1731220651
transform 1 0 240 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5555_6
timestamp 1731220651
transform 1 0 320 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5554_6
timestamp 1731220651
transform 1 0 408 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5553_6
timestamp 1731220651
transform 1 0 168 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5552_6
timestamp 1731220651
transform 1 0 128 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5551_6
timestamp 1731220651
transform 1 0 128 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5550_6
timestamp 1731220651
transform 1 0 168 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5549_6
timestamp 1731220651
transform 1 0 224 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5548_6
timestamp 1731220651
transform 1 0 296 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5547_6
timestamp 1731220651
transform 1 0 376 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5546_6
timestamp 1731220651
transform 1 0 128 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5545_6
timestamp 1731220651
transform 1 0 208 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5544_6
timestamp 1731220651
transform 1 0 296 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5543_6
timestamp 1731220651
transform 1 0 384 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5542_6
timestamp 1731220651
transform 1 0 192 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5541_6
timestamp 1731220651
transform 1 0 232 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5540_6
timestamp 1731220651
transform 1 0 280 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5539_6
timestamp 1731220651
transform 1 0 336 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5538_6
timestamp 1731220651
transform 1 0 384 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5537_6
timestamp 1731220651
transform 1 0 288 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5536_6
timestamp 1731220651
transform 1 0 336 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5535_6
timestamp 1731220651
transform 1 0 392 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5534_6
timestamp 1731220651
transform 1 0 464 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5533_6
timestamp 1731220651
transform 1 0 528 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5532_6
timestamp 1731220651
transform 1 0 448 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5531_6
timestamp 1731220651
transform 1 0 368 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5530_6
timestamp 1731220651
transform 1 0 248 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5529_6
timestamp 1731220651
transform 1 0 304 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5528_6
timestamp 1731220651
transform 1 0 304 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5527_6
timestamp 1731220651
transform 1 0 376 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5526_6
timestamp 1731220651
transform 1 0 184 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5525_6
timestamp 1731220651
transform 1 0 240 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5524_6
timestamp 1731220651
transform 1 0 272 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5523_6
timestamp 1731220651
transform 1 0 344 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5522_6
timestamp 1731220651
transform 1 0 208 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5521_6
timestamp 1731220651
transform 1 0 128 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5520_6
timestamp 1731220651
transform 1 0 168 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5519_6
timestamp 1731220651
transform 1 0 168 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5518_6
timestamp 1731220651
transform 1 0 224 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5517_6
timestamp 1731220651
transform 1 0 280 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5516_6
timestamp 1731220651
transform 1 0 128 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5515_6
timestamp 1731220651
transform 1 0 128 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5514_6
timestamp 1731220651
transform 1 0 176 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5513_6
timestamp 1731220651
transform 1 0 248 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5512_6
timestamp 1731220651
transform 1 0 320 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5511_6
timestamp 1731220651
transform 1 0 280 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5510_6
timestamp 1731220651
transform 1 0 144 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5509_6
timestamp 1731220651
transform 1 0 216 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5508_6
timestamp 1731220651
transform 1 0 232 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5507_6
timestamp 1731220651
transform 1 0 272 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5506_6
timestamp 1731220651
transform 1 0 320 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5505_6
timestamp 1731220651
transform 1 0 376 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5504_6
timestamp 1731220651
transform 1 0 264 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5503_6
timestamp 1731220651
transform 1 0 216 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5502_6
timestamp 1731220651
transform 1 0 176 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5501_6
timestamp 1731220651
transform 1 0 136 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5500_6
timestamp 1731220651
transform 1 0 168 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5499_6
timestamp 1731220651
transform 1 0 208 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5498_6
timestamp 1731220651
transform 1 0 248 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5497_6
timestamp 1731220651
transform 1 0 128 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5496_6
timestamp 1731220651
transform 1 0 128 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5495_6
timestamp 1731220651
transform 1 0 288 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5494_6
timestamp 1731220651
transform 1 0 328 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5493_6
timestamp 1731220651
transform 1 0 384 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5492_6
timestamp 1731220651
transform 1 0 440 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5491_6
timestamp 1731220651
transform 1 0 328 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5490_6
timestamp 1731220651
transform 1 0 392 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5489_6
timestamp 1731220651
transform 1 0 464 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5488_6
timestamp 1731220651
transform 1 0 536 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5487_6
timestamp 1731220651
transform 1 0 560 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5486_6
timestamp 1731220651
transform 1 0 496 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5485_6
timestamp 1731220651
transform 1 0 432 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5484_6
timestamp 1731220651
transform 1 0 344 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5483_6
timestamp 1731220651
transform 1 0 408 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5482_6
timestamp 1731220651
transform 1 0 472 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5481_6
timestamp 1731220651
transform 1 0 544 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5480_6
timestamp 1731220651
transform 1 0 552 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5479_6
timestamp 1731220651
transform 1 0 392 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5478_6
timestamp 1731220651
transform 1 0 472 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5477_6
timestamp 1731220651
transform 1 0 496 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5476_6
timestamp 1731220651
transform 1 0 448 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5475_6
timestamp 1731220651
transform 1 0 336 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5474_6
timestamp 1731220651
transform 1 0 392 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5473_6
timestamp 1731220651
transform 1 0 416 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5472_6
timestamp 1731220651
transform 1 0 488 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5471_6
timestamp 1731220651
transform 1 0 456 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5470_6
timestamp 1731220651
transform 1 0 536 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5469_6
timestamp 1731220651
transform 1 0 608 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5468_6
timestamp 1731220651
transform 1 0 616 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5467_6
timestamp 1731220651
transform 1 0 704 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5466_6
timestamp 1731220651
transform 1 0 720 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5465_6
timestamp 1731220651
transform 1 0 632 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5464_6
timestamp 1731220651
transform 1 0 544 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5463_6
timestamp 1731220651
transform 1 0 432 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5462_6
timestamp 1731220651
transform 1 0 480 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5461_6
timestamp 1731220651
transform 1 0 528 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5460_6
timestamp 1731220651
transform 1 0 552 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5459_6
timestamp 1731220651
transform 1 0 472 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5458_6
timestamp 1731220651
transform 1 0 464 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5457_6
timestamp 1731220651
transform 1 0 552 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5456_6
timestamp 1731220651
transform 1 0 632 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5455_6
timestamp 1731220651
transform 1 0 664 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5454_6
timestamp 1731220651
transform 1 0 584 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5453_6
timestamp 1731220651
transform 1 0 496 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5452_6
timestamp 1731220651
transform 1 0 576 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5451_6
timestamp 1731220651
transform 1 0 664 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5450_6
timestamp 1731220651
transform 1 0 752 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5449_6
timestamp 1731220651
transform 1 0 616 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5448_6
timestamp 1731220651
transform 1 0 680 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5447_6
timestamp 1731220651
transform 1 0 744 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5446_6
timestamp 1731220651
transform 1 0 808 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5445_6
timestamp 1731220651
transform 1 0 664 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5444_6
timestamp 1731220651
transform 1 0 728 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5443_6
timestamp 1731220651
transform 1 0 792 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5442_6
timestamp 1731220651
transform 1 0 848 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5441_6
timestamp 1731220651
transform 1 0 904 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5440_6
timestamp 1731220651
transform 1 0 960 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5439_6
timestamp 1731220651
transform 1 0 1016 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5438_6
timestamp 1731220651
transform 1 0 944 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5437_6
timestamp 1731220651
transform 1 0 872 0 -1 1412
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5436_6
timestamp 1731220651
transform 1 0 832 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5435_6
timestamp 1731220651
transform 1 0 912 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5434_6
timestamp 1731220651
transform 1 0 1000 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5433_6
timestamp 1731220651
transform 1 0 1088 0 1 1272
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5432_6
timestamp 1731220651
transform 1 0 1064 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5431_6
timestamp 1731220651
transform 1 0 1000 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5430_6
timestamp 1731220651
transform 1 0 936 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5429_6
timestamp 1731220651
transform 1 0 872 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5428_6
timestamp 1731220651
transform 1 0 736 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5427_6
timestamp 1731220651
transform 1 0 808 0 -1 1268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5426_6
timestamp 1731220651
transform 1 0 864 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5425_6
timestamp 1731220651
transform 1 0 792 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5424_6
timestamp 1731220651
transform 1 0 712 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5423_6
timestamp 1731220651
transform 1 0 704 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5422_6
timestamp 1731220651
transform 1 0 632 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5421_6
timestamp 1731220651
transform 1 0 576 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5420_6
timestamp 1731220651
transform 1 0 624 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5419_6
timestamp 1731220651
transform 1 0 672 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5418_6
timestamp 1731220651
transform 1 0 720 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5417_6
timestamp 1731220651
transform 1 0 776 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5416_6
timestamp 1731220651
transform 1 0 832 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5415_6
timestamp 1731220651
transform 1 0 888 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5414_6
timestamp 1731220651
transform 1 0 952 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5413_6
timestamp 1731220651
transform 1 0 768 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5412_6
timestamp 1731220651
transform 1 0 832 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5411_6
timestamp 1731220651
transform 1 0 896 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5410_6
timestamp 1731220651
transform 1 0 952 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5409_6
timestamp 1731220651
transform 1 0 1016 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5408_6
timestamp 1731220651
transform 1 0 928 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5407_6
timestamp 1731220651
transform 1 0 984 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5406_6
timestamp 1731220651
transform 1 0 1040 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5405_6
timestamp 1731220651
transform 1 0 1096 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5404_6
timestamp 1731220651
transform 1 0 1144 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5403_6
timestamp 1731220651
transform 1 0 1184 0 1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5402_6
timestamp 1731220651
transform 1 0 1080 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5401_6
timestamp 1731220651
transform 1 0 1144 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5400_6
timestamp 1731220651
transform 1 0 1184 0 -1 1124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5399_6
timestamp 1731220651
transform 1 0 1184 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5398_6
timestamp 1731220651
transform 1 0 1144 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5397_6
timestamp 1731220651
transform 1 0 1016 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5396_6
timestamp 1731220651
transform 1 0 1080 0 1 984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5395_6
timestamp 1731220651
transform 1 0 1080 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5394_6
timestamp 1731220651
transform 1 0 1144 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5393_6
timestamp 1731220651
transform 1 0 1184 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5392_6
timestamp 1731220651
transform 1 0 800 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5391_6
timestamp 1731220651
transform 1 0 880 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5390_6
timestamp 1731220651
transform 1 0 952 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5389_6
timestamp 1731220651
transform 1 0 1016 0 -1 972
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5388_6
timestamp 1731220651
transform 1 0 1048 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5387_6
timestamp 1731220651
transform 1 0 1112 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5386_6
timestamp 1731220651
transform 1 0 1176 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5385_6
timestamp 1731220651
transform 1 0 992 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5384_6
timestamp 1731220651
transform 1 0 928 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5383_6
timestamp 1731220651
transform 1 0 784 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5382_6
timestamp 1731220651
transform 1 0 856 0 1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5381_6
timestamp 1731220651
transform 1 0 920 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5380_6
timestamp 1731220651
transform 1 0 976 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5379_6
timestamp 1731220651
transform 1 0 1040 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5378_6
timestamp 1731220651
transform 1 0 864 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5377_6
timestamp 1731220651
transform 1 0 680 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5376_6
timestamp 1731220651
transform 1 0 744 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5375_6
timestamp 1731220651
transform 1 0 808 0 -1 828
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5374_6
timestamp 1731220651
transform 1 0 872 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5373_6
timestamp 1731220651
transform 1 0 976 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5372_6
timestamp 1731220651
transform 1 0 1088 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5371_6
timestamp 1731220651
transform 1 0 776 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5370_6
timestamp 1731220651
transform 1 0 552 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5369_6
timestamp 1731220651
transform 1 0 616 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5368_6
timestamp 1731220651
transform 1 0 688 0 1 692
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5367_6
timestamp 1731220651
transform 1 0 760 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5366_6
timestamp 1731220651
transform 1 0 832 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5365_6
timestamp 1731220651
transform 1 0 688 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5364_6
timestamp 1731220651
transform 1 0 552 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5363_6
timestamp 1731220651
transform 1 0 616 0 -1 684
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5362_6
timestamp 1731220651
transform 1 0 632 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5361_6
timestamp 1731220651
transform 1 0 712 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5360_6
timestamp 1731220651
transform 1 0 792 0 1 548
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5359_6
timestamp 1731220651
transform 1 0 616 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5358_6
timestamp 1731220651
transform 1 0 688 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5357_6
timestamp 1731220651
transform 1 0 760 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5356_6
timestamp 1731220651
transform 1 0 832 0 -1 544
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5355_6
timestamp 1731220651
transform 1 0 624 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5354_6
timestamp 1731220651
transform 1 0 688 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5353_6
timestamp 1731220651
transform 1 0 752 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5352_6
timestamp 1731220651
transform 1 0 816 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5351_6
timestamp 1731220651
transform 1 0 880 0 1 408
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5350_6
timestamp 1731220651
transform 1 0 856 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5349_6
timestamp 1731220651
transform 1 0 800 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5348_6
timestamp 1731220651
transform 1 0 744 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5347_6
timestamp 1731220651
transform 1 0 680 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5346_6
timestamp 1731220651
transform 1 0 608 0 -1 404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5345_6
timestamp 1731220651
transform 1 0 584 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5344_6
timestamp 1731220651
transform 1 0 632 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5343_6
timestamp 1731220651
transform 1 0 680 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5342_6
timestamp 1731220651
transform 1 0 728 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5341_6
timestamp 1731220651
transform 1 0 776 0 1 260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5340_6
timestamp 1731220651
transform 1 0 688 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5339_6
timestamp 1731220651
transform 1 0 728 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5338_6
timestamp 1731220651
transform 1 0 776 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5337_6
timestamp 1731220651
transform 1 0 824 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5336_6
timestamp 1731220651
transform 1 0 872 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5335_6
timestamp 1731220651
transform 1 0 920 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5334_6
timestamp 1731220651
transform 1 0 968 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5333_6
timestamp 1731220651
transform 1 0 1016 0 -1 252
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5332_6
timestamp 1731220651
transform 1 0 624 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5331_6
timestamp 1731220651
transform 1 0 664 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5330_6
timestamp 1731220651
transform 1 0 704 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5329_6
timestamp 1731220651
transform 1 0 744 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5328_6
timestamp 1731220651
transform 1 0 784 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5327_6
timestamp 1731220651
transform 1 0 824 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5326_6
timestamp 1731220651
transform 1 0 864 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5325_6
timestamp 1731220651
transform 1 0 904 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5324_6
timestamp 1731220651
transform 1 0 944 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5323_6
timestamp 1731220651
transform 1 0 984 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5322_6
timestamp 1731220651
transform 1 0 1024 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5321_6
timestamp 1731220651
transform 1 0 1064 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5320_6
timestamp 1731220651
transform 1 0 1104 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5319_6
timestamp 1731220651
transform 1 0 1144 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5318_6
timestamp 1731220651
transform 1 0 1184 0 1 84
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5317_6
timestamp 1731220651
transform 1 0 1296 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5316_6
timestamp 1731220651
transform 1 0 1336 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5315_6
timestamp 1731220651
transform 1 0 1376 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5314_6
timestamp 1731220651
transform 1 0 1416 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5313_6
timestamp 1731220651
transform 1 0 1456 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5312_6
timestamp 1731220651
transform 1 0 1512 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5311_6
timestamp 1731220651
transform 1 0 1576 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5310_6
timestamp 1731220651
transform 1 0 1640 0 1 100
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5309_6
timestamp 1731220651
transform 1 0 1360 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5308_6
timestamp 1731220651
transform 1 0 1400 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5307_6
timestamp 1731220651
transform 1 0 1448 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5306_6
timestamp 1731220651
transform 1 0 1504 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5305_6
timestamp 1731220651
transform 1 0 1560 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5304_6
timestamp 1731220651
transform 1 0 1624 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5303_6
timestamp 1731220651
transform 1 0 1696 0 -1 244
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5302_6
timestamp 1731220651
transform 1 0 1624 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5301_6
timestamp 1731220651
transform 1 0 1664 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5300_6
timestamp 1731220651
transform 1 0 1704 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5299_6
timestamp 1731220651
transform 1 0 1744 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5298_6
timestamp 1731220651
transform 1 0 1784 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5297_6
timestamp 1731220651
transform 1 0 1504 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5296_6
timestamp 1731220651
transform 1 0 1544 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5295_6
timestamp 1731220651
transform 1 0 1584 0 1 248
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5294_6
timestamp 1731220651
transform 1 0 1600 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5293_6
timestamp 1731220651
transform 1 0 1672 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5292_6
timestamp 1731220651
transform 1 0 1536 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5291_6
timestamp 1731220651
transform 1 0 1480 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5290_6
timestamp 1731220651
transform 1 0 1432 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5289_6
timestamp 1731220651
transform 1 0 1392 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5288_6
timestamp 1731220651
transform 1 0 1352 0 -1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5287_6
timestamp 1731220651
transform 1 0 1296 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5286_6
timestamp 1731220651
transform 1 0 1336 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5285_6
timestamp 1731220651
transform 1 0 1376 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5284_6
timestamp 1731220651
transform 1 0 1440 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5283_6
timestamp 1731220651
transform 1 0 1528 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5282_6
timestamp 1731220651
transform 1 0 1624 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5281_6
timestamp 1731220651
transform 1 0 1728 0 1 392
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5280_6
timestamp 1731220651
transform 1 0 1400 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5279_6
timestamp 1731220651
transform 1 0 1440 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5278_6
timestamp 1731220651
transform 1 0 1480 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5277_6
timestamp 1731220651
transform 1 0 1528 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5276_6
timestamp 1731220651
transform 1 0 1584 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5275_6
timestamp 1731220651
transform 1 0 1640 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5274_6
timestamp 1731220651
transform 1 0 1704 0 -1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5273_6
timestamp 1731220651
transform 1 0 1672 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5272_6
timestamp 1731220651
transform 1 0 1712 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5271_6
timestamp 1731220651
transform 1 0 1752 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5270_6
timestamp 1731220651
transform 1 0 1800 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5269_6
timestamp 1731220651
transform 1 0 1632 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5268_6
timestamp 1731220651
transform 1 0 1592 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5267_6
timestamp 1731220651
transform 1 0 1552 0 1 528
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5266_6
timestamp 1731220651
transform 1 0 1584 0 -1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5265_6
timestamp 1731220651
transform 1 0 1528 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5264_6
timestamp 1731220651
transform 1 0 1448 0 1 672
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5263_6
timestamp 1731220651
transform 1 0 1472 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5262_6
timestamp 1731220651
transform 1 0 1544 0 -1 808
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5261_6
timestamp 1731220651
transform 1 0 1528 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5260_6
timestamp 1731220651
transform 1 0 1464 0 1 812
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5259_6
timestamp 1731220651
transform 1 0 1456 0 -1 956
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5258_6
timestamp 1731220651
transform 1 0 1496 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5257_6
timestamp 1731220651
transform 1 0 1616 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5256_6
timestamp 1731220651
transform 1 0 1728 0 1 964
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5255_6
timestamp 1731220651
transform 1 0 1528 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5254_6
timestamp 1731220651
transform 1 0 1592 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5253_6
timestamp 1731220651
transform 1 0 1656 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5252_6
timestamp 1731220651
transform 1 0 1720 0 -1 1112
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5251_6
timestamp 1731220651
transform 1 0 1552 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5250_6
timestamp 1731220651
transform 1 0 1592 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5249_6
timestamp 1731220651
transform 1 0 1632 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5248_6
timestamp 1731220651
transform 1 0 1672 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5247_6
timestamp 1731220651
transform 1 0 1712 0 1 1120
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5246_6
timestamp 1731220651
transform 1 0 1744 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5245_6
timestamp 1731220651
transform 1 0 1704 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5244_6
timestamp 1731220651
transform 1 0 1664 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5243_6
timestamp 1731220651
transform 1 0 1624 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5242_6
timestamp 1731220651
transform 1 0 1504 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5241_6
timestamp 1731220651
transform 1 0 1544 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5240_6
timestamp 1731220651
transform 1 0 1584 0 -1 1260
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5239_6
timestamp 1731220651
transform 1 0 1608 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5238_6
timestamp 1731220651
transform 1 0 1664 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5237_6
timestamp 1731220651
transform 1 0 1712 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5236_6
timestamp 1731220651
transform 1 0 1560 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5235_6
timestamp 1731220651
transform 1 0 1440 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5234_6
timestamp 1731220651
transform 1 0 1480 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5233_6
timestamp 1731220651
transform 1 0 1520 0 1 1264
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5232_6
timestamp 1731220651
transform 1 0 1544 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5231_6
timestamp 1731220651
transform 1 0 1632 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5230_6
timestamp 1731220651
transform 1 0 1720 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5229_6
timestamp 1731220651
transform 1 0 1464 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5228_6
timestamp 1731220651
transform 1 0 1296 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5227_6
timestamp 1731220651
transform 1 0 1336 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5226_6
timestamp 1731220651
transform 1 0 1392 0 -1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5225_6
timestamp 1731220651
transform 1 0 1472 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5224_6
timestamp 1731220651
transform 1 0 1576 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5223_6
timestamp 1731220651
transform 1 0 1680 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5222_6
timestamp 1731220651
transform 1 0 1368 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5221_6
timestamp 1731220651
transform 1 0 1296 0 1 1404
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5220_6
timestamp 1731220651
transform 1 0 1184 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5219_6
timestamp 1731220651
transform 1 0 1016 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5218_6
timestamp 1731220651
transform 1 0 1080 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5217_6
timestamp 1731220651
transform 1 0 1144 0 1 1416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5216_6
timestamp 1731220651
transform 1 0 1184 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5215_6
timestamp 1731220651
transform 1 0 1112 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5214_6
timestamp 1731220651
transform 1 0 1040 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5213_6
timestamp 1731220651
transform 1 0 968 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5212_6
timestamp 1731220651
transform 1 0 728 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5211_6
timestamp 1731220651
transform 1 0 816 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5210_6
timestamp 1731220651
transform 1 0 896 0 -1 1556
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5209_6
timestamp 1731220651
transform 1 0 912 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5208_6
timestamp 1731220651
transform 1 0 976 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5207_6
timestamp 1731220651
transform 1 0 1040 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5206_6
timestamp 1731220651
transform 1 0 848 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5205_6
timestamp 1731220651
transform 1 0 632 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5204_6
timestamp 1731220651
transform 1 0 712 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5203_6
timestamp 1731220651
transform 1 0 784 0 1 1560
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5202_6
timestamp 1731220651
transform 1 0 832 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5201_6
timestamp 1731220651
transform 1 0 888 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5200_6
timestamp 1731220651
transform 1 0 776 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5199_6
timestamp 1731220651
transform 1 0 728 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5198_6
timestamp 1731220651
transform 1 0 680 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5197_6
timestamp 1731220651
transform 1 0 584 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5196_6
timestamp 1731220651
transform 1 0 632 0 -1 1700
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5195_6
timestamp 1731220651
transform 1 0 688 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5194_6
timestamp 1731220651
transform 1 0 744 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5193_6
timestamp 1731220651
transform 1 0 800 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5192_6
timestamp 1731220651
transform 1 0 864 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5191_6
timestamp 1731220651
transform 1 0 928 0 1 1704
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5190_6
timestamp 1731220651
transform 1 0 896 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5189_6
timestamp 1731220651
transform 1 0 752 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5188_6
timestamp 1731220651
transform 1 0 824 0 -1 1840
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5187_6
timestamp 1731220651
transform 1 0 848 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5186_6
timestamp 1731220651
transform 1 0 784 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5185_6
timestamp 1731220651
transform 1 0 720 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5184_6
timestamp 1731220651
transform 1 0 656 0 1 1844
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5183_6
timestamp 1731220651
transform 1 0 712 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5182_6
timestamp 1731220651
transform 1 0 640 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5181_6
timestamp 1731220651
transform 1 0 568 0 -1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5180_6
timestamp 1731220651
transform 1 0 608 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5179_6
timestamp 1731220651
transform 1 0 672 0 1 1984
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5178_6
timestamp 1731220651
transform 1 0 664 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5177_6
timestamp 1731220651
transform 1 0 600 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5176_6
timestamp 1731220651
transform 1 0 536 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5175_6
timestamp 1731220651
transform 1 0 592 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5174_6
timestamp 1731220651
transform 1 0 512 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5173_6
timestamp 1731220651
transform 1 0 472 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5172_6
timestamp 1731220651
transform 1 0 552 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5171_6
timestamp 1731220651
transform 1 0 544 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5170_6
timestamp 1731220651
transform 1 0 464 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5169_6
timestamp 1731220651
transform 1 0 264 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5168_6
timestamp 1731220651
transform 1 0 320 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5167_6
timestamp 1731220651
transform 1 0 392 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5166_6
timestamp 1731220651
transform 1 0 392 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5165_6
timestamp 1731220651
transform 1 0 320 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5164_6
timestamp 1731220651
transform 1 0 256 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5163_6
timestamp 1731220651
transform 1 0 192 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5162_6
timestamp 1731220651
transform 1 0 224 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5161_6
timestamp 1731220651
transform 1 0 264 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5160_6
timestamp 1731220651
transform 1 0 304 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5159_6
timestamp 1731220651
transform 1 0 344 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5158_6
timestamp 1731220651
transform 1 0 392 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5157_6
timestamp 1731220651
transform 1 0 448 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5156_6
timestamp 1731220651
transform 1 0 504 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5155_6
timestamp 1731220651
transform 1 0 568 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5154_6
timestamp 1731220651
transform 1 0 632 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5153_6
timestamp 1731220651
transform 1 0 464 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5152_6
timestamp 1731220651
transform 1 0 536 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5151_6
timestamp 1731220651
transform 1 0 608 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5150_6
timestamp 1731220651
transform 1 0 680 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5149_6
timestamp 1731220651
transform 1 0 704 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5148_6
timestamp 1731220651
transform 1 0 624 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5147_6
timestamp 1731220651
transform 1 0 640 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5146_6
timestamp 1731220651
transform 1 0 720 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5145_6
timestamp 1731220651
transform 1 0 800 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5144_6
timestamp 1731220651
transform 1 0 824 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5143_6
timestamp 1731220651
transform 1 0 752 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5142_6
timestamp 1731220651
transform 1 0 672 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5141_6
timestamp 1731220651
transform 1 0 728 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5140_6
timestamp 1731220651
transform 1 0 784 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5139_6
timestamp 1731220651
transform 1 0 832 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5138_6
timestamp 1731220651
transform 1 0 880 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5137_6
timestamp 1731220651
transform 1 0 928 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5136_6
timestamp 1731220651
transform 1 0 984 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5135_6
timestamp 1731220651
transform 1 0 1040 0 -1 2124
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5134_6
timestamp 1731220651
transform 1 0 896 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5133_6
timestamp 1731220651
transform 1 0 968 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5132_6
timestamp 1731220651
transform 1 0 1040 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5131_6
timestamp 1731220651
transform 1 0 1112 0 1 2132
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5130_6
timestamp 1731220651
transform 1 0 1120 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5129_6
timestamp 1731220651
transform 1 0 1040 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5128_6
timestamp 1731220651
transform 1 0 880 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5127_6
timestamp 1731220651
transform 1 0 960 0 -1 2268
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5126_6
timestamp 1731220651
transform 1 0 984 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5125_6
timestamp 1731220651
transform 1 0 1056 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5124_6
timestamp 1731220651
transform 1 0 912 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5123_6
timestamp 1731220651
transform 1 0 776 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5122_6
timestamp 1731220651
transform 1 0 848 0 1 2276
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5121_6
timestamp 1731220651
transform 1 0 888 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5120_6
timestamp 1731220651
transform 1 0 960 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5119_6
timestamp 1731220651
transform 1 0 816 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5118_6
timestamp 1731220651
transform 1 0 744 0 -1 2416
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5117_6
timestamp 1731220651
transform 1 0 696 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5116_6
timestamp 1731220651
transform 1 0 760 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5115_6
timestamp 1731220651
transform 1 0 816 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5114_6
timestamp 1731220651
transform 1 0 872 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5113_6
timestamp 1731220651
transform 1 0 920 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5112_6
timestamp 1731220651
transform 1 0 968 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5111_6
timestamp 1731220651
transform 1 0 1016 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5110_6
timestamp 1731220651
transform 1 0 1064 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5109_6
timestamp 1731220651
transform 1 0 1104 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5108_6
timestamp 1731220651
transform 1 0 1144 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5107_6
timestamp 1731220651
transform 1 0 1184 0 1 2424
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5106_6
timestamp 1731220651
transform 1 0 1296 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5105_6
timestamp 1731220651
transform 1 0 1336 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5104_6
timestamp 1731220651
transform 1 0 1376 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5103_6
timestamp 1731220651
transform 1 0 1432 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5102_6
timestamp 1731220651
transform 1 0 1504 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5101_6
timestamp 1731220651
transform 1 0 1576 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_5100_6
timestamp 1731220651
transform 1 0 1656 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_599_6
timestamp 1731220651
transform 1 0 1368 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_598_6
timestamp 1731220651
transform 1 0 1408 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_597_6
timestamp 1731220651
transform 1 0 1448 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_596_6
timestamp 1731220651
transform 1 0 1496 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_595_6
timestamp 1731220651
transform 1 0 1552 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_594_6
timestamp 1731220651
transform 1 0 1608 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_593_6
timestamp 1731220651
transform 1 0 1672 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_592_6
timestamp 1731220651
transform 1 0 1568 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_591_6
timestamp 1731220651
transform 1 0 1496 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_590_6
timestamp 1731220651
transform 1 0 1432 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_589_6
timestamp 1731220651
transform 1 0 1376 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_588_6
timestamp 1731220651
transform 1 0 1320 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_587_6
timestamp 1731220651
transform 1 0 1328 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_586_6
timestamp 1731220651
transform 1 0 1400 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_585_6
timestamp 1731220651
transform 1 0 1480 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_584_6
timestamp 1731220651
transform 1 0 1504 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_583_6
timestamp 1731220651
transform 1 0 1432 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_582_6
timestamp 1731220651
transform 1 0 1368 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_581_6
timestamp 1731220651
transform 1 0 1392 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_580_6
timestamp 1731220651
transform 1 0 1432 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_579_6
timestamp 1731220651
transform 1 0 1488 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_578_6
timestamp 1731220651
transform 1 0 1560 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_577_6
timestamp 1731220651
transform 1 0 1640 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_576_6
timestamp 1731220651
transform 1 0 1728 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_575_6
timestamp 1731220651
transform 1 0 1816 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_574_6
timestamp 1731220651
transform 1 0 1744 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_573_6
timestamp 1731220651
transform 1 0 1664 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_572_6
timestamp 1731220651
transform 1 0 1584 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_571_6
timestamp 1731220651
transform 1 0 1552 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_570_6
timestamp 1731220651
transform 1 0 1624 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_569_6
timestamp 1731220651
transform 1 0 1696 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_568_6
timestamp 1731220651
transform 1 0 1768 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_567_6
timestamp 1731220651
transform 1 0 1640 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_566_6
timestamp 1731220651
transform 1 0 1712 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_565_6
timestamp 1731220651
transform 1 0 1792 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_564_6
timestamp 1731220651
transform 1 0 1872 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_563_6
timestamp 1731220651
transform 1 0 1728 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_562_6
timestamp 1731220651
transform 1 0 1792 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_561_6
timestamp 1731220651
transform 1 0 1864 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_560_6
timestamp 1731220651
transform 1 0 1944 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_559_6
timestamp 1731220651
transform 1 0 1728 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_558_6
timestamp 1731220651
transform 1 0 1800 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_557_6
timestamp 1731220651
transform 1 0 1880 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_556_6
timestamp 1731220651
transform 1 0 1960 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_555_6
timestamp 1731220651
transform 1 0 2056 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_554_6
timestamp 1731220651
transform 1 0 2160 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_553_6
timestamp 1731220651
transform 1 0 2264 0 1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_552_6
timestamp 1731220651
transform 1 0 2256 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_551_6
timestamp 1731220651
transform 1 0 2040 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_550_6
timestamp 1731220651
transform 1 0 2144 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_549_6
timestamp 1731220651
transform 1 0 2160 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_548_6
timestamp 1731220651
transform 1 0 2056 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_547_6
timestamp 1731220651
transform 1 0 1960 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_546_6
timestamp 1731220651
transform 1 0 1832 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_545_6
timestamp 1731220651
transform 1 0 1904 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_544_6
timestamp 1731220651
transform 1 0 1984 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_543_6
timestamp 1731220651
transform 1 0 2072 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_542_6
timestamp 1731220651
transform 1 0 2168 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_541_6
timestamp 1731220651
transform 1 0 2272 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_540_6
timestamp 1731220651
transform 1 0 1824 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_539_6
timestamp 1731220651
transform 1 0 1896 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_538_6
timestamp 1731220651
transform 1 0 1960 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_537_6
timestamp 1731220651
transform 1 0 2024 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_536_6
timestamp 1731220651
transform 1 0 2088 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_535_6
timestamp 1731220651
transform 1 0 2160 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_534_6
timestamp 1731220651
transform 1 0 2232 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_533_6
timestamp 1731220651
transform 1 0 1904 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_532_6
timestamp 1731220651
transform 1 0 1992 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_531_6
timestamp 1731220651
transform 1 0 2080 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_530_6
timestamp 1731220651
transform 1 0 2168 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_529_6
timestamp 1731220651
transform 1 0 2264 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_528_6
timestamp 1731220651
transform 1 0 2072 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_527_6
timestamp 1731220651
transform 1 0 2032 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_526_6
timestamp 1731220651
transform 1 0 1912 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_525_6
timestamp 1731220651
transform 1 0 1960 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_524_6
timestamp 1731220651
transform 1 0 2008 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_523_6
timestamp 1731220651
transform 1 0 2144 0 1 1860
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_522_6
timestamp 1731220651
transform 1 0 2048 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_521_6
timestamp 1731220651
transform 1 0 2088 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_520_6
timestamp 1731220651
transform 1 0 2136 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_519_6
timestamp 1731220651
transform 1 0 2184 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_518_6
timestamp 1731220651
transform 1 0 2112 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_517_6
timestamp 1731220651
transform 1 0 2152 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_516_6
timestamp 1731220651
transform 1 0 2192 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_515_6
timestamp 1731220651
transform 1 0 2232 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_514_6
timestamp 1731220651
transform 1 0 2272 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_513_6
timestamp 1731220651
transform 1 0 2232 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_512_6
timestamp 1731220651
transform 1 0 2272 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_511_6
timestamp 1731220651
transform 1 0 2312 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_510_6
timestamp 1731220651
transform 1 0 2352 0 -1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_59_6
timestamp 1731220651
transform 1 0 2352 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_58_6
timestamp 1731220651
transform 1 0 2312 0 1 2000
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_57_6
timestamp 1731220651
transform 1 0 2352 0 -1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_56_6
timestamp 1731220651
transform 1 0 2304 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_55_6
timestamp 1731220651
transform 1 0 2352 0 1 2136
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_54_6
timestamp 1731220651
transform 1 0 2352 0 -1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_53_6
timestamp 1731220651
transform 1 0 2264 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_52_6
timestamp 1731220651
transform 1 0 2352 0 1 2280
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_51_6
timestamp 1731220651
transform 1 0 2352 0 -1 2420
box 4 6 36 64
use _0_0std_0_0cells_0_0NOR2X2  tst_50_6
timestamp 1731220651
transform 1 0 2352 0 1 2420
box 4 6 36 64
<< end >>
