magic
tech sky130l
timestamp 1730998298
<< ndiffusion >>
rect 8 6 13 16
rect 15 6 20 16
rect 22 10 27 16
rect 33 10 38 16
rect 40 10 47 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 43 6 47 10
rect 49 6 54 16
rect 60 6 65 16
rect 67 6 72 16
<< ndc >>
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 38 10 40 16
rect 47 6 49 16
rect 65 6 67 16
<< pdiffusion >>
rect 8 23 13 38
rect 15 31 19 38
rect 15 23 20 31
rect 22 23 27 31
rect 33 23 38 38
rect 40 23 47 38
rect 49 23 54 38
rect 60 23 65 38
rect 67 23 72 38
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 31
rect 38 23 40 38
rect 47 23 49 38
rect 65 23 67 38
<< polysilicon >>
rect 10 46 15 47
rect 10 43 11 46
rect 14 43 15 46
rect 10 42 15 43
rect 13 38 15 42
rect 20 46 25 47
rect 20 43 21 46
rect 24 43 25 46
rect 20 42 25 43
rect 38 46 43 47
rect 38 43 39 46
rect 42 43 43 46
rect 38 42 43 43
rect 20 31 22 42
rect 38 38 40 42
rect 47 38 49 40
rect 65 38 67 40
rect 13 16 15 23
rect 20 16 22 23
rect 38 16 40 23
rect 47 16 49 23
rect 65 21 67 23
rect 65 16 67 18
rect 38 8 40 10
rect 13 4 15 6
rect 20 4 22 6
rect 47 4 49 6
rect 65 4 67 6
<< pc >>
rect 11 43 14 46
rect 21 43 24 46
rect 39 43 42 46
<< m1 >>
rect 8 46 15 47
rect 8 43 11 46
rect 14 43 15 46
rect 8 42 15 43
rect 20 46 25 47
rect 20 43 21 46
rect 24 43 25 46
rect 20 42 25 43
rect 38 46 44 47
rect 38 43 39 46
rect 42 43 44 46
rect 38 42 44 43
rect 8 40 12 42
rect 40 40 44 42
rect 56 40 60 44
rect 72 40 76 44
rect 23 10 27 11
rect 8 4 12 8
rect 26 8 27 10
rect 33 8 37 14
rect 26 7 28 8
rect 23 4 28 7
rect 32 4 36 8
<< m2c >>
rect 21 43 24 46
rect 39 43 42 46
<< m2 >>
rect 20 46 44 47
rect 20 43 21 46
rect 24 43 39 46
rect 42 43 44 46
rect 20 42 44 43
<< labels >>
rlabel space 0 0 80 48 6 prboundary
rlabel pdiffusion 23 24 23 24 3 _S
rlabel ndiffusion 23 7 23 7 3 Y
rlabel polysilicon 21 17 21 17 3 S
rlabel polysilicon 21 22 21 22 3 S
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel polysilicon 14 17 14 17 3 A
rlabel polysilicon 14 22 14 22 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 #5
rlabel ndiffusion 50 7 50 7 3 #10
rlabel polysilicon 48 17 48 17 3 B
rlabel polysilicon 48 22 48 22 3 B
rlabel pdiffusion 50 24 50 24 3 Vdd
rlabel ndiffusion 41 11 41 11 3 GND
rlabel polysilicon 39 17 39 17 3 S
rlabel polysilicon 39 22 39 22 3 S
rlabel ndiffusion 34 11 34 11 3 _S
rlabel pdiffusion 34 24 34 24 3 Y
rlabel ndiffusion 68 7 68 7 3 #10
rlabel pdiffusion 68 24 68 24 3 Y
rlabel polysilicon 66 17 66 17 3 _S
rlabel polysilicon 66 22 66 22 3 _S
rlabel ndiffusion 61 7 61 7 3 Y
rlabel pdiffusion 61 24 61 24 3 #5
rlabel m1 73 41 73 41 3 GND
port 1 e
rlabel m1 57 41 57 41 3 Vdd
port 2 e
rlabel m1 41 41 41 41 3 S
port 3 e
rlabel m1 9 41 9 41 3 A
port 6 e
rlabel m1 24 5 24 5 1 Y
<< end >>
