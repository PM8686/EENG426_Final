magic
tech sky130l
timestamp 1731220342
<< m2 >>
rect 2046 4004 2052 4005
rect 3942 4004 3948 4005
rect 2046 4000 2047 4004
rect 2051 4000 2052 4004
rect 2046 3999 2052 4000
rect 2070 4003 2076 4004
rect 2070 3999 2071 4003
rect 2075 3999 2076 4003
rect 3942 4000 3943 4004
rect 3947 4000 3948 4004
rect 3942 3999 3948 4000
rect 2070 3998 2076 3999
rect 2046 3987 2052 3988
rect 110 3984 116 3985
rect 2006 3984 2012 3985
rect 110 3980 111 3984
rect 115 3980 116 3984
rect 110 3979 116 3980
rect 150 3983 156 3984
rect 150 3979 151 3983
rect 155 3979 156 3983
rect 150 3978 156 3979
rect 278 3983 284 3984
rect 278 3979 279 3983
rect 283 3979 284 3983
rect 278 3978 284 3979
rect 430 3983 436 3984
rect 430 3979 431 3983
rect 435 3979 436 3983
rect 430 3978 436 3979
rect 606 3983 612 3984
rect 606 3979 607 3983
rect 611 3979 612 3983
rect 606 3978 612 3979
rect 790 3983 796 3984
rect 790 3979 791 3983
rect 795 3979 796 3983
rect 790 3978 796 3979
rect 974 3983 980 3984
rect 974 3979 975 3983
rect 979 3979 980 3983
rect 974 3978 980 3979
rect 1150 3983 1156 3984
rect 1150 3979 1151 3983
rect 1155 3979 1156 3983
rect 1150 3978 1156 3979
rect 1310 3983 1316 3984
rect 1310 3979 1311 3983
rect 1315 3979 1316 3983
rect 1310 3978 1316 3979
rect 1470 3983 1476 3984
rect 1470 3979 1471 3983
rect 1475 3979 1476 3983
rect 1470 3978 1476 3979
rect 1622 3983 1628 3984
rect 1622 3979 1623 3983
rect 1627 3979 1628 3983
rect 1622 3978 1628 3979
rect 1774 3983 1780 3984
rect 1774 3979 1775 3983
rect 1779 3979 1780 3983
rect 1774 3978 1780 3979
rect 1902 3983 1908 3984
rect 1902 3979 1903 3983
rect 1907 3979 1908 3983
rect 2006 3980 2007 3984
rect 2011 3980 2012 3984
rect 2046 3983 2047 3987
rect 2051 3983 2052 3987
rect 3942 3987 3948 3988
rect 2046 3982 2052 3983
rect 2070 3984 2076 3985
rect 2006 3979 2012 3980
rect 2070 3980 2071 3984
rect 2075 3980 2076 3984
rect 3942 3983 3943 3987
rect 3947 3983 3948 3987
rect 3942 3982 3948 3983
rect 2070 3979 2076 3980
rect 1902 3978 1908 3979
rect 110 3967 116 3968
rect 110 3963 111 3967
rect 115 3963 116 3967
rect 2006 3967 2012 3968
rect 110 3962 116 3963
rect 150 3964 156 3965
rect 150 3960 151 3964
rect 155 3960 156 3964
rect 150 3959 156 3960
rect 278 3964 284 3965
rect 278 3960 279 3964
rect 283 3960 284 3964
rect 278 3959 284 3960
rect 430 3964 436 3965
rect 430 3960 431 3964
rect 435 3960 436 3964
rect 430 3959 436 3960
rect 606 3964 612 3965
rect 606 3960 607 3964
rect 611 3960 612 3964
rect 606 3959 612 3960
rect 790 3964 796 3965
rect 790 3960 791 3964
rect 795 3960 796 3964
rect 790 3959 796 3960
rect 974 3964 980 3965
rect 974 3960 975 3964
rect 979 3960 980 3964
rect 974 3959 980 3960
rect 1150 3964 1156 3965
rect 1150 3960 1151 3964
rect 1155 3960 1156 3964
rect 1150 3959 1156 3960
rect 1310 3964 1316 3965
rect 1310 3960 1311 3964
rect 1315 3960 1316 3964
rect 1310 3959 1316 3960
rect 1470 3964 1476 3965
rect 1470 3960 1471 3964
rect 1475 3960 1476 3964
rect 1470 3959 1476 3960
rect 1622 3964 1628 3965
rect 1622 3960 1623 3964
rect 1627 3960 1628 3964
rect 1622 3959 1628 3960
rect 1774 3964 1780 3965
rect 1774 3960 1775 3964
rect 1779 3960 1780 3964
rect 1774 3959 1780 3960
rect 1902 3964 1908 3965
rect 1902 3960 1903 3964
rect 1907 3960 1908 3964
rect 2006 3963 2007 3967
rect 2011 3963 2012 3967
rect 2006 3962 2012 3963
rect 1902 3959 1908 3960
rect 2078 3924 2084 3925
rect 2046 3921 2052 3922
rect 2046 3917 2047 3921
rect 2051 3917 2052 3921
rect 2078 3920 2079 3924
rect 2083 3920 2084 3924
rect 2078 3919 2084 3920
rect 2214 3924 2220 3925
rect 2214 3920 2215 3924
rect 2219 3920 2220 3924
rect 2214 3919 2220 3920
rect 2358 3924 2364 3925
rect 2358 3920 2359 3924
rect 2363 3920 2364 3924
rect 2358 3919 2364 3920
rect 2502 3924 2508 3925
rect 2502 3920 2503 3924
rect 2507 3920 2508 3924
rect 2502 3919 2508 3920
rect 2646 3924 2652 3925
rect 2646 3920 2647 3924
rect 2651 3920 2652 3924
rect 2646 3919 2652 3920
rect 2790 3924 2796 3925
rect 2790 3920 2791 3924
rect 2795 3920 2796 3924
rect 2790 3919 2796 3920
rect 2926 3924 2932 3925
rect 2926 3920 2927 3924
rect 2931 3920 2932 3924
rect 2926 3919 2932 3920
rect 3054 3924 3060 3925
rect 3054 3920 3055 3924
rect 3059 3920 3060 3924
rect 3054 3919 3060 3920
rect 3174 3924 3180 3925
rect 3174 3920 3175 3924
rect 3179 3920 3180 3924
rect 3174 3919 3180 3920
rect 3294 3924 3300 3925
rect 3294 3920 3295 3924
rect 3299 3920 3300 3924
rect 3294 3919 3300 3920
rect 3414 3924 3420 3925
rect 3414 3920 3415 3924
rect 3419 3920 3420 3924
rect 3414 3919 3420 3920
rect 3534 3924 3540 3925
rect 3534 3920 3535 3924
rect 3539 3920 3540 3924
rect 3534 3919 3540 3920
rect 3942 3921 3948 3922
rect 2046 3916 2052 3917
rect 3942 3917 3943 3921
rect 3947 3917 3948 3921
rect 3942 3916 3948 3917
rect 2078 3905 2084 3906
rect 302 3904 308 3905
rect 110 3901 116 3902
rect 110 3897 111 3901
rect 115 3897 116 3901
rect 302 3900 303 3904
rect 307 3900 308 3904
rect 302 3899 308 3900
rect 422 3904 428 3905
rect 422 3900 423 3904
rect 427 3900 428 3904
rect 422 3899 428 3900
rect 550 3904 556 3905
rect 550 3900 551 3904
rect 555 3900 556 3904
rect 550 3899 556 3900
rect 686 3904 692 3905
rect 686 3900 687 3904
rect 691 3900 692 3904
rect 686 3899 692 3900
rect 814 3904 820 3905
rect 814 3900 815 3904
rect 819 3900 820 3904
rect 814 3899 820 3900
rect 942 3904 948 3905
rect 942 3900 943 3904
rect 947 3900 948 3904
rect 942 3899 948 3900
rect 1070 3904 1076 3905
rect 1070 3900 1071 3904
rect 1075 3900 1076 3904
rect 1070 3899 1076 3900
rect 1198 3904 1204 3905
rect 1198 3900 1199 3904
rect 1203 3900 1204 3904
rect 1198 3899 1204 3900
rect 1326 3904 1332 3905
rect 1326 3900 1327 3904
rect 1331 3900 1332 3904
rect 1326 3899 1332 3900
rect 1462 3904 1468 3905
rect 1462 3900 1463 3904
rect 1467 3900 1468 3904
rect 2046 3904 2052 3905
rect 1462 3899 1468 3900
rect 2006 3901 2012 3902
rect 110 3896 116 3897
rect 2006 3897 2007 3901
rect 2011 3897 2012 3901
rect 2046 3900 2047 3904
rect 2051 3900 2052 3904
rect 2078 3901 2079 3905
rect 2083 3901 2084 3905
rect 2078 3900 2084 3901
rect 2214 3905 2220 3906
rect 2214 3901 2215 3905
rect 2219 3901 2220 3905
rect 2214 3900 2220 3901
rect 2358 3905 2364 3906
rect 2358 3901 2359 3905
rect 2363 3901 2364 3905
rect 2358 3900 2364 3901
rect 2502 3905 2508 3906
rect 2502 3901 2503 3905
rect 2507 3901 2508 3905
rect 2502 3900 2508 3901
rect 2646 3905 2652 3906
rect 2646 3901 2647 3905
rect 2651 3901 2652 3905
rect 2646 3900 2652 3901
rect 2790 3905 2796 3906
rect 2790 3901 2791 3905
rect 2795 3901 2796 3905
rect 2790 3900 2796 3901
rect 2926 3905 2932 3906
rect 2926 3901 2927 3905
rect 2931 3901 2932 3905
rect 2926 3900 2932 3901
rect 3054 3905 3060 3906
rect 3054 3901 3055 3905
rect 3059 3901 3060 3905
rect 3054 3900 3060 3901
rect 3174 3905 3180 3906
rect 3174 3901 3175 3905
rect 3179 3901 3180 3905
rect 3174 3900 3180 3901
rect 3294 3905 3300 3906
rect 3294 3901 3295 3905
rect 3299 3901 3300 3905
rect 3294 3900 3300 3901
rect 3414 3905 3420 3906
rect 3414 3901 3415 3905
rect 3419 3901 3420 3905
rect 3414 3900 3420 3901
rect 3534 3905 3540 3906
rect 3534 3901 3535 3905
rect 3539 3901 3540 3905
rect 3534 3900 3540 3901
rect 3942 3904 3948 3905
rect 3942 3900 3943 3904
rect 3947 3900 3948 3904
rect 2046 3899 2052 3900
rect 3942 3899 3948 3900
rect 2006 3896 2012 3897
rect 302 3885 308 3886
rect 110 3884 116 3885
rect 110 3880 111 3884
rect 115 3880 116 3884
rect 302 3881 303 3885
rect 307 3881 308 3885
rect 302 3880 308 3881
rect 422 3885 428 3886
rect 422 3881 423 3885
rect 427 3881 428 3885
rect 422 3880 428 3881
rect 550 3885 556 3886
rect 550 3881 551 3885
rect 555 3881 556 3885
rect 550 3880 556 3881
rect 686 3885 692 3886
rect 686 3881 687 3885
rect 691 3881 692 3885
rect 686 3880 692 3881
rect 814 3885 820 3886
rect 814 3881 815 3885
rect 819 3881 820 3885
rect 814 3880 820 3881
rect 942 3885 948 3886
rect 942 3881 943 3885
rect 947 3881 948 3885
rect 942 3880 948 3881
rect 1070 3885 1076 3886
rect 1070 3881 1071 3885
rect 1075 3881 1076 3885
rect 1070 3880 1076 3881
rect 1198 3885 1204 3886
rect 1198 3881 1199 3885
rect 1203 3881 1204 3885
rect 1198 3880 1204 3881
rect 1326 3885 1332 3886
rect 1326 3881 1327 3885
rect 1331 3881 1332 3885
rect 1326 3880 1332 3881
rect 1462 3885 1468 3886
rect 1462 3881 1463 3885
rect 1467 3881 1468 3885
rect 1462 3880 1468 3881
rect 2006 3884 2012 3885
rect 2006 3880 2007 3884
rect 2011 3880 2012 3884
rect 110 3879 116 3880
rect 2006 3879 2012 3880
rect 2046 3852 2052 3853
rect 3942 3852 3948 3853
rect 2046 3848 2047 3852
rect 2051 3848 2052 3852
rect 2046 3847 2052 3848
rect 2254 3851 2260 3852
rect 2254 3847 2255 3851
rect 2259 3847 2260 3851
rect 2254 3846 2260 3847
rect 2382 3851 2388 3852
rect 2382 3847 2383 3851
rect 2387 3847 2388 3851
rect 2382 3846 2388 3847
rect 2518 3851 2524 3852
rect 2518 3847 2519 3851
rect 2523 3847 2524 3851
rect 2518 3846 2524 3847
rect 2670 3851 2676 3852
rect 2670 3847 2671 3851
rect 2675 3847 2676 3851
rect 2670 3846 2676 3847
rect 2830 3851 2836 3852
rect 2830 3847 2831 3851
rect 2835 3847 2836 3851
rect 2830 3846 2836 3847
rect 2990 3851 2996 3852
rect 2990 3847 2991 3851
rect 2995 3847 2996 3851
rect 2990 3846 2996 3847
rect 3158 3851 3164 3852
rect 3158 3847 3159 3851
rect 3163 3847 3164 3851
rect 3158 3846 3164 3847
rect 3326 3851 3332 3852
rect 3326 3847 3327 3851
rect 3331 3847 3332 3851
rect 3326 3846 3332 3847
rect 3494 3851 3500 3852
rect 3494 3847 3495 3851
rect 3499 3847 3500 3851
rect 3494 3846 3500 3847
rect 3662 3851 3668 3852
rect 3662 3847 3663 3851
rect 3667 3847 3668 3851
rect 3942 3848 3943 3852
rect 3947 3848 3948 3852
rect 3942 3847 3948 3848
rect 3662 3846 3668 3847
rect 2046 3835 2052 3836
rect 2046 3831 2047 3835
rect 2051 3831 2052 3835
rect 3942 3835 3948 3836
rect 2046 3830 2052 3831
rect 2254 3832 2260 3833
rect 110 3828 116 3829
rect 2006 3828 2012 3829
rect 110 3824 111 3828
rect 115 3824 116 3828
rect 110 3823 116 3824
rect 414 3827 420 3828
rect 414 3823 415 3827
rect 419 3823 420 3827
rect 414 3822 420 3823
rect 566 3827 572 3828
rect 566 3823 567 3827
rect 571 3823 572 3827
rect 566 3822 572 3823
rect 726 3827 732 3828
rect 726 3823 727 3827
rect 731 3823 732 3827
rect 726 3822 732 3823
rect 886 3827 892 3828
rect 886 3823 887 3827
rect 891 3823 892 3827
rect 886 3822 892 3823
rect 1038 3827 1044 3828
rect 1038 3823 1039 3827
rect 1043 3823 1044 3827
rect 1038 3822 1044 3823
rect 1190 3827 1196 3828
rect 1190 3823 1191 3827
rect 1195 3823 1196 3827
rect 1190 3822 1196 3823
rect 1342 3827 1348 3828
rect 1342 3823 1343 3827
rect 1347 3823 1348 3827
rect 1342 3822 1348 3823
rect 1494 3827 1500 3828
rect 1494 3823 1495 3827
rect 1499 3823 1500 3827
rect 1494 3822 1500 3823
rect 1646 3827 1652 3828
rect 1646 3823 1647 3827
rect 1651 3823 1652 3827
rect 2006 3824 2007 3828
rect 2011 3824 2012 3828
rect 2254 3828 2255 3832
rect 2259 3828 2260 3832
rect 2254 3827 2260 3828
rect 2382 3832 2388 3833
rect 2382 3828 2383 3832
rect 2387 3828 2388 3832
rect 2382 3827 2388 3828
rect 2518 3832 2524 3833
rect 2518 3828 2519 3832
rect 2523 3828 2524 3832
rect 2518 3827 2524 3828
rect 2670 3832 2676 3833
rect 2670 3828 2671 3832
rect 2675 3828 2676 3832
rect 2670 3827 2676 3828
rect 2830 3832 2836 3833
rect 2830 3828 2831 3832
rect 2835 3828 2836 3832
rect 2830 3827 2836 3828
rect 2990 3832 2996 3833
rect 2990 3828 2991 3832
rect 2995 3828 2996 3832
rect 2990 3827 2996 3828
rect 3158 3832 3164 3833
rect 3158 3828 3159 3832
rect 3163 3828 3164 3832
rect 3158 3827 3164 3828
rect 3326 3832 3332 3833
rect 3326 3828 3327 3832
rect 3331 3828 3332 3832
rect 3326 3827 3332 3828
rect 3494 3832 3500 3833
rect 3494 3828 3495 3832
rect 3499 3828 3500 3832
rect 3494 3827 3500 3828
rect 3662 3832 3668 3833
rect 3662 3828 3663 3832
rect 3667 3828 3668 3832
rect 3942 3831 3943 3835
rect 3947 3831 3948 3835
rect 3942 3830 3948 3831
rect 3662 3827 3668 3828
rect 2006 3823 2012 3824
rect 1646 3822 1652 3823
rect 110 3811 116 3812
rect 110 3807 111 3811
rect 115 3807 116 3811
rect 2006 3811 2012 3812
rect 110 3806 116 3807
rect 414 3808 420 3809
rect 414 3804 415 3808
rect 419 3804 420 3808
rect 414 3803 420 3804
rect 566 3808 572 3809
rect 566 3804 567 3808
rect 571 3804 572 3808
rect 566 3803 572 3804
rect 726 3808 732 3809
rect 726 3804 727 3808
rect 731 3804 732 3808
rect 726 3803 732 3804
rect 886 3808 892 3809
rect 886 3804 887 3808
rect 891 3804 892 3808
rect 886 3803 892 3804
rect 1038 3808 1044 3809
rect 1038 3804 1039 3808
rect 1043 3804 1044 3808
rect 1038 3803 1044 3804
rect 1190 3808 1196 3809
rect 1190 3804 1191 3808
rect 1195 3804 1196 3808
rect 1190 3803 1196 3804
rect 1342 3808 1348 3809
rect 1342 3804 1343 3808
rect 1347 3804 1348 3808
rect 1342 3803 1348 3804
rect 1494 3808 1500 3809
rect 1494 3804 1495 3808
rect 1499 3804 1500 3808
rect 1494 3803 1500 3804
rect 1646 3808 1652 3809
rect 1646 3804 1647 3808
rect 1651 3804 1652 3808
rect 2006 3807 2007 3811
rect 2011 3807 2012 3811
rect 2006 3806 2012 3807
rect 1646 3803 1652 3804
rect 2070 3772 2076 3773
rect 2046 3769 2052 3770
rect 2046 3765 2047 3769
rect 2051 3765 2052 3769
rect 2070 3768 2071 3772
rect 2075 3768 2076 3772
rect 2070 3767 2076 3768
rect 2198 3772 2204 3773
rect 2198 3768 2199 3772
rect 2203 3768 2204 3772
rect 2198 3767 2204 3768
rect 2374 3772 2380 3773
rect 2374 3768 2375 3772
rect 2379 3768 2380 3772
rect 2374 3767 2380 3768
rect 2558 3772 2564 3773
rect 2558 3768 2559 3772
rect 2563 3768 2564 3772
rect 2558 3767 2564 3768
rect 2750 3772 2756 3773
rect 2750 3768 2751 3772
rect 2755 3768 2756 3772
rect 2750 3767 2756 3768
rect 2950 3772 2956 3773
rect 2950 3768 2951 3772
rect 2955 3768 2956 3772
rect 2950 3767 2956 3768
rect 3142 3772 3148 3773
rect 3142 3768 3143 3772
rect 3147 3768 3148 3772
rect 3142 3767 3148 3768
rect 3334 3772 3340 3773
rect 3334 3768 3335 3772
rect 3339 3768 3340 3772
rect 3334 3767 3340 3768
rect 3534 3772 3540 3773
rect 3534 3768 3535 3772
rect 3539 3768 3540 3772
rect 3534 3767 3540 3768
rect 3734 3772 3740 3773
rect 3734 3768 3735 3772
rect 3739 3768 3740 3772
rect 3734 3767 3740 3768
rect 3942 3769 3948 3770
rect 2046 3764 2052 3765
rect 3942 3765 3943 3769
rect 3947 3765 3948 3769
rect 3942 3764 3948 3765
rect 2070 3753 2076 3754
rect 2046 3752 2052 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2070 3749 2071 3753
rect 2075 3749 2076 3753
rect 2070 3748 2076 3749
rect 2198 3753 2204 3754
rect 2198 3749 2199 3753
rect 2203 3749 2204 3753
rect 2198 3748 2204 3749
rect 2374 3753 2380 3754
rect 2374 3749 2375 3753
rect 2379 3749 2380 3753
rect 2374 3748 2380 3749
rect 2558 3753 2564 3754
rect 2558 3749 2559 3753
rect 2563 3749 2564 3753
rect 2558 3748 2564 3749
rect 2750 3753 2756 3754
rect 2750 3749 2751 3753
rect 2755 3749 2756 3753
rect 2750 3748 2756 3749
rect 2950 3753 2956 3754
rect 2950 3749 2951 3753
rect 2955 3749 2956 3753
rect 2950 3748 2956 3749
rect 3142 3753 3148 3754
rect 3142 3749 3143 3753
rect 3147 3749 3148 3753
rect 3142 3748 3148 3749
rect 3334 3753 3340 3754
rect 3334 3749 3335 3753
rect 3339 3749 3340 3753
rect 3334 3748 3340 3749
rect 3534 3753 3540 3754
rect 3534 3749 3535 3753
rect 3539 3749 3540 3753
rect 3534 3748 3540 3749
rect 3734 3753 3740 3754
rect 3734 3749 3735 3753
rect 3739 3749 3740 3753
rect 3734 3748 3740 3749
rect 3942 3752 3948 3753
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 2046 3747 2052 3748
rect 3942 3747 3948 3748
rect 398 3744 404 3745
rect 110 3741 116 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 398 3740 399 3744
rect 403 3740 404 3744
rect 398 3739 404 3740
rect 566 3744 572 3745
rect 566 3740 567 3744
rect 571 3740 572 3744
rect 566 3739 572 3740
rect 750 3744 756 3745
rect 750 3740 751 3744
rect 755 3740 756 3744
rect 750 3739 756 3740
rect 934 3744 940 3745
rect 934 3740 935 3744
rect 939 3740 940 3744
rect 934 3739 940 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1310 3744 1316 3745
rect 1310 3740 1311 3744
rect 1315 3740 1316 3744
rect 1310 3739 1316 3740
rect 1502 3744 1508 3745
rect 1502 3740 1503 3744
rect 1507 3740 1508 3744
rect 1502 3739 1508 3740
rect 1694 3744 1700 3745
rect 1694 3740 1695 3744
rect 1699 3740 1700 3744
rect 1694 3739 1700 3740
rect 1886 3744 1892 3745
rect 1886 3740 1887 3744
rect 1891 3740 1892 3744
rect 1886 3739 1892 3740
rect 2006 3741 2012 3742
rect 110 3736 116 3737
rect 2006 3737 2007 3741
rect 2011 3737 2012 3741
rect 2006 3736 2012 3737
rect 398 3725 404 3726
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 398 3721 399 3725
rect 403 3721 404 3725
rect 398 3720 404 3721
rect 566 3725 572 3726
rect 566 3721 567 3725
rect 571 3721 572 3725
rect 566 3720 572 3721
rect 750 3725 756 3726
rect 750 3721 751 3725
rect 755 3721 756 3725
rect 750 3720 756 3721
rect 934 3725 940 3726
rect 934 3721 935 3725
rect 939 3721 940 3725
rect 934 3720 940 3721
rect 1126 3725 1132 3726
rect 1126 3721 1127 3725
rect 1131 3721 1132 3725
rect 1126 3720 1132 3721
rect 1310 3725 1316 3726
rect 1310 3721 1311 3725
rect 1315 3721 1316 3725
rect 1310 3720 1316 3721
rect 1502 3725 1508 3726
rect 1502 3721 1503 3725
rect 1507 3721 1508 3725
rect 1502 3720 1508 3721
rect 1694 3725 1700 3726
rect 1694 3721 1695 3725
rect 1699 3721 1700 3725
rect 1694 3720 1700 3721
rect 1886 3725 1892 3726
rect 1886 3721 1887 3725
rect 1891 3721 1892 3725
rect 1886 3720 1892 3721
rect 2006 3724 2012 3725
rect 2006 3720 2007 3724
rect 2011 3720 2012 3724
rect 110 3719 116 3720
rect 2006 3719 2012 3720
rect 2046 3688 2052 3689
rect 3942 3688 3948 3689
rect 2046 3684 2047 3688
rect 2051 3684 2052 3688
rect 2046 3683 2052 3684
rect 2070 3687 2076 3688
rect 2070 3683 2071 3687
rect 2075 3683 2076 3687
rect 2070 3682 2076 3683
rect 2262 3687 2268 3688
rect 2262 3683 2263 3687
rect 2267 3683 2268 3687
rect 2262 3682 2268 3683
rect 2478 3687 2484 3688
rect 2478 3683 2479 3687
rect 2483 3683 2484 3687
rect 2478 3682 2484 3683
rect 2694 3687 2700 3688
rect 2694 3683 2695 3687
rect 2699 3683 2700 3687
rect 2694 3682 2700 3683
rect 2910 3687 2916 3688
rect 2910 3683 2911 3687
rect 2915 3683 2916 3687
rect 2910 3682 2916 3683
rect 3118 3687 3124 3688
rect 3118 3683 3119 3687
rect 3123 3683 3124 3687
rect 3118 3682 3124 3683
rect 3318 3687 3324 3688
rect 3318 3683 3319 3687
rect 3323 3683 3324 3687
rect 3318 3682 3324 3683
rect 3518 3687 3524 3688
rect 3518 3683 3519 3687
rect 3523 3683 3524 3687
rect 3518 3682 3524 3683
rect 3726 3687 3732 3688
rect 3726 3683 3727 3687
rect 3731 3683 3732 3687
rect 3942 3684 3943 3688
rect 3947 3684 3948 3688
rect 3942 3683 3948 3684
rect 3726 3682 3732 3683
rect 2046 3671 2052 3672
rect 2046 3667 2047 3671
rect 2051 3667 2052 3671
rect 3942 3671 3948 3672
rect 2046 3666 2052 3667
rect 2070 3668 2076 3669
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 2262 3668 2268 3669
rect 2262 3664 2263 3668
rect 2267 3664 2268 3668
rect 2262 3663 2268 3664
rect 2478 3668 2484 3669
rect 2478 3664 2479 3668
rect 2483 3664 2484 3668
rect 2478 3663 2484 3664
rect 2694 3668 2700 3669
rect 2694 3664 2695 3668
rect 2699 3664 2700 3668
rect 2694 3663 2700 3664
rect 2910 3668 2916 3669
rect 2910 3664 2911 3668
rect 2915 3664 2916 3668
rect 2910 3663 2916 3664
rect 3118 3668 3124 3669
rect 3118 3664 3119 3668
rect 3123 3664 3124 3668
rect 3118 3663 3124 3664
rect 3318 3668 3324 3669
rect 3318 3664 3319 3668
rect 3323 3664 3324 3668
rect 3318 3663 3324 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3726 3668 3732 3669
rect 3726 3664 3727 3668
rect 3731 3664 3732 3668
rect 3942 3667 3943 3671
rect 3947 3667 3948 3671
rect 3942 3666 3948 3667
rect 3726 3663 3732 3664
rect 110 3660 116 3661
rect 2006 3660 2012 3661
rect 110 3656 111 3660
rect 115 3656 116 3660
rect 110 3655 116 3656
rect 366 3659 372 3660
rect 366 3655 367 3659
rect 371 3655 372 3659
rect 366 3654 372 3655
rect 518 3659 524 3660
rect 518 3655 519 3659
rect 523 3655 524 3659
rect 518 3654 524 3655
rect 678 3659 684 3660
rect 678 3655 679 3659
rect 683 3655 684 3659
rect 678 3654 684 3655
rect 846 3659 852 3660
rect 846 3655 847 3659
rect 851 3655 852 3659
rect 846 3654 852 3655
rect 1014 3659 1020 3660
rect 1014 3655 1015 3659
rect 1019 3655 1020 3659
rect 1014 3654 1020 3655
rect 1174 3659 1180 3660
rect 1174 3655 1175 3659
rect 1179 3655 1180 3659
rect 1174 3654 1180 3655
rect 1326 3659 1332 3660
rect 1326 3655 1327 3659
rect 1331 3655 1332 3659
rect 1326 3654 1332 3655
rect 1478 3659 1484 3660
rect 1478 3655 1479 3659
rect 1483 3655 1484 3659
rect 1478 3654 1484 3655
rect 1630 3659 1636 3660
rect 1630 3655 1631 3659
rect 1635 3655 1636 3659
rect 1630 3654 1636 3655
rect 1790 3659 1796 3660
rect 1790 3655 1791 3659
rect 1795 3655 1796 3659
rect 2006 3656 2007 3660
rect 2011 3656 2012 3660
rect 2006 3655 2012 3656
rect 1790 3654 1796 3655
rect 110 3643 116 3644
rect 110 3639 111 3643
rect 115 3639 116 3643
rect 2006 3643 2012 3644
rect 110 3638 116 3639
rect 366 3640 372 3641
rect 366 3636 367 3640
rect 371 3636 372 3640
rect 366 3635 372 3636
rect 518 3640 524 3641
rect 518 3636 519 3640
rect 523 3636 524 3640
rect 518 3635 524 3636
rect 678 3640 684 3641
rect 678 3636 679 3640
rect 683 3636 684 3640
rect 678 3635 684 3636
rect 846 3640 852 3641
rect 846 3636 847 3640
rect 851 3636 852 3640
rect 846 3635 852 3636
rect 1014 3640 1020 3641
rect 1014 3636 1015 3640
rect 1019 3636 1020 3640
rect 1014 3635 1020 3636
rect 1174 3640 1180 3641
rect 1174 3636 1175 3640
rect 1179 3636 1180 3640
rect 1174 3635 1180 3636
rect 1326 3640 1332 3641
rect 1326 3636 1327 3640
rect 1331 3636 1332 3640
rect 1326 3635 1332 3636
rect 1478 3640 1484 3641
rect 1478 3636 1479 3640
rect 1483 3636 1484 3640
rect 1478 3635 1484 3636
rect 1630 3640 1636 3641
rect 1630 3636 1631 3640
rect 1635 3636 1636 3640
rect 1630 3635 1636 3636
rect 1790 3640 1796 3641
rect 1790 3636 1791 3640
rect 1795 3636 1796 3640
rect 2006 3639 2007 3643
rect 2011 3639 2012 3643
rect 2006 3638 2012 3639
rect 1790 3635 1796 3636
rect 2110 3604 2116 3605
rect 2046 3601 2052 3602
rect 2046 3597 2047 3601
rect 2051 3597 2052 3601
rect 2110 3600 2111 3604
rect 2115 3600 2116 3604
rect 2110 3599 2116 3600
rect 2270 3604 2276 3605
rect 2270 3600 2271 3604
rect 2275 3600 2276 3604
rect 2270 3599 2276 3600
rect 2454 3604 2460 3605
rect 2454 3600 2455 3604
rect 2459 3600 2460 3604
rect 2454 3599 2460 3600
rect 2654 3604 2660 3605
rect 2654 3600 2655 3604
rect 2659 3600 2660 3604
rect 2654 3599 2660 3600
rect 2870 3604 2876 3605
rect 2870 3600 2871 3604
rect 2875 3600 2876 3604
rect 2870 3599 2876 3600
rect 3094 3604 3100 3605
rect 3094 3600 3095 3604
rect 3099 3600 3100 3604
rect 3094 3599 3100 3600
rect 3326 3604 3332 3605
rect 3326 3600 3327 3604
rect 3331 3600 3332 3604
rect 3326 3599 3332 3600
rect 3566 3604 3572 3605
rect 3566 3600 3567 3604
rect 3571 3600 3572 3604
rect 3566 3599 3572 3600
rect 3942 3601 3948 3602
rect 2046 3596 2052 3597
rect 3942 3597 3943 3601
rect 3947 3597 3948 3601
rect 3942 3596 3948 3597
rect 2110 3585 2116 3586
rect 2046 3584 2052 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2110 3581 2111 3585
rect 2115 3581 2116 3585
rect 2110 3580 2116 3581
rect 2270 3585 2276 3586
rect 2270 3581 2271 3585
rect 2275 3581 2276 3585
rect 2270 3580 2276 3581
rect 2454 3585 2460 3586
rect 2454 3581 2455 3585
rect 2459 3581 2460 3585
rect 2454 3580 2460 3581
rect 2654 3585 2660 3586
rect 2654 3581 2655 3585
rect 2659 3581 2660 3585
rect 2654 3580 2660 3581
rect 2870 3585 2876 3586
rect 2870 3581 2871 3585
rect 2875 3581 2876 3585
rect 2870 3580 2876 3581
rect 3094 3585 3100 3586
rect 3094 3581 3095 3585
rect 3099 3581 3100 3585
rect 3094 3580 3100 3581
rect 3326 3585 3332 3586
rect 3326 3581 3327 3585
rect 3331 3581 3332 3585
rect 3326 3580 3332 3581
rect 3566 3585 3572 3586
rect 3566 3581 3567 3585
rect 3571 3581 3572 3585
rect 3566 3580 3572 3581
rect 3942 3584 3948 3585
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 2046 3579 2052 3580
rect 3942 3579 3948 3580
rect 270 3572 276 3573
rect 110 3569 116 3570
rect 110 3565 111 3569
rect 115 3565 116 3569
rect 270 3568 271 3572
rect 275 3568 276 3572
rect 270 3567 276 3568
rect 414 3572 420 3573
rect 414 3568 415 3572
rect 419 3568 420 3572
rect 414 3567 420 3568
rect 574 3572 580 3573
rect 574 3568 575 3572
rect 579 3568 580 3572
rect 574 3567 580 3568
rect 734 3572 740 3573
rect 734 3568 735 3572
rect 739 3568 740 3572
rect 734 3567 740 3568
rect 894 3572 900 3573
rect 894 3568 895 3572
rect 899 3568 900 3572
rect 894 3567 900 3568
rect 1054 3572 1060 3573
rect 1054 3568 1055 3572
rect 1059 3568 1060 3572
rect 1054 3567 1060 3568
rect 1214 3572 1220 3573
rect 1214 3568 1215 3572
rect 1219 3568 1220 3572
rect 1214 3567 1220 3568
rect 1374 3572 1380 3573
rect 1374 3568 1375 3572
rect 1379 3568 1380 3572
rect 1374 3567 1380 3568
rect 1542 3572 1548 3573
rect 1542 3568 1543 3572
rect 1547 3568 1548 3572
rect 1542 3567 1548 3568
rect 2006 3569 2012 3570
rect 110 3564 116 3565
rect 2006 3565 2007 3569
rect 2011 3565 2012 3569
rect 2006 3564 2012 3565
rect 270 3553 276 3554
rect 110 3552 116 3553
rect 110 3548 111 3552
rect 115 3548 116 3552
rect 270 3549 271 3553
rect 275 3549 276 3553
rect 270 3548 276 3549
rect 414 3553 420 3554
rect 414 3549 415 3553
rect 419 3549 420 3553
rect 414 3548 420 3549
rect 574 3553 580 3554
rect 574 3549 575 3553
rect 579 3549 580 3553
rect 574 3548 580 3549
rect 734 3553 740 3554
rect 734 3549 735 3553
rect 739 3549 740 3553
rect 734 3548 740 3549
rect 894 3553 900 3554
rect 894 3549 895 3553
rect 899 3549 900 3553
rect 894 3548 900 3549
rect 1054 3553 1060 3554
rect 1054 3549 1055 3553
rect 1059 3549 1060 3553
rect 1054 3548 1060 3549
rect 1214 3553 1220 3554
rect 1214 3549 1215 3553
rect 1219 3549 1220 3553
rect 1214 3548 1220 3549
rect 1374 3553 1380 3554
rect 1374 3549 1375 3553
rect 1379 3549 1380 3553
rect 1374 3548 1380 3549
rect 1542 3553 1548 3554
rect 1542 3549 1543 3553
rect 1547 3549 1548 3553
rect 1542 3548 1548 3549
rect 2006 3552 2012 3553
rect 2006 3548 2007 3552
rect 2011 3548 2012 3552
rect 110 3547 116 3548
rect 2006 3547 2012 3548
rect 2046 3516 2052 3517
rect 3942 3516 3948 3517
rect 2046 3512 2047 3516
rect 2051 3512 2052 3516
rect 2046 3511 2052 3512
rect 2286 3515 2292 3516
rect 2286 3511 2287 3515
rect 2291 3511 2292 3515
rect 2286 3510 2292 3511
rect 2382 3515 2388 3516
rect 2382 3511 2383 3515
rect 2387 3511 2388 3515
rect 2382 3510 2388 3511
rect 2478 3515 2484 3516
rect 2478 3511 2479 3515
rect 2483 3511 2484 3515
rect 2478 3510 2484 3511
rect 2574 3515 2580 3516
rect 2574 3511 2575 3515
rect 2579 3511 2580 3515
rect 2574 3510 2580 3511
rect 2670 3515 2676 3516
rect 2670 3511 2671 3515
rect 2675 3511 2676 3515
rect 2670 3510 2676 3511
rect 2766 3515 2772 3516
rect 2766 3511 2767 3515
rect 2771 3511 2772 3515
rect 2766 3510 2772 3511
rect 2870 3515 2876 3516
rect 2870 3511 2871 3515
rect 2875 3511 2876 3515
rect 2870 3510 2876 3511
rect 2982 3515 2988 3516
rect 2982 3511 2983 3515
rect 2987 3511 2988 3515
rect 2982 3510 2988 3511
rect 3102 3515 3108 3516
rect 3102 3511 3103 3515
rect 3107 3511 3108 3515
rect 3102 3510 3108 3511
rect 3222 3515 3228 3516
rect 3222 3511 3223 3515
rect 3227 3511 3228 3515
rect 3222 3510 3228 3511
rect 3350 3515 3356 3516
rect 3350 3511 3351 3515
rect 3355 3511 3356 3515
rect 3350 3510 3356 3511
rect 3486 3515 3492 3516
rect 3486 3511 3487 3515
rect 3491 3511 3492 3515
rect 3942 3512 3943 3516
rect 3947 3512 3948 3516
rect 3942 3511 3948 3512
rect 3486 3510 3492 3511
rect 2046 3499 2052 3500
rect 2046 3495 2047 3499
rect 2051 3495 2052 3499
rect 3942 3499 3948 3500
rect 2046 3494 2052 3495
rect 2286 3496 2292 3497
rect 110 3492 116 3493
rect 2006 3492 2012 3493
rect 110 3488 111 3492
rect 115 3488 116 3492
rect 110 3487 116 3488
rect 158 3491 164 3492
rect 158 3487 159 3491
rect 163 3487 164 3491
rect 158 3486 164 3487
rect 286 3491 292 3492
rect 286 3487 287 3491
rect 291 3487 292 3491
rect 286 3486 292 3487
rect 422 3491 428 3492
rect 422 3487 423 3491
rect 427 3487 428 3491
rect 422 3486 428 3487
rect 558 3491 564 3492
rect 558 3487 559 3491
rect 563 3487 564 3491
rect 558 3486 564 3487
rect 694 3491 700 3492
rect 694 3487 695 3491
rect 699 3487 700 3491
rect 694 3486 700 3487
rect 830 3491 836 3492
rect 830 3487 831 3491
rect 835 3487 836 3491
rect 830 3486 836 3487
rect 966 3491 972 3492
rect 966 3487 967 3491
rect 971 3487 972 3491
rect 966 3486 972 3487
rect 1094 3491 1100 3492
rect 1094 3487 1095 3491
rect 1099 3487 1100 3491
rect 1094 3486 1100 3487
rect 1230 3491 1236 3492
rect 1230 3487 1231 3491
rect 1235 3487 1236 3491
rect 1230 3486 1236 3487
rect 1366 3491 1372 3492
rect 1366 3487 1367 3491
rect 1371 3487 1372 3491
rect 2006 3488 2007 3492
rect 2011 3488 2012 3492
rect 2286 3492 2287 3496
rect 2291 3492 2292 3496
rect 2286 3491 2292 3492
rect 2382 3496 2388 3497
rect 2382 3492 2383 3496
rect 2387 3492 2388 3496
rect 2382 3491 2388 3492
rect 2478 3496 2484 3497
rect 2478 3492 2479 3496
rect 2483 3492 2484 3496
rect 2478 3491 2484 3492
rect 2574 3496 2580 3497
rect 2574 3492 2575 3496
rect 2579 3492 2580 3496
rect 2574 3491 2580 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2766 3496 2772 3497
rect 2766 3492 2767 3496
rect 2771 3492 2772 3496
rect 2766 3491 2772 3492
rect 2870 3496 2876 3497
rect 2870 3492 2871 3496
rect 2875 3492 2876 3496
rect 2870 3491 2876 3492
rect 2982 3496 2988 3497
rect 2982 3492 2983 3496
rect 2987 3492 2988 3496
rect 2982 3491 2988 3492
rect 3102 3496 3108 3497
rect 3102 3492 3103 3496
rect 3107 3492 3108 3496
rect 3102 3491 3108 3492
rect 3222 3496 3228 3497
rect 3222 3492 3223 3496
rect 3227 3492 3228 3496
rect 3222 3491 3228 3492
rect 3350 3496 3356 3497
rect 3350 3492 3351 3496
rect 3355 3492 3356 3496
rect 3350 3491 3356 3492
rect 3486 3496 3492 3497
rect 3486 3492 3487 3496
rect 3491 3492 3492 3496
rect 3942 3495 3943 3499
rect 3947 3495 3948 3499
rect 3942 3494 3948 3495
rect 3486 3491 3492 3492
rect 2006 3487 2012 3488
rect 1366 3486 1372 3487
rect 110 3475 116 3476
rect 110 3471 111 3475
rect 115 3471 116 3475
rect 2006 3475 2012 3476
rect 110 3470 116 3471
rect 158 3472 164 3473
rect 158 3468 159 3472
rect 163 3468 164 3472
rect 158 3467 164 3468
rect 286 3472 292 3473
rect 286 3468 287 3472
rect 291 3468 292 3472
rect 286 3467 292 3468
rect 422 3472 428 3473
rect 422 3468 423 3472
rect 427 3468 428 3472
rect 422 3467 428 3468
rect 558 3472 564 3473
rect 558 3468 559 3472
rect 563 3468 564 3472
rect 558 3467 564 3468
rect 694 3472 700 3473
rect 694 3468 695 3472
rect 699 3468 700 3472
rect 694 3467 700 3468
rect 830 3472 836 3473
rect 830 3468 831 3472
rect 835 3468 836 3472
rect 830 3467 836 3468
rect 966 3472 972 3473
rect 966 3468 967 3472
rect 971 3468 972 3472
rect 966 3467 972 3468
rect 1094 3472 1100 3473
rect 1094 3468 1095 3472
rect 1099 3468 1100 3472
rect 1094 3467 1100 3468
rect 1230 3472 1236 3473
rect 1230 3468 1231 3472
rect 1235 3468 1236 3472
rect 1230 3467 1236 3468
rect 1366 3472 1372 3473
rect 1366 3468 1367 3472
rect 1371 3468 1372 3472
rect 2006 3471 2007 3475
rect 2011 3471 2012 3475
rect 2006 3470 2012 3471
rect 1366 3467 1372 3468
rect 2486 3436 2492 3437
rect 2046 3433 2052 3434
rect 2046 3429 2047 3433
rect 2051 3429 2052 3433
rect 2486 3432 2487 3436
rect 2491 3432 2492 3436
rect 2486 3431 2492 3432
rect 2582 3436 2588 3437
rect 2582 3432 2583 3436
rect 2587 3432 2588 3436
rect 2582 3431 2588 3432
rect 2678 3436 2684 3437
rect 2678 3432 2679 3436
rect 2683 3432 2684 3436
rect 2678 3431 2684 3432
rect 2782 3436 2788 3437
rect 2782 3432 2783 3436
rect 2787 3432 2788 3436
rect 2782 3431 2788 3432
rect 2894 3436 2900 3437
rect 2894 3432 2895 3436
rect 2899 3432 2900 3436
rect 2894 3431 2900 3432
rect 3014 3436 3020 3437
rect 3014 3432 3015 3436
rect 3019 3432 3020 3436
rect 3014 3431 3020 3432
rect 3142 3436 3148 3437
rect 3142 3432 3143 3436
rect 3147 3432 3148 3436
rect 3142 3431 3148 3432
rect 3270 3436 3276 3437
rect 3270 3432 3271 3436
rect 3275 3432 3276 3436
rect 3270 3431 3276 3432
rect 3406 3436 3412 3437
rect 3406 3432 3407 3436
rect 3411 3432 3412 3436
rect 3406 3431 3412 3432
rect 3942 3433 3948 3434
rect 2046 3428 2052 3429
rect 3942 3429 3943 3433
rect 3947 3429 3948 3433
rect 3942 3428 3948 3429
rect 2486 3417 2492 3418
rect 2046 3416 2052 3417
rect 2046 3412 2047 3416
rect 2051 3412 2052 3416
rect 2486 3413 2487 3417
rect 2491 3413 2492 3417
rect 2486 3412 2492 3413
rect 2582 3417 2588 3418
rect 2582 3413 2583 3417
rect 2587 3413 2588 3417
rect 2582 3412 2588 3413
rect 2678 3417 2684 3418
rect 2678 3413 2679 3417
rect 2683 3413 2684 3417
rect 2678 3412 2684 3413
rect 2782 3417 2788 3418
rect 2782 3413 2783 3417
rect 2787 3413 2788 3417
rect 2782 3412 2788 3413
rect 2894 3417 2900 3418
rect 2894 3413 2895 3417
rect 2899 3413 2900 3417
rect 2894 3412 2900 3413
rect 3014 3417 3020 3418
rect 3014 3413 3015 3417
rect 3019 3413 3020 3417
rect 3014 3412 3020 3413
rect 3142 3417 3148 3418
rect 3142 3413 3143 3417
rect 3147 3413 3148 3417
rect 3142 3412 3148 3413
rect 3270 3417 3276 3418
rect 3270 3413 3271 3417
rect 3275 3413 3276 3417
rect 3270 3412 3276 3413
rect 3406 3417 3412 3418
rect 3406 3413 3407 3417
rect 3411 3413 3412 3417
rect 3406 3412 3412 3413
rect 3942 3416 3948 3417
rect 3942 3412 3943 3416
rect 3947 3412 3948 3416
rect 2046 3411 2052 3412
rect 3942 3411 3948 3412
rect 134 3404 140 3405
rect 110 3401 116 3402
rect 110 3397 111 3401
rect 115 3397 116 3401
rect 134 3400 135 3404
rect 139 3400 140 3404
rect 134 3399 140 3400
rect 246 3404 252 3405
rect 246 3400 247 3404
rect 251 3400 252 3404
rect 246 3399 252 3400
rect 382 3404 388 3405
rect 382 3400 383 3404
rect 387 3400 388 3404
rect 382 3399 388 3400
rect 526 3404 532 3405
rect 526 3400 527 3404
rect 531 3400 532 3404
rect 526 3399 532 3400
rect 670 3404 676 3405
rect 670 3400 671 3404
rect 675 3400 676 3404
rect 670 3399 676 3400
rect 814 3404 820 3405
rect 814 3400 815 3404
rect 819 3400 820 3404
rect 814 3399 820 3400
rect 966 3404 972 3405
rect 966 3400 967 3404
rect 971 3400 972 3404
rect 966 3399 972 3400
rect 1118 3404 1124 3405
rect 1118 3400 1119 3404
rect 1123 3400 1124 3404
rect 1118 3399 1124 3400
rect 1270 3404 1276 3405
rect 1270 3400 1271 3404
rect 1275 3400 1276 3404
rect 1270 3399 1276 3400
rect 2006 3401 2012 3402
rect 110 3396 116 3397
rect 2006 3397 2007 3401
rect 2011 3397 2012 3401
rect 2006 3396 2012 3397
rect 134 3385 140 3386
rect 110 3384 116 3385
rect 110 3380 111 3384
rect 115 3380 116 3384
rect 134 3381 135 3385
rect 139 3381 140 3385
rect 134 3380 140 3381
rect 246 3385 252 3386
rect 246 3381 247 3385
rect 251 3381 252 3385
rect 246 3380 252 3381
rect 382 3385 388 3386
rect 382 3381 383 3385
rect 387 3381 388 3385
rect 382 3380 388 3381
rect 526 3385 532 3386
rect 526 3381 527 3385
rect 531 3381 532 3385
rect 526 3380 532 3381
rect 670 3385 676 3386
rect 670 3381 671 3385
rect 675 3381 676 3385
rect 670 3380 676 3381
rect 814 3385 820 3386
rect 814 3381 815 3385
rect 819 3381 820 3385
rect 814 3380 820 3381
rect 966 3385 972 3386
rect 966 3381 967 3385
rect 971 3381 972 3385
rect 966 3380 972 3381
rect 1118 3385 1124 3386
rect 1118 3381 1119 3385
rect 1123 3381 1124 3385
rect 1118 3380 1124 3381
rect 1270 3385 1276 3386
rect 1270 3381 1271 3385
rect 1275 3381 1276 3385
rect 1270 3380 1276 3381
rect 2006 3384 2012 3385
rect 2006 3380 2007 3384
rect 2011 3380 2012 3384
rect 110 3379 116 3380
rect 2006 3379 2012 3380
rect 2046 3356 2052 3357
rect 3942 3356 3948 3357
rect 2046 3352 2047 3356
rect 2051 3352 2052 3356
rect 2046 3351 2052 3352
rect 2350 3355 2356 3356
rect 2350 3351 2351 3355
rect 2355 3351 2356 3355
rect 2350 3350 2356 3351
rect 2478 3355 2484 3356
rect 2478 3351 2479 3355
rect 2483 3351 2484 3355
rect 2478 3350 2484 3351
rect 2614 3355 2620 3356
rect 2614 3351 2615 3355
rect 2619 3351 2620 3355
rect 2614 3350 2620 3351
rect 2750 3355 2756 3356
rect 2750 3351 2751 3355
rect 2755 3351 2756 3355
rect 2750 3350 2756 3351
rect 2886 3355 2892 3356
rect 2886 3351 2887 3355
rect 2891 3351 2892 3355
rect 2886 3350 2892 3351
rect 3022 3355 3028 3356
rect 3022 3351 3023 3355
rect 3027 3351 3028 3355
rect 3022 3350 3028 3351
rect 3158 3355 3164 3356
rect 3158 3351 3159 3355
rect 3163 3351 3164 3355
rect 3158 3350 3164 3351
rect 3302 3355 3308 3356
rect 3302 3351 3303 3355
rect 3307 3351 3308 3355
rect 3942 3352 3943 3356
rect 3947 3352 3948 3356
rect 3942 3351 3948 3352
rect 3302 3350 3308 3351
rect 2046 3339 2052 3340
rect 2046 3335 2047 3339
rect 2051 3335 2052 3339
rect 3942 3339 3948 3340
rect 2046 3334 2052 3335
rect 2350 3336 2356 3337
rect 2350 3332 2351 3336
rect 2355 3332 2356 3336
rect 2350 3331 2356 3332
rect 2478 3336 2484 3337
rect 2478 3332 2479 3336
rect 2483 3332 2484 3336
rect 2478 3331 2484 3332
rect 2614 3336 2620 3337
rect 2614 3332 2615 3336
rect 2619 3332 2620 3336
rect 2614 3331 2620 3332
rect 2750 3336 2756 3337
rect 2750 3332 2751 3336
rect 2755 3332 2756 3336
rect 2750 3331 2756 3332
rect 2886 3336 2892 3337
rect 2886 3332 2887 3336
rect 2891 3332 2892 3336
rect 2886 3331 2892 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3158 3336 3164 3337
rect 3158 3332 3159 3336
rect 3163 3332 3164 3336
rect 3158 3331 3164 3332
rect 3302 3336 3308 3337
rect 3302 3332 3303 3336
rect 3307 3332 3308 3336
rect 3942 3335 3943 3339
rect 3947 3335 3948 3339
rect 3942 3334 3948 3335
rect 3302 3331 3308 3332
rect 110 3324 116 3325
rect 2006 3324 2012 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 134 3323 140 3324
rect 134 3319 135 3323
rect 139 3319 140 3323
rect 134 3318 140 3319
rect 262 3323 268 3324
rect 262 3319 263 3323
rect 267 3319 268 3323
rect 262 3318 268 3319
rect 430 3323 436 3324
rect 430 3319 431 3323
rect 435 3319 436 3323
rect 430 3318 436 3319
rect 598 3323 604 3324
rect 598 3319 599 3323
rect 603 3319 604 3323
rect 598 3318 604 3319
rect 766 3323 772 3324
rect 766 3319 767 3323
rect 771 3319 772 3323
rect 766 3318 772 3319
rect 926 3323 932 3324
rect 926 3319 927 3323
rect 931 3319 932 3323
rect 926 3318 932 3319
rect 1086 3323 1092 3324
rect 1086 3319 1087 3323
rect 1091 3319 1092 3323
rect 1086 3318 1092 3319
rect 1238 3323 1244 3324
rect 1238 3319 1239 3323
rect 1243 3319 1244 3323
rect 1238 3318 1244 3319
rect 1390 3323 1396 3324
rect 1390 3319 1391 3323
rect 1395 3319 1396 3323
rect 1390 3318 1396 3319
rect 1550 3323 1556 3324
rect 1550 3319 1551 3323
rect 1555 3319 1556 3323
rect 2006 3320 2007 3324
rect 2011 3320 2012 3324
rect 2006 3319 2012 3320
rect 1550 3318 1556 3319
rect 110 3307 116 3308
rect 110 3303 111 3307
rect 115 3303 116 3307
rect 2006 3307 2012 3308
rect 110 3302 116 3303
rect 134 3304 140 3305
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 262 3304 268 3305
rect 262 3300 263 3304
rect 267 3300 268 3304
rect 262 3299 268 3300
rect 430 3304 436 3305
rect 430 3300 431 3304
rect 435 3300 436 3304
rect 430 3299 436 3300
rect 598 3304 604 3305
rect 598 3300 599 3304
rect 603 3300 604 3304
rect 598 3299 604 3300
rect 766 3304 772 3305
rect 766 3300 767 3304
rect 771 3300 772 3304
rect 766 3299 772 3300
rect 926 3304 932 3305
rect 926 3300 927 3304
rect 931 3300 932 3304
rect 926 3299 932 3300
rect 1086 3304 1092 3305
rect 1086 3300 1087 3304
rect 1091 3300 1092 3304
rect 1086 3299 1092 3300
rect 1238 3304 1244 3305
rect 1238 3300 1239 3304
rect 1243 3300 1244 3304
rect 1238 3299 1244 3300
rect 1390 3304 1396 3305
rect 1390 3300 1391 3304
rect 1395 3300 1396 3304
rect 1390 3299 1396 3300
rect 1550 3304 1556 3305
rect 1550 3300 1551 3304
rect 1555 3300 1556 3304
rect 2006 3303 2007 3307
rect 2011 3303 2012 3307
rect 2006 3302 2012 3303
rect 1550 3299 1556 3300
rect 2126 3272 2132 3273
rect 2046 3269 2052 3270
rect 2046 3265 2047 3269
rect 2051 3265 2052 3269
rect 2126 3268 2127 3272
rect 2131 3268 2132 3272
rect 2126 3267 2132 3268
rect 2294 3272 2300 3273
rect 2294 3268 2295 3272
rect 2299 3268 2300 3272
rect 2294 3267 2300 3268
rect 2454 3272 2460 3273
rect 2454 3268 2455 3272
rect 2459 3268 2460 3272
rect 2454 3267 2460 3268
rect 2614 3272 2620 3273
rect 2614 3268 2615 3272
rect 2619 3268 2620 3272
rect 2614 3267 2620 3268
rect 2774 3272 2780 3273
rect 2774 3268 2775 3272
rect 2779 3268 2780 3272
rect 2774 3267 2780 3268
rect 2934 3272 2940 3273
rect 2934 3268 2935 3272
rect 2939 3268 2940 3272
rect 2934 3267 2940 3268
rect 3094 3272 3100 3273
rect 3094 3268 3095 3272
rect 3099 3268 3100 3272
rect 3094 3267 3100 3268
rect 3262 3272 3268 3273
rect 3262 3268 3263 3272
rect 3267 3268 3268 3272
rect 3262 3267 3268 3268
rect 3942 3269 3948 3270
rect 2046 3264 2052 3265
rect 3942 3265 3943 3269
rect 3947 3265 3948 3269
rect 3942 3264 3948 3265
rect 2126 3253 2132 3254
rect 2046 3252 2052 3253
rect 2046 3248 2047 3252
rect 2051 3248 2052 3252
rect 2126 3249 2127 3253
rect 2131 3249 2132 3253
rect 2126 3248 2132 3249
rect 2294 3253 2300 3254
rect 2294 3249 2295 3253
rect 2299 3249 2300 3253
rect 2294 3248 2300 3249
rect 2454 3253 2460 3254
rect 2454 3249 2455 3253
rect 2459 3249 2460 3253
rect 2454 3248 2460 3249
rect 2614 3253 2620 3254
rect 2614 3249 2615 3253
rect 2619 3249 2620 3253
rect 2614 3248 2620 3249
rect 2774 3253 2780 3254
rect 2774 3249 2775 3253
rect 2779 3249 2780 3253
rect 2774 3248 2780 3249
rect 2934 3253 2940 3254
rect 2934 3249 2935 3253
rect 2939 3249 2940 3253
rect 2934 3248 2940 3249
rect 3094 3253 3100 3254
rect 3094 3249 3095 3253
rect 3099 3249 3100 3253
rect 3094 3248 3100 3249
rect 3262 3253 3268 3254
rect 3262 3249 3263 3253
rect 3267 3249 3268 3253
rect 3262 3248 3268 3249
rect 3942 3252 3948 3253
rect 3942 3248 3943 3252
rect 3947 3248 3948 3252
rect 2046 3247 2052 3248
rect 3942 3247 3948 3248
rect 142 3236 148 3237
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 142 3232 143 3236
rect 147 3232 148 3236
rect 142 3231 148 3232
rect 294 3236 300 3237
rect 294 3232 295 3236
rect 299 3232 300 3236
rect 294 3231 300 3232
rect 454 3236 460 3237
rect 454 3232 455 3236
rect 459 3232 460 3236
rect 454 3231 460 3232
rect 622 3236 628 3237
rect 622 3232 623 3236
rect 627 3232 628 3236
rect 622 3231 628 3232
rect 790 3236 796 3237
rect 790 3232 791 3236
rect 795 3232 796 3236
rect 790 3231 796 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 958 3231 964 3232
rect 1126 3236 1132 3237
rect 1126 3232 1127 3236
rect 1131 3232 1132 3236
rect 1126 3231 1132 3232
rect 1302 3236 1308 3237
rect 1302 3232 1303 3236
rect 1307 3232 1308 3236
rect 1302 3231 1308 3232
rect 1478 3236 1484 3237
rect 1478 3232 1479 3236
rect 1483 3232 1484 3236
rect 1478 3231 1484 3232
rect 2006 3233 2012 3234
rect 110 3228 116 3229
rect 2006 3229 2007 3233
rect 2011 3229 2012 3233
rect 2006 3228 2012 3229
rect 142 3217 148 3218
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 142 3213 143 3217
rect 147 3213 148 3217
rect 142 3212 148 3213
rect 294 3217 300 3218
rect 294 3213 295 3217
rect 299 3213 300 3217
rect 294 3212 300 3213
rect 454 3217 460 3218
rect 454 3213 455 3217
rect 459 3213 460 3217
rect 454 3212 460 3213
rect 622 3217 628 3218
rect 622 3213 623 3217
rect 627 3213 628 3217
rect 622 3212 628 3213
rect 790 3217 796 3218
rect 790 3213 791 3217
rect 795 3213 796 3217
rect 790 3212 796 3213
rect 958 3217 964 3218
rect 958 3213 959 3217
rect 963 3213 964 3217
rect 958 3212 964 3213
rect 1126 3217 1132 3218
rect 1126 3213 1127 3217
rect 1131 3213 1132 3217
rect 1126 3212 1132 3213
rect 1302 3217 1308 3218
rect 1302 3213 1303 3217
rect 1307 3213 1308 3217
rect 1302 3212 1308 3213
rect 1478 3217 1484 3218
rect 1478 3213 1479 3217
rect 1483 3213 1484 3217
rect 1478 3212 1484 3213
rect 2006 3216 2012 3217
rect 2006 3212 2007 3216
rect 2011 3212 2012 3216
rect 110 3211 116 3212
rect 2006 3211 2012 3212
rect 2046 3200 2052 3201
rect 3942 3200 3948 3201
rect 2046 3196 2047 3200
rect 2051 3196 2052 3200
rect 2046 3195 2052 3196
rect 2070 3199 2076 3200
rect 2070 3195 2071 3199
rect 2075 3195 2076 3199
rect 2070 3194 2076 3195
rect 2206 3199 2212 3200
rect 2206 3195 2207 3199
rect 2211 3195 2212 3199
rect 2206 3194 2212 3195
rect 2374 3199 2380 3200
rect 2374 3195 2375 3199
rect 2379 3195 2380 3199
rect 2374 3194 2380 3195
rect 2542 3199 2548 3200
rect 2542 3195 2543 3199
rect 2547 3195 2548 3199
rect 2542 3194 2548 3195
rect 2702 3199 2708 3200
rect 2702 3195 2703 3199
rect 2707 3195 2708 3199
rect 2702 3194 2708 3195
rect 2862 3199 2868 3200
rect 2862 3195 2863 3199
rect 2867 3195 2868 3199
rect 2862 3194 2868 3195
rect 3014 3199 3020 3200
rect 3014 3195 3015 3199
rect 3019 3195 3020 3199
rect 3014 3194 3020 3195
rect 3166 3199 3172 3200
rect 3166 3195 3167 3199
rect 3171 3195 3172 3199
rect 3166 3194 3172 3195
rect 3326 3199 3332 3200
rect 3326 3195 3327 3199
rect 3331 3195 3332 3199
rect 3942 3196 3943 3200
rect 3947 3196 3948 3200
rect 3942 3195 3948 3196
rect 3326 3194 3332 3195
rect 2046 3183 2052 3184
rect 2046 3179 2047 3183
rect 2051 3179 2052 3183
rect 3942 3183 3948 3184
rect 2046 3178 2052 3179
rect 2070 3180 2076 3181
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2206 3180 2212 3181
rect 2206 3176 2207 3180
rect 2211 3176 2212 3180
rect 2206 3175 2212 3176
rect 2374 3180 2380 3181
rect 2374 3176 2375 3180
rect 2379 3176 2380 3180
rect 2374 3175 2380 3176
rect 2542 3180 2548 3181
rect 2542 3176 2543 3180
rect 2547 3176 2548 3180
rect 2542 3175 2548 3176
rect 2702 3180 2708 3181
rect 2702 3176 2703 3180
rect 2707 3176 2708 3180
rect 2702 3175 2708 3176
rect 2862 3180 2868 3181
rect 2862 3176 2863 3180
rect 2867 3176 2868 3180
rect 2862 3175 2868 3176
rect 3014 3180 3020 3181
rect 3014 3176 3015 3180
rect 3019 3176 3020 3180
rect 3014 3175 3020 3176
rect 3166 3180 3172 3181
rect 3166 3176 3167 3180
rect 3171 3176 3172 3180
rect 3166 3175 3172 3176
rect 3326 3180 3332 3181
rect 3326 3176 3327 3180
rect 3331 3176 3332 3180
rect 3942 3179 3943 3183
rect 3947 3179 3948 3183
rect 3942 3178 3948 3179
rect 3326 3175 3332 3176
rect 110 3164 116 3165
rect 2006 3164 2012 3165
rect 110 3160 111 3164
rect 115 3160 116 3164
rect 110 3159 116 3160
rect 294 3163 300 3164
rect 294 3159 295 3163
rect 299 3159 300 3163
rect 294 3158 300 3159
rect 430 3163 436 3164
rect 430 3159 431 3163
rect 435 3159 436 3163
rect 430 3158 436 3159
rect 566 3163 572 3164
rect 566 3159 567 3163
rect 571 3159 572 3163
rect 566 3158 572 3159
rect 702 3163 708 3164
rect 702 3159 703 3163
rect 707 3159 708 3163
rect 702 3158 708 3159
rect 854 3163 860 3164
rect 854 3159 855 3163
rect 859 3159 860 3163
rect 854 3158 860 3159
rect 1030 3163 1036 3164
rect 1030 3159 1031 3163
rect 1035 3159 1036 3163
rect 1030 3158 1036 3159
rect 1230 3163 1236 3164
rect 1230 3159 1231 3163
rect 1235 3159 1236 3163
rect 1230 3158 1236 3159
rect 1454 3163 1460 3164
rect 1454 3159 1455 3163
rect 1459 3159 1460 3163
rect 1454 3158 1460 3159
rect 1686 3163 1692 3164
rect 1686 3159 1687 3163
rect 1691 3159 1692 3163
rect 1686 3158 1692 3159
rect 1902 3163 1908 3164
rect 1902 3159 1903 3163
rect 1907 3159 1908 3163
rect 2006 3160 2007 3164
rect 2011 3160 2012 3164
rect 2006 3159 2012 3160
rect 1902 3158 1908 3159
rect 110 3147 116 3148
rect 110 3143 111 3147
rect 115 3143 116 3147
rect 2006 3147 2012 3148
rect 110 3142 116 3143
rect 294 3144 300 3145
rect 294 3140 295 3144
rect 299 3140 300 3144
rect 294 3139 300 3140
rect 430 3144 436 3145
rect 430 3140 431 3144
rect 435 3140 436 3144
rect 430 3139 436 3140
rect 566 3144 572 3145
rect 566 3140 567 3144
rect 571 3140 572 3144
rect 566 3139 572 3140
rect 702 3144 708 3145
rect 702 3140 703 3144
rect 707 3140 708 3144
rect 702 3139 708 3140
rect 854 3144 860 3145
rect 854 3140 855 3144
rect 859 3140 860 3144
rect 854 3139 860 3140
rect 1030 3144 1036 3145
rect 1030 3140 1031 3144
rect 1035 3140 1036 3144
rect 1030 3139 1036 3140
rect 1230 3144 1236 3145
rect 1230 3140 1231 3144
rect 1235 3140 1236 3144
rect 1230 3139 1236 3140
rect 1454 3144 1460 3145
rect 1454 3140 1455 3144
rect 1459 3140 1460 3144
rect 1454 3139 1460 3140
rect 1686 3144 1692 3145
rect 1686 3140 1687 3144
rect 1691 3140 1692 3144
rect 1686 3139 1692 3140
rect 1902 3144 1908 3145
rect 1902 3140 1903 3144
rect 1907 3140 1908 3144
rect 2006 3143 2007 3147
rect 2011 3143 2012 3147
rect 2006 3142 2012 3143
rect 1902 3139 1908 3140
rect 2070 3116 2076 3117
rect 2046 3113 2052 3114
rect 2046 3109 2047 3113
rect 2051 3109 2052 3113
rect 2070 3112 2071 3116
rect 2075 3112 2076 3116
rect 2070 3111 2076 3112
rect 2342 3116 2348 3117
rect 2342 3112 2343 3116
rect 2347 3112 2348 3116
rect 2342 3111 2348 3112
rect 2630 3116 2636 3117
rect 2630 3112 2631 3116
rect 2635 3112 2636 3116
rect 2630 3111 2636 3112
rect 2902 3116 2908 3117
rect 2902 3112 2903 3116
rect 2907 3112 2908 3116
rect 2902 3111 2908 3112
rect 3174 3116 3180 3117
rect 3174 3112 3175 3116
rect 3179 3112 3180 3116
rect 3174 3111 3180 3112
rect 3446 3116 3452 3117
rect 3446 3112 3447 3116
rect 3451 3112 3452 3116
rect 3446 3111 3452 3112
rect 3942 3113 3948 3114
rect 2046 3108 2052 3109
rect 3942 3109 3943 3113
rect 3947 3109 3948 3113
rect 3942 3108 3948 3109
rect 2070 3097 2076 3098
rect 2046 3096 2052 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2070 3093 2071 3097
rect 2075 3093 2076 3097
rect 2070 3092 2076 3093
rect 2342 3097 2348 3098
rect 2342 3093 2343 3097
rect 2347 3093 2348 3097
rect 2342 3092 2348 3093
rect 2630 3097 2636 3098
rect 2630 3093 2631 3097
rect 2635 3093 2636 3097
rect 2630 3092 2636 3093
rect 2902 3097 2908 3098
rect 2902 3093 2903 3097
rect 2907 3093 2908 3097
rect 2902 3092 2908 3093
rect 3174 3097 3180 3098
rect 3174 3093 3175 3097
rect 3179 3093 3180 3097
rect 3174 3092 3180 3093
rect 3446 3097 3452 3098
rect 3446 3093 3447 3097
rect 3451 3093 3452 3097
rect 3446 3092 3452 3093
rect 3942 3096 3948 3097
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 2046 3091 2052 3092
rect 3942 3091 3948 3092
rect 310 3084 316 3085
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 310 3080 311 3084
rect 315 3080 316 3084
rect 310 3079 316 3080
rect 406 3084 412 3085
rect 406 3080 407 3084
rect 411 3080 412 3084
rect 406 3079 412 3080
rect 502 3084 508 3085
rect 502 3080 503 3084
rect 507 3080 508 3084
rect 502 3079 508 3080
rect 598 3084 604 3085
rect 598 3080 599 3084
rect 603 3080 604 3084
rect 598 3079 604 3080
rect 694 3084 700 3085
rect 694 3080 695 3084
rect 699 3080 700 3084
rect 694 3079 700 3080
rect 806 3084 812 3085
rect 806 3080 807 3084
rect 811 3080 812 3084
rect 806 3079 812 3080
rect 942 3084 948 3085
rect 942 3080 943 3084
rect 947 3080 948 3084
rect 942 3079 948 3080
rect 1086 3084 1092 3085
rect 1086 3080 1087 3084
rect 1091 3080 1092 3084
rect 1086 3079 1092 3080
rect 1246 3084 1252 3085
rect 1246 3080 1247 3084
rect 1251 3080 1252 3084
rect 1246 3079 1252 3080
rect 1406 3084 1412 3085
rect 1406 3080 1407 3084
rect 1411 3080 1412 3084
rect 1406 3079 1412 3080
rect 1574 3084 1580 3085
rect 1574 3080 1575 3084
rect 1579 3080 1580 3084
rect 1574 3079 1580 3080
rect 1750 3084 1756 3085
rect 1750 3080 1751 3084
rect 1755 3080 1756 3084
rect 1750 3079 1756 3080
rect 1902 3084 1908 3085
rect 1902 3080 1903 3084
rect 1907 3080 1908 3084
rect 1902 3079 1908 3080
rect 2006 3081 2012 3082
rect 110 3076 116 3077
rect 2006 3077 2007 3081
rect 2011 3077 2012 3081
rect 2006 3076 2012 3077
rect 310 3065 316 3066
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 310 3061 311 3065
rect 315 3061 316 3065
rect 310 3060 316 3061
rect 406 3065 412 3066
rect 406 3061 407 3065
rect 411 3061 412 3065
rect 406 3060 412 3061
rect 502 3065 508 3066
rect 502 3061 503 3065
rect 507 3061 508 3065
rect 502 3060 508 3061
rect 598 3065 604 3066
rect 598 3061 599 3065
rect 603 3061 604 3065
rect 598 3060 604 3061
rect 694 3065 700 3066
rect 694 3061 695 3065
rect 699 3061 700 3065
rect 694 3060 700 3061
rect 806 3065 812 3066
rect 806 3061 807 3065
rect 811 3061 812 3065
rect 806 3060 812 3061
rect 942 3065 948 3066
rect 942 3061 943 3065
rect 947 3061 948 3065
rect 942 3060 948 3061
rect 1086 3065 1092 3066
rect 1086 3061 1087 3065
rect 1091 3061 1092 3065
rect 1086 3060 1092 3061
rect 1246 3065 1252 3066
rect 1246 3061 1247 3065
rect 1251 3061 1252 3065
rect 1246 3060 1252 3061
rect 1406 3065 1412 3066
rect 1406 3061 1407 3065
rect 1411 3061 1412 3065
rect 1406 3060 1412 3061
rect 1574 3065 1580 3066
rect 1574 3061 1575 3065
rect 1579 3061 1580 3065
rect 1574 3060 1580 3061
rect 1750 3065 1756 3066
rect 1750 3061 1751 3065
rect 1755 3061 1756 3065
rect 1750 3060 1756 3061
rect 1902 3065 1908 3066
rect 1902 3061 1903 3065
rect 1907 3061 1908 3065
rect 1902 3060 1908 3061
rect 2006 3064 2012 3065
rect 2006 3060 2007 3064
rect 2011 3060 2012 3064
rect 110 3059 116 3060
rect 2006 3059 2012 3060
rect 2046 3040 2052 3041
rect 3942 3040 3948 3041
rect 2046 3036 2047 3040
rect 2051 3036 2052 3040
rect 2046 3035 2052 3036
rect 2486 3039 2492 3040
rect 2486 3035 2487 3039
rect 2491 3035 2492 3039
rect 2486 3034 2492 3035
rect 2614 3039 2620 3040
rect 2614 3035 2615 3039
rect 2619 3035 2620 3039
rect 2614 3034 2620 3035
rect 2742 3039 2748 3040
rect 2742 3035 2743 3039
rect 2747 3035 2748 3039
rect 2742 3034 2748 3035
rect 2862 3039 2868 3040
rect 2862 3035 2863 3039
rect 2867 3035 2868 3039
rect 2862 3034 2868 3035
rect 2982 3039 2988 3040
rect 2982 3035 2983 3039
rect 2987 3035 2988 3039
rect 2982 3034 2988 3035
rect 3102 3039 3108 3040
rect 3102 3035 3103 3039
rect 3107 3035 3108 3039
rect 3102 3034 3108 3035
rect 3214 3039 3220 3040
rect 3214 3035 3215 3039
rect 3219 3035 3220 3039
rect 3214 3034 3220 3035
rect 3326 3039 3332 3040
rect 3326 3035 3327 3039
rect 3331 3035 3332 3039
rect 3326 3034 3332 3035
rect 3430 3039 3436 3040
rect 3430 3035 3431 3039
rect 3435 3035 3436 3039
rect 3430 3034 3436 3035
rect 3534 3039 3540 3040
rect 3534 3035 3535 3039
rect 3539 3035 3540 3039
rect 3534 3034 3540 3035
rect 3638 3039 3644 3040
rect 3638 3035 3639 3039
rect 3643 3035 3644 3039
rect 3638 3034 3644 3035
rect 3742 3039 3748 3040
rect 3742 3035 3743 3039
rect 3747 3035 3748 3039
rect 3742 3034 3748 3035
rect 3838 3039 3844 3040
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3942 3036 3943 3040
rect 3947 3036 3948 3040
rect 3942 3035 3948 3036
rect 3838 3034 3844 3035
rect 2046 3023 2052 3024
rect 2046 3019 2047 3023
rect 2051 3019 2052 3023
rect 3942 3023 3948 3024
rect 2046 3018 2052 3019
rect 2486 3020 2492 3021
rect 2486 3016 2487 3020
rect 2491 3016 2492 3020
rect 2486 3015 2492 3016
rect 2614 3020 2620 3021
rect 2614 3016 2615 3020
rect 2619 3016 2620 3020
rect 2614 3015 2620 3016
rect 2742 3020 2748 3021
rect 2742 3016 2743 3020
rect 2747 3016 2748 3020
rect 2742 3015 2748 3016
rect 2862 3020 2868 3021
rect 2862 3016 2863 3020
rect 2867 3016 2868 3020
rect 2862 3015 2868 3016
rect 2982 3020 2988 3021
rect 2982 3016 2983 3020
rect 2987 3016 2988 3020
rect 2982 3015 2988 3016
rect 3102 3020 3108 3021
rect 3102 3016 3103 3020
rect 3107 3016 3108 3020
rect 3102 3015 3108 3016
rect 3214 3020 3220 3021
rect 3214 3016 3215 3020
rect 3219 3016 3220 3020
rect 3214 3015 3220 3016
rect 3326 3020 3332 3021
rect 3326 3016 3327 3020
rect 3331 3016 3332 3020
rect 3326 3015 3332 3016
rect 3430 3020 3436 3021
rect 3430 3016 3431 3020
rect 3435 3016 3436 3020
rect 3430 3015 3436 3016
rect 3534 3020 3540 3021
rect 3534 3016 3535 3020
rect 3539 3016 3540 3020
rect 3534 3015 3540 3016
rect 3638 3020 3644 3021
rect 3638 3016 3639 3020
rect 3643 3016 3644 3020
rect 3638 3015 3644 3016
rect 3742 3020 3748 3021
rect 3742 3016 3743 3020
rect 3747 3016 3748 3020
rect 3742 3015 3748 3016
rect 3838 3020 3844 3021
rect 3838 3016 3839 3020
rect 3843 3016 3844 3020
rect 3942 3019 3943 3023
rect 3947 3019 3948 3023
rect 3942 3018 3948 3019
rect 3838 3015 3844 3016
rect 110 3012 116 3013
rect 2006 3012 2012 3013
rect 110 3008 111 3012
rect 115 3008 116 3012
rect 110 3007 116 3008
rect 422 3011 428 3012
rect 422 3007 423 3011
rect 427 3007 428 3011
rect 422 3006 428 3007
rect 518 3011 524 3012
rect 518 3007 519 3011
rect 523 3007 524 3011
rect 518 3006 524 3007
rect 614 3011 620 3012
rect 614 3007 615 3011
rect 619 3007 620 3011
rect 614 3006 620 3007
rect 710 3011 716 3012
rect 710 3007 711 3011
rect 715 3007 716 3011
rect 710 3006 716 3007
rect 814 3011 820 3012
rect 814 3007 815 3011
rect 819 3007 820 3011
rect 814 3006 820 3007
rect 934 3011 940 3012
rect 934 3007 935 3011
rect 939 3007 940 3011
rect 934 3006 940 3007
rect 1054 3011 1060 3012
rect 1054 3007 1055 3011
rect 1059 3007 1060 3011
rect 1054 3006 1060 3007
rect 1182 3011 1188 3012
rect 1182 3007 1183 3011
rect 1187 3007 1188 3011
rect 1182 3006 1188 3007
rect 1310 3011 1316 3012
rect 1310 3007 1311 3011
rect 1315 3007 1316 3011
rect 1310 3006 1316 3007
rect 1430 3011 1436 3012
rect 1430 3007 1431 3011
rect 1435 3007 1436 3011
rect 1430 3006 1436 3007
rect 1550 3011 1556 3012
rect 1550 3007 1551 3011
rect 1555 3007 1556 3011
rect 1550 3006 1556 3007
rect 1670 3011 1676 3012
rect 1670 3007 1671 3011
rect 1675 3007 1676 3011
rect 1670 3006 1676 3007
rect 1798 3011 1804 3012
rect 1798 3007 1799 3011
rect 1803 3007 1804 3011
rect 1798 3006 1804 3007
rect 1902 3011 1908 3012
rect 1902 3007 1903 3011
rect 1907 3007 1908 3011
rect 2006 3008 2007 3012
rect 2011 3008 2012 3012
rect 2006 3007 2012 3008
rect 1902 3006 1908 3007
rect 110 2995 116 2996
rect 110 2991 111 2995
rect 115 2991 116 2995
rect 2006 2995 2012 2996
rect 110 2990 116 2991
rect 422 2992 428 2993
rect 422 2988 423 2992
rect 427 2988 428 2992
rect 422 2987 428 2988
rect 518 2992 524 2993
rect 518 2988 519 2992
rect 523 2988 524 2992
rect 518 2987 524 2988
rect 614 2992 620 2993
rect 614 2988 615 2992
rect 619 2988 620 2992
rect 614 2987 620 2988
rect 710 2992 716 2993
rect 710 2988 711 2992
rect 715 2988 716 2992
rect 710 2987 716 2988
rect 814 2992 820 2993
rect 814 2988 815 2992
rect 819 2988 820 2992
rect 814 2987 820 2988
rect 934 2992 940 2993
rect 934 2988 935 2992
rect 939 2988 940 2992
rect 934 2987 940 2988
rect 1054 2992 1060 2993
rect 1054 2988 1055 2992
rect 1059 2988 1060 2992
rect 1054 2987 1060 2988
rect 1182 2992 1188 2993
rect 1182 2988 1183 2992
rect 1187 2988 1188 2992
rect 1182 2987 1188 2988
rect 1310 2992 1316 2993
rect 1310 2988 1311 2992
rect 1315 2988 1316 2992
rect 1310 2987 1316 2988
rect 1430 2992 1436 2993
rect 1430 2988 1431 2992
rect 1435 2988 1436 2992
rect 1430 2987 1436 2988
rect 1550 2992 1556 2993
rect 1550 2988 1551 2992
rect 1555 2988 1556 2992
rect 1550 2987 1556 2988
rect 1670 2992 1676 2993
rect 1670 2988 1671 2992
rect 1675 2988 1676 2992
rect 1670 2987 1676 2988
rect 1798 2992 1804 2993
rect 1798 2988 1799 2992
rect 1803 2988 1804 2992
rect 1798 2987 1804 2988
rect 1902 2992 1908 2993
rect 1902 2988 1903 2992
rect 1907 2988 1908 2992
rect 2006 2991 2007 2995
rect 2011 2991 2012 2995
rect 2006 2990 2012 2991
rect 1902 2987 1908 2988
rect 2406 2956 2412 2957
rect 2046 2953 2052 2954
rect 2046 2949 2047 2953
rect 2051 2949 2052 2953
rect 2406 2952 2407 2956
rect 2411 2952 2412 2956
rect 2406 2951 2412 2952
rect 2574 2956 2580 2957
rect 2574 2952 2575 2956
rect 2579 2952 2580 2956
rect 2574 2951 2580 2952
rect 2766 2956 2772 2957
rect 2766 2952 2767 2956
rect 2771 2952 2772 2956
rect 2766 2951 2772 2952
rect 2966 2956 2972 2957
rect 2966 2952 2967 2956
rect 2971 2952 2972 2956
rect 2966 2951 2972 2952
rect 3182 2956 3188 2957
rect 3182 2952 3183 2956
rect 3187 2952 3188 2956
rect 3182 2951 3188 2952
rect 3398 2956 3404 2957
rect 3398 2952 3399 2956
rect 3403 2952 3404 2956
rect 3398 2951 3404 2952
rect 3622 2956 3628 2957
rect 3622 2952 3623 2956
rect 3627 2952 3628 2956
rect 3622 2951 3628 2952
rect 3838 2956 3844 2957
rect 3838 2952 3839 2956
rect 3843 2952 3844 2956
rect 3838 2951 3844 2952
rect 3942 2953 3948 2954
rect 2046 2948 2052 2949
rect 3942 2949 3943 2953
rect 3947 2949 3948 2953
rect 3942 2948 3948 2949
rect 2406 2937 2412 2938
rect 2046 2936 2052 2937
rect 2046 2932 2047 2936
rect 2051 2932 2052 2936
rect 2406 2933 2407 2937
rect 2411 2933 2412 2937
rect 2406 2932 2412 2933
rect 2574 2937 2580 2938
rect 2574 2933 2575 2937
rect 2579 2933 2580 2937
rect 2574 2932 2580 2933
rect 2766 2937 2772 2938
rect 2766 2933 2767 2937
rect 2771 2933 2772 2937
rect 2766 2932 2772 2933
rect 2966 2937 2972 2938
rect 2966 2933 2967 2937
rect 2971 2933 2972 2937
rect 2966 2932 2972 2933
rect 3182 2937 3188 2938
rect 3182 2933 3183 2937
rect 3187 2933 3188 2937
rect 3182 2932 3188 2933
rect 3398 2937 3404 2938
rect 3398 2933 3399 2937
rect 3403 2933 3404 2937
rect 3398 2932 3404 2933
rect 3622 2937 3628 2938
rect 3622 2933 3623 2937
rect 3627 2933 3628 2937
rect 3622 2932 3628 2933
rect 3838 2937 3844 2938
rect 3838 2933 3839 2937
rect 3843 2933 3844 2937
rect 3838 2932 3844 2933
rect 3942 2936 3948 2937
rect 3942 2932 3943 2936
rect 3947 2932 3948 2936
rect 2046 2931 2052 2932
rect 3942 2931 3948 2932
rect 1478 2908 1484 2909
rect 110 2905 116 2906
rect 110 2901 111 2905
rect 115 2901 116 2905
rect 1478 2904 1479 2908
rect 1483 2904 1484 2908
rect 1478 2903 1484 2904
rect 1574 2908 1580 2909
rect 1574 2904 1575 2908
rect 1579 2904 1580 2908
rect 1574 2903 1580 2904
rect 1670 2908 1676 2909
rect 1670 2904 1671 2908
rect 1675 2904 1676 2908
rect 1670 2903 1676 2904
rect 1766 2908 1772 2909
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1862 2908 1868 2909
rect 1862 2904 1863 2908
rect 1867 2904 1868 2908
rect 1862 2903 1868 2904
rect 2006 2905 2012 2906
rect 110 2900 116 2901
rect 2006 2901 2007 2905
rect 2011 2901 2012 2905
rect 2006 2900 2012 2901
rect 1478 2889 1484 2890
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 1478 2885 1479 2889
rect 1483 2885 1484 2889
rect 1478 2884 1484 2885
rect 1574 2889 1580 2890
rect 1574 2885 1575 2889
rect 1579 2885 1580 2889
rect 1574 2884 1580 2885
rect 1670 2889 1676 2890
rect 1670 2885 1671 2889
rect 1675 2885 1676 2889
rect 1670 2884 1676 2885
rect 1766 2889 1772 2890
rect 1766 2885 1767 2889
rect 1771 2885 1772 2889
rect 1766 2884 1772 2885
rect 1862 2889 1868 2890
rect 1862 2885 1863 2889
rect 1867 2885 1868 2889
rect 1862 2884 1868 2885
rect 2006 2888 2012 2889
rect 2006 2884 2007 2888
rect 2011 2884 2012 2888
rect 110 2883 116 2884
rect 2006 2883 2012 2884
rect 2046 2868 2052 2869
rect 3942 2868 3948 2869
rect 2046 2864 2047 2868
rect 2051 2864 2052 2868
rect 2046 2863 2052 2864
rect 2550 2867 2556 2868
rect 2550 2863 2551 2867
rect 2555 2863 2556 2867
rect 2550 2862 2556 2863
rect 2670 2867 2676 2868
rect 2670 2863 2671 2867
rect 2675 2863 2676 2867
rect 2670 2862 2676 2863
rect 2798 2867 2804 2868
rect 2798 2863 2799 2867
rect 2803 2863 2804 2867
rect 2798 2862 2804 2863
rect 2926 2867 2932 2868
rect 2926 2863 2927 2867
rect 2931 2863 2932 2867
rect 2926 2862 2932 2863
rect 3054 2867 3060 2868
rect 3054 2863 3055 2867
rect 3059 2863 3060 2867
rect 3054 2862 3060 2863
rect 3182 2867 3188 2868
rect 3182 2863 3183 2867
rect 3187 2863 3188 2867
rect 3182 2862 3188 2863
rect 3310 2867 3316 2868
rect 3310 2863 3311 2867
rect 3315 2863 3316 2867
rect 3310 2862 3316 2863
rect 3438 2867 3444 2868
rect 3438 2863 3439 2867
rect 3443 2863 3444 2867
rect 3438 2862 3444 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3942 2864 3943 2868
rect 3947 2864 3948 2868
rect 3942 2863 3948 2864
rect 3574 2862 3580 2863
rect 2046 2851 2052 2852
rect 2046 2847 2047 2851
rect 2051 2847 2052 2851
rect 3942 2851 3948 2852
rect 2046 2846 2052 2847
rect 2550 2848 2556 2849
rect 2550 2844 2551 2848
rect 2555 2844 2556 2848
rect 2550 2843 2556 2844
rect 2670 2848 2676 2849
rect 2670 2844 2671 2848
rect 2675 2844 2676 2848
rect 2670 2843 2676 2844
rect 2798 2848 2804 2849
rect 2798 2844 2799 2848
rect 2803 2844 2804 2848
rect 2798 2843 2804 2844
rect 2926 2848 2932 2849
rect 2926 2844 2927 2848
rect 2931 2844 2932 2848
rect 2926 2843 2932 2844
rect 3054 2848 3060 2849
rect 3054 2844 3055 2848
rect 3059 2844 3060 2848
rect 3054 2843 3060 2844
rect 3182 2848 3188 2849
rect 3182 2844 3183 2848
rect 3187 2844 3188 2848
rect 3182 2843 3188 2844
rect 3310 2848 3316 2849
rect 3310 2844 3311 2848
rect 3315 2844 3316 2848
rect 3310 2843 3316 2844
rect 3438 2848 3444 2849
rect 3438 2844 3439 2848
rect 3443 2844 3444 2848
rect 3438 2843 3444 2844
rect 3574 2848 3580 2849
rect 3574 2844 3575 2848
rect 3579 2844 3580 2848
rect 3942 2847 3943 2851
rect 3947 2847 3948 2851
rect 3942 2846 3948 2847
rect 3574 2843 3580 2844
rect 110 2828 116 2829
rect 2006 2828 2012 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 110 2823 116 2824
rect 278 2827 284 2828
rect 278 2823 279 2827
rect 283 2823 284 2827
rect 278 2822 284 2823
rect 446 2827 452 2828
rect 446 2823 447 2827
rect 451 2823 452 2827
rect 446 2822 452 2823
rect 630 2827 636 2828
rect 630 2823 631 2827
rect 635 2823 636 2827
rect 630 2822 636 2823
rect 814 2827 820 2828
rect 814 2823 815 2827
rect 819 2823 820 2827
rect 814 2822 820 2823
rect 998 2827 1004 2828
rect 998 2823 999 2827
rect 1003 2823 1004 2827
rect 998 2822 1004 2823
rect 1182 2827 1188 2828
rect 1182 2823 1183 2827
rect 1187 2823 1188 2827
rect 1182 2822 1188 2823
rect 1358 2827 1364 2828
rect 1358 2823 1359 2827
rect 1363 2823 1364 2827
rect 1358 2822 1364 2823
rect 1526 2827 1532 2828
rect 1526 2823 1527 2827
rect 1531 2823 1532 2827
rect 1526 2822 1532 2823
rect 1694 2827 1700 2828
rect 1694 2823 1695 2827
rect 1699 2823 1700 2827
rect 1694 2822 1700 2823
rect 1862 2827 1868 2828
rect 1862 2823 1863 2827
rect 1867 2823 1868 2827
rect 2006 2824 2007 2828
rect 2011 2824 2012 2828
rect 2006 2823 2012 2824
rect 1862 2822 1868 2823
rect 110 2811 116 2812
rect 110 2807 111 2811
rect 115 2807 116 2811
rect 2006 2811 2012 2812
rect 110 2806 116 2807
rect 278 2808 284 2809
rect 278 2804 279 2808
rect 283 2804 284 2808
rect 278 2803 284 2804
rect 446 2808 452 2809
rect 446 2804 447 2808
rect 451 2804 452 2808
rect 446 2803 452 2804
rect 630 2808 636 2809
rect 630 2804 631 2808
rect 635 2804 636 2808
rect 630 2803 636 2804
rect 814 2808 820 2809
rect 814 2804 815 2808
rect 819 2804 820 2808
rect 814 2803 820 2804
rect 998 2808 1004 2809
rect 998 2804 999 2808
rect 1003 2804 1004 2808
rect 998 2803 1004 2804
rect 1182 2808 1188 2809
rect 1182 2804 1183 2808
rect 1187 2804 1188 2808
rect 1182 2803 1188 2804
rect 1358 2808 1364 2809
rect 1358 2804 1359 2808
rect 1363 2804 1364 2808
rect 1358 2803 1364 2804
rect 1526 2808 1532 2809
rect 1526 2804 1527 2808
rect 1531 2804 1532 2808
rect 1526 2803 1532 2804
rect 1694 2808 1700 2809
rect 1694 2804 1695 2808
rect 1699 2804 1700 2808
rect 1694 2803 1700 2804
rect 1862 2808 1868 2809
rect 1862 2804 1863 2808
rect 1867 2804 1868 2808
rect 2006 2807 2007 2811
rect 2011 2807 2012 2811
rect 2006 2806 2012 2807
rect 1862 2803 1868 2804
rect 2438 2788 2444 2789
rect 2046 2785 2052 2786
rect 2046 2781 2047 2785
rect 2051 2781 2052 2785
rect 2438 2784 2439 2788
rect 2443 2784 2444 2788
rect 2438 2783 2444 2784
rect 2566 2788 2572 2789
rect 2566 2784 2567 2788
rect 2571 2784 2572 2788
rect 2566 2783 2572 2784
rect 2694 2788 2700 2789
rect 2694 2784 2695 2788
rect 2699 2784 2700 2788
rect 2694 2783 2700 2784
rect 2830 2788 2836 2789
rect 2830 2784 2831 2788
rect 2835 2784 2836 2788
rect 2830 2783 2836 2784
rect 2966 2788 2972 2789
rect 2966 2784 2967 2788
rect 2971 2784 2972 2788
rect 2966 2783 2972 2784
rect 3102 2788 3108 2789
rect 3102 2784 3103 2788
rect 3107 2784 3108 2788
rect 3102 2783 3108 2784
rect 3246 2788 3252 2789
rect 3246 2784 3247 2788
rect 3251 2784 3252 2788
rect 3246 2783 3252 2784
rect 3390 2788 3396 2789
rect 3390 2784 3391 2788
rect 3395 2784 3396 2788
rect 3390 2783 3396 2784
rect 3542 2788 3548 2789
rect 3542 2784 3543 2788
rect 3547 2784 3548 2788
rect 3542 2783 3548 2784
rect 3702 2788 3708 2789
rect 3702 2784 3703 2788
rect 3707 2784 3708 2788
rect 3702 2783 3708 2784
rect 3838 2788 3844 2789
rect 3838 2784 3839 2788
rect 3843 2784 3844 2788
rect 3838 2783 3844 2784
rect 3942 2785 3948 2786
rect 2046 2780 2052 2781
rect 3942 2781 3943 2785
rect 3947 2781 3948 2785
rect 3942 2780 3948 2781
rect 2438 2769 2444 2770
rect 2046 2768 2052 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2438 2765 2439 2769
rect 2443 2765 2444 2769
rect 2438 2764 2444 2765
rect 2566 2769 2572 2770
rect 2566 2765 2567 2769
rect 2571 2765 2572 2769
rect 2566 2764 2572 2765
rect 2694 2769 2700 2770
rect 2694 2765 2695 2769
rect 2699 2765 2700 2769
rect 2694 2764 2700 2765
rect 2830 2769 2836 2770
rect 2830 2765 2831 2769
rect 2835 2765 2836 2769
rect 2830 2764 2836 2765
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2966 2764 2972 2765
rect 3102 2769 3108 2770
rect 3102 2765 3103 2769
rect 3107 2765 3108 2769
rect 3102 2764 3108 2765
rect 3246 2769 3252 2770
rect 3246 2765 3247 2769
rect 3251 2765 3252 2769
rect 3246 2764 3252 2765
rect 3390 2769 3396 2770
rect 3390 2765 3391 2769
rect 3395 2765 3396 2769
rect 3390 2764 3396 2765
rect 3542 2769 3548 2770
rect 3542 2765 3543 2769
rect 3547 2765 3548 2769
rect 3542 2764 3548 2765
rect 3702 2769 3708 2770
rect 3702 2765 3703 2769
rect 3707 2765 3708 2769
rect 3702 2764 3708 2765
rect 3838 2769 3844 2770
rect 3838 2765 3839 2769
rect 3843 2765 3844 2769
rect 3838 2764 3844 2765
rect 3942 2768 3948 2769
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 2046 2763 2052 2764
rect 3942 2763 3948 2764
rect 238 2748 244 2749
rect 110 2745 116 2746
rect 110 2741 111 2745
rect 115 2741 116 2745
rect 238 2744 239 2748
rect 243 2744 244 2748
rect 238 2743 244 2744
rect 350 2748 356 2749
rect 350 2744 351 2748
rect 355 2744 356 2748
rect 350 2743 356 2744
rect 470 2748 476 2749
rect 470 2744 471 2748
rect 475 2744 476 2748
rect 470 2743 476 2744
rect 606 2748 612 2749
rect 606 2744 607 2748
rect 611 2744 612 2748
rect 606 2743 612 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 878 2748 884 2749
rect 878 2744 879 2748
rect 883 2744 884 2748
rect 878 2743 884 2744
rect 1014 2748 1020 2749
rect 1014 2744 1015 2748
rect 1019 2744 1020 2748
rect 1014 2743 1020 2744
rect 1150 2748 1156 2749
rect 1150 2744 1151 2748
rect 1155 2744 1156 2748
rect 1150 2743 1156 2744
rect 1286 2748 1292 2749
rect 1286 2744 1287 2748
rect 1291 2744 1292 2748
rect 1286 2743 1292 2744
rect 1422 2748 1428 2749
rect 1422 2744 1423 2748
rect 1427 2744 1428 2748
rect 1422 2743 1428 2744
rect 1566 2748 1572 2749
rect 1566 2744 1567 2748
rect 1571 2744 1572 2748
rect 1566 2743 1572 2744
rect 2006 2745 2012 2746
rect 110 2740 116 2741
rect 2006 2741 2007 2745
rect 2011 2741 2012 2745
rect 2006 2740 2012 2741
rect 238 2729 244 2730
rect 110 2728 116 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 238 2725 239 2729
rect 243 2725 244 2729
rect 238 2724 244 2725
rect 350 2729 356 2730
rect 350 2725 351 2729
rect 355 2725 356 2729
rect 350 2724 356 2725
rect 470 2729 476 2730
rect 470 2725 471 2729
rect 475 2725 476 2729
rect 470 2724 476 2725
rect 606 2729 612 2730
rect 606 2725 607 2729
rect 611 2725 612 2729
rect 606 2724 612 2725
rect 742 2729 748 2730
rect 742 2725 743 2729
rect 747 2725 748 2729
rect 742 2724 748 2725
rect 878 2729 884 2730
rect 878 2725 879 2729
rect 883 2725 884 2729
rect 878 2724 884 2725
rect 1014 2729 1020 2730
rect 1014 2725 1015 2729
rect 1019 2725 1020 2729
rect 1014 2724 1020 2725
rect 1150 2729 1156 2730
rect 1150 2725 1151 2729
rect 1155 2725 1156 2729
rect 1150 2724 1156 2725
rect 1286 2729 1292 2730
rect 1286 2725 1287 2729
rect 1291 2725 1292 2729
rect 1286 2724 1292 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1566 2729 1572 2730
rect 1566 2725 1567 2729
rect 1571 2725 1572 2729
rect 1566 2724 1572 2725
rect 2006 2728 2012 2729
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 110 2723 116 2724
rect 2006 2723 2012 2724
rect 2046 2708 2052 2709
rect 3942 2708 3948 2709
rect 2046 2704 2047 2708
rect 2051 2704 2052 2708
rect 2046 2703 2052 2704
rect 2334 2707 2340 2708
rect 2334 2703 2335 2707
rect 2339 2703 2340 2707
rect 2334 2702 2340 2703
rect 2494 2707 2500 2708
rect 2494 2703 2495 2707
rect 2499 2703 2500 2707
rect 2494 2702 2500 2703
rect 2662 2707 2668 2708
rect 2662 2703 2663 2707
rect 2667 2703 2668 2707
rect 2662 2702 2668 2703
rect 2830 2707 2836 2708
rect 2830 2703 2831 2707
rect 2835 2703 2836 2707
rect 2830 2702 2836 2703
rect 2998 2707 3004 2708
rect 2998 2703 2999 2707
rect 3003 2703 3004 2707
rect 2998 2702 3004 2703
rect 3166 2707 3172 2708
rect 3166 2703 3167 2707
rect 3171 2703 3172 2707
rect 3166 2702 3172 2703
rect 3334 2707 3340 2708
rect 3334 2703 3335 2707
rect 3339 2703 3340 2707
rect 3334 2702 3340 2703
rect 3510 2707 3516 2708
rect 3510 2703 3511 2707
rect 3515 2703 3516 2707
rect 3510 2702 3516 2703
rect 3686 2707 3692 2708
rect 3686 2703 3687 2707
rect 3691 2703 3692 2707
rect 3686 2702 3692 2703
rect 3838 2707 3844 2708
rect 3838 2703 3839 2707
rect 3843 2703 3844 2707
rect 3942 2704 3943 2708
rect 3947 2704 3948 2708
rect 3942 2703 3948 2704
rect 3838 2702 3844 2703
rect 2046 2691 2052 2692
rect 2046 2687 2047 2691
rect 2051 2687 2052 2691
rect 3942 2691 3948 2692
rect 2046 2686 2052 2687
rect 2334 2688 2340 2689
rect 2334 2684 2335 2688
rect 2339 2684 2340 2688
rect 2334 2683 2340 2684
rect 2494 2688 2500 2689
rect 2494 2684 2495 2688
rect 2499 2684 2500 2688
rect 2494 2683 2500 2684
rect 2662 2688 2668 2689
rect 2662 2684 2663 2688
rect 2667 2684 2668 2688
rect 2662 2683 2668 2684
rect 2830 2688 2836 2689
rect 2830 2684 2831 2688
rect 2835 2684 2836 2688
rect 2830 2683 2836 2684
rect 2998 2688 3004 2689
rect 2998 2684 2999 2688
rect 3003 2684 3004 2688
rect 2998 2683 3004 2684
rect 3166 2688 3172 2689
rect 3166 2684 3167 2688
rect 3171 2684 3172 2688
rect 3166 2683 3172 2684
rect 3334 2688 3340 2689
rect 3334 2684 3335 2688
rect 3339 2684 3340 2688
rect 3334 2683 3340 2684
rect 3510 2688 3516 2689
rect 3510 2684 3511 2688
rect 3515 2684 3516 2688
rect 3510 2683 3516 2684
rect 3686 2688 3692 2689
rect 3686 2684 3687 2688
rect 3691 2684 3692 2688
rect 3686 2683 3692 2684
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3942 2687 3943 2691
rect 3947 2687 3948 2691
rect 3942 2686 3948 2687
rect 3838 2683 3844 2684
rect 110 2676 116 2677
rect 2006 2676 2012 2677
rect 110 2672 111 2676
rect 115 2672 116 2676
rect 110 2671 116 2672
rect 222 2675 228 2676
rect 222 2671 223 2675
rect 227 2671 228 2675
rect 222 2670 228 2671
rect 366 2675 372 2676
rect 366 2671 367 2675
rect 371 2671 372 2675
rect 366 2670 372 2671
rect 502 2675 508 2676
rect 502 2671 503 2675
rect 507 2671 508 2675
rect 502 2670 508 2671
rect 638 2675 644 2676
rect 638 2671 639 2675
rect 643 2671 644 2675
rect 638 2670 644 2671
rect 766 2675 772 2676
rect 766 2671 767 2675
rect 771 2671 772 2675
rect 766 2670 772 2671
rect 886 2675 892 2676
rect 886 2671 887 2675
rect 891 2671 892 2675
rect 886 2670 892 2671
rect 998 2675 1004 2676
rect 998 2671 999 2675
rect 1003 2671 1004 2675
rect 998 2670 1004 2671
rect 1110 2675 1116 2676
rect 1110 2671 1111 2675
rect 1115 2671 1116 2675
rect 1110 2670 1116 2671
rect 1230 2675 1236 2676
rect 1230 2671 1231 2675
rect 1235 2671 1236 2675
rect 1230 2670 1236 2671
rect 1350 2675 1356 2676
rect 1350 2671 1351 2675
rect 1355 2671 1356 2675
rect 2006 2672 2007 2676
rect 2011 2672 2012 2676
rect 2006 2671 2012 2672
rect 1350 2670 1356 2671
rect 110 2659 116 2660
rect 110 2655 111 2659
rect 115 2655 116 2659
rect 2006 2659 2012 2660
rect 110 2654 116 2655
rect 222 2656 228 2657
rect 222 2652 223 2656
rect 227 2652 228 2656
rect 222 2651 228 2652
rect 366 2656 372 2657
rect 366 2652 367 2656
rect 371 2652 372 2656
rect 366 2651 372 2652
rect 502 2656 508 2657
rect 502 2652 503 2656
rect 507 2652 508 2656
rect 502 2651 508 2652
rect 638 2656 644 2657
rect 638 2652 639 2656
rect 643 2652 644 2656
rect 638 2651 644 2652
rect 766 2656 772 2657
rect 766 2652 767 2656
rect 771 2652 772 2656
rect 766 2651 772 2652
rect 886 2656 892 2657
rect 886 2652 887 2656
rect 891 2652 892 2656
rect 886 2651 892 2652
rect 998 2656 1004 2657
rect 998 2652 999 2656
rect 1003 2652 1004 2656
rect 998 2651 1004 2652
rect 1110 2656 1116 2657
rect 1110 2652 1111 2656
rect 1115 2652 1116 2656
rect 1110 2651 1116 2652
rect 1230 2656 1236 2657
rect 1230 2652 1231 2656
rect 1235 2652 1236 2656
rect 1230 2651 1236 2652
rect 1350 2656 1356 2657
rect 1350 2652 1351 2656
rect 1355 2652 1356 2656
rect 2006 2655 2007 2659
rect 2011 2655 2012 2659
rect 2006 2654 2012 2655
rect 1350 2651 1356 2652
rect 2126 2624 2132 2625
rect 2046 2621 2052 2622
rect 2046 2617 2047 2621
rect 2051 2617 2052 2621
rect 2126 2620 2127 2624
rect 2131 2620 2132 2624
rect 2126 2619 2132 2620
rect 2278 2624 2284 2625
rect 2278 2620 2279 2624
rect 2283 2620 2284 2624
rect 2278 2619 2284 2620
rect 2446 2624 2452 2625
rect 2446 2620 2447 2624
rect 2451 2620 2452 2624
rect 2446 2619 2452 2620
rect 2622 2624 2628 2625
rect 2622 2620 2623 2624
rect 2627 2620 2628 2624
rect 2622 2619 2628 2620
rect 2806 2624 2812 2625
rect 2806 2620 2807 2624
rect 2811 2620 2812 2624
rect 2806 2619 2812 2620
rect 2990 2624 2996 2625
rect 2990 2620 2991 2624
rect 2995 2620 2996 2624
rect 2990 2619 2996 2620
rect 3174 2624 3180 2625
rect 3174 2620 3175 2624
rect 3179 2620 3180 2624
rect 3174 2619 3180 2620
rect 3350 2624 3356 2625
rect 3350 2620 3351 2624
rect 3355 2620 3356 2624
rect 3350 2619 3356 2620
rect 3518 2624 3524 2625
rect 3518 2620 3519 2624
rect 3523 2620 3524 2624
rect 3518 2619 3524 2620
rect 3686 2624 3692 2625
rect 3686 2620 3687 2624
rect 3691 2620 3692 2624
rect 3686 2619 3692 2620
rect 3838 2624 3844 2625
rect 3838 2620 3839 2624
rect 3843 2620 3844 2624
rect 3838 2619 3844 2620
rect 3942 2621 3948 2622
rect 2046 2616 2052 2617
rect 3942 2617 3943 2621
rect 3947 2617 3948 2621
rect 3942 2616 3948 2617
rect 2126 2605 2132 2606
rect 2046 2604 2052 2605
rect 2046 2600 2047 2604
rect 2051 2600 2052 2604
rect 2126 2601 2127 2605
rect 2131 2601 2132 2605
rect 2126 2600 2132 2601
rect 2278 2605 2284 2606
rect 2278 2601 2279 2605
rect 2283 2601 2284 2605
rect 2278 2600 2284 2601
rect 2446 2605 2452 2606
rect 2446 2601 2447 2605
rect 2451 2601 2452 2605
rect 2446 2600 2452 2601
rect 2622 2605 2628 2606
rect 2622 2601 2623 2605
rect 2627 2601 2628 2605
rect 2622 2600 2628 2601
rect 2806 2605 2812 2606
rect 2806 2601 2807 2605
rect 2811 2601 2812 2605
rect 2806 2600 2812 2601
rect 2990 2605 2996 2606
rect 2990 2601 2991 2605
rect 2995 2601 2996 2605
rect 2990 2600 2996 2601
rect 3174 2605 3180 2606
rect 3174 2601 3175 2605
rect 3179 2601 3180 2605
rect 3174 2600 3180 2601
rect 3350 2605 3356 2606
rect 3350 2601 3351 2605
rect 3355 2601 3356 2605
rect 3350 2600 3356 2601
rect 3518 2605 3524 2606
rect 3518 2601 3519 2605
rect 3523 2601 3524 2605
rect 3518 2600 3524 2601
rect 3686 2605 3692 2606
rect 3686 2601 3687 2605
rect 3691 2601 3692 2605
rect 3686 2600 3692 2601
rect 3838 2605 3844 2606
rect 3838 2601 3839 2605
rect 3843 2601 3844 2605
rect 3838 2600 3844 2601
rect 3942 2604 3948 2605
rect 3942 2600 3943 2604
rect 3947 2600 3948 2604
rect 2046 2599 2052 2600
rect 3942 2599 3948 2600
rect 174 2596 180 2597
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 174 2592 175 2596
rect 179 2592 180 2596
rect 174 2591 180 2592
rect 366 2596 372 2597
rect 366 2592 367 2596
rect 371 2592 372 2596
rect 366 2591 372 2592
rect 542 2596 548 2597
rect 542 2592 543 2596
rect 547 2592 548 2596
rect 542 2591 548 2592
rect 710 2596 716 2597
rect 710 2592 711 2596
rect 715 2592 716 2596
rect 710 2591 716 2592
rect 862 2596 868 2597
rect 862 2592 863 2596
rect 867 2592 868 2596
rect 862 2591 868 2592
rect 1006 2596 1012 2597
rect 1006 2592 1007 2596
rect 1011 2592 1012 2596
rect 1006 2591 1012 2592
rect 1142 2596 1148 2597
rect 1142 2592 1143 2596
rect 1147 2592 1148 2596
rect 1142 2591 1148 2592
rect 1278 2596 1284 2597
rect 1278 2592 1279 2596
rect 1283 2592 1284 2596
rect 1278 2591 1284 2592
rect 1422 2596 1428 2597
rect 1422 2592 1423 2596
rect 1427 2592 1428 2596
rect 1422 2591 1428 2592
rect 2006 2593 2012 2594
rect 110 2588 116 2589
rect 2006 2589 2007 2593
rect 2011 2589 2012 2593
rect 2006 2588 2012 2589
rect 174 2577 180 2578
rect 110 2576 116 2577
rect 110 2572 111 2576
rect 115 2572 116 2576
rect 174 2573 175 2577
rect 179 2573 180 2577
rect 174 2572 180 2573
rect 366 2577 372 2578
rect 366 2573 367 2577
rect 371 2573 372 2577
rect 366 2572 372 2573
rect 542 2577 548 2578
rect 542 2573 543 2577
rect 547 2573 548 2577
rect 542 2572 548 2573
rect 710 2577 716 2578
rect 710 2573 711 2577
rect 715 2573 716 2577
rect 710 2572 716 2573
rect 862 2577 868 2578
rect 862 2573 863 2577
rect 867 2573 868 2577
rect 862 2572 868 2573
rect 1006 2577 1012 2578
rect 1006 2573 1007 2577
rect 1011 2573 1012 2577
rect 1006 2572 1012 2573
rect 1142 2577 1148 2578
rect 1142 2573 1143 2577
rect 1147 2573 1148 2577
rect 1142 2572 1148 2573
rect 1278 2577 1284 2578
rect 1278 2573 1279 2577
rect 1283 2573 1284 2577
rect 1278 2572 1284 2573
rect 1422 2577 1428 2578
rect 1422 2573 1423 2577
rect 1427 2573 1428 2577
rect 1422 2572 1428 2573
rect 2006 2576 2012 2577
rect 2006 2572 2007 2576
rect 2011 2572 2012 2576
rect 110 2571 116 2572
rect 2006 2571 2012 2572
rect 2046 2544 2052 2545
rect 3942 2544 3948 2545
rect 2046 2540 2047 2544
rect 2051 2540 2052 2544
rect 2046 2539 2052 2540
rect 2070 2543 2076 2544
rect 2070 2539 2071 2543
rect 2075 2539 2076 2543
rect 2070 2538 2076 2539
rect 2182 2543 2188 2544
rect 2182 2539 2183 2543
rect 2187 2539 2188 2543
rect 2182 2538 2188 2539
rect 2318 2543 2324 2544
rect 2318 2539 2319 2543
rect 2323 2539 2324 2543
rect 2318 2538 2324 2539
rect 2470 2543 2476 2544
rect 2470 2539 2471 2543
rect 2475 2539 2476 2543
rect 2470 2538 2476 2539
rect 2638 2543 2644 2544
rect 2638 2539 2639 2543
rect 2643 2539 2644 2543
rect 2638 2538 2644 2539
rect 2822 2543 2828 2544
rect 2822 2539 2823 2543
rect 2827 2539 2828 2543
rect 2822 2538 2828 2539
rect 3030 2543 3036 2544
rect 3030 2539 3031 2543
rect 3035 2539 3036 2543
rect 3030 2538 3036 2539
rect 3262 2543 3268 2544
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3502 2543 3508 2544
rect 3502 2539 3503 2543
rect 3507 2539 3508 2543
rect 3502 2538 3508 2539
rect 3742 2543 3748 2544
rect 3742 2539 3743 2543
rect 3747 2539 3748 2543
rect 3942 2540 3943 2544
rect 3947 2540 3948 2544
rect 3942 2539 3948 2540
rect 3742 2538 3748 2539
rect 2046 2527 2052 2528
rect 2046 2523 2047 2527
rect 2051 2523 2052 2527
rect 3942 2527 3948 2528
rect 2046 2522 2052 2523
rect 2070 2524 2076 2525
rect 110 2520 116 2521
rect 2006 2520 2012 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 134 2519 140 2520
rect 134 2515 135 2519
rect 139 2515 140 2519
rect 134 2514 140 2515
rect 270 2519 276 2520
rect 270 2515 271 2519
rect 275 2515 276 2519
rect 270 2514 276 2515
rect 438 2519 444 2520
rect 438 2515 439 2519
rect 443 2515 444 2519
rect 438 2514 444 2515
rect 606 2519 612 2520
rect 606 2515 607 2519
rect 611 2515 612 2519
rect 606 2514 612 2515
rect 774 2519 780 2520
rect 774 2515 775 2519
rect 779 2515 780 2519
rect 774 2514 780 2515
rect 926 2519 932 2520
rect 926 2515 927 2519
rect 931 2515 932 2519
rect 926 2514 932 2515
rect 1078 2519 1084 2520
rect 1078 2515 1079 2519
rect 1083 2515 1084 2519
rect 1078 2514 1084 2515
rect 1222 2519 1228 2520
rect 1222 2515 1223 2519
rect 1227 2515 1228 2519
rect 1222 2514 1228 2515
rect 1358 2519 1364 2520
rect 1358 2515 1359 2519
rect 1363 2515 1364 2519
rect 1358 2514 1364 2515
rect 1494 2519 1500 2520
rect 1494 2515 1495 2519
rect 1499 2515 1500 2519
rect 1494 2514 1500 2515
rect 1638 2519 1644 2520
rect 1638 2515 1639 2519
rect 1643 2515 1644 2519
rect 2006 2516 2007 2520
rect 2011 2516 2012 2520
rect 2070 2520 2071 2524
rect 2075 2520 2076 2524
rect 2070 2519 2076 2520
rect 2182 2524 2188 2525
rect 2182 2520 2183 2524
rect 2187 2520 2188 2524
rect 2182 2519 2188 2520
rect 2318 2524 2324 2525
rect 2318 2520 2319 2524
rect 2323 2520 2324 2524
rect 2318 2519 2324 2520
rect 2470 2524 2476 2525
rect 2470 2520 2471 2524
rect 2475 2520 2476 2524
rect 2470 2519 2476 2520
rect 2638 2524 2644 2525
rect 2638 2520 2639 2524
rect 2643 2520 2644 2524
rect 2638 2519 2644 2520
rect 2822 2524 2828 2525
rect 2822 2520 2823 2524
rect 2827 2520 2828 2524
rect 2822 2519 2828 2520
rect 3030 2524 3036 2525
rect 3030 2520 3031 2524
rect 3035 2520 3036 2524
rect 3030 2519 3036 2520
rect 3262 2524 3268 2525
rect 3262 2520 3263 2524
rect 3267 2520 3268 2524
rect 3262 2519 3268 2520
rect 3502 2524 3508 2525
rect 3502 2520 3503 2524
rect 3507 2520 3508 2524
rect 3502 2519 3508 2520
rect 3742 2524 3748 2525
rect 3742 2520 3743 2524
rect 3747 2520 3748 2524
rect 3942 2523 3943 2527
rect 3947 2523 3948 2527
rect 3942 2522 3948 2523
rect 3742 2519 3748 2520
rect 2006 2515 2012 2516
rect 1638 2514 1644 2515
rect 110 2503 116 2504
rect 110 2499 111 2503
rect 115 2499 116 2503
rect 2006 2503 2012 2504
rect 110 2498 116 2499
rect 134 2500 140 2501
rect 134 2496 135 2500
rect 139 2496 140 2500
rect 134 2495 140 2496
rect 270 2500 276 2501
rect 270 2496 271 2500
rect 275 2496 276 2500
rect 270 2495 276 2496
rect 438 2500 444 2501
rect 438 2496 439 2500
rect 443 2496 444 2500
rect 438 2495 444 2496
rect 606 2500 612 2501
rect 606 2496 607 2500
rect 611 2496 612 2500
rect 606 2495 612 2496
rect 774 2500 780 2501
rect 774 2496 775 2500
rect 779 2496 780 2500
rect 774 2495 780 2496
rect 926 2500 932 2501
rect 926 2496 927 2500
rect 931 2496 932 2500
rect 926 2495 932 2496
rect 1078 2500 1084 2501
rect 1078 2496 1079 2500
rect 1083 2496 1084 2500
rect 1078 2495 1084 2496
rect 1222 2500 1228 2501
rect 1222 2496 1223 2500
rect 1227 2496 1228 2500
rect 1222 2495 1228 2496
rect 1358 2500 1364 2501
rect 1358 2496 1359 2500
rect 1363 2496 1364 2500
rect 1358 2495 1364 2496
rect 1494 2500 1500 2501
rect 1494 2496 1495 2500
rect 1499 2496 1500 2500
rect 1494 2495 1500 2496
rect 1638 2500 1644 2501
rect 1638 2496 1639 2500
rect 1643 2496 1644 2500
rect 2006 2499 2007 2503
rect 2011 2499 2012 2503
rect 2006 2498 2012 2499
rect 1638 2495 1644 2496
rect 2070 2460 2076 2461
rect 2046 2457 2052 2458
rect 2046 2453 2047 2457
rect 2051 2453 2052 2457
rect 2070 2456 2071 2460
rect 2075 2456 2076 2460
rect 2070 2455 2076 2456
rect 2214 2460 2220 2461
rect 2214 2456 2215 2460
rect 2219 2456 2220 2460
rect 2214 2455 2220 2456
rect 2382 2460 2388 2461
rect 2382 2456 2383 2460
rect 2387 2456 2388 2460
rect 2382 2455 2388 2456
rect 2558 2460 2564 2461
rect 2558 2456 2559 2460
rect 2563 2456 2564 2460
rect 2558 2455 2564 2456
rect 2750 2460 2756 2461
rect 2750 2456 2751 2460
rect 2755 2456 2756 2460
rect 2750 2455 2756 2456
rect 2950 2460 2956 2461
rect 2950 2456 2951 2460
rect 2955 2456 2956 2460
rect 2950 2455 2956 2456
rect 3166 2460 3172 2461
rect 3166 2456 3167 2460
rect 3171 2456 3172 2460
rect 3166 2455 3172 2456
rect 3390 2460 3396 2461
rect 3390 2456 3391 2460
rect 3395 2456 3396 2460
rect 3390 2455 3396 2456
rect 3622 2460 3628 2461
rect 3622 2456 3623 2460
rect 3627 2456 3628 2460
rect 3622 2455 3628 2456
rect 3838 2460 3844 2461
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3838 2455 3844 2456
rect 3942 2457 3948 2458
rect 2046 2452 2052 2453
rect 3942 2453 3943 2457
rect 3947 2453 3948 2457
rect 3942 2452 3948 2453
rect 2070 2441 2076 2442
rect 2046 2440 2052 2441
rect 134 2436 140 2437
rect 110 2433 116 2434
rect 110 2429 111 2433
rect 115 2429 116 2433
rect 134 2432 135 2436
rect 139 2432 140 2436
rect 134 2431 140 2432
rect 310 2436 316 2437
rect 310 2432 311 2436
rect 315 2432 316 2436
rect 310 2431 316 2432
rect 510 2436 516 2437
rect 510 2432 511 2436
rect 515 2432 516 2436
rect 510 2431 516 2432
rect 710 2436 716 2437
rect 710 2432 711 2436
rect 715 2432 716 2436
rect 710 2431 716 2432
rect 902 2436 908 2437
rect 902 2432 903 2436
rect 907 2432 908 2436
rect 902 2431 908 2432
rect 1078 2436 1084 2437
rect 1078 2432 1079 2436
rect 1083 2432 1084 2436
rect 1078 2431 1084 2432
rect 1238 2436 1244 2437
rect 1238 2432 1239 2436
rect 1243 2432 1244 2436
rect 1238 2431 1244 2432
rect 1390 2436 1396 2437
rect 1390 2432 1391 2436
rect 1395 2432 1396 2436
rect 1390 2431 1396 2432
rect 1526 2436 1532 2437
rect 1526 2432 1527 2436
rect 1531 2432 1532 2436
rect 1526 2431 1532 2432
rect 1662 2436 1668 2437
rect 1662 2432 1663 2436
rect 1667 2432 1668 2436
rect 1662 2431 1668 2432
rect 1790 2436 1796 2437
rect 1790 2432 1791 2436
rect 1795 2432 1796 2436
rect 1790 2431 1796 2432
rect 1902 2436 1908 2437
rect 1902 2432 1903 2436
rect 1907 2432 1908 2436
rect 2046 2436 2047 2440
rect 2051 2436 2052 2440
rect 2070 2437 2071 2441
rect 2075 2437 2076 2441
rect 2070 2436 2076 2437
rect 2214 2441 2220 2442
rect 2214 2437 2215 2441
rect 2219 2437 2220 2441
rect 2214 2436 2220 2437
rect 2382 2441 2388 2442
rect 2382 2437 2383 2441
rect 2387 2437 2388 2441
rect 2382 2436 2388 2437
rect 2558 2441 2564 2442
rect 2558 2437 2559 2441
rect 2563 2437 2564 2441
rect 2558 2436 2564 2437
rect 2750 2441 2756 2442
rect 2750 2437 2751 2441
rect 2755 2437 2756 2441
rect 2750 2436 2756 2437
rect 2950 2441 2956 2442
rect 2950 2437 2951 2441
rect 2955 2437 2956 2441
rect 2950 2436 2956 2437
rect 3166 2441 3172 2442
rect 3166 2437 3167 2441
rect 3171 2437 3172 2441
rect 3166 2436 3172 2437
rect 3390 2441 3396 2442
rect 3390 2437 3391 2441
rect 3395 2437 3396 2441
rect 3390 2436 3396 2437
rect 3622 2441 3628 2442
rect 3622 2437 3623 2441
rect 3627 2437 3628 2441
rect 3622 2436 3628 2437
rect 3838 2441 3844 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3942 2440 3948 2441
rect 3942 2436 3943 2440
rect 3947 2436 3948 2440
rect 2046 2435 2052 2436
rect 3942 2435 3948 2436
rect 1902 2431 1908 2432
rect 2006 2433 2012 2434
rect 110 2428 116 2429
rect 2006 2429 2007 2433
rect 2011 2429 2012 2433
rect 2006 2428 2012 2429
rect 134 2417 140 2418
rect 110 2416 116 2417
rect 110 2412 111 2416
rect 115 2412 116 2416
rect 134 2413 135 2417
rect 139 2413 140 2417
rect 134 2412 140 2413
rect 310 2417 316 2418
rect 310 2413 311 2417
rect 315 2413 316 2417
rect 310 2412 316 2413
rect 510 2417 516 2418
rect 510 2413 511 2417
rect 515 2413 516 2417
rect 510 2412 516 2413
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 902 2417 908 2418
rect 902 2413 903 2417
rect 907 2413 908 2417
rect 902 2412 908 2413
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1238 2417 1244 2418
rect 1238 2413 1239 2417
rect 1243 2413 1244 2417
rect 1238 2412 1244 2413
rect 1390 2417 1396 2418
rect 1390 2413 1391 2417
rect 1395 2413 1396 2417
rect 1390 2412 1396 2413
rect 1526 2417 1532 2418
rect 1526 2413 1527 2417
rect 1531 2413 1532 2417
rect 1526 2412 1532 2413
rect 1662 2417 1668 2418
rect 1662 2413 1663 2417
rect 1667 2413 1668 2417
rect 1662 2412 1668 2413
rect 1790 2417 1796 2418
rect 1790 2413 1791 2417
rect 1795 2413 1796 2417
rect 1790 2412 1796 2413
rect 1902 2417 1908 2418
rect 1902 2413 1903 2417
rect 1907 2413 1908 2417
rect 1902 2412 1908 2413
rect 2006 2416 2012 2417
rect 2006 2412 2007 2416
rect 2011 2412 2012 2416
rect 110 2411 116 2412
rect 2006 2411 2012 2412
rect 2046 2372 2052 2373
rect 3942 2372 3948 2373
rect 2046 2368 2047 2372
rect 2051 2368 2052 2372
rect 2046 2367 2052 2368
rect 2070 2371 2076 2372
rect 2070 2367 2071 2371
rect 2075 2367 2076 2371
rect 2070 2366 2076 2367
rect 2246 2371 2252 2372
rect 2246 2367 2247 2371
rect 2251 2367 2252 2371
rect 2246 2366 2252 2367
rect 2430 2371 2436 2372
rect 2430 2367 2431 2371
rect 2435 2367 2436 2371
rect 2430 2366 2436 2367
rect 2606 2371 2612 2372
rect 2606 2367 2607 2371
rect 2611 2367 2612 2371
rect 2606 2366 2612 2367
rect 2774 2371 2780 2372
rect 2774 2367 2775 2371
rect 2779 2367 2780 2371
rect 2774 2366 2780 2367
rect 2934 2371 2940 2372
rect 2934 2367 2935 2371
rect 2939 2367 2940 2371
rect 2934 2366 2940 2367
rect 3102 2371 3108 2372
rect 3102 2367 3103 2371
rect 3107 2367 3108 2371
rect 3942 2368 3943 2372
rect 3947 2368 3948 2372
rect 3942 2367 3948 2368
rect 3102 2366 3108 2367
rect 110 2364 116 2365
rect 2006 2364 2012 2365
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 110 2359 116 2360
rect 134 2363 140 2364
rect 134 2359 135 2363
rect 139 2359 140 2363
rect 134 2358 140 2359
rect 326 2363 332 2364
rect 326 2359 327 2363
rect 331 2359 332 2363
rect 326 2358 332 2359
rect 550 2363 556 2364
rect 550 2359 551 2363
rect 555 2359 556 2363
rect 550 2358 556 2359
rect 766 2363 772 2364
rect 766 2359 767 2363
rect 771 2359 772 2363
rect 766 2358 772 2359
rect 974 2363 980 2364
rect 974 2359 975 2363
rect 979 2359 980 2363
rect 974 2358 980 2359
rect 1174 2363 1180 2364
rect 1174 2359 1175 2363
rect 1179 2359 1180 2363
rect 1174 2358 1180 2359
rect 1366 2363 1372 2364
rect 1366 2359 1367 2363
rect 1371 2359 1372 2363
rect 1366 2358 1372 2359
rect 1550 2363 1556 2364
rect 1550 2359 1551 2363
rect 1555 2359 1556 2363
rect 1550 2358 1556 2359
rect 1734 2363 1740 2364
rect 1734 2359 1735 2363
rect 1739 2359 1740 2363
rect 1734 2358 1740 2359
rect 1902 2363 1908 2364
rect 1902 2359 1903 2363
rect 1907 2359 1908 2363
rect 2006 2360 2007 2364
rect 2011 2360 2012 2364
rect 2006 2359 2012 2360
rect 1902 2358 1908 2359
rect 2046 2355 2052 2356
rect 2046 2351 2047 2355
rect 2051 2351 2052 2355
rect 3942 2355 3948 2356
rect 2046 2350 2052 2351
rect 2070 2352 2076 2353
rect 2070 2348 2071 2352
rect 2075 2348 2076 2352
rect 110 2347 116 2348
rect 110 2343 111 2347
rect 115 2343 116 2347
rect 2006 2347 2012 2348
rect 2070 2347 2076 2348
rect 2246 2352 2252 2353
rect 2246 2348 2247 2352
rect 2251 2348 2252 2352
rect 2246 2347 2252 2348
rect 2430 2352 2436 2353
rect 2430 2348 2431 2352
rect 2435 2348 2436 2352
rect 2430 2347 2436 2348
rect 2606 2352 2612 2353
rect 2606 2348 2607 2352
rect 2611 2348 2612 2352
rect 2606 2347 2612 2348
rect 2774 2352 2780 2353
rect 2774 2348 2775 2352
rect 2779 2348 2780 2352
rect 2774 2347 2780 2348
rect 2934 2352 2940 2353
rect 2934 2348 2935 2352
rect 2939 2348 2940 2352
rect 2934 2347 2940 2348
rect 3102 2352 3108 2353
rect 3102 2348 3103 2352
rect 3107 2348 3108 2352
rect 3942 2351 3943 2355
rect 3947 2351 3948 2355
rect 3942 2350 3948 2351
rect 3102 2347 3108 2348
rect 110 2342 116 2343
rect 134 2344 140 2345
rect 134 2340 135 2344
rect 139 2340 140 2344
rect 134 2339 140 2340
rect 326 2344 332 2345
rect 326 2340 327 2344
rect 331 2340 332 2344
rect 326 2339 332 2340
rect 550 2344 556 2345
rect 550 2340 551 2344
rect 555 2340 556 2344
rect 550 2339 556 2340
rect 766 2344 772 2345
rect 766 2340 767 2344
rect 771 2340 772 2344
rect 766 2339 772 2340
rect 974 2344 980 2345
rect 974 2340 975 2344
rect 979 2340 980 2344
rect 974 2339 980 2340
rect 1174 2344 1180 2345
rect 1174 2340 1175 2344
rect 1179 2340 1180 2344
rect 1174 2339 1180 2340
rect 1366 2344 1372 2345
rect 1366 2340 1367 2344
rect 1371 2340 1372 2344
rect 1366 2339 1372 2340
rect 1550 2344 1556 2345
rect 1550 2340 1551 2344
rect 1555 2340 1556 2344
rect 1550 2339 1556 2340
rect 1734 2344 1740 2345
rect 1734 2340 1735 2344
rect 1739 2340 1740 2344
rect 1734 2339 1740 2340
rect 1902 2344 1908 2345
rect 1902 2340 1903 2344
rect 1907 2340 1908 2344
rect 2006 2343 2007 2347
rect 2011 2343 2012 2347
rect 2006 2342 2012 2343
rect 1902 2339 1908 2340
rect 2070 2292 2076 2293
rect 2046 2289 2052 2290
rect 2046 2285 2047 2289
rect 2051 2285 2052 2289
rect 2070 2288 2071 2292
rect 2075 2288 2076 2292
rect 2070 2287 2076 2288
rect 2174 2292 2180 2293
rect 2174 2288 2175 2292
rect 2179 2288 2180 2292
rect 2174 2287 2180 2288
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2446 2292 2452 2293
rect 2446 2288 2447 2292
rect 2451 2288 2452 2292
rect 2446 2287 2452 2288
rect 2590 2292 2596 2293
rect 2590 2288 2591 2292
rect 2595 2288 2596 2292
rect 2590 2287 2596 2288
rect 2750 2292 2756 2293
rect 2750 2288 2751 2292
rect 2755 2288 2756 2292
rect 2750 2287 2756 2288
rect 2934 2292 2940 2293
rect 2934 2288 2935 2292
rect 2939 2288 2940 2292
rect 2934 2287 2940 2288
rect 3142 2292 3148 2293
rect 3142 2288 3143 2292
rect 3147 2288 3148 2292
rect 3142 2287 3148 2288
rect 3374 2292 3380 2293
rect 3374 2288 3375 2292
rect 3379 2288 3380 2292
rect 3374 2287 3380 2288
rect 3614 2292 3620 2293
rect 3614 2288 3615 2292
rect 3619 2288 3620 2292
rect 3614 2287 3620 2288
rect 3838 2292 3844 2293
rect 3838 2288 3839 2292
rect 3843 2288 3844 2292
rect 3838 2287 3844 2288
rect 3942 2289 3948 2290
rect 2046 2284 2052 2285
rect 3942 2285 3943 2289
rect 3947 2285 3948 2289
rect 3942 2284 3948 2285
rect 134 2276 140 2277
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 134 2272 135 2276
rect 139 2272 140 2276
rect 134 2271 140 2272
rect 270 2276 276 2277
rect 270 2272 271 2276
rect 275 2272 276 2276
rect 270 2271 276 2272
rect 430 2276 436 2277
rect 430 2272 431 2276
rect 435 2272 436 2276
rect 430 2271 436 2272
rect 590 2276 596 2277
rect 590 2272 591 2276
rect 595 2272 596 2276
rect 590 2271 596 2272
rect 750 2276 756 2277
rect 750 2272 751 2276
rect 755 2272 756 2276
rect 750 2271 756 2272
rect 918 2276 924 2277
rect 918 2272 919 2276
rect 923 2272 924 2276
rect 918 2271 924 2272
rect 1086 2276 1092 2277
rect 1086 2272 1087 2276
rect 1091 2272 1092 2276
rect 1086 2271 1092 2272
rect 1262 2276 1268 2277
rect 1262 2272 1263 2276
rect 1267 2272 1268 2276
rect 1262 2271 1268 2272
rect 1446 2276 1452 2277
rect 1446 2272 1447 2276
rect 1451 2272 1452 2276
rect 1446 2271 1452 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1814 2271 1820 2272
rect 2006 2273 2012 2274
rect 2070 2273 2076 2274
rect 110 2268 116 2269
rect 2006 2269 2007 2273
rect 2011 2269 2012 2273
rect 2006 2268 2012 2269
rect 2046 2272 2052 2273
rect 2046 2268 2047 2272
rect 2051 2268 2052 2272
rect 2070 2269 2071 2273
rect 2075 2269 2076 2273
rect 2070 2268 2076 2269
rect 2174 2273 2180 2274
rect 2174 2269 2175 2273
rect 2179 2269 2180 2273
rect 2174 2268 2180 2269
rect 2310 2273 2316 2274
rect 2310 2269 2311 2273
rect 2315 2269 2316 2273
rect 2310 2268 2316 2269
rect 2446 2273 2452 2274
rect 2446 2269 2447 2273
rect 2451 2269 2452 2273
rect 2446 2268 2452 2269
rect 2590 2273 2596 2274
rect 2590 2269 2591 2273
rect 2595 2269 2596 2273
rect 2590 2268 2596 2269
rect 2750 2273 2756 2274
rect 2750 2269 2751 2273
rect 2755 2269 2756 2273
rect 2750 2268 2756 2269
rect 2934 2273 2940 2274
rect 2934 2269 2935 2273
rect 2939 2269 2940 2273
rect 2934 2268 2940 2269
rect 3142 2273 3148 2274
rect 3142 2269 3143 2273
rect 3147 2269 3148 2273
rect 3142 2268 3148 2269
rect 3374 2273 3380 2274
rect 3374 2269 3375 2273
rect 3379 2269 3380 2273
rect 3374 2268 3380 2269
rect 3614 2273 3620 2274
rect 3614 2269 3615 2273
rect 3619 2269 3620 2273
rect 3614 2268 3620 2269
rect 3838 2273 3844 2274
rect 3838 2269 3839 2273
rect 3843 2269 3844 2273
rect 3838 2268 3844 2269
rect 3942 2272 3948 2273
rect 3942 2268 3943 2272
rect 3947 2268 3948 2272
rect 2046 2267 2052 2268
rect 3942 2267 3948 2268
rect 134 2257 140 2258
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 134 2253 135 2257
rect 139 2253 140 2257
rect 134 2252 140 2253
rect 270 2257 276 2258
rect 270 2253 271 2257
rect 275 2253 276 2257
rect 270 2252 276 2253
rect 430 2257 436 2258
rect 430 2253 431 2257
rect 435 2253 436 2257
rect 430 2252 436 2253
rect 590 2257 596 2258
rect 590 2253 591 2257
rect 595 2253 596 2257
rect 590 2252 596 2253
rect 750 2257 756 2258
rect 750 2253 751 2257
rect 755 2253 756 2257
rect 750 2252 756 2253
rect 918 2257 924 2258
rect 918 2253 919 2257
rect 923 2253 924 2257
rect 918 2252 924 2253
rect 1086 2257 1092 2258
rect 1086 2253 1087 2257
rect 1091 2253 1092 2257
rect 1086 2252 1092 2253
rect 1262 2257 1268 2258
rect 1262 2253 1263 2257
rect 1267 2253 1268 2257
rect 1262 2252 1268 2253
rect 1446 2257 1452 2258
rect 1446 2253 1447 2257
rect 1451 2253 1452 2257
rect 1446 2252 1452 2253
rect 1630 2257 1636 2258
rect 1630 2253 1631 2257
rect 1635 2253 1636 2257
rect 1630 2252 1636 2253
rect 1814 2257 1820 2258
rect 1814 2253 1815 2257
rect 1819 2253 1820 2257
rect 1814 2252 1820 2253
rect 2006 2256 2012 2257
rect 2006 2252 2007 2256
rect 2011 2252 2012 2256
rect 110 2251 116 2252
rect 2006 2251 2012 2252
rect 2046 2212 2052 2213
rect 3942 2212 3948 2213
rect 2046 2208 2047 2212
rect 2051 2208 2052 2212
rect 2046 2207 2052 2208
rect 2110 2211 2116 2212
rect 2110 2207 2111 2211
rect 2115 2207 2116 2211
rect 2110 2206 2116 2207
rect 2254 2211 2260 2212
rect 2254 2207 2255 2211
rect 2259 2207 2260 2211
rect 2254 2206 2260 2207
rect 2406 2211 2412 2212
rect 2406 2207 2407 2211
rect 2411 2207 2412 2211
rect 2406 2206 2412 2207
rect 2558 2211 2564 2212
rect 2558 2207 2559 2211
rect 2563 2207 2564 2211
rect 2558 2206 2564 2207
rect 2718 2211 2724 2212
rect 2718 2207 2719 2211
rect 2723 2207 2724 2211
rect 2718 2206 2724 2207
rect 2878 2211 2884 2212
rect 2878 2207 2879 2211
rect 2883 2207 2884 2211
rect 2878 2206 2884 2207
rect 3046 2211 3052 2212
rect 3046 2207 3047 2211
rect 3051 2207 3052 2211
rect 3046 2206 3052 2207
rect 3222 2211 3228 2212
rect 3222 2207 3223 2211
rect 3227 2207 3228 2211
rect 3222 2206 3228 2207
rect 3406 2211 3412 2212
rect 3406 2207 3407 2211
rect 3411 2207 3412 2211
rect 3406 2206 3412 2207
rect 3590 2211 3596 2212
rect 3590 2207 3591 2211
rect 3595 2207 3596 2211
rect 3590 2206 3596 2207
rect 3782 2211 3788 2212
rect 3782 2207 3783 2211
rect 3787 2207 3788 2211
rect 3942 2208 3943 2212
rect 3947 2208 3948 2212
rect 3942 2207 3948 2208
rect 3782 2206 3788 2207
rect 110 2204 116 2205
rect 2006 2204 2012 2205
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 110 2199 116 2200
rect 158 2203 164 2204
rect 158 2199 159 2203
rect 163 2199 164 2203
rect 158 2198 164 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 678 2203 684 2204
rect 678 2199 679 2203
rect 683 2199 684 2203
rect 678 2198 684 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 1094 2203 1100 2204
rect 1094 2199 1095 2203
rect 1099 2199 1100 2203
rect 1094 2198 1100 2199
rect 1326 2203 1332 2204
rect 1326 2199 1327 2203
rect 1331 2199 1332 2203
rect 1326 2198 1332 2199
rect 1566 2203 1572 2204
rect 1566 2199 1567 2203
rect 1571 2199 1572 2203
rect 1566 2198 1572 2199
rect 1814 2203 1820 2204
rect 1814 2199 1815 2203
rect 1819 2199 1820 2203
rect 2006 2200 2007 2204
rect 2011 2200 2012 2204
rect 2006 2199 2012 2200
rect 1814 2198 1820 2199
rect 2046 2195 2052 2196
rect 2046 2191 2047 2195
rect 2051 2191 2052 2195
rect 3942 2195 3948 2196
rect 2046 2190 2052 2191
rect 2110 2192 2116 2193
rect 2110 2188 2111 2192
rect 2115 2188 2116 2192
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 2006 2187 2012 2188
rect 2110 2187 2116 2188
rect 2254 2192 2260 2193
rect 2254 2188 2255 2192
rect 2259 2188 2260 2192
rect 2254 2187 2260 2188
rect 2406 2192 2412 2193
rect 2406 2188 2407 2192
rect 2411 2188 2412 2192
rect 2406 2187 2412 2188
rect 2558 2192 2564 2193
rect 2558 2188 2559 2192
rect 2563 2188 2564 2192
rect 2558 2187 2564 2188
rect 2718 2192 2724 2193
rect 2718 2188 2719 2192
rect 2723 2188 2724 2192
rect 2718 2187 2724 2188
rect 2878 2192 2884 2193
rect 2878 2188 2879 2192
rect 2883 2188 2884 2192
rect 2878 2187 2884 2188
rect 3046 2192 3052 2193
rect 3046 2188 3047 2192
rect 3051 2188 3052 2192
rect 3046 2187 3052 2188
rect 3222 2192 3228 2193
rect 3222 2188 3223 2192
rect 3227 2188 3228 2192
rect 3222 2187 3228 2188
rect 3406 2192 3412 2193
rect 3406 2188 3407 2192
rect 3411 2188 3412 2192
rect 3406 2187 3412 2188
rect 3590 2192 3596 2193
rect 3590 2188 3591 2192
rect 3595 2188 3596 2192
rect 3590 2187 3596 2188
rect 3782 2192 3788 2193
rect 3782 2188 3783 2192
rect 3787 2188 3788 2192
rect 3942 2191 3943 2195
rect 3947 2191 3948 2195
rect 3942 2190 3948 2191
rect 3782 2187 3788 2188
rect 110 2182 116 2183
rect 158 2184 164 2185
rect 158 2180 159 2184
rect 163 2180 164 2184
rect 158 2179 164 2180
rect 326 2184 332 2185
rect 326 2180 327 2184
rect 331 2180 332 2184
rect 326 2179 332 2180
rect 494 2184 500 2185
rect 494 2180 495 2184
rect 499 2180 500 2184
rect 494 2179 500 2180
rect 678 2184 684 2185
rect 678 2180 679 2184
rect 683 2180 684 2184
rect 678 2179 684 2180
rect 878 2184 884 2185
rect 878 2180 879 2184
rect 883 2180 884 2184
rect 878 2179 884 2180
rect 1094 2184 1100 2185
rect 1094 2180 1095 2184
rect 1099 2180 1100 2184
rect 1094 2179 1100 2180
rect 1326 2184 1332 2185
rect 1326 2180 1327 2184
rect 1331 2180 1332 2184
rect 1326 2179 1332 2180
rect 1566 2184 1572 2185
rect 1566 2180 1567 2184
rect 1571 2180 1572 2184
rect 1566 2179 1572 2180
rect 1814 2184 1820 2185
rect 1814 2180 1815 2184
rect 1819 2180 1820 2184
rect 2006 2183 2007 2187
rect 2011 2183 2012 2187
rect 2006 2182 2012 2183
rect 1814 2179 1820 2180
rect 222 2124 228 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 222 2120 223 2124
rect 227 2120 228 2124
rect 222 2119 228 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 494 2124 500 2125
rect 494 2120 495 2124
rect 499 2120 500 2124
rect 494 2119 500 2120
rect 638 2124 644 2125
rect 638 2120 639 2124
rect 643 2120 644 2124
rect 638 2119 644 2120
rect 782 2124 788 2125
rect 782 2120 783 2124
rect 787 2120 788 2124
rect 782 2119 788 2120
rect 934 2124 940 2125
rect 934 2120 935 2124
rect 939 2120 940 2124
rect 934 2119 940 2120
rect 1094 2124 1100 2125
rect 1094 2120 1095 2124
rect 1099 2120 1100 2124
rect 1094 2119 1100 2120
rect 1262 2124 1268 2125
rect 1262 2120 1263 2124
rect 1267 2120 1268 2124
rect 1262 2119 1268 2120
rect 1446 2124 1452 2125
rect 1446 2120 1447 2124
rect 1451 2120 1452 2124
rect 1446 2119 1452 2120
rect 1630 2124 1636 2125
rect 1630 2120 1631 2124
rect 1635 2120 1636 2124
rect 1630 2119 1636 2120
rect 1822 2124 1828 2125
rect 1822 2120 1823 2124
rect 1827 2120 1828 2124
rect 1822 2119 1828 2120
rect 2006 2121 2012 2122
rect 110 2116 116 2117
rect 2006 2117 2007 2121
rect 2011 2117 2012 2121
rect 2286 2120 2292 2121
rect 2006 2116 2012 2117
rect 2046 2117 2052 2118
rect 2046 2113 2047 2117
rect 2051 2113 2052 2117
rect 2286 2116 2287 2120
rect 2291 2116 2292 2120
rect 2286 2115 2292 2116
rect 2430 2120 2436 2121
rect 2430 2116 2431 2120
rect 2435 2116 2436 2120
rect 2430 2115 2436 2116
rect 2582 2120 2588 2121
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2734 2120 2740 2121
rect 2734 2116 2735 2120
rect 2739 2116 2740 2120
rect 2734 2115 2740 2116
rect 2886 2120 2892 2121
rect 2886 2116 2887 2120
rect 2891 2116 2892 2120
rect 2886 2115 2892 2116
rect 3046 2120 3052 2121
rect 3046 2116 3047 2120
rect 3051 2116 3052 2120
rect 3046 2115 3052 2116
rect 3206 2120 3212 2121
rect 3206 2116 3207 2120
rect 3211 2116 3212 2120
rect 3206 2115 3212 2116
rect 3366 2120 3372 2121
rect 3366 2116 3367 2120
rect 3371 2116 3372 2120
rect 3366 2115 3372 2116
rect 3526 2120 3532 2121
rect 3526 2116 3527 2120
rect 3531 2116 3532 2120
rect 3526 2115 3532 2116
rect 3694 2120 3700 2121
rect 3694 2116 3695 2120
rect 3699 2116 3700 2120
rect 3694 2115 3700 2116
rect 3838 2120 3844 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3838 2115 3844 2116
rect 3942 2117 3948 2118
rect 2046 2112 2052 2113
rect 3942 2113 3943 2117
rect 3947 2113 3948 2117
rect 3942 2112 3948 2113
rect 222 2105 228 2106
rect 110 2104 116 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 222 2101 223 2105
rect 227 2101 228 2105
rect 222 2100 228 2101
rect 358 2105 364 2106
rect 358 2101 359 2105
rect 363 2101 364 2105
rect 358 2100 364 2101
rect 494 2105 500 2106
rect 494 2101 495 2105
rect 499 2101 500 2105
rect 494 2100 500 2101
rect 638 2105 644 2106
rect 638 2101 639 2105
rect 643 2101 644 2105
rect 638 2100 644 2101
rect 782 2105 788 2106
rect 782 2101 783 2105
rect 787 2101 788 2105
rect 782 2100 788 2101
rect 934 2105 940 2106
rect 934 2101 935 2105
rect 939 2101 940 2105
rect 934 2100 940 2101
rect 1094 2105 1100 2106
rect 1094 2101 1095 2105
rect 1099 2101 1100 2105
rect 1094 2100 1100 2101
rect 1262 2105 1268 2106
rect 1262 2101 1263 2105
rect 1267 2101 1268 2105
rect 1262 2100 1268 2101
rect 1446 2105 1452 2106
rect 1446 2101 1447 2105
rect 1451 2101 1452 2105
rect 1446 2100 1452 2101
rect 1630 2105 1636 2106
rect 1630 2101 1631 2105
rect 1635 2101 1636 2105
rect 1630 2100 1636 2101
rect 1822 2105 1828 2106
rect 1822 2101 1823 2105
rect 1827 2101 1828 2105
rect 1822 2100 1828 2101
rect 2006 2104 2012 2105
rect 2006 2100 2007 2104
rect 2011 2100 2012 2104
rect 2286 2101 2292 2102
rect 110 2099 116 2100
rect 2006 2099 2012 2100
rect 2046 2100 2052 2101
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2286 2097 2287 2101
rect 2291 2097 2292 2101
rect 2286 2096 2292 2097
rect 2430 2101 2436 2102
rect 2430 2097 2431 2101
rect 2435 2097 2436 2101
rect 2430 2096 2436 2097
rect 2582 2101 2588 2102
rect 2582 2097 2583 2101
rect 2587 2097 2588 2101
rect 2582 2096 2588 2097
rect 2734 2101 2740 2102
rect 2734 2097 2735 2101
rect 2739 2097 2740 2101
rect 2734 2096 2740 2097
rect 2886 2101 2892 2102
rect 2886 2097 2887 2101
rect 2891 2097 2892 2101
rect 2886 2096 2892 2097
rect 3046 2101 3052 2102
rect 3046 2097 3047 2101
rect 3051 2097 3052 2101
rect 3046 2096 3052 2097
rect 3206 2101 3212 2102
rect 3206 2097 3207 2101
rect 3211 2097 3212 2101
rect 3206 2096 3212 2097
rect 3366 2101 3372 2102
rect 3366 2097 3367 2101
rect 3371 2097 3372 2101
rect 3366 2096 3372 2097
rect 3526 2101 3532 2102
rect 3526 2097 3527 2101
rect 3531 2097 3532 2101
rect 3526 2096 3532 2097
rect 3694 2101 3700 2102
rect 3694 2097 3695 2101
rect 3699 2097 3700 2101
rect 3694 2096 3700 2097
rect 3838 2101 3844 2102
rect 3838 2097 3839 2101
rect 3843 2097 3844 2101
rect 3838 2096 3844 2097
rect 3942 2100 3948 2101
rect 3942 2096 3943 2100
rect 3947 2096 3948 2100
rect 2046 2095 2052 2096
rect 3942 2095 3948 2096
rect 110 2044 116 2045
rect 2006 2044 2012 2045
rect 110 2040 111 2044
rect 115 2040 116 2044
rect 110 2039 116 2040
rect 374 2043 380 2044
rect 374 2039 375 2043
rect 379 2039 380 2043
rect 374 2038 380 2039
rect 494 2043 500 2044
rect 494 2039 495 2043
rect 499 2039 500 2043
rect 494 2038 500 2039
rect 614 2043 620 2044
rect 614 2039 615 2043
rect 619 2039 620 2043
rect 614 2038 620 2039
rect 750 2043 756 2044
rect 750 2039 751 2043
rect 755 2039 756 2043
rect 750 2038 756 2039
rect 894 2043 900 2044
rect 894 2039 895 2043
rect 899 2039 900 2043
rect 894 2038 900 2039
rect 1046 2043 1052 2044
rect 1046 2039 1047 2043
rect 1051 2039 1052 2043
rect 1046 2038 1052 2039
rect 1214 2043 1220 2044
rect 1214 2039 1215 2043
rect 1219 2039 1220 2043
rect 1214 2038 1220 2039
rect 1398 2043 1404 2044
rect 1398 2039 1399 2043
rect 1403 2039 1404 2043
rect 1398 2038 1404 2039
rect 1582 2043 1588 2044
rect 1582 2039 1583 2043
rect 1587 2039 1588 2043
rect 1582 2038 1588 2039
rect 1774 2043 1780 2044
rect 1774 2039 1775 2043
rect 1779 2039 1780 2043
rect 2006 2040 2007 2044
rect 2011 2040 2012 2044
rect 2006 2039 2012 2040
rect 2046 2040 2052 2041
rect 3942 2040 3948 2041
rect 1774 2038 1780 2039
rect 2046 2036 2047 2040
rect 2051 2036 2052 2040
rect 2046 2035 2052 2036
rect 2502 2039 2508 2040
rect 2502 2035 2503 2039
rect 2507 2035 2508 2039
rect 2502 2034 2508 2035
rect 2670 2039 2676 2040
rect 2670 2035 2671 2039
rect 2675 2035 2676 2039
rect 2670 2034 2676 2035
rect 2838 2039 2844 2040
rect 2838 2035 2839 2039
rect 2843 2035 2844 2039
rect 2838 2034 2844 2035
rect 3006 2039 3012 2040
rect 3006 2035 3007 2039
rect 3011 2035 3012 2039
rect 3006 2034 3012 2035
rect 3166 2039 3172 2040
rect 3166 2035 3167 2039
rect 3171 2035 3172 2039
rect 3166 2034 3172 2035
rect 3310 2039 3316 2040
rect 3310 2035 3311 2039
rect 3315 2035 3316 2039
rect 3310 2034 3316 2035
rect 3454 2039 3460 2040
rect 3454 2035 3455 2039
rect 3459 2035 3460 2039
rect 3454 2034 3460 2035
rect 3590 2039 3596 2040
rect 3590 2035 3591 2039
rect 3595 2035 3596 2039
rect 3590 2034 3596 2035
rect 3726 2039 3732 2040
rect 3726 2035 3727 2039
rect 3731 2035 3732 2039
rect 3726 2034 3732 2035
rect 3838 2039 3844 2040
rect 3838 2035 3839 2039
rect 3843 2035 3844 2039
rect 3942 2036 3943 2040
rect 3947 2036 3948 2040
rect 3942 2035 3948 2036
rect 3838 2034 3844 2035
rect 110 2027 116 2028
rect 110 2023 111 2027
rect 115 2023 116 2027
rect 2006 2027 2012 2028
rect 110 2022 116 2023
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 494 2024 500 2025
rect 494 2020 495 2024
rect 499 2020 500 2024
rect 494 2019 500 2020
rect 614 2024 620 2025
rect 614 2020 615 2024
rect 619 2020 620 2024
rect 614 2019 620 2020
rect 750 2024 756 2025
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 894 2024 900 2025
rect 894 2020 895 2024
rect 899 2020 900 2024
rect 894 2019 900 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1214 2024 1220 2025
rect 1214 2020 1215 2024
rect 1219 2020 1220 2024
rect 1214 2019 1220 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1582 2024 1588 2025
rect 1582 2020 1583 2024
rect 1587 2020 1588 2024
rect 1582 2019 1588 2020
rect 1774 2024 1780 2025
rect 1774 2020 1775 2024
rect 1779 2020 1780 2024
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2006 2022 2012 2023
rect 2046 2023 2052 2024
rect 1774 2019 1780 2020
rect 2046 2019 2047 2023
rect 2051 2019 2052 2023
rect 3942 2023 3948 2024
rect 2046 2018 2052 2019
rect 2502 2020 2508 2021
rect 2502 2016 2503 2020
rect 2507 2016 2508 2020
rect 2502 2015 2508 2016
rect 2670 2020 2676 2021
rect 2670 2016 2671 2020
rect 2675 2016 2676 2020
rect 2670 2015 2676 2016
rect 2838 2020 2844 2021
rect 2838 2016 2839 2020
rect 2843 2016 2844 2020
rect 2838 2015 2844 2016
rect 3006 2020 3012 2021
rect 3006 2016 3007 2020
rect 3011 2016 3012 2020
rect 3006 2015 3012 2016
rect 3166 2020 3172 2021
rect 3166 2016 3167 2020
rect 3171 2016 3172 2020
rect 3166 2015 3172 2016
rect 3310 2020 3316 2021
rect 3310 2016 3311 2020
rect 3315 2016 3316 2020
rect 3310 2015 3316 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3590 2020 3596 2021
rect 3590 2016 3591 2020
rect 3595 2016 3596 2020
rect 3590 2015 3596 2016
rect 3726 2020 3732 2021
rect 3726 2016 3727 2020
rect 3731 2016 3732 2020
rect 3726 2015 3732 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3942 2019 3943 2023
rect 3947 2019 3948 2023
rect 3942 2018 3948 2019
rect 3838 2015 3844 2016
rect 510 1956 516 1957
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 510 1952 511 1956
rect 515 1952 516 1956
rect 510 1951 516 1952
rect 622 1956 628 1957
rect 622 1952 623 1956
rect 627 1952 628 1956
rect 622 1951 628 1952
rect 742 1956 748 1957
rect 742 1952 743 1956
rect 747 1952 748 1956
rect 742 1951 748 1952
rect 870 1956 876 1957
rect 870 1952 871 1956
rect 875 1952 876 1956
rect 870 1951 876 1952
rect 1006 1956 1012 1957
rect 1006 1952 1007 1956
rect 1011 1952 1012 1956
rect 1006 1951 1012 1952
rect 1142 1956 1148 1957
rect 1142 1952 1143 1956
rect 1147 1952 1148 1956
rect 1142 1951 1148 1952
rect 1278 1956 1284 1957
rect 1278 1952 1279 1956
rect 1283 1952 1284 1956
rect 1278 1951 1284 1952
rect 1414 1956 1420 1957
rect 1414 1952 1415 1956
rect 1419 1952 1420 1956
rect 1414 1951 1420 1952
rect 1558 1956 1564 1957
rect 1558 1952 1559 1956
rect 1563 1952 1564 1956
rect 1558 1951 1564 1952
rect 1702 1956 1708 1957
rect 1702 1952 1703 1956
rect 1707 1952 1708 1956
rect 2494 1956 2500 1957
rect 1702 1951 1708 1952
rect 2006 1953 2012 1954
rect 110 1948 116 1949
rect 2006 1949 2007 1953
rect 2011 1949 2012 1953
rect 2006 1948 2012 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2494 1952 2495 1956
rect 2499 1952 2500 1956
rect 2494 1951 2500 1952
rect 2590 1956 2596 1957
rect 2590 1952 2591 1956
rect 2595 1952 2596 1956
rect 2590 1951 2596 1952
rect 2694 1956 2700 1957
rect 2694 1952 2695 1956
rect 2699 1952 2700 1956
rect 2694 1951 2700 1952
rect 2806 1956 2812 1957
rect 2806 1952 2807 1956
rect 2811 1952 2812 1956
rect 2806 1951 2812 1952
rect 2926 1956 2932 1957
rect 2926 1952 2927 1956
rect 2931 1952 2932 1956
rect 2926 1951 2932 1952
rect 3046 1956 3052 1957
rect 3046 1952 3047 1956
rect 3051 1952 3052 1956
rect 3046 1951 3052 1952
rect 3174 1956 3180 1957
rect 3174 1952 3175 1956
rect 3179 1952 3180 1956
rect 3174 1951 3180 1952
rect 3294 1956 3300 1957
rect 3294 1952 3295 1956
rect 3299 1952 3300 1956
rect 3294 1951 3300 1952
rect 3414 1956 3420 1957
rect 3414 1952 3415 1956
rect 3419 1952 3420 1956
rect 3414 1951 3420 1952
rect 3542 1956 3548 1957
rect 3542 1952 3543 1956
rect 3547 1952 3548 1956
rect 3542 1951 3548 1952
rect 3670 1956 3676 1957
rect 3670 1952 3671 1956
rect 3675 1952 3676 1956
rect 3670 1951 3676 1952
rect 3798 1956 3804 1957
rect 3798 1952 3799 1956
rect 3803 1952 3804 1956
rect 3798 1951 3804 1952
rect 3942 1953 3948 1954
rect 2046 1948 2052 1949
rect 3942 1949 3943 1953
rect 3947 1949 3948 1953
rect 3942 1948 3948 1949
rect 510 1937 516 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 510 1933 511 1937
rect 515 1933 516 1937
rect 510 1932 516 1933
rect 622 1937 628 1938
rect 622 1933 623 1937
rect 627 1933 628 1937
rect 622 1932 628 1933
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 870 1937 876 1938
rect 870 1933 871 1937
rect 875 1933 876 1937
rect 870 1932 876 1933
rect 1006 1937 1012 1938
rect 1006 1933 1007 1937
rect 1011 1933 1012 1937
rect 1006 1932 1012 1933
rect 1142 1937 1148 1938
rect 1142 1933 1143 1937
rect 1147 1933 1148 1937
rect 1142 1932 1148 1933
rect 1278 1937 1284 1938
rect 1278 1933 1279 1937
rect 1283 1933 1284 1937
rect 1278 1932 1284 1933
rect 1414 1937 1420 1938
rect 1414 1933 1415 1937
rect 1419 1933 1420 1937
rect 1414 1932 1420 1933
rect 1558 1937 1564 1938
rect 1558 1933 1559 1937
rect 1563 1933 1564 1937
rect 1558 1932 1564 1933
rect 1702 1937 1708 1938
rect 2494 1937 2500 1938
rect 1702 1933 1703 1937
rect 1707 1933 1708 1937
rect 1702 1932 1708 1933
rect 2006 1936 2012 1937
rect 2006 1932 2007 1936
rect 2011 1932 2012 1936
rect 110 1931 116 1932
rect 2006 1931 2012 1932
rect 2046 1936 2052 1937
rect 2046 1932 2047 1936
rect 2051 1932 2052 1936
rect 2494 1933 2495 1937
rect 2499 1933 2500 1937
rect 2494 1932 2500 1933
rect 2590 1937 2596 1938
rect 2590 1933 2591 1937
rect 2595 1933 2596 1937
rect 2590 1932 2596 1933
rect 2694 1937 2700 1938
rect 2694 1933 2695 1937
rect 2699 1933 2700 1937
rect 2694 1932 2700 1933
rect 2806 1937 2812 1938
rect 2806 1933 2807 1937
rect 2811 1933 2812 1937
rect 2806 1932 2812 1933
rect 2926 1937 2932 1938
rect 2926 1933 2927 1937
rect 2931 1933 2932 1937
rect 2926 1932 2932 1933
rect 3046 1937 3052 1938
rect 3046 1933 3047 1937
rect 3051 1933 3052 1937
rect 3046 1932 3052 1933
rect 3174 1937 3180 1938
rect 3174 1933 3175 1937
rect 3179 1933 3180 1937
rect 3174 1932 3180 1933
rect 3294 1937 3300 1938
rect 3294 1933 3295 1937
rect 3299 1933 3300 1937
rect 3294 1932 3300 1933
rect 3414 1937 3420 1938
rect 3414 1933 3415 1937
rect 3419 1933 3420 1937
rect 3414 1932 3420 1933
rect 3542 1937 3548 1938
rect 3542 1933 3543 1937
rect 3547 1933 3548 1937
rect 3542 1932 3548 1933
rect 3670 1937 3676 1938
rect 3670 1933 3671 1937
rect 3675 1933 3676 1937
rect 3670 1932 3676 1933
rect 3798 1937 3804 1938
rect 3798 1933 3799 1937
rect 3803 1933 3804 1937
rect 3798 1932 3804 1933
rect 3942 1936 3948 1937
rect 3942 1932 3943 1936
rect 3947 1932 3948 1936
rect 2046 1931 2052 1932
rect 3942 1931 3948 1932
rect 2046 1880 2052 1881
rect 3942 1880 3948 1881
rect 110 1876 116 1877
rect 2006 1876 2012 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 550 1875 556 1876
rect 550 1871 551 1875
rect 555 1871 556 1875
rect 550 1870 556 1871
rect 662 1875 668 1876
rect 662 1871 663 1875
rect 667 1871 668 1875
rect 662 1870 668 1871
rect 782 1875 788 1876
rect 782 1871 783 1875
rect 787 1871 788 1875
rect 782 1870 788 1871
rect 910 1875 916 1876
rect 910 1871 911 1875
rect 915 1871 916 1875
rect 910 1870 916 1871
rect 1046 1875 1052 1876
rect 1046 1871 1047 1875
rect 1051 1871 1052 1875
rect 1046 1870 1052 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1174 1870 1180 1871
rect 1310 1875 1316 1876
rect 1310 1871 1311 1875
rect 1315 1871 1316 1875
rect 1310 1870 1316 1871
rect 1446 1875 1452 1876
rect 1446 1871 1447 1875
rect 1451 1871 1452 1875
rect 1446 1870 1452 1871
rect 1582 1875 1588 1876
rect 1582 1871 1583 1875
rect 1587 1871 1588 1875
rect 1582 1870 1588 1871
rect 1718 1875 1724 1876
rect 1718 1871 1719 1875
rect 1723 1871 1724 1875
rect 2006 1872 2007 1876
rect 2011 1872 2012 1876
rect 2046 1876 2047 1880
rect 2051 1876 2052 1880
rect 2046 1875 2052 1876
rect 2070 1879 2076 1880
rect 2070 1875 2071 1879
rect 2075 1875 2076 1879
rect 2070 1874 2076 1875
rect 2246 1879 2252 1880
rect 2246 1875 2247 1879
rect 2251 1875 2252 1879
rect 2246 1874 2252 1875
rect 2438 1879 2444 1880
rect 2438 1875 2439 1879
rect 2443 1875 2444 1879
rect 2438 1874 2444 1875
rect 2622 1879 2628 1880
rect 2622 1875 2623 1879
rect 2627 1875 2628 1879
rect 2622 1874 2628 1875
rect 2790 1879 2796 1880
rect 2790 1875 2791 1879
rect 2795 1875 2796 1879
rect 2790 1874 2796 1875
rect 2958 1879 2964 1880
rect 2958 1875 2959 1879
rect 2963 1875 2964 1879
rect 2958 1874 2964 1875
rect 3126 1879 3132 1880
rect 3126 1875 3127 1879
rect 3131 1875 3132 1879
rect 3126 1874 3132 1875
rect 3302 1879 3308 1880
rect 3302 1875 3303 1879
rect 3307 1875 3308 1879
rect 3302 1874 3308 1875
rect 3486 1879 3492 1880
rect 3486 1875 3487 1879
rect 3491 1875 3492 1879
rect 3486 1874 3492 1875
rect 3670 1879 3676 1880
rect 3670 1875 3671 1879
rect 3675 1875 3676 1879
rect 3670 1874 3676 1875
rect 3838 1879 3844 1880
rect 3838 1875 3839 1879
rect 3843 1875 3844 1879
rect 3942 1876 3943 1880
rect 3947 1876 3948 1880
rect 3942 1875 3948 1876
rect 3838 1874 3844 1875
rect 2006 1871 2012 1872
rect 1718 1870 1724 1871
rect 2046 1863 2052 1864
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 2006 1859 2012 1860
rect 110 1854 116 1855
rect 550 1856 556 1857
rect 550 1852 551 1856
rect 555 1852 556 1856
rect 550 1851 556 1852
rect 662 1856 668 1857
rect 662 1852 663 1856
rect 667 1852 668 1856
rect 662 1851 668 1852
rect 782 1856 788 1857
rect 782 1852 783 1856
rect 787 1852 788 1856
rect 782 1851 788 1852
rect 910 1856 916 1857
rect 910 1852 911 1856
rect 915 1852 916 1856
rect 910 1851 916 1852
rect 1046 1856 1052 1857
rect 1046 1852 1047 1856
rect 1051 1852 1052 1856
rect 1046 1851 1052 1852
rect 1174 1856 1180 1857
rect 1174 1852 1175 1856
rect 1179 1852 1180 1856
rect 1174 1851 1180 1852
rect 1310 1856 1316 1857
rect 1310 1852 1311 1856
rect 1315 1852 1316 1856
rect 1310 1851 1316 1852
rect 1446 1856 1452 1857
rect 1446 1852 1447 1856
rect 1451 1852 1452 1856
rect 1446 1851 1452 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1718 1856 1724 1857
rect 1718 1852 1719 1856
rect 1723 1852 1724 1856
rect 2006 1855 2007 1859
rect 2011 1855 2012 1859
rect 2046 1859 2047 1863
rect 2051 1859 2052 1863
rect 3942 1863 3948 1864
rect 2046 1858 2052 1859
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2070 1855 2076 1856
rect 2246 1860 2252 1861
rect 2246 1856 2247 1860
rect 2251 1856 2252 1860
rect 2246 1855 2252 1856
rect 2438 1860 2444 1861
rect 2438 1856 2439 1860
rect 2443 1856 2444 1860
rect 2438 1855 2444 1856
rect 2622 1860 2628 1861
rect 2622 1856 2623 1860
rect 2627 1856 2628 1860
rect 2622 1855 2628 1856
rect 2790 1860 2796 1861
rect 2790 1856 2791 1860
rect 2795 1856 2796 1860
rect 2790 1855 2796 1856
rect 2958 1860 2964 1861
rect 2958 1856 2959 1860
rect 2963 1856 2964 1860
rect 2958 1855 2964 1856
rect 3126 1860 3132 1861
rect 3126 1856 3127 1860
rect 3131 1856 3132 1860
rect 3126 1855 3132 1856
rect 3302 1860 3308 1861
rect 3302 1856 3303 1860
rect 3307 1856 3308 1860
rect 3302 1855 3308 1856
rect 3486 1860 3492 1861
rect 3486 1856 3487 1860
rect 3491 1856 3492 1860
rect 3486 1855 3492 1856
rect 3670 1860 3676 1861
rect 3670 1856 3671 1860
rect 3675 1856 3676 1860
rect 3670 1855 3676 1856
rect 3838 1860 3844 1861
rect 3838 1856 3839 1860
rect 3843 1856 3844 1860
rect 3942 1859 3943 1863
rect 3947 1859 3948 1863
rect 3942 1858 3948 1859
rect 3838 1855 3844 1856
rect 2006 1854 2012 1855
rect 1718 1851 1724 1852
rect 2094 1800 2100 1801
rect 2046 1797 2052 1798
rect 502 1796 508 1797
rect 110 1793 116 1794
rect 110 1789 111 1793
rect 115 1789 116 1793
rect 502 1792 503 1796
rect 507 1792 508 1796
rect 502 1791 508 1792
rect 614 1796 620 1797
rect 614 1792 615 1796
rect 619 1792 620 1796
rect 614 1791 620 1792
rect 734 1796 740 1797
rect 734 1792 735 1796
rect 739 1792 740 1796
rect 734 1791 740 1792
rect 862 1796 868 1797
rect 862 1792 863 1796
rect 867 1792 868 1796
rect 862 1791 868 1792
rect 998 1796 1004 1797
rect 998 1792 999 1796
rect 1003 1792 1004 1796
rect 998 1791 1004 1792
rect 1150 1796 1156 1797
rect 1150 1792 1151 1796
rect 1155 1792 1156 1796
rect 1150 1791 1156 1792
rect 1318 1796 1324 1797
rect 1318 1792 1319 1796
rect 1323 1792 1324 1796
rect 1318 1791 1324 1792
rect 1486 1796 1492 1797
rect 1486 1792 1487 1796
rect 1491 1792 1492 1796
rect 1486 1791 1492 1792
rect 1662 1796 1668 1797
rect 1662 1792 1663 1796
rect 1667 1792 1668 1796
rect 1662 1791 1668 1792
rect 1846 1796 1852 1797
rect 1846 1792 1847 1796
rect 1851 1792 1852 1796
rect 1846 1791 1852 1792
rect 2006 1793 2012 1794
rect 110 1788 116 1789
rect 2006 1789 2007 1793
rect 2011 1789 2012 1793
rect 2046 1793 2047 1797
rect 2051 1793 2052 1797
rect 2094 1796 2095 1800
rect 2099 1796 2100 1800
rect 2094 1795 2100 1796
rect 2230 1800 2236 1801
rect 2230 1796 2231 1800
rect 2235 1796 2236 1800
rect 2230 1795 2236 1796
rect 2366 1800 2372 1801
rect 2366 1796 2367 1800
rect 2371 1796 2372 1800
rect 2366 1795 2372 1796
rect 2510 1800 2516 1801
rect 2510 1796 2511 1800
rect 2515 1796 2516 1800
rect 2510 1795 2516 1796
rect 2670 1800 2676 1801
rect 2670 1796 2671 1800
rect 2675 1796 2676 1800
rect 2670 1795 2676 1796
rect 2854 1800 2860 1801
rect 2854 1796 2855 1800
rect 2859 1796 2860 1800
rect 2854 1795 2860 1796
rect 3070 1800 3076 1801
rect 3070 1796 3071 1800
rect 3075 1796 3076 1800
rect 3070 1795 3076 1796
rect 3302 1800 3308 1801
rect 3302 1796 3303 1800
rect 3307 1796 3308 1800
rect 3302 1795 3308 1796
rect 3542 1800 3548 1801
rect 3542 1796 3543 1800
rect 3547 1796 3548 1800
rect 3542 1795 3548 1796
rect 3790 1800 3796 1801
rect 3790 1796 3791 1800
rect 3795 1796 3796 1800
rect 3790 1795 3796 1796
rect 3942 1797 3948 1798
rect 2046 1792 2052 1793
rect 3942 1793 3943 1797
rect 3947 1793 3948 1797
rect 3942 1792 3948 1793
rect 2006 1788 2012 1789
rect 2094 1781 2100 1782
rect 2046 1780 2052 1781
rect 502 1777 508 1778
rect 110 1776 116 1777
rect 110 1772 111 1776
rect 115 1772 116 1776
rect 502 1773 503 1777
rect 507 1773 508 1777
rect 502 1772 508 1773
rect 614 1777 620 1778
rect 614 1773 615 1777
rect 619 1773 620 1777
rect 614 1772 620 1773
rect 734 1777 740 1778
rect 734 1773 735 1777
rect 739 1773 740 1777
rect 734 1772 740 1773
rect 862 1777 868 1778
rect 862 1773 863 1777
rect 867 1773 868 1777
rect 862 1772 868 1773
rect 998 1777 1004 1778
rect 998 1773 999 1777
rect 1003 1773 1004 1777
rect 998 1772 1004 1773
rect 1150 1777 1156 1778
rect 1150 1773 1151 1777
rect 1155 1773 1156 1777
rect 1150 1772 1156 1773
rect 1318 1777 1324 1778
rect 1318 1773 1319 1777
rect 1323 1773 1324 1777
rect 1318 1772 1324 1773
rect 1486 1777 1492 1778
rect 1486 1773 1487 1777
rect 1491 1773 1492 1777
rect 1486 1772 1492 1773
rect 1662 1777 1668 1778
rect 1662 1773 1663 1777
rect 1667 1773 1668 1777
rect 1662 1772 1668 1773
rect 1846 1777 1852 1778
rect 1846 1773 1847 1777
rect 1851 1773 1852 1777
rect 1846 1772 1852 1773
rect 2006 1776 2012 1777
rect 2006 1772 2007 1776
rect 2011 1772 2012 1776
rect 2046 1776 2047 1780
rect 2051 1776 2052 1780
rect 2094 1777 2095 1781
rect 2099 1777 2100 1781
rect 2094 1776 2100 1777
rect 2230 1781 2236 1782
rect 2230 1777 2231 1781
rect 2235 1777 2236 1781
rect 2230 1776 2236 1777
rect 2366 1781 2372 1782
rect 2366 1777 2367 1781
rect 2371 1777 2372 1781
rect 2366 1776 2372 1777
rect 2510 1781 2516 1782
rect 2510 1777 2511 1781
rect 2515 1777 2516 1781
rect 2510 1776 2516 1777
rect 2670 1781 2676 1782
rect 2670 1777 2671 1781
rect 2675 1777 2676 1781
rect 2670 1776 2676 1777
rect 2854 1781 2860 1782
rect 2854 1777 2855 1781
rect 2859 1777 2860 1781
rect 2854 1776 2860 1777
rect 3070 1781 3076 1782
rect 3070 1777 3071 1781
rect 3075 1777 3076 1781
rect 3070 1776 3076 1777
rect 3302 1781 3308 1782
rect 3302 1777 3303 1781
rect 3307 1777 3308 1781
rect 3302 1776 3308 1777
rect 3542 1781 3548 1782
rect 3542 1777 3543 1781
rect 3547 1777 3548 1781
rect 3542 1776 3548 1777
rect 3790 1781 3796 1782
rect 3790 1777 3791 1781
rect 3795 1777 3796 1781
rect 3790 1776 3796 1777
rect 3942 1780 3948 1781
rect 3942 1776 3943 1780
rect 3947 1776 3948 1780
rect 2046 1775 2052 1776
rect 3942 1775 3948 1776
rect 110 1771 116 1772
rect 2006 1771 2012 1772
rect 2046 1728 2052 1729
rect 3942 1728 3948 1729
rect 110 1724 116 1725
rect 2006 1724 2012 1725
rect 110 1720 111 1724
rect 115 1720 116 1724
rect 110 1719 116 1720
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1719 348 1723
rect 342 1718 348 1719
rect 462 1723 468 1724
rect 462 1719 463 1723
rect 467 1719 468 1723
rect 462 1718 468 1719
rect 590 1723 596 1724
rect 590 1719 591 1723
rect 595 1719 596 1723
rect 590 1718 596 1719
rect 718 1723 724 1724
rect 718 1719 719 1723
rect 723 1719 724 1723
rect 718 1718 724 1719
rect 846 1723 852 1724
rect 846 1719 847 1723
rect 851 1719 852 1723
rect 846 1718 852 1719
rect 982 1723 988 1724
rect 982 1719 983 1723
rect 987 1719 988 1723
rect 982 1718 988 1719
rect 1126 1723 1132 1724
rect 1126 1719 1127 1723
rect 1131 1719 1132 1723
rect 1126 1718 1132 1719
rect 1278 1723 1284 1724
rect 1278 1719 1279 1723
rect 1283 1719 1284 1723
rect 1278 1718 1284 1719
rect 1438 1723 1444 1724
rect 1438 1719 1439 1723
rect 1443 1719 1444 1723
rect 1438 1718 1444 1719
rect 1598 1723 1604 1724
rect 1598 1719 1599 1723
rect 1603 1719 1604 1723
rect 2006 1720 2007 1724
rect 2011 1720 2012 1724
rect 2046 1724 2047 1728
rect 2051 1724 2052 1728
rect 2046 1723 2052 1724
rect 2182 1727 2188 1728
rect 2182 1723 2183 1727
rect 2187 1723 2188 1727
rect 2182 1722 2188 1723
rect 2286 1727 2292 1728
rect 2286 1723 2287 1727
rect 2291 1723 2292 1727
rect 2286 1722 2292 1723
rect 2390 1727 2396 1728
rect 2390 1723 2391 1727
rect 2395 1723 2396 1727
rect 2390 1722 2396 1723
rect 2494 1727 2500 1728
rect 2494 1723 2495 1727
rect 2499 1723 2500 1727
rect 2494 1722 2500 1723
rect 2598 1727 2604 1728
rect 2598 1723 2599 1727
rect 2603 1723 2604 1727
rect 2598 1722 2604 1723
rect 2702 1727 2708 1728
rect 2702 1723 2703 1727
rect 2707 1723 2708 1727
rect 2702 1722 2708 1723
rect 2806 1727 2812 1728
rect 2806 1723 2807 1727
rect 2811 1723 2812 1727
rect 2806 1722 2812 1723
rect 2910 1727 2916 1728
rect 2910 1723 2911 1727
rect 2915 1723 2916 1727
rect 2910 1722 2916 1723
rect 3014 1727 3020 1728
rect 3014 1723 3015 1727
rect 3019 1723 3020 1727
rect 3014 1722 3020 1723
rect 3126 1727 3132 1728
rect 3126 1723 3127 1727
rect 3131 1723 3132 1727
rect 3942 1724 3943 1728
rect 3947 1724 3948 1728
rect 3942 1723 3948 1724
rect 3126 1722 3132 1723
rect 2006 1719 2012 1720
rect 1598 1718 1604 1719
rect 2046 1711 2052 1712
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 2006 1707 2012 1708
rect 110 1702 116 1703
rect 342 1704 348 1705
rect 342 1700 343 1704
rect 347 1700 348 1704
rect 342 1699 348 1700
rect 462 1704 468 1705
rect 462 1700 463 1704
rect 467 1700 468 1704
rect 462 1699 468 1700
rect 590 1704 596 1705
rect 590 1700 591 1704
rect 595 1700 596 1704
rect 590 1699 596 1700
rect 718 1704 724 1705
rect 718 1700 719 1704
rect 723 1700 724 1704
rect 718 1699 724 1700
rect 846 1704 852 1705
rect 846 1700 847 1704
rect 851 1700 852 1704
rect 846 1699 852 1700
rect 982 1704 988 1705
rect 982 1700 983 1704
rect 987 1700 988 1704
rect 982 1699 988 1700
rect 1126 1704 1132 1705
rect 1126 1700 1127 1704
rect 1131 1700 1132 1704
rect 1126 1699 1132 1700
rect 1278 1704 1284 1705
rect 1278 1700 1279 1704
rect 1283 1700 1284 1704
rect 1278 1699 1284 1700
rect 1438 1704 1444 1705
rect 1438 1700 1439 1704
rect 1443 1700 1444 1704
rect 1438 1699 1444 1700
rect 1598 1704 1604 1705
rect 1598 1700 1599 1704
rect 1603 1700 1604 1704
rect 2006 1703 2007 1707
rect 2011 1703 2012 1707
rect 2046 1707 2047 1711
rect 2051 1707 2052 1711
rect 3942 1711 3948 1712
rect 2046 1706 2052 1707
rect 2182 1708 2188 1709
rect 2182 1704 2183 1708
rect 2187 1704 2188 1708
rect 2182 1703 2188 1704
rect 2286 1708 2292 1709
rect 2286 1704 2287 1708
rect 2291 1704 2292 1708
rect 2286 1703 2292 1704
rect 2390 1708 2396 1709
rect 2390 1704 2391 1708
rect 2395 1704 2396 1708
rect 2390 1703 2396 1704
rect 2494 1708 2500 1709
rect 2494 1704 2495 1708
rect 2499 1704 2500 1708
rect 2494 1703 2500 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2702 1708 2708 1709
rect 2702 1704 2703 1708
rect 2707 1704 2708 1708
rect 2702 1703 2708 1704
rect 2806 1708 2812 1709
rect 2806 1704 2807 1708
rect 2811 1704 2812 1708
rect 2806 1703 2812 1704
rect 2910 1708 2916 1709
rect 2910 1704 2911 1708
rect 2915 1704 2916 1708
rect 2910 1703 2916 1704
rect 3014 1708 3020 1709
rect 3014 1704 3015 1708
rect 3019 1704 3020 1708
rect 3014 1703 3020 1704
rect 3126 1708 3132 1709
rect 3126 1704 3127 1708
rect 3131 1704 3132 1708
rect 3942 1707 3943 1711
rect 3947 1707 3948 1711
rect 3942 1706 3948 1707
rect 3126 1703 3132 1704
rect 2006 1702 2012 1703
rect 1598 1699 1604 1700
rect 2230 1648 2236 1649
rect 2046 1645 2052 1646
rect 2046 1641 2047 1645
rect 2051 1641 2052 1645
rect 2230 1644 2231 1648
rect 2235 1644 2236 1648
rect 2230 1643 2236 1644
rect 2366 1648 2372 1649
rect 2366 1644 2367 1648
rect 2371 1644 2372 1648
rect 2366 1643 2372 1644
rect 2518 1648 2524 1649
rect 2518 1644 2519 1648
rect 2523 1644 2524 1648
rect 2518 1643 2524 1644
rect 2678 1648 2684 1649
rect 2678 1644 2679 1648
rect 2683 1644 2684 1648
rect 2678 1643 2684 1644
rect 2846 1648 2852 1649
rect 2846 1644 2847 1648
rect 2851 1644 2852 1648
rect 2846 1643 2852 1644
rect 3022 1648 3028 1649
rect 3022 1644 3023 1648
rect 3027 1644 3028 1648
rect 3022 1643 3028 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3526 1648 3532 1649
rect 3526 1644 3527 1648
rect 3531 1644 3532 1648
rect 3526 1643 3532 1644
rect 3694 1648 3700 1649
rect 3694 1644 3695 1648
rect 3699 1644 3700 1648
rect 3694 1643 3700 1644
rect 3838 1648 3844 1649
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3838 1643 3844 1644
rect 3942 1645 3948 1646
rect 158 1640 164 1641
rect 110 1637 116 1638
rect 110 1633 111 1637
rect 115 1633 116 1637
rect 158 1636 159 1640
rect 163 1636 164 1640
rect 158 1635 164 1636
rect 294 1640 300 1641
rect 294 1636 295 1640
rect 299 1636 300 1640
rect 294 1635 300 1636
rect 454 1640 460 1641
rect 454 1636 455 1640
rect 459 1636 460 1640
rect 454 1635 460 1636
rect 622 1640 628 1641
rect 622 1636 623 1640
rect 627 1636 628 1640
rect 622 1635 628 1636
rect 798 1640 804 1641
rect 798 1636 799 1640
rect 803 1636 804 1640
rect 798 1635 804 1636
rect 982 1640 988 1641
rect 982 1636 983 1640
rect 987 1636 988 1640
rect 982 1635 988 1636
rect 1166 1640 1172 1641
rect 1166 1636 1167 1640
rect 1171 1636 1172 1640
rect 1166 1635 1172 1636
rect 1350 1640 1356 1641
rect 1350 1636 1351 1640
rect 1355 1636 1356 1640
rect 1350 1635 1356 1636
rect 1542 1640 1548 1641
rect 1542 1636 1543 1640
rect 1547 1636 1548 1640
rect 1542 1635 1548 1636
rect 1734 1640 1740 1641
rect 2046 1640 2052 1641
rect 3942 1641 3943 1645
rect 3947 1641 3948 1645
rect 3942 1640 3948 1641
rect 1734 1636 1735 1640
rect 1739 1636 1740 1640
rect 1734 1635 1740 1636
rect 2006 1637 2012 1638
rect 110 1632 116 1633
rect 2006 1633 2007 1637
rect 2011 1633 2012 1637
rect 2006 1632 2012 1633
rect 2230 1629 2236 1630
rect 2046 1628 2052 1629
rect 2046 1624 2047 1628
rect 2051 1624 2052 1628
rect 2230 1625 2231 1629
rect 2235 1625 2236 1629
rect 2230 1624 2236 1625
rect 2366 1629 2372 1630
rect 2366 1625 2367 1629
rect 2371 1625 2372 1629
rect 2366 1624 2372 1625
rect 2518 1629 2524 1630
rect 2518 1625 2519 1629
rect 2523 1625 2524 1629
rect 2518 1624 2524 1625
rect 2678 1629 2684 1630
rect 2678 1625 2679 1629
rect 2683 1625 2684 1629
rect 2678 1624 2684 1625
rect 2846 1629 2852 1630
rect 2846 1625 2847 1629
rect 2851 1625 2852 1629
rect 2846 1624 2852 1625
rect 3022 1629 3028 1630
rect 3022 1625 3023 1629
rect 3027 1625 3028 1629
rect 3022 1624 3028 1625
rect 3190 1629 3196 1630
rect 3190 1625 3191 1629
rect 3195 1625 3196 1629
rect 3190 1624 3196 1625
rect 3358 1629 3364 1630
rect 3358 1625 3359 1629
rect 3363 1625 3364 1629
rect 3358 1624 3364 1625
rect 3526 1629 3532 1630
rect 3526 1625 3527 1629
rect 3531 1625 3532 1629
rect 3526 1624 3532 1625
rect 3694 1629 3700 1630
rect 3694 1625 3695 1629
rect 3699 1625 3700 1629
rect 3694 1624 3700 1625
rect 3838 1629 3844 1630
rect 3838 1625 3839 1629
rect 3843 1625 3844 1629
rect 3838 1624 3844 1625
rect 3942 1628 3948 1629
rect 3942 1624 3943 1628
rect 3947 1624 3948 1628
rect 2046 1623 2052 1624
rect 3942 1623 3948 1624
rect 158 1621 164 1622
rect 110 1620 116 1621
rect 110 1616 111 1620
rect 115 1616 116 1620
rect 158 1617 159 1621
rect 163 1617 164 1621
rect 158 1616 164 1617
rect 294 1621 300 1622
rect 294 1617 295 1621
rect 299 1617 300 1621
rect 294 1616 300 1617
rect 454 1621 460 1622
rect 454 1617 455 1621
rect 459 1617 460 1621
rect 454 1616 460 1617
rect 622 1621 628 1622
rect 622 1617 623 1621
rect 627 1617 628 1621
rect 622 1616 628 1617
rect 798 1621 804 1622
rect 798 1617 799 1621
rect 803 1617 804 1621
rect 798 1616 804 1617
rect 982 1621 988 1622
rect 982 1617 983 1621
rect 987 1617 988 1621
rect 982 1616 988 1617
rect 1166 1621 1172 1622
rect 1166 1617 1167 1621
rect 1171 1617 1172 1621
rect 1166 1616 1172 1617
rect 1350 1621 1356 1622
rect 1350 1617 1351 1621
rect 1355 1617 1356 1621
rect 1350 1616 1356 1617
rect 1542 1621 1548 1622
rect 1542 1617 1543 1621
rect 1547 1617 1548 1621
rect 1542 1616 1548 1617
rect 1734 1621 1740 1622
rect 1734 1617 1735 1621
rect 1739 1617 1740 1621
rect 1734 1616 1740 1617
rect 2006 1620 2012 1621
rect 2006 1616 2007 1620
rect 2011 1616 2012 1620
rect 110 1615 116 1616
rect 2006 1615 2012 1616
rect 110 1568 116 1569
rect 2006 1568 2012 1569
rect 110 1564 111 1568
rect 115 1564 116 1568
rect 110 1563 116 1564
rect 134 1567 140 1568
rect 134 1563 135 1567
rect 139 1563 140 1567
rect 134 1562 140 1563
rect 254 1567 260 1568
rect 254 1563 255 1567
rect 259 1563 260 1567
rect 254 1562 260 1563
rect 422 1567 428 1568
rect 422 1563 423 1567
rect 427 1563 428 1567
rect 422 1562 428 1563
rect 606 1567 612 1568
rect 606 1563 607 1567
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 798 1567 804 1568
rect 798 1563 799 1567
rect 803 1563 804 1567
rect 798 1562 804 1563
rect 990 1567 996 1568
rect 990 1563 991 1567
rect 995 1563 996 1567
rect 990 1562 996 1563
rect 1182 1567 1188 1568
rect 1182 1563 1183 1567
rect 1187 1563 1188 1567
rect 1182 1562 1188 1563
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 1550 1567 1556 1568
rect 1550 1563 1551 1567
rect 1555 1563 1556 1567
rect 1550 1562 1556 1563
rect 1734 1567 1740 1568
rect 1734 1563 1735 1567
rect 1739 1563 1740 1567
rect 1734 1562 1740 1563
rect 1902 1567 1908 1568
rect 1902 1563 1903 1567
rect 1907 1563 1908 1567
rect 2006 1564 2007 1568
rect 2011 1564 2012 1568
rect 2006 1563 2012 1564
rect 2046 1568 2052 1569
rect 3942 1568 3948 1569
rect 2046 1564 2047 1568
rect 2051 1564 2052 1568
rect 2046 1563 2052 1564
rect 2070 1567 2076 1568
rect 2070 1563 2071 1567
rect 2075 1563 2076 1567
rect 1902 1562 1908 1563
rect 2070 1562 2076 1563
rect 2270 1567 2276 1568
rect 2270 1563 2271 1567
rect 2275 1563 2276 1567
rect 2270 1562 2276 1563
rect 2494 1567 2500 1568
rect 2494 1563 2495 1567
rect 2499 1563 2500 1567
rect 2494 1562 2500 1563
rect 2710 1567 2716 1568
rect 2710 1563 2711 1567
rect 2715 1563 2716 1567
rect 2710 1562 2716 1563
rect 2910 1567 2916 1568
rect 2910 1563 2911 1567
rect 2915 1563 2916 1567
rect 2910 1562 2916 1563
rect 3094 1567 3100 1568
rect 3094 1563 3095 1567
rect 3099 1563 3100 1567
rect 3094 1562 3100 1563
rect 3262 1567 3268 1568
rect 3262 1563 3263 1567
rect 3267 1563 3268 1567
rect 3262 1562 3268 1563
rect 3422 1567 3428 1568
rect 3422 1563 3423 1567
rect 3427 1563 3428 1567
rect 3422 1562 3428 1563
rect 3566 1567 3572 1568
rect 3566 1563 3567 1567
rect 3571 1563 3572 1567
rect 3566 1562 3572 1563
rect 3710 1567 3716 1568
rect 3710 1563 3711 1567
rect 3715 1563 3716 1567
rect 3710 1562 3716 1563
rect 3838 1567 3844 1568
rect 3838 1563 3839 1567
rect 3843 1563 3844 1567
rect 3942 1564 3943 1568
rect 3947 1564 3948 1568
rect 3942 1563 3948 1564
rect 3838 1562 3844 1563
rect 110 1551 116 1552
rect 110 1547 111 1551
rect 115 1547 116 1551
rect 2006 1551 2012 1552
rect 110 1546 116 1547
rect 134 1548 140 1549
rect 134 1544 135 1548
rect 139 1544 140 1548
rect 134 1543 140 1544
rect 254 1548 260 1549
rect 254 1544 255 1548
rect 259 1544 260 1548
rect 254 1543 260 1544
rect 422 1548 428 1549
rect 422 1544 423 1548
rect 427 1544 428 1548
rect 422 1543 428 1544
rect 606 1548 612 1549
rect 606 1544 607 1548
rect 611 1544 612 1548
rect 606 1543 612 1544
rect 798 1548 804 1549
rect 798 1544 799 1548
rect 803 1544 804 1548
rect 798 1543 804 1544
rect 990 1548 996 1549
rect 990 1544 991 1548
rect 995 1544 996 1548
rect 990 1543 996 1544
rect 1182 1548 1188 1549
rect 1182 1544 1183 1548
rect 1187 1544 1188 1548
rect 1182 1543 1188 1544
rect 1366 1548 1372 1549
rect 1366 1544 1367 1548
rect 1371 1544 1372 1548
rect 1366 1543 1372 1544
rect 1550 1548 1556 1549
rect 1550 1544 1551 1548
rect 1555 1544 1556 1548
rect 1550 1543 1556 1544
rect 1734 1548 1740 1549
rect 1734 1544 1735 1548
rect 1739 1544 1740 1548
rect 1734 1543 1740 1544
rect 1902 1548 1908 1549
rect 1902 1544 1903 1548
rect 1907 1544 1908 1548
rect 2006 1547 2007 1551
rect 2011 1547 2012 1551
rect 2006 1546 2012 1547
rect 2046 1551 2052 1552
rect 2046 1547 2047 1551
rect 2051 1547 2052 1551
rect 3942 1551 3948 1552
rect 2046 1546 2052 1547
rect 2070 1548 2076 1549
rect 1902 1543 1908 1544
rect 2070 1544 2071 1548
rect 2075 1544 2076 1548
rect 2070 1543 2076 1544
rect 2270 1548 2276 1549
rect 2270 1544 2271 1548
rect 2275 1544 2276 1548
rect 2270 1543 2276 1544
rect 2494 1548 2500 1549
rect 2494 1544 2495 1548
rect 2499 1544 2500 1548
rect 2494 1543 2500 1544
rect 2710 1548 2716 1549
rect 2710 1544 2711 1548
rect 2715 1544 2716 1548
rect 2710 1543 2716 1544
rect 2910 1548 2916 1549
rect 2910 1544 2911 1548
rect 2915 1544 2916 1548
rect 2910 1543 2916 1544
rect 3094 1548 3100 1549
rect 3094 1544 3095 1548
rect 3099 1544 3100 1548
rect 3094 1543 3100 1544
rect 3262 1548 3268 1549
rect 3262 1544 3263 1548
rect 3267 1544 3268 1548
rect 3262 1543 3268 1544
rect 3422 1548 3428 1549
rect 3422 1544 3423 1548
rect 3427 1544 3428 1548
rect 3422 1543 3428 1544
rect 3566 1548 3572 1549
rect 3566 1544 3567 1548
rect 3571 1544 3572 1548
rect 3566 1543 3572 1544
rect 3710 1548 3716 1549
rect 3710 1544 3711 1548
rect 3715 1544 3716 1548
rect 3710 1543 3716 1544
rect 3838 1548 3844 1549
rect 3838 1544 3839 1548
rect 3843 1544 3844 1548
rect 3942 1547 3943 1551
rect 3947 1547 3948 1551
rect 3942 1546 3948 1547
rect 3838 1543 3844 1544
rect 2070 1488 2076 1489
rect 2046 1485 2052 1486
rect 134 1484 140 1485
rect 110 1481 116 1482
rect 110 1477 111 1481
rect 115 1477 116 1481
rect 134 1480 135 1484
rect 139 1480 140 1484
rect 134 1479 140 1480
rect 246 1484 252 1485
rect 246 1480 247 1484
rect 251 1480 252 1484
rect 246 1479 252 1480
rect 398 1484 404 1485
rect 398 1480 399 1484
rect 403 1480 404 1484
rect 398 1479 404 1480
rect 558 1484 564 1485
rect 558 1480 559 1484
rect 563 1480 564 1484
rect 558 1479 564 1480
rect 718 1484 724 1485
rect 718 1480 719 1484
rect 723 1480 724 1484
rect 718 1479 724 1480
rect 878 1484 884 1485
rect 878 1480 879 1484
rect 883 1480 884 1484
rect 878 1479 884 1480
rect 1038 1484 1044 1485
rect 1038 1480 1039 1484
rect 1043 1480 1044 1484
rect 1038 1479 1044 1480
rect 1182 1484 1188 1485
rect 1182 1480 1183 1484
rect 1187 1480 1188 1484
rect 1182 1479 1188 1480
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1446 1484 1452 1485
rect 1446 1480 1447 1484
rect 1451 1480 1452 1484
rect 1446 1479 1452 1480
rect 1566 1484 1572 1485
rect 1566 1480 1567 1484
rect 1571 1480 1572 1484
rect 1566 1479 1572 1480
rect 1686 1484 1692 1485
rect 1686 1480 1687 1484
rect 1691 1480 1692 1484
rect 1686 1479 1692 1480
rect 1806 1484 1812 1485
rect 1806 1480 1807 1484
rect 1811 1480 1812 1484
rect 1806 1479 1812 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 2006 1481 2012 1482
rect 110 1476 116 1477
rect 2006 1477 2007 1481
rect 2011 1477 2012 1481
rect 2046 1481 2047 1485
rect 2051 1481 2052 1485
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 2430 1488 2436 1489
rect 2430 1484 2431 1488
rect 2435 1484 2436 1488
rect 2430 1483 2436 1484
rect 2790 1488 2796 1489
rect 2790 1484 2791 1488
rect 2795 1484 2796 1488
rect 2790 1483 2796 1484
rect 3126 1488 3132 1489
rect 3126 1484 3127 1488
rect 3131 1484 3132 1488
rect 3126 1483 3132 1484
rect 3462 1488 3468 1489
rect 3462 1484 3463 1488
rect 3467 1484 3468 1488
rect 3462 1483 3468 1484
rect 3798 1488 3804 1489
rect 3798 1484 3799 1488
rect 3803 1484 3804 1488
rect 3798 1483 3804 1484
rect 3942 1485 3948 1486
rect 2046 1480 2052 1481
rect 3942 1481 3943 1485
rect 3947 1481 3948 1485
rect 3942 1480 3948 1481
rect 2006 1476 2012 1477
rect 2070 1469 2076 1470
rect 2046 1468 2052 1469
rect 134 1465 140 1466
rect 110 1464 116 1465
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 134 1461 135 1465
rect 139 1461 140 1465
rect 134 1460 140 1461
rect 246 1465 252 1466
rect 246 1461 247 1465
rect 251 1461 252 1465
rect 246 1460 252 1461
rect 398 1465 404 1466
rect 398 1461 399 1465
rect 403 1461 404 1465
rect 398 1460 404 1461
rect 558 1465 564 1466
rect 558 1461 559 1465
rect 563 1461 564 1465
rect 558 1460 564 1461
rect 718 1465 724 1466
rect 718 1461 719 1465
rect 723 1461 724 1465
rect 718 1460 724 1461
rect 878 1465 884 1466
rect 878 1461 879 1465
rect 883 1461 884 1465
rect 878 1460 884 1461
rect 1038 1465 1044 1466
rect 1038 1461 1039 1465
rect 1043 1461 1044 1465
rect 1038 1460 1044 1461
rect 1182 1465 1188 1466
rect 1182 1461 1183 1465
rect 1187 1461 1188 1465
rect 1182 1460 1188 1461
rect 1318 1465 1324 1466
rect 1318 1461 1319 1465
rect 1323 1461 1324 1465
rect 1318 1460 1324 1461
rect 1446 1465 1452 1466
rect 1446 1461 1447 1465
rect 1451 1461 1452 1465
rect 1446 1460 1452 1461
rect 1566 1465 1572 1466
rect 1566 1461 1567 1465
rect 1571 1461 1572 1465
rect 1566 1460 1572 1461
rect 1686 1465 1692 1466
rect 1686 1461 1687 1465
rect 1691 1461 1692 1465
rect 1686 1460 1692 1461
rect 1806 1465 1812 1466
rect 1806 1461 1807 1465
rect 1811 1461 1812 1465
rect 1806 1460 1812 1461
rect 1902 1465 1908 1466
rect 1902 1461 1903 1465
rect 1907 1461 1908 1465
rect 1902 1460 1908 1461
rect 2006 1464 2012 1465
rect 2006 1460 2007 1464
rect 2011 1460 2012 1464
rect 2046 1464 2047 1468
rect 2051 1464 2052 1468
rect 2070 1465 2071 1469
rect 2075 1465 2076 1469
rect 2070 1464 2076 1465
rect 2430 1469 2436 1470
rect 2430 1465 2431 1469
rect 2435 1465 2436 1469
rect 2430 1464 2436 1465
rect 2790 1469 2796 1470
rect 2790 1465 2791 1469
rect 2795 1465 2796 1469
rect 2790 1464 2796 1465
rect 3126 1469 3132 1470
rect 3126 1465 3127 1469
rect 3131 1465 3132 1469
rect 3126 1464 3132 1465
rect 3462 1469 3468 1470
rect 3462 1465 3463 1469
rect 3467 1465 3468 1469
rect 3462 1464 3468 1465
rect 3798 1469 3804 1470
rect 3798 1465 3799 1469
rect 3803 1465 3804 1469
rect 3798 1464 3804 1465
rect 3942 1468 3948 1469
rect 3942 1464 3943 1468
rect 3947 1464 3948 1468
rect 2046 1463 2052 1464
rect 3942 1463 3948 1464
rect 110 1459 116 1460
rect 2006 1459 2012 1460
rect 110 1412 116 1413
rect 2006 1412 2012 1413
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 110 1407 116 1408
rect 134 1411 140 1412
rect 134 1407 135 1411
rect 139 1407 140 1411
rect 134 1406 140 1407
rect 262 1411 268 1412
rect 262 1407 263 1411
rect 267 1407 268 1411
rect 262 1406 268 1407
rect 430 1411 436 1412
rect 430 1407 431 1411
rect 435 1407 436 1411
rect 430 1406 436 1407
rect 606 1411 612 1412
rect 606 1407 607 1411
rect 611 1407 612 1411
rect 606 1406 612 1407
rect 790 1411 796 1412
rect 790 1407 791 1411
rect 795 1407 796 1411
rect 790 1406 796 1407
rect 974 1411 980 1412
rect 974 1407 975 1411
rect 979 1407 980 1411
rect 974 1406 980 1407
rect 1158 1411 1164 1412
rect 1158 1407 1159 1411
rect 1163 1407 1164 1411
rect 1158 1406 1164 1407
rect 1350 1411 1356 1412
rect 1350 1407 1351 1411
rect 1355 1407 1356 1411
rect 1350 1406 1356 1407
rect 1542 1411 1548 1412
rect 1542 1407 1543 1411
rect 1547 1407 1548 1411
rect 1542 1406 1548 1407
rect 1734 1411 1740 1412
rect 1734 1407 1735 1411
rect 1739 1407 1740 1411
rect 1734 1406 1740 1407
rect 1902 1411 1908 1412
rect 1902 1407 1903 1411
rect 1907 1407 1908 1411
rect 2006 1408 2007 1412
rect 2011 1408 2012 1412
rect 2006 1407 2012 1408
rect 2046 1408 2052 1409
rect 3942 1408 3948 1409
rect 1902 1406 1908 1407
rect 2046 1404 2047 1408
rect 2051 1404 2052 1408
rect 2046 1403 2052 1404
rect 2070 1407 2076 1408
rect 2070 1403 2071 1407
rect 2075 1403 2076 1407
rect 2070 1402 2076 1403
rect 2270 1407 2276 1408
rect 2270 1403 2271 1407
rect 2275 1403 2276 1407
rect 2270 1402 2276 1403
rect 2494 1407 2500 1408
rect 2494 1403 2495 1407
rect 2499 1403 2500 1407
rect 2494 1402 2500 1403
rect 2710 1407 2716 1408
rect 2710 1403 2711 1407
rect 2715 1403 2716 1407
rect 2710 1402 2716 1403
rect 2910 1407 2916 1408
rect 2910 1403 2911 1407
rect 2915 1403 2916 1407
rect 2910 1402 2916 1403
rect 3094 1407 3100 1408
rect 3094 1403 3095 1407
rect 3099 1403 3100 1407
rect 3094 1402 3100 1403
rect 3270 1407 3276 1408
rect 3270 1403 3271 1407
rect 3275 1403 3276 1407
rect 3270 1402 3276 1403
rect 3438 1407 3444 1408
rect 3438 1403 3439 1407
rect 3443 1403 3444 1407
rect 3438 1402 3444 1403
rect 3606 1407 3612 1408
rect 3606 1403 3607 1407
rect 3611 1403 3612 1407
rect 3606 1402 3612 1403
rect 3782 1407 3788 1408
rect 3782 1403 3783 1407
rect 3787 1403 3788 1407
rect 3942 1404 3943 1408
rect 3947 1404 3948 1408
rect 3942 1403 3948 1404
rect 3782 1402 3788 1403
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 2006 1395 2012 1396
rect 110 1390 116 1391
rect 134 1392 140 1393
rect 134 1388 135 1392
rect 139 1388 140 1392
rect 134 1387 140 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 430 1392 436 1393
rect 430 1388 431 1392
rect 435 1388 436 1392
rect 430 1387 436 1388
rect 606 1392 612 1393
rect 606 1388 607 1392
rect 611 1388 612 1392
rect 606 1387 612 1388
rect 790 1392 796 1393
rect 790 1388 791 1392
rect 795 1388 796 1392
rect 790 1387 796 1388
rect 974 1392 980 1393
rect 974 1388 975 1392
rect 979 1388 980 1392
rect 974 1387 980 1388
rect 1158 1392 1164 1393
rect 1158 1388 1159 1392
rect 1163 1388 1164 1392
rect 1158 1387 1164 1388
rect 1350 1392 1356 1393
rect 1350 1388 1351 1392
rect 1355 1388 1356 1392
rect 1350 1387 1356 1388
rect 1542 1392 1548 1393
rect 1542 1388 1543 1392
rect 1547 1388 1548 1392
rect 1542 1387 1548 1388
rect 1734 1392 1740 1393
rect 1734 1388 1735 1392
rect 1739 1388 1740 1392
rect 1734 1387 1740 1388
rect 1902 1392 1908 1393
rect 1902 1388 1903 1392
rect 1907 1388 1908 1392
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2006 1390 2012 1391
rect 2046 1391 2052 1392
rect 1902 1387 1908 1388
rect 2046 1387 2047 1391
rect 2051 1387 2052 1391
rect 3942 1391 3948 1392
rect 2046 1386 2052 1387
rect 2070 1388 2076 1389
rect 2070 1384 2071 1388
rect 2075 1384 2076 1388
rect 2070 1383 2076 1384
rect 2270 1388 2276 1389
rect 2270 1384 2271 1388
rect 2275 1384 2276 1388
rect 2270 1383 2276 1384
rect 2494 1388 2500 1389
rect 2494 1384 2495 1388
rect 2499 1384 2500 1388
rect 2494 1383 2500 1384
rect 2710 1388 2716 1389
rect 2710 1384 2711 1388
rect 2715 1384 2716 1388
rect 2710 1383 2716 1384
rect 2910 1388 2916 1389
rect 2910 1384 2911 1388
rect 2915 1384 2916 1388
rect 2910 1383 2916 1384
rect 3094 1388 3100 1389
rect 3094 1384 3095 1388
rect 3099 1384 3100 1388
rect 3094 1383 3100 1384
rect 3270 1388 3276 1389
rect 3270 1384 3271 1388
rect 3275 1384 3276 1388
rect 3270 1383 3276 1384
rect 3438 1388 3444 1389
rect 3438 1384 3439 1388
rect 3443 1384 3444 1388
rect 3438 1383 3444 1384
rect 3606 1388 3612 1389
rect 3606 1384 3607 1388
rect 3611 1384 3612 1388
rect 3606 1383 3612 1384
rect 3782 1388 3788 1389
rect 3782 1384 3783 1388
rect 3787 1384 3788 1388
rect 3942 1387 3943 1391
rect 3947 1387 3948 1391
rect 3942 1386 3948 1387
rect 3782 1383 3788 1384
rect 158 1328 164 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 158 1324 159 1328
rect 163 1324 164 1328
rect 158 1323 164 1324
rect 310 1328 316 1329
rect 310 1324 311 1328
rect 315 1324 316 1328
rect 310 1323 316 1324
rect 478 1328 484 1329
rect 478 1324 479 1328
rect 483 1324 484 1328
rect 478 1323 484 1324
rect 662 1328 668 1329
rect 662 1324 663 1328
rect 667 1324 668 1328
rect 662 1323 668 1324
rect 854 1328 860 1329
rect 854 1324 855 1328
rect 859 1324 860 1328
rect 854 1323 860 1324
rect 1046 1328 1052 1329
rect 1046 1324 1047 1328
rect 1051 1324 1052 1328
rect 1046 1323 1052 1324
rect 1246 1328 1252 1329
rect 1246 1324 1247 1328
rect 1251 1324 1252 1328
rect 1246 1323 1252 1324
rect 1446 1328 1452 1329
rect 1446 1324 1447 1328
rect 1451 1324 1452 1328
rect 1446 1323 1452 1324
rect 1654 1328 1660 1329
rect 1654 1324 1655 1328
rect 1659 1324 1660 1328
rect 1654 1323 1660 1324
rect 1862 1328 1868 1329
rect 1862 1324 1863 1328
rect 1867 1324 1868 1328
rect 2070 1328 2076 1329
rect 1862 1323 1868 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2046 1325 2052 1326
rect 2046 1321 2047 1325
rect 2051 1321 2052 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2206 1328 2212 1329
rect 2206 1324 2207 1328
rect 2211 1324 2212 1328
rect 2206 1323 2212 1324
rect 2382 1328 2388 1329
rect 2382 1324 2383 1328
rect 2387 1324 2388 1328
rect 2382 1323 2388 1324
rect 2566 1328 2572 1329
rect 2566 1324 2567 1328
rect 2571 1324 2572 1328
rect 2566 1323 2572 1324
rect 2750 1328 2756 1329
rect 2750 1324 2751 1328
rect 2755 1324 2756 1328
rect 2750 1323 2756 1324
rect 2934 1328 2940 1329
rect 2934 1324 2935 1328
rect 2939 1324 2940 1328
rect 2934 1323 2940 1324
rect 3110 1328 3116 1329
rect 3110 1324 3111 1328
rect 3115 1324 3116 1328
rect 3110 1323 3116 1324
rect 3278 1328 3284 1329
rect 3278 1324 3279 1328
rect 3283 1324 3284 1328
rect 3278 1323 3284 1324
rect 3446 1328 3452 1329
rect 3446 1324 3447 1328
rect 3451 1324 3452 1328
rect 3446 1323 3452 1324
rect 3622 1328 3628 1329
rect 3622 1324 3623 1328
rect 3627 1324 3628 1328
rect 3622 1323 3628 1324
rect 3942 1325 3948 1326
rect 2046 1320 2052 1321
rect 3942 1321 3943 1325
rect 3947 1321 3948 1325
rect 3942 1320 3948 1321
rect 158 1309 164 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 158 1305 159 1309
rect 163 1305 164 1309
rect 158 1304 164 1305
rect 310 1309 316 1310
rect 310 1305 311 1309
rect 315 1305 316 1309
rect 310 1304 316 1305
rect 478 1309 484 1310
rect 478 1305 479 1309
rect 483 1305 484 1309
rect 478 1304 484 1305
rect 662 1309 668 1310
rect 662 1305 663 1309
rect 667 1305 668 1309
rect 662 1304 668 1305
rect 854 1309 860 1310
rect 854 1305 855 1309
rect 859 1305 860 1309
rect 854 1304 860 1305
rect 1046 1309 1052 1310
rect 1046 1305 1047 1309
rect 1051 1305 1052 1309
rect 1046 1304 1052 1305
rect 1246 1309 1252 1310
rect 1246 1305 1247 1309
rect 1251 1305 1252 1309
rect 1246 1304 1252 1305
rect 1446 1309 1452 1310
rect 1446 1305 1447 1309
rect 1451 1305 1452 1309
rect 1446 1304 1452 1305
rect 1654 1309 1660 1310
rect 1654 1305 1655 1309
rect 1659 1305 1660 1309
rect 1654 1304 1660 1305
rect 1862 1309 1868 1310
rect 2070 1309 2076 1310
rect 1862 1305 1863 1309
rect 1867 1305 1868 1309
rect 1862 1304 1868 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 110 1303 116 1304
rect 2006 1303 2012 1304
rect 2046 1308 2052 1309
rect 2046 1304 2047 1308
rect 2051 1304 2052 1308
rect 2070 1305 2071 1309
rect 2075 1305 2076 1309
rect 2070 1304 2076 1305
rect 2206 1309 2212 1310
rect 2206 1305 2207 1309
rect 2211 1305 2212 1309
rect 2206 1304 2212 1305
rect 2382 1309 2388 1310
rect 2382 1305 2383 1309
rect 2387 1305 2388 1309
rect 2382 1304 2388 1305
rect 2566 1309 2572 1310
rect 2566 1305 2567 1309
rect 2571 1305 2572 1309
rect 2566 1304 2572 1305
rect 2750 1309 2756 1310
rect 2750 1305 2751 1309
rect 2755 1305 2756 1309
rect 2750 1304 2756 1305
rect 2934 1309 2940 1310
rect 2934 1305 2935 1309
rect 2939 1305 2940 1309
rect 2934 1304 2940 1305
rect 3110 1309 3116 1310
rect 3110 1305 3111 1309
rect 3115 1305 3116 1309
rect 3110 1304 3116 1305
rect 3278 1309 3284 1310
rect 3278 1305 3279 1309
rect 3283 1305 3284 1309
rect 3278 1304 3284 1305
rect 3446 1309 3452 1310
rect 3446 1305 3447 1309
rect 3451 1305 3452 1309
rect 3446 1304 3452 1305
rect 3622 1309 3628 1310
rect 3622 1305 3623 1309
rect 3627 1305 3628 1309
rect 3622 1304 3628 1305
rect 3942 1308 3948 1309
rect 3942 1304 3943 1308
rect 3947 1304 3948 1308
rect 2046 1303 2052 1304
rect 3942 1303 3948 1304
rect 2046 1256 2052 1257
rect 3942 1256 3948 1257
rect 110 1252 116 1253
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 406 1251 412 1252
rect 406 1247 407 1251
rect 411 1247 412 1251
rect 406 1246 412 1247
rect 542 1251 548 1252
rect 542 1247 543 1251
rect 547 1247 548 1251
rect 542 1246 548 1247
rect 694 1251 700 1252
rect 694 1247 695 1251
rect 699 1247 700 1251
rect 694 1246 700 1247
rect 854 1251 860 1252
rect 854 1247 855 1251
rect 859 1247 860 1251
rect 854 1246 860 1247
rect 1022 1251 1028 1252
rect 1022 1247 1023 1251
rect 1027 1247 1028 1251
rect 1022 1246 1028 1247
rect 1190 1251 1196 1252
rect 1190 1247 1191 1251
rect 1195 1247 1196 1251
rect 1190 1246 1196 1247
rect 1366 1251 1372 1252
rect 1366 1247 1367 1251
rect 1371 1247 1372 1251
rect 1366 1246 1372 1247
rect 1542 1251 1548 1252
rect 1542 1247 1543 1251
rect 1547 1247 1548 1251
rect 1542 1246 1548 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 1718 1246 1724 1247
rect 1894 1251 1900 1252
rect 1894 1247 1895 1251
rect 1899 1247 1900 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2046 1252 2047 1256
rect 2051 1252 2052 1256
rect 2046 1251 2052 1252
rect 2150 1255 2156 1256
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2286 1255 2292 1256
rect 2286 1251 2287 1255
rect 2291 1251 2292 1255
rect 2286 1250 2292 1251
rect 2430 1255 2436 1256
rect 2430 1251 2431 1255
rect 2435 1251 2436 1255
rect 2430 1250 2436 1251
rect 2582 1255 2588 1256
rect 2582 1251 2583 1255
rect 2587 1251 2588 1255
rect 2582 1250 2588 1251
rect 2742 1255 2748 1256
rect 2742 1251 2743 1255
rect 2747 1251 2748 1255
rect 2742 1250 2748 1251
rect 2902 1255 2908 1256
rect 2902 1251 2903 1255
rect 2907 1251 2908 1255
rect 2902 1250 2908 1251
rect 3070 1255 3076 1256
rect 3070 1251 3071 1255
rect 3075 1251 3076 1255
rect 3070 1250 3076 1251
rect 3246 1255 3252 1256
rect 3246 1251 3247 1255
rect 3251 1251 3252 1255
rect 3246 1250 3252 1251
rect 3430 1255 3436 1256
rect 3430 1251 3431 1255
rect 3435 1251 3436 1255
rect 3430 1250 3436 1251
rect 3614 1255 3620 1256
rect 3614 1251 3615 1255
rect 3619 1251 3620 1255
rect 3614 1250 3620 1251
rect 3806 1255 3812 1256
rect 3806 1251 3807 1255
rect 3811 1251 3812 1255
rect 3942 1252 3943 1256
rect 3947 1252 3948 1256
rect 3942 1251 3948 1252
rect 3806 1250 3812 1251
rect 2006 1247 2012 1248
rect 1894 1246 1900 1247
rect 2046 1239 2052 1240
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 406 1232 412 1233
rect 406 1228 407 1232
rect 411 1228 412 1232
rect 406 1227 412 1228
rect 542 1232 548 1233
rect 542 1228 543 1232
rect 547 1228 548 1232
rect 542 1227 548 1228
rect 694 1232 700 1233
rect 694 1228 695 1232
rect 699 1228 700 1232
rect 694 1227 700 1228
rect 854 1232 860 1233
rect 854 1228 855 1232
rect 859 1228 860 1232
rect 854 1227 860 1228
rect 1022 1232 1028 1233
rect 1022 1228 1023 1232
rect 1027 1228 1028 1232
rect 1022 1227 1028 1228
rect 1190 1232 1196 1233
rect 1190 1228 1191 1232
rect 1195 1228 1196 1232
rect 1190 1227 1196 1228
rect 1366 1232 1372 1233
rect 1366 1228 1367 1232
rect 1371 1228 1372 1232
rect 1366 1227 1372 1228
rect 1542 1232 1548 1233
rect 1542 1228 1543 1232
rect 1547 1228 1548 1232
rect 1542 1227 1548 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 1718 1227 1724 1228
rect 1894 1232 1900 1233
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2046 1235 2047 1239
rect 2051 1235 2052 1239
rect 3942 1239 3948 1240
rect 2046 1234 2052 1235
rect 2150 1236 2156 1237
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2286 1236 2292 1237
rect 2286 1232 2287 1236
rect 2291 1232 2292 1236
rect 2286 1231 2292 1232
rect 2430 1236 2436 1237
rect 2430 1232 2431 1236
rect 2435 1232 2436 1236
rect 2430 1231 2436 1232
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 2582 1231 2588 1232
rect 2742 1236 2748 1237
rect 2742 1232 2743 1236
rect 2747 1232 2748 1236
rect 2742 1231 2748 1232
rect 2902 1236 2908 1237
rect 2902 1232 2903 1236
rect 2907 1232 2908 1236
rect 2902 1231 2908 1232
rect 3070 1236 3076 1237
rect 3070 1232 3071 1236
rect 3075 1232 3076 1236
rect 3070 1231 3076 1232
rect 3246 1236 3252 1237
rect 3246 1232 3247 1236
rect 3251 1232 3252 1236
rect 3246 1231 3252 1232
rect 3430 1236 3436 1237
rect 3430 1232 3431 1236
rect 3435 1232 3436 1236
rect 3430 1231 3436 1232
rect 3614 1236 3620 1237
rect 3614 1232 3615 1236
rect 3619 1232 3620 1236
rect 3614 1231 3620 1232
rect 3806 1236 3812 1237
rect 3806 1232 3807 1236
rect 3811 1232 3812 1236
rect 3942 1235 3943 1239
rect 3947 1235 3948 1239
rect 3942 1234 3948 1235
rect 3806 1231 3812 1232
rect 2006 1230 2012 1231
rect 1894 1227 1900 1228
rect 2310 1176 2316 1177
rect 2046 1173 2052 1174
rect 422 1172 428 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 422 1168 423 1172
rect 427 1168 428 1172
rect 422 1167 428 1168
rect 590 1172 596 1173
rect 590 1168 591 1172
rect 595 1168 596 1172
rect 590 1167 596 1168
rect 758 1172 764 1173
rect 758 1168 759 1172
rect 763 1168 764 1172
rect 758 1167 764 1168
rect 926 1172 932 1173
rect 926 1168 927 1172
rect 931 1168 932 1172
rect 926 1167 932 1168
rect 1094 1172 1100 1173
rect 1094 1168 1095 1172
rect 1099 1168 1100 1172
rect 1094 1167 1100 1168
rect 1246 1172 1252 1173
rect 1246 1168 1247 1172
rect 1251 1168 1252 1172
rect 1246 1167 1252 1168
rect 1398 1172 1404 1173
rect 1398 1168 1399 1172
rect 1403 1168 1404 1172
rect 1398 1167 1404 1168
rect 1542 1172 1548 1173
rect 1542 1168 1543 1172
rect 1547 1168 1548 1172
rect 1542 1167 1548 1168
rect 1686 1172 1692 1173
rect 1686 1168 1687 1172
rect 1691 1168 1692 1172
rect 1686 1167 1692 1168
rect 1838 1172 1844 1173
rect 1838 1168 1839 1172
rect 1843 1168 1844 1172
rect 1838 1167 1844 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2046 1169 2047 1173
rect 2051 1169 2052 1173
rect 2310 1172 2311 1176
rect 2315 1172 2316 1176
rect 2310 1171 2316 1172
rect 2414 1176 2420 1177
rect 2414 1172 2415 1176
rect 2419 1172 2420 1176
rect 2414 1171 2420 1172
rect 2526 1176 2532 1177
rect 2526 1172 2527 1176
rect 2531 1172 2532 1176
rect 2526 1171 2532 1172
rect 2638 1176 2644 1177
rect 2638 1172 2639 1176
rect 2643 1172 2644 1176
rect 2638 1171 2644 1172
rect 2766 1176 2772 1177
rect 2766 1172 2767 1176
rect 2771 1172 2772 1176
rect 2766 1171 2772 1172
rect 2910 1176 2916 1177
rect 2910 1172 2911 1176
rect 2915 1172 2916 1176
rect 2910 1171 2916 1172
rect 3070 1176 3076 1177
rect 3070 1172 3071 1176
rect 3075 1172 3076 1176
rect 3070 1171 3076 1172
rect 3246 1176 3252 1177
rect 3246 1172 3247 1176
rect 3251 1172 3252 1176
rect 3246 1171 3252 1172
rect 3438 1176 3444 1177
rect 3438 1172 3439 1176
rect 3443 1172 3444 1176
rect 3438 1171 3444 1172
rect 3630 1176 3636 1177
rect 3630 1172 3631 1176
rect 3635 1172 3636 1176
rect 3630 1171 3636 1172
rect 3830 1176 3836 1177
rect 3830 1172 3831 1176
rect 3835 1172 3836 1176
rect 3830 1171 3836 1172
rect 3942 1173 3948 1174
rect 2046 1168 2052 1169
rect 3942 1169 3943 1173
rect 3947 1169 3948 1173
rect 3942 1168 3948 1169
rect 2006 1164 2012 1165
rect 2310 1157 2316 1158
rect 2046 1156 2052 1157
rect 422 1153 428 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 422 1149 423 1153
rect 427 1149 428 1153
rect 422 1148 428 1149
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 758 1153 764 1154
rect 758 1149 759 1153
rect 763 1149 764 1153
rect 758 1148 764 1149
rect 926 1153 932 1154
rect 926 1149 927 1153
rect 931 1149 932 1153
rect 926 1148 932 1149
rect 1094 1153 1100 1154
rect 1094 1149 1095 1153
rect 1099 1149 1100 1153
rect 1094 1148 1100 1149
rect 1246 1153 1252 1154
rect 1246 1149 1247 1153
rect 1251 1149 1252 1153
rect 1246 1148 1252 1149
rect 1398 1153 1404 1154
rect 1398 1149 1399 1153
rect 1403 1149 1404 1153
rect 1398 1148 1404 1149
rect 1542 1153 1548 1154
rect 1542 1149 1543 1153
rect 1547 1149 1548 1153
rect 1542 1148 1548 1149
rect 1686 1153 1692 1154
rect 1686 1149 1687 1153
rect 1691 1149 1692 1153
rect 1686 1148 1692 1149
rect 1838 1153 1844 1154
rect 1838 1149 1839 1153
rect 1843 1149 1844 1153
rect 1838 1148 1844 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2046 1152 2047 1156
rect 2051 1152 2052 1156
rect 2310 1153 2311 1157
rect 2315 1153 2316 1157
rect 2310 1152 2316 1153
rect 2414 1157 2420 1158
rect 2414 1153 2415 1157
rect 2419 1153 2420 1157
rect 2414 1152 2420 1153
rect 2526 1157 2532 1158
rect 2526 1153 2527 1157
rect 2531 1153 2532 1157
rect 2526 1152 2532 1153
rect 2638 1157 2644 1158
rect 2638 1153 2639 1157
rect 2643 1153 2644 1157
rect 2638 1152 2644 1153
rect 2766 1157 2772 1158
rect 2766 1153 2767 1157
rect 2771 1153 2772 1157
rect 2766 1152 2772 1153
rect 2910 1157 2916 1158
rect 2910 1153 2911 1157
rect 2915 1153 2916 1157
rect 2910 1152 2916 1153
rect 3070 1157 3076 1158
rect 3070 1153 3071 1157
rect 3075 1153 3076 1157
rect 3070 1152 3076 1153
rect 3246 1157 3252 1158
rect 3246 1153 3247 1157
rect 3251 1153 3252 1157
rect 3246 1152 3252 1153
rect 3438 1157 3444 1158
rect 3438 1153 3439 1157
rect 3443 1153 3444 1157
rect 3438 1152 3444 1153
rect 3630 1157 3636 1158
rect 3630 1153 3631 1157
rect 3635 1153 3636 1157
rect 3630 1152 3636 1153
rect 3830 1157 3836 1158
rect 3830 1153 3831 1157
rect 3835 1153 3836 1157
rect 3830 1152 3836 1153
rect 3942 1156 3948 1157
rect 3942 1152 3943 1156
rect 3947 1152 3948 1156
rect 2046 1151 2052 1152
rect 3942 1151 3948 1152
rect 110 1147 116 1148
rect 2006 1147 2012 1148
rect 2046 1100 2052 1101
rect 3942 1100 3948 1101
rect 110 1096 116 1097
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 486 1095 492 1096
rect 486 1091 487 1095
rect 491 1091 492 1095
rect 486 1090 492 1091
rect 598 1095 604 1096
rect 598 1091 599 1095
rect 603 1091 604 1095
rect 598 1090 604 1091
rect 710 1095 716 1096
rect 710 1091 711 1095
rect 715 1091 716 1095
rect 710 1090 716 1091
rect 830 1095 836 1096
rect 830 1091 831 1095
rect 835 1091 836 1095
rect 830 1090 836 1091
rect 966 1095 972 1096
rect 966 1091 967 1095
rect 971 1091 972 1095
rect 966 1090 972 1091
rect 1118 1095 1124 1096
rect 1118 1091 1119 1095
rect 1123 1091 1124 1095
rect 1118 1090 1124 1091
rect 1278 1095 1284 1096
rect 1278 1091 1279 1095
rect 1283 1091 1284 1095
rect 1278 1090 1284 1091
rect 1446 1095 1452 1096
rect 1446 1091 1447 1095
rect 1451 1091 1452 1095
rect 1446 1090 1452 1091
rect 1622 1095 1628 1096
rect 1622 1091 1623 1095
rect 1627 1091 1628 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2046 1096 2047 1100
rect 2051 1096 2052 1100
rect 2046 1095 2052 1096
rect 2406 1099 2412 1100
rect 2406 1095 2407 1099
rect 2411 1095 2412 1099
rect 2406 1094 2412 1095
rect 2502 1099 2508 1100
rect 2502 1095 2503 1099
rect 2507 1095 2508 1099
rect 2502 1094 2508 1095
rect 2598 1099 2604 1100
rect 2598 1095 2599 1099
rect 2603 1095 2604 1099
rect 2598 1094 2604 1095
rect 2694 1099 2700 1100
rect 2694 1095 2695 1099
rect 2699 1095 2700 1099
rect 2694 1094 2700 1095
rect 2806 1099 2812 1100
rect 2806 1095 2807 1099
rect 2811 1095 2812 1099
rect 2806 1094 2812 1095
rect 2942 1099 2948 1100
rect 2942 1095 2943 1099
rect 2947 1095 2948 1099
rect 2942 1094 2948 1095
rect 3094 1099 3100 1100
rect 3094 1095 3095 1099
rect 3099 1095 3100 1099
rect 3094 1094 3100 1095
rect 3262 1099 3268 1100
rect 3262 1095 3263 1099
rect 3267 1095 3268 1099
rect 3262 1094 3268 1095
rect 3446 1099 3452 1100
rect 3446 1095 3447 1099
rect 3451 1095 3452 1099
rect 3446 1094 3452 1095
rect 3638 1099 3644 1100
rect 3638 1095 3639 1099
rect 3643 1095 3644 1099
rect 3638 1094 3644 1095
rect 3838 1099 3844 1100
rect 3838 1095 3839 1099
rect 3843 1095 3844 1099
rect 3942 1096 3943 1100
rect 3947 1096 3948 1100
rect 3942 1095 3948 1096
rect 3838 1094 3844 1095
rect 2006 1091 2012 1092
rect 1622 1090 1628 1091
rect 2046 1083 2052 1084
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 374 1076 380 1077
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 486 1076 492 1077
rect 486 1072 487 1076
rect 491 1072 492 1076
rect 486 1071 492 1072
rect 598 1076 604 1077
rect 598 1072 599 1076
rect 603 1072 604 1076
rect 598 1071 604 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 830 1076 836 1077
rect 830 1072 831 1076
rect 835 1072 836 1076
rect 830 1071 836 1072
rect 966 1076 972 1077
rect 966 1072 967 1076
rect 971 1072 972 1076
rect 966 1071 972 1072
rect 1118 1076 1124 1077
rect 1118 1072 1119 1076
rect 1123 1072 1124 1076
rect 1118 1071 1124 1072
rect 1278 1076 1284 1077
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 1446 1076 1452 1077
rect 1446 1072 1447 1076
rect 1451 1072 1452 1076
rect 1446 1071 1452 1072
rect 1622 1076 1628 1077
rect 1622 1072 1623 1076
rect 1627 1072 1628 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2046 1079 2047 1083
rect 2051 1079 2052 1083
rect 3942 1083 3948 1084
rect 2046 1078 2052 1079
rect 2406 1080 2412 1081
rect 2406 1076 2407 1080
rect 2411 1076 2412 1080
rect 2406 1075 2412 1076
rect 2502 1080 2508 1081
rect 2502 1076 2503 1080
rect 2507 1076 2508 1080
rect 2502 1075 2508 1076
rect 2598 1080 2604 1081
rect 2598 1076 2599 1080
rect 2603 1076 2604 1080
rect 2598 1075 2604 1076
rect 2694 1080 2700 1081
rect 2694 1076 2695 1080
rect 2699 1076 2700 1080
rect 2694 1075 2700 1076
rect 2806 1080 2812 1081
rect 2806 1076 2807 1080
rect 2811 1076 2812 1080
rect 2806 1075 2812 1076
rect 2942 1080 2948 1081
rect 2942 1076 2943 1080
rect 2947 1076 2948 1080
rect 2942 1075 2948 1076
rect 3094 1080 3100 1081
rect 3094 1076 3095 1080
rect 3099 1076 3100 1080
rect 3094 1075 3100 1076
rect 3262 1080 3268 1081
rect 3262 1076 3263 1080
rect 3267 1076 3268 1080
rect 3262 1075 3268 1076
rect 3446 1080 3452 1081
rect 3446 1076 3447 1080
rect 3451 1076 3452 1080
rect 3446 1075 3452 1076
rect 3638 1080 3644 1081
rect 3638 1076 3639 1080
rect 3643 1076 3644 1080
rect 3638 1075 3644 1076
rect 3838 1080 3844 1081
rect 3838 1076 3839 1080
rect 3843 1076 3844 1080
rect 3942 1079 3943 1083
rect 3947 1079 3948 1083
rect 3942 1078 3948 1079
rect 3838 1075 3844 1076
rect 2006 1074 2012 1075
rect 1622 1071 1628 1072
rect 302 1016 308 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 302 1012 303 1016
rect 307 1012 308 1016
rect 302 1011 308 1012
rect 446 1016 452 1017
rect 446 1012 447 1016
rect 451 1012 452 1016
rect 446 1011 452 1012
rect 590 1016 596 1017
rect 590 1012 591 1016
rect 595 1012 596 1016
rect 590 1011 596 1012
rect 726 1016 732 1017
rect 726 1012 727 1016
rect 731 1012 732 1016
rect 726 1011 732 1012
rect 854 1016 860 1017
rect 854 1012 855 1016
rect 859 1012 860 1016
rect 854 1011 860 1012
rect 974 1016 980 1017
rect 974 1012 975 1016
rect 979 1012 980 1016
rect 974 1011 980 1012
rect 1086 1016 1092 1017
rect 1086 1012 1087 1016
rect 1091 1012 1092 1016
rect 1086 1011 1092 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1310 1016 1316 1017
rect 1310 1012 1311 1016
rect 1315 1012 1316 1016
rect 1310 1011 1316 1012
rect 1430 1016 1436 1017
rect 1430 1012 1431 1016
rect 1435 1012 1436 1016
rect 2454 1016 2460 1017
rect 1430 1011 1436 1012
rect 2006 1013 2012 1014
rect 110 1008 116 1009
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1013 2052 1014
rect 2046 1009 2047 1013
rect 2051 1009 2052 1013
rect 2454 1012 2455 1016
rect 2459 1012 2460 1016
rect 2454 1011 2460 1012
rect 2550 1016 2556 1017
rect 2550 1012 2551 1016
rect 2555 1012 2556 1016
rect 2550 1011 2556 1012
rect 2646 1016 2652 1017
rect 2646 1012 2647 1016
rect 2651 1012 2652 1016
rect 2646 1011 2652 1012
rect 2758 1016 2764 1017
rect 2758 1012 2759 1016
rect 2763 1012 2764 1016
rect 2758 1011 2764 1012
rect 2886 1016 2892 1017
rect 2886 1012 2887 1016
rect 2891 1012 2892 1016
rect 2886 1011 2892 1012
rect 3030 1016 3036 1017
rect 3030 1012 3031 1016
rect 3035 1012 3036 1016
rect 3030 1011 3036 1012
rect 3182 1016 3188 1017
rect 3182 1012 3183 1016
rect 3187 1012 3188 1016
rect 3182 1011 3188 1012
rect 3342 1016 3348 1017
rect 3342 1012 3343 1016
rect 3347 1012 3348 1016
rect 3342 1011 3348 1012
rect 3502 1016 3508 1017
rect 3502 1012 3503 1016
rect 3507 1012 3508 1016
rect 3502 1011 3508 1012
rect 3670 1016 3676 1017
rect 3670 1012 3671 1016
rect 3675 1012 3676 1016
rect 3670 1011 3676 1012
rect 3838 1016 3844 1017
rect 3838 1012 3839 1016
rect 3843 1012 3844 1016
rect 3838 1011 3844 1012
rect 3942 1013 3948 1014
rect 2046 1008 2052 1009
rect 3942 1009 3943 1013
rect 3947 1009 3948 1013
rect 3942 1008 3948 1009
rect 302 997 308 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 302 993 303 997
rect 307 993 308 997
rect 302 992 308 993
rect 446 997 452 998
rect 446 993 447 997
rect 451 993 452 997
rect 446 992 452 993
rect 590 997 596 998
rect 590 993 591 997
rect 595 993 596 997
rect 590 992 596 993
rect 726 997 732 998
rect 726 993 727 997
rect 731 993 732 997
rect 726 992 732 993
rect 854 997 860 998
rect 854 993 855 997
rect 859 993 860 997
rect 854 992 860 993
rect 974 997 980 998
rect 974 993 975 997
rect 979 993 980 997
rect 974 992 980 993
rect 1086 997 1092 998
rect 1086 993 1087 997
rect 1091 993 1092 997
rect 1086 992 1092 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1310 997 1316 998
rect 1310 993 1311 997
rect 1315 993 1316 997
rect 1310 992 1316 993
rect 1430 997 1436 998
rect 2454 997 2460 998
rect 1430 993 1431 997
rect 1435 993 1436 997
rect 1430 992 1436 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 2006 991 2012 992
rect 2046 996 2052 997
rect 2046 992 2047 996
rect 2051 992 2052 996
rect 2454 993 2455 997
rect 2459 993 2460 997
rect 2454 992 2460 993
rect 2550 997 2556 998
rect 2550 993 2551 997
rect 2555 993 2556 997
rect 2550 992 2556 993
rect 2646 997 2652 998
rect 2646 993 2647 997
rect 2651 993 2652 997
rect 2646 992 2652 993
rect 2758 997 2764 998
rect 2758 993 2759 997
rect 2763 993 2764 997
rect 2758 992 2764 993
rect 2886 997 2892 998
rect 2886 993 2887 997
rect 2891 993 2892 997
rect 2886 992 2892 993
rect 3030 997 3036 998
rect 3030 993 3031 997
rect 3035 993 3036 997
rect 3030 992 3036 993
rect 3182 997 3188 998
rect 3182 993 3183 997
rect 3187 993 3188 997
rect 3182 992 3188 993
rect 3342 997 3348 998
rect 3342 993 3343 997
rect 3347 993 3348 997
rect 3342 992 3348 993
rect 3502 997 3508 998
rect 3502 993 3503 997
rect 3507 993 3508 997
rect 3502 992 3508 993
rect 3670 997 3676 998
rect 3670 993 3671 997
rect 3675 993 3676 997
rect 3670 992 3676 993
rect 3838 997 3844 998
rect 3838 993 3839 997
rect 3843 993 3844 997
rect 3838 992 3844 993
rect 3942 996 3948 997
rect 3942 992 3943 996
rect 3947 992 3948 996
rect 2046 991 2052 992
rect 3942 991 3948 992
rect 110 944 116 945
rect 2006 944 2012 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 254 943 260 944
rect 254 939 255 943
rect 259 939 260 943
rect 254 938 260 939
rect 446 943 452 944
rect 446 939 447 943
rect 451 939 452 943
rect 446 938 452 939
rect 630 943 636 944
rect 630 939 631 943
rect 635 939 636 943
rect 630 938 636 939
rect 806 943 812 944
rect 806 939 807 943
rect 811 939 812 943
rect 806 938 812 939
rect 974 943 980 944
rect 974 939 975 943
rect 979 939 980 943
rect 974 938 980 939
rect 1126 943 1132 944
rect 1126 939 1127 943
rect 1131 939 1132 943
rect 1126 938 1132 939
rect 1270 943 1276 944
rect 1270 939 1271 943
rect 1275 939 1276 943
rect 1270 938 1276 939
rect 1414 943 1420 944
rect 1414 939 1415 943
rect 1419 939 1420 943
rect 1414 938 1420 939
rect 1550 943 1556 944
rect 1550 939 1551 943
rect 1555 939 1556 943
rect 1550 938 1556 939
rect 1694 943 1700 944
rect 1694 939 1695 943
rect 1699 939 1700 943
rect 2006 940 2007 944
rect 2011 940 2012 944
rect 2006 939 2012 940
rect 2046 940 2052 941
rect 3942 940 3948 941
rect 1694 938 1700 939
rect 2046 936 2047 940
rect 2051 936 2052 940
rect 2046 935 2052 936
rect 2422 939 2428 940
rect 2422 935 2423 939
rect 2427 935 2428 939
rect 2422 934 2428 935
rect 2518 939 2524 940
rect 2518 935 2519 939
rect 2523 935 2524 939
rect 2518 934 2524 935
rect 2614 939 2620 940
rect 2614 935 2615 939
rect 2619 935 2620 939
rect 2614 934 2620 935
rect 2710 939 2716 940
rect 2710 935 2711 939
rect 2715 935 2716 939
rect 2710 934 2716 935
rect 2822 939 2828 940
rect 2822 935 2823 939
rect 2827 935 2828 939
rect 2822 934 2828 935
rect 2950 939 2956 940
rect 2950 935 2951 939
rect 2955 935 2956 939
rect 2950 934 2956 935
rect 3102 939 3108 940
rect 3102 935 3103 939
rect 3107 935 3108 939
rect 3102 934 3108 935
rect 3270 939 3276 940
rect 3270 935 3271 939
rect 3275 935 3276 939
rect 3270 934 3276 935
rect 3454 939 3460 940
rect 3454 935 3455 939
rect 3459 935 3460 939
rect 3454 934 3460 935
rect 3646 939 3652 940
rect 3646 935 3647 939
rect 3651 935 3652 939
rect 3646 934 3652 935
rect 3838 939 3844 940
rect 3838 935 3839 939
rect 3843 935 3844 939
rect 3942 936 3943 940
rect 3947 936 3948 940
rect 3942 935 3948 936
rect 3838 934 3844 935
rect 110 927 116 928
rect 110 923 111 927
rect 115 923 116 927
rect 2006 927 2012 928
rect 110 922 116 923
rect 254 924 260 925
rect 254 920 255 924
rect 259 920 260 924
rect 254 919 260 920
rect 446 924 452 925
rect 446 920 447 924
rect 451 920 452 924
rect 446 919 452 920
rect 630 924 636 925
rect 630 920 631 924
rect 635 920 636 924
rect 630 919 636 920
rect 806 924 812 925
rect 806 920 807 924
rect 811 920 812 924
rect 806 919 812 920
rect 974 924 980 925
rect 974 920 975 924
rect 979 920 980 924
rect 974 919 980 920
rect 1126 924 1132 925
rect 1126 920 1127 924
rect 1131 920 1132 924
rect 1126 919 1132 920
rect 1270 924 1276 925
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1414 924 1420 925
rect 1414 920 1415 924
rect 1419 920 1420 924
rect 1414 919 1420 920
rect 1550 924 1556 925
rect 1550 920 1551 924
rect 1555 920 1556 924
rect 1550 919 1556 920
rect 1694 924 1700 925
rect 1694 920 1695 924
rect 1699 920 1700 924
rect 2006 923 2007 927
rect 2011 923 2012 927
rect 2006 922 2012 923
rect 2046 923 2052 924
rect 1694 919 1700 920
rect 2046 919 2047 923
rect 2051 919 2052 923
rect 3942 923 3948 924
rect 2046 918 2052 919
rect 2422 920 2428 921
rect 2422 916 2423 920
rect 2427 916 2428 920
rect 2422 915 2428 916
rect 2518 920 2524 921
rect 2518 916 2519 920
rect 2523 916 2524 920
rect 2518 915 2524 916
rect 2614 920 2620 921
rect 2614 916 2615 920
rect 2619 916 2620 920
rect 2614 915 2620 916
rect 2710 920 2716 921
rect 2710 916 2711 920
rect 2715 916 2716 920
rect 2710 915 2716 916
rect 2822 920 2828 921
rect 2822 916 2823 920
rect 2827 916 2828 920
rect 2822 915 2828 916
rect 2950 920 2956 921
rect 2950 916 2951 920
rect 2955 916 2956 920
rect 2950 915 2956 916
rect 3102 920 3108 921
rect 3102 916 3103 920
rect 3107 916 3108 920
rect 3102 915 3108 916
rect 3270 920 3276 921
rect 3270 916 3271 920
rect 3275 916 3276 920
rect 3270 915 3276 916
rect 3454 920 3460 921
rect 3454 916 3455 920
rect 3459 916 3460 920
rect 3454 915 3460 916
rect 3646 920 3652 921
rect 3646 916 3647 920
rect 3651 916 3652 920
rect 3646 915 3652 916
rect 3838 920 3844 921
rect 3838 916 3839 920
rect 3843 916 3844 920
rect 3942 919 3943 923
rect 3947 919 3948 923
rect 3942 918 3948 919
rect 3838 915 3844 916
rect 254 860 260 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 254 856 255 860
rect 259 856 260 860
rect 254 855 260 856
rect 446 860 452 861
rect 446 856 447 860
rect 451 856 452 860
rect 446 855 452 856
rect 638 860 644 861
rect 638 856 639 860
rect 643 856 644 860
rect 638 855 644 856
rect 822 860 828 861
rect 822 856 823 860
rect 827 856 828 860
rect 822 855 828 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1166 860 1172 861
rect 1166 856 1167 860
rect 1171 856 1172 860
rect 1166 855 1172 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1478 860 1484 861
rect 1478 856 1479 860
rect 1483 856 1484 860
rect 1478 855 1484 856
rect 1630 860 1636 861
rect 1630 856 1631 860
rect 1635 856 1636 860
rect 1630 855 1636 856
rect 1782 860 1788 861
rect 1782 856 1783 860
rect 1787 856 1788 860
rect 2342 860 2348 861
rect 1782 855 1788 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2006 852 2012 853
rect 2046 857 2052 858
rect 2046 853 2047 857
rect 2051 853 2052 857
rect 2342 856 2343 860
rect 2347 856 2348 860
rect 2342 855 2348 856
rect 2438 860 2444 861
rect 2438 856 2439 860
rect 2443 856 2444 860
rect 2438 855 2444 856
rect 2534 860 2540 861
rect 2534 856 2535 860
rect 2539 856 2540 860
rect 2534 855 2540 856
rect 2630 860 2636 861
rect 2630 856 2631 860
rect 2635 856 2636 860
rect 2630 855 2636 856
rect 2734 860 2740 861
rect 2734 856 2735 860
rect 2739 856 2740 860
rect 2734 855 2740 856
rect 2862 860 2868 861
rect 2862 856 2863 860
rect 2867 856 2868 860
rect 2862 855 2868 856
rect 3014 860 3020 861
rect 3014 856 3015 860
rect 3019 856 3020 860
rect 3014 855 3020 856
rect 3190 860 3196 861
rect 3190 856 3191 860
rect 3195 856 3196 860
rect 3190 855 3196 856
rect 3390 860 3396 861
rect 3390 856 3391 860
rect 3395 856 3396 860
rect 3390 855 3396 856
rect 3606 860 3612 861
rect 3606 856 3607 860
rect 3611 856 3612 860
rect 3606 855 3612 856
rect 3822 860 3828 861
rect 3822 856 3823 860
rect 3827 856 3828 860
rect 3822 855 3828 856
rect 3942 857 3948 858
rect 2046 852 2052 853
rect 3942 853 3943 857
rect 3947 853 3948 857
rect 3942 852 3948 853
rect 254 841 260 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 254 837 255 841
rect 259 837 260 841
rect 254 836 260 837
rect 446 841 452 842
rect 446 837 447 841
rect 451 837 452 841
rect 446 836 452 837
rect 638 841 644 842
rect 638 837 639 841
rect 643 837 644 841
rect 638 836 644 837
rect 822 841 828 842
rect 822 837 823 841
rect 827 837 828 841
rect 822 836 828 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1166 841 1172 842
rect 1166 837 1167 841
rect 1171 837 1172 841
rect 1166 836 1172 837
rect 1326 841 1332 842
rect 1326 837 1327 841
rect 1331 837 1332 841
rect 1326 836 1332 837
rect 1478 841 1484 842
rect 1478 837 1479 841
rect 1483 837 1484 841
rect 1478 836 1484 837
rect 1630 841 1636 842
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1782 841 1788 842
rect 2342 841 2348 842
rect 1782 837 1783 841
rect 1787 837 1788 841
rect 1782 836 1788 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 110 835 116 836
rect 2006 835 2012 836
rect 2046 840 2052 841
rect 2046 836 2047 840
rect 2051 836 2052 840
rect 2342 837 2343 841
rect 2347 837 2348 841
rect 2342 836 2348 837
rect 2438 841 2444 842
rect 2438 837 2439 841
rect 2443 837 2444 841
rect 2438 836 2444 837
rect 2534 841 2540 842
rect 2534 837 2535 841
rect 2539 837 2540 841
rect 2534 836 2540 837
rect 2630 841 2636 842
rect 2630 837 2631 841
rect 2635 837 2636 841
rect 2630 836 2636 837
rect 2734 841 2740 842
rect 2734 837 2735 841
rect 2739 837 2740 841
rect 2734 836 2740 837
rect 2862 841 2868 842
rect 2862 837 2863 841
rect 2867 837 2868 841
rect 2862 836 2868 837
rect 3014 841 3020 842
rect 3014 837 3015 841
rect 3019 837 3020 841
rect 3014 836 3020 837
rect 3190 841 3196 842
rect 3190 837 3191 841
rect 3195 837 3196 841
rect 3190 836 3196 837
rect 3390 841 3396 842
rect 3390 837 3391 841
rect 3395 837 3396 841
rect 3390 836 3396 837
rect 3606 841 3612 842
rect 3606 837 3607 841
rect 3611 837 3612 841
rect 3606 836 3612 837
rect 3822 841 3828 842
rect 3822 837 3823 841
rect 3827 837 3828 841
rect 3822 836 3828 837
rect 3942 840 3948 841
rect 3942 836 3943 840
rect 3947 836 3948 840
rect 2046 835 2052 836
rect 3942 835 3948 836
rect 2046 788 2052 789
rect 3942 788 3948 789
rect 110 784 116 785
rect 2006 784 2012 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 158 783 164 784
rect 158 779 159 783
rect 163 779 164 783
rect 158 778 164 779
rect 310 783 316 784
rect 310 779 311 783
rect 315 779 316 783
rect 310 778 316 779
rect 470 783 476 784
rect 470 779 471 783
rect 475 779 476 783
rect 470 778 476 779
rect 622 783 628 784
rect 622 779 623 783
rect 627 779 628 783
rect 622 778 628 779
rect 774 783 780 784
rect 774 779 775 783
rect 779 779 780 783
rect 774 778 780 779
rect 934 783 940 784
rect 934 779 935 783
rect 939 779 940 783
rect 934 778 940 779
rect 1094 783 1100 784
rect 1094 779 1095 783
rect 1099 779 1100 783
rect 1094 778 1100 779
rect 1254 783 1260 784
rect 1254 779 1255 783
rect 1259 779 1260 783
rect 1254 778 1260 779
rect 1414 783 1420 784
rect 1414 779 1415 783
rect 1419 779 1420 783
rect 1414 778 1420 779
rect 1582 783 1588 784
rect 1582 779 1583 783
rect 1587 779 1588 783
rect 1582 778 1588 779
rect 1750 783 1756 784
rect 1750 779 1751 783
rect 1755 779 1756 783
rect 1750 778 1756 779
rect 1902 783 1908 784
rect 1902 779 1903 783
rect 1907 779 1908 783
rect 2006 780 2007 784
rect 2011 780 2012 784
rect 2046 784 2047 788
rect 2051 784 2052 788
rect 2046 783 2052 784
rect 2310 787 2316 788
rect 2310 783 2311 787
rect 2315 783 2316 787
rect 2310 782 2316 783
rect 2494 787 2500 788
rect 2494 783 2495 787
rect 2499 783 2500 787
rect 2494 782 2500 783
rect 2686 787 2692 788
rect 2686 783 2687 787
rect 2691 783 2692 787
rect 2686 782 2692 783
rect 2878 787 2884 788
rect 2878 783 2879 787
rect 2883 783 2884 787
rect 2878 782 2884 783
rect 3078 787 3084 788
rect 3078 783 3079 787
rect 3083 783 3084 787
rect 3078 782 3084 783
rect 3286 787 3292 788
rect 3286 783 3287 787
rect 3291 783 3292 787
rect 3286 782 3292 783
rect 3502 787 3508 788
rect 3502 783 3503 787
rect 3507 783 3508 787
rect 3502 782 3508 783
rect 3718 787 3724 788
rect 3718 783 3719 787
rect 3723 783 3724 787
rect 3942 784 3943 788
rect 3947 784 3948 788
rect 3942 783 3948 784
rect 3718 782 3724 783
rect 2006 779 2012 780
rect 1902 778 1908 779
rect 2046 771 2052 772
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 2006 767 2012 768
rect 110 762 116 763
rect 158 764 164 765
rect 158 760 159 764
rect 163 760 164 764
rect 158 759 164 760
rect 310 764 316 765
rect 310 760 311 764
rect 315 760 316 764
rect 310 759 316 760
rect 470 764 476 765
rect 470 760 471 764
rect 475 760 476 764
rect 470 759 476 760
rect 622 764 628 765
rect 622 760 623 764
rect 627 760 628 764
rect 622 759 628 760
rect 774 764 780 765
rect 774 760 775 764
rect 779 760 780 764
rect 774 759 780 760
rect 934 764 940 765
rect 934 760 935 764
rect 939 760 940 764
rect 934 759 940 760
rect 1094 764 1100 765
rect 1094 760 1095 764
rect 1099 760 1100 764
rect 1094 759 1100 760
rect 1254 764 1260 765
rect 1254 760 1255 764
rect 1259 760 1260 764
rect 1254 759 1260 760
rect 1414 764 1420 765
rect 1414 760 1415 764
rect 1419 760 1420 764
rect 1414 759 1420 760
rect 1582 764 1588 765
rect 1582 760 1583 764
rect 1587 760 1588 764
rect 1582 759 1588 760
rect 1750 764 1756 765
rect 1750 760 1751 764
rect 1755 760 1756 764
rect 1750 759 1756 760
rect 1902 764 1908 765
rect 1902 760 1903 764
rect 1907 760 1908 764
rect 2006 763 2007 767
rect 2011 763 2012 767
rect 2046 767 2047 771
rect 2051 767 2052 771
rect 3942 771 3948 772
rect 2046 766 2052 767
rect 2310 768 2316 769
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2494 768 2500 769
rect 2494 764 2495 768
rect 2499 764 2500 768
rect 2494 763 2500 764
rect 2686 768 2692 769
rect 2686 764 2687 768
rect 2691 764 2692 768
rect 2686 763 2692 764
rect 2878 768 2884 769
rect 2878 764 2879 768
rect 2883 764 2884 768
rect 2878 763 2884 764
rect 3078 768 3084 769
rect 3078 764 3079 768
rect 3083 764 3084 768
rect 3078 763 3084 764
rect 3286 768 3292 769
rect 3286 764 3287 768
rect 3291 764 3292 768
rect 3286 763 3292 764
rect 3502 768 3508 769
rect 3502 764 3503 768
rect 3507 764 3508 768
rect 3502 763 3508 764
rect 3718 768 3724 769
rect 3718 764 3719 768
rect 3723 764 3724 768
rect 3942 767 3943 771
rect 3947 767 3948 771
rect 3942 766 3948 767
rect 3718 763 3724 764
rect 2006 762 2012 763
rect 1902 759 1908 760
rect 134 704 140 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 134 700 135 704
rect 139 700 140 704
rect 134 699 140 700
rect 262 704 268 705
rect 262 700 263 704
rect 267 700 268 704
rect 262 699 268 700
rect 430 704 436 705
rect 430 700 431 704
rect 435 700 436 704
rect 430 699 436 700
rect 622 704 628 705
rect 622 700 623 704
rect 627 700 628 704
rect 622 699 628 700
rect 822 704 828 705
rect 822 700 823 704
rect 827 700 828 704
rect 822 699 828 700
rect 1014 704 1020 705
rect 1014 700 1015 704
rect 1019 700 1020 704
rect 1014 699 1020 700
rect 1206 704 1212 705
rect 1206 700 1207 704
rect 1211 700 1212 704
rect 1206 699 1212 700
rect 1390 704 1396 705
rect 1390 700 1391 704
rect 1395 700 1396 704
rect 1390 699 1396 700
rect 1566 704 1572 705
rect 1566 700 1567 704
rect 1571 700 1572 704
rect 1566 699 1572 700
rect 1742 704 1748 705
rect 1742 700 1743 704
rect 1747 700 1748 704
rect 1742 699 1748 700
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2070 704 2076 705
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2046 701 2052 702
rect 2046 697 2047 701
rect 2051 697 2052 701
rect 2070 700 2071 704
rect 2075 700 2076 704
rect 2070 699 2076 700
rect 2254 704 2260 705
rect 2254 700 2255 704
rect 2259 700 2260 704
rect 2254 699 2260 700
rect 2454 704 2460 705
rect 2454 700 2455 704
rect 2459 700 2460 704
rect 2454 699 2460 700
rect 2654 704 2660 705
rect 2654 700 2655 704
rect 2659 700 2660 704
rect 2654 699 2660 700
rect 2854 704 2860 705
rect 2854 700 2855 704
rect 2859 700 2860 704
rect 2854 699 2860 700
rect 3046 704 3052 705
rect 3046 700 3047 704
rect 3051 700 3052 704
rect 3046 699 3052 700
rect 3238 704 3244 705
rect 3238 700 3239 704
rect 3243 700 3244 704
rect 3238 699 3244 700
rect 3438 704 3444 705
rect 3438 700 3439 704
rect 3443 700 3444 704
rect 3438 699 3444 700
rect 3638 704 3644 705
rect 3638 700 3639 704
rect 3643 700 3644 704
rect 3638 699 3644 700
rect 3838 704 3844 705
rect 3838 700 3839 704
rect 3843 700 3844 704
rect 3838 699 3844 700
rect 3942 701 3948 702
rect 2046 696 2052 697
rect 3942 697 3943 701
rect 3947 697 3948 701
rect 3942 696 3948 697
rect 134 685 140 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 134 681 135 685
rect 139 681 140 685
rect 134 680 140 681
rect 262 685 268 686
rect 262 681 263 685
rect 267 681 268 685
rect 262 680 268 681
rect 430 685 436 686
rect 430 681 431 685
rect 435 681 436 685
rect 430 680 436 681
rect 622 685 628 686
rect 622 681 623 685
rect 627 681 628 685
rect 622 680 628 681
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 1014 685 1020 686
rect 1014 681 1015 685
rect 1019 681 1020 685
rect 1014 680 1020 681
rect 1206 685 1212 686
rect 1206 681 1207 685
rect 1211 681 1212 685
rect 1206 680 1212 681
rect 1390 685 1396 686
rect 1390 681 1391 685
rect 1395 681 1396 685
rect 1390 680 1396 681
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 1742 685 1748 686
rect 1742 681 1743 685
rect 1747 681 1748 685
rect 1742 680 1748 681
rect 1902 685 1908 686
rect 2070 685 2076 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 2006 679 2012 680
rect 2046 684 2052 685
rect 2046 680 2047 684
rect 2051 680 2052 684
rect 2070 681 2071 685
rect 2075 681 2076 685
rect 2070 680 2076 681
rect 2254 685 2260 686
rect 2254 681 2255 685
rect 2259 681 2260 685
rect 2254 680 2260 681
rect 2454 685 2460 686
rect 2454 681 2455 685
rect 2459 681 2460 685
rect 2454 680 2460 681
rect 2654 685 2660 686
rect 2654 681 2655 685
rect 2659 681 2660 685
rect 2654 680 2660 681
rect 2854 685 2860 686
rect 2854 681 2855 685
rect 2859 681 2860 685
rect 2854 680 2860 681
rect 3046 685 3052 686
rect 3046 681 3047 685
rect 3051 681 3052 685
rect 3046 680 3052 681
rect 3238 685 3244 686
rect 3238 681 3239 685
rect 3243 681 3244 685
rect 3238 680 3244 681
rect 3438 685 3444 686
rect 3438 681 3439 685
rect 3443 681 3444 685
rect 3438 680 3444 681
rect 3638 685 3644 686
rect 3638 681 3639 685
rect 3643 681 3644 685
rect 3638 680 3644 681
rect 3838 685 3844 686
rect 3838 681 3839 685
rect 3843 681 3844 685
rect 3838 680 3844 681
rect 3942 684 3948 685
rect 3942 680 3943 684
rect 3947 680 3948 684
rect 2046 679 2052 680
rect 3942 679 3948 680
rect 110 632 116 633
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 134 631 140 632
rect 134 627 135 631
rect 139 627 140 631
rect 134 626 140 627
rect 246 631 252 632
rect 246 627 247 631
rect 251 627 252 631
rect 246 626 252 627
rect 382 631 388 632
rect 382 627 383 631
rect 387 627 388 631
rect 382 626 388 627
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 870 631 876 632
rect 870 627 871 631
rect 875 627 876 631
rect 870 626 876 627
rect 1078 631 1084 632
rect 1078 627 1079 631
rect 1083 627 1084 631
rect 1078 626 1084 627
rect 1302 631 1308 632
rect 1302 627 1303 631
rect 1307 627 1308 631
rect 1302 626 1308 627
rect 1542 631 1548 632
rect 1542 627 1543 631
rect 1547 627 1548 631
rect 1542 626 1548 627
rect 1782 631 1788 632
rect 1782 627 1783 631
rect 1787 627 1788 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 632 2052 633
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2070 631 2076 632
rect 2070 627 2071 631
rect 2075 627 2076 631
rect 1782 626 1788 627
rect 2070 626 2076 627
rect 2230 631 2236 632
rect 2230 627 2231 631
rect 2235 627 2236 631
rect 2230 626 2236 627
rect 2430 631 2436 632
rect 2430 627 2431 631
rect 2435 627 2436 631
rect 2430 626 2436 627
rect 2630 631 2636 632
rect 2630 627 2631 631
rect 2635 627 2636 631
rect 2630 626 2636 627
rect 2830 631 2836 632
rect 2830 627 2831 631
rect 2835 627 2836 631
rect 2830 626 2836 627
rect 3022 631 3028 632
rect 3022 627 3023 631
rect 3027 627 3028 631
rect 3022 626 3028 627
rect 3206 631 3212 632
rect 3206 627 3207 631
rect 3211 627 3212 631
rect 3206 626 3212 627
rect 3374 631 3380 632
rect 3374 627 3375 631
rect 3379 627 3380 631
rect 3374 626 3380 627
rect 3534 631 3540 632
rect 3534 627 3535 631
rect 3539 627 3540 631
rect 3534 626 3540 627
rect 3694 631 3700 632
rect 3694 627 3695 631
rect 3699 627 3700 631
rect 3694 626 3700 627
rect 3838 631 3844 632
rect 3838 627 3839 631
rect 3843 627 3844 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3838 626 3844 627
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 2006 615 2012 616
rect 110 610 116 611
rect 134 612 140 613
rect 134 608 135 612
rect 139 608 140 612
rect 134 607 140 608
rect 246 612 252 613
rect 246 608 247 612
rect 251 608 252 612
rect 246 607 252 608
rect 382 612 388 613
rect 382 608 383 612
rect 387 608 388 612
rect 382 607 388 608
rect 526 612 532 613
rect 526 608 527 612
rect 531 608 532 612
rect 526 607 532 608
rect 686 612 692 613
rect 686 608 687 612
rect 691 608 692 612
rect 686 607 692 608
rect 870 612 876 613
rect 870 608 871 612
rect 875 608 876 612
rect 870 607 876 608
rect 1078 612 1084 613
rect 1078 608 1079 612
rect 1083 608 1084 612
rect 1078 607 1084 608
rect 1302 612 1308 613
rect 1302 608 1303 612
rect 1307 608 1308 612
rect 1302 607 1308 608
rect 1542 612 1548 613
rect 1542 608 1543 612
rect 1547 608 1548 612
rect 1542 607 1548 608
rect 1782 612 1788 613
rect 1782 608 1783 612
rect 1787 608 1788 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 615 2052 616
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2070 612 2076 613
rect 1782 607 1788 608
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 2230 612 2236 613
rect 2230 608 2231 612
rect 2235 608 2236 612
rect 2230 607 2236 608
rect 2430 612 2436 613
rect 2430 608 2431 612
rect 2435 608 2436 612
rect 2430 607 2436 608
rect 2630 612 2636 613
rect 2630 608 2631 612
rect 2635 608 2636 612
rect 2630 607 2636 608
rect 2830 612 2836 613
rect 2830 608 2831 612
rect 2835 608 2836 612
rect 2830 607 2836 608
rect 3022 612 3028 613
rect 3022 608 3023 612
rect 3027 608 3028 612
rect 3022 607 3028 608
rect 3206 612 3212 613
rect 3206 608 3207 612
rect 3211 608 3212 612
rect 3206 607 3212 608
rect 3374 612 3380 613
rect 3374 608 3375 612
rect 3379 608 3380 612
rect 3374 607 3380 608
rect 3534 612 3540 613
rect 3534 608 3535 612
rect 3539 608 3540 612
rect 3534 607 3540 608
rect 3694 612 3700 613
rect 3694 608 3695 612
rect 3699 608 3700 612
rect 3694 607 3700 608
rect 3838 612 3844 613
rect 3838 608 3839 612
rect 3843 608 3844 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3838 607 3844 608
rect 134 548 140 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 134 544 135 548
rect 139 544 140 548
rect 134 543 140 544
rect 294 548 300 549
rect 294 544 295 548
rect 299 544 300 548
rect 294 543 300 544
rect 478 548 484 549
rect 478 544 479 548
rect 483 544 484 548
rect 478 543 484 544
rect 662 548 668 549
rect 662 544 663 548
rect 667 544 668 548
rect 662 543 668 544
rect 846 548 852 549
rect 846 544 847 548
rect 851 544 852 548
rect 846 543 852 544
rect 1030 548 1036 549
rect 1030 544 1031 548
rect 1035 544 1036 548
rect 1030 543 1036 544
rect 1214 548 1220 549
rect 1214 544 1215 548
rect 1219 544 1220 548
rect 1214 543 1220 544
rect 1398 548 1404 549
rect 1398 544 1399 548
rect 1403 544 1404 548
rect 1398 543 1404 544
rect 1590 548 1596 549
rect 1590 544 1591 548
rect 1595 544 1596 548
rect 1590 543 1596 544
rect 1782 548 1788 549
rect 1782 544 1783 548
rect 1787 544 1788 548
rect 2070 548 2076 549
rect 1782 543 1788 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2214 548 2220 549
rect 2214 544 2215 548
rect 2219 544 2220 548
rect 2214 543 2220 544
rect 2398 548 2404 549
rect 2398 544 2399 548
rect 2403 544 2404 548
rect 2398 543 2404 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2774 548 2780 549
rect 2774 544 2775 548
rect 2779 544 2780 548
rect 2774 543 2780 544
rect 2958 548 2964 549
rect 2958 544 2959 548
rect 2963 544 2964 548
rect 2958 543 2964 544
rect 3142 548 3148 549
rect 3142 544 3143 548
rect 3147 544 3148 548
rect 3142 543 3148 544
rect 3318 548 3324 549
rect 3318 544 3319 548
rect 3323 544 3324 548
rect 3318 543 3324 544
rect 3494 548 3500 549
rect 3494 544 3495 548
rect 3499 544 3500 548
rect 3494 543 3500 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3678 543 3684 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 134 529 140 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 134 525 135 529
rect 139 525 140 529
rect 134 524 140 525
rect 294 529 300 530
rect 294 525 295 529
rect 299 525 300 529
rect 294 524 300 525
rect 478 529 484 530
rect 478 525 479 529
rect 483 525 484 529
rect 478 524 484 525
rect 662 529 668 530
rect 662 525 663 529
rect 667 525 668 529
rect 662 524 668 525
rect 846 529 852 530
rect 846 525 847 529
rect 851 525 852 529
rect 846 524 852 525
rect 1030 529 1036 530
rect 1030 525 1031 529
rect 1035 525 1036 529
rect 1030 524 1036 525
rect 1214 529 1220 530
rect 1214 525 1215 529
rect 1219 525 1220 529
rect 1214 524 1220 525
rect 1398 529 1404 530
rect 1398 525 1399 529
rect 1403 525 1404 529
rect 1398 524 1404 525
rect 1590 529 1596 530
rect 1590 525 1591 529
rect 1595 525 1596 529
rect 1590 524 1596 525
rect 1782 529 1788 530
rect 2070 529 2076 530
rect 1782 525 1783 529
rect 1787 525 1788 529
rect 1782 524 1788 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2214 529 2220 530
rect 2214 525 2215 529
rect 2219 525 2220 529
rect 2214 524 2220 525
rect 2398 529 2404 530
rect 2398 525 2399 529
rect 2403 525 2404 529
rect 2398 524 2404 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2774 529 2780 530
rect 2774 525 2775 529
rect 2779 525 2780 529
rect 2774 524 2780 525
rect 2958 529 2964 530
rect 2958 525 2959 529
rect 2963 525 2964 529
rect 2958 524 2964 525
rect 3142 529 3148 530
rect 3142 525 3143 529
rect 3147 525 3148 529
rect 3142 524 3148 525
rect 3318 529 3324 530
rect 3318 525 3319 529
rect 3323 525 3324 529
rect 3318 524 3324 525
rect 3494 529 3500 530
rect 3494 525 3495 529
rect 3499 525 3500 529
rect 3494 524 3500 525
rect 3678 529 3684 530
rect 3678 525 3679 529
rect 3683 525 3684 529
rect 3678 524 3684 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 3942 523 3948 524
rect 110 476 116 477
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 454 475 460 476
rect 454 471 455 475
rect 459 471 460 475
rect 454 470 460 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 766 475 772 476
rect 766 471 767 475
rect 771 471 772 475
rect 766 470 772 471
rect 902 475 908 476
rect 902 471 903 475
rect 907 471 908 475
rect 902 470 908 471
rect 1030 475 1036 476
rect 1030 471 1031 475
rect 1035 471 1036 475
rect 1030 470 1036 471
rect 1158 475 1164 476
rect 1158 471 1159 475
rect 1163 471 1164 475
rect 1158 470 1164 471
rect 1286 475 1292 476
rect 1286 471 1287 475
rect 1291 471 1292 475
rect 1286 470 1292 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2006 471 2012 472
rect 2046 472 2052 473
rect 3942 472 3948 473
rect 1414 470 1420 471
rect 2046 468 2047 472
rect 2051 468 2052 472
rect 2046 467 2052 468
rect 2070 471 2076 472
rect 2070 467 2071 471
rect 2075 467 2076 471
rect 2070 466 2076 467
rect 2222 471 2228 472
rect 2222 467 2223 471
rect 2227 467 2228 471
rect 2222 466 2228 467
rect 2390 471 2396 472
rect 2390 467 2391 471
rect 2395 467 2396 471
rect 2390 466 2396 467
rect 2558 471 2564 472
rect 2558 467 2559 471
rect 2563 467 2564 471
rect 2558 466 2564 467
rect 2726 471 2732 472
rect 2726 467 2727 471
rect 2731 467 2732 471
rect 2726 466 2732 467
rect 2894 471 2900 472
rect 2894 467 2895 471
rect 2899 467 2900 471
rect 2894 466 2900 467
rect 3062 471 3068 472
rect 3062 467 3063 471
rect 3067 467 3068 471
rect 3062 466 3068 467
rect 3222 471 3228 472
rect 3222 467 3223 471
rect 3227 467 3228 471
rect 3222 466 3228 467
rect 3382 471 3388 472
rect 3382 467 3383 471
rect 3387 467 3388 471
rect 3382 466 3388 467
rect 3542 471 3548 472
rect 3542 467 3543 471
rect 3547 467 3548 471
rect 3542 466 3548 467
rect 3702 471 3708 472
rect 3702 467 3703 471
rect 3707 467 3708 471
rect 3702 466 3708 467
rect 3838 471 3844 472
rect 3838 467 3839 471
rect 3843 467 3844 471
rect 3942 468 3943 472
rect 3947 468 3948 472
rect 3942 467 3948 468
rect 3838 466 3844 467
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 454 456 460 457
rect 454 452 455 456
rect 459 452 460 456
rect 454 451 460 452
rect 614 456 620 457
rect 614 452 615 456
rect 619 452 620 456
rect 614 451 620 452
rect 766 456 772 457
rect 766 452 767 456
rect 771 452 772 456
rect 766 451 772 452
rect 902 456 908 457
rect 902 452 903 456
rect 907 452 908 456
rect 902 451 908 452
rect 1030 456 1036 457
rect 1030 452 1031 456
rect 1035 452 1036 456
rect 1030 451 1036 452
rect 1158 456 1164 457
rect 1158 452 1159 456
rect 1163 452 1164 456
rect 1158 451 1164 452
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1286 451 1292 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 455 2052 456
rect 1414 451 1420 452
rect 2046 451 2047 455
rect 2051 451 2052 455
rect 3942 455 3948 456
rect 2046 450 2052 451
rect 2070 452 2076 453
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 2222 452 2228 453
rect 2222 448 2223 452
rect 2227 448 2228 452
rect 2222 447 2228 448
rect 2390 452 2396 453
rect 2390 448 2391 452
rect 2395 448 2396 452
rect 2390 447 2396 448
rect 2558 452 2564 453
rect 2558 448 2559 452
rect 2563 448 2564 452
rect 2558 447 2564 448
rect 2726 452 2732 453
rect 2726 448 2727 452
rect 2731 448 2732 452
rect 2726 447 2732 448
rect 2894 452 2900 453
rect 2894 448 2895 452
rect 2899 448 2900 452
rect 2894 447 2900 448
rect 3062 452 3068 453
rect 3062 448 3063 452
rect 3067 448 3068 452
rect 3062 447 3068 448
rect 3222 452 3228 453
rect 3222 448 3223 452
rect 3227 448 3228 452
rect 3222 447 3228 448
rect 3382 452 3388 453
rect 3382 448 3383 452
rect 3387 448 3388 452
rect 3382 447 3388 448
rect 3542 452 3548 453
rect 3542 448 3543 452
rect 3547 448 3548 452
rect 3542 447 3548 448
rect 3702 452 3708 453
rect 3702 448 3703 452
rect 3707 448 3708 452
rect 3702 447 3708 448
rect 3838 452 3844 453
rect 3838 448 3839 452
rect 3843 448 3844 452
rect 3942 451 3943 455
rect 3947 451 3948 455
rect 3942 450 3948 451
rect 3838 447 3844 448
rect 134 396 140 397
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 134 392 135 396
rect 139 392 140 396
rect 134 391 140 392
rect 286 396 292 397
rect 286 392 287 396
rect 291 392 292 396
rect 286 391 292 392
rect 446 396 452 397
rect 446 392 447 396
rect 451 392 452 396
rect 446 391 452 392
rect 598 396 604 397
rect 598 392 599 396
rect 603 392 604 396
rect 598 391 604 392
rect 750 396 756 397
rect 750 392 751 396
rect 755 392 756 396
rect 750 391 756 392
rect 902 396 908 397
rect 902 392 903 396
rect 907 392 908 396
rect 902 391 908 392
rect 1078 396 1084 397
rect 1078 392 1079 396
rect 1083 392 1084 396
rect 1078 391 1084 392
rect 1270 396 1276 397
rect 1270 392 1271 396
rect 1275 392 1276 396
rect 1270 391 1276 392
rect 1478 396 1484 397
rect 1478 392 1479 396
rect 1483 392 1484 396
rect 1478 391 1484 392
rect 1702 396 1708 397
rect 1702 392 1703 396
rect 1707 392 1708 396
rect 1702 391 1708 392
rect 1902 396 1908 397
rect 1902 392 1903 396
rect 1907 392 1908 396
rect 1902 391 1908 392
rect 2006 393 2012 394
rect 110 388 116 389
rect 2006 389 2007 393
rect 2011 389 2012 393
rect 2462 392 2468 393
rect 2006 388 2012 389
rect 2046 389 2052 390
rect 2046 385 2047 389
rect 2051 385 2052 389
rect 2462 388 2463 392
rect 2467 388 2468 392
rect 2462 387 2468 388
rect 2558 392 2564 393
rect 2558 388 2559 392
rect 2563 388 2564 392
rect 2558 387 2564 388
rect 2654 392 2660 393
rect 2654 388 2655 392
rect 2659 388 2660 392
rect 2654 387 2660 388
rect 2750 392 2756 393
rect 2750 388 2751 392
rect 2755 388 2756 392
rect 2750 387 2756 388
rect 2846 392 2852 393
rect 2846 388 2847 392
rect 2851 388 2852 392
rect 2846 387 2852 388
rect 2942 392 2948 393
rect 2942 388 2943 392
rect 2947 388 2948 392
rect 2942 387 2948 388
rect 3038 392 3044 393
rect 3038 388 3039 392
rect 3043 388 3044 392
rect 3038 387 3044 388
rect 3134 392 3140 393
rect 3134 388 3135 392
rect 3139 388 3140 392
rect 3134 387 3140 388
rect 3230 392 3236 393
rect 3230 388 3231 392
rect 3235 388 3236 392
rect 3230 387 3236 388
rect 3942 389 3948 390
rect 2046 384 2052 385
rect 3942 385 3943 389
rect 3947 385 3948 389
rect 3942 384 3948 385
rect 134 377 140 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 134 373 135 377
rect 139 373 140 377
rect 134 372 140 373
rect 286 377 292 378
rect 286 373 287 377
rect 291 373 292 377
rect 286 372 292 373
rect 446 377 452 378
rect 446 373 447 377
rect 451 373 452 377
rect 446 372 452 373
rect 598 377 604 378
rect 598 373 599 377
rect 603 373 604 377
rect 598 372 604 373
rect 750 377 756 378
rect 750 373 751 377
rect 755 373 756 377
rect 750 372 756 373
rect 902 377 908 378
rect 902 373 903 377
rect 907 373 908 377
rect 902 372 908 373
rect 1078 377 1084 378
rect 1078 373 1079 377
rect 1083 373 1084 377
rect 1078 372 1084 373
rect 1270 377 1276 378
rect 1270 373 1271 377
rect 1275 373 1276 377
rect 1270 372 1276 373
rect 1478 377 1484 378
rect 1478 373 1479 377
rect 1483 373 1484 377
rect 1478 372 1484 373
rect 1702 377 1708 378
rect 1702 373 1703 377
rect 1707 373 1708 377
rect 1702 372 1708 373
rect 1902 377 1908 378
rect 1902 373 1903 377
rect 1907 373 1908 377
rect 1902 372 1908 373
rect 2006 376 2012 377
rect 2006 372 2007 376
rect 2011 372 2012 376
rect 2462 373 2468 374
rect 110 371 116 372
rect 2006 371 2012 372
rect 2046 372 2052 373
rect 2046 368 2047 372
rect 2051 368 2052 372
rect 2462 369 2463 373
rect 2467 369 2468 373
rect 2462 368 2468 369
rect 2558 373 2564 374
rect 2558 369 2559 373
rect 2563 369 2564 373
rect 2558 368 2564 369
rect 2654 373 2660 374
rect 2654 369 2655 373
rect 2659 369 2660 373
rect 2654 368 2660 369
rect 2750 373 2756 374
rect 2750 369 2751 373
rect 2755 369 2756 373
rect 2750 368 2756 369
rect 2846 373 2852 374
rect 2846 369 2847 373
rect 2851 369 2852 373
rect 2846 368 2852 369
rect 2942 373 2948 374
rect 2942 369 2943 373
rect 2947 369 2948 373
rect 2942 368 2948 369
rect 3038 373 3044 374
rect 3038 369 3039 373
rect 3043 369 3044 373
rect 3038 368 3044 369
rect 3134 373 3140 374
rect 3134 369 3135 373
rect 3139 369 3140 373
rect 3134 368 3140 369
rect 3230 373 3236 374
rect 3230 369 3231 373
rect 3235 369 3236 373
rect 3230 368 3236 369
rect 3942 372 3948 373
rect 3942 368 3943 372
rect 3947 368 3948 372
rect 2046 367 2052 368
rect 3942 367 3948 368
rect 110 320 116 321
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 158 319 164 320
rect 158 315 159 319
rect 163 315 164 319
rect 158 314 164 315
rect 350 319 356 320
rect 350 315 351 319
rect 355 315 356 319
rect 350 314 356 315
rect 550 319 556 320
rect 550 315 551 319
rect 555 315 556 319
rect 550 314 556 315
rect 758 319 764 320
rect 758 315 759 319
rect 763 315 764 319
rect 758 314 764 315
rect 958 319 964 320
rect 958 315 959 319
rect 963 315 964 319
rect 958 314 964 315
rect 1158 319 1164 320
rect 1158 315 1159 319
rect 1163 315 1164 319
rect 1158 314 1164 315
rect 1342 319 1348 320
rect 1342 315 1343 319
rect 1347 315 1348 319
rect 1342 314 1348 315
rect 1526 319 1532 320
rect 1526 315 1527 319
rect 1531 315 1532 319
rect 1526 314 1532 315
rect 1710 319 1716 320
rect 1710 315 1711 319
rect 1715 315 1716 319
rect 1710 314 1716 315
rect 1894 319 1900 320
rect 1894 315 1895 319
rect 1899 315 1900 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2398 319 2404 320
rect 2398 315 2399 319
rect 2403 315 2404 319
rect 1894 314 1900 315
rect 2398 314 2404 315
rect 2502 319 2508 320
rect 2502 315 2503 319
rect 2507 315 2508 319
rect 2502 314 2508 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2758 319 2764 320
rect 2758 315 2759 319
rect 2763 315 2764 319
rect 2758 314 2764 315
rect 2910 319 2916 320
rect 2910 315 2911 319
rect 2915 315 2916 319
rect 2910 314 2916 315
rect 3070 319 3076 320
rect 3070 315 3071 319
rect 3075 315 3076 319
rect 3070 314 3076 315
rect 3246 319 3252 320
rect 3246 315 3247 319
rect 3251 315 3252 319
rect 3246 314 3252 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3606 319 3612 320
rect 3606 315 3607 319
rect 3611 315 3612 319
rect 3606 314 3612 315
rect 3790 319 3796 320
rect 3790 315 3791 319
rect 3795 315 3796 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3790 314 3796 315
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 158 300 164 301
rect 158 296 159 300
rect 163 296 164 300
rect 158 295 164 296
rect 350 300 356 301
rect 350 296 351 300
rect 355 296 356 300
rect 350 295 356 296
rect 550 300 556 301
rect 550 296 551 300
rect 555 296 556 300
rect 550 295 556 296
rect 758 300 764 301
rect 758 296 759 300
rect 763 296 764 300
rect 758 295 764 296
rect 958 300 964 301
rect 958 296 959 300
rect 963 296 964 300
rect 958 295 964 296
rect 1158 300 1164 301
rect 1158 296 1159 300
rect 1163 296 1164 300
rect 1158 295 1164 296
rect 1342 300 1348 301
rect 1342 296 1343 300
rect 1347 296 1348 300
rect 1342 295 1348 296
rect 1526 300 1532 301
rect 1526 296 1527 300
rect 1531 296 1532 300
rect 1526 295 1532 296
rect 1710 300 1716 301
rect 1710 296 1711 300
rect 1715 296 1716 300
rect 1710 295 1716 296
rect 1894 300 1900 301
rect 1894 296 1895 300
rect 1899 296 1900 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2398 300 2404 301
rect 1894 295 1900 296
rect 2398 296 2399 300
rect 2403 296 2404 300
rect 2398 295 2404 296
rect 2502 300 2508 301
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2758 300 2764 301
rect 2758 296 2759 300
rect 2763 296 2764 300
rect 2758 295 2764 296
rect 2910 300 2916 301
rect 2910 296 2911 300
rect 2915 296 2916 300
rect 2910 295 2916 296
rect 3070 300 3076 301
rect 3070 296 3071 300
rect 3075 296 3076 300
rect 3070 295 3076 296
rect 3246 300 3252 301
rect 3246 296 3247 300
rect 3251 296 3252 300
rect 3246 295 3252 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3606 300 3612 301
rect 3606 296 3607 300
rect 3611 296 3612 300
rect 3606 295 3612 296
rect 3790 300 3796 301
rect 3790 296 3791 300
rect 3795 296 3796 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3790 295 3796 296
rect 2190 240 2196 241
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2190 236 2191 240
rect 2195 236 2196 240
rect 2190 235 2196 236
rect 2350 240 2356 241
rect 2350 236 2351 240
rect 2355 236 2356 240
rect 2350 235 2356 236
rect 2518 240 2524 241
rect 2518 236 2519 240
rect 2523 236 2524 240
rect 2518 235 2524 236
rect 2686 240 2692 241
rect 2686 236 2687 240
rect 2691 236 2692 240
rect 2686 235 2692 236
rect 2854 240 2860 241
rect 2854 236 2855 240
rect 2859 236 2860 240
rect 2854 235 2860 236
rect 3030 240 3036 241
rect 3030 236 3031 240
rect 3035 236 3036 240
rect 3030 235 3036 236
rect 3214 240 3220 241
rect 3214 236 3215 240
rect 3219 236 3220 240
rect 3214 235 3220 236
rect 3406 240 3412 241
rect 3406 236 3407 240
rect 3411 236 3412 240
rect 3406 235 3412 236
rect 3606 240 3612 241
rect 3606 236 3607 240
rect 3611 236 3612 240
rect 3606 235 3612 236
rect 3806 240 3812 241
rect 3806 236 3807 240
rect 3811 236 3812 240
rect 3806 235 3812 236
rect 3942 237 3948 238
rect 222 232 228 233
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 222 228 223 232
rect 227 228 228 232
rect 222 227 228 228
rect 382 232 388 233
rect 382 228 383 232
rect 387 228 388 232
rect 382 227 388 228
rect 542 232 548 233
rect 542 228 543 232
rect 547 228 548 232
rect 542 227 548 228
rect 702 232 708 233
rect 702 228 703 232
rect 707 228 708 232
rect 702 227 708 228
rect 862 232 868 233
rect 862 228 863 232
rect 867 228 868 232
rect 862 227 868 228
rect 1030 232 1036 233
rect 1030 228 1031 232
rect 1035 228 1036 232
rect 1030 227 1036 228
rect 1198 232 1204 233
rect 1198 228 1199 232
rect 1203 228 1204 232
rect 1198 227 1204 228
rect 1366 232 1372 233
rect 1366 228 1367 232
rect 1371 228 1372 232
rect 1366 227 1372 228
rect 1542 232 1548 233
rect 1542 228 1543 232
rect 1547 228 1548 232
rect 1542 227 1548 228
rect 1726 232 1732 233
rect 1726 228 1727 232
rect 1731 228 1732 232
rect 1726 227 1732 228
rect 1902 232 1908 233
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 1902 228 1903 232
rect 1907 228 1908 232
rect 1902 227 1908 228
rect 2006 229 2012 230
rect 110 224 116 225
rect 2006 225 2007 229
rect 2011 225 2012 229
rect 2006 224 2012 225
rect 2190 221 2196 222
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2190 217 2191 221
rect 2195 217 2196 221
rect 2190 216 2196 217
rect 2350 221 2356 222
rect 2350 217 2351 221
rect 2355 217 2356 221
rect 2350 216 2356 217
rect 2518 221 2524 222
rect 2518 217 2519 221
rect 2523 217 2524 221
rect 2518 216 2524 217
rect 2686 221 2692 222
rect 2686 217 2687 221
rect 2691 217 2692 221
rect 2686 216 2692 217
rect 2854 221 2860 222
rect 2854 217 2855 221
rect 2859 217 2860 221
rect 2854 216 2860 217
rect 3030 221 3036 222
rect 3030 217 3031 221
rect 3035 217 3036 221
rect 3030 216 3036 217
rect 3214 221 3220 222
rect 3214 217 3215 221
rect 3219 217 3220 221
rect 3214 216 3220 217
rect 3406 221 3412 222
rect 3406 217 3407 221
rect 3411 217 3412 221
rect 3406 216 3412 217
rect 3606 221 3612 222
rect 3606 217 3607 221
rect 3611 217 3612 221
rect 3606 216 3612 217
rect 3806 221 3812 222
rect 3806 217 3807 221
rect 3811 217 3812 221
rect 3806 216 3812 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 3942 215 3948 216
rect 222 213 228 214
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 222 209 223 213
rect 227 209 228 213
rect 222 208 228 209
rect 382 213 388 214
rect 382 209 383 213
rect 387 209 388 213
rect 382 208 388 209
rect 542 213 548 214
rect 542 209 543 213
rect 547 209 548 213
rect 542 208 548 209
rect 702 213 708 214
rect 702 209 703 213
rect 707 209 708 213
rect 702 208 708 209
rect 862 213 868 214
rect 862 209 863 213
rect 867 209 868 213
rect 862 208 868 209
rect 1030 213 1036 214
rect 1030 209 1031 213
rect 1035 209 1036 213
rect 1030 208 1036 209
rect 1198 213 1204 214
rect 1198 209 1199 213
rect 1203 209 1204 213
rect 1198 208 1204 209
rect 1366 213 1372 214
rect 1366 209 1367 213
rect 1371 209 1372 213
rect 1366 208 1372 209
rect 1542 213 1548 214
rect 1542 209 1543 213
rect 1547 209 1548 213
rect 1542 208 1548 209
rect 1726 213 1732 214
rect 1726 209 1727 213
rect 1731 209 1732 213
rect 1726 208 1732 209
rect 1902 213 1908 214
rect 1902 209 1903 213
rect 1907 209 1908 213
rect 1902 208 1908 209
rect 2006 212 2012 213
rect 2006 208 2007 212
rect 2011 208 2012 212
rect 110 207 116 208
rect 2006 207 2012 208
rect 110 140 116 141
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2006 135 2012 136
rect 2046 136 2052 137
rect 3942 136 3948 137
rect 1902 134 1908 135
rect 2046 132 2047 136
rect 2051 132 2052 136
rect 2046 131 2052 132
rect 2070 135 2076 136
rect 2070 131 2071 135
rect 2075 131 2076 135
rect 2070 130 2076 131
rect 2166 135 2172 136
rect 2166 131 2167 135
rect 2171 131 2172 135
rect 2166 130 2172 131
rect 2262 135 2268 136
rect 2262 131 2263 135
rect 2267 131 2268 135
rect 2262 130 2268 131
rect 2366 135 2372 136
rect 2366 131 2367 135
rect 2371 131 2372 135
rect 2366 130 2372 131
rect 2486 135 2492 136
rect 2486 131 2487 135
rect 2491 131 2492 135
rect 2486 130 2492 131
rect 2614 135 2620 136
rect 2614 131 2615 135
rect 2619 131 2620 135
rect 2614 130 2620 131
rect 2742 135 2748 136
rect 2742 131 2743 135
rect 2747 131 2748 135
rect 2742 130 2748 131
rect 2870 135 2876 136
rect 2870 131 2871 135
rect 2875 131 2876 135
rect 2870 130 2876 131
rect 2990 135 2996 136
rect 2990 131 2991 135
rect 2995 131 2996 135
rect 2990 130 2996 131
rect 3110 135 3116 136
rect 3110 131 3111 135
rect 3115 131 3116 135
rect 3110 130 3116 131
rect 3222 135 3228 136
rect 3222 131 3223 135
rect 3227 131 3228 135
rect 3222 130 3228 131
rect 3326 135 3332 136
rect 3326 131 3327 135
rect 3331 131 3332 135
rect 3326 130 3332 131
rect 3430 135 3436 136
rect 3430 131 3431 135
rect 3435 131 3436 135
rect 3430 130 3436 131
rect 3534 135 3540 136
rect 3534 131 3535 135
rect 3539 131 3540 135
rect 3534 130 3540 131
rect 3638 135 3644 136
rect 3638 131 3639 135
rect 3643 131 3644 135
rect 3638 130 3644 131
rect 3742 135 3748 136
rect 3742 131 3743 135
rect 3747 131 3748 135
rect 3742 130 3748 131
rect 3838 135 3844 136
rect 3838 131 3839 135
rect 3843 131 3844 135
rect 3942 132 3943 136
rect 3947 132 3948 136
rect 3942 131 3948 132
rect 3838 130 3844 131
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2006 118 2012 119
rect 2046 119 2052 120
rect 1902 115 1908 116
rect 2046 115 2047 119
rect 2051 115 2052 119
rect 3942 119 3948 120
rect 2046 114 2052 115
rect 2070 116 2076 117
rect 2070 112 2071 116
rect 2075 112 2076 116
rect 2070 111 2076 112
rect 2166 116 2172 117
rect 2166 112 2167 116
rect 2171 112 2172 116
rect 2166 111 2172 112
rect 2262 116 2268 117
rect 2262 112 2263 116
rect 2267 112 2268 116
rect 2262 111 2268 112
rect 2366 116 2372 117
rect 2366 112 2367 116
rect 2371 112 2372 116
rect 2366 111 2372 112
rect 2486 116 2492 117
rect 2486 112 2487 116
rect 2491 112 2492 116
rect 2486 111 2492 112
rect 2614 116 2620 117
rect 2614 112 2615 116
rect 2619 112 2620 116
rect 2614 111 2620 112
rect 2742 116 2748 117
rect 2742 112 2743 116
rect 2747 112 2748 116
rect 2742 111 2748 112
rect 2870 116 2876 117
rect 2870 112 2871 116
rect 2875 112 2876 116
rect 2870 111 2876 112
rect 2990 116 2996 117
rect 2990 112 2991 116
rect 2995 112 2996 116
rect 2990 111 2996 112
rect 3110 116 3116 117
rect 3110 112 3111 116
rect 3115 112 3116 116
rect 3110 111 3116 112
rect 3222 116 3228 117
rect 3222 112 3223 116
rect 3227 112 3228 116
rect 3222 111 3228 112
rect 3326 116 3332 117
rect 3326 112 3327 116
rect 3331 112 3332 116
rect 3326 111 3332 112
rect 3430 116 3436 117
rect 3430 112 3431 116
rect 3435 112 3436 116
rect 3430 111 3436 112
rect 3534 116 3540 117
rect 3534 112 3535 116
rect 3539 112 3540 116
rect 3534 111 3540 112
rect 3638 116 3644 117
rect 3638 112 3639 116
rect 3643 112 3644 116
rect 3638 111 3644 112
rect 3742 116 3748 117
rect 3742 112 3743 116
rect 3747 112 3748 116
rect 3742 111 3748 112
rect 3838 116 3844 117
rect 3838 112 3839 116
rect 3843 112 3844 116
rect 3942 115 3943 119
rect 3947 115 3948 119
rect 3942 114 3948 115
rect 3838 111 3844 112
<< m3c >>
rect 2047 4000 2051 4004
rect 2071 3999 2075 4003
rect 3943 4000 3947 4004
rect 111 3980 115 3984
rect 151 3979 155 3983
rect 279 3979 283 3983
rect 431 3979 435 3983
rect 607 3979 611 3983
rect 791 3979 795 3983
rect 975 3979 979 3983
rect 1151 3979 1155 3983
rect 1311 3979 1315 3983
rect 1471 3979 1475 3983
rect 1623 3979 1627 3983
rect 1775 3979 1779 3983
rect 1903 3979 1907 3983
rect 2007 3980 2011 3984
rect 2047 3983 2051 3987
rect 2071 3980 2075 3984
rect 3943 3983 3947 3987
rect 111 3963 115 3967
rect 151 3960 155 3964
rect 279 3960 283 3964
rect 431 3960 435 3964
rect 607 3960 611 3964
rect 791 3960 795 3964
rect 975 3960 979 3964
rect 1151 3960 1155 3964
rect 1311 3960 1315 3964
rect 1471 3960 1475 3964
rect 1623 3960 1627 3964
rect 1775 3960 1779 3964
rect 1903 3960 1907 3964
rect 2007 3963 2011 3967
rect 2047 3917 2051 3921
rect 2079 3920 2083 3924
rect 2215 3920 2219 3924
rect 2359 3920 2363 3924
rect 2503 3920 2507 3924
rect 2647 3920 2651 3924
rect 2791 3920 2795 3924
rect 2927 3920 2931 3924
rect 3055 3920 3059 3924
rect 3175 3920 3179 3924
rect 3295 3920 3299 3924
rect 3415 3920 3419 3924
rect 3535 3920 3539 3924
rect 3943 3917 3947 3921
rect 111 3897 115 3901
rect 303 3900 307 3904
rect 423 3900 427 3904
rect 551 3900 555 3904
rect 687 3900 691 3904
rect 815 3900 819 3904
rect 943 3900 947 3904
rect 1071 3900 1075 3904
rect 1199 3900 1203 3904
rect 1327 3900 1331 3904
rect 1463 3900 1467 3904
rect 2007 3897 2011 3901
rect 2047 3900 2051 3904
rect 2079 3901 2083 3905
rect 2215 3901 2219 3905
rect 2359 3901 2363 3905
rect 2503 3901 2507 3905
rect 2647 3901 2651 3905
rect 2791 3901 2795 3905
rect 2927 3901 2931 3905
rect 3055 3901 3059 3905
rect 3175 3901 3179 3905
rect 3295 3901 3299 3905
rect 3415 3901 3419 3905
rect 3535 3901 3539 3905
rect 3943 3900 3947 3904
rect 111 3880 115 3884
rect 303 3881 307 3885
rect 423 3881 427 3885
rect 551 3881 555 3885
rect 687 3881 691 3885
rect 815 3881 819 3885
rect 943 3881 947 3885
rect 1071 3881 1075 3885
rect 1199 3881 1203 3885
rect 1327 3881 1331 3885
rect 1463 3881 1467 3885
rect 2007 3880 2011 3884
rect 2047 3848 2051 3852
rect 2255 3847 2259 3851
rect 2383 3847 2387 3851
rect 2519 3847 2523 3851
rect 2671 3847 2675 3851
rect 2831 3847 2835 3851
rect 2991 3847 2995 3851
rect 3159 3847 3163 3851
rect 3327 3847 3331 3851
rect 3495 3847 3499 3851
rect 3663 3847 3667 3851
rect 3943 3848 3947 3852
rect 2047 3831 2051 3835
rect 111 3824 115 3828
rect 415 3823 419 3827
rect 567 3823 571 3827
rect 727 3823 731 3827
rect 887 3823 891 3827
rect 1039 3823 1043 3827
rect 1191 3823 1195 3827
rect 1343 3823 1347 3827
rect 1495 3823 1499 3827
rect 1647 3823 1651 3827
rect 2007 3824 2011 3828
rect 2255 3828 2259 3832
rect 2383 3828 2387 3832
rect 2519 3828 2523 3832
rect 2671 3828 2675 3832
rect 2831 3828 2835 3832
rect 2991 3828 2995 3832
rect 3159 3828 3163 3832
rect 3327 3828 3331 3832
rect 3495 3828 3499 3832
rect 3663 3828 3667 3832
rect 3943 3831 3947 3835
rect 111 3807 115 3811
rect 415 3804 419 3808
rect 567 3804 571 3808
rect 727 3804 731 3808
rect 887 3804 891 3808
rect 1039 3804 1043 3808
rect 1191 3804 1195 3808
rect 1343 3804 1347 3808
rect 1495 3804 1499 3808
rect 1647 3804 1651 3808
rect 2007 3807 2011 3811
rect 2047 3765 2051 3769
rect 2071 3768 2075 3772
rect 2199 3768 2203 3772
rect 2375 3768 2379 3772
rect 2559 3768 2563 3772
rect 2751 3768 2755 3772
rect 2951 3768 2955 3772
rect 3143 3768 3147 3772
rect 3335 3768 3339 3772
rect 3535 3768 3539 3772
rect 3735 3768 3739 3772
rect 3943 3765 3947 3769
rect 2047 3748 2051 3752
rect 2071 3749 2075 3753
rect 2199 3749 2203 3753
rect 2375 3749 2379 3753
rect 2559 3749 2563 3753
rect 2751 3749 2755 3753
rect 2951 3749 2955 3753
rect 3143 3749 3147 3753
rect 3335 3749 3339 3753
rect 3535 3749 3539 3753
rect 3735 3749 3739 3753
rect 3943 3748 3947 3752
rect 111 3737 115 3741
rect 399 3740 403 3744
rect 567 3740 571 3744
rect 751 3740 755 3744
rect 935 3740 939 3744
rect 1127 3740 1131 3744
rect 1311 3740 1315 3744
rect 1503 3740 1507 3744
rect 1695 3740 1699 3744
rect 1887 3740 1891 3744
rect 2007 3737 2011 3741
rect 111 3720 115 3724
rect 399 3721 403 3725
rect 567 3721 571 3725
rect 751 3721 755 3725
rect 935 3721 939 3725
rect 1127 3721 1131 3725
rect 1311 3721 1315 3725
rect 1503 3721 1507 3725
rect 1695 3721 1699 3725
rect 1887 3721 1891 3725
rect 2007 3720 2011 3724
rect 2047 3684 2051 3688
rect 2071 3683 2075 3687
rect 2263 3683 2267 3687
rect 2479 3683 2483 3687
rect 2695 3683 2699 3687
rect 2911 3683 2915 3687
rect 3119 3683 3123 3687
rect 3319 3683 3323 3687
rect 3519 3683 3523 3687
rect 3727 3683 3731 3687
rect 3943 3684 3947 3688
rect 2047 3667 2051 3671
rect 2071 3664 2075 3668
rect 2263 3664 2267 3668
rect 2479 3664 2483 3668
rect 2695 3664 2699 3668
rect 2911 3664 2915 3668
rect 3119 3664 3123 3668
rect 3319 3664 3323 3668
rect 3519 3664 3523 3668
rect 3727 3664 3731 3668
rect 3943 3667 3947 3671
rect 111 3656 115 3660
rect 367 3655 371 3659
rect 519 3655 523 3659
rect 679 3655 683 3659
rect 847 3655 851 3659
rect 1015 3655 1019 3659
rect 1175 3655 1179 3659
rect 1327 3655 1331 3659
rect 1479 3655 1483 3659
rect 1631 3655 1635 3659
rect 1791 3655 1795 3659
rect 2007 3656 2011 3660
rect 111 3639 115 3643
rect 367 3636 371 3640
rect 519 3636 523 3640
rect 679 3636 683 3640
rect 847 3636 851 3640
rect 1015 3636 1019 3640
rect 1175 3636 1179 3640
rect 1327 3636 1331 3640
rect 1479 3636 1483 3640
rect 1631 3636 1635 3640
rect 1791 3636 1795 3640
rect 2007 3639 2011 3643
rect 2047 3597 2051 3601
rect 2111 3600 2115 3604
rect 2271 3600 2275 3604
rect 2455 3600 2459 3604
rect 2655 3600 2659 3604
rect 2871 3600 2875 3604
rect 3095 3600 3099 3604
rect 3327 3600 3331 3604
rect 3567 3600 3571 3604
rect 3943 3597 3947 3601
rect 2047 3580 2051 3584
rect 2111 3581 2115 3585
rect 2271 3581 2275 3585
rect 2455 3581 2459 3585
rect 2655 3581 2659 3585
rect 2871 3581 2875 3585
rect 3095 3581 3099 3585
rect 3327 3581 3331 3585
rect 3567 3581 3571 3585
rect 3943 3580 3947 3584
rect 111 3565 115 3569
rect 271 3568 275 3572
rect 415 3568 419 3572
rect 575 3568 579 3572
rect 735 3568 739 3572
rect 895 3568 899 3572
rect 1055 3568 1059 3572
rect 1215 3568 1219 3572
rect 1375 3568 1379 3572
rect 1543 3568 1547 3572
rect 2007 3565 2011 3569
rect 111 3548 115 3552
rect 271 3549 275 3553
rect 415 3549 419 3553
rect 575 3549 579 3553
rect 735 3549 739 3553
rect 895 3549 899 3553
rect 1055 3549 1059 3553
rect 1215 3549 1219 3553
rect 1375 3549 1379 3553
rect 1543 3549 1547 3553
rect 2007 3548 2011 3552
rect 2047 3512 2051 3516
rect 2287 3511 2291 3515
rect 2383 3511 2387 3515
rect 2479 3511 2483 3515
rect 2575 3511 2579 3515
rect 2671 3511 2675 3515
rect 2767 3511 2771 3515
rect 2871 3511 2875 3515
rect 2983 3511 2987 3515
rect 3103 3511 3107 3515
rect 3223 3511 3227 3515
rect 3351 3511 3355 3515
rect 3487 3511 3491 3515
rect 3943 3512 3947 3516
rect 2047 3495 2051 3499
rect 111 3488 115 3492
rect 159 3487 163 3491
rect 287 3487 291 3491
rect 423 3487 427 3491
rect 559 3487 563 3491
rect 695 3487 699 3491
rect 831 3487 835 3491
rect 967 3487 971 3491
rect 1095 3487 1099 3491
rect 1231 3487 1235 3491
rect 1367 3487 1371 3491
rect 2007 3488 2011 3492
rect 2287 3492 2291 3496
rect 2383 3492 2387 3496
rect 2479 3492 2483 3496
rect 2575 3492 2579 3496
rect 2671 3492 2675 3496
rect 2767 3492 2771 3496
rect 2871 3492 2875 3496
rect 2983 3492 2987 3496
rect 3103 3492 3107 3496
rect 3223 3492 3227 3496
rect 3351 3492 3355 3496
rect 3487 3492 3491 3496
rect 3943 3495 3947 3499
rect 111 3471 115 3475
rect 159 3468 163 3472
rect 287 3468 291 3472
rect 423 3468 427 3472
rect 559 3468 563 3472
rect 695 3468 699 3472
rect 831 3468 835 3472
rect 967 3468 971 3472
rect 1095 3468 1099 3472
rect 1231 3468 1235 3472
rect 1367 3468 1371 3472
rect 2007 3471 2011 3475
rect 2047 3429 2051 3433
rect 2487 3432 2491 3436
rect 2583 3432 2587 3436
rect 2679 3432 2683 3436
rect 2783 3432 2787 3436
rect 2895 3432 2899 3436
rect 3015 3432 3019 3436
rect 3143 3432 3147 3436
rect 3271 3432 3275 3436
rect 3407 3432 3411 3436
rect 3943 3429 3947 3433
rect 2047 3412 2051 3416
rect 2487 3413 2491 3417
rect 2583 3413 2587 3417
rect 2679 3413 2683 3417
rect 2783 3413 2787 3417
rect 2895 3413 2899 3417
rect 3015 3413 3019 3417
rect 3143 3413 3147 3417
rect 3271 3413 3275 3417
rect 3407 3413 3411 3417
rect 3943 3412 3947 3416
rect 111 3397 115 3401
rect 135 3400 139 3404
rect 247 3400 251 3404
rect 383 3400 387 3404
rect 527 3400 531 3404
rect 671 3400 675 3404
rect 815 3400 819 3404
rect 967 3400 971 3404
rect 1119 3400 1123 3404
rect 1271 3400 1275 3404
rect 2007 3397 2011 3401
rect 111 3380 115 3384
rect 135 3381 139 3385
rect 247 3381 251 3385
rect 383 3381 387 3385
rect 527 3381 531 3385
rect 671 3381 675 3385
rect 815 3381 819 3385
rect 967 3381 971 3385
rect 1119 3381 1123 3385
rect 1271 3381 1275 3385
rect 2007 3380 2011 3384
rect 2047 3352 2051 3356
rect 2351 3351 2355 3355
rect 2479 3351 2483 3355
rect 2615 3351 2619 3355
rect 2751 3351 2755 3355
rect 2887 3351 2891 3355
rect 3023 3351 3027 3355
rect 3159 3351 3163 3355
rect 3303 3351 3307 3355
rect 3943 3352 3947 3356
rect 2047 3335 2051 3339
rect 2351 3332 2355 3336
rect 2479 3332 2483 3336
rect 2615 3332 2619 3336
rect 2751 3332 2755 3336
rect 2887 3332 2891 3336
rect 3023 3332 3027 3336
rect 3159 3332 3163 3336
rect 3303 3332 3307 3336
rect 3943 3335 3947 3339
rect 111 3320 115 3324
rect 135 3319 139 3323
rect 263 3319 267 3323
rect 431 3319 435 3323
rect 599 3319 603 3323
rect 767 3319 771 3323
rect 927 3319 931 3323
rect 1087 3319 1091 3323
rect 1239 3319 1243 3323
rect 1391 3319 1395 3323
rect 1551 3319 1555 3323
rect 2007 3320 2011 3324
rect 111 3303 115 3307
rect 135 3300 139 3304
rect 263 3300 267 3304
rect 431 3300 435 3304
rect 599 3300 603 3304
rect 767 3300 771 3304
rect 927 3300 931 3304
rect 1087 3300 1091 3304
rect 1239 3300 1243 3304
rect 1391 3300 1395 3304
rect 1551 3300 1555 3304
rect 2007 3303 2011 3307
rect 2047 3265 2051 3269
rect 2127 3268 2131 3272
rect 2295 3268 2299 3272
rect 2455 3268 2459 3272
rect 2615 3268 2619 3272
rect 2775 3268 2779 3272
rect 2935 3268 2939 3272
rect 3095 3268 3099 3272
rect 3263 3268 3267 3272
rect 3943 3265 3947 3269
rect 2047 3248 2051 3252
rect 2127 3249 2131 3253
rect 2295 3249 2299 3253
rect 2455 3249 2459 3253
rect 2615 3249 2619 3253
rect 2775 3249 2779 3253
rect 2935 3249 2939 3253
rect 3095 3249 3099 3253
rect 3263 3249 3267 3253
rect 3943 3248 3947 3252
rect 111 3229 115 3233
rect 143 3232 147 3236
rect 295 3232 299 3236
rect 455 3232 459 3236
rect 623 3232 627 3236
rect 791 3232 795 3236
rect 959 3232 963 3236
rect 1127 3232 1131 3236
rect 1303 3232 1307 3236
rect 1479 3232 1483 3236
rect 2007 3229 2011 3233
rect 111 3212 115 3216
rect 143 3213 147 3217
rect 295 3213 299 3217
rect 455 3213 459 3217
rect 623 3213 627 3217
rect 791 3213 795 3217
rect 959 3213 963 3217
rect 1127 3213 1131 3217
rect 1303 3213 1307 3217
rect 1479 3213 1483 3217
rect 2007 3212 2011 3216
rect 2047 3196 2051 3200
rect 2071 3195 2075 3199
rect 2207 3195 2211 3199
rect 2375 3195 2379 3199
rect 2543 3195 2547 3199
rect 2703 3195 2707 3199
rect 2863 3195 2867 3199
rect 3015 3195 3019 3199
rect 3167 3195 3171 3199
rect 3327 3195 3331 3199
rect 3943 3196 3947 3200
rect 2047 3179 2051 3183
rect 2071 3176 2075 3180
rect 2207 3176 2211 3180
rect 2375 3176 2379 3180
rect 2543 3176 2547 3180
rect 2703 3176 2707 3180
rect 2863 3176 2867 3180
rect 3015 3176 3019 3180
rect 3167 3176 3171 3180
rect 3327 3176 3331 3180
rect 3943 3179 3947 3183
rect 111 3160 115 3164
rect 295 3159 299 3163
rect 431 3159 435 3163
rect 567 3159 571 3163
rect 703 3159 707 3163
rect 855 3159 859 3163
rect 1031 3159 1035 3163
rect 1231 3159 1235 3163
rect 1455 3159 1459 3163
rect 1687 3159 1691 3163
rect 1903 3159 1907 3163
rect 2007 3160 2011 3164
rect 111 3143 115 3147
rect 295 3140 299 3144
rect 431 3140 435 3144
rect 567 3140 571 3144
rect 703 3140 707 3144
rect 855 3140 859 3144
rect 1031 3140 1035 3144
rect 1231 3140 1235 3144
rect 1455 3140 1459 3144
rect 1687 3140 1691 3144
rect 1903 3140 1907 3144
rect 2007 3143 2011 3147
rect 2047 3109 2051 3113
rect 2071 3112 2075 3116
rect 2343 3112 2347 3116
rect 2631 3112 2635 3116
rect 2903 3112 2907 3116
rect 3175 3112 3179 3116
rect 3447 3112 3451 3116
rect 3943 3109 3947 3113
rect 2047 3092 2051 3096
rect 2071 3093 2075 3097
rect 2343 3093 2347 3097
rect 2631 3093 2635 3097
rect 2903 3093 2907 3097
rect 3175 3093 3179 3097
rect 3447 3093 3451 3097
rect 3943 3092 3947 3096
rect 111 3077 115 3081
rect 311 3080 315 3084
rect 407 3080 411 3084
rect 503 3080 507 3084
rect 599 3080 603 3084
rect 695 3080 699 3084
rect 807 3080 811 3084
rect 943 3080 947 3084
rect 1087 3080 1091 3084
rect 1247 3080 1251 3084
rect 1407 3080 1411 3084
rect 1575 3080 1579 3084
rect 1751 3080 1755 3084
rect 1903 3080 1907 3084
rect 2007 3077 2011 3081
rect 111 3060 115 3064
rect 311 3061 315 3065
rect 407 3061 411 3065
rect 503 3061 507 3065
rect 599 3061 603 3065
rect 695 3061 699 3065
rect 807 3061 811 3065
rect 943 3061 947 3065
rect 1087 3061 1091 3065
rect 1247 3061 1251 3065
rect 1407 3061 1411 3065
rect 1575 3061 1579 3065
rect 1751 3061 1755 3065
rect 1903 3061 1907 3065
rect 2007 3060 2011 3064
rect 2047 3036 2051 3040
rect 2487 3035 2491 3039
rect 2615 3035 2619 3039
rect 2743 3035 2747 3039
rect 2863 3035 2867 3039
rect 2983 3035 2987 3039
rect 3103 3035 3107 3039
rect 3215 3035 3219 3039
rect 3327 3035 3331 3039
rect 3431 3035 3435 3039
rect 3535 3035 3539 3039
rect 3639 3035 3643 3039
rect 3743 3035 3747 3039
rect 3839 3035 3843 3039
rect 3943 3036 3947 3040
rect 2047 3019 2051 3023
rect 2487 3016 2491 3020
rect 2615 3016 2619 3020
rect 2743 3016 2747 3020
rect 2863 3016 2867 3020
rect 2983 3016 2987 3020
rect 3103 3016 3107 3020
rect 3215 3016 3219 3020
rect 3327 3016 3331 3020
rect 3431 3016 3435 3020
rect 3535 3016 3539 3020
rect 3639 3016 3643 3020
rect 3743 3016 3747 3020
rect 3839 3016 3843 3020
rect 3943 3019 3947 3023
rect 111 3008 115 3012
rect 423 3007 427 3011
rect 519 3007 523 3011
rect 615 3007 619 3011
rect 711 3007 715 3011
rect 815 3007 819 3011
rect 935 3007 939 3011
rect 1055 3007 1059 3011
rect 1183 3007 1187 3011
rect 1311 3007 1315 3011
rect 1431 3007 1435 3011
rect 1551 3007 1555 3011
rect 1671 3007 1675 3011
rect 1799 3007 1803 3011
rect 1903 3007 1907 3011
rect 2007 3008 2011 3012
rect 111 2991 115 2995
rect 423 2988 427 2992
rect 519 2988 523 2992
rect 615 2988 619 2992
rect 711 2988 715 2992
rect 815 2988 819 2992
rect 935 2988 939 2992
rect 1055 2988 1059 2992
rect 1183 2988 1187 2992
rect 1311 2988 1315 2992
rect 1431 2988 1435 2992
rect 1551 2988 1555 2992
rect 1671 2988 1675 2992
rect 1799 2988 1803 2992
rect 1903 2988 1907 2992
rect 2007 2991 2011 2995
rect 2047 2949 2051 2953
rect 2407 2952 2411 2956
rect 2575 2952 2579 2956
rect 2767 2952 2771 2956
rect 2967 2952 2971 2956
rect 3183 2952 3187 2956
rect 3399 2952 3403 2956
rect 3623 2952 3627 2956
rect 3839 2952 3843 2956
rect 3943 2949 3947 2953
rect 2047 2932 2051 2936
rect 2407 2933 2411 2937
rect 2575 2933 2579 2937
rect 2767 2933 2771 2937
rect 2967 2933 2971 2937
rect 3183 2933 3187 2937
rect 3399 2933 3403 2937
rect 3623 2933 3627 2937
rect 3839 2933 3843 2937
rect 3943 2932 3947 2936
rect 111 2901 115 2905
rect 1479 2904 1483 2908
rect 1575 2904 1579 2908
rect 1671 2904 1675 2908
rect 1767 2904 1771 2908
rect 1863 2904 1867 2908
rect 2007 2901 2011 2905
rect 111 2884 115 2888
rect 1479 2885 1483 2889
rect 1575 2885 1579 2889
rect 1671 2885 1675 2889
rect 1767 2885 1771 2889
rect 1863 2885 1867 2889
rect 2007 2884 2011 2888
rect 2047 2864 2051 2868
rect 2551 2863 2555 2867
rect 2671 2863 2675 2867
rect 2799 2863 2803 2867
rect 2927 2863 2931 2867
rect 3055 2863 3059 2867
rect 3183 2863 3187 2867
rect 3311 2863 3315 2867
rect 3439 2863 3443 2867
rect 3575 2863 3579 2867
rect 3943 2864 3947 2868
rect 2047 2847 2051 2851
rect 2551 2844 2555 2848
rect 2671 2844 2675 2848
rect 2799 2844 2803 2848
rect 2927 2844 2931 2848
rect 3055 2844 3059 2848
rect 3183 2844 3187 2848
rect 3311 2844 3315 2848
rect 3439 2844 3443 2848
rect 3575 2844 3579 2848
rect 3943 2847 3947 2851
rect 111 2824 115 2828
rect 279 2823 283 2827
rect 447 2823 451 2827
rect 631 2823 635 2827
rect 815 2823 819 2827
rect 999 2823 1003 2827
rect 1183 2823 1187 2827
rect 1359 2823 1363 2827
rect 1527 2823 1531 2827
rect 1695 2823 1699 2827
rect 1863 2823 1867 2827
rect 2007 2824 2011 2828
rect 111 2807 115 2811
rect 279 2804 283 2808
rect 447 2804 451 2808
rect 631 2804 635 2808
rect 815 2804 819 2808
rect 999 2804 1003 2808
rect 1183 2804 1187 2808
rect 1359 2804 1363 2808
rect 1527 2804 1531 2808
rect 1695 2804 1699 2808
rect 1863 2804 1867 2808
rect 2007 2807 2011 2811
rect 2047 2781 2051 2785
rect 2439 2784 2443 2788
rect 2567 2784 2571 2788
rect 2695 2784 2699 2788
rect 2831 2784 2835 2788
rect 2967 2784 2971 2788
rect 3103 2784 3107 2788
rect 3247 2784 3251 2788
rect 3391 2784 3395 2788
rect 3543 2784 3547 2788
rect 3703 2784 3707 2788
rect 3839 2784 3843 2788
rect 3943 2781 3947 2785
rect 2047 2764 2051 2768
rect 2439 2765 2443 2769
rect 2567 2765 2571 2769
rect 2695 2765 2699 2769
rect 2831 2765 2835 2769
rect 2967 2765 2971 2769
rect 3103 2765 3107 2769
rect 3247 2765 3251 2769
rect 3391 2765 3395 2769
rect 3543 2765 3547 2769
rect 3703 2765 3707 2769
rect 3839 2765 3843 2769
rect 3943 2764 3947 2768
rect 111 2741 115 2745
rect 239 2744 243 2748
rect 351 2744 355 2748
rect 471 2744 475 2748
rect 607 2744 611 2748
rect 743 2744 747 2748
rect 879 2744 883 2748
rect 1015 2744 1019 2748
rect 1151 2744 1155 2748
rect 1287 2744 1291 2748
rect 1423 2744 1427 2748
rect 1567 2744 1571 2748
rect 2007 2741 2011 2745
rect 111 2724 115 2728
rect 239 2725 243 2729
rect 351 2725 355 2729
rect 471 2725 475 2729
rect 607 2725 611 2729
rect 743 2725 747 2729
rect 879 2725 883 2729
rect 1015 2725 1019 2729
rect 1151 2725 1155 2729
rect 1287 2725 1291 2729
rect 1423 2725 1427 2729
rect 1567 2725 1571 2729
rect 2007 2724 2011 2728
rect 2047 2704 2051 2708
rect 2335 2703 2339 2707
rect 2495 2703 2499 2707
rect 2663 2703 2667 2707
rect 2831 2703 2835 2707
rect 2999 2703 3003 2707
rect 3167 2703 3171 2707
rect 3335 2703 3339 2707
rect 3511 2703 3515 2707
rect 3687 2703 3691 2707
rect 3839 2703 3843 2707
rect 3943 2704 3947 2708
rect 2047 2687 2051 2691
rect 2335 2684 2339 2688
rect 2495 2684 2499 2688
rect 2663 2684 2667 2688
rect 2831 2684 2835 2688
rect 2999 2684 3003 2688
rect 3167 2684 3171 2688
rect 3335 2684 3339 2688
rect 3511 2684 3515 2688
rect 3687 2684 3691 2688
rect 3839 2684 3843 2688
rect 3943 2687 3947 2691
rect 111 2672 115 2676
rect 223 2671 227 2675
rect 367 2671 371 2675
rect 503 2671 507 2675
rect 639 2671 643 2675
rect 767 2671 771 2675
rect 887 2671 891 2675
rect 999 2671 1003 2675
rect 1111 2671 1115 2675
rect 1231 2671 1235 2675
rect 1351 2671 1355 2675
rect 2007 2672 2011 2676
rect 111 2655 115 2659
rect 223 2652 227 2656
rect 367 2652 371 2656
rect 503 2652 507 2656
rect 639 2652 643 2656
rect 767 2652 771 2656
rect 887 2652 891 2656
rect 999 2652 1003 2656
rect 1111 2652 1115 2656
rect 1231 2652 1235 2656
rect 1351 2652 1355 2656
rect 2007 2655 2011 2659
rect 2047 2617 2051 2621
rect 2127 2620 2131 2624
rect 2279 2620 2283 2624
rect 2447 2620 2451 2624
rect 2623 2620 2627 2624
rect 2807 2620 2811 2624
rect 2991 2620 2995 2624
rect 3175 2620 3179 2624
rect 3351 2620 3355 2624
rect 3519 2620 3523 2624
rect 3687 2620 3691 2624
rect 3839 2620 3843 2624
rect 3943 2617 3947 2621
rect 2047 2600 2051 2604
rect 2127 2601 2131 2605
rect 2279 2601 2283 2605
rect 2447 2601 2451 2605
rect 2623 2601 2627 2605
rect 2807 2601 2811 2605
rect 2991 2601 2995 2605
rect 3175 2601 3179 2605
rect 3351 2601 3355 2605
rect 3519 2601 3523 2605
rect 3687 2601 3691 2605
rect 3839 2601 3843 2605
rect 3943 2600 3947 2604
rect 111 2589 115 2593
rect 175 2592 179 2596
rect 367 2592 371 2596
rect 543 2592 547 2596
rect 711 2592 715 2596
rect 863 2592 867 2596
rect 1007 2592 1011 2596
rect 1143 2592 1147 2596
rect 1279 2592 1283 2596
rect 1423 2592 1427 2596
rect 2007 2589 2011 2593
rect 111 2572 115 2576
rect 175 2573 179 2577
rect 367 2573 371 2577
rect 543 2573 547 2577
rect 711 2573 715 2577
rect 863 2573 867 2577
rect 1007 2573 1011 2577
rect 1143 2573 1147 2577
rect 1279 2573 1283 2577
rect 1423 2573 1427 2577
rect 2007 2572 2011 2576
rect 2047 2540 2051 2544
rect 2071 2539 2075 2543
rect 2183 2539 2187 2543
rect 2319 2539 2323 2543
rect 2471 2539 2475 2543
rect 2639 2539 2643 2543
rect 2823 2539 2827 2543
rect 3031 2539 3035 2543
rect 3263 2539 3267 2543
rect 3503 2539 3507 2543
rect 3743 2539 3747 2543
rect 3943 2540 3947 2544
rect 2047 2523 2051 2527
rect 111 2516 115 2520
rect 135 2515 139 2519
rect 271 2515 275 2519
rect 439 2515 443 2519
rect 607 2515 611 2519
rect 775 2515 779 2519
rect 927 2515 931 2519
rect 1079 2515 1083 2519
rect 1223 2515 1227 2519
rect 1359 2515 1363 2519
rect 1495 2515 1499 2519
rect 1639 2515 1643 2519
rect 2007 2516 2011 2520
rect 2071 2520 2075 2524
rect 2183 2520 2187 2524
rect 2319 2520 2323 2524
rect 2471 2520 2475 2524
rect 2639 2520 2643 2524
rect 2823 2520 2827 2524
rect 3031 2520 3035 2524
rect 3263 2520 3267 2524
rect 3503 2520 3507 2524
rect 3743 2520 3747 2524
rect 3943 2523 3947 2527
rect 111 2499 115 2503
rect 135 2496 139 2500
rect 271 2496 275 2500
rect 439 2496 443 2500
rect 607 2496 611 2500
rect 775 2496 779 2500
rect 927 2496 931 2500
rect 1079 2496 1083 2500
rect 1223 2496 1227 2500
rect 1359 2496 1363 2500
rect 1495 2496 1499 2500
rect 1639 2496 1643 2500
rect 2007 2499 2011 2503
rect 2047 2453 2051 2457
rect 2071 2456 2075 2460
rect 2215 2456 2219 2460
rect 2383 2456 2387 2460
rect 2559 2456 2563 2460
rect 2751 2456 2755 2460
rect 2951 2456 2955 2460
rect 3167 2456 3171 2460
rect 3391 2456 3395 2460
rect 3623 2456 3627 2460
rect 3839 2456 3843 2460
rect 3943 2453 3947 2457
rect 111 2429 115 2433
rect 135 2432 139 2436
rect 311 2432 315 2436
rect 511 2432 515 2436
rect 711 2432 715 2436
rect 903 2432 907 2436
rect 1079 2432 1083 2436
rect 1239 2432 1243 2436
rect 1391 2432 1395 2436
rect 1527 2432 1531 2436
rect 1663 2432 1667 2436
rect 1791 2432 1795 2436
rect 1903 2432 1907 2436
rect 2047 2436 2051 2440
rect 2071 2437 2075 2441
rect 2215 2437 2219 2441
rect 2383 2437 2387 2441
rect 2559 2437 2563 2441
rect 2751 2437 2755 2441
rect 2951 2437 2955 2441
rect 3167 2437 3171 2441
rect 3391 2437 3395 2441
rect 3623 2437 3627 2441
rect 3839 2437 3843 2441
rect 3943 2436 3947 2440
rect 2007 2429 2011 2433
rect 111 2412 115 2416
rect 135 2413 139 2417
rect 311 2413 315 2417
rect 511 2413 515 2417
rect 711 2413 715 2417
rect 903 2413 907 2417
rect 1079 2413 1083 2417
rect 1239 2413 1243 2417
rect 1391 2413 1395 2417
rect 1527 2413 1531 2417
rect 1663 2413 1667 2417
rect 1791 2413 1795 2417
rect 1903 2413 1907 2417
rect 2007 2412 2011 2416
rect 2047 2368 2051 2372
rect 2071 2367 2075 2371
rect 2247 2367 2251 2371
rect 2431 2367 2435 2371
rect 2607 2367 2611 2371
rect 2775 2367 2779 2371
rect 2935 2367 2939 2371
rect 3103 2367 3107 2371
rect 3943 2368 3947 2372
rect 111 2360 115 2364
rect 135 2359 139 2363
rect 327 2359 331 2363
rect 551 2359 555 2363
rect 767 2359 771 2363
rect 975 2359 979 2363
rect 1175 2359 1179 2363
rect 1367 2359 1371 2363
rect 1551 2359 1555 2363
rect 1735 2359 1739 2363
rect 1903 2359 1907 2363
rect 2007 2360 2011 2364
rect 2047 2351 2051 2355
rect 2071 2348 2075 2352
rect 111 2343 115 2347
rect 2247 2348 2251 2352
rect 2431 2348 2435 2352
rect 2607 2348 2611 2352
rect 2775 2348 2779 2352
rect 2935 2348 2939 2352
rect 3103 2348 3107 2352
rect 3943 2351 3947 2355
rect 135 2340 139 2344
rect 327 2340 331 2344
rect 551 2340 555 2344
rect 767 2340 771 2344
rect 975 2340 979 2344
rect 1175 2340 1179 2344
rect 1367 2340 1371 2344
rect 1551 2340 1555 2344
rect 1735 2340 1739 2344
rect 1903 2340 1907 2344
rect 2007 2343 2011 2347
rect 2047 2285 2051 2289
rect 2071 2288 2075 2292
rect 2175 2288 2179 2292
rect 2311 2288 2315 2292
rect 2447 2288 2451 2292
rect 2591 2288 2595 2292
rect 2751 2288 2755 2292
rect 2935 2288 2939 2292
rect 3143 2288 3147 2292
rect 3375 2288 3379 2292
rect 3615 2288 3619 2292
rect 3839 2288 3843 2292
rect 3943 2285 3947 2289
rect 111 2269 115 2273
rect 135 2272 139 2276
rect 271 2272 275 2276
rect 431 2272 435 2276
rect 591 2272 595 2276
rect 751 2272 755 2276
rect 919 2272 923 2276
rect 1087 2272 1091 2276
rect 1263 2272 1267 2276
rect 1447 2272 1451 2276
rect 1631 2272 1635 2276
rect 1815 2272 1819 2276
rect 2007 2269 2011 2273
rect 2047 2268 2051 2272
rect 2071 2269 2075 2273
rect 2175 2269 2179 2273
rect 2311 2269 2315 2273
rect 2447 2269 2451 2273
rect 2591 2269 2595 2273
rect 2751 2269 2755 2273
rect 2935 2269 2939 2273
rect 3143 2269 3147 2273
rect 3375 2269 3379 2273
rect 3615 2269 3619 2273
rect 3839 2269 3843 2273
rect 3943 2268 3947 2272
rect 111 2252 115 2256
rect 135 2253 139 2257
rect 271 2253 275 2257
rect 431 2253 435 2257
rect 591 2253 595 2257
rect 751 2253 755 2257
rect 919 2253 923 2257
rect 1087 2253 1091 2257
rect 1263 2253 1267 2257
rect 1447 2253 1451 2257
rect 1631 2253 1635 2257
rect 1815 2253 1819 2257
rect 2007 2252 2011 2256
rect 2047 2208 2051 2212
rect 2111 2207 2115 2211
rect 2255 2207 2259 2211
rect 2407 2207 2411 2211
rect 2559 2207 2563 2211
rect 2719 2207 2723 2211
rect 2879 2207 2883 2211
rect 3047 2207 3051 2211
rect 3223 2207 3227 2211
rect 3407 2207 3411 2211
rect 3591 2207 3595 2211
rect 3783 2207 3787 2211
rect 3943 2208 3947 2212
rect 111 2200 115 2204
rect 159 2199 163 2203
rect 327 2199 331 2203
rect 495 2199 499 2203
rect 679 2199 683 2203
rect 879 2199 883 2203
rect 1095 2199 1099 2203
rect 1327 2199 1331 2203
rect 1567 2199 1571 2203
rect 1815 2199 1819 2203
rect 2007 2200 2011 2204
rect 2047 2191 2051 2195
rect 2111 2188 2115 2192
rect 111 2183 115 2187
rect 2255 2188 2259 2192
rect 2407 2188 2411 2192
rect 2559 2188 2563 2192
rect 2719 2188 2723 2192
rect 2879 2188 2883 2192
rect 3047 2188 3051 2192
rect 3223 2188 3227 2192
rect 3407 2188 3411 2192
rect 3591 2188 3595 2192
rect 3783 2188 3787 2192
rect 3943 2191 3947 2195
rect 159 2180 163 2184
rect 327 2180 331 2184
rect 495 2180 499 2184
rect 679 2180 683 2184
rect 879 2180 883 2184
rect 1095 2180 1099 2184
rect 1327 2180 1331 2184
rect 1567 2180 1571 2184
rect 1815 2180 1819 2184
rect 2007 2183 2011 2187
rect 111 2117 115 2121
rect 223 2120 227 2124
rect 359 2120 363 2124
rect 495 2120 499 2124
rect 639 2120 643 2124
rect 783 2120 787 2124
rect 935 2120 939 2124
rect 1095 2120 1099 2124
rect 1263 2120 1267 2124
rect 1447 2120 1451 2124
rect 1631 2120 1635 2124
rect 1823 2120 1827 2124
rect 2007 2117 2011 2121
rect 2047 2113 2051 2117
rect 2287 2116 2291 2120
rect 2431 2116 2435 2120
rect 2583 2116 2587 2120
rect 2735 2116 2739 2120
rect 2887 2116 2891 2120
rect 3047 2116 3051 2120
rect 3207 2116 3211 2120
rect 3367 2116 3371 2120
rect 3527 2116 3531 2120
rect 3695 2116 3699 2120
rect 3839 2116 3843 2120
rect 3943 2113 3947 2117
rect 111 2100 115 2104
rect 223 2101 227 2105
rect 359 2101 363 2105
rect 495 2101 499 2105
rect 639 2101 643 2105
rect 783 2101 787 2105
rect 935 2101 939 2105
rect 1095 2101 1099 2105
rect 1263 2101 1267 2105
rect 1447 2101 1451 2105
rect 1631 2101 1635 2105
rect 1823 2101 1827 2105
rect 2007 2100 2011 2104
rect 2047 2096 2051 2100
rect 2287 2097 2291 2101
rect 2431 2097 2435 2101
rect 2583 2097 2587 2101
rect 2735 2097 2739 2101
rect 2887 2097 2891 2101
rect 3047 2097 3051 2101
rect 3207 2097 3211 2101
rect 3367 2097 3371 2101
rect 3527 2097 3531 2101
rect 3695 2097 3699 2101
rect 3839 2097 3843 2101
rect 3943 2096 3947 2100
rect 111 2040 115 2044
rect 375 2039 379 2043
rect 495 2039 499 2043
rect 615 2039 619 2043
rect 751 2039 755 2043
rect 895 2039 899 2043
rect 1047 2039 1051 2043
rect 1215 2039 1219 2043
rect 1399 2039 1403 2043
rect 1583 2039 1587 2043
rect 1775 2039 1779 2043
rect 2007 2040 2011 2044
rect 2047 2036 2051 2040
rect 2503 2035 2507 2039
rect 2671 2035 2675 2039
rect 2839 2035 2843 2039
rect 3007 2035 3011 2039
rect 3167 2035 3171 2039
rect 3311 2035 3315 2039
rect 3455 2035 3459 2039
rect 3591 2035 3595 2039
rect 3727 2035 3731 2039
rect 3839 2035 3843 2039
rect 3943 2036 3947 2040
rect 111 2023 115 2027
rect 375 2020 379 2024
rect 495 2020 499 2024
rect 615 2020 619 2024
rect 751 2020 755 2024
rect 895 2020 899 2024
rect 1047 2020 1051 2024
rect 1215 2020 1219 2024
rect 1399 2020 1403 2024
rect 1583 2020 1587 2024
rect 1775 2020 1779 2024
rect 2007 2023 2011 2027
rect 2047 2019 2051 2023
rect 2503 2016 2507 2020
rect 2671 2016 2675 2020
rect 2839 2016 2843 2020
rect 3007 2016 3011 2020
rect 3167 2016 3171 2020
rect 3311 2016 3315 2020
rect 3455 2016 3459 2020
rect 3591 2016 3595 2020
rect 3727 2016 3731 2020
rect 3839 2016 3843 2020
rect 3943 2019 3947 2023
rect 111 1949 115 1953
rect 511 1952 515 1956
rect 623 1952 627 1956
rect 743 1952 747 1956
rect 871 1952 875 1956
rect 1007 1952 1011 1956
rect 1143 1952 1147 1956
rect 1279 1952 1283 1956
rect 1415 1952 1419 1956
rect 1559 1952 1563 1956
rect 1703 1952 1707 1956
rect 2007 1949 2011 1953
rect 2047 1949 2051 1953
rect 2495 1952 2499 1956
rect 2591 1952 2595 1956
rect 2695 1952 2699 1956
rect 2807 1952 2811 1956
rect 2927 1952 2931 1956
rect 3047 1952 3051 1956
rect 3175 1952 3179 1956
rect 3295 1952 3299 1956
rect 3415 1952 3419 1956
rect 3543 1952 3547 1956
rect 3671 1952 3675 1956
rect 3799 1952 3803 1956
rect 3943 1949 3947 1953
rect 111 1932 115 1936
rect 511 1933 515 1937
rect 623 1933 627 1937
rect 743 1933 747 1937
rect 871 1933 875 1937
rect 1007 1933 1011 1937
rect 1143 1933 1147 1937
rect 1279 1933 1283 1937
rect 1415 1933 1419 1937
rect 1559 1933 1563 1937
rect 1703 1933 1707 1937
rect 2007 1932 2011 1936
rect 2047 1932 2051 1936
rect 2495 1933 2499 1937
rect 2591 1933 2595 1937
rect 2695 1933 2699 1937
rect 2807 1933 2811 1937
rect 2927 1933 2931 1937
rect 3047 1933 3051 1937
rect 3175 1933 3179 1937
rect 3295 1933 3299 1937
rect 3415 1933 3419 1937
rect 3543 1933 3547 1937
rect 3671 1933 3675 1937
rect 3799 1933 3803 1937
rect 3943 1932 3947 1936
rect 111 1872 115 1876
rect 551 1871 555 1875
rect 663 1871 667 1875
rect 783 1871 787 1875
rect 911 1871 915 1875
rect 1047 1871 1051 1875
rect 1175 1871 1179 1875
rect 1311 1871 1315 1875
rect 1447 1871 1451 1875
rect 1583 1871 1587 1875
rect 1719 1871 1723 1875
rect 2007 1872 2011 1876
rect 2047 1876 2051 1880
rect 2071 1875 2075 1879
rect 2247 1875 2251 1879
rect 2439 1875 2443 1879
rect 2623 1875 2627 1879
rect 2791 1875 2795 1879
rect 2959 1875 2963 1879
rect 3127 1875 3131 1879
rect 3303 1875 3307 1879
rect 3487 1875 3491 1879
rect 3671 1875 3675 1879
rect 3839 1875 3843 1879
rect 3943 1876 3947 1880
rect 111 1855 115 1859
rect 551 1852 555 1856
rect 663 1852 667 1856
rect 783 1852 787 1856
rect 911 1852 915 1856
rect 1047 1852 1051 1856
rect 1175 1852 1179 1856
rect 1311 1852 1315 1856
rect 1447 1852 1451 1856
rect 1583 1852 1587 1856
rect 1719 1852 1723 1856
rect 2007 1855 2011 1859
rect 2047 1859 2051 1863
rect 2071 1856 2075 1860
rect 2247 1856 2251 1860
rect 2439 1856 2443 1860
rect 2623 1856 2627 1860
rect 2791 1856 2795 1860
rect 2959 1856 2963 1860
rect 3127 1856 3131 1860
rect 3303 1856 3307 1860
rect 3487 1856 3491 1860
rect 3671 1856 3675 1860
rect 3839 1856 3843 1860
rect 3943 1859 3947 1863
rect 111 1789 115 1793
rect 503 1792 507 1796
rect 615 1792 619 1796
rect 735 1792 739 1796
rect 863 1792 867 1796
rect 999 1792 1003 1796
rect 1151 1792 1155 1796
rect 1319 1792 1323 1796
rect 1487 1792 1491 1796
rect 1663 1792 1667 1796
rect 1847 1792 1851 1796
rect 2007 1789 2011 1793
rect 2047 1793 2051 1797
rect 2095 1796 2099 1800
rect 2231 1796 2235 1800
rect 2367 1796 2371 1800
rect 2511 1796 2515 1800
rect 2671 1796 2675 1800
rect 2855 1796 2859 1800
rect 3071 1796 3075 1800
rect 3303 1796 3307 1800
rect 3543 1796 3547 1800
rect 3791 1796 3795 1800
rect 3943 1793 3947 1797
rect 111 1772 115 1776
rect 503 1773 507 1777
rect 615 1773 619 1777
rect 735 1773 739 1777
rect 863 1773 867 1777
rect 999 1773 1003 1777
rect 1151 1773 1155 1777
rect 1319 1773 1323 1777
rect 1487 1773 1491 1777
rect 1663 1773 1667 1777
rect 1847 1773 1851 1777
rect 2007 1772 2011 1776
rect 2047 1776 2051 1780
rect 2095 1777 2099 1781
rect 2231 1777 2235 1781
rect 2367 1777 2371 1781
rect 2511 1777 2515 1781
rect 2671 1777 2675 1781
rect 2855 1777 2859 1781
rect 3071 1777 3075 1781
rect 3303 1777 3307 1781
rect 3543 1777 3547 1781
rect 3791 1777 3795 1781
rect 3943 1776 3947 1780
rect 111 1720 115 1724
rect 343 1719 347 1723
rect 463 1719 467 1723
rect 591 1719 595 1723
rect 719 1719 723 1723
rect 847 1719 851 1723
rect 983 1719 987 1723
rect 1127 1719 1131 1723
rect 1279 1719 1283 1723
rect 1439 1719 1443 1723
rect 1599 1719 1603 1723
rect 2007 1720 2011 1724
rect 2047 1724 2051 1728
rect 2183 1723 2187 1727
rect 2287 1723 2291 1727
rect 2391 1723 2395 1727
rect 2495 1723 2499 1727
rect 2599 1723 2603 1727
rect 2703 1723 2707 1727
rect 2807 1723 2811 1727
rect 2911 1723 2915 1727
rect 3015 1723 3019 1727
rect 3127 1723 3131 1727
rect 3943 1724 3947 1728
rect 111 1703 115 1707
rect 343 1700 347 1704
rect 463 1700 467 1704
rect 591 1700 595 1704
rect 719 1700 723 1704
rect 847 1700 851 1704
rect 983 1700 987 1704
rect 1127 1700 1131 1704
rect 1279 1700 1283 1704
rect 1439 1700 1443 1704
rect 1599 1700 1603 1704
rect 2007 1703 2011 1707
rect 2047 1707 2051 1711
rect 2183 1704 2187 1708
rect 2287 1704 2291 1708
rect 2391 1704 2395 1708
rect 2495 1704 2499 1708
rect 2599 1704 2603 1708
rect 2703 1704 2707 1708
rect 2807 1704 2811 1708
rect 2911 1704 2915 1708
rect 3015 1704 3019 1708
rect 3127 1704 3131 1708
rect 3943 1707 3947 1711
rect 2047 1641 2051 1645
rect 2231 1644 2235 1648
rect 2367 1644 2371 1648
rect 2519 1644 2523 1648
rect 2679 1644 2683 1648
rect 2847 1644 2851 1648
rect 3023 1644 3027 1648
rect 3191 1644 3195 1648
rect 3359 1644 3363 1648
rect 3527 1644 3531 1648
rect 3695 1644 3699 1648
rect 3839 1644 3843 1648
rect 111 1633 115 1637
rect 159 1636 163 1640
rect 295 1636 299 1640
rect 455 1636 459 1640
rect 623 1636 627 1640
rect 799 1636 803 1640
rect 983 1636 987 1640
rect 1167 1636 1171 1640
rect 1351 1636 1355 1640
rect 1543 1636 1547 1640
rect 3943 1641 3947 1645
rect 1735 1636 1739 1640
rect 2007 1633 2011 1637
rect 2047 1624 2051 1628
rect 2231 1625 2235 1629
rect 2367 1625 2371 1629
rect 2519 1625 2523 1629
rect 2679 1625 2683 1629
rect 2847 1625 2851 1629
rect 3023 1625 3027 1629
rect 3191 1625 3195 1629
rect 3359 1625 3363 1629
rect 3527 1625 3531 1629
rect 3695 1625 3699 1629
rect 3839 1625 3843 1629
rect 3943 1624 3947 1628
rect 111 1616 115 1620
rect 159 1617 163 1621
rect 295 1617 299 1621
rect 455 1617 459 1621
rect 623 1617 627 1621
rect 799 1617 803 1621
rect 983 1617 987 1621
rect 1167 1617 1171 1621
rect 1351 1617 1355 1621
rect 1543 1617 1547 1621
rect 1735 1617 1739 1621
rect 2007 1616 2011 1620
rect 111 1564 115 1568
rect 135 1563 139 1567
rect 255 1563 259 1567
rect 423 1563 427 1567
rect 607 1563 611 1567
rect 799 1563 803 1567
rect 991 1563 995 1567
rect 1183 1563 1187 1567
rect 1367 1563 1371 1567
rect 1551 1563 1555 1567
rect 1735 1563 1739 1567
rect 1903 1563 1907 1567
rect 2007 1564 2011 1568
rect 2047 1564 2051 1568
rect 2071 1563 2075 1567
rect 2271 1563 2275 1567
rect 2495 1563 2499 1567
rect 2711 1563 2715 1567
rect 2911 1563 2915 1567
rect 3095 1563 3099 1567
rect 3263 1563 3267 1567
rect 3423 1563 3427 1567
rect 3567 1563 3571 1567
rect 3711 1563 3715 1567
rect 3839 1563 3843 1567
rect 3943 1564 3947 1568
rect 111 1547 115 1551
rect 135 1544 139 1548
rect 255 1544 259 1548
rect 423 1544 427 1548
rect 607 1544 611 1548
rect 799 1544 803 1548
rect 991 1544 995 1548
rect 1183 1544 1187 1548
rect 1367 1544 1371 1548
rect 1551 1544 1555 1548
rect 1735 1544 1739 1548
rect 1903 1544 1907 1548
rect 2007 1547 2011 1551
rect 2047 1547 2051 1551
rect 2071 1544 2075 1548
rect 2271 1544 2275 1548
rect 2495 1544 2499 1548
rect 2711 1544 2715 1548
rect 2911 1544 2915 1548
rect 3095 1544 3099 1548
rect 3263 1544 3267 1548
rect 3423 1544 3427 1548
rect 3567 1544 3571 1548
rect 3711 1544 3715 1548
rect 3839 1544 3843 1548
rect 3943 1547 3947 1551
rect 111 1477 115 1481
rect 135 1480 139 1484
rect 247 1480 251 1484
rect 399 1480 403 1484
rect 559 1480 563 1484
rect 719 1480 723 1484
rect 879 1480 883 1484
rect 1039 1480 1043 1484
rect 1183 1480 1187 1484
rect 1319 1480 1323 1484
rect 1447 1480 1451 1484
rect 1567 1480 1571 1484
rect 1687 1480 1691 1484
rect 1807 1480 1811 1484
rect 1903 1480 1907 1484
rect 2007 1477 2011 1481
rect 2047 1481 2051 1485
rect 2071 1484 2075 1488
rect 2431 1484 2435 1488
rect 2791 1484 2795 1488
rect 3127 1484 3131 1488
rect 3463 1484 3467 1488
rect 3799 1484 3803 1488
rect 3943 1481 3947 1485
rect 111 1460 115 1464
rect 135 1461 139 1465
rect 247 1461 251 1465
rect 399 1461 403 1465
rect 559 1461 563 1465
rect 719 1461 723 1465
rect 879 1461 883 1465
rect 1039 1461 1043 1465
rect 1183 1461 1187 1465
rect 1319 1461 1323 1465
rect 1447 1461 1451 1465
rect 1567 1461 1571 1465
rect 1687 1461 1691 1465
rect 1807 1461 1811 1465
rect 1903 1461 1907 1465
rect 2007 1460 2011 1464
rect 2047 1464 2051 1468
rect 2071 1465 2075 1469
rect 2431 1465 2435 1469
rect 2791 1465 2795 1469
rect 3127 1465 3131 1469
rect 3463 1465 3467 1469
rect 3799 1465 3803 1469
rect 3943 1464 3947 1468
rect 111 1408 115 1412
rect 135 1407 139 1411
rect 263 1407 267 1411
rect 431 1407 435 1411
rect 607 1407 611 1411
rect 791 1407 795 1411
rect 975 1407 979 1411
rect 1159 1407 1163 1411
rect 1351 1407 1355 1411
rect 1543 1407 1547 1411
rect 1735 1407 1739 1411
rect 1903 1407 1907 1411
rect 2007 1408 2011 1412
rect 2047 1404 2051 1408
rect 2071 1403 2075 1407
rect 2271 1403 2275 1407
rect 2495 1403 2499 1407
rect 2711 1403 2715 1407
rect 2911 1403 2915 1407
rect 3095 1403 3099 1407
rect 3271 1403 3275 1407
rect 3439 1403 3443 1407
rect 3607 1403 3611 1407
rect 3783 1403 3787 1407
rect 3943 1404 3947 1408
rect 111 1391 115 1395
rect 135 1388 139 1392
rect 263 1388 267 1392
rect 431 1388 435 1392
rect 607 1388 611 1392
rect 791 1388 795 1392
rect 975 1388 979 1392
rect 1159 1388 1163 1392
rect 1351 1388 1355 1392
rect 1543 1388 1547 1392
rect 1735 1388 1739 1392
rect 1903 1388 1907 1392
rect 2007 1391 2011 1395
rect 2047 1387 2051 1391
rect 2071 1384 2075 1388
rect 2271 1384 2275 1388
rect 2495 1384 2499 1388
rect 2711 1384 2715 1388
rect 2911 1384 2915 1388
rect 3095 1384 3099 1388
rect 3271 1384 3275 1388
rect 3439 1384 3443 1388
rect 3607 1384 3611 1388
rect 3783 1384 3787 1388
rect 3943 1387 3947 1391
rect 111 1321 115 1325
rect 159 1324 163 1328
rect 311 1324 315 1328
rect 479 1324 483 1328
rect 663 1324 667 1328
rect 855 1324 859 1328
rect 1047 1324 1051 1328
rect 1247 1324 1251 1328
rect 1447 1324 1451 1328
rect 1655 1324 1659 1328
rect 1863 1324 1867 1328
rect 2007 1321 2011 1325
rect 2047 1321 2051 1325
rect 2071 1324 2075 1328
rect 2207 1324 2211 1328
rect 2383 1324 2387 1328
rect 2567 1324 2571 1328
rect 2751 1324 2755 1328
rect 2935 1324 2939 1328
rect 3111 1324 3115 1328
rect 3279 1324 3283 1328
rect 3447 1324 3451 1328
rect 3623 1324 3627 1328
rect 3943 1321 3947 1325
rect 111 1304 115 1308
rect 159 1305 163 1309
rect 311 1305 315 1309
rect 479 1305 483 1309
rect 663 1305 667 1309
rect 855 1305 859 1309
rect 1047 1305 1051 1309
rect 1247 1305 1251 1309
rect 1447 1305 1451 1309
rect 1655 1305 1659 1309
rect 1863 1305 1867 1309
rect 2007 1304 2011 1308
rect 2047 1304 2051 1308
rect 2071 1305 2075 1309
rect 2207 1305 2211 1309
rect 2383 1305 2387 1309
rect 2567 1305 2571 1309
rect 2751 1305 2755 1309
rect 2935 1305 2939 1309
rect 3111 1305 3115 1309
rect 3279 1305 3283 1309
rect 3447 1305 3451 1309
rect 3623 1305 3627 1309
rect 3943 1304 3947 1308
rect 111 1248 115 1252
rect 407 1247 411 1251
rect 543 1247 547 1251
rect 695 1247 699 1251
rect 855 1247 859 1251
rect 1023 1247 1027 1251
rect 1191 1247 1195 1251
rect 1367 1247 1371 1251
rect 1543 1247 1547 1251
rect 1719 1247 1723 1251
rect 1895 1247 1899 1251
rect 2007 1248 2011 1252
rect 2047 1252 2051 1256
rect 2151 1251 2155 1255
rect 2287 1251 2291 1255
rect 2431 1251 2435 1255
rect 2583 1251 2587 1255
rect 2743 1251 2747 1255
rect 2903 1251 2907 1255
rect 3071 1251 3075 1255
rect 3247 1251 3251 1255
rect 3431 1251 3435 1255
rect 3615 1251 3619 1255
rect 3807 1251 3811 1255
rect 3943 1252 3947 1256
rect 111 1231 115 1235
rect 407 1228 411 1232
rect 543 1228 547 1232
rect 695 1228 699 1232
rect 855 1228 859 1232
rect 1023 1228 1027 1232
rect 1191 1228 1195 1232
rect 1367 1228 1371 1232
rect 1543 1228 1547 1232
rect 1719 1228 1723 1232
rect 1895 1228 1899 1232
rect 2007 1231 2011 1235
rect 2047 1235 2051 1239
rect 2151 1232 2155 1236
rect 2287 1232 2291 1236
rect 2431 1232 2435 1236
rect 2583 1232 2587 1236
rect 2743 1232 2747 1236
rect 2903 1232 2907 1236
rect 3071 1232 3075 1236
rect 3247 1232 3251 1236
rect 3431 1232 3435 1236
rect 3615 1232 3619 1236
rect 3807 1232 3811 1236
rect 3943 1235 3947 1239
rect 111 1165 115 1169
rect 423 1168 427 1172
rect 591 1168 595 1172
rect 759 1168 763 1172
rect 927 1168 931 1172
rect 1095 1168 1099 1172
rect 1247 1168 1251 1172
rect 1399 1168 1403 1172
rect 1543 1168 1547 1172
rect 1687 1168 1691 1172
rect 1839 1168 1843 1172
rect 2007 1165 2011 1169
rect 2047 1169 2051 1173
rect 2311 1172 2315 1176
rect 2415 1172 2419 1176
rect 2527 1172 2531 1176
rect 2639 1172 2643 1176
rect 2767 1172 2771 1176
rect 2911 1172 2915 1176
rect 3071 1172 3075 1176
rect 3247 1172 3251 1176
rect 3439 1172 3443 1176
rect 3631 1172 3635 1176
rect 3831 1172 3835 1176
rect 3943 1169 3947 1173
rect 111 1148 115 1152
rect 423 1149 427 1153
rect 591 1149 595 1153
rect 759 1149 763 1153
rect 927 1149 931 1153
rect 1095 1149 1099 1153
rect 1247 1149 1251 1153
rect 1399 1149 1403 1153
rect 1543 1149 1547 1153
rect 1687 1149 1691 1153
rect 1839 1149 1843 1153
rect 2007 1148 2011 1152
rect 2047 1152 2051 1156
rect 2311 1153 2315 1157
rect 2415 1153 2419 1157
rect 2527 1153 2531 1157
rect 2639 1153 2643 1157
rect 2767 1153 2771 1157
rect 2911 1153 2915 1157
rect 3071 1153 3075 1157
rect 3247 1153 3251 1157
rect 3439 1153 3443 1157
rect 3631 1153 3635 1157
rect 3831 1153 3835 1157
rect 3943 1152 3947 1156
rect 111 1092 115 1096
rect 375 1091 379 1095
rect 487 1091 491 1095
rect 599 1091 603 1095
rect 711 1091 715 1095
rect 831 1091 835 1095
rect 967 1091 971 1095
rect 1119 1091 1123 1095
rect 1279 1091 1283 1095
rect 1447 1091 1451 1095
rect 1623 1091 1627 1095
rect 2007 1092 2011 1096
rect 2047 1096 2051 1100
rect 2407 1095 2411 1099
rect 2503 1095 2507 1099
rect 2599 1095 2603 1099
rect 2695 1095 2699 1099
rect 2807 1095 2811 1099
rect 2943 1095 2947 1099
rect 3095 1095 3099 1099
rect 3263 1095 3267 1099
rect 3447 1095 3451 1099
rect 3639 1095 3643 1099
rect 3839 1095 3843 1099
rect 3943 1096 3947 1100
rect 111 1075 115 1079
rect 375 1072 379 1076
rect 487 1072 491 1076
rect 599 1072 603 1076
rect 711 1072 715 1076
rect 831 1072 835 1076
rect 967 1072 971 1076
rect 1119 1072 1123 1076
rect 1279 1072 1283 1076
rect 1447 1072 1451 1076
rect 1623 1072 1627 1076
rect 2007 1075 2011 1079
rect 2047 1079 2051 1083
rect 2407 1076 2411 1080
rect 2503 1076 2507 1080
rect 2599 1076 2603 1080
rect 2695 1076 2699 1080
rect 2807 1076 2811 1080
rect 2943 1076 2947 1080
rect 3095 1076 3099 1080
rect 3263 1076 3267 1080
rect 3447 1076 3451 1080
rect 3639 1076 3643 1080
rect 3839 1076 3843 1080
rect 3943 1079 3947 1083
rect 111 1009 115 1013
rect 303 1012 307 1016
rect 447 1012 451 1016
rect 591 1012 595 1016
rect 727 1012 731 1016
rect 855 1012 859 1016
rect 975 1012 979 1016
rect 1087 1012 1091 1016
rect 1199 1012 1203 1016
rect 1311 1012 1315 1016
rect 1431 1012 1435 1016
rect 2007 1009 2011 1013
rect 2047 1009 2051 1013
rect 2455 1012 2459 1016
rect 2551 1012 2555 1016
rect 2647 1012 2651 1016
rect 2759 1012 2763 1016
rect 2887 1012 2891 1016
rect 3031 1012 3035 1016
rect 3183 1012 3187 1016
rect 3343 1012 3347 1016
rect 3503 1012 3507 1016
rect 3671 1012 3675 1016
rect 3839 1012 3843 1016
rect 3943 1009 3947 1013
rect 111 992 115 996
rect 303 993 307 997
rect 447 993 451 997
rect 591 993 595 997
rect 727 993 731 997
rect 855 993 859 997
rect 975 993 979 997
rect 1087 993 1091 997
rect 1199 993 1203 997
rect 1311 993 1315 997
rect 1431 993 1435 997
rect 2007 992 2011 996
rect 2047 992 2051 996
rect 2455 993 2459 997
rect 2551 993 2555 997
rect 2647 993 2651 997
rect 2759 993 2763 997
rect 2887 993 2891 997
rect 3031 993 3035 997
rect 3183 993 3187 997
rect 3343 993 3347 997
rect 3503 993 3507 997
rect 3671 993 3675 997
rect 3839 993 3843 997
rect 3943 992 3947 996
rect 111 940 115 944
rect 255 939 259 943
rect 447 939 451 943
rect 631 939 635 943
rect 807 939 811 943
rect 975 939 979 943
rect 1127 939 1131 943
rect 1271 939 1275 943
rect 1415 939 1419 943
rect 1551 939 1555 943
rect 1695 939 1699 943
rect 2007 940 2011 944
rect 2047 936 2051 940
rect 2423 935 2427 939
rect 2519 935 2523 939
rect 2615 935 2619 939
rect 2711 935 2715 939
rect 2823 935 2827 939
rect 2951 935 2955 939
rect 3103 935 3107 939
rect 3271 935 3275 939
rect 3455 935 3459 939
rect 3647 935 3651 939
rect 3839 935 3843 939
rect 3943 936 3947 940
rect 111 923 115 927
rect 255 920 259 924
rect 447 920 451 924
rect 631 920 635 924
rect 807 920 811 924
rect 975 920 979 924
rect 1127 920 1131 924
rect 1271 920 1275 924
rect 1415 920 1419 924
rect 1551 920 1555 924
rect 1695 920 1699 924
rect 2007 923 2011 927
rect 2047 919 2051 923
rect 2423 916 2427 920
rect 2519 916 2523 920
rect 2615 916 2619 920
rect 2711 916 2715 920
rect 2823 916 2827 920
rect 2951 916 2955 920
rect 3103 916 3107 920
rect 3271 916 3275 920
rect 3455 916 3459 920
rect 3647 916 3651 920
rect 3839 916 3843 920
rect 3943 919 3947 923
rect 111 853 115 857
rect 255 856 259 860
rect 447 856 451 860
rect 639 856 643 860
rect 823 856 827 860
rect 999 856 1003 860
rect 1167 856 1171 860
rect 1327 856 1331 860
rect 1479 856 1483 860
rect 1631 856 1635 860
rect 1783 856 1787 860
rect 2007 853 2011 857
rect 2047 853 2051 857
rect 2343 856 2347 860
rect 2439 856 2443 860
rect 2535 856 2539 860
rect 2631 856 2635 860
rect 2735 856 2739 860
rect 2863 856 2867 860
rect 3015 856 3019 860
rect 3191 856 3195 860
rect 3391 856 3395 860
rect 3607 856 3611 860
rect 3823 856 3827 860
rect 3943 853 3947 857
rect 111 836 115 840
rect 255 837 259 841
rect 447 837 451 841
rect 639 837 643 841
rect 823 837 827 841
rect 999 837 1003 841
rect 1167 837 1171 841
rect 1327 837 1331 841
rect 1479 837 1483 841
rect 1631 837 1635 841
rect 1783 837 1787 841
rect 2007 836 2011 840
rect 2047 836 2051 840
rect 2343 837 2347 841
rect 2439 837 2443 841
rect 2535 837 2539 841
rect 2631 837 2635 841
rect 2735 837 2739 841
rect 2863 837 2867 841
rect 3015 837 3019 841
rect 3191 837 3195 841
rect 3391 837 3395 841
rect 3607 837 3611 841
rect 3823 837 3827 841
rect 3943 836 3947 840
rect 111 780 115 784
rect 159 779 163 783
rect 311 779 315 783
rect 471 779 475 783
rect 623 779 627 783
rect 775 779 779 783
rect 935 779 939 783
rect 1095 779 1099 783
rect 1255 779 1259 783
rect 1415 779 1419 783
rect 1583 779 1587 783
rect 1751 779 1755 783
rect 1903 779 1907 783
rect 2007 780 2011 784
rect 2047 784 2051 788
rect 2311 783 2315 787
rect 2495 783 2499 787
rect 2687 783 2691 787
rect 2879 783 2883 787
rect 3079 783 3083 787
rect 3287 783 3291 787
rect 3503 783 3507 787
rect 3719 783 3723 787
rect 3943 784 3947 788
rect 111 763 115 767
rect 159 760 163 764
rect 311 760 315 764
rect 471 760 475 764
rect 623 760 627 764
rect 775 760 779 764
rect 935 760 939 764
rect 1095 760 1099 764
rect 1255 760 1259 764
rect 1415 760 1419 764
rect 1583 760 1587 764
rect 1751 760 1755 764
rect 1903 760 1907 764
rect 2007 763 2011 767
rect 2047 767 2051 771
rect 2311 764 2315 768
rect 2495 764 2499 768
rect 2687 764 2691 768
rect 2879 764 2883 768
rect 3079 764 3083 768
rect 3287 764 3291 768
rect 3503 764 3507 768
rect 3719 764 3723 768
rect 3943 767 3947 771
rect 111 697 115 701
rect 135 700 139 704
rect 263 700 267 704
rect 431 700 435 704
rect 623 700 627 704
rect 823 700 827 704
rect 1015 700 1019 704
rect 1207 700 1211 704
rect 1391 700 1395 704
rect 1567 700 1571 704
rect 1743 700 1747 704
rect 1903 700 1907 704
rect 2007 697 2011 701
rect 2047 697 2051 701
rect 2071 700 2075 704
rect 2255 700 2259 704
rect 2455 700 2459 704
rect 2655 700 2659 704
rect 2855 700 2859 704
rect 3047 700 3051 704
rect 3239 700 3243 704
rect 3439 700 3443 704
rect 3639 700 3643 704
rect 3839 700 3843 704
rect 3943 697 3947 701
rect 111 680 115 684
rect 135 681 139 685
rect 263 681 267 685
rect 431 681 435 685
rect 623 681 627 685
rect 823 681 827 685
rect 1015 681 1019 685
rect 1207 681 1211 685
rect 1391 681 1395 685
rect 1567 681 1571 685
rect 1743 681 1747 685
rect 1903 681 1907 685
rect 2007 680 2011 684
rect 2047 680 2051 684
rect 2071 681 2075 685
rect 2255 681 2259 685
rect 2455 681 2459 685
rect 2655 681 2659 685
rect 2855 681 2859 685
rect 3047 681 3051 685
rect 3239 681 3243 685
rect 3439 681 3443 685
rect 3639 681 3643 685
rect 3839 681 3843 685
rect 3943 680 3947 684
rect 111 628 115 632
rect 135 627 139 631
rect 247 627 251 631
rect 383 627 387 631
rect 527 627 531 631
rect 687 627 691 631
rect 871 627 875 631
rect 1079 627 1083 631
rect 1303 627 1307 631
rect 1543 627 1547 631
rect 1783 627 1787 631
rect 2007 628 2011 632
rect 2047 628 2051 632
rect 2071 627 2075 631
rect 2231 627 2235 631
rect 2431 627 2435 631
rect 2631 627 2635 631
rect 2831 627 2835 631
rect 3023 627 3027 631
rect 3207 627 3211 631
rect 3375 627 3379 631
rect 3535 627 3539 631
rect 3695 627 3699 631
rect 3839 627 3843 631
rect 3943 628 3947 632
rect 111 611 115 615
rect 135 608 139 612
rect 247 608 251 612
rect 383 608 387 612
rect 527 608 531 612
rect 687 608 691 612
rect 871 608 875 612
rect 1079 608 1083 612
rect 1303 608 1307 612
rect 1543 608 1547 612
rect 1783 608 1787 612
rect 2007 611 2011 615
rect 2047 611 2051 615
rect 2071 608 2075 612
rect 2231 608 2235 612
rect 2431 608 2435 612
rect 2631 608 2635 612
rect 2831 608 2835 612
rect 3023 608 3027 612
rect 3207 608 3211 612
rect 3375 608 3379 612
rect 3535 608 3539 612
rect 3695 608 3699 612
rect 3839 608 3843 612
rect 3943 611 3947 615
rect 111 541 115 545
rect 135 544 139 548
rect 295 544 299 548
rect 479 544 483 548
rect 663 544 667 548
rect 847 544 851 548
rect 1031 544 1035 548
rect 1215 544 1219 548
rect 1399 544 1403 548
rect 1591 544 1595 548
rect 1783 544 1787 548
rect 2007 541 2011 545
rect 2047 541 2051 545
rect 2071 544 2075 548
rect 2215 544 2219 548
rect 2399 544 2403 548
rect 2583 544 2587 548
rect 2775 544 2779 548
rect 2959 544 2963 548
rect 3143 544 3147 548
rect 3319 544 3323 548
rect 3495 544 3499 548
rect 3679 544 3683 548
rect 3839 544 3843 548
rect 3943 541 3947 545
rect 111 524 115 528
rect 135 525 139 529
rect 295 525 299 529
rect 479 525 483 529
rect 663 525 667 529
rect 847 525 851 529
rect 1031 525 1035 529
rect 1215 525 1219 529
rect 1399 525 1403 529
rect 1591 525 1595 529
rect 1783 525 1787 529
rect 2007 524 2011 528
rect 2047 524 2051 528
rect 2071 525 2075 529
rect 2215 525 2219 529
rect 2399 525 2403 529
rect 2583 525 2587 529
rect 2775 525 2779 529
rect 2959 525 2963 529
rect 3143 525 3147 529
rect 3319 525 3323 529
rect 3495 525 3499 529
rect 3679 525 3683 529
rect 3839 525 3843 529
rect 3943 524 3947 528
rect 111 472 115 476
rect 135 471 139 475
rect 287 471 291 475
rect 455 471 459 475
rect 615 471 619 475
rect 767 471 771 475
rect 903 471 907 475
rect 1031 471 1035 475
rect 1159 471 1163 475
rect 1287 471 1291 475
rect 1415 471 1419 475
rect 2007 472 2011 476
rect 2047 468 2051 472
rect 2071 467 2075 471
rect 2223 467 2227 471
rect 2391 467 2395 471
rect 2559 467 2563 471
rect 2727 467 2731 471
rect 2895 467 2899 471
rect 3063 467 3067 471
rect 3223 467 3227 471
rect 3383 467 3387 471
rect 3543 467 3547 471
rect 3703 467 3707 471
rect 3839 467 3843 471
rect 3943 468 3947 472
rect 111 455 115 459
rect 135 452 139 456
rect 287 452 291 456
rect 455 452 459 456
rect 615 452 619 456
rect 767 452 771 456
rect 903 452 907 456
rect 1031 452 1035 456
rect 1159 452 1163 456
rect 1287 452 1291 456
rect 1415 452 1419 456
rect 2007 455 2011 459
rect 2047 451 2051 455
rect 2071 448 2075 452
rect 2223 448 2227 452
rect 2391 448 2395 452
rect 2559 448 2563 452
rect 2727 448 2731 452
rect 2895 448 2899 452
rect 3063 448 3067 452
rect 3223 448 3227 452
rect 3383 448 3387 452
rect 3543 448 3547 452
rect 3703 448 3707 452
rect 3839 448 3843 452
rect 3943 451 3947 455
rect 111 389 115 393
rect 135 392 139 396
rect 287 392 291 396
rect 447 392 451 396
rect 599 392 603 396
rect 751 392 755 396
rect 903 392 907 396
rect 1079 392 1083 396
rect 1271 392 1275 396
rect 1479 392 1483 396
rect 1703 392 1707 396
rect 1903 392 1907 396
rect 2007 389 2011 393
rect 2047 385 2051 389
rect 2463 388 2467 392
rect 2559 388 2563 392
rect 2655 388 2659 392
rect 2751 388 2755 392
rect 2847 388 2851 392
rect 2943 388 2947 392
rect 3039 388 3043 392
rect 3135 388 3139 392
rect 3231 388 3235 392
rect 3943 385 3947 389
rect 111 372 115 376
rect 135 373 139 377
rect 287 373 291 377
rect 447 373 451 377
rect 599 373 603 377
rect 751 373 755 377
rect 903 373 907 377
rect 1079 373 1083 377
rect 1271 373 1275 377
rect 1479 373 1483 377
rect 1703 373 1707 377
rect 1903 373 1907 377
rect 2007 372 2011 376
rect 2047 368 2051 372
rect 2463 369 2467 373
rect 2559 369 2563 373
rect 2655 369 2659 373
rect 2751 369 2755 373
rect 2847 369 2851 373
rect 2943 369 2947 373
rect 3039 369 3043 373
rect 3135 369 3139 373
rect 3231 369 3235 373
rect 3943 368 3947 372
rect 111 316 115 320
rect 159 315 163 319
rect 351 315 355 319
rect 551 315 555 319
rect 759 315 763 319
rect 959 315 963 319
rect 1159 315 1163 319
rect 1343 315 1347 319
rect 1527 315 1531 319
rect 1711 315 1715 319
rect 1895 315 1899 319
rect 2007 316 2011 320
rect 2047 316 2051 320
rect 2399 315 2403 319
rect 2503 315 2507 319
rect 2623 315 2627 319
rect 2759 315 2763 319
rect 2911 315 2915 319
rect 3071 315 3075 319
rect 3247 315 3251 319
rect 3423 315 3427 319
rect 3607 315 3611 319
rect 3791 315 3795 319
rect 3943 316 3947 320
rect 111 299 115 303
rect 159 296 163 300
rect 351 296 355 300
rect 551 296 555 300
rect 759 296 763 300
rect 959 296 963 300
rect 1159 296 1163 300
rect 1343 296 1347 300
rect 1527 296 1531 300
rect 1711 296 1715 300
rect 1895 296 1899 300
rect 2007 299 2011 303
rect 2047 299 2051 303
rect 2399 296 2403 300
rect 2503 296 2507 300
rect 2623 296 2627 300
rect 2759 296 2763 300
rect 2911 296 2915 300
rect 3071 296 3075 300
rect 3247 296 3251 300
rect 3423 296 3427 300
rect 3607 296 3611 300
rect 3791 296 3795 300
rect 3943 299 3947 303
rect 2047 233 2051 237
rect 2191 236 2195 240
rect 2351 236 2355 240
rect 2519 236 2523 240
rect 2687 236 2691 240
rect 2855 236 2859 240
rect 3031 236 3035 240
rect 3215 236 3219 240
rect 3407 236 3411 240
rect 3607 236 3611 240
rect 3807 236 3811 240
rect 111 225 115 229
rect 223 228 227 232
rect 383 228 387 232
rect 543 228 547 232
rect 703 228 707 232
rect 863 228 867 232
rect 1031 228 1035 232
rect 1199 228 1203 232
rect 1367 228 1371 232
rect 1543 228 1547 232
rect 1727 228 1731 232
rect 3943 233 3947 237
rect 1903 228 1907 232
rect 2007 225 2011 229
rect 2047 216 2051 220
rect 2191 217 2195 221
rect 2351 217 2355 221
rect 2519 217 2523 221
rect 2687 217 2691 221
rect 2855 217 2859 221
rect 3031 217 3035 221
rect 3215 217 3219 221
rect 3407 217 3411 221
rect 3607 217 3611 221
rect 3807 217 3811 221
rect 3943 216 3947 220
rect 111 208 115 212
rect 223 209 227 213
rect 383 209 387 213
rect 543 209 547 213
rect 703 209 707 213
rect 863 209 867 213
rect 1031 209 1035 213
rect 1199 209 1203 213
rect 1367 209 1371 213
rect 1543 209 1547 213
rect 1727 209 1731 213
rect 1903 209 1907 213
rect 2007 208 2011 212
rect 111 136 115 140
rect 135 135 139 139
rect 231 135 235 139
rect 327 135 331 139
rect 423 135 427 139
rect 527 135 531 139
rect 647 135 651 139
rect 775 135 779 139
rect 903 135 907 139
rect 1031 135 1035 139
rect 1151 135 1155 139
rect 1271 135 1275 139
rect 1383 135 1387 139
rect 1487 135 1491 139
rect 1591 135 1595 139
rect 1703 135 1707 139
rect 1807 135 1811 139
rect 1903 135 1907 139
rect 2007 136 2011 140
rect 2047 132 2051 136
rect 2071 131 2075 135
rect 2167 131 2171 135
rect 2263 131 2267 135
rect 2367 131 2371 135
rect 2487 131 2491 135
rect 2615 131 2619 135
rect 2743 131 2747 135
rect 2871 131 2875 135
rect 2991 131 2995 135
rect 3111 131 3115 135
rect 3223 131 3227 135
rect 3327 131 3331 135
rect 3431 131 3435 135
rect 3535 131 3539 135
rect 3639 131 3643 135
rect 3743 131 3747 135
rect 3839 131 3843 135
rect 3943 132 3947 136
rect 111 119 115 123
rect 135 116 139 120
rect 231 116 235 120
rect 327 116 331 120
rect 423 116 427 120
rect 527 116 531 120
rect 647 116 651 120
rect 775 116 779 120
rect 903 116 907 120
rect 1031 116 1035 120
rect 1151 116 1155 120
rect 1271 116 1275 120
rect 1383 116 1387 120
rect 1487 116 1491 120
rect 1591 116 1595 120
rect 1703 116 1707 120
rect 1807 116 1811 120
rect 1903 116 1907 120
rect 2007 119 2011 123
rect 2047 115 2051 119
rect 2071 112 2075 116
rect 2167 112 2171 116
rect 2263 112 2267 116
rect 2367 112 2371 116
rect 2487 112 2491 116
rect 2615 112 2619 116
rect 2743 112 2747 116
rect 2871 112 2875 116
rect 2991 112 2995 116
rect 3111 112 3115 116
rect 3223 112 3227 116
rect 3327 112 3331 116
rect 3431 112 3435 116
rect 3535 112 3539 116
rect 3639 112 3643 116
rect 3743 112 3747 116
rect 3839 112 3843 116
rect 3943 115 3947 119
<< m3 >>
rect 2047 4030 2051 4031
rect 2047 4025 2051 4026
rect 2071 4030 2075 4031
rect 2071 4025 2075 4026
rect 3943 4030 3947 4031
rect 3943 4025 3947 4026
rect 111 4010 115 4011
rect 111 4005 115 4006
rect 151 4010 155 4011
rect 151 4005 155 4006
rect 279 4010 283 4011
rect 279 4005 283 4006
rect 431 4010 435 4011
rect 431 4005 435 4006
rect 607 4010 611 4011
rect 607 4005 611 4006
rect 791 4010 795 4011
rect 791 4005 795 4006
rect 975 4010 979 4011
rect 975 4005 979 4006
rect 1151 4010 1155 4011
rect 1151 4005 1155 4006
rect 1311 4010 1315 4011
rect 1311 4005 1315 4006
rect 1471 4010 1475 4011
rect 1471 4005 1475 4006
rect 1623 4010 1627 4011
rect 1623 4005 1627 4006
rect 1775 4010 1779 4011
rect 1775 4005 1779 4006
rect 1903 4010 1907 4011
rect 1903 4005 1907 4006
rect 2007 4010 2011 4011
rect 2007 4005 2011 4006
rect 2048 4005 2050 4025
rect 112 3985 114 4005
rect 110 3984 116 3985
rect 152 3984 154 4005
rect 280 3984 282 4005
rect 432 3984 434 4005
rect 608 3984 610 4005
rect 792 3984 794 4005
rect 976 3984 978 4005
rect 1152 3984 1154 4005
rect 1312 3984 1314 4005
rect 1472 3984 1474 4005
rect 1624 3984 1626 4005
rect 1776 3984 1778 4005
rect 1904 3984 1906 4005
rect 2008 3985 2010 4005
rect 2046 4004 2052 4005
rect 2072 4004 2074 4025
rect 3944 4005 3946 4025
rect 3942 4004 3948 4005
rect 2046 4000 2047 4004
rect 2051 4000 2052 4004
rect 2046 3999 2052 4000
rect 2070 4003 2076 4004
rect 2070 3999 2071 4003
rect 2075 3999 2076 4003
rect 3942 4000 3943 4004
rect 3947 4000 3948 4004
rect 3942 3999 3948 4000
rect 2070 3998 2076 3999
rect 2046 3987 2052 3988
rect 2006 3984 2012 3985
rect 110 3980 111 3984
rect 115 3980 116 3984
rect 110 3979 116 3980
rect 150 3983 156 3984
rect 150 3979 151 3983
rect 155 3979 156 3983
rect 150 3978 156 3979
rect 278 3983 284 3984
rect 278 3979 279 3983
rect 283 3979 284 3983
rect 278 3978 284 3979
rect 430 3983 436 3984
rect 430 3979 431 3983
rect 435 3979 436 3983
rect 430 3978 436 3979
rect 606 3983 612 3984
rect 606 3979 607 3983
rect 611 3979 612 3983
rect 606 3978 612 3979
rect 790 3983 796 3984
rect 790 3979 791 3983
rect 795 3979 796 3983
rect 790 3978 796 3979
rect 974 3983 980 3984
rect 974 3979 975 3983
rect 979 3979 980 3983
rect 974 3978 980 3979
rect 1150 3983 1156 3984
rect 1150 3979 1151 3983
rect 1155 3979 1156 3983
rect 1150 3978 1156 3979
rect 1310 3983 1316 3984
rect 1310 3979 1311 3983
rect 1315 3979 1316 3983
rect 1310 3978 1316 3979
rect 1470 3983 1476 3984
rect 1470 3979 1471 3983
rect 1475 3979 1476 3983
rect 1470 3978 1476 3979
rect 1622 3983 1628 3984
rect 1622 3979 1623 3983
rect 1627 3979 1628 3983
rect 1622 3978 1628 3979
rect 1774 3983 1780 3984
rect 1774 3979 1775 3983
rect 1779 3979 1780 3983
rect 1774 3978 1780 3979
rect 1902 3983 1908 3984
rect 1902 3979 1903 3983
rect 1907 3979 1908 3983
rect 2006 3980 2007 3984
rect 2011 3980 2012 3984
rect 2046 3983 2047 3987
rect 2051 3983 2052 3987
rect 3942 3987 3948 3988
rect 2046 3982 2052 3983
rect 2070 3984 2076 3985
rect 2006 3979 2012 3980
rect 1902 3978 1908 3979
rect 110 3967 116 3968
rect 110 3963 111 3967
rect 115 3963 116 3967
rect 2006 3967 2012 3968
rect 110 3962 116 3963
rect 150 3964 156 3965
rect 112 3935 114 3962
rect 150 3960 151 3964
rect 155 3960 156 3964
rect 150 3959 156 3960
rect 278 3964 284 3965
rect 278 3960 279 3964
rect 283 3960 284 3964
rect 278 3959 284 3960
rect 430 3964 436 3965
rect 430 3960 431 3964
rect 435 3960 436 3964
rect 430 3959 436 3960
rect 606 3964 612 3965
rect 606 3960 607 3964
rect 611 3960 612 3964
rect 606 3959 612 3960
rect 790 3964 796 3965
rect 790 3960 791 3964
rect 795 3960 796 3964
rect 790 3959 796 3960
rect 974 3964 980 3965
rect 974 3960 975 3964
rect 979 3960 980 3964
rect 974 3959 980 3960
rect 1150 3964 1156 3965
rect 1150 3960 1151 3964
rect 1155 3960 1156 3964
rect 1150 3959 1156 3960
rect 1310 3964 1316 3965
rect 1310 3960 1311 3964
rect 1315 3960 1316 3964
rect 1310 3959 1316 3960
rect 1470 3964 1476 3965
rect 1470 3960 1471 3964
rect 1475 3960 1476 3964
rect 1470 3959 1476 3960
rect 1622 3964 1628 3965
rect 1622 3960 1623 3964
rect 1627 3960 1628 3964
rect 1622 3959 1628 3960
rect 1774 3964 1780 3965
rect 1774 3960 1775 3964
rect 1779 3960 1780 3964
rect 1774 3959 1780 3960
rect 1902 3964 1908 3965
rect 1902 3960 1903 3964
rect 1907 3960 1908 3964
rect 2006 3963 2007 3967
rect 2011 3963 2012 3967
rect 2006 3962 2012 3963
rect 1902 3959 1908 3960
rect 152 3935 154 3959
rect 280 3935 282 3959
rect 432 3935 434 3959
rect 608 3935 610 3959
rect 792 3935 794 3959
rect 976 3935 978 3959
rect 1152 3935 1154 3959
rect 1312 3935 1314 3959
rect 1472 3935 1474 3959
rect 1624 3935 1626 3959
rect 1776 3935 1778 3959
rect 1904 3935 1906 3959
rect 2008 3935 2010 3962
rect 2048 3955 2050 3982
rect 2070 3980 2071 3984
rect 2075 3980 2076 3984
rect 3942 3983 3943 3987
rect 3947 3983 3948 3987
rect 3942 3982 3948 3983
rect 2070 3979 2076 3980
rect 2072 3955 2074 3979
rect 3944 3955 3946 3982
rect 2047 3954 2051 3955
rect 2047 3949 2051 3950
rect 2071 3954 2075 3955
rect 2071 3949 2075 3950
rect 2079 3954 2083 3955
rect 2079 3949 2083 3950
rect 2215 3954 2219 3955
rect 2215 3949 2219 3950
rect 2359 3954 2363 3955
rect 2359 3949 2363 3950
rect 2503 3954 2507 3955
rect 2503 3949 2507 3950
rect 2647 3954 2651 3955
rect 2647 3949 2651 3950
rect 2791 3954 2795 3955
rect 2791 3949 2795 3950
rect 2927 3954 2931 3955
rect 2927 3949 2931 3950
rect 3055 3954 3059 3955
rect 3055 3949 3059 3950
rect 3175 3954 3179 3955
rect 3175 3949 3179 3950
rect 3295 3954 3299 3955
rect 3295 3949 3299 3950
rect 3415 3954 3419 3955
rect 3415 3949 3419 3950
rect 3535 3954 3539 3955
rect 3535 3949 3539 3950
rect 3943 3954 3947 3955
rect 3943 3949 3947 3950
rect 111 3934 115 3935
rect 111 3929 115 3930
rect 151 3934 155 3935
rect 151 3929 155 3930
rect 279 3934 283 3935
rect 279 3929 283 3930
rect 303 3934 307 3935
rect 303 3929 307 3930
rect 423 3934 427 3935
rect 423 3929 427 3930
rect 431 3934 435 3935
rect 431 3929 435 3930
rect 551 3934 555 3935
rect 551 3929 555 3930
rect 607 3934 611 3935
rect 607 3929 611 3930
rect 687 3934 691 3935
rect 687 3929 691 3930
rect 791 3934 795 3935
rect 791 3929 795 3930
rect 815 3934 819 3935
rect 815 3929 819 3930
rect 943 3934 947 3935
rect 943 3929 947 3930
rect 975 3934 979 3935
rect 975 3929 979 3930
rect 1071 3934 1075 3935
rect 1071 3929 1075 3930
rect 1151 3934 1155 3935
rect 1151 3929 1155 3930
rect 1199 3934 1203 3935
rect 1199 3929 1203 3930
rect 1311 3934 1315 3935
rect 1311 3929 1315 3930
rect 1327 3934 1331 3935
rect 1327 3929 1331 3930
rect 1463 3934 1467 3935
rect 1463 3929 1467 3930
rect 1471 3934 1475 3935
rect 1471 3929 1475 3930
rect 1623 3934 1627 3935
rect 1623 3929 1627 3930
rect 1775 3934 1779 3935
rect 1775 3929 1779 3930
rect 1903 3934 1907 3935
rect 1903 3929 1907 3930
rect 2007 3934 2011 3935
rect 2007 3929 2011 3930
rect 112 3902 114 3929
rect 304 3905 306 3929
rect 424 3905 426 3929
rect 552 3905 554 3929
rect 688 3905 690 3929
rect 816 3905 818 3929
rect 944 3905 946 3929
rect 1072 3905 1074 3929
rect 1200 3905 1202 3929
rect 1328 3905 1330 3929
rect 1464 3905 1466 3929
rect 302 3904 308 3905
rect 110 3901 116 3902
rect 110 3897 111 3901
rect 115 3897 116 3901
rect 302 3900 303 3904
rect 307 3900 308 3904
rect 302 3899 308 3900
rect 422 3904 428 3905
rect 422 3900 423 3904
rect 427 3900 428 3904
rect 422 3899 428 3900
rect 550 3904 556 3905
rect 550 3900 551 3904
rect 555 3900 556 3904
rect 550 3899 556 3900
rect 686 3904 692 3905
rect 686 3900 687 3904
rect 691 3900 692 3904
rect 686 3899 692 3900
rect 814 3904 820 3905
rect 814 3900 815 3904
rect 819 3900 820 3904
rect 814 3899 820 3900
rect 942 3904 948 3905
rect 942 3900 943 3904
rect 947 3900 948 3904
rect 942 3899 948 3900
rect 1070 3904 1076 3905
rect 1070 3900 1071 3904
rect 1075 3900 1076 3904
rect 1070 3899 1076 3900
rect 1198 3904 1204 3905
rect 1198 3900 1199 3904
rect 1203 3900 1204 3904
rect 1198 3899 1204 3900
rect 1326 3904 1332 3905
rect 1326 3900 1327 3904
rect 1331 3900 1332 3904
rect 1326 3899 1332 3900
rect 1462 3904 1468 3905
rect 1462 3900 1463 3904
rect 1467 3900 1468 3904
rect 2008 3902 2010 3929
rect 2048 3922 2050 3949
rect 2080 3925 2082 3949
rect 2216 3925 2218 3949
rect 2360 3925 2362 3949
rect 2504 3925 2506 3949
rect 2648 3925 2650 3949
rect 2792 3925 2794 3949
rect 2928 3925 2930 3949
rect 3056 3925 3058 3949
rect 3176 3925 3178 3949
rect 3296 3925 3298 3949
rect 3416 3925 3418 3949
rect 3536 3925 3538 3949
rect 2078 3924 2084 3925
rect 2046 3921 2052 3922
rect 2046 3917 2047 3921
rect 2051 3917 2052 3921
rect 2078 3920 2079 3924
rect 2083 3920 2084 3924
rect 2078 3919 2084 3920
rect 2214 3924 2220 3925
rect 2214 3920 2215 3924
rect 2219 3920 2220 3924
rect 2214 3919 2220 3920
rect 2358 3924 2364 3925
rect 2358 3920 2359 3924
rect 2363 3920 2364 3924
rect 2358 3919 2364 3920
rect 2502 3924 2508 3925
rect 2502 3920 2503 3924
rect 2507 3920 2508 3924
rect 2502 3919 2508 3920
rect 2646 3924 2652 3925
rect 2646 3920 2647 3924
rect 2651 3920 2652 3924
rect 2646 3919 2652 3920
rect 2790 3924 2796 3925
rect 2790 3920 2791 3924
rect 2795 3920 2796 3924
rect 2790 3919 2796 3920
rect 2926 3924 2932 3925
rect 2926 3920 2927 3924
rect 2931 3920 2932 3924
rect 2926 3919 2932 3920
rect 3054 3924 3060 3925
rect 3054 3920 3055 3924
rect 3059 3920 3060 3924
rect 3054 3919 3060 3920
rect 3174 3924 3180 3925
rect 3174 3920 3175 3924
rect 3179 3920 3180 3924
rect 3174 3919 3180 3920
rect 3294 3924 3300 3925
rect 3294 3920 3295 3924
rect 3299 3920 3300 3924
rect 3294 3919 3300 3920
rect 3414 3924 3420 3925
rect 3414 3920 3415 3924
rect 3419 3920 3420 3924
rect 3414 3919 3420 3920
rect 3534 3924 3540 3925
rect 3534 3920 3535 3924
rect 3539 3920 3540 3924
rect 3944 3922 3946 3949
rect 3534 3919 3540 3920
rect 3942 3921 3948 3922
rect 2046 3916 2052 3917
rect 3942 3917 3943 3921
rect 3947 3917 3948 3921
rect 3942 3916 3948 3917
rect 2078 3905 2084 3906
rect 2046 3904 2052 3905
rect 1462 3899 1468 3900
rect 2006 3901 2012 3902
rect 110 3896 116 3897
rect 2006 3897 2007 3901
rect 2011 3897 2012 3901
rect 2046 3900 2047 3904
rect 2051 3900 2052 3904
rect 2078 3901 2079 3905
rect 2083 3901 2084 3905
rect 2078 3900 2084 3901
rect 2214 3905 2220 3906
rect 2214 3901 2215 3905
rect 2219 3901 2220 3905
rect 2214 3900 2220 3901
rect 2358 3905 2364 3906
rect 2358 3901 2359 3905
rect 2363 3901 2364 3905
rect 2358 3900 2364 3901
rect 2502 3905 2508 3906
rect 2502 3901 2503 3905
rect 2507 3901 2508 3905
rect 2502 3900 2508 3901
rect 2646 3905 2652 3906
rect 2646 3901 2647 3905
rect 2651 3901 2652 3905
rect 2646 3900 2652 3901
rect 2790 3905 2796 3906
rect 2790 3901 2791 3905
rect 2795 3901 2796 3905
rect 2790 3900 2796 3901
rect 2926 3905 2932 3906
rect 2926 3901 2927 3905
rect 2931 3901 2932 3905
rect 2926 3900 2932 3901
rect 3054 3905 3060 3906
rect 3054 3901 3055 3905
rect 3059 3901 3060 3905
rect 3054 3900 3060 3901
rect 3174 3905 3180 3906
rect 3174 3901 3175 3905
rect 3179 3901 3180 3905
rect 3174 3900 3180 3901
rect 3294 3905 3300 3906
rect 3294 3901 3295 3905
rect 3299 3901 3300 3905
rect 3294 3900 3300 3901
rect 3414 3905 3420 3906
rect 3414 3901 3415 3905
rect 3419 3901 3420 3905
rect 3414 3900 3420 3901
rect 3534 3905 3540 3906
rect 3534 3901 3535 3905
rect 3539 3901 3540 3905
rect 3534 3900 3540 3901
rect 3942 3904 3948 3905
rect 3942 3900 3943 3904
rect 3947 3900 3948 3904
rect 2046 3899 2052 3900
rect 2006 3896 2012 3897
rect 302 3885 308 3886
rect 110 3884 116 3885
rect 110 3880 111 3884
rect 115 3880 116 3884
rect 302 3881 303 3885
rect 307 3881 308 3885
rect 302 3880 308 3881
rect 422 3885 428 3886
rect 422 3881 423 3885
rect 427 3881 428 3885
rect 422 3880 428 3881
rect 550 3885 556 3886
rect 550 3881 551 3885
rect 555 3881 556 3885
rect 550 3880 556 3881
rect 686 3885 692 3886
rect 686 3881 687 3885
rect 691 3881 692 3885
rect 686 3880 692 3881
rect 814 3885 820 3886
rect 814 3881 815 3885
rect 819 3881 820 3885
rect 814 3880 820 3881
rect 942 3885 948 3886
rect 942 3881 943 3885
rect 947 3881 948 3885
rect 942 3880 948 3881
rect 1070 3885 1076 3886
rect 1070 3881 1071 3885
rect 1075 3881 1076 3885
rect 1070 3880 1076 3881
rect 1198 3885 1204 3886
rect 1198 3881 1199 3885
rect 1203 3881 1204 3885
rect 1198 3880 1204 3881
rect 1326 3885 1332 3886
rect 1326 3881 1327 3885
rect 1331 3881 1332 3885
rect 1326 3880 1332 3881
rect 1462 3885 1468 3886
rect 1462 3881 1463 3885
rect 1467 3881 1468 3885
rect 1462 3880 1468 3881
rect 2006 3884 2012 3885
rect 2006 3880 2007 3884
rect 2011 3880 2012 3884
rect 110 3879 116 3880
rect 112 3855 114 3879
rect 304 3855 306 3880
rect 424 3855 426 3880
rect 552 3855 554 3880
rect 688 3855 690 3880
rect 816 3855 818 3880
rect 944 3855 946 3880
rect 1072 3855 1074 3880
rect 1200 3855 1202 3880
rect 1328 3855 1330 3880
rect 1464 3855 1466 3880
rect 2006 3879 2012 3880
rect 2048 3879 2050 3899
rect 2080 3879 2082 3900
rect 2216 3879 2218 3900
rect 2360 3879 2362 3900
rect 2504 3879 2506 3900
rect 2648 3879 2650 3900
rect 2792 3879 2794 3900
rect 2928 3879 2930 3900
rect 3056 3879 3058 3900
rect 3176 3879 3178 3900
rect 3296 3879 3298 3900
rect 3416 3879 3418 3900
rect 3536 3879 3538 3900
rect 3942 3899 3948 3900
rect 3944 3879 3946 3899
rect 2008 3855 2010 3879
rect 2047 3878 2051 3879
rect 2047 3873 2051 3874
rect 2079 3878 2083 3879
rect 2079 3873 2083 3874
rect 2215 3878 2219 3879
rect 2215 3873 2219 3874
rect 2255 3878 2259 3879
rect 2255 3873 2259 3874
rect 2359 3878 2363 3879
rect 2359 3873 2363 3874
rect 2383 3878 2387 3879
rect 2383 3873 2387 3874
rect 2503 3878 2507 3879
rect 2503 3873 2507 3874
rect 2519 3878 2523 3879
rect 2519 3873 2523 3874
rect 2647 3878 2651 3879
rect 2647 3873 2651 3874
rect 2671 3878 2675 3879
rect 2671 3873 2675 3874
rect 2791 3878 2795 3879
rect 2791 3873 2795 3874
rect 2831 3878 2835 3879
rect 2831 3873 2835 3874
rect 2927 3878 2931 3879
rect 2927 3873 2931 3874
rect 2991 3878 2995 3879
rect 2991 3873 2995 3874
rect 3055 3878 3059 3879
rect 3055 3873 3059 3874
rect 3159 3878 3163 3879
rect 3159 3873 3163 3874
rect 3175 3878 3179 3879
rect 3175 3873 3179 3874
rect 3295 3878 3299 3879
rect 3295 3873 3299 3874
rect 3327 3878 3331 3879
rect 3327 3873 3331 3874
rect 3415 3878 3419 3879
rect 3415 3873 3419 3874
rect 3495 3878 3499 3879
rect 3495 3873 3499 3874
rect 3535 3878 3539 3879
rect 3535 3873 3539 3874
rect 3663 3878 3667 3879
rect 3663 3873 3667 3874
rect 3943 3878 3947 3879
rect 3943 3873 3947 3874
rect 111 3854 115 3855
rect 111 3849 115 3850
rect 303 3854 307 3855
rect 303 3849 307 3850
rect 415 3854 419 3855
rect 415 3849 419 3850
rect 423 3854 427 3855
rect 423 3849 427 3850
rect 551 3854 555 3855
rect 551 3849 555 3850
rect 567 3854 571 3855
rect 567 3849 571 3850
rect 687 3854 691 3855
rect 687 3849 691 3850
rect 727 3854 731 3855
rect 727 3849 731 3850
rect 815 3854 819 3855
rect 815 3849 819 3850
rect 887 3854 891 3855
rect 887 3849 891 3850
rect 943 3854 947 3855
rect 943 3849 947 3850
rect 1039 3854 1043 3855
rect 1039 3849 1043 3850
rect 1071 3854 1075 3855
rect 1071 3849 1075 3850
rect 1191 3854 1195 3855
rect 1191 3849 1195 3850
rect 1199 3854 1203 3855
rect 1199 3849 1203 3850
rect 1327 3854 1331 3855
rect 1327 3849 1331 3850
rect 1343 3854 1347 3855
rect 1343 3849 1347 3850
rect 1463 3854 1467 3855
rect 1463 3849 1467 3850
rect 1495 3854 1499 3855
rect 1495 3849 1499 3850
rect 1647 3854 1651 3855
rect 1647 3849 1651 3850
rect 2007 3854 2011 3855
rect 2048 3853 2050 3873
rect 2007 3849 2011 3850
rect 2046 3852 2052 3853
rect 2256 3852 2258 3873
rect 2384 3852 2386 3873
rect 2520 3852 2522 3873
rect 2672 3852 2674 3873
rect 2832 3852 2834 3873
rect 2992 3852 2994 3873
rect 3160 3852 3162 3873
rect 3328 3852 3330 3873
rect 3496 3852 3498 3873
rect 3664 3852 3666 3873
rect 3944 3853 3946 3873
rect 3942 3852 3948 3853
rect 112 3829 114 3849
rect 110 3828 116 3829
rect 416 3828 418 3849
rect 568 3828 570 3849
rect 728 3828 730 3849
rect 888 3828 890 3849
rect 1040 3828 1042 3849
rect 1192 3828 1194 3849
rect 1344 3828 1346 3849
rect 1496 3828 1498 3849
rect 1648 3828 1650 3849
rect 2008 3829 2010 3849
rect 2046 3848 2047 3852
rect 2051 3848 2052 3852
rect 2046 3847 2052 3848
rect 2254 3851 2260 3852
rect 2254 3847 2255 3851
rect 2259 3847 2260 3851
rect 2254 3846 2260 3847
rect 2382 3851 2388 3852
rect 2382 3847 2383 3851
rect 2387 3847 2388 3851
rect 2382 3846 2388 3847
rect 2518 3851 2524 3852
rect 2518 3847 2519 3851
rect 2523 3847 2524 3851
rect 2518 3846 2524 3847
rect 2670 3851 2676 3852
rect 2670 3847 2671 3851
rect 2675 3847 2676 3851
rect 2670 3846 2676 3847
rect 2830 3851 2836 3852
rect 2830 3847 2831 3851
rect 2835 3847 2836 3851
rect 2830 3846 2836 3847
rect 2990 3851 2996 3852
rect 2990 3847 2991 3851
rect 2995 3847 2996 3851
rect 2990 3846 2996 3847
rect 3158 3851 3164 3852
rect 3158 3847 3159 3851
rect 3163 3847 3164 3851
rect 3158 3846 3164 3847
rect 3326 3851 3332 3852
rect 3326 3847 3327 3851
rect 3331 3847 3332 3851
rect 3326 3846 3332 3847
rect 3494 3851 3500 3852
rect 3494 3847 3495 3851
rect 3499 3847 3500 3851
rect 3494 3846 3500 3847
rect 3662 3851 3668 3852
rect 3662 3847 3663 3851
rect 3667 3847 3668 3851
rect 3942 3848 3943 3852
rect 3947 3848 3948 3852
rect 3942 3847 3948 3848
rect 3662 3846 3668 3847
rect 2046 3835 2052 3836
rect 2046 3831 2047 3835
rect 2051 3831 2052 3835
rect 3942 3835 3948 3836
rect 2046 3830 2052 3831
rect 2254 3832 2260 3833
rect 2006 3828 2012 3829
rect 110 3824 111 3828
rect 115 3824 116 3828
rect 110 3823 116 3824
rect 414 3827 420 3828
rect 414 3823 415 3827
rect 419 3823 420 3827
rect 414 3822 420 3823
rect 566 3827 572 3828
rect 566 3823 567 3827
rect 571 3823 572 3827
rect 566 3822 572 3823
rect 726 3827 732 3828
rect 726 3823 727 3827
rect 731 3823 732 3827
rect 726 3822 732 3823
rect 886 3827 892 3828
rect 886 3823 887 3827
rect 891 3823 892 3827
rect 886 3822 892 3823
rect 1038 3827 1044 3828
rect 1038 3823 1039 3827
rect 1043 3823 1044 3827
rect 1038 3822 1044 3823
rect 1190 3827 1196 3828
rect 1190 3823 1191 3827
rect 1195 3823 1196 3827
rect 1190 3822 1196 3823
rect 1342 3827 1348 3828
rect 1342 3823 1343 3827
rect 1347 3823 1348 3827
rect 1342 3822 1348 3823
rect 1494 3827 1500 3828
rect 1494 3823 1495 3827
rect 1499 3823 1500 3827
rect 1494 3822 1500 3823
rect 1646 3827 1652 3828
rect 1646 3823 1647 3827
rect 1651 3823 1652 3827
rect 2006 3824 2007 3828
rect 2011 3824 2012 3828
rect 2006 3823 2012 3824
rect 1646 3822 1652 3823
rect 110 3811 116 3812
rect 110 3807 111 3811
rect 115 3807 116 3811
rect 2006 3811 2012 3812
rect 110 3806 116 3807
rect 414 3808 420 3809
rect 112 3775 114 3806
rect 414 3804 415 3808
rect 419 3804 420 3808
rect 414 3803 420 3804
rect 566 3808 572 3809
rect 566 3804 567 3808
rect 571 3804 572 3808
rect 566 3803 572 3804
rect 726 3808 732 3809
rect 726 3804 727 3808
rect 731 3804 732 3808
rect 726 3803 732 3804
rect 886 3808 892 3809
rect 886 3804 887 3808
rect 891 3804 892 3808
rect 886 3803 892 3804
rect 1038 3808 1044 3809
rect 1038 3804 1039 3808
rect 1043 3804 1044 3808
rect 1038 3803 1044 3804
rect 1190 3808 1196 3809
rect 1190 3804 1191 3808
rect 1195 3804 1196 3808
rect 1190 3803 1196 3804
rect 1342 3808 1348 3809
rect 1342 3804 1343 3808
rect 1347 3804 1348 3808
rect 1342 3803 1348 3804
rect 1494 3808 1500 3809
rect 1494 3804 1495 3808
rect 1499 3804 1500 3808
rect 1494 3803 1500 3804
rect 1646 3808 1652 3809
rect 1646 3804 1647 3808
rect 1651 3804 1652 3808
rect 2006 3807 2007 3811
rect 2011 3807 2012 3811
rect 2006 3806 2012 3807
rect 1646 3803 1652 3804
rect 416 3775 418 3803
rect 568 3775 570 3803
rect 728 3775 730 3803
rect 888 3775 890 3803
rect 1040 3775 1042 3803
rect 1192 3775 1194 3803
rect 1344 3775 1346 3803
rect 1496 3775 1498 3803
rect 1648 3775 1650 3803
rect 2008 3775 2010 3806
rect 2048 3803 2050 3830
rect 2254 3828 2255 3832
rect 2259 3828 2260 3832
rect 2254 3827 2260 3828
rect 2382 3832 2388 3833
rect 2382 3828 2383 3832
rect 2387 3828 2388 3832
rect 2382 3827 2388 3828
rect 2518 3832 2524 3833
rect 2518 3828 2519 3832
rect 2523 3828 2524 3832
rect 2518 3827 2524 3828
rect 2670 3832 2676 3833
rect 2670 3828 2671 3832
rect 2675 3828 2676 3832
rect 2670 3827 2676 3828
rect 2830 3832 2836 3833
rect 2830 3828 2831 3832
rect 2835 3828 2836 3832
rect 2830 3827 2836 3828
rect 2990 3832 2996 3833
rect 2990 3828 2991 3832
rect 2995 3828 2996 3832
rect 2990 3827 2996 3828
rect 3158 3832 3164 3833
rect 3158 3828 3159 3832
rect 3163 3828 3164 3832
rect 3158 3827 3164 3828
rect 3326 3832 3332 3833
rect 3326 3828 3327 3832
rect 3331 3828 3332 3832
rect 3326 3827 3332 3828
rect 3494 3832 3500 3833
rect 3494 3828 3495 3832
rect 3499 3828 3500 3832
rect 3494 3827 3500 3828
rect 3662 3832 3668 3833
rect 3662 3828 3663 3832
rect 3667 3828 3668 3832
rect 3942 3831 3943 3835
rect 3947 3831 3948 3835
rect 3942 3830 3948 3831
rect 3662 3827 3668 3828
rect 2256 3803 2258 3827
rect 2384 3803 2386 3827
rect 2520 3803 2522 3827
rect 2672 3803 2674 3827
rect 2832 3803 2834 3827
rect 2992 3803 2994 3827
rect 3160 3803 3162 3827
rect 3328 3803 3330 3827
rect 3496 3803 3498 3827
rect 3664 3803 3666 3827
rect 3944 3803 3946 3830
rect 2047 3802 2051 3803
rect 2047 3797 2051 3798
rect 2071 3802 2075 3803
rect 2071 3797 2075 3798
rect 2199 3802 2203 3803
rect 2199 3797 2203 3798
rect 2255 3802 2259 3803
rect 2255 3797 2259 3798
rect 2375 3802 2379 3803
rect 2375 3797 2379 3798
rect 2383 3802 2387 3803
rect 2383 3797 2387 3798
rect 2519 3802 2523 3803
rect 2519 3797 2523 3798
rect 2559 3802 2563 3803
rect 2559 3797 2563 3798
rect 2671 3802 2675 3803
rect 2671 3797 2675 3798
rect 2751 3802 2755 3803
rect 2751 3797 2755 3798
rect 2831 3802 2835 3803
rect 2831 3797 2835 3798
rect 2951 3802 2955 3803
rect 2951 3797 2955 3798
rect 2991 3802 2995 3803
rect 2991 3797 2995 3798
rect 3143 3802 3147 3803
rect 3143 3797 3147 3798
rect 3159 3802 3163 3803
rect 3159 3797 3163 3798
rect 3327 3802 3331 3803
rect 3327 3797 3331 3798
rect 3335 3802 3339 3803
rect 3335 3797 3339 3798
rect 3495 3802 3499 3803
rect 3495 3797 3499 3798
rect 3535 3802 3539 3803
rect 3535 3797 3539 3798
rect 3663 3802 3667 3803
rect 3663 3797 3667 3798
rect 3735 3802 3739 3803
rect 3735 3797 3739 3798
rect 3943 3802 3947 3803
rect 3943 3797 3947 3798
rect 111 3774 115 3775
rect 111 3769 115 3770
rect 399 3774 403 3775
rect 399 3769 403 3770
rect 415 3774 419 3775
rect 415 3769 419 3770
rect 567 3774 571 3775
rect 567 3769 571 3770
rect 727 3774 731 3775
rect 727 3769 731 3770
rect 751 3774 755 3775
rect 751 3769 755 3770
rect 887 3774 891 3775
rect 887 3769 891 3770
rect 935 3774 939 3775
rect 935 3769 939 3770
rect 1039 3774 1043 3775
rect 1039 3769 1043 3770
rect 1127 3774 1131 3775
rect 1127 3769 1131 3770
rect 1191 3774 1195 3775
rect 1191 3769 1195 3770
rect 1311 3774 1315 3775
rect 1311 3769 1315 3770
rect 1343 3774 1347 3775
rect 1343 3769 1347 3770
rect 1495 3774 1499 3775
rect 1495 3769 1499 3770
rect 1503 3774 1507 3775
rect 1503 3769 1507 3770
rect 1647 3774 1651 3775
rect 1647 3769 1651 3770
rect 1695 3774 1699 3775
rect 1695 3769 1699 3770
rect 1887 3774 1891 3775
rect 1887 3769 1891 3770
rect 2007 3774 2011 3775
rect 2048 3770 2050 3797
rect 2072 3773 2074 3797
rect 2200 3773 2202 3797
rect 2376 3773 2378 3797
rect 2560 3773 2562 3797
rect 2752 3773 2754 3797
rect 2952 3773 2954 3797
rect 3144 3773 3146 3797
rect 3336 3773 3338 3797
rect 3536 3773 3538 3797
rect 3736 3773 3738 3797
rect 2070 3772 2076 3773
rect 2007 3769 2011 3770
rect 2046 3769 2052 3770
rect 112 3742 114 3769
rect 400 3745 402 3769
rect 568 3745 570 3769
rect 752 3745 754 3769
rect 936 3745 938 3769
rect 1128 3745 1130 3769
rect 1312 3745 1314 3769
rect 1504 3745 1506 3769
rect 1696 3745 1698 3769
rect 1888 3745 1890 3769
rect 398 3744 404 3745
rect 110 3741 116 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 398 3740 399 3744
rect 403 3740 404 3744
rect 398 3739 404 3740
rect 566 3744 572 3745
rect 566 3740 567 3744
rect 571 3740 572 3744
rect 566 3739 572 3740
rect 750 3744 756 3745
rect 750 3740 751 3744
rect 755 3740 756 3744
rect 750 3739 756 3740
rect 934 3744 940 3745
rect 934 3740 935 3744
rect 939 3740 940 3744
rect 934 3739 940 3740
rect 1126 3744 1132 3745
rect 1126 3740 1127 3744
rect 1131 3740 1132 3744
rect 1126 3739 1132 3740
rect 1310 3744 1316 3745
rect 1310 3740 1311 3744
rect 1315 3740 1316 3744
rect 1310 3739 1316 3740
rect 1502 3744 1508 3745
rect 1502 3740 1503 3744
rect 1507 3740 1508 3744
rect 1502 3739 1508 3740
rect 1694 3744 1700 3745
rect 1694 3740 1695 3744
rect 1699 3740 1700 3744
rect 1694 3739 1700 3740
rect 1886 3744 1892 3745
rect 1886 3740 1887 3744
rect 1891 3740 1892 3744
rect 2008 3742 2010 3769
rect 2046 3765 2047 3769
rect 2051 3765 2052 3769
rect 2070 3768 2071 3772
rect 2075 3768 2076 3772
rect 2070 3767 2076 3768
rect 2198 3772 2204 3773
rect 2198 3768 2199 3772
rect 2203 3768 2204 3772
rect 2198 3767 2204 3768
rect 2374 3772 2380 3773
rect 2374 3768 2375 3772
rect 2379 3768 2380 3772
rect 2374 3767 2380 3768
rect 2558 3772 2564 3773
rect 2558 3768 2559 3772
rect 2563 3768 2564 3772
rect 2558 3767 2564 3768
rect 2750 3772 2756 3773
rect 2750 3768 2751 3772
rect 2755 3768 2756 3772
rect 2750 3767 2756 3768
rect 2950 3772 2956 3773
rect 2950 3768 2951 3772
rect 2955 3768 2956 3772
rect 2950 3767 2956 3768
rect 3142 3772 3148 3773
rect 3142 3768 3143 3772
rect 3147 3768 3148 3772
rect 3142 3767 3148 3768
rect 3334 3772 3340 3773
rect 3334 3768 3335 3772
rect 3339 3768 3340 3772
rect 3334 3767 3340 3768
rect 3534 3772 3540 3773
rect 3534 3768 3535 3772
rect 3539 3768 3540 3772
rect 3534 3767 3540 3768
rect 3734 3772 3740 3773
rect 3734 3768 3735 3772
rect 3739 3768 3740 3772
rect 3944 3770 3946 3797
rect 3734 3767 3740 3768
rect 3942 3769 3948 3770
rect 2046 3764 2052 3765
rect 3942 3765 3943 3769
rect 3947 3765 3948 3769
rect 3942 3764 3948 3765
rect 2070 3753 2076 3754
rect 2046 3752 2052 3753
rect 2046 3748 2047 3752
rect 2051 3748 2052 3752
rect 2070 3749 2071 3753
rect 2075 3749 2076 3753
rect 2070 3748 2076 3749
rect 2198 3753 2204 3754
rect 2198 3749 2199 3753
rect 2203 3749 2204 3753
rect 2198 3748 2204 3749
rect 2374 3753 2380 3754
rect 2374 3749 2375 3753
rect 2379 3749 2380 3753
rect 2374 3748 2380 3749
rect 2558 3753 2564 3754
rect 2558 3749 2559 3753
rect 2563 3749 2564 3753
rect 2558 3748 2564 3749
rect 2750 3753 2756 3754
rect 2750 3749 2751 3753
rect 2755 3749 2756 3753
rect 2750 3748 2756 3749
rect 2950 3753 2956 3754
rect 2950 3749 2951 3753
rect 2955 3749 2956 3753
rect 2950 3748 2956 3749
rect 3142 3753 3148 3754
rect 3142 3749 3143 3753
rect 3147 3749 3148 3753
rect 3142 3748 3148 3749
rect 3334 3753 3340 3754
rect 3334 3749 3335 3753
rect 3339 3749 3340 3753
rect 3334 3748 3340 3749
rect 3534 3753 3540 3754
rect 3534 3749 3535 3753
rect 3539 3749 3540 3753
rect 3534 3748 3540 3749
rect 3734 3753 3740 3754
rect 3734 3749 3735 3753
rect 3739 3749 3740 3753
rect 3734 3748 3740 3749
rect 3942 3752 3948 3753
rect 3942 3748 3943 3752
rect 3947 3748 3948 3752
rect 2046 3747 2052 3748
rect 1886 3739 1892 3740
rect 2006 3741 2012 3742
rect 110 3736 116 3737
rect 2006 3737 2007 3741
rect 2011 3737 2012 3741
rect 2006 3736 2012 3737
rect 398 3725 404 3726
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 398 3721 399 3725
rect 403 3721 404 3725
rect 398 3720 404 3721
rect 566 3725 572 3726
rect 566 3721 567 3725
rect 571 3721 572 3725
rect 566 3720 572 3721
rect 750 3725 756 3726
rect 750 3721 751 3725
rect 755 3721 756 3725
rect 750 3720 756 3721
rect 934 3725 940 3726
rect 934 3721 935 3725
rect 939 3721 940 3725
rect 934 3720 940 3721
rect 1126 3725 1132 3726
rect 1126 3721 1127 3725
rect 1131 3721 1132 3725
rect 1126 3720 1132 3721
rect 1310 3725 1316 3726
rect 1310 3721 1311 3725
rect 1315 3721 1316 3725
rect 1310 3720 1316 3721
rect 1502 3725 1508 3726
rect 1502 3721 1503 3725
rect 1507 3721 1508 3725
rect 1502 3720 1508 3721
rect 1694 3725 1700 3726
rect 1694 3721 1695 3725
rect 1699 3721 1700 3725
rect 1694 3720 1700 3721
rect 1886 3725 1892 3726
rect 1886 3721 1887 3725
rect 1891 3721 1892 3725
rect 1886 3720 1892 3721
rect 2006 3724 2012 3725
rect 2006 3720 2007 3724
rect 2011 3720 2012 3724
rect 110 3719 116 3720
rect 112 3687 114 3719
rect 400 3687 402 3720
rect 568 3687 570 3720
rect 752 3687 754 3720
rect 936 3687 938 3720
rect 1128 3687 1130 3720
rect 1312 3687 1314 3720
rect 1504 3687 1506 3720
rect 1696 3687 1698 3720
rect 1888 3687 1890 3720
rect 2006 3719 2012 3720
rect 2008 3687 2010 3719
rect 2048 3715 2050 3747
rect 2072 3715 2074 3748
rect 2200 3715 2202 3748
rect 2376 3715 2378 3748
rect 2560 3715 2562 3748
rect 2752 3715 2754 3748
rect 2952 3715 2954 3748
rect 3144 3715 3146 3748
rect 3336 3715 3338 3748
rect 3536 3715 3538 3748
rect 3736 3715 3738 3748
rect 3942 3747 3948 3748
rect 3944 3715 3946 3747
rect 2047 3714 2051 3715
rect 2047 3709 2051 3710
rect 2071 3714 2075 3715
rect 2071 3709 2075 3710
rect 2199 3714 2203 3715
rect 2199 3709 2203 3710
rect 2263 3714 2267 3715
rect 2263 3709 2267 3710
rect 2375 3714 2379 3715
rect 2375 3709 2379 3710
rect 2479 3714 2483 3715
rect 2479 3709 2483 3710
rect 2559 3714 2563 3715
rect 2559 3709 2563 3710
rect 2695 3714 2699 3715
rect 2695 3709 2699 3710
rect 2751 3714 2755 3715
rect 2751 3709 2755 3710
rect 2911 3714 2915 3715
rect 2911 3709 2915 3710
rect 2951 3714 2955 3715
rect 2951 3709 2955 3710
rect 3119 3714 3123 3715
rect 3119 3709 3123 3710
rect 3143 3714 3147 3715
rect 3143 3709 3147 3710
rect 3319 3714 3323 3715
rect 3319 3709 3323 3710
rect 3335 3714 3339 3715
rect 3335 3709 3339 3710
rect 3519 3714 3523 3715
rect 3519 3709 3523 3710
rect 3535 3714 3539 3715
rect 3535 3709 3539 3710
rect 3727 3714 3731 3715
rect 3727 3709 3731 3710
rect 3735 3714 3739 3715
rect 3735 3709 3739 3710
rect 3943 3714 3947 3715
rect 3943 3709 3947 3710
rect 2048 3689 2050 3709
rect 2046 3688 2052 3689
rect 2072 3688 2074 3709
rect 2264 3688 2266 3709
rect 2480 3688 2482 3709
rect 2696 3688 2698 3709
rect 2912 3688 2914 3709
rect 3120 3688 3122 3709
rect 3320 3688 3322 3709
rect 3520 3688 3522 3709
rect 3728 3688 3730 3709
rect 3944 3689 3946 3709
rect 3942 3688 3948 3689
rect 111 3686 115 3687
rect 111 3681 115 3682
rect 367 3686 371 3687
rect 367 3681 371 3682
rect 399 3686 403 3687
rect 399 3681 403 3682
rect 519 3686 523 3687
rect 519 3681 523 3682
rect 567 3686 571 3687
rect 567 3681 571 3682
rect 679 3686 683 3687
rect 679 3681 683 3682
rect 751 3686 755 3687
rect 751 3681 755 3682
rect 847 3686 851 3687
rect 847 3681 851 3682
rect 935 3686 939 3687
rect 935 3681 939 3682
rect 1015 3686 1019 3687
rect 1015 3681 1019 3682
rect 1127 3686 1131 3687
rect 1127 3681 1131 3682
rect 1175 3686 1179 3687
rect 1175 3681 1179 3682
rect 1311 3686 1315 3687
rect 1311 3681 1315 3682
rect 1327 3686 1331 3687
rect 1327 3681 1331 3682
rect 1479 3686 1483 3687
rect 1479 3681 1483 3682
rect 1503 3686 1507 3687
rect 1503 3681 1507 3682
rect 1631 3686 1635 3687
rect 1631 3681 1635 3682
rect 1695 3686 1699 3687
rect 1695 3681 1699 3682
rect 1791 3686 1795 3687
rect 1791 3681 1795 3682
rect 1887 3686 1891 3687
rect 1887 3681 1891 3682
rect 2007 3686 2011 3687
rect 2046 3684 2047 3688
rect 2051 3684 2052 3688
rect 2046 3683 2052 3684
rect 2070 3687 2076 3688
rect 2070 3683 2071 3687
rect 2075 3683 2076 3687
rect 2070 3682 2076 3683
rect 2262 3687 2268 3688
rect 2262 3683 2263 3687
rect 2267 3683 2268 3687
rect 2262 3682 2268 3683
rect 2478 3687 2484 3688
rect 2478 3683 2479 3687
rect 2483 3683 2484 3687
rect 2478 3682 2484 3683
rect 2694 3687 2700 3688
rect 2694 3683 2695 3687
rect 2699 3683 2700 3687
rect 2694 3682 2700 3683
rect 2910 3687 2916 3688
rect 2910 3683 2911 3687
rect 2915 3683 2916 3687
rect 2910 3682 2916 3683
rect 3118 3687 3124 3688
rect 3118 3683 3119 3687
rect 3123 3683 3124 3687
rect 3118 3682 3124 3683
rect 3318 3687 3324 3688
rect 3318 3683 3319 3687
rect 3323 3683 3324 3687
rect 3318 3682 3324 3683
rect 3518 3687 3524 3688
rect 3518 3683 3519 3687
rect 3523 3683 3524 3687
rect 3518 3682 3524 3683
rect 3726 3687 3732 3688
rect 3726 3683 3727 3687
rect 3731 3683 3732 3687
rect 3942 3684 3943 3688
rect 3947 3684 3948 3688
rect 3942 3683 3948 3684
rect 3726 3682 3732 3683
rect 2007 3681 2011 3682
rect 112 3661 114 3681
rect 110 3660 116 3661
rect 368 3660 370 3681
rect 520 3660 522 3681
rect 680 3660 682 3681
rect 848 3660 850 3681
rect 1016 3660 1018 3681
rect 1176 3660 1178 3681
rect 1328 3660 1330 3681
rect 1480 3660 1482 3681
rect 1632 3660 1634 3681
rect 1792 3660 1794 3681
rect 2008 3661 2010 3681
rect 2046 3671 2052 3672
rect 2046 3667 2047 3671
rect 2051 3667 2052 3671
rect 3942 3671 3948 3672
rect 2046 3666 2052 3667
rect 2070 3668 2076 3669
rect 2006 3660 2012 3661
rect 110 3656 111 3660
rect 115 3656 116 3660
rect 110 3655 116 3656
rect 366 3659 372 3660
rect 366 3655 367 3659
rect 371 3655 372 3659
rect 366 3654 372 3655
rect 518 3659 524 3660
rect 518 3655 519 3659
rect 523 3655 524 3659
rect 518 3654 524 3655
rect 678 3659 684 3660
rect 678 3655 679 3659
rect 683 3655 684 3659
rect 678 3654 684 3655
rect 846 3659 852 3660
rect 846 3655 847 3659
rect 851 3655 852 3659
rect 846 3654 852 3655
rect 1014 3659 1020 3660
rect 1014 3655 1015 3659
rect 1019 3655 1020 3659
rect 1014 3654 1020 3655
rect 1174 3659 1180 3660
rect 1174 3655 1175 3659
rect 1179 3655 1180 3659
rect 1174 3654 1180 3655
rect 1326 3659 1332 3660
rect 1326 3655 1327 3659
rect 1331 3655 1332 3659
rect 1326 3654 1332 3655
rect 1478 3659 1484 3660
rect 1478 3655 1479 3659
rect 1483 3655 1484 3659
rect 1478 3654 1484 3655
rect 1630 3659 1636 3660
rect 1630 3655 1631 3659
rect 1635 3655 1636 3659
rect 1630 3654 1636 3655
rect 1790 3659 1796 3660
rect 1790 3655 1791 3659
rect 1795 3655 1796 3659
rect 2006 3656 2007 3660
rect 2011 3656 2012 3660
rect 2006 3655 2012 3656
rect 1790 3654 1796 3655
rect 110 3643 116 3644
rect 110 3639 111 3643
rect 115 3639 116 3643
rect 2006 3643 2012 3644
rect 110 3638 116 3639
rect 366 3640 372 3641
rect 112 3603 114 3638
rect 366 3636 367 3640
rect 371 3636 372 3640
rect 366 3635 372 3636
rect 518 3640 524 3641
rect 518 3636 519 3640
rect 523 3636 524 3640
rect 518 3635 524 3636
rect 678 3640 684 3641
rect 678 3636 679 3640
rect 683 3636 684 3640
rect 678 3635 684 3636
rect 846 3640 852 3641
rect 846 3636 847 3640
rect 851 3636 852 3640
rect 846 3635 852 3636
rect 1014 3640 1020 3641
rect 1014 3636 1015 3640
rect 1019 3636 1020 3640
rect 1014 3635 1020 3636
rect 1174 3640 1180 3641
rect 1174 3636 1175 3640
rect 1179 3636 1180 3640
rect 1174 3635 1180 3636
rect 1326 3640 1332 3641
rect 1326 3636 1327 3640
rect 1331 3636 1332 3640
rect 1326 3635 1332 3636
rect 1478 3640 1484 3641
rect 1478 3636 1479 3640
rect 1483 3636 1484 3640
rect 1478 3635 1484 3636
rect 1630 3640 1636 3641
rect 1630 3636 1631 3640
rect 1635 3636 1636 3640
rect 1630 3635 1636 3636
rect 1790 3640 1796 3641
rect 1790 3636 1791 3640
rect 1795 3636 1796 3640
rect 2006 3639 2007 3643
rect 2011 3639 2012 3643
rect 2006 3638 2012 3639
rect 1790 3635 1796 3636
rect 368 3603 370 3635
rect 520 3603 522 3635
rect 680 3603 682 3635
rect 848 3603 850 3635
rect 1016 3603 1018 3635
rect 1176 3603 1178 3635
rect 1328 3603 1330 3635
rect 1480 3603 1482 3635
rect 1632 3603 1634 3635
rect 1792 3603 1794 3635
rect 2008 3603 2010 3638
rect 2048 3635 2050 3666
rect 2070 3664 2071 3668
rect 2075 3664 2076 3668
rect 2070 3663 2076 3664
rect 2262 3668 2268 3669
rect 2262 3664 2263 3668
rect 2267 3664 2268 3668
rect 2262 3663 2268 3664
rect 2478 3668 2484 3669
rect 2478 3664 2479 3668
rect 2483 3664 2484 3668
rect 2478 3663 2484 3664
rect 2694 3668 2700 3669
rect 2694 3664 2695 3668
rect 2699 3664 2700 3668
rect 2694 3663 2700 3664
rect 2910 3668 2916 3669
rect 2910 3664 2911 3668
rect 2915 3664 2916 3668
rect 2910 3663 2916 3664
rect 3118 3668 3124 3669
rect 3118 3664 3119 3668
rect 3123 3664 3124 3668
rect 3118 3663 3124 3664
rect 3318 3668 3324 3669
rect 3318 3664 3319 3668
rect 3323 3664 3324 3668
rect 3318 3663 3324 3664
rect 3518 3668 3524 3669
rect 3518 3664 3519 3668
rect 3523 3664 3524 3668
rect 3518 3663 3524 3664
rect 3726 3668 3732 3669
rect 3726 3664 3727 3668
rect 3731 3664 3732 3668
rect 3942 3667 3943 3671
rect 3947 3667 3948 3671
rect 3942 3666 3948 3667
rect 3726 3663 3732 3664
rect 2072 3635 2074 3663
rect 2264 3635 2266 3663
rect 2480 3635 2482 3663
rect 2696 3635 2698 3663
rect 2912 3635 2914 3663
rect 3120 3635 3122 3663
rect 3320 3635 3322 3663
rect 3520 3635 3522 3663
rect 3728 3635 3730 3663
rect 3944 3635 3946 3666
rect 2047 3634 2051 3635
rect 2047 3629 2051 3630
rect 2071 3634 2075 3635
rect 2071 3629 2075 3630
rect 2111 3634 2115 3635
rect 2111 3629 2115 3630
rect 2263 3634 2267 3635
rect 2263 3629 2267 3630
rect 2271 3634 2275 3635
rect 2271 3629 2275 3630
rect 2455 3634 2459 3635
rect 2455 3629 2459 3630
rect 2479 3634 2483 3635
rect 2479 3629 2483 3630
rect 2655 3634 2659 3635
rect 2655 3629 2659 3630
rect 2695 3634 2699 3635
rect 2695 3629 2699 3630
rect 2871 3634 2875 3635
rect 2871 3629 2875 3630
rect 2911 3634 2915 3635
rect 2911 3629 2915 3630
rect 3095 3634 3099 3635
rect 3095 3629 3099 3630
rect 3119 3634 3123 3635
rect 3119 3629 3123 3630
rect 3319 3634 3323 3635
rect 3319 3629 3323 3630
rect 3327 3634 3331 3635
rect 3327 3629 3331 3630
rect 3519 3634 3523 3635
rect 3519 3629 3523 3630
rect 3567 3634 3571 3635
rect 3567 3629 3571 3630
rect 3727 3634 3731 3635
rect 3727 3629 3731 3630
rect 3943 3634 3947 3635
rect 3943 3629 3947 3630
rect 111 3602 115 3603
rect 111 3597 115 3598
rect 271 3602 275 3603
rect 271 3597 275 3598
rect 367 3602 371 3603
rect 367 3597 371 3598
rect 415 3602 419 3603
rect 415 3597 419 3598
rect 519 3602 523 3603
rect 519 3597 523 3598
rect 575 3602 579 3603
rect 575 3597 579 3598
rect 679 3602 683 3603
rect 679 3597 683 3598
rect 735 3602 739 3603
rect 735 3597 739 3598
rect 847 3602 851 3603
rect 847 3597 851 3598
rect 895 3602 899 3603
rect 895 3597 899 3598
rect 1015 3602 1019 3603
rect 1015 3597 1019 3598
rect 1055 3602 1059 3603
rect 1055 3597 1059 3598
rect 1175 3602 1179 3603
rect 1175 3597 1179 3598
rect 1215 3602 1219 3603
rect 1215 3597 1219 3598
rect 1327 3602 1331 3603
rect 1327 3597 1331 3598
rect 1375 3602 1379 3603
rect 1375 3597 1379 3598
rect 1479 3602 1483 3603
rect 1479 3597 1483 3598
rect 1543 3602 1547 3603
rect 1543 3597 1547 3598
rect 1631 3602 1635 3603
rect 1631 3597 1635 3598
rect 1791 3602 1795 3603
rect 1791 3597 1795 3598
rect 2007 3602 2011 3603
rect 2048 3602 2050 3629
rect 2112 3605 2114 3629
rect 2272 3605 2274 3629
rect 2456 3605 2458 3629
rect 2656 3605 2658 3629
rect 2872 3605 2874 3629
rect 3096 3605 3098 3629
rect 3328 3605 3330 3629
rect 3568 3605 3570 3629
rect 2110 3604 2116 3605
rect 2007 3597 2011 3598
rect 2046 3601 2052 3602
rect 2046 3597 2047 3601
rect 2051 3597 2052 3601
rect 2110 3600 2111 3604
rect 2115 3600 2116 3604
rect 2110 3599 2116 3600
rect 2270 3604 2276 3605
rect 2270 3600 2271 3604
rect 2275 3600 2276 3604
rect 2270 3599 2276 3600
rect 2454 3604 2460 3605
rect 2454 3600 2455 3604
rect 2459 3600 2460 3604
rect 2454 3599 2460 3600
rect 2654 3604 2660 3605
rect 2654 3600 2655 3604
rect 2659 3600 2660 3604
rect 2654 3599 2660 3600
rect 2870 3604 2876 3605
rect 2870 3600 2871 3604
rect 2875 3600 2876 3604
rect 2870 3599 2876 3600
rect 3094 3604 3100 3605
rect 3094 3600 3095 3604
rect 3099 3600 3100 3604
rect 3094 3599 3100 3600
rect 3326 3604 3332 3605
rect 3326 3600 3327 3604
rect 3331 3600 3332 3604
rect 3326 3599 3332 3600
rect 3566 3604 3572 3605
rect 3566 3600 3567 3604
rect 3571 3600 3572 3604
rect 3944 3602 3946 3629
rect 3566 3599 3572 3600
rect 3942 3601 3948 3602
rect 112 3570 114 3597
rect 272 3573 274 3597
rect 416 3573 418 3597
rect 576 3573 578 3597
rect 736 3573 738 3597
rect 896 3573 898 3597
rect 1056 3573 1058 3597
rect 1216 3573 1218 3597
rect 1376 3573 1378 3597
rect 1544 3573 1546 3597
rect 270 3572 276 3573
rect 110 3569 116 3570
rect 110 3565 111 3569
rect 115 3565 116 3569
rect 270 3568 271 3572
rect 275 3568 276 3572
rect 270 3567 276 3568
rect 414 3572 420 3573
rect 414 3568 415 3572
rect 419 3568 420 3572
rect 414 3567 420 3568
rect 574 3572 580 3573
rect 574 3568 575 3572
rect 579 3568 580 3572
rect 574 3567 580 3568
rect 734 3572 740 3573
rect 734 3568 735 3572
rect 739 3568 740 3572
rect 734 3567 740 3568
rect 894 3572 900 3573
rect 894 3568 895 3572
rect 899 3568 900 3572
rect 894 3567 900 3568
rect 1054 3572 1060 3573
rect 1054 3568 1055 3572
rect 1059 3568 1060 3572
rect 1054 3567 1060 3568
rect 1214 3572 1220 3573
rect 1214 3568 1215 3572
rect 1219 3568 1220 3572
rect 1214 3567 1220 3568
rect 1374 3572 1380 3573
rect 1374 3568 1375 3572
rect 1379 3568 1380 3572
rect 1374 3567 1380 3568
rect 1542 3572 1548 3573
rect 1542 3568 1543 3572
rect 1547 3568 1548 3572
rect 2008 3570 2010 3597
rect 2046 3596 2052 3597
rect 3942 3597 3943 3601
rect 3947 3597 3948 3601
rect 3942 3596 3948 3597
rect 2110 3585 2116 3586
rect 2046 3584 2052 3585
rect 2046 3580 2047 3584
rect 2051 3580 2052 3584
rect 2110 3581 2111 3585
rect 2115 3581 2116 3585
rect 2110 3580 2116 3581
rect 2270 3585 2276 3586
rect 2270 3581 2271 3585
rect 2275 3581 2276 3585
rect 2270 3580 2276 3581
rect 2454 3585 2460 3586
rect 2454 3581 2455 3585
rect 2459 3581 2460 3585
rect 2454 3580 2460 3581
rect 2654 3585 2660 3586
rect 2654 3581 2655 3585
rect 2659 3581 2660 3585
rect 2654 3580 2660 3581
rect 2870 3585 2876 3586
rect 2870 3581 2871 3585
rect 2875 3581 2876 3585
rect 2870 3580 2876 3581
rect 3094 3585 3100 3586
rect 3094 3581 3095 3585
rect 3099 3581 3100 3585
rect 3094 3580 3100 3581
rect 3326 3585 3332 3586
rect 3326 3581 3327 3585
rect 3331 3581 3332 3585
rect 3326 3580 3332 3581
rect 3566 3585 3572 3586
rect 3566 3581 3567 3585
rect 3571 3581 3572 3585
rect 3566 3580 3572 3581
rect 3942 3584 3948 3585
rect 3942 3580 3943 3584
rect 3947 3580 3948 3584
rect 2046 3579 2052 3580
rect 1542 3567 1548 3568
rect 2006 3569 2012 3570
rect 110 3564 116 3565
rect 2006 3565 2007 3569
rect 2011 3565 2012 3569
rect 2006 3564 2012 3565
rect 270 3553 276 3554
rect 110 3552 116 3553
rect 110 3548 111 3552
rect 115 3548 116 3552
rect 270 3549 271 3553
rect 275 3549 276 3553
rect 270 3548 276 3549
rect 414 3553 420 3554
rect 414 3549 415 3553
rect 419 3549 420 3553
rect 414 3548 420 3549
rect 574 3553 580 3554
rect 574 3549 575 3553
rect 579 3549 580 3553
rect 574 3548 580 3549
rect 734 3553 740 3554
rect 734 3549 735 3553
rect 739 3549 740 3553
rect 734 3548 740 3549
rect 894 3553 900 3554
rect 894 3549 895 3553
rect 899 3549 900 3553
rect 894 3548 900 3549
rect 1054 3553 1060 3554
rect 1054 3549 1055 3553
rect 1059 3549 1060 3553
rect 1054 3548 1060 3549
rect 1214 3553 1220 3554
rect 1214 3549 1215 3553
rect 1219 3549 1220 3553
rect 1214 3548 1220 3549
rect 1374 3553 1380 3554
rect 1374 3549 1375 3553
rect 1379 3549 1380 3553
rect 1374 3548 1380 3549
rect 1542 3553 1548 3554
rect 1542 3549 1543 3553
rect 1547 3549 1548 3553
rect 1542 3548 1548 3549
rect 2006 3552 2012 3553
rect 2006 3548 2007 3552
rect 2011 3548 2012 3552
rect 110 3547 116 3548
rect 112 3519 114 3547
rect 272 3519 274 3548
rect 416 3519 418 3548
rect 576 3519 578 3548
rect 736 3519 738 3548
rect 896 3519 898 3548
rect 1056 3519 1058 3548
rect 1216 3519 1218 3548
rect 1376 3519 1378 3548
rect 1544 3519 1546 3548
rect 2006 3547 2012 3548
rect 2008 3519 2010 3547
rect 2048 3543 2050 3579
rect 2112 3543 2114 3580
rect 2272 3543 2274 3580
rect 2456 3543 2458 3580
rect 2656 3543 2658 3580
rect 2872 3543 2874 3580
rect 3096 3543 3098 3580
rect 3328 3543 3330 3580
rect 3568 3543 3570 3580
rect 3942 3579 3948 3580
rect 3944 3543 3946 3579
rect 2047 3542 2051 3543
rect 2047 3537 2051 3538
rect 2111 3542 2115 3543
rect 2111 3537 2115 3538
rect 2271 3542 2275 3543
rect 2271 3537 2275 3538
rect 2287 3542 2291 3543
rect 2287 3537 2291 3538
rect 2383 3542 2387 3543
rect 2383 3537 2387 3538
rect 2455 3542 2459 3543
rect 2455 3537 2459 3538
rect 2479 3542 2483 3543
rect 2479 3537 2483 3538
rect 2575 3542 2579 3543
rect 2575 3537 2579 3538
rect 2655 3542 2659 3543
rect 2655 3537 2659 3538
rect 2671 3542 2675 3543
rect 2671 3537 2675 3538
rect 2767 3542 2771 3543
rect 2767 3537 2771 3538
rect 2871 3542 2875 3543
rect 2871 3537 2875 3538
rect 2983 3542 2987 3543
rect 2983 3537 2987 3538
rect 3095 3542 3099 3543
rect 3095 3537 3099 3538
rect 3103 3542 3107 3543
rect 3103 3537 3107 3538
rect 3223 3542 3227 3543
rect 3223 3537 3227 3538
rect 3327 3542 3331 3543
rect 3327 3537 3331 3538
rect 3351 3542 3355 3543
rect 3351 3537 3355 3538
rect 3487 3542 3491 3543
rect 3487 3537 3491 3538
rect 3567 3542 3571 3543
rect 3567 3537 3571 3538
rect 3943 3542 3947 3543
rect 3943 3537 3947 3538
rect 111 3518 115 3519
rect 111 3513 115 3514
rect 159 3518 163 3519
rect 159 3513 163 3514
rect 271 3518 275 3519
rect 271 3513 275 3514
rect 287 3518 291 3519
rect 287 3513 291 3514
rect 415 3518 419 3519
rect 415 3513 419 3514
rect 423 3518 427 3519
rect 423 3513 427 3514
rect 559 3518 563 3519
rect 559 3513 563 3514
rect 575 3518 579 3519
rect 575 3513 579 3514
rect 695 3518 699 3519
rect 695 3513 699 3514
rect 735 3518 739 3519
rect 735 3513 739 3514
rect 831 3518 835 3519
rect 831 3513 835 3514
rect 895 3518 899 3519
rect 895 3513 899 3514
rect 967 3518 971 3519
rect 967 3513 971 3514
rect 1055 3518 1059 3519
rect 1055 3513 1059 3514
rect 1095 3518 1099 3519
rect 1095 3513 1099 3514
rect 1215 3518 1219 3519
rect 1215 3513 1219 3514
rect 1231 3518 1235 3519
rect 1231 3513 1235 3514
rect 1367 3518 1371 3519
rect 1367 3513 1371 3514
rect 1375 3518 1379 3519
rect 1375 3513 1379 3514
rect 1543 3518 1547 3519
rect 1543 3513 1547 3514
rect 2007 3518 2011 3519
rect 2048 3517 2050 3537
rect 2007 3513 2011 3514
rect 2046 3516 2052 3517
rect 2288 3516 2290 3537
rect 2384 3516 2386 3537
rect 2480 3516 2482 3537
rect 2576 3516 2578 3537
rect 2672 3516 2674 3537
rect 2768 3516 2770 3537
rect 2872 3516 2874 3537
rect 2984 3516 2986 3537
rect 3104 3516 3106 3537
rect 3224 3516 3226 3537
rect 3352 3516 3354 3537
rect 3488 3516 3490 3537
rect 3944 3517 3946 3537
rect 3942 3516 3948 3517
rect 112 3493 114 3513
rect 110 3492 116 3493
rect 160 3492 162 3513
rect 288 3492 290 3513
rect 424 3492 426 3513
rect 560 3492 562 3513
rect 696 3492 698 3513
rect 832 3492 834 3513
rect 968 3492 970 3513
rect 1096 3492 1098 3513
rect 1232 3492 1234 3513
rect 1368 3492 1370 3513
rect 2008 3493 2010 3513
rect 2046 3512 2047 3516
rect 2051 3512 2052 3516
rect 2046 3511 2052 3512
rect 2286 3515 2292 3516
rect 2286 3511 2287 3515
rect 2291 3511 2292 3515
rect 2286 3510 2292 3511
rect 2382 3515 2388 3516
rect 2382 3511 2383 3515
rect 2387 3511 2388 3515
rect 2382 3510 2388 3511
rect 2478 3515 2484 3516
rect 2478 3511 2479 3515
rect 2483 3511 2484 3515
rect 2478 3510 2484 3511
rect 2574 3515 2580 3516
rect 2574 3511 2575 3515
rect 2579 3511 2580 3515
rect 2574 3510 2580 3511
rect 2670 3515 2676 3516
rect 2670 3511 2671 3515
rect 2675 3511 2676 3515
rect 2670 3510 2676 3511
rect 2766 3515 2772 3516
rect 2766 3511 2767 3515
rect 2771 3511 2772 3515
rect 2766 3510 2772 3511
rect 2870 3515 2876 3516
rect 2870 3511 2871 3515
rect 2875 3511 2876 3515
rect 2870 3510 2876 3511
rect 2982 3515 2988 3516
rect 2982 3511 2983 3515
rect 2987 3511 2988 3515
rect 2982 3510 2988 3511
rect 3102 3515 3108 3516
rect 3102 3511 3103 3515
rect 3107 3511 3108 3515
rect 3102 3510 3108 3511
rect 3222 3515 3228 3516
rect 3222 3511 3223 3515
rect 3227 3511 3228 3515
rect 3222 3510 3228 3511
rect 3350 3515 3356 3516
rect 3350 3511 3351 3515
rect 3355 3511 3356 3515
rect 3350 3510 3356 3511
rect 3486 3515 3492 3516
rect 3486 3511 3487 3515
rect 3491 3511 3492 3515
rect 3942 3512 3943 3516
rect 3947 3512 3948 3516
rect 3942 3511 3948 3512
rect 3486 3510 3492 3511
rect 2046 3499 2052 3500
rect 2046 3495 2047 3499
rect 2051 3495 2052 3499
rect 3942 3499 3948 3500
rect 2046 3494 2052 3495
rect 2286 3496 2292 3497
rect 2006 3492 2012 3493
rect 110 3488 111 3492
rect 115 3488 116 3492
rect 110 3487 116 3488
rect 158 3491 164 3492
rect 158 3487 159 3491
rect 163 3487 164 3491
rect 158 3486 164 3487
rect 286 3491 292 3492
rect 286 3487 287 3491
rect 291 3487 292 3491
rect 286 3486 292 3487
rect 422 3491 428 3492
rect 422 3487 423 3491
rect 427 3487 428 3491
rect 422 3486 428 3487
rect 558 3491 564 3492
rect 558 3487 559 3491
rect 563 3487 564 3491
rect 558 3486 564 3487
rect 694 3491 700 3492
rect 694 3487 695 3491
rect 699 3487 700 3491
rect 694 3486 700 3487
rect 830 3491 836 3492
rect 830 3487 831 3491
rect 835 3487 836 3491
rect 830 3486 836 3487
rect 966 3491 972 3492
rect 966 3487 967 3491
rect 971 3487 972 3491
rect 966 3486 972 3487
rect 1094 3491 1100 3492
rect 1094 3487 1095 3491
rect 1099 3487 1100 3491
rect 1094 3486 1100 3487
rect 1230 3491 1236 3492
rect 1230 3487 1231 3491
rect 1235 3487 1236 3491
rect 1230 3486 1236 3487
rect 1366 3491 1372 3492
rect 1366 3487 1367 3491
rect 1371 3487 1372 3491
rect 2006 3488 2007 3492
rect 2011 3488 2012 3492
rect 2006 3487 2012 3488
rect 1366 3486 1372 3487
rect 110 3475 116 3476
rect 110 3471 111 3475
rect 115 3471 116 3475
rect 2006 3475 2012 3476
rect 110 3470 116 3471
rect 158 3472 164 3473
rect 112 3435 114 3470
rect 158 3468 159 3472
rect 163 3468 164 3472
rect 158 3467 164 3468
rect 286 3472 292 3473
rect 286 3468 287 3472
rect 291 3468 292 3472
rect 286 3467 292 3468
rect 422 3472 428 3473
rect 422 3468 423 3472
rect 427 3468 428 3472
rect 422 3467 428 3468
rect 558 3472 564 3473
rect 558 3468 559 3472
rect 563 3468 564 3472
rect 558 3467 564 3468
rect 694 3472 700 3473
rect 694 3468 695 3472
rect 699 3468 700 3472
rect 694 3467 700 3468
rect 830 3472 836 3473
rect 830 3468 831 3472
rect 835 3468 836 3472
rect 830 3467 836 3468
rect 966 3472 972 3473
rect 966 3468 967 3472
rect 971 3468 972 3472
rect 966 3467 972 3468
rect 1094 3472 1100 3473
rect 1094 3468 1095 3472
rect 1099 3468 1100 3472
rect 1094 3467 1100 3468
rect 1230 3472 1236 3473
rect 1230 3468 1231 3472
rect 1235 3468 1236 3472
rect 1230 3467 1236 3468
rect 1366 3472 1372 3473
rect 1366 3468 1367 3472
rect 1371 3468 1372 3472
rect 2006 3471 2007 3475
rect 2011 3471 2012 3475
rect 2006 3470 2012 3471
rect 1366 3467 1372 3468
rect 160 3435 162 3467
rect 288 3435 290 3467
rect 424 3435 426 3467
rect 560 3435 562 3467
rect 696 3435 698 3467
rect 832 3435 834 3467
rect 968 3435 970 3467
rect 1096 3435 1098 3467
rect 1232 3435 1234 3467
rect 1368 3435 1370 3467
rect 2008 3435 2010 3470
rect 2048 3467 2050 3494
rect 2286 3492 2287 3496
rect 2291 3492 2292 3496
rect 2286 3491 2292 3492
rect 2382 3496 2388 3497
rect 2382 3492 2383 3496
rect 2387 3492 2388 3496
rect 2382 3491 2388 3492
rect 2478 3496 2484 3497
rect 2478 3492 2479 3496
rect 2483 3492 2484 3496
rect 2478 3491 2484 3492
rect 2574 3496 2580 3497
rect 2574 3492 2575 3496
rect 2579 3492 2580 3496
rect 2574 3491 2580 3492
rect 2670 3496 2676 3497
rect 2670 3492 2671 3496
rect 2675 3492 2676 3496
rect 2670 3491 2676 3492
rect 2766 3496 2772 3497
rect 2766 3492 2767 3496
rect 2771 3492 2772 3496
rect 2766 3491 2772 3492
rect 2870 3496 2876 3497
rect 2870 3492 2871 3496
rect 2875 3492 2876 3496
rect 2870 3491 2876 3492
rect 2982 3496 2988 3497
rect 2982 3492 2983 3496
rect 2987 3492 2988 3496
rect 2982 3491 2988 3492
rect 3102 3496 3108 3497
rect 3102 3492 3103 3496
rect 3107 3492 3108 3496
rect 3102 3491 3108 3492
rect 3222 3496 3228 3497
rect 3222 3492 3223 3496
rect 3227 3492 3228 3496
rect 3222 3491 3228 3492
rect 3350 3496 3356 3497
rect 3350 3492 3351 3496
rect 3355 3492 3356 3496
rect 3350 3491 3356 3492
rect 3486 3496 3492 3497
rect 3486 3492 3487 3496
rect 3491 3492 3492 3496
rect 3942 3495 3943 3499
rect 3947 3495 3948 3499
rect 3942 3494 3948 3495
rect 3486 3491 3492 3492
rect 2288 3467 2290 3491
rect 2384 3467 2386 3491
rect 2480 3467 2482 3491
rect 2576 3467 2578 3491
rect 2672 3467 2674 3491
rect 2768 3467 2770 3491
rect 2872 3467 2874 3491
rect 2984 3467 2986 3491
rect 3104 3467 3106 3491
rect 3224 3467 3226 3491
rect 3352 3467 3354 3491
rect 3488 3467 3490 3491
rect 3944 3467 3946 3494
rect 2047 3466 2051 3467
rect 2047 3461 2051 3462
rect 2287 3466 2291 3467
rect 2287 3461 2291 3462
rect 2383 3466 2387 3467
rect 2383 3461 2387 3462
rect 2479 3466 2483 3467
rect 2479 3461 2483 3462
rect 2487 3466 2491 3467
rect 2487 3461 2491 3462
rect 2575 3466 2579 3467
rect 2575 3461 2579 3462
rect 2583 3466 2587 3467
rect 2583 3461 2587 3462
rect 2671 3466 2675 3467
rect 2671 3461 2675 3462
rect 2679 3466 2683 3467
rect 2679 3461 2683 3462
rect 2767 3466 2771 3467
rect 2767 3461 2771 3462
rect 2783 3466 2787 3467
rect 2783 3461 2787 3462
rect 2871 3466 2875 3467
rect 2871 3461 2875 3462
rect 2895 3466 2899 3467
rect 2895 3461 2899 3462
rect 2983 3466 2987 3467
rect 2983 3461 2987 3462
rect 3015 3466 3019 3467
rect 3015 3461 3019 3462
rect 3103 3466 3107 3467
rect 3103 3461 3107 3462
rect 3143 3466 3147 3467
rect 3143 3461 3147 3462
rect 3223 3466 3227 3467
rect 3223 3461 3227 3462
rect 3271 3466 3275 3467
rect 3271 3461 3275 3462
rect 3351 3466 3355 3467
rect 3351 3461 3355 3462
rect 3407 3466 3411 3467
rect 3407 3461 3411 3462
rect 3487 3466 3491 3467
rect 3487 3461 3491 3462
rect 3943 3466 3947 3467
rect 3943 3461 3947 3462
rect 111 3434 115 3435
rect 111 3429 115 3430
rect 135 3434 139 3435
rect 135 3429 139 3430
rect 159 3434 163 3435
rect 159 3429 163 3430
rect 247 3434 251 3435
rect 247 3429 251 3430
rect 287 3434 291 3435
rect 287 3429 291 3430
rect 383 3434 387 3435
rect 383 3429 387 3430
rect 423 3434 427 3435
rect 423 3429 427 3430
rect 527 3434 531 3435
rect 527 3429 531 3430
rect 559 3434 563 3435
rect 559 3429 563 3430
rect 671 3434 675 3435
rect 671 3429 675 3430
rect 695 3434 699 3435
rect 695 3429 699 3430
rect 815 3434 819 3435
rect 815 3429 819 3430
rect 831 3434 835 3435
rect 831 3429 835 3430
rect 967 3434 971 3435
rect 967 3429 971 3430
rect 1095 3434 1099 3435
rect 1095 3429 1099 3430
rect 1119 3434 1123 3435
rect 1119 3429 1123 3430
rect 1231 3434 1235 3435
rect 1231 3429 1235 3430
rect 1271 3434 1275 3435
rect 1271 3429 1275 3430
rect 1367 3434 1371 3435
rect 1367 3429 1371 3430
rect 2007 3434 2011 3435
rect 2048 3434 2050 3461
rect 2488 3437 2490 3461
rect 2584 3437 2586 3461
rect 2680 3437 2682 3461
rect 2784 3437 2786 3461
rect 2896 3437 2898 3461
rect 3016 3437 3018 3461
rect 3144 3437 3146 3461
rect 3272 3437 3274 3461
rect 3408 3437 3410 3461
rect 2486 3436 2492 3437
rect 2007 3429 2011 3430
rect 2046 3433 2052 3434
rect 2046 3429 2047 3433
rect 2051 3429 2052 3433
rect 2486 3432 2487 3436
rect 2491 3432 2492 3436
rect 2486 3431 2492 3432
rect 2582 3436 2588 3437
rect 2582 3432 2583 3436
rect 2587 3432 2588 3436
rect 2582 3431 2588 3432
rect 2678 3436 2684 3437
rect 2678 3432 2679 3436
rect 2683 3432 2684 3436
rect 2678 3431 2684 3432
rect 2782 3436 2788 3437
rect 2782 3432 2783 3436
rect 2787 3432 2788 3436
rect 2782 3431 2788 3432
rect 2894 3436 2900 3437
rect 2894 3432 2895 3436
rect 2899 3432 2900 3436
rect 2894 3431 2900 3432
rect 3014 3436 3020 3437
rect 3014 3432 3015 3436
rect 3019 3432 3020 3436
rect 3014 3431 3020 3432
rect 3142 3436 3148 3437
rect 3142 3432 3143 3436
rect 3147 3432 3148 3436
rect 3142 3431 3148 3432
rect 3270 3436 3276 3437
rect 3270 3432 3271 3436
rect 3275 3432 3276 3436
rect 3270 3431 3276 3432
rect 3406 3436 3412 3437
rect 3406 3432 3407 3436
rect 3411 3432 3412 3436
rect 3944 3434 3946 3461
rect 3406 3431 3412 3432
rect 3942 3433 3948 3434
rect 112 3402 114 3429
rect 136 3405 138 3429
rect 248 3405 250 3429
rect 384 3405 386 3429
rect 528 3405 530 3429
rect 672 3405 674 3429
rect 816 3405 818 3429
rect 968 3405 970 3429
rect 1120 3405 1122 3429
rect 1272 3405 1274 3429
rect 134 3404 140 3405
rect 110 3401 116 3402
rect 110 3397 111 3401
rect 115 3397 116 3401
rect 134 3400 135 3404
rect 139 3400 140 3404
rect 134 3399 140 3400
rect 246 3404 252 3405
rect 246 3400 247 3404
rect 251 3400 252 3404
rect 246 3399 252 3400
rect 382 3404 388 3405
rect 382 3400 383 3404
rect 387 3400 388 3404
rect 382 3399 388 3400
rect 526 3404 532 3405
rect 526 3400 527 3404
rect 531 3400 532 3404
rect 526 3399 532 3400
rect 670 3404 676 3405
rect 670 3400 671 3404
rect 675 3400 676 3404
rect 670 3399 676 3400
rect 814 3404 820 3405
rect 814 3400 815 3404
rect 819 3400 820 3404
rect 814 3399 820 3400
rect 966 3404 972 3405
rect 966 3400 967 3404
rect 971 3400 972 3404
rect 966 3399 972 3400
rect 1118 3404 1124 3405
rect 1118 3400 1119 3404
rect 1123 3400 1124 3404
rect 1118 3399 1124 3400
rect 1270 3404 1276 3405
rect 1270 3400 1271 3404
rect 1275 3400 1276 3404
rect 2008 3402 2010 3429
rect 2046 3428 2052 3429
rect 3942 3429 3943 3433
rect 3947 3429 3948 3433
rect 3942 3428 3948 3429
rect 2486 3417 2492 3418
rect 2046 3416 2052 3417
rect 2046 3412 2047 3416
rect 2051 3412 2052 3416
rect 2486 3413 2487 3417
rect 2491 3413 2492 3417
rect 2486 3412 2492 3413
rect 2582 3417 2588 3418
rect 2582 3413 2583 3417
rect 2587 3413 2588 3417
rect 2582 3412 2588 3413
rect 2678 3417 2684 3418
rect 2678 3413 2679 3417
rect 2683 3413 2684 3417
rect 2678 3412 2684 3413
rect 2782 3417 2788 3418
rect 2782 3413 2783 3417
rect 2787 3413 2788 3417
rect 2782 3412 2788 3413
rect 2894 3417 2900 3418
rect 2894 3413 2895 3417
rect 2899 3413 2900 3417
rect 2894 3412 2900 3413
rect 3014 3417 3020 3418
rect 3014 3413 3015 3417
rect 3019 3413 3020 3417
rect 3014 3412 3020 3413
rect 3142 3417 3148 3418
rect 3142 3413 3143 3417
rect 3147 3413 3148 3417
rect 3142 3412 3148 3413
rect 3270 3417 3276 3418
rect 3270 3413 3271 3417
rect 3275 3413 3276 3417
rect 3270 3412 3276 3413
rect 3406 3417 3412 3418
rect 3406 3413 3407 3417
rect 3411 3413 3412 3417
rect 3406 3412 3412 3413
rect 3942 3416 3948 3417
rect 3942 3412 3943 3416
rect 3947 3412 3948 3416
rect 2046 3411 2052 3412
rect 1270 3399 1276 3400
rect 2006 3401 2012 3402
rect 110 3396 116 3397
rect 2006 3397 2007 3401
rect 2011 3397 2012 3401
rect 2006 3396 2012 3397
rect 134 3385 140 3386
rect 110 3384 116 3385
rect 110 3380 111 3384
rect 115 3380 116 3384
rect 134 3381 135 3385
rect 139 3381 140 3385
rect 134 3380 140 3381
rect 246 3385 252 3386
rect 246 3381 247 3385
rect 251 3381 252 3385
rect 246 3380 252 3381
rect 382 3385 388 3386
rect 382 3381 383 3385
rect 387 3381 388 3385
rect 382 3380 388 3381
rect 526 3385 532 3386
rect 526 3381 527 3385
rect 531 3381 532 3385
rect 526 3380 532 3381
rect 670 3385 676 3386
rect 670 3381 671 3385
rect 675 3381 676 3385
rect 670 3380 676 3381
rect 814 3385 820 3386
rect 814 3381 815 3385
rect 819 3381 820 3385
rect 814 3380 820 3381
rect 966 3385 972 3386
rect 966 3381 967 3385
rect 971 3381 972 3385
rect 966 3380 972 3381
rect 1118 3385 1124 3386
rect 1118 3381 1119 3385
rect 1123 3381 1124 3385
rect 1118 3380 1124 3381
rect 1270 3385 1276 3386
rect 1270 3381 1271 3385
rect 1275 3381 1276 3385
rect 1270 3380 1276 3381
rect 2006 3384 2012 3385
rect 2006 3380 2007 3384
rect 2011 3380 2012 3384
rect 2048 3383 2050 3411
rect 2488 3383 2490 3412
rect 2584 3383 2586 3412
rect 2680 3383 2682 3412
rect 2784 3383 2786 3412
rect 2896 3383 2898 3412
rect 3016 3383 3018 3412
rect 3144 3383 3146 3412
rect 3272 3383 3274 3412
rect 3408 3383 3410 3412
rect 3942 3411 3948 3412
rect 3944 3383 3946 3411
rect 110 3379 116 3380
rect 112 3351 114 3379
rect 136 3351 138 3380
rect 248 3351 250 3380
rect 384 3351 386 3380
rect 528 3351 530 3380
rect 672 3351 674 3380
rect 816 3351 818 3380
rect 968 3351 970 3380
rect 1120 3351 1122 3380
rect 1272 3351 1274 3380
rect 2006 3379 2012 3380
rect 2047 3382 2051 3383
rect 2008 3351 2010 3379
rect 2047 3377 2051 3378
rect 2351 3382 2355 3383
rect 2351 3377 2355 3378
rect 2479 3382 2483 3383
rect 2479 3377 2483 3378
rect 2487 3382 2491 3383
rect 2487 3377 2491 3378
rect 2583 3382 2587 3383
rect 2583 3377 2587 3378
rect 2615 3382 2619 3383
rect 2615 3377 2619 3378
rect 2679 3382 2683 3383
rect 2679 3377 2683 3378
rect 2751 3382 2755 3383
rect 2751 3377 2755 3378
rect 2783 3382 2787 3383
rect 2783 3377 2787 3378
rect 2887 3382 2891 3383
rect 2887 3377 2891 3378
rect 2895 3382 2899 3383
rect 2895 3377 2899 3378
rect 3015 3382 3019 3383
rect 3015 3377 3019 3378
rect 3023 3382 3027 3383
rect 3023 3377 3027 3378
rect 3143 3382 3147 3383
rect 3143 3377 3147 3378
rect 3159 3382 3163 3383
rect 3159 3377 3163 3378
rect 3271 3382 3275 3383
rect 3271 3377 3275 3378
rect 3303 3382 3307 3383
rect 3303 3377 3307 3378
rect 3407 3382 3411 3383
rect 3407 3377 3411 3378
rect 3943 3382 3947 3383
rect 3943 3377 3947 3378
rect 2048 3357 2050 3377
rect 2046 3356 2052 3357
rect 2352 3356 2354 3377
rect 2480 3356 2482 3377
rect 2616 3356 2618 3377
rect 2752 3356 2754 3377
rect 2888 3356 2890 3377
rect 3024 3356 3026 3377
rect 3160 3356 3162 3377
rect 3304 3356 3306 3377
rect 3944 3357 3946 3377
rect 3942 3356 3948 3357
rect 2046 3352 2047 3356
rect 2051 3352 2052 3356
rect 2046 3351 2052 3352
rect 2350 3355 2356 3356
rect 2350 3351 2351 3355
rect 2355 3351 2356 3355
rect 111 3350 115 3351
rect 111 3345 115 3346
rect 135 3350 139 3351
rect 135 3345 139 3346
rect 247 3350 251 3351
rect 247 3345 251 3346
rect 263 3350 267 3351
rect 263 3345 267 3346
rect 383 3350 387 3351
rect 383 3345 387 3346
rect 431 3350 435 3351
rect 431 3345 435 3346
rect 527 3350 531 3351
rect 527 3345 531 3346
rect 599 3350 603 3351
rect 599 3345 603 3346
rect 671 3350 675 3351
rect 671 3345 675 3346
rect 767 3350 771 3351
rect 767 3345 771 3346
rect 815 3350 819 3351
rect 815 3345 819 3346
rect 927 3350 931 3351
rect 927 3345 931 3346
rect 967 3350 971 3351
rect 967 3345 971 3346
rect 1087 3350 1091 3351
rect 1087 3345 1091 3346
rect 1119 3350 1123 3351
rect 1119 3345 1123 3346
rect 1239 3350 1243 3351
rect 1239 3345 1243 3346
rect 1271 3350 1275 3351
rect 1271 3345 1275 3346
rect 1391 3350 1395 3351
rect 1391 3345 1395 3346
rect 1551 3350 1555 3351
rect 1551 3345 1555 3346
rect 2007 3350 2011 3351
rect 2350 3350 2356 3351
rect 2478 3355 2484 3356
rect 2478 3351 2479 3355
rect 2483 3351 2484 3355
rect 2478 3350 2484 3351
rect 2614 3355 2620 3356
rect 2614 3351 2615 3355
rect 2619 3351 2620 3355
rect 2614 3350 2620 3351
rect 2750 3355 2756 3356
rect 2750 3351 2751 3355
rect 2755 3351 2756 3355
rect 2750 3350 2756 3351
rect 2886 3355 2892 3356
rect 2886 3351 2887 3355
rect 2891 3351 2892 3355
rect 2886 3350 2892 3351
rect 3022 3355 3028 3356
rect 3022 3351 3023 3355
rect 3027 3351 3028 3355
rect 3022 3350 3028 3351
rect 3158 3355 3164 3356
rect 3158 3351 3159 3355
rect 3163 3351 3164 3355
rect 3158 3350 3164 3351
rect 3302 3355 3308 3356
rect 3302 3351 3303 3355
rect 3307 3351 3308 3355
rect 3942 3352 3943 3356
rect 3947 3352 3948 3356
rect 3942 3351 3948 3352
rect 3302 3350 3308 3351
rect 2007 3345 2011 3346
rect 112 3325 114 3345
rect 110 3324 116 3325
rect 136 3324 138 3345
rect 264 3324 266 3345
rect 432 3324 434 3345
rect 600 3324 602 3345
rect 768 3324 770 3345
rect 928 3324 930 3345
rect 1088 3324 1090 3345
rect 1240 3324 1242 3345
rect 1392 3324 1394 3345
rect 1552 3324 1554 3345
rect 2008 3325 2010 3345
rect 2046 3339 2052 3340
rect 2046 3335 2047 3339
rect 2051 3335 2052 3339
rect 3942 3339 3948 3340
rect 2046 3334 2052 3335
rect 2350 3336 2356 3337
rect 2006 3324 2012 3325
rect 110 3320 111 3324
rect 115 3320 116 3324
rect 110 3319 116 3320
rect 134 3323 140 3324
rect 134 3319 135 3323
rect 139 3319 140 3323
rect 134 3318 140 3319
rect 262 3323 268 3324
rect 262 3319 263 3323
rect 267 3319 268 3323
rect 262 3318 268 3319
rect 430 3323 436 3324
rect 430 3319 431 3323
rect 435 3319 436 3323
rect 430 3318 436 3319
rect 598 3323 604 3324
rect 598 3319 599 3323
rect 603 3319 604 3323
rect 598 3318 604 3319
rect 766 3323 772 3324
rect 766 3319 767 3323
rect 771 3319 772 3323
rect 766 3318 772 3319
rect 926 3323 932 3324
rect 926 3319 927 3323
rect 931 3319 932 3323
rect 926 3318 932 3319
rect 1086 3323 1092 3324
rect 1086 3319 1087 3323
rect 1091 3319 1092 3323
rect 1086 3318 1092 3319
rect 1238 3323 1244 3324
rect 1238 3319 1239 3323
rect 1243 3319 1244 3323
rect 1238 3318 1244 3319
rect 1390 3323 1396 3324
rect 1390 3319 1391 3323
rect 1395 3319 1396 3323
rect 1390 3318 1396 3319
rect 1550 3323 1556 3324
rect 1550 3319 1551 3323
rect 1555 3319 1556 3323
rect 2006 3320 2007 3324
rect 2011 3320 2012 3324
rect 2006 3319 2012 3320
rect 1550 3318 1556 3319
rect 110 3307 116 3308
rect 110 3303 111 3307
rect 115 3303 116 3307
rect 2006 3307 2012 3308
rect 110 3302 116 3303
rect 134 3304 140 3305
rect 112 3267 114 3302
rect 134 3300 135 3304
rect 139 3300 140 3304
rect 134 3299 140 3300
rect 262 3304 268 3305
rect 262 3300 263 3304
rect 267 3300 268 3304
rect 262 3299 268 3300
rect 430 3304 436 3305
rect 430 3300 431 3304
rect 435 3300 436 3304
rect 430 3299 436 3300
rect 598 3304 604 3305
rect 598 3300 599 3304
rect 603 3300 604 3304
rect 598 3299 604 3300
rect 766 3304 772 3305
rect 766 3300 767 3304
rect 771 3300 772 3304
rect 766 3299 772 3300
rect 926 3304 932 3305
rect 926 3300 927 3304
rect 931 3300 932 3304
rect 926 3299 932 3300
rect 1086 3304 1092 3305
rect 1086 3300 1087 3304
rect 1091 3300 1092 3304
rect 1086 3299 1092 3300
rect 1238 3304 1244 3305
rect 1238 3300 1239 3304
rect 1243 3300 1244 3304
rect 1238 3299 1244 3300
rect 1390 3304 1396 3305
rect 1390 3300 1391 3304
rect 1395 3300 1396 3304
rect 1390 3299 1396 3300
rect 1550 3304 1556 3305
rect 1550 3300 1551 3304
rect 1555 3300 1556 3304
rect 2006 3303 2007 3307
rect 2011 3303 2012 3307
rect 2048 3303 2050 3334
rect 2350 3332 2351 3336
rect 2355 3332 2356 3336
rect 2350 3331 2356 3332
rect 2478 3336 2484 3337
rect 2478 3332 2479 3336
rect 2483 3332 2484 3336
rect 2478 3331 2484 3332
rect 2614 3336 2620 3337
rect 2614 3332 2615 3336
rect 2619 3332 2620 3336
rect 2614 3331 2620 3332
rect 2750 3336 2756 3337
rect 2750 3332 2751 3336
rect 2755 3332 2756 3336
rect 2750 3331 2756 3332
rect 2886 3336 2892 3337
rect 2886 3332 2887 3336
rect 2891 3332 2892 3336
rect 2886 3331 2892 3332
rect 3022 3336 3028 3337
rect 3022 3332 3023 3336
rect 3027 3332 3028 3336
rect 3022 3331 3028 3332
rect 3158 3336 3164 3337
rect 3158 3332 3159 3336
rect 3163 3332 3164 3336
rect 3158 3331 3164 3332
rect 3302 3336 3308 3337
rect 3302 3332 3303 3336
rect 3307 3332 3308 3336
rect 3942 3335 3943 3339
rect 3947 3335 3948 3339
rect 3942 3334 3948 3335
rect 3302 3331 3308 3332
rect 2352 3303 2354 3331
rect 2480 3303 2482 3331
rect 2616 3303 2618 3331
rect 2752 3303 2754 3331
rect 2888 3303 2890 3331
rect 3024 3303 3026 3331
rect 3160 3303 3162 3331
rect 3304 3303 3306 3331
rect 3944 3303 3946 3334
rect 2006 3302 2012 3303
rect 2047 3302 2051 3303
rect 1550 3299 1556 3300
rect 136 3267 138 3299
rect 264 3267 266 3299
rect 432 3267 434 3299
rect 600 3267 602 3299
rect 768 3267 770 3299
rect 928 3267 930 3299
rect 1088 3267 1090 3299
rect 1240 3267 1242 3299
rect 1392 3267 1394 3299
rect 1552 3267 1554 3299
rect 2008 3267 2010 3302
rect 2047 3297 2051 3298
rect 2127 3302 2131 3303
rect 2127 3297 2131 3298
rect 2295 3302 2299 3303
rect 2295 3297 2299 3298
rect 2351 3302 2355 3303
rect 2351 3297 2355 3298
rect 2455 3302 2459 3303
rect 2455 3297 2459 3298
rect 2479 3302 2483 3303
rect 2479 3297 2483 3298
rect 2615 3302 2619 3303
rect 2615 3297 2619 3298
rect 2751 3302 2755 3303
rect 2751 3297 2755 3298
rect 2775 3302 2779 3303
rect 2775 3297 2779 3298
rect 2887 3302 2891 3303
rect 2887 3297 2891 3298
rect 2935 3302 2939 3303
rect 2935 3297 2939 3298
rect 3023 3302 3027 3303
rect 3023 3297 3027 3298
rect 3095 3302 3099 3303
rect 3095 3297 3099 3298
rect 3159 3302 3163 3303
rect 3159 3297 3163 3298
rect 3263 3302 3267 3303
rect 3263 3297 3267 3298
rect 3303 3302 3307 3303
rect 3303 3297 3307 3298
rect 3943 3302 3947 3303
rect 3943 3297 3947 3298
rect 2048 3270 2050 3297
rect 2128 3273 2130 3297
rect 2296 3273 2298 3297
rect 2456 3273 2458 3297
rect 2616 3273 2618 3297
rect 2776 3273 2778 3297
rect 2936 3273 2938 3297
rect 3096 3273 3098 3297
rect 3264 3273 3266 3297
rect 2126 3272 2132 3273
rect 2046 3269 2052 3270
rect 111 3266 115 3267
rect 111 3261 115 3262
rect 135 3266 139 3267
rect 135 3261 139 3262
rect 143 3266 147 3267
rect 143 3261 147 3262
rect 263 3266 267 3267
rect 263 3261 267 3262
rect 295 3266 299 3267
rect 295 3261 299 3262
rect 431 3266 435 3267
rect 431 3261 435 3262
rect 455 3266 459 3267
rect 455 3261 459 3262
rect 599 3266 603 3267
rect 599 3261 603 3262
rect 623 3266 627 3267
rect 623 3261 627 3262
rect 767 3266 771 3267
rect 767 3261 771 3262
rect 791 3266 795 3267
rect 791 3261 795 3262
rect 927 3266 931 3267
rect 927 3261 931 3262
rect 959 3266 963 3267
rect 959 3261 963 3262
rect 1087 3266 1091 3267
rect 1087 3261 1091 3262
rect 1127 3266 1131 3267
rect 1127 3261 1131 3262
rect 1239 3266 1243 3267
rect 1239 3261 1243 3262
rect 1303 3266 1307 3267
rect 1303 3261 1307 3262
rect 1391 3266 1395 3267
rect 1391 3261 1395 3262
rect 1479 3266 1483 3267
rect 1479 3261 1483 3262
rect 1551 3266 1555 3267
rect 1551 3261 1555 3262
rect 2007 3266 2011 3267
rect 2046 3265 2047 3269
rect 2051 3265 2052 3269
rect 2126 3268 2127 3272
rect 2131 3268 2132 3272
rect 2126 3267 2132 3268
rect 2294 3272 2300 3273
rect 2294 3268 2295 3272
rect 2299 3268 2300 3272
rect 2294 3267 2300 3268
rect 2454 3272 2460 3273
rect 2454 3268 2455 3272
rect 2459 3268 2460 3272
rect 2454 3267 2460 3268
rect 2614 3272 2620 3273
rect 2614 3268 2615 3272
rect 2619 3268 2620 3272
rect 2614 3267 2620 3268
rect 2774 3272 2780 3273
rect 2774 3268 2775 3272
rect 2779 3268 2780 3272
rect 2774 3267 2780 3268
rect 2934 3272 2940 3273
rect 2934 3268 2935 3272
rect 2939 3268 2940 3272
rect 2934 3267 2940 3268
rect 3094 3272 3100 3273
rect 3094 3268 3095 3272
rect 3099 3268 3100 3272
rect 3094 3267 3100 3268
rect 3262 3272 3268 3273
rect 3262 3268 3263 3272
rect 3267 3268 3268 3272
rect 3944 3270 3946 3297
rect 3262 3267 3268 3268
rect 3942 3269 3948 3270
rect 2046 3264 2052 3265
rect 3942 3265 3943 3269
rect 3947 3265 3948 3269
rect 3942 3264 3948 3265
rect 2007 3261 2011 3262
rect 112 3234 114 3261
rect 144 3237 146 3261
rect 296 3237 298 3261
rect 456 3237 458 3261
rect 624 3237 626 3261
rect 792 3237 794 3261
rect 960 3237 962 3261
rect 1128 3237 1130 3261
rect 1304 3237 1306 3261
rect 1480 3237 1482 3261
rect 142 3236 148 3237
rect 110 3233 116 3234
rect 110 3229 111 3233
rect 115 3229 116 3233
rect 142 3232 143 3236
rect 147 3232 148 3236
rect 142 3231 148 3232
rect 294 3236 300 3237
rect 294 3232 295 3236
rect 299 3232 300 3236
rect 294 3231 300 3232
rect 454 3236 460 3237
rect 454 3232 455 3236
rect 459 3232 460 3236
rect 454 3231 460 3232
rect 622 3236 628 3237
rect 622 3232 623 3236
rect 627 3232 628 3236
rect 622 3231 628 3232
rect 790 3236 796 3237
rect 790 3232 791 3236
rect 795 3232 796 3236
rect 790 3231 796 3232
rect 958 3236 964 3237
rect 958 3232 959 3236
rect 963 3232 964 3236
rect 958 3231 964 3232
rect 1126 3236 1132 3237
rect 1126 3232 1127 3236
rect 1131 3232 1132 3236
rect 1126 3231 1132 3232
rect 1302 3236 1308 3237
rect 1302 3232 1303 3236
rect 1307 3232 1308 3236
rect 1302 3231 1308 3232
rect 1478 3236 1484 3237
rect 1478 3232 1479 3236
rect 1483 3232 1484 3236
rect 2008 3234 2010 3261
rect 2126 3253 2132 3254
rect 2046 3252 2052 3253
rect 2046 3248 2047 3252
rect 2051 3248 2052 3252
rect 2126 3249 2127 3253
rect 2131 3249 2132 3253
rect 2126 3248 2132 3249
rect 2294 3253 2300 3254
rect 2294 3249 2295 3253
rect 2299 3249 2300 3253
rect 2294 3248 2300 3249
rect 2454 3253 2460 3254
rect 2454 3249 2455 3253
rect 2459 3249 2460 3253
rect 2454 3248 2460 3249
rect 2614 3253 2620 3254
rect 2614 3249 2615 3253
rect 2619 3249 2620 3253
rect 2614 3248 2620 3249
rect 2774 3253 2780 3254
rect 2774 3249 2775 3253
rect 2779 3249 2780 3253
rect 2774 3248 2780 3249
rect 2934 3253 2940 3254
rect 2934 3249 2935 3253
rect 2939 3249 2940 3253
rect 2934 3248 2940 3249
rect 3094 3253 3100 3254
rect 3094 3249 3095 3253
rect 3099 3249 3100 3253
rect 3094 3248 3100 3249
rect 3262 3253 3268 3254
rect 3262 3249 3263 3253
rect 3267 3249 3268 3253
rect 3262 3248 3268 3249
rect 3942 3252 3948 3253
rect 3942 3248 3943 3252
rect 3947 3248 3948 3252
rect 2046 3247 2052 3248
rect 1478 3231 1484 3232
rect 2006 3233 2012 3234
rect 110 3228 116 3229
rect 2006 3229 2007 3233
rect 2011 3229 2012 3233
rect 2006 3228 2012 3229
rect 2048 3227 2050 3247
rect 2128 3227 2130 3248
rect 2296 3227 2298 3248
rect 2456 3227 2458 3248
rect 2616 3227 2618 3248
rect 2776 3227 2778 3248
rect 2936 3227 2938 3248
rect 3096 3227 3098 3248
rect 3264 3227 3266 3248
rect 3942 3247 3948 3248
rect 3944 3227 3946 3247
rect 2047 3226 2051 3227
rect 2047 3221 2051 3222
rect 2071 3226 2075 3227
rect 2071 3221 2075 3222
rect 2127 3226 2131 3227
rect 2127 3221 2131 3222
rect 2207 3226 2211 3227
rect 2207 3221 2211 3222
rect 2295 3226 2299 3227
rect 2295 3221 2299 3222
rect 2375 3226 2379 3227
rect 2375 3221 2379 3222
rect 2455 3226 2459 3227
rect 2455 3221 2459 3222
rect 2543 3226 2547 3227
rect 2543 3221 2547 3222
rect 2615 3226 2619 3227
rect 2615 3221 2619 3222
rect 2703 3226 2707 3227
rect 2703 3221 2707 3222
rect 2775 3226 2779 3227
rect 2775 3221 2779 3222
rect 2863 3226 2867 3227
rect 2863 3221 2867 3222
rect 2935 3226 2939 3227
rect 2935 3221 2939 3222
rect 3015 3226 3019 3227
rect 3015 3221 3019 3222
rect 3095 3226 3099 3227
rect 3095 3221 3099 3222
rect 3167 3226 3171 3227
rect 3167 3221 3171 3222
rect 3263 3226 3267 3227
rect 3263 3221 3267 3222
rect 3327 3226 3331 3227
rect 3327 3221 3331 3222
rect 3943 3226 3947 3227
rect 3943 3221 3947 3222
rect 142 3217 148 3218
rect 110 3216 116 3217
rect 110 3212 111 3216
rect 115 3212 116 3216
rect 142 3213 143 3217
rect 147 3213 148 3217
rect 142 3212 148 3213
rect 294 3217 300 3218
rect 294 3213 295 3217
rect 299 3213 300 3217
rect 294 3212 300 3213
rect 454 3217 460 3218
rect 454 3213 455 3217
rect 459 3213 460 3217
rect 454 3212 460 3213
rect 622 3217 628 3218
rect 622 3213 623 3217
rect 627 3213 628 3217
rect 622 3212 628 3213
rect 790 3217 796 3218
rect 790 3213 791 3217
rect 795 3213 796 3217
rect 790 3212 796 3213
rect 958 3217 964 3218
rect 958 3213 959 3217
rect 963 3213 964 3217
rect 958 3212 964 3213
rect 1126 3217 1132 3218
rect 1126 3213 1127 3217
rect 1131 3213 1132 3217
rect 1126 3212 1132 3213
rect 1302 3217 1308 3218
rect 1302 3213 1303 3217
rect 1307 3213 1308 3217
rect 1302 3212 1308 3213
rect 1478 3217 1484 3218
rect 1478 3213 1479 3217
rect 1483 3213 1484 3217
rect 1478 3212 1484 3213
rect 2006 3216 2012 3217
rect 2006 3212 2007 3216
rect 2011 3212 2012 3216
rect 110 3211 116 3212
rect 112 3191 114 3211
rect 144 3191 146 3212
rect 296 3191 298 3212
rect 456 3191 458 3212
rect 624 3191 626 3212
rect 792 3191 794 3212
rect 960 3191 962 3212
rect 1128 3191 1130 3212
rect 1304 3191 1306 3212
rect 1480 3191 1482 3212
rect 2006 3211 2012 3212
rect 2008 3191 2010 3211
rect 2048 3201 2050 3221
rect 2046 3200 2052 3201
rect 2072 3200 2074 3221
rect 2208 3200 2210 3221
rect 2376 3200 2378 3221
rect 2544 3200 2546 3221
rect 2704 3200 2706 3221
rect 2864 3200 2866 3221
rect 3016 3200 3018 3221
rect 3168 3200 3170 3221
rect 3328 3200 3330 3221
rect 3944 3201 3946 3221
rect 3942 3200 3948 3201
rect 2046 3196 2047 3200
rect 2051 3196 2052 3200
rect 2046 3195 2052 3196
rect 2070 3199 2076 3200
rect 2070 3195 2071 3199
rect 2075 3195 2076 3199
rect 2070 3194 2076 3195
rect 2206 3199 2212 3200
rect 2206 3195 2207 3199
rect 2211 3195 2212 3199
rect 2206 3194 2212 3195
rect 2374 3199 2380 3200
rect 2374 3195 2375 3199
rect 2379 3195 2380 3199
rect 2374 3194 2380 3195
rect 2542 3199 2548 3200
rect 2542 3195 2543 3199
rect 2547 3195 2548 3199
rect 2542 3194 2548 3195
rect 2702 3199 2708 3200
rect 2702 3195 2703 3199
rect 2707 3195 2708 3199
rect 2702 3194 2708 3195
rect 2862 3199 2868 3200
rect 2862 3195 2863 3199
rect 2867 3195 2868 3199
rect 2862 3194 2868 3195
rect 3014 3199 3020 3200
rect 3014 3195 3015 3199
rect 3019 3195 3020 3199
rect 3014 3194 3020 3195
rect 3166 3199 3172 3200
rect 3166 3195 3167 3199
rect 3171 3195 3172 3199
rect 3166 3194 3172 3195
rect 3326 3199 3332 3200
rect 3326 3195 3327 3199
rect 3331 3195 3332 3199
rect 3942 3196 3943 3200
rect 3947 3196 3948 3200
rect 3942 3195 3948 3196
rect 3326 3194 3332 3195
rect 111 3190 115 3191
rect 111 3185 115 3186
rect 143 3190 147 3191
rect 143 3185 147 3186
rect 295 3190 299 3191
rect 295 3185 299 3186
rect 431 3190 435 3191
rect 431 3185 435 3186
rect 455 3190 459 3191
rect 455 3185 459 3186
rect 567 3190 571 3191
rect 567 3185 571 3186
rect 623 3190 627 3191
rect 623 3185 627 3186
rect 703 3190 707 3191
rect 703 3185 707 3186
rect 791 3190 795 3191
rect 791 3185 795 3186
rect 855 3190 859 3191
rect 855 3185 859 3186
rect 959 3190 963 3191
rect 959 3185 963 3186
rect 1031 3190 1035 3191
rect 1031 3185 1035 3186
rect 1127 3190 1131 3191
rect 1127 3185 1131 3186
rect 1231 3190 1235 3191
rect 1231 3185 1235 3186
rect 1303 3190 1307 3191
rect 1303 3185 1307 3186
rect 1455 3190 1459 3191
rect 1455 3185 1459 3186
rect 1479 3190 1483 3191
rect 1479 3185 1483 3186
rect 1687 3190 1691 3191
rect 1687 3185 1691 3186
rect 1903 3190 1907 3191
rect 1903 3185 1907 3186
rect 2007 3190 2011 3191
rect 2007 3185 2011 3186
rect 112 3165 114 3185
rect 110 3164 116 3165
rect 296 3164 298 3185
rect 432 3164 434 3185
rect 568 3164 570 3185
rect 704 3164 706 3185
rect 856 3164 858 3185
rect 1032 3164 1034 3185
rect 1232 3164 1234 3185
rect 1456 3164 1458 3185
rect 1688 3164 1690 3185
rect 1904 3164 1906 3185
rect 2008 3165 2010 3185
rect 2046 3183 2052 3184
rect 2046 3179 2047 3183
rect 2051 3179 2052 3183
rect 3942 3183 3948 3184
rect 2046 3178 2052 3179
rect 2070 3180 2076 3181
rect 2006 3164 2012 3165
rect 110 3160 111 3164
rect 115 3160 116 3164
rect 110 3159 116 3160
rect 294 3163 300 3164
rect 294 3159 295 3163
rect 299 3159 300 3163
rect 294 3158 300 3159
rect 430 3163 436 3164
rect 430 3159 431 3163
rect 435 3159 436 3163
rect 430 3158 436 3159
rect 566 3163 572 3164
rect 566 3159 567 3163
rect 571 3159 572 3163
rect 566 3158 572 3159
rect 702 3163 708 3164
rect 702 3159 703 3163
rect 707 3159 708 3163
rect 702 3158 708 3159
rect 854 3163 860 3164
rect 854 3159 855 3163
rect 859 3159 860 3163
rect 854 3158 860 3159
rect 1030 3163 1036 3164
rect 1030 3159 1031 3163
rect 1035 3159 1036 3163
rect 1030 3158 1036 3159
rect 1230 3163 1236 3164
rect 1230 3159 1231 3163
rect 1235 3159 1236 3163
rect 1230 3158 1236 3159
rect 1454 3163 1460 3164
rect 1454 3159 1455 3163
rect 1459 3159 1460 3163
rect 1454 3158 1460 3159
rect 1686 3163 1692 3164
rect 1686 3159 1687 3163
rect 1691 3159 1692 3163
rect 1686 3158 1692 3159
rect 1902 3163 1908 3164
rect 1902 3159 1903 3163
rect 1907 3159 1908 3163
rect 2006 3160 2007 3164
rect 2011 3160 2012 3164
rect 2006 3159 2012 3160
rect 1902 3158 1908 3159
rect 110 3147 116 3148
rect 110 3143 111 3147
rect 115 3143 116 3147
rect 2006 3147 2012 3148
rect 2048 3147 2050 3178
rect 2070 3176 2071 3180
rect 2075 3176 2076 3180
rect 2070 3175 2076 3176
rect 2206 3180 2212 3181
rect 2206 3176 2207 3180
rect 2211 3176 2212 3180
rect 2206 3175 2212 3176
rect 2374 3180 2380 3181
rect 2374 3176 2375 3180
rect 2379 3176 2380 3180
rect 2374 3175 2380 3176
rect 2542 3180 2548 3181
rect 2542 3176 2543 3180
rect 2547 3176 2548 3180
rect 2542 3175 2548 3176
rect 2702 3180 2708 3181
rect 2702 3176 2703 3180
rect 2707 3176 2708 3180
rect 2702 3175 2708 3176
rect 2862 3180 2868 3181
rect 2862 3176 2863 3180
rect 2867 3176 2868 3180
rect 2862 3175 2868 3176
rect 3014 3180 3020 3181
rect 3014 3176 3015 3180
rect 3019 3176 3020 3180
rect 3014 3175 3020 3176
rect 3166 3180 3172 3181
rect 3166 3176 3167 3180
rect 3171 3176 3172 3180
rect 3166 3175 3172 3176
rect 3326 3180 3332 3181
rect 3326 3176 3327 3180
rect 3331 3176 3332 3180
rect 3942 3179 3943 3183
rect 3947 3179 3948 3183
rect 3942 3178 3948 3179
rect 3326 3175 3332 3176
rect 2072 3147 2074 3175
rect 2208 3147 2210 3175
rect 2376 3147 2378 3175
rect 2544 3147 2546 3175
rect 2704 3147 2706 3175
rect 2864 3147 2866 3175
rect 3016 3147 3018 3175
rect 3168 3147 3170 3175
rect 3328 3147 3330 3175
rect 3944 3147 3946 3178
rect 110 3142 116 3143
rect 294 3144 300 3145
rect 112 3115 114 3142
rect 294 3140 295 3144
rect 299 3140 300 3144
rect 294 3139 300 3140
rect 430 3144 436 3145
rect 430 3140 431 3144
rect 435 3140 436 3144
rect 430 3139 436 3140
rect 566 3144 572 3145
rect 566 3140 567 3144
rect 571 3140 572 3144
rect 566 3139 572 3140
rect 702 3144 708 3145
rect 702 3140 703 3144
rect 707 3140 708 3144
rect 702 3139 708 3140
rect 854 3144 860 3145
rect 854 3140 855 3144
rect 859 3140 860 3144
rect 854 3139 860 3140
rect 1030 3144 1036 3145
rect 1030 3140 1031 3144
rect 1035 3140 1036 3144
rect 1030 3139 1036 3140
rect 1230 3144 1236 3145
rect 1230 3140 1231 3144
rect 1235 3140 1236 3144
rect 1230 3139 1236 3140
rect 1454 3144 1460 3145
rect 1454 3140 1455 3144
rect 1459 3140 1460 3144
rect 1454 3139 1460 3140
rect 1686 3144 1692 3145
rect 1686 3140 1687 3144
rect 1691 3140 1692 3144
rect 1686 3139 1692 3140
rect 1902 3144 1908 3145
rect 1902 3140 1903 3144
rect 1907 3140 1908 3144
rect 2006 3143 2007 3147
rect 2011 3143 2012 3147
rect 2006 3142 2012 3143
rect 2047 3146 2051 3147
rect 1902 3139 1908 3140
rect 296 3115 298 3139
rect 432 3115 434 3139
rect 568 3115 570 3139
rect 704 3115 706 3139
rect 856 3115 858 3139
rect 1032 3115 1034 3139
rect 1232 3115 1234 3139
rect 1456 3115 1458 3139
rect 1688 3115 1690 3139
rect 1904 3115 1906 3139
rect 2008 3115 2010 3142
rect 2047 3141 2051 3142
rect 2071 3146 2075 3147
rect 2071 3141 2075 3142
rect 2207 3146 2211 3147
rect 2207 3141 2211 3142
rect 2343 3146 2347 3147
rect 2343 3141 2347 3142
rect 2375 3146 2379 3147
rect 2375 3141 2379 3142
rect 2543 3146 2547 3147
rect 2543 3141 2547 3142
rect 2631 3146 2635 3147
rect 2631 3141 2635 3142
rect 2703 3146 2707 3147
rect 2703 3141 2707 3142
rect 2863 3146 2867 3147
rect 2863 3141 2867 3142
rect 2903 3146 2907 3147
rect 2903 3141 2907 3142
rect 3015 3146 3019 3147
rect 3015 3141 3019 3142
rect 3167 3146 3171 3147
rect 3167 3141 3171 3142
rect 3175 3146 3179 3147
rect 3175 3141 3179 3142
rect 3327 3146 3331 3147
rect 3327 3141 3331 3142
rect 3447 3146 3451 3147
rect 3447 3141 3451 3142
rect 3943 3146 3947 3147
rect 3943 3141 3947 3142
rect 111 3114 115 3115
rect 111 3109 115 3110
rect 295 3114 299 3115
rect 295 3109 299 3110
rect 311 3114 315 3115
rect 311 3109 315 3110
rect 407 3114 411 3115
rect 407 3109 411 3110
rect 431 3114 435 3115
rect 431 3109 435 3110
rect 503 3114 507 3115
rect 503 3109 507 3110
rect 567 3114 571 3115
rect 567 3109 571 3110
rect 599 3114 603 3115
rect 599 3109 603 3110
rect 695 3114 699 3115
rect 695 3109 699 3110
rect 703 3114 707 3115
rect 703 3109 707 3110
rect 807 3114 811 3115
rect 807 3109 811 3110
rect 855 3114 859 3115
rect 855 3109 859 3110
rect 943 3114 947 3115
rect 943 3109 947 3110
rect 1031 3114 1035 3115
rect 1031 3109 1035 3110
rect 1087 3114 1091 3115
rect 1087 3109 1091 3110
rect 1231 3114 1235 3115
rect 1231 3109 1235 3110
rect 1247 3114 1251 3115
rect 1247 3109 1251 3110
rect 1407 3114 1411 3115
rect 1407 3109 1411 3110
rect 1455 3114 1459 3115
rect 1455 3109 1459 3110
rect 1575 3114 1579 3115
rect 1575 3109 1579 3110
rect 1687 3114 1691 3115
rect 1687 3109 1691 3110
rect 1751 3114 1755 3115
rect 1751 3109 1755 3110
rect 1903 3114 1907 3115
rect 1903 3109 1907 3110
rect 2007 3114 2011 3115
rect 2048 3114 2050 3141
rect 2072 3117 2074 3141
rect 2344 3117 2346 3141
rect 2632 3117 2634 3141
rect 2904 3117 2906 3141
rect 3176 3117 3178 3141
rect 3448 3117 3450 3141
rect 2070 3116 2076 3117
rect 2007 3109 2011 3110
rect 2046 3113 2052 3114
rect 2046 3109 2047 3113
rect 2051 3109 2052 3113
rect 2070 3112 2071 3116
rect 2075 3112 2076 3116
rect 2070 3111 2076 3112
rect 2342 3116 2348 3117
rect 2342 3112 2343 3116
rect 2347 3112 2348 3116
rect 2342 3111 2348 3112
rect 2630 3116 2636 3117
rect 2630 3112 2631 3116
rect 2635 3112 2636 3116
rect 2630 3111 2636 3112
rect 2902 3116 2908 3117
rect 2902 3112 2903 3116
rect 2907 3112 2908 3116
rect 2902 3111 2908 3112
rect 3174 3116 3180 3117
rect 3174 3112 3175 3116
rect 3179 3112 3180 3116
rect 3174 3111 3180 3112
rect 3446 3116 3452 3117
rect 3446 3112 3447 3116
rect 3451 3112 3452 3116
rect 3944 3114 3946 3141
rect 3446 3111 3452 3112
rect 3942 3113 3948 3114
rect 112 3082 114 3109
rect 312 3085 314 3109
rect 408 3085 410 3109
rect 504 3085 506 3109
rect 600 3085 602 3109
rect 696 3085 698 3109
rect 808 3085 810 3109
rect 944 3085 946 3109
rect 1088 3085 1090 3109
rect 1248 3085 1250 3109
rect 1408 3085 1410 3109
rect 1576 3085 1578 3109
rect 1752 3085 1754 3109
rect 1904 3085 1906 3109
rect 310 3084 316 3085
rect 110 3081 116 3082
rect 110 3077 111 3081
rect 115 3077 116 3081
rect 310 3080 311 3084
rect 315 3080 316 3084
rect 310 3079 316 3080
rect 406 3084 412 3085
rect 406 3080 407 3084
rect 411 3080 412 3084
rect 406 3079 412 3080
rect 502 3084 508 3085
rect 502 3080 503 3084
rect 507 3080 508 3084
rect 502 3079 508 3080
rect 598 3084 604 3085
rect 598 3080 599 3084
rect 603 3080 604 3084
rect 598 3079 604 3080
rect 694 3084 700 3085
rect 694 3080 695 3084
rect 699 3080 700 3084
rect 694 3079 700 3080
rect 806 3084 812 3085
rect 806 3080 807 3084
rect 811 3080 812 3084
rect 806 3079 812 3080
rect 942 3084 948 3085
rect 942 3080 943 3084
rect 947 3080 948 3084
rect 942 3079 948 3080
rect 1086 3084 1092 3085
rect 1086 3080 1087 3084
rect 1091 3080 1092 3084
rect 1086 3079 1092 3080
rect 1246 3084 1252 3085
rect 1246 3080 1247 3084
rect 1251 3080 1252 3084
rect 1246 3079 1252 3080
rect 1406 3084 1412 3085
rect 1406 3080 1407 3084
rect 1411 3080 1412 3084
rect 1406 3079 1412 3080
rect 1574 3084 1580 3085
rect 1574 3080 1575 3084
rect 1579 3080 1580 3084
rect 1574 3079 1580 3080
rect 1750 3084 1756 3085
rect 1750 3080 1751 3084
rect 1755 3080 1756 3084
rect 1750 3079 1756 3080
rect 1902 3084 1908 3085
rect 1902 3080 1903 3084
rect 1907 3080 1908 3084
rect 2008 3082 2010 3109
rect 2046 3108 2052 3109
rect 3942 3109 3943 3113
rect 3947 3109 3948 3113
rect 3942 3108 3948 3109
rect 2070 3097 2076 3098
rect 2046 3096 2052 3097
rect 2046 3092 2047 3096
rect 2051 3092 2052 3096
rect 2070 3093 2071 3097
rect 2075 3093 2076 3097
rect 2070 3092 2076 3093
rect 2342 3097 2348 3098
rect 2342 3093 2343 3097
rect 2347 3093 2348 3097
rect 2342 3092 2348 3093
rect 2630 3097 2636 3098
rect 2630 3093 2631 3097
rect 2635 3093 2636 3097
rect 2630 3092 2636 3093
rect 2902 3097 2908 3098
rect 2902 3093 2903 3097
rect 2907 3093 2908 3097
rect 2902 3092 2908 3093
rect 3174 3097 3180 3098
rect 3174 3093 3175 3097
rect 3179 3093 3180 3097
rect 3174 3092 3180 3093
rect 3446 3097 3452 3098
rect 3446 3093 3447 3097
rect 3451 3093 3452 3097
rect 3446 3092 3452 3093
rect 3942 3096 3948 3097
rect 3942 3092 3943 3096
rect 3947 3092 3948 3096
rect 2046 3091 2052 3092
rect 1902 3079 1908 3080
rect 2006 3081 2012 3082
rect 110 3076 116 3077
rect 2006 3077 2007 3081
rect 2011 3077 2012 3081
rect 2006 3076 2012 3077
rect 2048 3067 2050 3091
rect 2072 3067 2074 3092
rect 2344 3067 2346 3092
rect 2632 3067 2634 3092
rect 2904 3067 2906 3092
rect 3176 3067 3178 3092
rect 3448 3067 3450 3092
rect 3942 3091 3948 3092
rect 3944 3067 3946 3091
rect 2047 3066 2051 3067
rect 310 3065 316 3066
rect 110 3064 116 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 310 3061 311 3065
rect 315 3061 316 3065
rect 310 3060 316 3061
rect 406 3065 412 3066
rect 406 3061 407 3065
rect 411 3061 412 3065
rect 406 3060 412 3061
rect 502 3065 508 3066
rect 502 3061 503 3065
rect 507 3061 508 3065
rect 502 3060 508 3061
rect 598 3065 604 3066
rect 598 3061 599 3065
rect 603 3061 604 3065
rect 598 3060 604 3061
rect 694 3065 700 3066
rect 694 3061 695 3065
rect 699 3061 700 3065
rect 694 3060 700 3061
rect 806 3065 812 3066
rect 806 3061 807 3065
rect 811 3061 812 3065
rect 806 3060 812 3061
rect 942 3065 948 3066
rect 942 3061 943 3065
rect 947 3061 948 3065
rect 942 3060 948 3061
rect 1086 3065 1092 3066
rect 1086 3061 1087 3065
rect 1091 3061 1092 3065
rect 1086 3060 1092 3061
rect 1246 3065 1252 3066
rect 1246 3061 1247 3065
rect 1251 3061 1252 3065
rect 1246 3060 1252 3061
rect 1406 3065 1412 3066
rect 1406 3061 1407 3065
rect 1411 3061 1412 3065
rect 1406 3060 1412 3061
rect 1574 3065 1580 3066
rect 1574 3061 1575 3065
rect 1579 3061 1580 3065
rect 1574 3060 1580 3061
rect 1750 3065 1756 3066
rect 1750 3061 1751 3065
rect 1755 3061 1756 3065
rect 1750 3060 1756 3061
rect 1902 3065 1908 3066
rect 1902 3061 1903 3065
rect 1907 3061 1908 3065
rect 1902 3060 1908 3061
rect 2006 3064 2012 3065
rect 2006 3060 2007 3064
rect 2011 3060 2012 3064
rect 2047 3061 2051 3062
rect 2071 3066 2075 3067
rect 2071 3061 2075 3062
rect 2343 3066 2347 3067
rect 2343 3061 2347 3062
rect 2487 3066 2491 3067
rect 2487 3061 2491 3062
rect 2615 3066 2619 3067
rect 2615 3061 2619 3062
rect 2631 3066 2635 3067
rect 2631 3061 2635 3062
rect 2743 3066 2747 3067
rect 2743 3061 2747 3062
rect 2863 3066 2867 3067
rect 2863 3061 2867 3062
rect 2903 3066 2907 3067
rect 2903 3061 2907 3062
rect 2983 3066 2987 3067
rect 2983 3061 2987 3062
rect 3103 3066 3107 3067
rect 3103 3061 3107 3062
rect 3175 3066 3179 3067
rect 3175 3061 3179 3062
rect 3215 3066 3219 3067
rect 3215 3061 3219 3062
rect 3327 3066 3331 3067
rect 3327 3061 3331 3062
rect 3431 3066 3435 3067
rect 3431 3061 3435 3062
rect 3447 3066 3451 3067
rect 3447 3061 3451 3062
rect 3535 3066 3539 3067
rect 3535 3061 3539 3062
rect 3639 3066 3643 3067
rect 3639 3061 3643 3062
rect 3743 3066 3747 3067
rect 3743 3061 3747 3062
rect 3839 3066 3843 3067
rect 3839 3061 3843 3062
rect 3943 3066 3947 3067
rect 3943 3061 3947 3062
rect 110 3059 116 3060
rect 112 3039 114 3059
rect 312 3039 314 3060
rect 408 3039 410 3060
rect 504 3039 506 3060
rect 600 3039 602 3060
rect 696 3039 698 3060
rect 808 3039 810 3060
rect 944 3039 946 3060
rect 1088 3039 1090 3060
rect 1248 3039 1250 3060
rect 1408 3039 1410 3060
rect 1576 3039 1578 3060
rect 1752 3039 1754 3060
rect 1904 3039 1906 3060
rect 2006 3059 2012 3060
rect 2008 3039 2010 3059
rect 2048 3041 2050 3061
rect 2046 3040 2052 3041
rect 2488 3040 2490 3061
rect 2616 3040 2618 3061
rect 2744 3040 2746 3061
rect 2864 3040 2866 3061
rect 2984 3040 2986 3061
rect 3104 3040 3106 3061
rect 3216 3040 3218 3061
rect 3328 3040 3330 3061
rect 3432 3040 3434 3061
rect 3536 3040 3538 3061
rect 3640 3040 3642 3061
rect 3744 3040 3746 3061
rect 3840 3040 3842 3061
rect 3944 3041 3946 3061
rect 3942 3040 3948 3041
rect 111 3038 115 3039
rect 111 3033 115 3034
rect 311 3038 315 3039
rect 311 3033 315 3034
rect 407 3038 411 3039
rect 407 3033 411 3034
rect 423 3038 427 3039
rect 423 3033 427 3034
rect 503 3038 507 3039
rect 503 3033 507 3034
rect 519 3038 523 3039
rect 519 3033 523 3034
rect 599 3038 603 3039
rect 599 3033 603 3034
rect 615 3038 619 3039
rect 615 3033 619 3034
rect 695 3038 699 3039
rect 695 3033 699 3034
rect 711 3038 715 3039
rect 711 3033 715 3034
rect 807 3038 811 3039
rect 807 3033 811 3034
rect 815 3038 819 3039
rect 815 3033 819 3034
rect 935 3038 939 3039
rect 935 3033 939 3034
rect 943 3038 947 3039
rect 943 3033 947 3034
rect 1055 3038 1059 3039
rect 1055 3033 1059 3034
rect 1087 3038 1091 3039
rect 1087 3033 1091 3034
rect 1183 3038 1187 3039
rect 1183 3033 1187 3034
rect 1247 3038 1251 3039
rect 1247 3033 1251 3034
rect 1311 3038 1315 3039
rect 1311 3033 1315 3034
rect 1407 3038 1411 3039
rect 1407 3033 1411 3034
rect 1431 3038 1435 3039
rect 1431 3033 1435 3034
rect 1551 3038 1555 3039
rect 1551 3033 1555 3034
rect 1575 3038 1579 3039
rect 1575 3033 1579 3034
rect 1671 3038 1675 3039
rect 1671 3033 1675 3034
rect 1751 3038 1755 3039
rect 1751 3033 1755 3034
rect 1799 3038 1803 3039
rect 1799 3033 1803 3034
rect 1903 3038 1907 3039
rect 1903 3033 1907 3034
rect 2007 3038 2011 3039
rect 2046 3036 2047 3040
rect 2051 3036 2052 3040
rect 2046 3035 2052 3036
rect 2486 3039 2492 3040
rect 2486 3035 2487 3039
rect 2491 3035 2492 3039
rect 2486 3034 2492 3035
rect 2614 3039 2620 3040
rect 2614 3035 2615 3039
rect 2619 3035 2620 3039
rect 2614 3034 2620 3035
rect 2742 3039 2748 3040
rect 2742 3035 2743 3039
rect 2747 3035 2748 3039
rect 2742 3034 2748 3035
rect 2862 3039 2868 3040
rect 2862 3035 2863 3039
rect 2867 3035 2868 3039
rect 2862 3034 2868 3035
rect 2982 3039 2988 3040
rect 2982 3035 2983 3039
rect 2987 3035 2988 3039
rect 2982 3034 2988 3035
rect 3102 3039 3108 3040
rect 3102 3035 3103 3039
rect 3107 3035 3108 3039
rect 3102 3034 3108 3035
rect 3214 3039 3220 3040
rect 3214 3035 3215 3039
rect 3219 3035 3220 3039
rect 3214 3034 3220 3035
rect 3326 3039 3332 3040
rect 3326 3035 3327 3039
rect 3331 3035 3332 3039
rect 3326 3034 3332 3035
rect 3430 3039 3436 3040
rect 3430 3035 3431 3039
rect 3435 3035 3436 3039
rect 3430 3034 3436 3035
rect 3534 3039 3540 3040
rect 3534 3035 3535 3039
rect 3539 3035 3540 3039
rect 3534 3034 3540 3035
rect 3638 3039 3644 3040
rect 3638 3035 3639 3039
rect 3643 3035 3644 3039
rect 3638 3034 3644 3035
rect 3742 3039 3748 3040
rect 3742 3035 3743 3039
rect 3747 3035 3748 3039
rect 3742 3034 3748 3035
rect 3838 3039 3844 3040
rect 3838 3035 3839 3039
rect 3843 3035 3844 3039
rect 3942 3036 3943 3040
rect 3947 3036 3948 3040
rect 3942 3035 3948 3036
rect 3838 3034 3844 3035
rect 2007 3033 2011 3034
rect 112 3013 114 3033
rect 110 3012 116 3013
rect 424 3012 426 3033
rect 520 3012 522 3033
rect 616 3012 618 3033
rect 712 3012 714 3033
rect 816 3012 818 3033
rect 936 3012 938 3033
rect 1056 3012 1058 3033
rect 1184 3012 1186 3033
rect 1312 3012 1314 3033
rect 1432 3012 1434 3033
rect 1552 3012 1554 3033
rect 1672 3012 1674 3033
rect 1800 3012 1802 3033
rect 1904 3012 1906 3033
rect 2008 3013 2010 3033
rect 2046 3023 2052 3024
rect 2046 3019 2047 3023
rect 2051 3019 2052 3023
rect 3942 3023 3948 3024
rect 2046 3018 2052 3019
rect 2486 3020 2492 3021
rect 2006 3012 2012 3013
rect 110 3008 111 3012
rect 115 3008 116 3012
rect 110 3007 116 3008
rect 422 3011 428 3012
rect 422 3007 423 3011
rect 427 3007 428 3011
rect 422 3006 428 3007
rect 518 3011 524 3012
rect 518 3007 519 3011
rect 523 3007 524 3011
rect 518 3006 524 3007
rect 614 3011 620 3012
rect 614 3007 615 3011
rect 619 3007 620 3011
rect 614 3006 620 3007
rect 710 3011 716 3012
rect 710 3007 711 3011
rect 715 3007 716 3011
rect 710 3006 716 3007
rect 814 3011 820 3012
rect 814 3007 815 3011
rect 819 3007 820 3011
rect 814 3006 820 3007
rect 934 3011 940 3012
rect 934 3007 935 3011
rect 939 3007 940 3011
rect 934 3006 940 3007
rect 1054 3011 1060 3012
rect 1054 3007 1055 3011
rect 1059 3007 1060 3011
rect 1054 3006 1060 3007
rect 1182 3011 1188 3012
rect 1182 3007 1183 3011
rect 1187 3007 1188 3011
rect 1182 3006 1188 3007
rect 1310 3011 1316 3012
rect 1310 3007 1311 3011
rect 1315 3007 1316 3011
rect 1310 3006 1316 3007
rect 1430 3011 1436 3012
rect 1430 3007 1431 3011
rect 1435 3007 1436 3011
rect 1430 3006 1436 3007
rect 1550 3011 1556 3012
rect 1550 3007 1551 3011
rect 1555 3007 1556 3011
rect 1550 3006 1556 3007
rect 1670 3011 1676 3012
rect 1670 3007 1671 3011
rect 1675 3007 1676 3011
rect 1670 3006 1676 3007
rect 1798 3011 1804 3012
rect 1798 3007 1799 3011
rect 1803 3007 1804 3011
rect 1798 3006 1804 3007
rect 1902 3011 1908 3012
rect 1902 3007 1903 3011
rect 1907 3007 1908 3011
rect 2006 3008 2007 3012
rect 2011 3008 2012 3012
rect 2006 3007 2012 3008
rect 1902 3006 1908 3007
rect 110 2995 116 2996
rect 110 2991 111 2995
rect 115 2991 116 2995
rect 2006 2995 2012 2996
rect 110 2990 116 2991
rect 422 2992 428 2993
rect 112 2939 114 2990
rect 422 2988 423 2992
rect 427 2988 428 2992
rect 422 2987 428 2988
rect 518 2992 524 2993
rect 518 2988 519 2992
rect 523 2988 524 2992
rect 518 2987 524 2988
rect 614 2992 620 2993
rect 614 2988 615 2992
rect 619 2988 620 2992
rect 614 2987 620 2988
rect 710 2992 716 2993
rect 710 2988 711 2992
rect 715 2988 716 2992
rect 710 2987 716 2988
rect 814 2992 820 2993
rect 814 2988 815 2992
rect 819 2988 820 2992
rect 814 2987 820 2988
rect 934 2992 940 2993
rect 934 2988 935 2992
rect 939 2988 940 2992
rect 934 2987 940 2988
rect 1054 2992 1060 2993
rect 1054 2988 1055 2992
rect 1059 2988 1060 2992
rect 1054 2987 1060 2988
rect 1182 2992 1188 2993
rect 1182 2988 1183 2992
rect 1187 2988 1188 2992
rect 1182 2987 1188 2988
rect 1310 2992 1316 2993
rect 1310 2988 1311 2992
rect 1315 2988 1316 2992
rect 1310 2987 1316 2988
rect 1430 2992 1436 2993
rect 1430 2988 1431 2992
rect 1435 2988 1436 2992
rect 1430 2987 1436 2988
rect 1550 2992 1556 2993
rect 1550 2988 1551 2992
rect 1555 2988 1556 2992
rect 1550 2987 1556 2988
rect 1670 2992 1676 2993
rect 1670 2988 1671 2992
rect 1675 2988 1676 2992
rect 1670 2987 1676 2988
rect 1798 2992 1804 2993
rect 1798 2988 1799 2992
rect 1803 2988 1804 2992
rect 1798 2987 1804 2988
rect 1902 2992 1908 2993
rect 1902 2988 1903 2992
rect 1907 2988 1908 2992
rect 2006 2991 2007 2995
rect 2011 2991 2012 2995
rect 2006 2990 2012 2991
rect 1902 2987 1908 2988
rect 424 2939 426 2987
rect 520 2939 522 2987
rect 616 2939 618 2987
rect 712 2939 714 2987
rect 816 2939 818 2987
rect 936 2939 938 2987
rect 1056 2939 1058 2987
rect 1184 2939 1186 2987
rect 1312 2939 1314 2987
rect 1432 2939 1434 2987
rect 1552 2939 1554 2987
rect 1672 2939 1674 2987
rect 1800 2939 1802 2987
rect 1904 2939 1906 2987
rect 2008 2939 2010 2990
rect 2048 2987 2050 3018
rect 2486 3016 2487 3020
rect 2491 3016 2492 3020
rect 2486 3015 2492 3016
rect 2614 3020 2620 3021
rect 2614 3016 2615 3020
rect 2619 3016 2620 3020
rect 2614 3015 2620 3016
rect 2742 3020 2748 3021
rect 2742 3016 2743 3020
rect 2747 3016 2748 3020
rect 2742 3015 2748 3016
rect 2862 3020 2868 3021
rect 2862 3016 2863 3020
rect 2867 3016 2868 3020
rect 2862 3015 2868 3016
rect 2982 3020 2988 3021
rect 2982 3016 2983 3020
rect 2987 3016 2988 3020
rect 2982 3015 2988 3016
rect 3102 3020 3108 3021
rect 3102 3016 3103 3020
rect 3107 3016 3108 3020
rect 3102 3015 3108 3016
rect 3214 3020 3220 3021
rect 3214 3016 3215 3020
rect 3219 3016 3220 3020
rect 3214 3015 3220 3016
rect 3326 3020 3332 3021
rect 3326 3016 3327 3020
rect 3331 3016 3332 3020
rect 3326 3015 3332 3016
rect 3430 3020 3436 3021
rect 3430 3016 3431 3020
rect 3435 3016 3436 3020
rect 3430 3015 3436 3016
rect 3534 3020 3540 3021
rect 3534 3016 3535 3020
rect 3539 3016 3540 3020
rect 3534 3015 3540 3016
rect 3638 3020 3644 3021
rect 3638 3016 3639 3020
rect 3643 3016 3644 3020
rect 3638 3015 3644 3016
rect 3742 3020 3748 3021
rect 3742 3016 3743 3020
rect 3747 3016 3748 3020
rect 3742 3015 3748 3016
rect 3838 3020 3844 3021
rect 3838 3016 3839 3020
rect 3843 3016 3844 3020
rect 3942 3019 3943 3023
rect 3947 3019 3948 3023
rect 3942 3018 3948 3019
rect 3838 3015 3844 3016
rect 2488 2987 2490 3015
rect 2616 2987 2618 3015
rect 2744 2987 2746 3015
rect 2864 2987 2866 3015
rect 2984 2987 2986 3015
rect 3104 2987 3106 3015
rect 3216 2987 3218 3015
rect 3328 2987 3330 3015
rect 3432 2987 3434 3015
rect 3536 2987 3538 3015
rect 3640 2987 3642 3015
rect 3744 2987 3746 3015
rect 3840 2987 3842 3015
rect 3944 2987 3946 3018
rect 2047 2986 2051 2987
rect 2047 2981 2051 2982
rect 2407 2986 2411 2987
rect 2407 2981 2411 2982
rect 2487 2986 2491 2987
rect 2487 2981 2491 2982
rect 2575 2986 2579 2987
rect 2575 2981 2579 2982
rect 2615 2986 2619 2987
rect 2615 2981 2619 2982
rect 2743 2986 2747 2987
rect 2743 2981 2747 2982
rect 2767 2986 2771 2987
rect 2767 2981 2771 2982
rect 2863 2986 2867 2987
rect 2863 2981 2867 2982
rect 2967 2986 2971 2987
rect 2967 2981 2971 2982
rect 2983 2986 2987 2987
rect 2983 2981 2987 2982
rect 3103 2986 3107 2987
rect 3103 2981 3107 2982
rect 3183 2986 3187 2987
rect 3183 2981 3187 2982
rect 3215 2986 3219 2987
rect 3215 2981 3219 2982
rect 3327 2986 3331 2987
rect 3327 2981 3331 2982
rect 3399 2986 3403 2987
rect 3399 2981 3403 2982
rect 3431 2986 3435 2987
rect 3431 2981 3435 2982
rect 3535 2986 3539 2987
rect 3535 2981 3539 2982
rect 3623 2986 3627 2987
rect 3623 2981 3627 2982
rect 3639 2986 3643 2987
rect 3639 2981 3643 2982
rect 3743 2986 3747 2987
rect 3743 2981 3747 2982
rect 3839 2986 3843 2987
rect 3839 2981 3843 2982
rect 3943 2986 3947 2987
rect 3943 2981 3947 2982
rect 2048 2954 2050 2981
rect 2408 2957 2410 2981
rect 2576 2957 2578 2981
rect 2768 2957 2770 2981
rect 2968 2957 2970 2981
rect 3184 2957 3186 2981
rect 3400 2957 3402 2981
rect 3624 2957 3626 2981
rect 3840 2957 3842 2981
rect 2406 2956 2412 2957
rect 2046 2953 2052 2954
rect 2046 2949 2047 2953
rect 2051 2949 2052 2953
rect 2406 2952 2407 2956
rect 2411 2952 2412 2956
rect 2406 2951 2412 2952
rect 2574 2956 2580 2957
rect 2574 2952 2575 2956
rect 2579 2952 2580 2956
rect 2574 2951 2580 2952
rect 2766 2956 2772 2957
rect 2766 2952 2767 2956
rect 2771 2952 2772 2956
rect 2766 2951 2772 2952
rect 2966 2956 2972 2957
rect 2966 2952 2967 2956
rect 2971 2952 2972 2956
rect 2966 2951 2972 2952
rect 3182 2956 3188 2957
rect 3182 2952 3183 2956
rect 3187 2952 3188 2956
rect 3182 2951 3188 2952
rect 3398 2956 3404 2957
rect 3398 2952 3399 2956
rect 3403 2952 3404 2956
rect 3398 2951 3404 2952
rect 3622 2956 3628 2957
rect 3622 2952 3623 2956
rect 3627 2952 3628 2956
rect 3622 2951 3628 2952
rect 3838 2956 3844 2957
rect 3838 2952 3839 2956
rect 3843 2952 3844 2956
rect 3944 2954 3946 2981
rect 3838 2951 3844 2952
rect 3942 2953 3948 2954
rect 2046 2948 2052 2949
rect 3942 2949 3943 2953
rect 3947 2949 3948 2953
rect 3942 2948 3948 2949
rect 111 2938 115 2939
rect 111 2933 115 2934
rect 423 2938 427 2939
rect 423 2933 427 2934
rect 519 2938 523 2939
rect 519 2933 523 2934
rect 615 2938 619 2939
rect 615 2933 619 2934
rect 711 2938 715 2939
rect 711 2933 715 2934
rect 815 2938 819 2939
rect 815 2933 819 2934
rect 935 2938 939 2939
rect 935 2933 939 2934
rect 1055 2938 1059 2939
rect 1055 2933 1059 2934
rect 1183 2938 1187 2939
rect 1183 2933 1187 2934
rect 1311 2938 1315 2939
rect 1311 2933 1315 2934
rect 1431 2938 1435 2939
rect 1431 2933 1435 2934
rect 1479 2938 1483 2939
rect 1479 2933 1483 2934
rect 1551 2938 1555 2939
rect 1551 2933 1555 2934
rect 1575 2938 1579 2939
rect 1575 2933 1579 2934
rect 1671 2938 1675 2939
rect 1671 2933 1675 2934
rect 1767 2938 1771 2939
rect 1767 2933 1771 2934
rect 1799 2938 1803 2939
rect 1799 2933 1803 2934
rect 1863 2938 1867 2939
rect 1863 2933 1867 2934
rect 1903 2938 1907 2939
rect 1903 2933 1907 2934
rect 2007 2938 2011 2939
rect 2406 2937 2412 2938
rect 2007 2933 2011 2934
rect 2046 2936 2052 2937
rect 112 2906 114 2933
rect 1480 2909 1482 2933
rect 1576 2909 1578 2933
rect 1672 2909 1674 2933
rect 1768 2909 1770 2933
rect 1864 2909 1866 2933
rect 1478 2908 1484 2909
rect 110 2905 116 2906
rect 110 2901 111 2905
rect 115 2901 116 2905
rect 1478 2904 1479 2908
rect 1483 2904 1484 2908
rect 1478 2903 1484 2904
rect 1574 2908 1580 2909
rect 1574 2904 1575 2908
rect 1579 2904 1580 2908
rect 1574 2903 1580 2904
rect 1670 2908 1676 2909
rect 1670 2904 1671 2908
rect 1675 2904 1676 2908
rect 1670 2903 1676 2904
rect 1766 2908 1772 2909
rect 1766 2904 1767 2908
rect 1771 2904 1772 2908
rect 1766 2903 1772 2904
rect 1862 2908 1868 2909
rect 1862 2904 1863 2908
rect 1867 2904 1868 2908
rect 2008 2906 2010 2933
rect 2046 2932 2047 2936
rect 2051 2932 2052 2936
rect 2406 2933 2407 2937
rect 2411 2933 2412 2937
rect 2406 2932 2412 2933
rect 2574 2937 2580 2938
rect 2574 2933 2575 2937
rect 2579 2933 2580 2937
rect 2574 2932 2580 2933
rect 2766 2937 2772 2938
rect 2766 2933 2767 2937
rect 2771 2933 2772 2937
rect 2766 2932 2772 2933
rect 2966 2937 2972 2938
rect 2966 2933 2967 2937
rect 2971 2933 2972 2937
rect 2966 2932 2972 2933
rect 3182 2937 3188 2938
rect 3182 2933 3183 2937
rect 3187 2933 3188 2937
rect 3182 2932 3188 2933
rect 3398 2937 3404 2938
rect 3398 2933 3399 2937
rect 3403 2933 3404 2937
rect 3398 2932 3404 2933
rect 3622 2937 3628 2938
rect 3622 2933 3623 2937
rect 3627 2933 3628 2937
rect 3622 2932 3628 2933
rect 3838 2937 3844 2938
rect 3838 2933 3839 2937
rect 3843 2933 3844 2937
rect 3838 2932 3844 2933
rect 3942 2936 3948 2937
rect 3942 2932 3943 2936
rect 3947 2932 3948 2936
rect 2046 2931 2052 2932
rect 1862 2903 1868 2904
rect 2006 2905 2012 2906
rect 110 2900 116 2901
rect 2006 2901 2007 2905
rect 2011 2901 2012 2905
rect 2006 2900 2012 2901
rect 2048 2895 2050 2931
rect 2408 2895 2410 2932
rect 2576 2895 2578 2932
rect 2768 2895 2770 2932
rect 2968 2895 2970 2932
rect 3184 2895 3186 2932
rect 3400 2895 3402 2932
rect 3624 2895 3626 2932
rect 3840 2895 3842 2932
rect 3942 2931 3948 2932
rect 3944 2895 3946 2931
rect 2047 2894 2051 2895
rect 1478 2889 1484 2890
rect 110 2888 116 2889
rect 110 2884 111 2888
rect 115 2884 116 2888
rect 1478 2885 1479 2889
rect 1483 2885 1484 2889
rect 1478 2884 1484 2885
rect 1574 2889 1580 2890
rect 1574 2885 1575 2889
rect 1579 2885 1580 2889
rect 1574 2884 1580 2885
rect 1670 2889 1676 2890
rect 1670 2885 1671 2889
rect 1675 2885 1676 2889
rect 1670 2884 1676 2885
rect 1766 2889 1772 2890
rect 1766 2885 1767 2889
rect 1771 2885 1772 2889
rect 1766 2884 1772 2885
rect 1862 2889 1868 2890
rect 2047 2889 2051 2890
rect 2407 2894 2411 2895
rect 2407 2889 2411 2890
rect 2551 2894 2555 2895
rect 2551 2889 2555 2890
rect 2575 2894 2579 2895
rect 2575 2889 2579 2890
rect 2671 2894 2675 2895
rect 2671 2889 2675 2890
rect 2767 2894 2771 2895
rect 2767 2889 2771 2890
rect 2799 2894 2803 2895
rect 2799 2889 2803 2890
rect 2927 2894 2931 2895
rect 2927 2889 2931 2890
rect 2967 2894 2971 2895
rect 2967 2889 2971 2890
rect 3055 2894 3059 2895
rect 3055 2889 3059 2890
rect 3183 2894 3187 2895
rect 3183 2889 3187 2890
rect 3311 2894 3315 2895
rect 3311 2889 3315 2890
rect 3399 2894 3403 2895
rect 3399 2889 3403 2890
rect 3439 2894 3443 2895
rect 3439 2889 3443 2890
rect 3575 2894 3579 2895
rect 3575 2889 3579 2890
rect 3623 2894 3627 2895
rect 3623 2889 3627 2890
rect 3839 2894 3843 2895
rect 3839 2889 3843 2890
rect 3943 2894 3947 2895
rect 3943 2889 3947 2890
rect 1862 2885 1863 2889
rect 1867 2885 1868 2889
rect 1862 2884 1868 2885
rect 2006 2888 2012 2889
rect 2006 2884 2007 2888
rect 2011 2884 2012 2888
rect 110 2883 116 2884
rect 112 2855 114 2883
rect 1480 2855 1482 2884
rect 1576 2855 1578 2884
rect 1672 2855 1674 2884
rect 1768 2855 1770 2884
rect 1864 2855 1866 2884
rect 2006 2883 2012 2884
rect 2008 2855 2010 2883
rect 2048 2869 2050 2889
rect 2046 2868 2052 2869
rect 2552 2868 2554 2889
rect 2672 2868 2674 2889
rect 2800 2868 2802 2889
rect 2928 2868 2930 2889
rect 3056 2868 3058 2889
rect 3184 2868 3186 2889
rect 3312 2868 3314 2889
rect 3440 2868 3442 2889
rect 3576 2868 3578 2889
rect 3944 2869 3946 2889
rect 3942 2868 3948 2869
rect 2046 2864 2047 2868
rect 2051 2864 2052 2868
rect 2046 2863 2052 2864
rect 2550 2867 2556 2868
rect 2550 2863 2551 2867
rect 2555 2863 2556 2867
rect 2550 2862 2556 2863
rect 2670 2867 2676 2868
rect 2670 2863 2671 2867
rect 2675 2863 2676 2867
rect 2670 2862 2676 2863
rect 2798 2867 2804 2868
rect 2798 2863 2799 2867
rect 2803 2863 2804 2867
rect 2798 2862 2804 2863
rect 2926 2867 2932 2868
rect 2926 2863 2927 2867
rect 2931 2863 2932 2867
rect 2926 2862 2932 2863
rect 3054 2867 3060 2868
rect 3054 2863 3055 2867
rect 3059 2863 3060 2867
rect 3054 2862 3060 2863
rect 3182 2867 3188 2868
rect 3182 2863 3183 2867
rect 3187 2863 3188 2867
rect 3182 2862 3188 2863
rect 3310 2867 3316 2868
rect 3310 2863 3311 2867
rect 3315 2863 3316 2867
rect 3310 2862 3316 2863
rect 3438 2867 3444 2868
rect 3438 2863 3439 2867
rect 3443 2863 3444 2867
rect 3438 2862 3444 2863
rect 3574 2867 3580 2868
rect 3574 2863 3575 2867
rect 3579 2863 3580 2867
rect 3942 2864 3943 2868
rect 3947 2864 3948 2868
rect 3942 2863 3948 2864
rect 3574 2862 3580 2863
rect 111 2854 115 2855
rect 111 2849 115 2850
rect 279 2854 283 2855
rect 279 2849 283 2850
rect 447 2854 451 2855
rect 447 2849 451 2850
rect 631 2854 635 2855
rect 631 2849 635 2850
rect 815 2854 819 2855
rect 815 2849 819 2850
rect 999 2854 1003 2855
rect 999 2849 1003 2850
rect 1183 2854 1187 2855
rect 1183 2849 1187 2850
rect 1359 2854 1363 2855
rect 1359 2849 1363 2850
rect 1479 2854 1483 2855
rect 1479 2849 1483 2850
rect 1527 2854 1531 2855
rect 1527 2849 1531 2850
rect 1575 2854 1579 2855
rect 1575 2849 1579 2850
rect 1671 2854 1675 2855
rect 1671 2849 1675 2850
rect 1695 2854 1699 2855
rect 1695 2849 1699 2850
rect 1767 2854 1771 2855
rect 1767 2849 1771 2850
rect 1863 2854 1867 2855
rect 1863 2849 1867 2850
rect 2007 2854 2011 2855
rect 2007 2849 2011 2850
rect 2046 2851 2052 2852
rect 112 2829 114 2849
rect 110 2828 116 2829
rect 280 2828 282 2849
rect 448 2828 450 2849
rect 632 2828 634 2849
rect 816 2828 818 2849
rect 1000 2828 1002 2849
rect 1184 2828 1186 2849
rect 1360 2828 1362 2849
rect 1528 2828 1530 2849
rect 1696 2828 1698 2849
rect 1864 2828 1866 2849
rect 2008 2829 2010 2849
rect 2046 2847 2047 2851
rect 2051 2847 2052 2851
rect 3942 2851 3948 2852
rect 2046 2846 2052 2847
rect 2550 2848 2556 2849
rect 2006 2828 2012 2829
rect 110 2824 111 2828
rect 115 2824 116 2828
rect 110 2823 116 2824
rect 278 2827 284 2828
rect 278 2823 279 2827
rect 283 2823 284 2827
rect 278 2822 284 2823
rect 446 2827 452 2828
rect 446 2823 447 2827
rect 451 2823 452 2827
rect 446 2822 452 2823
rect 630 2827 636 2828
rect 630 2823 631 2827
rect 635 2823 636 2827
rect 630 2822 636 2823
rect 814 2827 820 2828
rect 814 2823 815 2827
rect 819 2823 820 2827
rect 814 2822 820 2823
rect 998 2827 1004 2828
rect 998 2823 999 2827
rect 1003 2823 1004 2827
rect 998 2822 1004 2823
rect 1182 2827 1188 2828
rect 1182 2823 1183 2827
rect 1187 2823 1188 2827
rect 1182 2822 1188 2823
rect 1358 2827 1364 2828
rect 1358 2823 1359 2827
rect 1363 2823 1364 2827
rect 1358 2822 1364 2823
rect 1526 2827 1532 2828
rect 1526 2823 1527 2827
rect 1531 2823 1532 2827
rect 1526 2822 1532 2823
rect 1694 2827 1700 2828
rect 1694 2823 1695 2827
rect 1699 2823 1700 2827
rect 1694 2822 1700 2823
rect 1862 2827 1868 2828
rect 1862 2823 1863 2827
rect 1867 2823 1868 2827
rect 2006 2824 2007 2828
rect 2011 2824 2012 2828
rect 2006 2823 2012 2824
rect 1862 2822 1868 2823
rect 2048 2819 2050 2846
rect 2550 2844 2551 2848
rect 2555 2844 2556 2848
rect 2550 2843 2556 2844
rect 2670 2848 2676 2849
rect 2670 2844 2671 2848
rect 2675 2844 2676 2848
rect 2670 2843 2676 2844
rect 2798 2848 2804 2849
rect 2798 2844 2799 2848
rect 2803 2844 2804 2848
rect 2798 2843 2804 2844
rect 2926 2848 2932 2849
rect 2926 2844 2927 2848
rect 2931 2844 2932 2848
rect 2926 2843 2932 2844
rect 3054 2848 3060 2849
rect 3054 2844 3055 2848
rect 3059 2844 3060 2848
rect 3054 2843 3060 2844
rect 3182 2848 3188 2849
rect 3182 2844 3183 2848
rect 3187 2844 3188 2848
rect 3182 2843 3188 2844
rect 3310 2848 3316 2849
rect 3310 2844 3311 2848
rect 3315 2844 3316 2848
rect 3310 2843 3316 2844
rect 3438 2848 3444 2849
rect 3438 2844 3439 2848
rect 3443 2844 3444 2848
rect 3438 2843 3444 2844
rect 3574 2848 3580 2849
rect 3574 2844 3575 2848
rect 3579 2844 3580 2848
rect 3942 2847 3943 2851
rect 3947 2847 3948 2851
rect 3942 2846 3948 2847
rect 3574 2843 3580 2844
rect 2552 2819 2554 2843
rect 2672 2819 2674 2843
rect 2800 2819 2802 2843
rect 2928 2819 2930 2843
rect 3056 2819 3058 2843
rect 3184 2819 3186 2843
rect 3312 2819 3314 2843
rect 3440 2819 3442 2843
rect 3576 2819 3578 2843
rect 3944 2819 3946 2846
rect 2047 2818 2051 2819
rect 2047 2813 2051 2814
rect 2439 2818 2443 2819
rect 2439 2813 2443 2814
rect 2551 2818 2555 2819
rect 2551 2813 2555 2814
rect 2567 2818 2571 2819
rect 2567 2813 2571 2814
rect 2671 2818 2675 2819
rect 2671 2813 2675 2814
rect 2695 2818 2699 2819
rect 2695 2813 2699 2814
rect 2799 2818 2803 2819
rect 2799 2813 2803 2814
rect 2831 2818 2835 2819
rect 2831 2813 2835 2814
rect 2927 2818 2931 2819
rect 2927 2813 2931 2814
rect 2967 2818 2971 2819
rect 2967 2813 2971 2814
rect 3055 2818 3059 2819
rect 3055 2813 3059 2814
rect 3103 2818 3107 2819
rect 3103 2813 3107 2814
rect 3183 2818 3187 2819
rect 3183 2813 3187 2814
rect 3247 2818 3251 2819
rect 3247 2813 3251 2814
rect 3311 2818 3315 2819
rect 3311 2813 3315 2814
rect 3391 2818 3395 2819
rect 3391 2813 3395 2814
rect 3439 2818 3443 2819
rect 3439 2813 3443 2814
rect 3543 2818 3547 2819
rect 3543 2813 3547 2814
rect 3575 2818 3579 2819
rect 3575 2813 3579 2814
rect 3703 2818 3707 2819
rect 3703 2813 3707 2814
rect 3839 2818 3843 2819
rect 3839 2813 3843 2814
rect 3943 2818 3947 2819
rect 3943 2813 3947 2814
rect 110 2811 116 2812
rect 110 2807 111 2811
rect 115 2807 116 2811
rect 2006 2811 2012 2812
rect 110 2806 116 2807
rect 278 2808 284 2809
rect 112 2779 114 2806
rect 278 2804 279 2808
rect 283 2804 284 2808
rect 278 2803 284 2804
rect 446 2808 452 2809
rect 446 2804 447 2808
rect 451 2804 452 2808
rect 446 2803 452 2804
rect 630 2808 636 2809
rect 630 2804 631 2808
rect 635 2804 636 2808
rect 630 2803 636 2804
rect 814 2808 820 2809
rect 814 2804 815 2808
rect 819 2804 820 2808
rect 814 2803 820 2804
rect 998 2808 1004 2809
rect 998 2804 999 2808
rect 1003 2804 1004 2808
rect 998 2803 1004 2804
rect 1182 2808 1188 2809
rect 1182 2804 1183 2808
rect 1187 2804 1188 2808
rect 1182 2803 1188 2804
rect 1358 2808 1364 2809
rect 1358 2804 1359 2808
rect 1363 2804 1364 2808
rect 1358 2803 1364 2804
rect 1526 2808 1532 2809
rect 1526 2804 1527 2808
rect 1531 2804 1532 2808
rect 1526 2803 1532 2804
rect 1694 2808 1700 2809
rect 1694 2804 1695 2808
rect 1699 2804 1700 2808
rect 1694 2803 1700 2804
rect 1862 2808 1868 2809
rect 1862 2804 1863 2808
rect 1867 2804 1868 2808
rect 2006 2807 2007 2811
rect 2011 2807 2012 2811
rect 2006 2806 2012 2807
rect 1862 2803 1868 2804
rect 280 2779 282 2803
rect 448 2779 450 2803
rect 632 2779 634 2803
rect 816 2779 818 2803
rect 1000 2779 1002 2803
rect 1184 2779 1186 2803
rect 1360 2779 1362 2803
rect 1528 2779 1530 2803
rect 1696 2779 1698 2803
rect 1864 2779 1866 2803
rect 2008 2779 2010 2806
rect 2048 2786 2050 2813
rect 2440 2789 2442 2813
rect 2568 2789 2570 2813
rect 2696 2789 2698 2813
rect 2832 2789 2834 2813
rect 2968 2789 2970 2813
rect 3104 2789 3106 2813
rect 3248 2789 3250 2813
rect 3392 2789 3394 2813
rect 3544 2789 3546 2813
rect 3704 2789 3706 2813
rect 3840 2789 3842 2813
rect 2438 2788 2444 2789
rect 2046 2785 2052 2786
rect 2046 2781 2047 2785
rect 2051 2781 2052 2785
rect 2438 2784 2439 2788
rect 2443 2784 2444 2788
rect 2438 2783 2444 2784
rect 2566 2788 2572 2789
rect 2566 2784 2567 2788
rect 2571 2784 2572 2788
rect 2566 2783 2572 2784
rect 2694 2788 2700 2789
rect 2694 2784 2695 2788
rect 2699 2784 2700 2788
rect 2694 2783 2700 2784
rect 2830 2788 2836 2789
rect 2830 2784 2831 2788
rect 2835 2784 2836 2788
rect 2830 2783 2836 2784
rect 2966 2788 2972 2789
rect 2966 2784 2967 2788
rect 2971 2784 2972 2788
rect 2966 2783 2972 2784
rect 3102 2788 3108 2789
rect 3102 2784 3103 2788
rect 3107 2784 3108 2788
rect 3102 2783 3108 2784
rect 3246 2788 3252 2789
rect 3246 2784 3247 2788
rect 3251 2784 3252 2788
rect 3246 2783 3252 2784
rect 3390 2788 3396 2789
rect 3390 2784 3391 2788
rect 3395 2784 3396 2788
rect 3390 2783 3396 2784
rect 3542 2788 3548 2789
rect 3542 2784 3543 2788
rect 3547 2784 3548 2788
rect 3542 2783 3548 2784
rect 3702 2788 3708 2789
rect 3702 2784 3703 2788
rect 3707 2784 3708 2788
rect 3702 2783 3708 2784
rect 3838 2788 3844 2789
rect 3838 2784 3839 2788
rect 3843 2784 3844 2788
rect 3944 2786 3946 2813
rect 3838 2783 3844 2784
rect 3942 2785 3948 2786
rect 2046 2780 2052 2781
rect 3942 2781 3943 2785
rect 3947 2781 3948 2785
rect 3942 2780 3948 2781
rect 111 2778 115 2779
rect 111 2773 115 2774
rect 239 2778 243 2779
rect 239 2773 243 2774
rect 279 2778 283 2779
rect 279 2773 283 2774
rect 351 2778 355 2779
rect 351 2773 355 2774
rect 447 2778 451 2779
rect 447 2773 451 2774
rect 471 2778 475 2779
rect 471 2773 475 2774
rect 607 2778 611 2779
rect 607 2773 611 2774
rect 631 2778 635 2779
rect 631 2773 635 2774
rect 743 2778 747 2779
rect 743 2773 747 2774
rect 815 2778 819 2779
rect 815 2773 819 2774
rect 879 2778 883 2779
rect 879 2773 883 2774
rect 999 2778 1003 2779
rect 999 2773 1003 2774
rect 1015 2778 1019 2779
rect 1015 2773 1019 2774
rect 1151 2778 1155 2779
rect 1151 2773 1155 2774
rect 1183 2778 1187 2779
rect 1183 2773 1187 2774
rect 1287 2778 1291 2779
rect 1287 2773 1291 2774
rect 1359 2778 1363 2779
rect 1359 2773 1363 2774
rect 1423 2778 1427 2779
rect 1423 2773 1427 2774
rect 1527 2778 1531 2779
rect 1527 2773 1531 2774
rect 1567 2778 1571 2779
rect 1567 2773 1571 2774
rect 1695 2778 1699 2779
rect 1695 2773 1699 2774
rect 1863 2778 1867 2779
rect 1863 2773 1867 2774
rect 2007 2778 2011 2779
rect 2007 2773 2011 2774
rect 112 2746 114 2773
rect 240 2749 242 2773
rect 352 2749 354 2773
rect 472 2749 474 2773
rect 608 2749 610 2773
rect 744 2749 746 2773
rect 880 2749 882 2773
rect 1016 2749 1018 2773
rect 1152 2749 1154 2773
rect 1288 2749 1290 2773
rect 1424 2749 1426 2773
rect 1568 2749 1570 2773
rect 238 2748 244 2749
rect 110 2745 116 2746
rect 110 2741 111 2745
rect 115 2741 116 2745
rect 238 2744 239 2748
rect 243 2744 244 2748
rect 238 2743 244 2744
rect 350 2748 356 2749
rect 350 2744 351 2748
rect 355 2744 356 2748
rect 350 2743 356 2744
rect 470 2748 476 2749
rect 470 2744 471 2748
rect 475 2744 476 2748
rect 470 2743 476 2744
rect 606 2748 612 2749
rect 606 2744 607 2748
rect 611 2744 612 2748
rect 606 2743 612 2744
rect 742 2748 748 2749
rect 742 2744 743 2748
rect 747 2744 748 2748
rect 742 2743 748 2744
rect 878 2748 884 2749
rect 878 2744 879 2748
rect 883 2744 884 2748
rect 878 2743 884 2744
rect 1014 2748 1020 2749
rect 1014 2744 1015 2748
rect 1019 2744 1020 2748
rect 1014 2743 1020 2744
rect 1150 2748 1156 2749
rect 1150 2744 1151 2748
rect 1155 2744 1156 2748
rect 1150 2743 1156 2744
rect 1286 2748 1292 2749
rect 1286 2744 1287 2748
rect 1291 2744 1292 2748
rect 1286 2743 1292 2744
rect 1422 2748 1428 2749
rect 1422 2744 1423 2748
rect 1427 2744 1428 2748
rect 1422 2743 1428 2744
rect 1566 2748 1572 2749
rect 1566 2744 1567 2748
rect 1571 2744 1572 2748
rect 2008 2746 2010 2773
rect 2438 2769 2444 2770
rect 2046 2768 2052 2769
rect 2046 2764 2047 2768
rect 2051 2764 2052 2768
rect 2438 2765 2439 2769
rect 2443 2765 2444 2769
rect 2438 2764 2444 2765
rect 2566 2769 2572 2770
rect 2566 2765 2567 2769
rect 2571 2765 2572 2769
rect 2566 2764 2572 2765
rect 2694 2769 2700 2770
rect 2694 2765 2695 2769
rect 2699 2765 2700 2769
rect 2694 2764 2700 2765
rect 2830 2769 2836 2770
rect 2830 2765 2831 2769
rect 2835 2765 2836 2769
rect 2830 2764 2836 2765
rect 2966 2769 2972 2770
rect 2966 2765 2967 2769
rect 2971 2765 2972 2769
rect 2966 2764 2972 2765
rect 3102 2769 3108 2770
rect 3102 2765 3103 2769
rect 3107 2765 3108 2769
rect 3102 2764 3108 2765
rect 3246 2769 3252 2770
rect 3246 2765 3247 2769
rect 3251 2765 3252 2769
rect 3246 2764 3252 2765
rect 3390 2769 3396 2770
rect 3390 2765 3391 2769
rect 3395 2765 3396 2769
rect 3390 2764 3396 2765
rect 3542 2769 3548 2770
rect 3542 2765 3543 2769
rect 3547 2765 3548 2769
rect 3542 2764 3548 2765
rect 3702 2769 3708 2770
rect 3702 2765 3703 2769
rect 3707 2765 3708 2769
rect 3702 2764 3708 2765
rect 3838 2769 3844 2770
rect 3838 2765 3839 2769
rect 3843 2765 3844 2769
rect 3838 2764 3844 2765
rect 3942 2768 3948 2769
rect 3942 2764 3943 2768
rect 3947 2764 3948 2768
rect 2046 2763 2052 2764
rect 1566 2743 1572 2744
rect 2006 2745 2012 2746
rect 110 2740 116 2741
rect 2006 2741 2007 2745
rect 2011 2741 2012 2745
rect 2006 2740 2012 2741
rect 2048 2735 2050 2763
rect 2440 2735 2442 2764
rect 2568 2735 2570 2764
rect 2696 2735 2698 2764
rect 2832 2735 2834 2764
rect 2968 2735 2970 2764
rect 3104 2735 3106 2764
rect 3248 2735 3250 2764
rect 3392 2735 3394 2764
rect 3544 2735 3546 2764
rect 3704 2735 3706 2764
rect 3840 2735 3842 2764
rect 3942 2763 3948 2764
rect 3944 2735 3946 2763
rect 2047 2734 2051 2735
rect 238 2729 244 2730
rect 110 2728 116 2729
rect 110 2724 111 2728
rect 115 2724 116 2728
rect 238 2725 239 2729
rect 243 2725 244 2729
rect 238 2724 244 2725
rect 350 2729 356 2730
rect 350 2725 351 2729
rect 355 2725 356 2729
rect 350 2724 356 2725
rect 470 2729 476 2730
rect 470 2725 471 2729
rect 475 2725 476 2729
rect 470 2724 476 2725
rect 606 2729 612 2730
rect 606 2725 607 2729
rect 611 2725 612 2729
rect 606 2724 612 2725
rect 742 2729 748 2730
rect 742 2725 743 2729
rect 747 2725 748 2729
rect 742 2724 748 2725
rect 878 2729 884 2730
rect 878 2725 879 2729
rect 883 2725 884 2729
rect 878 2724 884 2725
rect 1014 2729 1020 2730
rect 1014 2725 1015 2729
rect 1019 2725 1020 2729
rect 1014 2724 1020 2725
rect 1150 2729 1156 2730
rect 1150 2725 1151 2729
rect 1155 2725 1156 2729
rect 1150 2724 1156 2725
rect 1286 2729 1292 2730
rect 1286 2725 1287 2729
rect 1291 2725 1292 2729
rect 1286 2724 1292 2725
rect 1422 2729 1428 2730
rect 1422 2725 1423 2729
rect 1427 2725 1428 2729
rect 1422 2724 1428 2725
rect 1566 2729 1572 2730
rect 2047 2729 2051 2730
rect 2335 2734 2339 2735
rect 2335 2729 2339 2730
rect 2439 2734 2443 2735
rect 2439 2729 2443 2730
rect 2495 2734 2499 2735
rect 2495 2729 2499 2730
rect 2567 2734 2571 2735
rect 2567 2729 2571 2730
rect 2663 2734 2667 2735
rect 2663 2729 2667 2730
rect 2695 2734 2699 2735
rect 2695 2729 2699 2730
rect 2831 2734 2835 2735
rect 2831 2729 2835 2730
rect 2967 2734 2971 2735
rect 2967 2729 2971 2730
rect 2999 2734 3003 2735
rect 2999 2729 3003 2730
rect 3103 2734 3107 2735
rect 3103 2729 3107 2730
rect 3167 2734 3171 2735
rect 3167 2729 3171 2730
rect 3247 2734 3251 2735
rect 3247 2729 3251 2730
rect 3335 2734 3339 2735
rect 3335 2729 3339 2730
rect 3391 2734 3395 2735
rect 3391 2729 3395 2730
rect 3511 2734 3515 2735
rect 3511 2729 3515 2730
rect 3543 2734 3547 2735
rect 3543 2729 3547 2730
rect 3687 2734 3691 2735
rect 3687 2729 3691 2730
rect 3703 2734 3707 2735
rect 3703 2729 3707 2730
rect 3839 2734 3843 2735
rect 3839 2729 3843 2730
rect 3943 2734 3947 2735
rect 3943 2729 3947 2730
rect 1566 2725 1567 2729
rect 1571 2725 1572 2729
rect 1566 2724 1572 2725
rect 2006 2728 2012 2729
rect 2006 2724 2007 2728
rect 2011 2724 2012 2728
rect 110 2723 116 2724
rect 112 2703 114 2723
rect 240 2703 242 2724
rect 352 2703 354 2724
rect 472 2703 474 2724
rect 608 2703 610 2724
rect 744 2703 746 2724
rect 880 2703 882 2724
rect 1016 2703 1018 2724
rect 1152 2703 1154 2724
rect 1288 2703 1290 2724
rect 1424 2703 1426 2724
rect 1568 2703 1570 2724
rect 2006 2723 2012 2724
rect 2008 2703 2010 2723
rect 2048 2709 2050 2729
rect 2046 2708 2052 2709
rect 2336 2708 2338 2729
rect 2496 2708 2498 2729
rect 2664 2708 2666 2729
rect 2832 2708 2834 2729
rect 3000 2708 3002 2729
rect 3168 2708 3170 2729
rect 3336 2708 3338 2729
rect 3512 2708 3514 2729
rect 3688 2708 3690 2729
rect 3840 2708 3842 2729
rect 3944 2709 3946 2729
rect 3942 2708 3948 2709
rect 2046 2704 2047 2708
rect 2051 2704 2052 2708
rect 2046 2703 2052 2704
rect 2334 2707 2340 2708
rect 2334 2703 2335 2707
rect 2339 2703 2340 2707
rect 111 2702 115 2703
rect 111 2697 115 2698
rect 223 2702 227 2703
rect 223 2697 227 2698
rect 239 2702 243 2703
rect 239 2697 243 2698
rect 351 2702 355 2703
rect 351 2697 355 2698
rect 367 2702 371 2703
rect 367 2697 371 2698
rect 471 2702 475 2703
rect 471 2697 475 2698
rect 503 2702 507 2703
rect 503 2697 507 2698
rect 607 2702 611 2703
rect 607 2697 611 2698
rect 639 2702 643 2703
rect 639 2697 643 2698
rect 743 2702 747 2703
rect 743 2697 747 2698
rect 767 2702 771 2703
rect 767 2697 771 2698
rect 879 2702 883 2703
rect 879 2697 883 2698
rect 887 2702 891 2703
rect 887 2697 891 2698
rect 999 2702 1003 2703
rect 999 2697 1003 2698
rect 1015 2702 1019 2703
rect 1015 2697 1019 2698
rect 1111 2702 1115 2703
rect 1111 2697 1115 2698
rect 1151 2702 1155 2703
rect 1151 2697 1155 2698
rect 1231 2702 1235 2703
rect 1231 2697 1235 2698
rect 1287 2702 1291 2703
rect 1287 2697 1291 2698
rect 1351 2702 1355 2703
rect 1351 2697 1355 2698
rect 1423 2702 1427 2703
rect 1423 2697 1427 2698
rect 1567 2702 1571 2703
rect 1567 2697 1571 2698
rect 2007 2702 2011 2703
rect 2334 2702 2340 2703
rect 2494 2707 2500 2708
rect 2494 2703 2495 2707
rect 2499 2703 2500 2707
rect 2494 2702 2500 2703
rect 2662 2707 2668 2708
rect 2662 2703 2663 2707
rect 2667 2703 2668 2707
rect 2662 2702 2668 2703
rect 2830 2707 2836 2708
rect 2830 2703 2831 2707
rect 2835 2703 2836 2707
rect 2830 2702 2836 2703
rect 2998 2707 3004 2708
rect 2998 2703 2999 2707
rect 3003 2703 3004 2707
rect 2998 2702 3004 2703
rect 3166 2707 3172 2708
rect 3166 2703 3167 2707
rect 3171 2703 3172 2707
rect 3166 2702 3172 2703
rect 3334 2707 3340 2708
rect 3334 2703 3335 2707
rect 3339 2703 3340 2707
rect 3334 2702 3340 2703
rect 3510 2707 3516 2708
rect 3510 2703 3511 2707
rect 3515 2703 3516 2707
rect 3510 2702 3516 2703
rect 3686 2707 3692 2708
rect 3686 2703 3687 2707
rect 3691 2703 3692 2707
rect 3686 2702 3692 2703
rect 3838 2707 3844 2708
rect 3838 2703 3839 2707
rect 3843 2703 3844 2707
rect 3942 2704 3943 2708
rect 3947 2704 3948 2708
rect 3942 2703 3948 2704
rect 3838 2702 3844 2703
rect 2007 2697 2011 2698
rect 112 2677 114 2697
rect 110 2676 116 2677
rect 224 2676 226 2697
rect 368 2676 370 2697
rect 504 2676 506 2697
rect 640 2676 642 2697
rect 768 2676 770 2697
rect 888 2676 890 2697
rect 1000 2676 1002 2697
rect 1112 2676 1114 2697
rect 1232 2676 1234 2697
rect 1352 2676 1354 2697
rect 2008 2677 2010 2697
rect 2046 2691 2052 2692
rect 2046 2687 2047 2691
rect 2051 2687 2052 2691
rect 3942 2691 3948 2692
rect 2046 2686 2052 2687
rect 2334 2688 2340 2689
rect 2006 2676 2012 2677
rect 110 2672 111 2676
rect 115 2672 116 2676
rect 110 2671 116 2672
rect 222 2675 228 2676
rect 222 2671 223 2675
rect 227 2671 228 2675
rect 222 2670 228 2671
rect 366 2675 372 2676
rect 366 2671 367 2675
rect 371 2671 372 2675
rect 366 2670 372 2671
rect 502 2675 508 2676
rect 502 2671 503 2675
rect 507 2671 508 2675
rect 502 2670 508 2671
rect 638 2675 644 2676
rect 638 2671 639 2675
rect 643 2671 644 2675
rect 638 2670 644 2671
rect 766 2675 772 2676
rect 766 2671 767 2675
rect 771 2671 772 2675
rect 766 2670 772 2671
rect 886 2675 892 2676
rect 886 2671 887 2675
rect 891 2671 892 2675
rect 886 2670 892 2671
rect 998 2675 1004 2676
rect 998 2671 999 2675
rect 1003 2671 1004 2675
rect 998 2670 1004 2671
rect 1110 2675 1116 2676
rect 1110 2671 1111 2675
rect 1115 2671 1116 2675
rect 1110 2670 1116 2671
rect 1230 2675 1236 2676
rect 1230 2671 1231 2675
rect 1235 2671 1236 2675
rect 1230 2670 1236 2671
rect 1350 2675 1356 2676
rect 1350 2671 1351 2675
rect 1355 2671 1356 2675
rect 2006 2672 2007 2676
rect 2011 2672 2012 2676
rect 2006 2671 2012 2672
rect 1350 2670 1356 2671
rect 110 2659 116 2660
rect 110 2655 111 2659
rect 115 2655 116 2659
rect 2006 2659 2012 2660
rect 110 2654 116 2655
rect 222 2656 228 2657
rect 112 2627 114 2654
rect 222 2652 223 2656
rect 227 2652 228 2656
rect 222 2651 228 2652
rect 366 2656 372 2657
rect 366 2652 367 2656
rect 371 2652 372 2656
rect 366 2651 372 2652
rect 502 2656 508 2657
rect 502 2652 503 2656
rect 507 2652 508 2656
rect 502 2651 508 2652
rect 638 2656 644 2657
rect 638 2652 639 2656
rect 643 2652 644 2656
rect 638 2651 644 2652
rect 766 2656 772 2657
rect 766 2652 767 2656
rect 771 2652 772 2656
rect 766 2651 772 2652
rect 886 2656 892 2657
rect 886 2652 887 2656
rect 891 2652 892 2656
rect 886 2651 892 2652
rect 998 2656 1004 2657
rect 998 2652 999 2656
rect 1003 2652 1004 2656
rect 998 2651 1004 2652
rect 1110 2656 1116 2657
rect 1110 2652 1111 2656
rect 1115 2652 1116 2656
rect 1110 2651 1116 2652
rect 1230 2656 1236 2657
rect 1230 2652 1231 2656
rect 1235 2652 1236 2656
rect 1230 2651 1236 2652
rect 1350 2656 1356 2657
rect 1350 2652 1351 2656
rect 1355 2652 1356 2656
rect 2006 2655 2007 2659
rect 2011 2655 2012 2659
rect 2048 2655 2050 2686
rect 2334 2684 2335 2688
rect 2339 2684 2340 2688
rect 2334 2683 2340 2684
rect 2494 2688 2500 2689
rect 2494 2684 2495 2688
rect 2499 2684 2500 2688
rect 2494 2683 2500 2684
rect 2662 2688 2668 2689
rect 2662 2684 2663 2688
rect 2667 2684 2668 2688
rect 2662 2683 2668 2684
rect 2830 2688 2836 2689
rect 2830 2684 2831 2688
rect 2835 2684 2836 2688
rect 2830 2683 2836 2684
rect 2998 2688 3004 2689
rect 2998 2684 2999 2688
rect 3003 2684 3004 2688
rect 2998 2683 3004 2684
rect 3166 2688 3172 2689
rect 3166 2684 3167 2688
rect 3171 2684 3172 2688
rect 3166 2683 3172 2684
rect 3334 2688 3340 2689
rect 3334 2684 3335 2688
rect 3339 2684 3340 2688
rect 3334 2683 3340 2684
rect 3510 2688 3516 2689
rect 3510 2684 3511 2688
rect 3515 2684 3516 2688
rect 3510 2683 3516 2684
rect 3686 2688 3692 2689
rect 3686 2684 3687 2688
rect 3691 2684 3692 2688
rect 3686 2683 3692 2684
rect 3838 2688 3844 2689
rect 3838 2684 3839 2688
rect 3843 2684 3844 2688
rect 3942 2687 3943 2691
rect 3947 2687 3948 2691
rect 3942 2686 3948 2687
rect 3838 2683 3844 2684
rect 2336 2655 2338 2683
rect 2496 2655 2498 2683
rect 2664 2655 2666 2683
rect 2832 2655 2834 2683
rect 3000 2655 3002 2683
rect 3168 2655 3170 2683
rect 3336 2655 3338 2683
rect 3512 2655 3514 2683
rect 3688 2655 3690 2683
rect 3840 2655 3842 2683
rect 3944 2655 3946 2686
rect 2006 2654 2012 2655
rect 2047 2654 2051 2655
rect 1350 2651 1356 2652
rect 224 2627 226 2651
rect 368 2627 370 2651
rect 504 2627 506 2651
rect 640 2627 642 2651
rect 768 2627 770 2651
rect 888 2627 890 2651
rect 1000 2627 1002 2651
rect 1112 2627 1114 2651
rect 1232 2627 1234 2651
rect 1352 2627 1354 2651
rect 2008 2627 2010 2654
rect 2047 2649 2051 2650
rect 2127 2654 2131 2655
rect 2127 2649 2131 2650
rect 2279 2654 2283 2655
rect 2279 2649 2283 2650
rect 2335 2654 2339 2655
rect 2335 2649 2339 2650
rect 2447 2654 2451 2655
rect 2447 2649 2451 2650
rect 2495 2654 2499 2655
rect 2495 2649 2499 2650
rect 2623 2654 2627 2655
rect 2623 2649 2627 2650
rect 2663 2654 2667 2655
rect 2663 2649 2667 2650
rect 2807 2654 2811 2655
rect 2807 2649 2811 2650
rect 2831 2654 2835 2655
rect 2831 2649 2835 2650
rect 2991 2654 2995 2655
rect 2991 2649 2995 2650
rect 2999 2654 3003 2655
rect 2999 2649 3003 2650
rect 3167 2654 3171 2655
rect 3167 2649 3171 2650
rect 3175 2654 3179 2655
rect 3175 2649 3179 2650
rect 3335 2654 3339 2655
rect 3335 2649 3339 2650
rect 3351 2654 3355 2655
rect 3351 2649 3355 2650
rect 3511 2654 3515 2655
rect 3511 2649 3515 2650
rect 3519 2654 3523 2655
rect 3519 2649 3523 2650
rect 3687 2654 3691 2655
rect 3687 2649 3691 2650
rect 3839 2654 3843 2655
rect 3839 2649 3843 2650
rect 3943 2654 3947 2655
rect 3943 2649 3947 2650
rect 111 2626 115 2627
rect 111 2621 115 2622
rect 175 2626 179 2627
rect 175 2621 179 2622
rect 223 2626 227 2627
rect 223 2621 227 2622
rect 367 2626 371 2627
rect 367 2621 371 2622
rect 503 2626 507 2627
rect 503 2621 507 2622
rect 543 2626 547 2627
rect 543 2621 547 2622
rect 639 2626 643 2627
rect 639 2621 643 2622
rect 711 2626 715 2627
rect 711 2621 715 2622
rect 767 2626 771 2627
rect 767 2621 771 2622
rect 863 2626 867 2627
rect 863 2621 867 2622
rect 887 2626 891 2627
rect 887 2621 891 2622
rect 999 2626 1003 2627
rect 999 2621 1003 2622
rect 1007 2626 1011 2627
rect 1007 2621 1011 2622
rect 1111 2626 1115 2627
rect 1111 2621 1115 2622
rect 1143 2626 1147 2627
rect 1143 2621 1147 2622
rect 1231 2626 1235 2627
rect 1231 2621 1235 2622
rect 1279 2626 1283 2627
rect 1279 2621 1283 2622
rect 1351 2626 1355 2627
rect 1351 2621 1355 2622
rect 1423 2626 1427 2627
rect 1423 2621 1427 2622
rect 2007 2626 2011 2627
rect 2048 2622 2050 2649
rect 2128 2625 2130 2649
rect 2280 2625 2282 2649
rect 2448 2625 2450 2649
rect 2624 2625 2626 2649
rect 2808 2625 2810 2649
rect 2992 2625 2994 2649
rect 3176 2625 3178 2649
rect 3352 2625 3354 2649
rect 3520 2625 3522 2649
rect 3688 2625 3690 2649
rect 3840 2625 3842 2649
rect 2126 2624 2132 2625
rect 2007 2621 2011 2622
rect 2046 2621 2052 2622
rect 112 2594 114 2621
rect 176 2597 178 2621
rect 368 2597 370 2621
rect 544 2597 546 2621
rect 712 2597 714 2621
rect 864 2597 866 2621
rect 1008 2597 1010 2621
rect 1144 2597 1146 2621
rect 1280 2597 1282 2621
rect 1424 2597 1426 2621
rect 174 2596 180 2597
rect 110 2593 116 2594
rect 110 2589 111 2593
rect 115 2589 116 2593
rect 174 2592 175 2596
rect 179 2592 180 2596
rect 174 2591 180 2592
rect 366 2596 372 2597
rect 366 2592 367 2596
rect 371 2592 372 2596
rect 366 2591 372 2592
rect 542 2596 548 2597
rect 542 2592 543 2596
rect 547 2592 548 2596
rect 542 2591 548 2592
rect 710 2596 716 2597
rect 710 2592 711 2596
rect 715 2592 716 2596
rect 710 2591 716 2592
rect 862 2596 868 2597
rect 862 2592 863 2596
rect 867 2592 868 2596
rect 862 2591 868 2592
rect 1006 2596 1012 2597
rect 1006 2592 1007 2596
rect 1011 2592 1012 2596
rect 1006 2591 1012 2592
rect 1142 2596 1148 2597
rect 1142 2592 1143 2596
rect 1147 2592 1148 2596
rect 1142 2591 1148 2592
rect 1278 2596 1284 2597
rect 1278 2592 1279 2596
rect 1283 2592 1284 2596
rect 1278 2591 1284 2592
rect 1422 2596 1428 2597
rect 1422 2592 1423 2596
rect 1427 2592 1428 2596
rect 2008 2594 2010 2621
rect 2046 2617 2047 2621
rect 2051 2617 2052 2621
rect 2126 2620 2127 2624
rect 2131 2620 2132 2624
rect 2126 2619 2132 2620
rect 2278 2624 2284 2625
rect 2278 2620 2279 2624
rect 2283 2620 2284 2624
rect 2278 2619 2284 2620
rect 2446 2624 2452 2625
rect 2446 2620 2447 2624
rect 2451 2620 2452 2624
rect 2446 2619 2452 2620
rect 2622 2624 2628 2625
rect 2622 2620 2623 2624
rect 2627 2620 2628 2624
rect 2622 2619 2628 2620
rect 2806 2624 2812 2625
rect 2806 2620 2807 2624
rect 2811 2620 2812 2624
rect 2806 2619 2812 2620
rect 2990 2624 2996 2625
rect 2990 2620 2991 2624
rect 2995 2620 2996 2624
rect 2990 2619 2996 2620
rect 3174 2624 3180 2625
rect 3174 2620 3175 2624
rect 3179 2620 3180 2624
rect 3174 2619 3180 2620
rect 3350 2624 3356 2625
rect 3350 2620 3351 2624
rect 3355 2620 3356 2624
rect 3350 2619 3356 2620
rect 3518 2624 3524 2625
rect 3518 2620 3519 2624
rect 3523 2620 3524 2624
rect 3518 2619 3524 2620
rect 3686 2624 3692 2625
rect 3686 2620 3687 2624
rect 3691 2620 3692 2624
rect 3686 2619 3692 2620
rect 3838 2624 3844 2625
rect 3838 2620 3839 2624
rect 3843 2620 3844 2624
rect 3944 2622 3946 2649
rect 3838 2619 3844 2620
rect 3942 2621 3948 2622
rect 2046 2616 2052 2617
rect 3942 2617 3943 2621
rect 3947 2617 3948 2621
rect 3942 2616 3948 2617
rect 2126 2605 2132 2606
rect 2046 2604 2052 2605
rect 2046 2600 2047 2604
rect 2051 2600 2052 2604
rect 2126 2601 2127 2605
rect 2131 2601 2132 2605
rect 2126 2600 2132 2601
rect 2278 2605 2284 2606
rect 2278 2601 2279 2605
rect 2283 2601 2284 2605
rect 2278 2600 2284 2601
rect 2446 2605 2452 2606
rect 2446 2601 2447 2605
rect 2451 2601 2452 2605
rect 2446 2600 2452 2601
rect 2622 2605 2628 2606
rect 2622 2601 2623 2605
rect 2627 2601 2628 2605
rect 2622 2600 2628 2601
rect 2806 2605 2812 2606
rect 2806 2601 2807 2605
rect 2811 2601 2812 2605
rect 2806 2600 2812 2601
rect 2990 2605 2996 2606
rect 2990 2601 2991 2605
rect 2995 2601 2996 2605
rect 2990 2600 2996 2601
rect 3174 2605 3180 2606
rect 3174 2601 3175 2605
rect 3179 2601 3180 2605
rect 3174 2600 3180 2601
rect 3350 2605 3356 2606
rect 3350 2601 3351 2605
rect 3355 2601 3356 2605
rect 3350 2600 3356 2601
rect 3518 2605 3524 2606
rect 3518 2601 3519 2605
rect 3523 2601 3524 2605
rect 3518 2600 3524 2601
rect 3686 2605 3692 2606
rect 3686 2601 3687 2605
rect 3691 2601 3692 2605
rect 3686 2600 3692 2601
rect 3838 2605 3844 2606
rect 3838 2601 3839 2605
rect 3843 2601 3844 2605
rect 3838 2600 3844 2601
rect 3942 2604 3948 2605
rect 3942 2600 3943 2604
rect 3947 2600 3948 2604
rect 2046 2599 2052 2600
rect 1422 2591 1428 2592
rect 2006 2593 2012 2594
rect 110 2588 116 2589
rect 2006 2589 2007 2593
rect 2011 2589 2012 2593
rect 2006 2588 2012 2589
rect 174 2577 180 2578
rect 110 2576 116 2577
rect 110 2572 111 2576
rect 115 2572 116 2576
rect 174 2573 175 2577
rect 179 2573 180 2577
rect 174 2572 180 2573
rect 366 2577 372 2578
rect 366 2573 367 2577
rect 371 2573 372 2577
rect 366 2572 372 2573
rect 542 2577 548 2578
rect 542 2573 543 2577
rect 547 2573 548 2577
rect 542 2572 548 2573
rect 710 2577 716 2578
rect 710 2573 711 2577
rect 715 2573 716 2577
rect 710 2572 716 2573
rect 862 2577 868 2578
rect 862 2573 863 2577
rect 867 2573 868 2577
rect 862 2572 868 2573
rect 1006 2577 1012 2578
rect 1006 2573 1007 2577
rect 1011 2573 1012 2577
rect 1006 2572 1012 2573
rect 1142 2577 1148 2578
rect 1142 2573 1143 2577
rect 1147 2573 1148 2577
rect 1142 2572 1148 2573
rect 1278 2577 1284 2578
rect 1278 2573 1279 2577
rect 1283 2573 1284 2577
rect 1278 2572 1284 2573
rect 1422 2577 1428 2578
rect 1422 2573 1423 2577
rect 1427 2573 1428 2577
rect 1422 2572 1428 2573
rect 2006 2576 2012 2577
rect 2006 2572 2007 2576
rect 2011 2572 2012 2576
rect 110 2571 116 2572
rect 112 2547 114 2571
rect 176 2547 178 2572
rect 368 2547 370 2572
rect 544 2547 546 2572
rect 712 2547 714 2572
rect 864 2547 866 2572
rect 1008 2547 1010 2572
rect 1144 2547 1146 2572
rect 1280 2547 1282 2572
rect 1424 2547 1426 2572
rect 2006 2571 2012 2572
rect 2048 2571 2050 2599
rect 2128 2571 2130 2600
rect 2280 2571 2282 2600
rect 2448 2571 2450 2600
rect 2624 2571 2626 2600
rect 2808 2571 2810 2600
rect 2992 2571 2994 2600
rect 3176 2571 3178 2600
rect 3352 2571 3354 2600
rect 3520 2571 3522 2600
rect 3688 2571 3690 2600
rect 3840 2571 3842 2600
rect 3942 2599 3948 2600
rect 3944 2571 3946 2599
rect 2008 2547 2010 2571
rect 2047 2570 2051 2571
rect 2047 2565 2051 2566
rect 2071 2570 2075 2571
rect 2071 2565 2075 2566
rect 2127 2570 2131 2571
rect 2127 2565 2131 2566
rect 2183 2570 2187 2571
rect 2183 2565 2187 2566
rect 2279 2570 2283 2571
rect 2279 2565 2283 2566
rect 2319 2570 2323 2571
rect 2319 2565 2323 2566
rect 2447 2570 2451 2571
rect 2447 2565 2451 2566
rect 2471 2570 2475 2571
rect 2471 2565 2475 2566
rect 2623 2570 2627 2571
rect 2623 2565 2627 2566
rect 2639 2570 2643 2571
rect 2639 2565 2643 2566
rect 2807 2570 2811 2571
rect 2807 2565 2811 2566
rect 2823 2570 2827 2571
rect 2823 2565 2827 2566
rect 2991 2570 2995 2571
rect 2991 2565 2995 2566
rect 3031 2570 3035 2571
rect 3031 2565 3035 2566
rect 3175 2570 3179 2571
rect 3175 2565 3179 2566
rect 3263 2570 3267 2571
rect 3263 2565 3267 2566
rect 3351 2570 3355 2571
rect 3351 2565 3355 2566
rect 3503 2570 3507 2571
rect 3503 2565 3507 2566
rect 3519 2570 3523 2571
rect 3519 2565 3523 2566
rect 3687 2570 3691 2571
rect 3687 2565 3691 2566
rect 3743 2570 3747 2571
rect 3743 2565 3747 2566
rect 3839 2570 3843 2571
rect 3839 2565 3843 2566
rect 3943 2570 3947 2571
rect 3943 2565 3947 2566
rect 111 2546 115 2547
rect 111 2541 115 2542
rect 135 2546 139 2547
rect 135 2541 139 2542
rect 175 2546 179 2547
rect 175 2541 179 2542
rect 271 2546 275 2547
rect 271 2541 275 2542
rect 367 2546 371 2547
rect 367 2541 371 2542
rect 439 2546 443 2547
rect 439 2541 443 2542
rect 543 2546 547 2547
rect 543 2541 547 2542
rect 607 2546 611 2547
rect 607 2541 611 2542
rect 711 2546 715 2547
rect 711 2541 715 2542
rect 775 2546 779 2547
rect 775 2541 779 2542
rect 863 2546 867 2547
rect 863 2541 867 2542
rect 927 2546 931 2547
rect 927 2541 931 2542
rect 1007 2546 1011 2547
rect 1007 2541 1011 2542
rect 1079 2546 1083 2547
rect 1079 2541 1083 2542
rect 1143 2546 1147 2547
rect 1143 2541 1147 2542
rect 1223 2546 1227 2547
rect 1223 2541 1227 2542
rect 1279 2546 1283 2547
rect 1279 2541 1283 2542
rect 1359 2546 1363 2547
rect 1359 2541 1363 2542
rect 1423 2546 1427 2547
rect 1423 2541 1427 2542
rect 1495 2546 1499 2547
rect 1495 2541 1499 2542
rect 1639 2546 1643 2547
rect 1639 2541 1643 2542
rect 2007 2546 2011 2547
rect 2048 2545 2050 2565
rect 2007 2541 2011 2542
rect 2046 2544 2052 2545
rect 2072 2544 2074 2565
rect 2184 2544 2186 2565
rect 2320 2544 2322 2565
rect 2472 2544 2474 2565
rect 2640 2544 2642 2565
rect 2824 2544 2826 2565
rect 3032 2544 3034 2565
rect 3264 2544 3266 2565
rect 3504 2544 3506 2565
rect 3744 2544 3746 2565
rect 3944 2545 3946 2565
rect 3942 2544 3948 2545
rect 112 2521 114 2541
rect 110 2520 116 2521
rect 136 2520 138 2541
rect 272 2520 274 2541
rect 440 2520 442 2541
rect 608 2520 610 2541
rect 776 2520 778 2541
rect 928 2520 930 2541
rect 1080 2520 1082 2541
rect 1224 2520 1226 2541
rect 1360 2520 1362 2541
rect 1496 2520 1498 2541
rect 1640 2520 1642 2541
rect 2008 2521 2010 2541
rect 2046 2540 2047 2544
rect 2051 2540 2052 2544
rect 2046 2539 2052 2540
rect 2070 2543 2076 2544
rect 2070 2539 2071 2543
rect 2075 2539 2076 2543
rect 2070 2538 2076 2539
rect 2182 2543 2188 2544
rect 2182 2539 2183 2543
rect 2187 2539 2188 2543
rect 2182 2538 2188 2539
rect 2318 2543 2324 2544
rect 2318 2539 2319 2543
rect 2323 2539 2324 2543
rect 2318 2538 2324 2539
rect 2470 2543 2476 2544
rect 2470 2539 2471 2543
rect 2475 2539 2476 2543
rect 2470 2538 2476 2539
rect 2638 2543 2644 2544
rect 2638 2539 2639 2543
rect 2643 2539 2644 2543
rect 2638 2538 2644 2539
rect 2822 2543 2828 2544
rect 2822 2539 2823 2543
rect 2827 2539 2828 2543
rect 2822 2538 2828 2539
rect 3030 2543 3036 2544
rect 3030 2539 3031 2543
rect 3035 2539 3036 2543
rect 3030 2538 3036 2539
rect 3262 2543 3268 2544
rect 3262 2539 3263 2543
rect 3267 2539 3268 2543
rect 3262 2538 3268 2539
rect 3502 2543 3508 2544
rect 3502 2539 3503 2543
rect 3507 2539 3508 2543
rect 3502 2538 3508 2539
rect 3742 2543 3748 2544
rect 3742 2539 3743 2543
rect 3747 2539 3748 2543
rect 3942 2540 3943 2544
rect 3947 2540 3948 2544
rect 3942 2539 3948 2540
rect 3742 2538 3748 2539
rect 2046 2527 2052 2528
rect 2046 2523 2047 2527
rect 2051 2523 2052 2527
rect 3942 2527 3948 2528
rect 2046 2522 2052 2523
rect 2070 2524 2076 2525
rect 2006 2520 2012 2521
rect 110 2516 111 2520
rect 115 2516 116 2520
rect 110 2515 116 2516
rect 134 2519 140 2520
rect 134 2515 135 2519
rect 139 2515 140 2519
rect 134 2514 140 2515
rect 270 2519 276 2520
rect 270 2515 271 2519
rect 275 2515 276 2519
rect 270 2514 276 2515
rect 438 2519 444 2520
rect 438 2515 439 2519
rect 443 2515 444 2519
rect 438 2514 444 2515
rect 606 2519 612 2520
rect 606 2515 607 2519
rect 611 2515 612 2519
rect 606 2514 612 2515
rect 774 2519 780 2520
rect 774 2515 775 2519
rect 779 2515 780 2519
rect 774 2514 780 2515
rect 926 2519 932 2520
rect 926 2515 927 2519
rect 931 2515 932 2519
rect 926 2514 932 2515
rect 1078 2519 1084 2520
rect 1078 2515 1079 2519
rect 1083 2515 1084 2519
rect 1078 2514 1084 2515
rect 1222 2519 1228 2520
rect 1222 2515 1223 2519
rect 1227 2515 1228 2519
rect 1222 2514 1228 2515
rect 1358 2519 1364 2520
rect 1358 2515 1359 2519
rect 1363 2515 1364 2519
rect 1358 2514 1364 2515
rect 1494 2519 1500 2520
rect 1494 2515 1495 2519
rect 1499 2515 1500 2519
rect 1494 2514 1500 2515
rect 1638 2519 1644 2520
rect 1638 2515 1639 2519
rect 1643 2515 1644 2519
rect 2006 2516 2007 2520
rect 2011 2516 2012 2520
rect 2006 2515 2012 2516
rect 1638 2514 1644 2515
rect 110 2503 116 2504
rect 110 2499 111 2503
rect 115 2499 116 2503
rect 2006 2503 2012 2504
rect 110 2498 116 2499
rect 134 2500 140 2501
rect 112 2467 114 2498
rect 134 2496 135 2500
rect 139 2496 140 2500
rect 134 2495 140 2496
rect 270 2500 276 2501
rect 270 2496 271 2500
rect 275 2496 276 2500
rect 270 2495 276 2496
rect 438 2500 444 2501
rect 438 2496 439 2500
rect 443 2496 444 2500
rect 438 2495 444 2496
rect 606 2500 612 2501
rect 606 2496 607 2500
rect 611 2496 612 2500
rect 606 2495 612 2496
rect 774 2500 780 2501
rect 774 2496 775 2500
rect 779 2496 780 2500
rect 774 2495 780 2496
rect 926 2500 932 2501
rect 926 2496 927 2500
rect 931 2496 932 2500
rect 926 2495 932 2496
rect 1078 2500 1084 2501
rect 1078 2496 1079 2500
rect 1083 2496 1084 2500
rect 1078 2495 1084 2496
rect 1222 2500 1228 2501
rect 1222 2496 1223 2500
rect 1227 2496 1228 2500
rect 1222 2495 1228 2496
rect 1358 2500 1364 2501
rect 1358 2496 1359 2500
rect 1363 2496 1364 2500
rect 1358 2495 1364 2496
rect 1494 2500 1500 2501
rect 1494 2496 1495 2500
rect 1499 2496 1500 2500
rect 1494 2495 1500 2496
rect 1638 2500 1644 2501
rect 1638 2496 1639 2500
rect 1643 2496 1644 2500
rect 2006 2499 2007 2503
rect 2011 2499 2012 2503
rect 2006 2498 2012 2499
rect 1638 2495 1644 2496
rect 136 2467 138 2495
rect 272 2467 274 2495
rect 440 2467 442 2495
rect 608 2467 610 2495
rect 776 2467 778 2495
rect 928 2467 930 2495
rect 1080 2467 1082 2495
rect 1224 2467 1226 2495
rect 1360 2467 1362 2495
rect 1496 2467 1498 2495
rect 1640 2467 1642 2495
rect 2008 2467 2010 2498
rect 2048 2491 2050 2522
rect 2070 2520 2071 2524
rect 2075 2520 2076 2524
rect 2070 2519 2076 2520
rect 2182 2524 2188 2525
rect 2182 2520 2183 2524
rect 2187 2520 2188 2524
rect 2182 2519 2188 2520
rect 2318 2524 2324 2525
rect 2318 2520 2319 2524
rect 2323 2520 2324 2524
rect 2318 2519 2324 2520
rect 2470 2524 2476 2525
rect 2470 2520 2471 2524
rect 2475 2520 2476 2524
rect 2470 2519 2476 2520
rect 2638 2524 2644 2525
rect 2638 2520 2639 2524
rect 2643 2520 2644 2524
rect 2638 2519 2644 2520
rect 2822 2524 2828 2525
rect 2822 2520 2823 2524
rect 2827 2520 2828 2524
rect 2822 2519 2828 2520
rect 3030 2524 3036 2525
rect 3030 2520 3031 2524
rect 3035 2520 3036 2524
rect 3030 2519 3036 2520
rect 3262 2524 3268 2525
rect 3262 2520 3263 2524
rect 3267 2520 3268 2524
rect 3262 2519 3268 2520
rect 3502 2524 3508 2525
rect 3502 2520 3503 2524
rect 3507 2520 3508 2524
rect 3502 2519 3508 2520
rect 3742 2524 3748 2525
rect 3742 2520 3743 2524
rect 3747 2520 3748 2524
rect 3942 2523 3943 2527
rect 3947 2523 3948 2527
rect 3942 2522 3948 2523
rect 3742 2519 3748 2520
rect 2072 2491 2074 2519
rect 2184 2491 2186 2519
rect 2320 2491 2322 2519
rect 2472 2491 2474 2519
rect 2640 2491 2642 2519
rect 2824 2491 2826 2519
rect 3032 2491 3034 2519
rect 3264 2491 3266 2519
rect 3504 2491 3506 2519
rect 3744 2491 3746 2519
rect 3944 2491 3946 2522
rect 2047 2490 2051 2491
rect 2047 2485 2051 2486
rect 2071 2490 2075 2491
rect 2071 2485 2075 2486
rect 2183 2490 2187 2491
rect 2183 2485 2187 2486
rect 2215 2490 2219 2491
rect 2215 2485 2219 2486
rect 2319 2490 2323 2491
rect 2319 2485 2323 2486
rect 2383 2490 2387 2491
rect 2383 2485 2387 2486
rect 2471 2490 2475 2491
rect 2471 2485 2475 2486
rect 2559 2490 2563 2491
rect 2559 2485 2563 2486
rect 2639 2490 2643 2491
rect 2639 2485 2643 2486
rect 2751 2490 2755 2491
rect 2751 2485 2755 2486
rect 2823 2490 2827 2491
rect 2823 2485 2827 2486
rect 2951 2490 2955 2491
rect 2951 2485 2955 2486
rect 3031 2490 3035 2491
rect 3031 2485 3035 2486
rect 3167 2490 3171 2491
rect 3167 2485 3171 2486
rect 3263 2490 3267 2491
rect 3263 2485 3267 2486
rect 3391 2490 3395 2491
rect 3391 2485 3395 2486
rect 3503 2490 3507 2491
rect 3503 2485 3507 2486
rect 3623 2490 3627 2491
rect 3623 2485 3627 2486
rect 3743 2490 3747 2491
rect 3743 2485 3747 2486
rect 3839 2490 3843 2491
rect 3839 2485 3843 2486
rect 3943 2490 3947 2491
rect 3943 2485 3947 2486
rect 111 2466 115 2467
rect 111 2461 115 2462
rect 135 2466 139 2467
rect 135 2461 139 2462
rect 271 2466 275 2467
rect 271 2461 275 2462
rect 311 2466 315 2467
rect 311 2461 315 2462
rect 439 2466 443 2467
rect 439 2461 443 2462
rect 511 2466 515 2467
rect 511 2461 515 2462
rect 607 2466 611 2467
rect 607 2461 611 2462
rect 711 2466 715 2467
rect 711 2461 715 2462
rect 775 2466 779 2467
rect 775 2461 779 2462
rect 903 2466 907 2467
rect 903 2461 907 2462
rect 927 2466 931 2467
rect 927 2461 931 2462
rect 1079 2466 1083 2467
rect 1079 2461 1083 2462
rect 1223 2466 1227 2467
rect 1223 2461 1227 2462
rect 1239 2466 1243 2467
rect 1239 2461 1243 2462
rect 1359 2466 1363 2467
rect 1359 2461 1363 2462
rect 1391 2466 1395 2467
rect 1391 2461 1395 2462
rect 1495 2466 1499 2467
rect 1495 2461 1499 2462
rect 1527 2466 1531 2467
rect 1527 2461 1531 2462
rect 1639 2466 1643 2467
rect 1639 2461 1643 2462
rect 1663 2466 1667 2467
rect 1663 2461 1667 2462
rect 1791 2466 1795 2467
rect 1791 2461 1795 2462
rect 1903 2466 1907 2467
rect 1903 2461 1907 2462
rect 2007 2466 2011 2467
rect 2007 2461 2011 2462
rect 112 2434 114 2461
rect 136 2437 138 2461
rect 312 2437 314 2461
rect 512 2437 514 2461
rect 712 2437 714 2461
rect 904 2437 906 2461
rect 1080 2437 1082 2461
rect 1240 2437 1242 2461
rect 1392 2437 1394 2461
rect 1528 2437 1530 2461
rect 1664 2437 1666 2461
rect 1792 2437 1794 2461
rect 1904 2437 1906 2461
rect 134 2436 140 2437
rect 110 2433 116 2434
rect 110 2429 111 2433
rect 115 2429 116 2433
rect 134 2432 135 2436
rect 139 2432 140 2436
rect 134 2431 140 2432
rect 310 2436 316 2437
rect 310 2432 311 2436
rect 315 2432 316 2436
rect 310 2431 316 2432
rect 510 2436 516 2437
rect 510 2432 511 2436
rect 515 2432 516 2436
rect 510 2431 516 2432
rect 710 2436 716 2437
rect 710 2432 711 2436
rect 715 2432 716 2436
rect 710 2431 716 2432
rect 902 2436 908 2437
rect 902 2432 903 2436
rect 907 2432 908 2436
rect 902 2431 908 2432
rect 1078 2436 1084 2437
rect 1078 2432 1079 2436
rect 1083 2432 1084 2436
rect 1078 2431 1084 2432
rect 1238 2436 1244 2437
rect 1238 2432 1239 2436
rect 1243 2432 1244 2436
rect 1238 2431 1244 2432
rect 1390 2436 1396 2437
rect 1390 2432 1391 2436
rect 1395 2432 1396 2436
rect 1390 2431 1396 2432
rect 1526 2436 1532 2437
rect 1526 2432 1527 2436
rect 1531 2432 1532 2436
rect 1526 2431 1532 2432
rect 1662 2436 1668 2437
rect 1662 2432 1663 2436
rect 1667 2432 1668 2436
rect 1662 2431 1668 2432
rect 1790 2436 1796 2437
rect 1790 2432 1791 2436
rect 1795 2432 1796 2436
rect 1790 2431 1796 2432
rect 1902 2436 1908 2437
rect 1902 2432 1903 2436
rect 1907 2432 1908 2436
rect 2008 2434 2010 2461
rect 2048 2458 2050 2485
rect 2072 2461 2074 2485
rect 2216 2461 2218 2485
rect 2384 2461 2386 2485
rect 2560 2461 2562 2485
rect 2752 2461 2754 2485
rect 2952 2461 2954 2485
rect 3168 2461 3170 2485
rect 3392 2461 3394 2485
rect 3624 2461 3626 2485
rect 3840 2461 3842 2485
rect 2070 2460 2076 2461
rect 2046 2457 2052 2458
rect 2046 2453 2047 2457
rect 2051 2453 2052 2457
rect 2070 2456 2071 2460
rect 2075 2456 2076 2460
rect 2070 2455 2076 2456
rect 2214 2460 2220 2461
rect 2214 2456 2215 2460
rect 2219 2456 2220 2460
rect 2214 2455 2220 2456
rect 2382 2460 2388 2461
rect 2382 2456 2383 2460
rect 2387 2456 2388 2460
rect 2382 2455 2388 2456
rect 2558 2460 2564 2461
rect 2558 2456 2559 2460
rect 2563 2456 2564 2460
rect 2558 2455 2564 2456
rect 2750 2460 2756 2461
rect 2750 2456 2751 2460
rect 2755 2456 2756 2460
rect 2750 2455 2756 2456
rect 2950 2460 2956 2461
rect 2950 2456 2951 2460
rect 2955 2456 2956 2460
rect 2950 2455 2956 2456
rect 3166 2460 3172 2461
rect 3166 2456 3167 2460
rect 3171 2456 3172 2460
rect 3166 2455 3172 2456
rect 3390 2460 3396 2461
rect 3390 2456 3391 2460
rect 3395 2456 3396 2460
rect 3390 2455 3396 2456
rect 3622 2460 3628 2461
rect 3622 2456 3623 2460
rect 3627 2456 3628 2460
rect 3622 2455 3628 2456
rect 3838 2460 3844 2461
rect 3838 2456 3839 2460
rect 3843 2456 3844 2460
rect 3944 2458 3946 2485
rect 3838 2455 3844 2456
rect 3942 2457 3948 2458
rect 2046 2452 2052 2453
rect 3942 2453 3943 2457
rect 3947 2453 3948 2457
rect 3942 2452 3948 2453
rect 2070 2441 2076 2442
rect 2046 2440 2052 2441
rect 2046 2436 2047 2440
rect 2051 2436 2052 2440
rect 2070 2437 2071 2441
rect 2075 2437 2076 2441
rect 2070 2436 2076 2437
rect 2214 2441 2220 2442
rect 2214 2437 2215 2441
rect 2219 2437 2220 2441
rect 2214 2436 2220 2437
rect 2382 2441 2388 2442
rect 2382 2437 2383 2441
rect 2387 2437 2388 2441
rect 2382 2436 2388 2437
rect 2558 2441 2564 2442
rect 2558 2437 2559 2441
rect 2563 2437 2564 2441
rect 2558 2436 2564 2437
rect 2750 2441 2756 2442
rect 2750 2437 2751 2441
rect 2755 2437 2756 2441
rect 2750 2436 2756 2437
rect 2950 2441 2956 2442
rect 2950 2437 2951 2441
rect 2955 2437 2956 2441
rect 2950 2436 2956 2437
rect 3166 2441 3172 2442
rect 3166 2437 3167 2441
rect 3171 2437 3172 2441
rect 3166 2436 3172 2437
rect 3390 2441 3396 2442
rect 3390 2437 3391 2441
rect 3395 2437 3396 2441
rect 3390 2436 3396 2437
rect 3622 2441 3628 2442
rect 3622 2437 3623 2441
rect 3627 2437 3628 2441
rect 3622 2436 3628 2437
rect 3838 2441 3844 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3942 2440 3948 2441
rect 3942 2436 3943 2440
rect 3947 2436 3948 2440
rect 2046 2435 2052 2436
rect 1902 2431 1908 2432
rect 2006 2433 2012 2434
rect 110 2428 116 2429
rect 2006 2429 2007 2433
rect 2011 2429 2012 2433
rect 2006 2428 2012 2429
rect 134 2417 140 2418
rect 110 2416 116 2417
rect 110 2412 111 2416
rect 115 2412 116 2416
rect 134 2413 135 2417
rect 139 2413 140 2417
rect 134 2412 140 2413
rect 310 2417 316 2418
rect 310 2413 311 2417
rect 315 2413 316 2417
rect 310 2412 316 2413
rect 510 2417 516 2418
rect 510 2413 511 2417
rect 515 2413 516 2417
rect 510 2412 516 2413
rect 710 2417 716 2418
rect 710 2413 711 2417
rect 715 2413 716 2417
rect 710 2412 716 2413
rect 902 2417 908 2418
rect 902 2413 903 2417
rect 907 2413 908 2417
rect 902 2412 908 2413
rect 1078 2417 1084 2418
rect 1078 2413 1079 2417
rect 1083 2413 1084 2417
rect 1078 2412 1084 2413
rect 1238 2417 1244 2418
rect 1238 2413 1239 2417
rect 1243 2413 1244 2417
rect 1238 2412 1244 2413
rect 1390 2417 1396 2418
rect 1390 2413 1391 2417
rect 1395 2413 1396 2417
rect 1390 2412 1396 2413
rect 1526 2417 1532 2418
rect 1526 2413 1527 2417
rect 1531 2413 1532 2417
rect 1526 2412 1532 2413
rect 1662 2417 1668 2418
rect 1662 2413 1663 2417
rect 1667 2413 1668 2417
rect 1662 2412 1668 2413
rect 1790 2417 1796 2418
rect 1790 2413 1791 2417
rect 1795 2413 1796 2417
rect 1790 2412 1796 2413
rect 1902 2417 1908 2418
rect 1902 2413 1903 2417
rect 1907 2413 1908 2417
rect 1902 2412 1908 2413
rect 2006 2416 2012 2417
rect 2006 2412 2007 2416
rect 2011 2412 2012 2416
rect 110 2411 116 2412
rect 112 2391 114 2411
rect 136 2391 138 2412
rect 312 2391 314 2412
rect 512 2391 514 2412
rect 712 2391 714 2412
rect 904 2391 906 2412
rect 1080 2391 1082 2412
rect 1240 2391 1242 2412
rect 1392 2391 1394 2412
rect 1528 2391 1530 2412
rect 1664 2391 1666 2412
rect 1792 2391 1794 2412
rect 1904 2391 1906 2412
rect 2006 2411 2012 2412
rect 2008 2391 2010 2411
rect 2048 2399 2050 2435
rect 2072 2399 2074 2436
rect 2216 2399 2218 2436
rect 2384 2399 2386 2436
rect 2560 2399 2562 2436
rect 2752 2399 2754 2436
rect 2952 2399 2954 2436
rect 3168 2399 3170 2436
rect 3392 2399 3394 2436
rect 3624 2399 3626 2436
rect 3840 2399 3842 2436
rect 3942 2435 3948 2436
rect 3944 2399 3946 2435
rect 2047 2398 2051 2399
rect 2047 2393 2051 2394
rect 2071 2398 2075 2399
rect 2071 2393 2075 2394
rect 2215 2398 2219 2399
rect 2215 2393 2219 2394
rect 2247 2398 2251 2399
rect 2247 2393 2251 2394
rect 2383 2398 2387 2399
rect 2383 2393 2387 2394
rect 2431 2398 2435 2399
rect 2431 2393 2435 2394
rect 2559 2398 2563 2399
rect 2559 2393 2563 2394
rect 2607 2398 2611 2399
rect 2607 2393 2611 2394
rect 2751 2398 2755 2399
rect 2751 2393 2755 2394
rect 2775 2398 2779 2399
rect 2775 2393 2779 2394
rect 2935 2398 2939 2399
rect 2935 2393 2939 2394
rect 2951 2398 2955 2399
rect 2951 2393 2955 2394
rect 3103 2398 3107 2399
rect 3103 2393 3107 2394
rect 3167 2398 3171 2399
rect 3167 2393 3171 2394
rect 3391 2398 3395 2399
rect 3391 2393 3395 2394
rect 3623 2398 3627 2399
rect 3623 2393 3627 2394
rect 3839 2398 3843 2399
rect 3839 2393 3843 2394
rect 3943 2398 3947 2399
rect 3943 2393 3947 2394
rect 111 2390 115 2391
rect 111 2385 115 2386
rect 135 2390 139 2391
rect 135 2385 139 2386
rect 311 2390 315 2391
rect 311 2385 315 2386
rect 327 2390 331 2391
rect 327 2385 331 2386
rect 511 2390 515 2391
rect 511 2385 515 2386
rect 551 2390 555 2391
rect 551 2385 555 2386
rect 711 2390 715 2391
rect 711 2385 715 2386
rect 767 2390 771 2391
rect 767 2385 771 2386
rect 903 2390 907 2391
rect 903 2385 907 2386
rect 975 2390 979 2391
rect 975 2385 979 2386
rect 1079 2390 1083 2391
rect 1079 2385 1083 2386
rect 1175 2390 1179 2391
rect 1175 2385 1179 2386
rect 1239 2390 1243 2391
rect 1239 2385 1243 2386
rect 1367 2390 1371 2391
rect 1367 2385 1371 2386
rect 1391 2390 1395 2391
rect 1391 2385 1395 2386
rect 1527 2390 1531 2391
rect 1527 2385 1531 2386
rect 1551 2390 1555 2391
rect 1551 2385 1555 2386
rect 1663 2390 1667 2391
rect 1663 2385 1667 2386
rect 1735 2390 1739 2391
rect 1735 2385 1739 2386
rect 1791 2390 1795 2391
rect 1791 2385 1795 2386
rect 1903 2390 1907 2391
rect 1903 2385 1907 2386
rect 2007 2390 2011 2391
rect 2007 2385 2011 2386
rect 112 2365 114 2385
rect 110 2364 116 2365
rect 136 2364 138 2385
rect 328 2364 330 2385
rect 552 2364 554 2385
rect 768 2364 770 2385
rect 976 2364 978 2385
rect 1176 2364 1178 2385
rect 1368 2364 1370 2385
rect 1552 2364 1554 2385
rect 1736 2364 1738 2385
rect 1904 2364 1906 2385
rect 2008 2365 2010 2385
rect 2048 2373 2050 2393
rect 2046 2372 2052 2373
rect 2072 2372 2074 2393
rect 2248 2372 2250 2393
rect 2432 2372 2434 2393
rect 2608 2372 2610 2393
rect 2776 2372 2778 2393
rect 2936 2372 2938 2393
rect 3104 2372 3106 2393
rect 3944 2373 3946 2393
rect 3942 2372 3948 2373
rect 2046 2368 2047 2372
rect 2051 2368 2052 2372
rect 2046 2367 2052 2368
rect 2070 2371 2076 2372
rect 2070 2367 2071 2371
rect 2075 2367 2076 2371
rect 2070 2366 2076 2367
rect 2246 2371 2252 2372
rect 2246 2367 2247 2371
rect 2251 2367 2252 2371
rect 2246 2366 2252 2367
rect 2430 2371 2436 2372
rect 2430 2367 2431 2371
rect 2435 2367 2436 2371
rect 2430 2366 2436 2367
rect 2606 2371 2612 2372
rect 2606 2367 2607 2371
rect 2611 2367 2612 2371
rect 2606 2366 2612 2367
rect 2774 2371 2780 2372
rect 2774 2367 2775 2371
rect 2779 2367 2780 2371
rect 2774 2366 2780 2367
rect 2934 2371 2940 2372
rect 2934 2367 2935 2371
rect 2939 2367 2940 2371
rect 2934 2366 2940 2367
rect 3102 2371 3108 2372
rect 3102 2367 3103 2371
rect 3107 2367 3108 2371
rect 3942 2368 3943 2372
rect 3947 2368 3948 2372
rect 3942 2367 3948 2368
rect 3102 2366 3108 2367
rect 2006 2364 2012 2365
rect 110 2360 111 2364
rect 115 2360 116 2364
rect 110 2359 116 2360
rect 134 2363 140 2364
rect 134 2359 135 2363
rect 139 2359 140 2363
rect 134 2358 140 2359
rect 326 2363 332 2364
rect 326 2359 327 2363
rect 331 2359 332 2363
rect 326 2358 332 2359
rect 550 2363 556 2364
rect 550 2359 551 2363
rect 555 2359 556 2363
rect 550 2358 556 2359
rect 766 2363 772 2364
rect 766 2359 767 2363
rect 771 2359 772 2363
rect 766 2358 772 2359
rect 974 2363 980 2364
rect 974 2359 975 2363
rect 979 2359 980 2363
rect 974 2358 980 2359
rect 1174 2363 1180 2364
rect 1174 2359 1175 2363
rect 1179 2359 1180 2363
rect 1174 2358 1180 2359
rect 1366 2363 1372 2364
rect 1366 2359 1367 2363
rect 1371 2359 1372 2363
rect 1366 2358 1372 2359
rect 1550 2363 1556 2364
rect 1550 2359 1551 2363
rect 1555 2359 1556 2363
rect 1550 2358 1556 2359
rect 1734 2363 1740 2364
rect 1734 2359 1735 2363
rect 1739 2359 1740 2363
rect 1734 2358 1740 2359
rect 1902 2363 1908 2364
rect 1902 2359 1903 2363
rect 1907 2359 1908 2363
rect 2006 2360 2007 2364
rect 2011 2360 2012 2364
rect 2006 2359 2012 2360
rect 1902 2358 1908 2359
rect 2046 2355 2052 2356
rect 2046 2351 2047 2355
rect 2051 2351 2052 2355
rect 3942 2355 3948 2356
rect 2046 2350 2052 2351
rect 2070 2352 2076 2353
rect 110 2347 116 2348
rect 110 2343 111 2347
rect 115 2343 116 2347
rect 2006 2347 2012 2348
rect 110 2342 116 2343
rect 134 2344 140 2345
rect 112 2307 114 2342
rect 134 2340 135 2344
rect 139 2340 140 2344
rect 134 2339 140 2340
rect 326 2344 332 2345
rect 326 2340 327 2344
rect 331 2340 332 2344
rect 326 2339 332 2340
rect 550 2344 556 2345
rect 550 2340 551 2344
rect 555 2340 556 2344
rect 550 2339 556 2340
rect 766 2344 772 2345
rect 766 2340 767 2344
rect 771 2340 772 2344
rect 766 2339 772 2340
rect 974 2344 980 2345
rect 974 2340 975 2344
rect 979 2340 980 2344
rect 974 2339 980 2340
rect 1174 2344 1180 2345
rect 1174 2340 1175 2344
rect 1179 2340 1180 2344
rect 1174 2339 1180 2340
rect 1366 2344 1372 2345
rect 1366 2340 1367 2344
rect 1371 2340 1372 2344
rect 1366 2339 1372 2340
rect 1550 2344 1556 2345
rect 1550 2340 1551 2344
rect 1555 2340 1556 2344
rect 1550 2339 1556 2340
rect 1734 2344 1740 2345
rect 1734 2340 1735 2344
rect 1739 2340 1740 2344
rect 1734 2339 1740 2340
rect 1902 2344 1908 2345
rect 1902 2340 1903 2344
rect 1907 2340 1908 2344
rect 2006 2343 2007 2347
rect 2011 2343 2012 2347
rect 2006 2342 2012 2343
rect 1902 2339 1908 2340
rect 136 2307 138 2339
rect 328 2307 330 2339
rect 552 2307 554 2339
rect 768 2307 770 2339
rect 976 2307 978 2339
rect 1176 2307 1178 2339
rect 1368 2307 1370 2339
rect 1552 2307 1554 2339
rect 1736 2307 1738 2339
rect 1904 2307 1906 2339
rect 2008 2307 2010 2342
rect 2048 2323 2050 2350
rect 2070 2348 2071 2352
rect 2075 2348 2076 2352
rect 2070 2347 2076 2348
rect 2246 2352 2252 2353
rect 2246 2348 2247 2352
rect 2251 2348 2252 2352
rect 2246 2347 2252 2348
rect 2430 2352 2436 2353
rect 2430 2348 2431 2352
rect 2435 2348 2436 2352
rect 2430 2347 2436 2348
rect 2606 2352 2612 2353
rect 2606 2348 2607 2352
rect 2611 2348 2612 2352
rect 2606 2347 2612 2348
rect 2774 2352 2780 2353
rect 2774 2348 2775 2352
rect 2779 2348 2780 2352
rect 2774 2347 2780 2348
rect 2934 2352 2940 2353
rect 2934 2348 2935 2352
rect 2939 2348 2940 2352
rect 2934 2347 2940 2348
rect 3102 2352 3108 2353
rect 3102 2348 3103 2352
rect 3107 2348 3108 2352
rect 3942 2351 3943 2355
rect 3947 2351 3948 2355
rect 3942 2350 3948 2351
rect 3102 2347 3108 2348
rect 2072 2323 2074 2347
rect 2248 2323 2250 2347
rect 2432 2323 2434 2347
rect 2608 2323 2610 2347
rect 2776 2323 2778 2347
rect 2936 2323 2938 2347
rect 3104 2323 3106 2347
rect 3944 2323 3946 2350
rect 2047 2322 2051 2323
rect 2047 2317 2051 2318
rect 2071 2322 2075 2323
rect 2071 2317 2075 2318
rect 2175 2322 2179 2323
rect 2175 2317 2179 2318
rect 2247 2322 2251 2323
rect 2247 2317 2251 2318
rect 2311 2322 2315 2323
rect 2311 2317 2315 2318
rect 2431 2322 2435 2323
rect 2431 2317 2435 2318
rect 2447 2322 2451 2323
rect 2447 2317 2451 2318
rect 2591 2322 2595 2323
rect 2591 2317 2595 2318
rect 2607 2322 2611 2323
rect 2607 2317 2611 2318
rect 2751 2322 2755 2323
rect 2751 2317 2755 2318
rect 2775 2322 2779 2323
rect 2775 2317 2779 2318
rect 2935 2322 2939 2323
rect 2935 2317 2939 2318
rect 3103 2322 3107 2323
rect 3103 2317 3107 2318
rect 3143 2322 3147 2323
rect 3143 2317 3147 2318
rect 3375 2322 3379 2323
rect 3375 2317 3379 2318
rect 3615 2322 3619 2323
rect 3615 2317 3619 2318
rect 3839 2322 3843 2323
rect 3839 2317 3843 2318
rect 3943 2322 3947 2323
rect 3943 2317 3947 2318
rect 111 2306 115 2307
rect 111 2301 115 2302
rect 135 2306 139 2307
rect 135 2301 139 2302
rect 271 2306 275 2307
rect 271 2301 275 2302
rect 327 2306 331 2307
rect 327 2301 331 2302
rect 431 2306 435 2307
rect 431 2301 435 2302
rect 551 2306 555 2307
rect 551 2301 555 2302
rect 591 2306 595 2307
rect 591 2301 595 2302
rect 751 2306 755 2307
rect 751 2301 755 2302
rect 767 2306 771 2307
rect 767 2301 771 2302
rect 919 2306 923 2307
rect 919 2301 923 2302
rect 975 2306 979 2307
rect 975 2301 979 2302
rect 1087 2306 1091 2307
rect 1087 2301 1091 2302
rect 1175 2306 1179 2307
rect 1175 2301 1179 2302
rect 1263 2306 1267 2307
rect 1263 2301 1267 2302
rect 1367 2306 1371 2307
rect 1367 2301 1371 2302
rect 1447 2306 1451 2307
rect 1447 2301 1451 2302
rect 1551 2306 1555 2307
rect 1551 2301 1555 2302
rect 1631 2306 1635 2307
rect 1631 2301 1635 2302
rect 1735 2306 1739 2307
rect 1735 2301 1739 2302
rect 1815 2306 1819 2307
rect 1815 2301 1819 2302
rect 1903 2306 1907 2307
rect 1903 2301 1907 2302
rect 2007 2306 2011 2307
rect 2007 2301 2011 2302
rect 112 2274 114 2301
rect 136 2277 138 2301
rect 272 2277 274 2301
rect 432 2277 434 2301
rect 592 2277 594 2301
rect 752 2277 754 2301
rect 920 2277 922 2301
rect 1088 2277 1090 2301
rect 1264 2277 1266 2301
rect 1448 2277 1450 2301
rect 1632 2277 1634 2301
rect 1816 2277 1818 2301
rect 134 2276 140 2277
rect 110 2273 116 2274
rect 110 2269 111 2273
rect 115 2269 116 2273
rect 134 2272 135 2276
rect 139 2272 140 2276
rect 134 2271 140 2272
rect 270 2276 276 2277
rect 270 2272 271 2276
rect 275 2272 276 2276
rect 270 2271 276 2272
rect 430 2276 436 2277
rect 430 2272 431 2276
rect 435 2272 436 2276
rect 430 2271 436 2272
rect 590 2276 596 2277
rect 590 2272 591 2276
rect 595 2272 596 2276
rect 590 2271 596 2272
rect 750 2276 756 2277
rect 750 2272 751 2276
rect 755 2272 756 2276
rect 750 2271 756 2272
rect 918 2276 924 2277
rect 918 2272 919 2276
rect 923 2272 924 2276
rect 918 2271 924 2272
rect 1086 2276 1092 2277
rect 1086 2272 1087 2276
rect 1091 2272 1092 2276
rect 1086 2271 1092 2272
rect 1262 2276 1268 2277
rect 1262 2272 1263 2276
rect 1267 2272 1268 2276
rect 1262 2271 1268 2272
rect 1446 2276 1452 2277
rect 1446 2272 1447 2276
rect 1451 2272 1452 2276
rect 1446 2271 1452 2272
rect 1630 2276 1636 2277
rect 1630 2272 1631 2276
rect 1635 2272 1636 2276
rect 1630 2271 1636 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 2008 2274 2010 2301
rect 2048 2290 2050 2317
rect 2072 2293 2074 2317
rect 2176 2293 2178 2317
rect 2312 2293 2314 2317
rect 2448 2293 2450 2317
rect 2592 2293 2594 2317
rect 2752 2293 2754 2317
rect 2936 2293 2938 2317
rect 3144 2293 3146 2317
rect 3376 2293 3378 2317
rect 3616 2293 3618 2317
rect 3840 2293 3842 2317
rect 2070 2292 2076 2293
rect 2046 2289 2052 2290
rect 2046 2285 2047 2289
rect 2051 2285 2052 2289
rect 2070 2288 2071 2292
rect 2075 2288 2076 2292
rect 2070 2287 2076 2288
rect 2174 2292 2180 2293
rect 2174 2288 2175 2292
rect 2179 2288 2180 2292
rect 2174 2287 2180 2288
rect 2310 2292 2316 2293
rect 2310 2288 2311 2292
rect 2315 2288 2316 2292
rect 2310 2287 2316 2288
rect 2446 2292 2452 2293
rect 2446 2288 2447 2292
rect 2451 2288 2452 2292
rect 2446 2287 2452 2288
rect 2590 2292 2596 2293
rect 2590 2288 2591 2292
rect 2595 2288 2596 2292
rect 2590 2287 2596 2288
rect 2750 2292 2756 2293
rect 2750 2288 2751 2292
rect 2755 2288 2756 2292
rect 2750 2287 2756 2288
rect 2934 2292 2940 2293
rect 2934 2288 2935 2292
rect 2939 2288 2940 2292
rect 2934 2287 2940 2288
rect 3142 2292 3148 2293
rect 3142 2288 3143 2292
rect 3147 2288 3148 2292
rect 3142 2287 3148 2288
rect 3374 2292 3380 2293
rect 3374 2288 3375 2292
rect 3379 2288 3380 2292
rect 3374 2287 3380 2288
rect 3614 2292 3620 2293
rect 3614 2288 3615 2292
rect 3619 2288 3620 2292
rect 3614 2287 3620 2288
rect 3838 2292 3844 2293
rect 3838 2288 3839 2292
rect 3843 2288 3844 2292
rect 3944 2290 3946 2317
rect 3838 2287 3844 2288
rect 3942 2289 3948 2290
rect 2046 2284 2052 2285
rect 3942 2285 3943 2289
rect 3947 2285 3948 2289
rect 3942 2284 3948 2285
rect 1814 2271 1820 2272
rect 2006 2273 2012 2274
rect 2070 2273 2076 2274
rect 110 2268 116 2269
rect 2006 2269 2007 2273
rect 2011 2269 2012 2273
rect 2006 2268 2012 2269
rect 2046 2272 2052 2273
rect 2046 2268 2047 2272
rect 2051 2268 2052 2272
rect 2070 2269 2071 2273
rect 2075 2269 2076 2273
rect 2070 2268 2076 2269
rect 2174 2273 2180 2274
rect 2174 2269 2175 2273
rect 2179 2269 2180 2273
rect 2174 2268 2180 2269
rect 2310 2273 2316 2274
rect 2310 2269 2311 2273
rect 2315 2269 2316 2273
rect 2310 2268 2316 2269
rect 2446 2273 2452 2274
rect 2446 2269 2447 2273
rect 2451 2269 2452 2273
rect 2446 2268 2452 2269
rect 2590 2273 2596 2274
rect 2590 2269 2591 2273
rect 2595 2269 2596 2273
rect 2590 2268 2596 2269
rect 2750 2273 2756 2274
rect 2750 2269 2751 2273
rect 2755 2269 2756 2273
rect 2750 2268 2756 2269
rect 2934 2273 2940 2274
rect 2934 2269 2935 2273
rect 2939 2269 2940 2273
rect 2934 2268 2940 2269
rect 3142 2273 3148 2274
rect 3142 2269 3143 2273
rect 3147 2269 3148 2273
rect 3142 2268 3148 2269
rect 3374 2273 3380 2274
rect 3374 2269 3375 2273
rect 3379 2269 3380 2273
rect 3374 2268 3380 2269
rect 3614 2273 3620 2274
rect 3614 2269 3615 2273
rect 3619 2269 3620 2273
rect 3614 2268 3620 2269
rect 3838 2273 3844 2274
rect 3838 2269 3839 2273
rect 3843 2269 3844 2273
rect 3838 2268 3844 2269
rect 3942 2272 3948 2273
rect 3942 2268 3943 2272
rect 3947 2268 3948 2272
rect 2046 2267 2052 2268
rect 134 2257 140 2258
rect 110 2256 116 2257
rect 110 2252 111 2256
rect 115 2252 116 2256
rect 134 2253 135 2257
rect 139 2253 140 2257
rect 134 2252 140 2253
rect 270 2257 276 2258
rect 270 2253 271 2257
rect 275 2253 276 2257
rect 270 2252 276 2253
rect 430 2257 436 2258
rect 430 2253 431 2257
rect 435 2253 436 2257
rect 430 2252 436 2253
rect 590 2257 596 2258
rect 590 2253 591 2257
rect 595 2253 596 2257
rect 590 2252 596 2253
rect 750 2257 756 2258
rect 750 2253 751 2257
rect 755 2253 756 2257
rect 750 2252 756 2253
rect 918 2257 924 2258
rect 918 2253 919 2257
rect 923 2253 924 2257
rect 918 2252 924 2253
rect 1086 2257 1092 2258
rect 1086 2253 1087 2257
rect 1091 2253 1092 2257
rect 1086 2252 1092 2253
rect 1262 2257 1268 2258
rect 1262 2253 1263 2257
rect 1267 2253 1268 2257
rect 1262 2252 1268 2253
rect 1446 2257 1452 2258
rect 1446 2253 1447 2257
rect 1451 2253 1452 2257
rect 1446 2252 1452 2253
rect 1630 2257 1636 2258
rect 1630 2253 1631 2257
rect 1635 2253 1636 2257
rect 1630 2252 1636 2253
rect 1814 2257 1820 2258
rect 1814 2253 1815 2257
rect 1819 2253 1820 2257
rect 1814 2252 1820 2253
rect 2006 2256 2012 2257
rect 2006 2252 2007 2256
rect 2011 2252 2012 2256
rect 110 2251 116 2252
rect 112 2231 114 2251
rect 136 2231 138 2252
rect 272 2231 274 2252
rect 432 2231 434 2252
rect 592 2231 594 2252
rect 752 2231 754 2252
rect 920 2231 922 2252
rect 1088 2231 1090 2252
rect 1264 2231 1266 2252
rect 1448 2231 1450 2252
rect 1632 2231 1634 2252
rect 1816 2231 1818 2252
rect 2006 2251 2012 2252
rect 2008 2231 2010 2251
rect 2048 2239 2050 2267
rect 2072 2239 2074 2268
rect 2176 2239 2178 2268
rect 2312 2239 2314 2268
rect 2448 2239 2450 2268
rect 2592 2239 2594 2268
rect 2752 2239 2754 2268
rect 2936 2239 2938 2268
rect 3144 2239 3146 2268
rect 3376 2239 3378 2268
rect 3616 2239 3618 2268
rect 3840 2239 3842 2268
rect 3942 2267 3948 2268
rect 3944 2239 3946 2267
rect 2047 2238 2051 2239
rect 2047 2233 2051 2234
rect 2071 2238 2075 2239
rect 2071 2233 2075 2234
rect 2111 2238 2115 2239
rect 2111 2233 2115 2234
rect 2175 2238 2179 2239
rect 2175 2233 2179 2234
rect 2255 2238 2259 2239
rect 2255 2233 2259 2234
rect 2311 2238 2315 2239
rect 2311 2233 2315 2234
rect 2407 2238 2411 2239
rect 2407 2233 2411 2234
rect 2447 2238 2451 2239
rect 2447 2233 2451 2234
rect 2559 2238 2563 2239
rect 2559 2233 2563 2234
rect 2591 2238 2595 2239
rect 2591 2233 2595 2234
rect 2719 2238 2723 2239
rect 2719 2233 2723 2234
rect 2751 2238 2755 2239
rect 2751 2233 2755 2234
rect 2879 2238 2883 2239
rect 2879 2233 2883 2234
rect 2935 2238 2939 2239
rect 2935 2233 2939 2234
rect 3047 2238 3051 2239
rect 3047 2233 3051 2234
rect 3143 2238 3147 2239
rect 3143 2233 3147 2234
rect 3223 2238 3227 2239
rect 3223 2233 3227 2234
rect 3375 2238 3379 2239
rect 3375 2233 3379 2234
rect 3407 2238 3411 2239
rect 3407 2233 3411 2234
rect 3591 2238 3595 2239
rect 3591 2233 3595 2234
rect 3615 2238 3619 2239
rect 3615 2233 3619 2234
rect 3783 2238 3787 2239
rect 3783 2233 3787 2234
rect 3839 2238 3843 2239
rect 3839 2233 3843 2234
rect 3943 2238 3947 2239
rect 3943 2233 3947 2234
rect 111 2230 115 2231
rect 111 2225 115 2226
rect 135 2230 139 2231
rect 135 2225 139 2226
rect 159 2230 163 2231
rect 159 2225 163 2226
rect 271 2230 275 2231
rect 271 2225 275 2226
rect 327 2230 331 2231
rect 327 2225 331 2226
rect 431 2230 435 2231
rect 431 2225 435 2226
rect 495 2230 499 2231
rect 495 2225 499 2226
rect 591 2230 595 2231
rect 591 2225 595 2226
rect 679 2230 683 2231
rect 679 2225 683 2226
rect 751 2230 755 2231
rect 751 2225 755 2226
rect 879 2230 883 2231
rect 879 2225 883 2226
rect 919 2230 923 2231
rect 919 2225 923 2226
rect 1087 2230 1091 2231
rect 1087 2225 1091 2226
rect 1095 2230 1099 2231
rect 1095 2225 1099 2226
rect 1263 2230 1267 2231
rect 1263 2225 1267 2226
rect 1327 2230 1331 2231
rect 1327 2225 1331 2226
rect 1447 2230 1451 2231
rect 1447 2225 1451 2226
rect 1567 2230 1571 2231
rect 1567 2225 1571 2226
rect 1631 2230 1635 2231
rect 1631 2225 1635 2226
rect 1815 2230 1819 2231
rect 1815 2225 1819 2226
rect 2007 2230 2011 2231
rect 2007 2225 2011 2226
rect 112 2205 114 2225
rect 110 2204 116 2205
rect 160 2204 162 2225
rect 328 2204 330 2225
rect 496 2204 498 2225
rect 680 2204 682 2225
rect 880 2204 882 2225
rect 1096 2204 1098 2225
rect 1328 2204 1330 2225
rect 1568 2204 1570 2225
rect 1816 2204 1818 2225
rect 2008 2205 2010 2225
rect 2048 2213 2050 2233
rect 2046 2212 2052 2213
rect 2112 2212 2114 2233
rect 2256 2212 2258 2233
rect 2408 2212 2410 2233
rect 2560 2212 2562 2233
rect 2720 2212 2722 2233
rect 2880 2212 2882 2233
rect 3048 2212 3050 2233
rect 3224 2212 3226 2233
rect 3408 2212 3410 2233
rect 3592 2212 3594 2233
rect 3784 2212 3786 2233
rect 3944 2213 3946 2233
rect 3942 2212 3948 2213
rect 2046 2208 2047 2212
rect 2051 2208 2052 2212
rect 2046 2207 2052 2208
rect 2110 2211 2116 2212
rect 2110 2207 2111 2211
rect 2115 2207 2116 2211
rect 2110 2206 2116 2207
rect 2254 2211 2260 2212
rect 2254 2207 2255 2211
rect 2259 2207 2260 2211
rect 2254 2206 2260 2207
rect 2406 2211 2412 2212
rect 2406 2207 2407 2211
rect 2411 2207 2412 2211
rect 2406 2206 2412 2207
rect 2558 2211 2564 2212
rect 2558 2207 2559 2211
rect 2563 2207 2564 2211
rect 2558 2206 2564 2207
rect 2718 2211 2724 2212
rect 2718 2207 2719 2211
rect 2723 2207 2724 2211
rect 2718 2206 2724 2207
rect 2878 2211 2884 2212
rect 2878 2207 2879 2211
rect 2883 2207 2884 2211
rect 2878 2206 2884 2207
rect 3046 2211 3052 2212
rect 3046 2207 3047 2211
rect 3051 2207 3052 2211
rect 3046 2206 3052 2207
rect 3222 2211 3228 2212
rect 3222 2207 3223 2211
rect 3227 2207 3228 2211
rect 3222 2206 3228 2207
rect 3406 2211 3412 2212
rect 3406 2207 3407 2211
rect 3411 2207 3412 2211
rect 3406 2206 3412 2207
rect 3590 2211 3596 2212
rect 3590 2207 3591 2211
rect 3595 2207 3596 2211
rect 3590 2206 3596 2207
rect 3782 2211 3788 2212
rect 3782 2207 3783 2211
rect 3787 2207 3788 2211
rect 3942 2208 3943 2212
rect 3947 2208 3948 2212
rect 3942 2207 3948 2208
rect 3782 2206 3788 2207
rect 2006 2204 2012 2205
rect 110 2200 111 2204
rect 115 2200 116 2204
rect 110 2199 116 2200
rect 158 2203 164 2204
rect 158 2199 159 2203
rect 163 2199 164 2203
rect 158 2198 164 2199
rect 326 2203 332 2204
rect 326 2199 327 2203
rect 331 2199 332 2203
rect 326 2198 332 2199
rect 494 2203 500 2204
rect 494 2199 495 2203
rect 499 2199 500 2203
rect 494 2198 500 2199
rect 678 2203 684 2204
rect 678 2199 679 2203
rect 683 2199 684 2203
rect 678 2198 684 2199
rect 878 2203 884 2204
rect 878 2199 879 2203
rect 883 2199 884 2203
rect 878 2198 884 2199
rect 1094 2203 1100 2204
rect 1094 2199 1095 2203
rect 1099 2199 1100 2203
rect 1094 2198 1100 2199
rect 1326 2203 1332 2204
rect 1326 2199 1327 2203
rect 1331 2199 1332 2203
rect 1326 2198 1332 2199
rect 1566 2203 1572 2204
rect 1566 2199 1567 2203
rect 1571 2199 1572 2203
rect 1566 2198 1572 2199
rect 1814 2203 1820 2204
rect 1814 2199 1815 2203
rect 1819 2199 1820 2203
rect 2006 2200 2007 2204
rect 2011 2200 2012 2204
rect 2006 2199 2012 2200
rect 1814 2198 1820 2199
rect 2046 2195 2052 2196
rect 2046 2191 2047 2195
rect 2051 2191 2052 2195
rect 3942 2195 3948 2196
rect 2046 2190 2052 2191
rect 2110 2192 2116 2193
rect 110 2187 116 2188
rect 110 2183 111 2187
rect 115 2183 116 2187
rect 2006 2187 2012 2188
rect 110 2182 116 2183
rect 158 2184 164 2185
rect 112 2155 114 2182
rect 158 2180 159 2184
rect 163 2180 164 2184
rect 158 2179 164 2180
rect 326 2184 332 2185
rect 326 2180 327 2184
rect 331 2180 332 2184
rect 326 2179 332 2180
rect 494 2184 500 2185
rect 494 2180 495 2184
rect 499 2180 500 2184
rect 494 2179 500 2180
rect 678 2184 684 2185
rect 678 2180 679 2184
rect 683 2180 684 2184
rect 678 2179 684 2180
rect 878 2184 884 2185
rect 878 2180 879 2184
rect 883 2180 884 2184
rect 878 2179 884 2180
rect 1094 2184 1100 2185
rect 1094 2180 1095 2184
rect 1099 2180 1100 2184
rect 1094 2179 1100 2180
rect 1326 2184 1332 2185
rect 1326 2180 1327 2184
rect 1331 2180 1332 2184
rect 1326 2179 1332 2180
rect 1566 2184 1572 2185
rect 1566 2180 1567 2184
rect 1571 2180 1572 2184
rect 1566 2179 1572 2180
rect 1814 2184 1820 2185
rect 1814 2180 1815 2184
rect 1819 2180 1820 2184
rect 2006 2183 2007 2187
rect 2011 2183 2012 2187
rect 2006 2182 2012 2183
rect 1814 2179 1820 2180
rect 160 2155 162 2179
rect 328 2155 330 2179
rect 496 2155 498 2179
rect 680 2155 682 2179
rect 880 2155 882 2179
rect 1096 2155 1098 2179
rect 1328 2155 1330 2179
rect 1568 2155 1570 2179
rect 1816 2155 1818 2179
rect 2008 2155 2010 2182
rect 111 2154 115 2155
rect 111 2149 115 2150
rect 159 2154 163 2155
rect 159 2149 163 2150
rect 223 2154 227 2155
rect 223 2149 227 2150
rect 327 2154 331 2155
rect 327 2149 331 2150
rect 359 2154 363 2155
rect 359 2149 363 2150
rect 495 2154 499 2155
rect 495 2149 499 2150
rect 639 2154 643 2155
rect 639 2149 643 2150
rect 679 2154 683 2155
rect 679 2149 683 2150
rect 783 2154 787 2155
rect 783 2149 787 2150
rect 879 2154 883 2155
rect 879 2149 883 2150
rect 935 2154 939 2155
rect 935 2149 939 2150
rect 1095 2154 1099 2155
rect 1095 2149 1099 2150
rect 1263 2154 1267 2155
rect 1263 2149 1267 2150
rect 1327 2154 1331 2155
rect 1327 2149 1331 2150
rect 1447 2154 1451 2155
rect 1447 2149 1451 2150
rect 1567 2154 1571 2155
rect 1567 2149 1571 2150
rect 1631 2154 1635 2155
rect 1631 2149 1635 2150
rect 1815 2154 1819 2155
rect 1815 2149 1819 2150
rect 1823 2154 1827 2155
rect 1823 2149 1827 2150
rect 2007 2154 2011 2155
rect 2048 2151 2050 2190
rect 2110 2188 2111 2192
rect 2115 2188 2116 2192
rect 2110 2187 2116 2188
rect 2254 2192 2260 2193
rect 2254 2188 2255 2192
rect 2259 2188 2260 2192
rect 2254 2187 2260 2188
rect 2406 2192 2412 2193
rect 2406 2188 2407 2192
rect 2411 2188 2412 2192
rect 2406 2187 2412 2188
rect 2558 2192 2564 2193
rect 2558 2188 2559 2192
rect 2563 2188 2564 2192
rect 2558 2187 2564 2188
rect 2718 2192 2724 2193
rect 2718 2188 2719 2192
rect 2723 2188 2724 2192
rect 2718 2187 2724 2188
rect 2878 2192 2884 2193
rect 2878 2188 2879 2192
rect 2883 2188 2884 2192
rect 2878 2187 2884 2188
rect 3046 2192 3052 2193
rect 3046 2188 3047 2192
rect 3051 2188 3052 2192
rect 3046 2187 3052 2188
rect 3222 2192 3228 2193
rect 3222 2188 3223 2192
rect 3227 2188 3228 2192
rect 3222 2187 3228 2188
rect 3406 2192 3412 2193
rect 3406 2188 3407 2192
rect 3411 2188 3412 2192
rect 3406 2187 3412 2188
rect 3590 2192 3596 2193
rect 3590 2188 3591 2192
rect 3595 2188 3596 2192
rect 3590 2187 3596 2188
rect 3782 2192 3788 2193
rect 3782 2188 3783 2192
rect 3787 2188 3788 2192
rect 3942 2191 3943 2195
rect 3947 2191 3948 2195
rect 3942 2190 3948 2191
rect 3782 2187 3788 2188
rect 2112 2151 2114 2187
rect 2256 2151 2258 2187
rect 2408 2151 2410 2187
rect 2560 2151 2562 2187
rect 2720 2151 2722 2187
rect 2880 2151 2882 2187
rect 3048 2151 3050 2187
rect 3224 2151 3226 2187
rect 3408 2151 3410 2187
rect 3592 2151 3594 2187
rect 3784 2151 3786 2187
rect 3944 2151 3946 2190
rect 2007 2149 2011 2150
rect 2047 2150 2051 2151
rect 112 2122 114 2149
rect 224 2125 226 2149
rect 360 2125 362 2149
rect 496 2125 498 2149
rect 640 2125 642 2149
rect 784 2125 786 2149
rect 936 2125 938 2149
rect 1096 2125 1098 2149
rect 1264 2125 1266 2149
rect 1448 2125 1450 2149
rect 1632 2125 1634 2149
rect 1824 2125 1826 2149
rect 222 2124 228 2125
rect 110 2121 116 2122
rect 110 2117 111 2121
rect 115 2117 116 2121
rect 222 2120 223 2124
rect 227 2120 228 2124
rect 222 2119 228 2120
rect 358 2124 364 2125
rect 358 2120 359 2124
rect 363 2120 364 2124
rect 358 2119 364 2120
rect 494 2124 500 2125
rect 494 2120 495 2124
rect 499 2120 500 2124
rect 494 2119 500 2120
rect 638 2124 644 2125
rect 638 2120 639 2124
rect 643 2120 644 2124
rect 638 2119 644 2120
rect 782 2124 788 2125
rect 782 2120 783 2124
rect 787 2120 788 2124
rect 782 2119 788 2120
rect 934 2124 940 2125
rect 934 2120 935 2124
rect 939 2120 940 2124
rect 934 2119 940 2120
rect 1094 2124 1100 2125
rect 1094 2120 1095 2124
rect 1099 2120 1100 2124
rect 1094 2119 1100 2120
rect 1262 2124 1268 2125
rect 1262 2120 1263 2124
rect 1267 2120 1268 2124
rect 1262 2119 1268 2120
rect 1446 2124 1452 2125
rect 1446 2120 1447 2124
rect 1451 2120 1452 2124
rect 1446 2119 1452 2120
rect 1630 2124 1636 2125
rect 1630 2120 1631 2124
rect 1635 2120 1636 2124
rect 1630 2119 1636 2120
rect 1822 2124 1828 2125
rect 1822 2120 1823 2124
rect 1827 2120 1828 2124
rect 2008 2122 2010 2149
rect 2047 2145 2051 2146
rect 2111 2150 2115 2151
rect 2111 2145 2115 2146
rect 2255 2150 2259 2151
rect 2255 2145 2259 2146
rect 2287 2150 2291 2151
rect 2287 2145 2291 2146
rect 2407 2150 2411 2151
rect 2407 2145 2411 2146
rect 2431 2150 2435 2151
rect 2431 2145 2435 2146
rect 2559 2150 2563 2151
rect 2559 2145 2563 2146
rect 2583 2150 2587 2151
rect 2583 2145 2587 2146
rect 2719 2150 2723 2151
rect 2719 2145 2723 2146
rect 2735 2150 2739 2151
rect 2735 2145 2739 2146
rect 2879 2150 2883 2151
rect 2879 2145 2883 2146
rect 2887 2150 2891 2151
rect 2887 2145 2891 2146
rect 3047 2150 3051 2151
rect 3047 2145 3051 2146
rect 3207 2150 3211 2151
rect 3207 2145 3211 2146
rect 3223 2150 3227 2151
rect 3223 2145 3227 2146
rect 3367 2150 3371 2151
rect 3367 2145 3371 2146
rect 3407 2150 3411 2151
rect 3407 2145 3411 2146
rect 3527 2150 3531 2151
rect 3527 2145 3531 2146
rect 3591 2150 3595 2151
rect 3591 2145 3595 2146
rect 3695 2150 3699 2151
rect 3695 2145 3699 2146
rect 3783 2150 3787 2151
rect 3783 2145 3787 2146
rect 3839 2150 3843 2151
rect 3839 2145 3843 2146
rect 3943 2150 3947 2151
rect 3943 2145 3947 2146
rect 1822 2119 1828 2120
rect 2006 2121 2012 2122
rect 110 2116 116 2117
rect 2006 2117 2007 2121
rect 2011 2117 2012 2121
rect 2048 2118 2050 2145
rect 2288 2121 2290 2145
rect 2432 2121 2434 2145
rect 2584 2121 2586 2145
rect 2736 2121 2738 2145
rect 2888 2121 2890 2145
rect 3048 2121 3050 2145
rect 3208 2121 3210 2145
rect 3368 2121 3370 2145
rect 3528 2121 3530 2145
rect 3696 2121 3698 2145
rect 3840 2121 3842 2145
rect 2286 2120 2292 2121
rect 2006 2116 2012 2117
rect 2046 2117 2052 2118
rect 2046 2113 2047 2117
rect 2051 2113 2052 2117
rect 2286 2116 2287 2120
rect 2291 2116 2292 2120
rect 2286 2115 2292 2116
rect 2430 2120 2436 2121
rect 2430 2116 2431 2120
rect 2435 2116 2436 2120
rect 2430 2115 2436 2116
rect 2582 2120 2588 2121
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2582 2115 2588 2116
rect 2734 2120 2740 2121
rect 2734 2116 2735 2120
rect 2739 2116 2740 2120
rect 2734 2115 2740 2116
rect 2886 2120 2892 2121
rect 2886 2116 2887 2120
rect 2891 2116 2892 2120
rect 2886 2115 2892 2116
rect 3046 2120 3052 2121
rect 3046 2116 3047 2120
rect 3051 2116 3052 2120
rect 3046 2115 3052 2116
rect 3206 2120 3212 2121
rect 3206 2116 3207 2120
rect 3211 2116 3212 2120
rect 3206 2115 3212 2116
rect 3366 2120 3372 2121
rect 3366 2116 3367 2120
rect 3371 2116 3372 2120
rect 3366 2115 3372 2116
rect 3526 2120 3532 2121
rect 3526 2116 3527 2120
rect 3531 2116 3532 2120
rect 3526 2115 3532 2116
rect 3694 2120 3700 2121
rect 3694 2116 3695 2120
rect 3699 2116 3700 2120
rect 3694 2115 3700 2116
rect 3838 2120 3844 2121
rect 3838 2116 3839 2120
rect 3843 2116 3844 2120
rect 3944 2118 3946 2145
rect 3838 2115 3844 2116
rect 3942 2117 3948 2118
rect 2046 2112 2052 2113
rect 3942 2113 3943 2117
rect 3947 2113 3948 2117
rect 3942 2112 3948 2113
rect 222 2105 228 2106
rect 110 2104 116 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 222 2101 223 2105
rect 227 2101 228 2105
rect 222 2100 228 2101
rect 358 2105 364 2106
rect 358 2101 359 2105
rect 363 2101 364 2105
rect 358 2100 364 2101
rect 494 2105 500 2106
rect 494 2101 495 2105
rect 499 2101 500 2105
rect 494 2100 500 2101
rect 638 2105 644 2106
rect 638 2101 639 2105
rect 643 2101 644 2105
rect 638 2100 644 2101
rect 782 2105 788 2106
rect 782 2101 783 2105
rect 787 2101 788 2105
rect 782 2100 788 2101
rect 934 2105 940 2106
rect 934 2101 935 2105
rect 939 2101 940 2105
rect 934 2100 940 2101
rect 1094 2105 1100 2106
rect 1094 2101 1095 2105
rect 1099 2101 1100 2105
rect 1094 2100 1100 2101
rect 1262 2105 1268 2106
rect 1262 2101 1263 2105
rect 1267 2101 1268 2105
rect 1262 2100 1268 2101
rect 1446 2105 1452 2106
rect 1446 2101 1447 2105
rect 1451 2101 1452 2105
rect 1446 2100 1452 2101
rect 1630 2105 1636 2106
rect 1630 2101 1631 2105
rect 1635 2101 1636 2105
rect 1630 2100 1636 2101
rect 1822 2105 1828 2106
rect 1822 2101 1823 2105
rect 1827 2101 1828 2105
rect 1822 2100 1828 2101
rect 2006 2104 2012 2105
rect 2006 2100 2007 2104
rect 2011 2100 2012 2104
rect 2286 2101 2292 2102
rect 110 2099 116 2100
rect 112 2071 114 2099
rect 224 2071 226 2100
rect 360 2071 362 2100
rect 496 2071 498 2100
rect 640 2071 642 2100
rect 784 2071 786 2100
rect 936 2071 938 2100
rect 1096 2071 1098 2100
rect 1264 2071 1266 2100
rect 1448 2071 1450 2100
rect 1632 2071 1634 2100
rect 1824 2071 1826 2100
rect 2006 2099 2012 2100
rect 2046 2100 2052 2101
rect 2008 2071 2010 2099
rect 2046 2096 2047 2100
rect 2051 2096 2052 2100
rect 2286 2097 2287 2101
rect 2291 2097 2292 2101
rect 2286 2096 2292 2097
rect 2430 2101 2436 2102
rect 2430 2097 2431 2101
rect 2435 2097 2436 2101
rect 2430 2096 2436 2097
rect 2582 2101 2588 2102
rect 2582 2097 2583 2101
rect 2587 2097 2588 2101
rect 2582 2096 2588 2097
rect 2734 2101 2740 2102
rect 2734 2097 2735 2101
rect 2739 2097 2740 2101
rect 2734 2096 2740 2097
rect 2886 2101 2892 2102
rect 2886 2097 2887 2101
rect 2891 2097 2892 2101
rect 2886 2096 2892 2097
rect 3046 2101 3052 2102
rect 3046 2097 3047 2101
rect 3051 2097 3052 2101
rect 3046 2096 3052 2097
rect 3206 2101 3212 2102
rect 3206 2097 3207 2101
rect 3211 2097 3212 2101
rect 3206 2096 3212 2097
rect 3366 2101 3372 2102
rect 3366 2097 3367 2101
rect 3371 2097 3372 2101
rect 3366 2096 3372 2097
rect 3526 2101 3532 2102
rect 3526 2097 3527 2101
rect 3531 2097 3532 2101
rect 3526 2096 3532 2097
rect 3694 2101 3700 2102
rect 3694 2097 3695 2101
rect 3699 2097 3700 2101
rect 3694 2096 3700 2097
rect 3838 2101 3844 2102
rect 3838 2097 3839 2101
rect 3843 2097 3844 2101
rect 3838 2096 3844 2097
rect 3942 2100 3948 2101
rect 3942 2096 3943 2100
rect 3947 2096 3948 2100
rect 2046 2095 2052 2096
rect 111 2070 115 2071
rect 111 2065 115 2066
rect 223 2070 227 2071
rect 223 2065 227 2066
rect 359 2070 363 2071
rect 359 2065 363 2066
rect 375 2070 379 2071
rect 375 2065 379 2066
rect 495 2070 499 2071
rect 495 2065 499 2066
rect 615 2070 619 2071
rect 615 2065 619 2066
rect 639 2070 643 2071
rect 639 2065 643 2066
rect 751 2070 755 2071
rect 751 2065 755 2066
rect 783 2070 787 2071
rect 783 2065 787 2066
rect 895 2070 899 2071
rect 895 2065 899 2066
rect 935 2070 939 2071
rect 935 2065 939 2066
rect 1047 2070 1051 2071
rect 1047 2065 1051 2066
rect 1095 2070 1099 2071
rect 1095 2065 1099 2066
rect 1215 2070 1219 2071
rect 1215 2065 1219 2066
rect 1263 2070 1267 2071
rect 1263 2065 1267 2066
rect 1399 2070 1403 2071
rect 1399 2065 1403 2066
rect 1447 2070 1451 2071
rect 1447 2065 1451 2066
rect 1583 2070 1587 2071
rect 1583 2065 1587 2066
rect 1631 2070 1635 2071
rect 1631 2065 1635 2066
rect 1775 2070 1779 2071
rect 1775 2065 1779 2066
rect 1823 2070 1827 2071
rect 1823 2065 1827 2066
rect 2007 2070 2011 2071
rect 2048 2067 2050 2095
rect 2288 2067 2290 2096
rect 2432 2067 2434 2096
rect 2584 2067 2586 2096
rect 2736 2067 2738 2096
rect 2888 2067 2890 2096
rect 3048 2067 3050 2096
rect 3208 2067 3210 2096
rect 3368 2067 3370 2096
rect 3528 2067 3530 2096
rect 3696 2067 3698 2096
rect 3840 2067 3842 2096
rect 3942 2095 3948 2096
rect 3944 2067 3946 2095
rect 2007 2065 2011 2066
rect 2047 2066 2051 2067
rect 112 2045 114 2065
rect 110 2044 116 2045
rect 376 2044 378 2065
rect 496 2044 498 2065
rect 616 2044 618 2065
rect 752 2044 754 2065
rect 896 2044 898 2065
rect 1048 2044 1050 2065
rect 1216 2044 1218 2065
rect 1400 2044 1402 2065
rect 1584 2044 1586 2065
rect 1776 2044 1778 2065
rect 2008 2045 2010 2065
rect 2047 2061 2051 2062
rect 2287 2066 2291 2067
rect 2287 2061 2291 2062
rect 2431 2066 2435 2067
rect 2431 2061 2435 2062
rect 2503 2066 2507 2067
rect 2503 2061 2507 2062
rect 2583 2066 2587 2067
rect 2583 2061 2587 2062
rect 2671 2066 2675 2067
rect 2671 2061 2675 2062
rect 2735 2066 2739 2067
rect 2735 2061 2739 2062
rect 2839 2066 2843 2067
rect 2839 2061 2843 2062
rect 2887 2066 2891 2067
rect 2887 2061 2891 2062
rect 3007 2066 3011 2067
rect 3007 2061 3011 2062
rect 3047 2066 3051 2067
rect 3047 2061 3051 2062
rect 3167 2066 3171 2067
rect 3167 2061 3171 2062
rect 3207 2066 3211 2067
rect 3207 2061 3211 2062
rect 3311 2066 3315 2067
rect 3311 2061 3315 2062
rect 3367 2066 3371 2067
rect 3367 2061 3371 2062
rect 3455 2066 3459 2067
rect 3455 2061 3459 2062
rect 3527 2066 3531 2067
rect 3527 2061 3531 2062
rect 3591 2066 3595 2067
rect 3591 2061 3595 2062
rect 3695 2066 3699 2067
rect 3695 2061 3699 2062
rect 3727 2066 3731 2067
rect 3727 2061 3731 2062
rect 3839 2066 3843 2067
rect 3839 2061 3843 2062
rect 3943 2066 3947 2067
rect 3943 2061 3947 2062
rect 2006 2044 2012 2045
rect 110 2040 111 2044
rect 115 2040 116 2044
rect 110 2039 116 2040
rect 374 2043 380 2044
rect 374 2039 375 2043
rect 379 2039 380 2043
rect 374 2038 380 2039
rect 494 2043 500 2044
rect 494 2039 495 2043
rect 499 2039 500 2043
rect 494 2038 500 2039
rect 614 2043 620 2044
rect 614 2039 615 2043
rect 619 2039 620 2043
rect 614 2038 620 2039
rect 750 2043 756 2044
rect 750 2039 751 2043
rect 755 2039 756 2043
rect 750 2038 756 2039
rect 894 2043 900 2044
rect 894 2039 895 2043
rect 899 2039 900 2043
rect 894 2038 900 2039
rect 1046 2043 1052 2044
rect 1046 2039 1047 2043
rect 1051 2039 1052 2043
rect 1046 2038 1052 2039
rect 1214 2043 1220 2044
rect 1214 2039 1215 2043
rect 1219 2039 1220 2043
rect 1214 2038 1220 2039
rect 1398 2043 1404 2044
rect 1398 2039 1399 2043
rect 1403 2039 1404 2043
rect 1398 2038 1404 2039
rect 1582 2043 1588 2044
rect 1582 2039 1583 2043
rect 1587 2039 1588 2043
rect 1582 2038 1588 2039
rect 1774 2043 1780 2044
rect 1774 2039 1775 2043
rect 1779 2039 1780 2043
rect 2006 2040 2007 2044
rect 2011 2040 2012 2044
rect 2048 2041 2050 2061
rect 2006 2039 2012 2040
rect 2046 2040 2052 2041
rect 2504 2040 2506 2061
rect 2672 2040 2674 2061
rect 2840 2040 2842 2061
rect 3008 2040 3010 2061
rect 3168 2040 3170 2061
rect 3312 2040 3314 2061
rect 3456 2040 3458 2061
rect 3592 2040 3594 2061
rect 3728 2040 3730 2061
rect 3840 2040 3842 2061
rect 3944 2041 3946 2061
rect 3942 2040 3948 2041
rect 1774 2038 1780 2039
rect 2046 2036 2047 2040
rect 2051 2036 2052 2040
rect 2046 2035 2052 2036
rect 2502 2039 2508 2040
rect 2502 2035 2503 2039
rect 2507 2035 2508 2039
rect 2502 2034 2508 2035
rect 2670 2039 2676 2040
rect 2670 2035 2671 2039
rect 2675 2035 2676 2039
rect 2670 2034 2676 2035
rect 2838 2039 2844 2040
rect 2838 2035 2839 2039
rect 2843 2035 2844 2039
rect 2838 2034 2844 2035
rect 3006 2039 3012 2040
rect 3006 2035 3007 2039
rect 3011 2035 3012 2039
rect 3006 2034 3012 2035
rect 3166 2039 3172 2040
rect 3166 2035 3167 2039
rect 3171 2035 3172 2039
rect 3166 2034 3172 2035
rect 3310 2039 3316 2040
rect 3310 2035 3311 2039
rect 3315 2035 3316 2039
rect 3310 2034 3316 2035
rect 3454 2039 3460 2040
rect 3454 2035 3455 2039
rect 3459 2035 3460 2039
rect 3454 2034 3460 2035
rect 3590 2039 3596 2040
rect 3590 2035 3591 2039
rect 3595 2035 3596 2039
rect 3590 2034 3596 2035
rect 3726 2039 3732 2040
rect 3726 2035 3727 2039
rect 3731 2035 3732 2039
rect 3726 2034 3732 2035
rect 3838 2039 3844 2040
rect 3838 2035 3839 2039
rect 3843 2035 3844 2039
rect 3942 2036 3943 2040
rect 3947 2036 3948 2040
rect 3942 2035 3948 2036
rect 3838 2034 3844 2035
rect 110 2027 116 2028
rect 110 2023 111 2027
rect 115 2023 116 2027
rect 2006 2027 2012 2028
rect 110 2022 116 2023
rect 374 2024 380 2025
rect 112 1987 114 2022
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 494 2024 500 2025
rect 494 2020 495 2024
rect 499 2020 500 2024
rect 494 2019 500 2020
rect 614 2024 620 2025
rect 614 2020 615 2024
rect 619 2020 620 2024
rect 614 2019 620 2020
rect 750 2024 756 2025
rect 750 2020 751 2024
rect 755 2020 756 2024
rect 750 2019 756 2020
rect 894 2024 900 2025
rect 894 2020 895 2024
rect 899 2020 900 2024
rect 894 2019 900 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1214 2024 1220 2025
rect 1214 2020 1215 2024
rect 1219 2020 1220 2024
rect 1214 2019 1220 2020
rect 1398 2024 1404 2025
rect 1398 2020 1399 2024
rect 1403 2020 1404 2024
rect 1398 2019 1404 2020
rect 1582 2024 1588 2025
rect 1582 2020 1583 2024
rect 1587 2020 1588 2024
rect 1582 2019 1588 2020
rect 1774 2024 1780 2025
rect 1774 2020 1775 2024
rect 1779 2020 1780 2024
rect 2006 2023 2007 2027
rect 2011 2023 2012 2027
rect 2006 2022 2012 2023
rect 2046 2023 2052 2024
rect 1774 2019 1780 2020
rect 376 1987 378 2019
rect 496 1987 498 2019
rect 616 1987 618 2019
rect 752 1987 754 2019
rect 896 1987 898 2019
rect 1048 1987 1050 2019
rect 1216 1987 1218 2019
rect 1400 1987 1402 2019
rect 1584 1987 1586 2019
rect 1776 1987 1778 2019
rect 2008 1987 2010 2022
rect 2046 2019 2047 2023
rect 2051 2019 2052 2023
rect 3942 2023 3948 2024
rect 2046 2018 2052 2019
rect 2502 2020 2508 2021
rect 2048 1987 2050 2018
rect 2502 2016 2503 2020
rect 2507 2016 2508 2020
rect 2502 2015 2508 2016
rect 2670 2020 2676 2021
rect 2670 2016 2671 2020
rect 2675 2016 2676 2020
rect 2670 2015 2676 2016
rect 2838 2020 2844 2021
rect 2838 2016 2839 2020
rect 2843 2016 2844 2020
rect 2838 2015 2844 2016
rect 3006 2020 3012 2021
rect 3006 2016 3007 2020
rect 3011 2016 3012 2020
rect 3006 2015 3012 2016
rect 3166 2020 3172 2021
rect 3166 2016 3167 2020
rect 3171 2016 3172 2020
rect 3166 2015 3172 2016
rect 3310 2020 3316 2021
rect 3310 2016 3311 2020
rect 3315 2016 3316 2020
rect 3310 2015 3316 2016
rect 3454 2020 3460 2021
rect 3454 2016 3455 2020
rect 3459 2016 3460 2020
rect 3454 2015 3460 2016
rect 3590 2020 3596 2021
rect 3590 2016 3591 2020
rect 3595 2016 3596 2020
rect 3590 2015 3596 2016
rect 3726 2020 3732 2021
rect 3726 2016 3727 2020
rect 3731 2016 3732 2020
rect 3726 2015 3732 2016
rect 3838 2020 3844 2021
rect 3838 2016 3839 2020
rect 3843 2016 3844 2020
rect 3942 2019 3943 2023
rect 3947 2019 3948 2023
rect 3942 2018 3948 2019
rect 3838 2015 3844 2016
rect 2504 1987 2506 2015
rect 2672 1987 2674 2015
rect 2840 1987 2842 2015
rect 3008 1987 3010 2015
rect 3168 1987 3170 2015
rect 3312 1987 3314 2015
rect 3456 1987 3458 2015
rect 3592 1987 3594 2015
rect 3728 1987 3730 2015
rect 3840 1987 3842 2015
rect 3944 1987 3946 2018
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 375 1986 379 1987
rect 375 1981 379 1982
rect 495 1986 499 1987
rect 495 1981 499 1982
rect 511 1986 515 1987
rect 511 1981 515 1982
rect 615 1986 619 1987
rect 615 1981 619 1982
rect 623 1986 627 1987
rect 623 1981 627 1982
rect 743 1986 747 1987
rect 743 1981 747 1982
rect 751 1986 755 1987
rect 751 1981 755 1982
rect 871 1986 875 1987
rect 871 1981 875 1982
rect 895 1986 899 1987
rect 895 1981 899 1982
rect 1007 1986 1011 1987
rect 1007 1981 1011 1982
rect 1047 1986 1051 1987
rect 1047 1981 1051 1982
rect 1143 1986 1147 1987
rect 1143 1981 1147 1982
rect 1215 1986 1219 1987
rect 1215 1981 1219 1982
rect 1279 1986 1283 1987
rect 1279 1981 1283 1982
rect 1399 1986 1403 1987
rect 1399 1981 1403 1982
rect 1415 1986 1419 1987
rect 1415 1981 1419 1982
rect 1559 1986 1563 1987
rect 1559 1981 1563 1982
rect 1583 1986 1587 1987
rect 1583 1981 1587 1982
rect 1703 1986 1707 1987
rect 1703 1981 1707 1982
rect 1775 1986 1779 1987
rect 1775 1981 1779 1982
rect 2007 1986 2011 1987
rect 2007 1981 2011 1982
rect 2047 1986 2051 1987
rect 2047 1981 2051 1982
rect 2495 1986 2499 1987
rect 2495 1981 2499 1982
rect 2503 1986 2507 1987
rect 2503 1981 2507 1982
rect 2591 1986 2595 1987
rect 2591 1981 2595 1982
rect 2671 1986 2675 1987
rect 2671 1981 2675 1982
rect 2695 1986 2699 1987
rect 2695 1981 2699 1982
rect 2807 1986 2811 1987
rect 2807 1981 2811 1982
rect 2839 1986 2843 1987
rect 2839 1981 2843 1982
rect 2927 1986 2931 1987
rect 2927 1981 2931 1982
rect 3007 1986 3011 1987
rect 3007 1981 3011 1982
rect 3047 1986 3051 1987
rect 3047 1981 3051 1982
rect 3167 1986 3171 1987
rect 3167 1981 3171 1982
rect 3175 1986 3179 1987
rect 3175 1981 3179 1982
rect 3295 1986 3299 1987
rect 3295 1981 3299 1982
rect 3311 1986 3315 1987
rect 3311 1981 3315 1982
rect 3415 1986 3419 1987
rect 3415 1981 3419 1982
rect 3455 1986 3459 1987
rect 3455 1981 3459 1982
rect 3543 1986 3547 1987
rect 3543 1981 3547 1982
rect 3591 1986 3595 1987
rect 3591 1981 3595 1982
rect 3671 1986 3675 1987
rect 3671 1981 3675 1982
rect 3727 1986 3731 1987
rect 3727 1981 3731 1982
rect 3799 1986 3803 1987
rect 3799 1981 3803 1982
rect 3839 1986 3843 1987
rect 3839 1981 3843 1982
rect 3943 1986 3947 1987
rect 3943 1981 3947 1982
rect 112 1954 114 1981
rect 512 1957 514 1981
rect 624 1957 626 1981
rect 744 1957 746 1981
rect 872 1957 874 1981
rect 1008 1957 1010 1981
rect 1144 1957 1146 1981
rect 1280 1957 1282 1981
rect 1416 1957 1418 1981
rect 1560 1957 1562 1981
rect 1704 1957 1706 1981
rect 510 1956 516 1957
rect 110 1953 116 1954
rect 110 1949 111 1953
rect 115 1949 116 1953
rect 510 1952 511 1956
rect 515 1952 516 1956
rect 510 1951 516 1952
rect 622 1956 628 1957
rect 622 1952 623 1956
rect 627 1952 628 1956
rect 622 1951 628 1952
rect 742 1956 748 1957
rect 742 1952 743 1956
rect 747 1952 748 1956
rect 742 1951 748 1952
rect 870 1956 876 1957
rect 870 1952 871 1956
rect 875 1952 876 1956
rect 870 1951 876 1952
rect 1006 1956 1012 1957
rect 1006 1952 1007 1956
rect 1011 1952 1012 1956
rect 1006 1951 1012 1952
rect 1142 1956 1148 1957
rect 1142 1952 1143 1956
rect 1147 1952 1148 1956
rect 1142 1951 1148 1952
rect 1278 1956 1284 1957
rect 1278 1952 1279 1956
rect 1283 1952 1284 1956
rect 1278 1951 1284 1952
rect 1414 1956 1420 1957
rect 1414 1952 1415 1956
rect 1419 1952 1420 1956
rect 1414 1951 1420 1952
rect 1558 1956 1564 1957
rect 1558 1952 1559 1956
rect 1563 1952 1564 1956
rect 1558 1951 1564 1952
rect 1702 1956 1708 1957
rect 1702 1952 1703 1956
rect 1707 1952 1708 1956
rect 2008 1954 2010 1981
rect 2048 1954 2050 1981
rect 2496 1957 2498 1981
rect 2592 1957 2594 1981
rect 2696 1957 2698 1981
rect 2808 1957 2810 1981
rect 2928 1957 2930 1981
rect 3048 1957 3050 1981
rect 3176 1957 3178 1981
rect 3296 1957 3298 1981
rect 3416 1957 3418 1981
rect 3544 1957 3546 1981
rect 3672 1957 3674 1981
rect 3800 1957 3802 1981
rect 2494 1956 2500 1957
rect 1702 1951 1708 1952
rect 2006 1953 2012 1954
rect 110 1948 116 1949
rect 2006 1949 2007 1953
rect 2011 1949 2012 1953
rect 2006 1948 2012 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2494 1952 2495 1956
rect 2499 1952 2500 1956
rect 2494 1951 2500 1952
rect 2590 1956 2596 1957
rect 2590 1952 2591 1956
rect 2595 1952 2596 1956
rect 2590 1951 2596 1952
rect 2694 1956 2700 1957
rect 2694 1952 2695 1956
rect 2699 1952 2700 1956
rect 2694 1951 2700 1952
rect 2806 1956 2812 1957
rect 2806 1952 2807 1956
rect 2811 1952 2812 1956
rect 2806 1951 2812 1952
rect 2926 1956 2932 1957
rect 2926 1952 2927 1956
rect 2931 1952 2932 1956
rect 2926 1951 2932 1952
rect 3046 1956 3052 1957
rect 3046 1952 3047 1956
rect 3051 1952 3052 1956
rect 3046 1951 3052 1952
rect 3174 1956 3180 1957
rect 3174 1952 3175 1956
rect 3179 1952 3180 1956
rect 3174 1951 3180 1952
rect 3294 1956 3300 1957
rect 3294 1952 3295 1956
rect 3299 1952 3300 1956
rect 3294 1951 3300 1952
rect 3414 1956 3420 1957
rect 3414 1952 3415 1956
rect 3419 1952 3420 1956
rect 3414 1951 3420 1952
rect 3542 1956 3548 1957
rect 3542 1952 3543 1956
rect 3547 1952 3548 1956
rect 3542 1951 3548 1952
rect 3670 1956 3676 1957
rect 3670 1952 3671 1956
rect 3675 1952 3676 1956
rect 3670 1951 3676 1952
rect 3798 1956 3804 1957
rect 3798 1952 3799 1956
rect 3803 1952 3804 1956
rect 3944 1954 3946 1981
rect 3798 1951 3804 1952
rect 3942 1953 3948 1954
rect 2046 1948 2052 1949
rect 3942 1949 3943 1953
rect 3947 1949 3948 1953
rect 3942 1948 3948 1949
rect 510 1937 516 1938
rect 110 1936 116 1937
rect 110 1932 111 1936
rect 115 1932 116 1936
rect 510 1933 511 1937
rect 515 1933 516 1937
rect 510 1932 516 1933
rect 622 1937 628 1938
rect 622 1933 623 1937
rect 627 1933 628 1937
rect 622 1932 628 1933
rect 742 1937 748 1938
rect 742 1933 743 1937
rect 747 1933 748 1937
rect 742 1932 748 1933
rect 870 1937 876 1938
rect 870 1933 871 1937
rect 875 1933 876 1937
rect 870 1932 876 1933
rect 1006 1937 1012 1938
rect 1006 1933 1007 1937
rect 1011 1933 1012 1937
rect 1006 1932 1012 1933
rect 1142 1937 1148 1938
rect 1142 1933 1143 1937
rect 1147 1933 1148 1937
rect 1142 1932 1148 1933
rect 1278 1937 1284 1938
rect 1278 1933 1279 1937
rect 1283 1933 1284 1937
rect 1278 1932 1284 1933
rect 1414 1937 1420 1938
rect 1414 1933 1415 1937
rect 1419 1933 1420 1937
rect 1414 1932 1420 1933
rect 1558 1937 1564 1938
rect 1558 1933 1559 1937
rect 1563 1933 1564 1937
rect 1558 1932 1564 1933
rect 1702 1937 1708 1938
rect 2494 1937 2500 1938
rect 1702 1933 1703 1937
rect 1707 1933 1708 1937
rect 1702 1932 1708 1933
rect 2006 1936 2012 1937
rect 2006 1932 2007 1936
rect 2011 1932 2012 1936
rect 110 1931 116 1932
rect 112 1903 114 1931
rect 512 1903 514 1932
rect 624 1903 626 1932
rect 744 1903 746 1932
rect 872 1903 874 1932
rect 1008 1903 1010 1932
rect 1144 1903 1146 1932
rect 1280 1903 1282 1932
rect 1416 1903 1418 1932
rect 1560 1903 1562 1932
rect 1704 1903 1706 1932
rect 2006 1931 2012 1932
rect 2046 1936 2052 1937
rect 2046 1932 2047 1936
rect 2051 1932 2052 1936
rect 2494 1933 2495 1937
rect 2499 1933 2500 1937
rect 2494 1932 2500 1933
rect 2590 1937 2596 1938
rect 2590 1933 2591 1937
rect 2595 1933 2596 1937
rect 2590 1932 2596 1933
rect 2694 1937 2700 1938
rect 2694 1933 2695 1937
rect 2699 1933 2700 1937
rect 2694 1932 2700 1933
rect 2806 1937 2812 1938
rect 2806 1933 2807 1937
rect 2811 1933 2812 1937
rect 2806 1932 2812 1933
rect 2926 1937 2932 1938
rect 2926 1933 2927 1937
rect 2931 1933 2932 1937
rect 2926 1932 2932 1933
rect 3046 1937 3052 1938
rect 3046 1933 3047 1937
rect 3051 1933 3052 1937
rect 3046 1932 3052 1933
rect 3174 1937 3180 1938
rect 3174 1933 3175 1937
rect 3179 1933 3180 1937
rect 3174 1932 3180 1933
rect 3294 1937 3300 1938
rect 3294 1933 3295 1937
rect 3299 1933 3300 1937
rect 3294 1932 3300 1933
rect 3414 1937 3420 1938
rect 3414 1933 3415 1937
rect 3419 1933 3420 1937
rect 3414 1932 3420 1933
rect 3542 1937 3548 1938
rect 3542 1933 3543 1937
rect 3547 1933 3548 1937
rect 3542 1932 3548 1933
rect 3670 1937 3676 1938
rect 3670 1933 3671 1937
rect 3675 1933 3676 1937
rect 3670 1932 3676 1933
rect 3798 1937 3804 1938
rect 3798 1933 3799 1937
rect 3803 1933 3804 1937
rect 3798 1932 3804 1933
rect 3942 1936 3948 1937
rect 3942 1932 3943 1936
rect 3947 1932 3948 1936
rect 2046 1931 2052 1932
rect 2008 1903 2010 1931
rect 2048 1907 2050 1931
rect 2496 1907 2498 1932
rect 2592 1907 2594 1932
rect 2696 1907 2698 1932
rect 2808 1907 2810 1932
rect 2928 1907 2930 1932
rect 3048 1907 3050 1932
rect 3176 1907 3178 1932
rect 3296 1907 3298 1932
rect 3416 1907 3418 1932
rect 3544 1907 3546 1932
rect 3672 1907 3674 1932
rect 3800 1907 3802 1932
rect 3942 1931 3948 1932
rect 3944 1907 3946 1931
rect 2047 1906 2051 1907
rect 111 1902 115 1903
rect 111 1897 115 1898
rect 511 1902 515 1903
rect 511 1897 515 1898
rect 551 1902 555 1903
rect 551 1897 555 1898
rect 623 1902 627 1903
rect 623 1897 627 1898
rect 663 1902 667 1903
rect 663 1897 667 1898
rect 743 1902 747 1903
rect 743 1897 747 1898
rect 783 1902 787 1903
rect 783 1897 787 1898
rect 871 1902 875 1903
rect 871 1897 875 1898
rect 911 1902 915 1903
rect 911 1897 915 1898
rect 1007 1902 1011 1903
rect 1007 1897 1011 1898
rect 1047 1902 1051 1903
rect 1047 1897 1051 1898
rect 1143 1902 1147 1903
rect 1143 1897 1147 1898
rect 1175 1902 1179 1903
rect 1175 1897 1179 1898
rect 1279 1902 1283 1903
rect 1279 1897 1283 1898
rect 1311 1902 1315 1903
rect 1311 1897 1315 1898
rect 1415 1902 1419 1903
rect 1415 1897 1419 1898
rect 1447 1902 1451 1903
rect 1447 1897 1451 1898
rect 1559 1902 1563 1903
rect 1559 1897 1563 1898
rect 1583 1902 1587 1903
rect 1583 1897 1587 1898
rect 1703 1902 1707 1903
rect 1703 1897 1707 1898
rect 1719 1902 1723 1903
rect 1719 1897 1723 1898
rect 2007 1902 2011 1903
rect 2047 1901 2051 1902
rect 2071 1906 2075 1907
rect 2071 1901 2075 1902
rect 2247 1906 2251 1907
rect 2247 1901 2251 1902
rect 2439 1906 2443 1907
rect 2439 1901 2443 1902
rect 2495 1906 2499 1907
rect 2495 1901 2499 1902
rect 2591 1906 2595 1907
rect 2591 1901 2595 1902
rect 2623 1906 2627 1907
rect 2623 1901 2627 1902
rect 2695 1906 2699 1907
rect 2695 1901 2699 1902
rect 2791 1906 2795 1907
rect 2791 1901 2795 1902
rect 2807 1906 2811 1907
rect 2807 1901 2811 1902
rect 2927 1906 2931 1907
rect 2927 1901 2931 1902
rect 2959 1906 2963 1907
rect 2959 1901 2963 1902
rect 3047 1906 3051 1907
rect 3047 1901 3051 1902
rect 3127 1906 3131 1907
rect 3127 1901 3131 1902
rect 3175 1906 3179 1907
rect 3175 1901 3179 1902
rect 3295 1906 3299 1907
rect 3295 1901 3299 1902
rect 3303 1906 3307 1907
rect 3303 1901 3307 1902
rect 3415 1906 3419 1907
rect 3415 1901 3419 1902
rect 3487 1906 3491 1907
rect 3487 1901 3491 1902
rect 3543 1906 3547 1907
rect 3543 1901 3547 1902
rect 3671 1906 3675 1907
rect 3671 1901 3675 1902
rect 3799 1906 3803 1907
rect 3799 1901 3803 1902
rect 3839 1906 3843 1907
rect 3839 1901 3843 1902
rect 3943 1906 3947 1907
rect 3943 1901 3947 1902
rect 2007 1897 2011 1898
rect 112 1877 114 1897
rect 110 1876 116 1877
rect 552 1876 554 1897
rect 664 1876 666 1897
rect 784 1876 786 1897
rect 912 1876 914 1897
rect 1048 1876 1050 1897
rect 1176 1876 1178 1897
rect 1312 1876 1314 1897
rect 1448 1876 1450 1897
rect 1584 1876 1586 1897
rect 1720 1876 1722 1897
rect 2008 1877 2010 1897
rect 2048 1881 2050 1901
rect 2046 1880 2052 1881
rect 2072 1880 2074 1901
rect 2248 1880 2250 1901
rect 2440 1880 2442 1901
rect 2624 1880 2626 1901
rect 2792 1880 2794 1901
rect 2960 1880 2962 1901
rect 3128 1880 3130 1901
rect 3304 1880 3306 1901
rect 3488 1880 3490 1901
rect 3672 1880 3674 1901
rect 3840 1880 3842 1901
rect 3944 1881 3946 1901
rect 3942 1880 3948 1881
rect 2006 1876 2012 1877
rect 110 1872 111 1876
rect 115 1872 116 1876
rect 110 1871 116 1872
rect 550 1875 556 1876
rect 550 1871 551 1875
rect 555 1871 556 1875
rect 550 1870 556 1871
rect 662 1875 668 1876
rect 662 1871 663 1875
rect 667 1871 668 1875
rect 662 1870 668 1871
rect 782 1875 788 1876
rect 782 1871 783 1875
rect 787 1871 788 1875
rect 782 1870 788 1871
rect 910 1875 916 1876
rect 910 1871 911 1875
rect 915 1871 916 1875
rect 910 1870 916 1871
rect 1046 1875 1052 1876
rect 1046 1871 1047 1875
rect 1051 1871 1052 1875
rect 1046 1870 1052 1871
rect 1174 1875 1180 1876
rect 1174 1871 1175 1875
rect 1179 1871 1180 1875
rect 1174 1870 1180 1871
rect 1310 1875 1316 1876
rect 1310 1871 1311 1875
rect 1315 1871 1316 1875
rect 1310 1870 1316 1871
rect 1446 1875 1452 1876
rect 1446 1871 1447 1875
rect 1451 1871 1452 1875
rect 1446 1870 1452 1871
rect 1582 1875 1588 1876
rect 1582 1871 1583 1875
rect 1587 1871 1588 1875
rect 1582 1870 1588 1871
rect 1718 1875 1724 1876
rect 1718 1871 1719 1875
rect 1723 1871 1724 1875
rect 2006 1872 2007 1876
rect 2011 1872 2012 1876
rect 2046 1876 2047 1880
rect 2051 1876 2052 1880
rect 2046 1875 2052 1876
rect 2070 1879 2076 1880
rect 2070 1875 2071 1879
rect 2075 1875 2076 1879
rect 2070 1874 2076 1875
rect 2246 1879 2252 1880
rect 2246 1875 2247 1879
rect 2251 1875 2252 1879
rect 2246 1874 2252 1875
rect 2438 1879 2444 1880
rect 2438 1875 2439 1879
rect 2443 1875 2444 1879
rect 2438 1874 2444 1875
rect 2622 1879 2628 1880
rect 2622 1875 2623 1879
rect 2627 1875 2628 1879
rect 2622 1874 2628 1875
rect 2790 1879 2796 1880
rect 2790 1875 2791 1879
rect 2795 1875 2796 1879
rect 2790 1874 2796 1875
rect 2958 1879 2964 1880
rect 2958 1875 2959 1879
rect 2963 1875 2964 1879
rect 2958 1874 2964 1875
rect 3126 1879 3132 1880
rect 3126 1875 3127 1879
rect 3131 1875 3132 1879
rect 3126 1874 3132 1875
rect 3302 1879 3308 1880
rect 3302 1875 3303 1879
rect 3307 1875 3308 1879
rect 3302 1874 3308 1875
rect 3486 1879 3492 1880
rect 3486 1875 3487 1879
rect 3491 1875 3492 1879
rect 3486 1874 3492 1875
rect 3670 1879 3676 1880
rect 3670 1875 3671 1879
rect 3675 1875 3676 1879
rect 3670 1874 3676 1875
rect 3838 1879 3844 1880
rect 3838 1875 3839 1879
rect 3843 1875 3844 1879
rect 3942 1876 3943 1880
rect 3947 1876 3948 1880
rect 3942 1875 3948 1876
rect 3838 1874 3844 1875
rect 2006 1871 2012 1872
rect 1718 1870 1724 1871
rect 2046 1863 2052 1864
rect 110 1859 116 1860
rect 110 1855 111 1859
rect 115 1855 116 1859
rect 2006 1859 2012 1860
rect 110 1854 116 1855
rect 550 1856 556 1857
rect 112 1827 114 1854
rect 550 1852 551 1856
rect 555 1852 556 1856
rect 550 1851 556 1852
rect 662 1856 668 1857
rect 662 1852 663 1856
rect 667 1852 668 1856
rect 662 1851 668 1852
rect 782 1856 788 1857
rect 782 1852 783 1856
rect 787 1852 788 1856
rect 782 1851 788 1852
rect 910 1856 916 1857
rect 910 1852 911 1856
rect 915 1852 916 1856
rect 910 1851 916 1852
rect 1046 1856 1052 1857
rect 1046 1852 1047 1856
rect 1051 1852 1052 1856
rect 1046 1851 1052 1852
rect 1174 1856 1180 1857
rect 1174 1852 1175 1856
rect 1179 1852 1180 1856
rect 1174 1851 1180 1852
rect 1310 1856 1316 1857
rect 1310 1852 1311 1856
rect 1315 1852 1316 1856
rect 1310 1851 1316 1852
rect 1446 1856 1452 1857
rect 1446 1852 1447 1856
rect 1451 1852 1452 1856
rect 1446 1851 1452 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1718 1856 1724 1857
rect 1718 1852 1719 1856
rect 1723 1852 1724 1856
rect 2006 1855 2007 1859
rect 2011 1855 2012 1859
rect 2046 1859 2047 1863
rect 2051 1859 2052 1863
rect 3942 1863 3948 1864
rect 2046 1858 2052 1859
rect 2070 1860 2076 1861
rect 2006 1854 2012 1855
rect 1718 1851 1724 1852
rect 552 1827 554 1851
rect 664 1827 666 1851
rect 784 1827 786 1851
rect 912 1827 914 1851
rect 1048 1827 1050 1851
rect 1176 1827 1178 1851
rect 1312 1827 1314 1851
rect 1448 1827 1450 1851
rect 1584 1827 1586 1851
rect 1720 1827 1722 1851
rect 2008 1827 2010 1854
rect 2048 1831 2050 1858
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2070 1855 2076 1856
rect 2246 1860 2252 1861
rect 2246 1856 2247 1860
rect 2251 1856 2252 1860
rect 2246 1855 2252 1856
rect 2438 1860 2444 1861
rect 2438 1856 2439 1860
rect 2443 1856 2444 1860
rect 2438 1855 2444 1856
rect 2622 1860 2628 1861
rect 2622 1856 2623 1860
rect 2627 1856 2628 1860
rect 2622 1855 2628 1856
rect 2790 1860 2796 1861
rect 2790 1856 2791 1860
rect 2795 1856 2796 1860
rect 2790 1855 2796 1856
rect 2958 1860 2964 1861
rect 2958 1856 2959 1860
rect 2963 1856 2964 1860
rect 2958 1855 2964 1856
rect 3126 1860 3132 1861
rect 3126 1856 3127 1860
rect 3131 1856 3132 1860
rect 3126 1855 3132 1856
rect 3302 1860 3308 1861
rect 3302 1856 3303 1860
rect 3307 1856 3308 1860
rect 3302 1855 3308 1856
rect 3486 1860 3492 1861
rect 3486 1856 3487 1860
rect 3491 1856 3492 1860
rect 3486 1855 3492 1856
rect 3670 1860 3676 1861
rect 3670 1856 3671 1860
rect 3675 1856 3676 1860
rect 3670 1855 3676 1856
rect 3838 1860 3844 1861
rect 3838 1856 3839 1860
rect 3843 1856 3844 1860
rect 3942 1859 3943 1863
rect 3947 1859 3948 1863
rect 3942 1858 3948 1859
rect 3838 1855 3844 1856
rect 2072 1831 2074 1855
rect 2248 1831 2250 1855
rect 2440 1831 2442 1855
rect 2624 1831 2626 1855
rect 2792 1831 2794 1855
rect 2960 1831 2962 1855
rect 3128 1831 3130 1855
rect 3304 1831 3306 1855
rect 3488 1831 3490 1855
rect 3672 1831 3674 1855
rect 3840 1831 3842 1855
rect 3944 1831 3946 1858
rect 2047 1830 2051 1831
rect 111 1826 115 1827
rect 111 1821 115 1822
rect 503 1826 507 1827
rect 503 1821 507 1822
rect 551 1826 555 1827
rect 551 1821 555 1822
rect 615 1826 619 1827
rect 615 1821 619 1822
rect 663 1826 667 1827
rect 663 1821 667 1822
rect 735 1826 739 1827
rect 735 1821 739 1822
rect 783 1826 787 1827
rect 783 1821 787 1822
rect 863 1826 867 1827
rect 863 1821 867 1822
rect 911 1826 915 1827
rect 911 1821 915 1822
rect 999 1826 1003 1827
rect 999 1821 1003 1822
rect 1047 1826 1051 1827
rect 1047 1821 1051 1822
rect 1151 1826 1155 1827
rect 1151 1821 1155 1822
rect 1175 1826 1179 1827
rect 1175 1821 1179 1822
rect 1311 1826 1315 1827
rect 1311 1821 1315 1822
rect 1319 1826 1323 1827
rect 1319 1821 1323 1822
rect 1447 1826 1451 1827
rect 1447 1821 1451 1822
rect 1487 1826 1491 1827
rect 1487 1821 1491 1822
rect 1583 1826 1587 1827
rect 1583 1821 1587 1822
rect 1663 1826 1667 1827
rect 1663 1821 1667 1822
rect 1719 1826 1723 1827
rect 1719 1821 1723 1822
rect 1847 1826 1851 1827
rect 1847 1821 1851 1822
rect 2007 1826 2011 1827
rect 2047 1825 2051 1826
rect 2071 1830 2075 1831
rect 2071 1825 2075 1826
rect 2095 1830 2099 1831
rect 2095 1825 2099 1826
rect 2231 1830 2235 1831
rect 2231 1825 2235 1826
rect 2247 1830 2251 1831
rect 2247 1825 2251 1826
rect 2367 1830 2371 1831
rect 2367 1825 2371 1826
rect 2439 1830 2443 1831
rect 2439 1825 2443 1826
rect 2511 1830 2515 1831
rect 2511 1825 2515 1826
rect 2623 1830 2627 1831
rect 2623 1825 2627 1826
rect 2671 1830 2675 1831
rect 2671 1825 2675 1826
rect 2791 1830 2795 1831
rect 2791 1825 2795 1826
rect 2855 1830 2859 1831
rect 2855 1825 2859 1826
rect 2959 1830 2963 1831
rect 2959 1825 2963 1826
rect 3071 1830 3075 1831
rect 3071 1825 3075 1826
rect 3127 1830 3131 1831
rect 3127 1825 3131 1826
rect 3303 1830 3307 1831
rect 3303 1825 3307 1826
rect 3487 1830 3491 1831
rect 3487 1825 3491 1826
rect 3543 1830 3547 1831
rect 3543 1825 3547 1826
rect 3671 1830 3675 1831
rect 3671 1825 3675 1826
rect 3791 1830 3795 1831
rect 3791 1825 3795 1826
rect 3839 1830 3843 1831
rect 3839 1825 3843 1826
rect 3943 1830 3947 1831
rect 3943 1825 3947 1826
rect 2007 1821 2011 1822
rect 112 1794 114 1821
rect 504 1797 506 1821
rect 616 1797 618 1821
rect 736 1797 738 1821
rect 864 1797 866 1821
rect 1000 1797 1002 1821
rect 1152 1797 1154 1821
rect 1320 1797 1322 1821
rect 1488 1797 1490 1821
rect 1664 1797 1666 1821
rect 1848 1797 1850 1821
rect 502 1796 508 1797
rect 110 1793 116 1794
rect 110 1789 111 1793
rect 115 1789 116 1793
rect 502 1792 503 1796
rect 507 1792 508 1796
rect 502 1791 508 1792
rect 614 1796 620 1797
rect 614 1792 615 1796
rect 619 1792 620 1796
rect 614 1791 620 1792
rect 734 1796 740 1797
rect 734 1792 735 1796
rect 739 1792 740 1796
rect 734 1791 740 1792
rect 862 1796 868 1797
rect 862 1792 863 1796
rect 867 1792 868 1796
rect 862 1791 868 1792
rect 998 1796 1004 1797
rect 998 1792 999 1796
rect 1003 1792 1004 1796
rect 998 1791 1004 1792
rect 1150 1796 1156 1797
rect 1150 1792 1151 1796
rect 1155 1792 1156 1796
rect 1150 1791 1156 1792
rect 1318 1796 1324 1797
rect 1318 1792 1319 1796
rect 1323 1792 1324 1796
rect 1318 1791 1324 1792
rect 1486 1796 1492 1797
rect 1486 1792 1487 1796
rect 1491 1792 1492 1796
rect 1486 1791 1492 1792
rect 1662 1796 1668 1797
rect 1662 1792 1663 1796
rect 1667 1792 1668 1796
rect 1662 1791 1668 1792
rect 1846 1796 1852 1797
rect 1846 1792 1847 1796
rect 1851 1792 1852 1796
rect 2008 1794 2010 1821
rect 2048 1798 2050 1825
rect 2096 1801 2098 1825
rect 2232 1801 2234 1825
rect 2368 1801 2370 1825
rect 2512 1801 2514 1825
rect 2672 1801 2674 1825
rect 2856 1801 2858 1825
rect 3072 1801 3074 1825
rect 3304 1801 3306 1825
rect 3544 1801 3546 1825
rect 3792 1801 3794 1825
rect 2094 1800 2100 1801
rect 2046 1797 2052 1798
rect 1846 1791 1852 1792
rect 2006 1793 2012 1794
rect 110 1788 116 1789
rect 2006 1789 2007 1793
rect 2011 1789 2012 1793
rect 2046 1793 2047 1797
rect 2051 1793 2052 1797
rect 2094 1796 2095 1800
rect 2099 1796 2100 1800
rect 2094 1795 2100 1796
rect 2230 1800 2236 1801
rect 2230 1796 2231 1800
rect 2235 1796 2236 1800
rect 2230 1795 2236 1796
rect 2366 1800 2372 1801
rect 2366 1796 2367 1800
rect 2371 1796 2372 1800
rect 2366 1795 2372 1796
rect 2510 1800 2516 1801
rect 2510 1796 2511 1800
rect 2515 1796 2516 1800
rect 2510 1795 2516 1796
rect 2670 1800 2676 1801
rect 2670 1796 2671 1800
rect 2675 1796 2676 1800
rect 2670 1795 2676 1796
rect 2854 1800 2860 1801
rect 2854 1796 2855 1800
rect 2859 1796 2860 1800
rect 2854 1795 2860 1796
rect 3070 1800 3076 1801
rect 3070 1796 3071 1800
rect 3075 1796 3076 1800
rect 3070 1795 3076 1796
rect 3302 1800 3308 1801
rect 3302 1796 3303 1800
rect 3307 1796 3308 1800
rect 3302 1795 3308 1796
rect 3542 1800 3548 1801
rect 3542 1796 3543 1800
rect 3547 1796 3548 1800
rect 3542 1795 3548 1796
rect 3790 1800 3796 1801
rect 3790 1796 3791 1800
rect 3795 1796 3796 1800
rect 3944 1798 3946 1825
rect 3790 1795 3796 1796
rect 3942 1797 3948 1798
rect 2046 1792 2052 1793
rect 3942 1793 3943 1797
rect 3947 1793 3948 1797
rect 3942 1792 3948 1793
rect 2006 1788 2012 1789
rect 2094 1781 2100 1782
rect 2046 1780 2052 1781
rect 502 1777 508 1778
rect 110 1776 116 1777
rect 110 1772 111 1776
rect 115 1772 116 1776
rect 502 1773 503 1777
rect 507 1773 508 1777
rect 502 1772 508 1773
rect 614 1777 620 1778
rect 614 1773 615 1777
rect 619 1773 620 1777
rect 614 1772 620 1773
rect 734 1777 740 1778
rect 734 1773 735 1777
rect 739 1773 740 1777
rect 734 1772 740 1773
rect 862 1777 868 1778
rect 862 1773 863 1777
rect 867 1773 868 1777
rect 862 1772 868 1773
rect 998 1777 1004 1778
rect 998 1773 999 1777
rect 1003 1773 1004 1777
rect 998 1772 1004 1773
rect 1150 1777 1156 1778
rect 1150 1773 1151 1777
rect 1155 1773 1156 1777
rect 1150 1772 1156 1773
rect 1318 1777 1324 1778
rect 1318 1773 1319 1777
rect 1323 1773 1324 1777
rect 1318 1772 1324 1773
rect 1486 1777 1492 1778
rect 1486 1773 1487 1777
rect 1491 1773 1492 1777
rect 1486 1772 1492 1773
rect 1662 1777 1668 1778
rect 1662 1773 1663 1777
rect 1667 1773 1668 1777
rect 1662 1772 1668 1773
rect 1846 1777 1852 1778
rect 1846 1773 1847 1777
rect 1851 1773 1852 1777
rect 1846 1772 1852 1773
rect 2006 1776 2012 1777
rect 2006 1772 2007 1776
rect 2011 1772 2012 1776
rect 2046 1776 2047 1780
rect 2051 1776 2052 1780
rect 2094 1777 2095 1781
rect 2099 1777 2100 1781
rect 2094 1776 2100 1777
rect 2230 1781 2236 1782
rect 2230 1777 2231 1781
rect 2235 1777 2236 1781
rect 2230 1776 2236 1777
rect 2366 1781 2372 1782
rect 2366 1777 2367 1781
rect 2371 1777 2372 1781
rect 2366 1776 2372 1777
rect 2510 1781 2516 1782
rect 2510 1777 2511 1781
rect 2515 1777 2516 1781
rect 2510 1776 2516 1777
rect 2670 1781 2676 1782
rect 2670 1777 2671 1781
rect 2675 1777 2676 1781
rect 2670 1776 2676 1777
rect 2854 1781 2860 1782
rect 2854 1777 2855 1781
rect 2859 1777 2860 1781
rect 2854 1776 2860 1777
rect 3070 1781 3076 1782
rect 3070 1777 3071 1781
rect 3075 1777 3076 1781
rect 3070 1776 3076 1777
rect 3302 1781 3308 1782
rect 3302 1777 3303 1781
rect 3307 1777 3308 1781
rect 3302 1776 3308 1777
rect 3542 1781 3548 1782
rect 3542 1777 3543 1781
rect 3547 1777 3548 1781
rect 3542 1776 3548 1777
rect 3790 1781 3796 1782
rect 3790 1777 3791 1781
rect 3795 1777 3796 1781
rect 3790 1776 3796 1777
rect 3942 1780 3948 1781
rect 3942 1776 3943 1780
rect 3947 1776 3948 1780
rect 2046 1775 2052 1776
rect 110 1771 116 1772
rect 112 1751 114 1771
rect 504 1751 506 1772
rect 616 1751 618 1772
rect 736 1751 738 1772
rect 864 1751 866 1772
rect 1000 1751 1002 1772
rect 1152 1751 1154 1772
rect 1320 1751 1322 1772
rect 1488 1751 1490 1772
rect 1664 1751 1666 1772
rect 1848 1751 1850 1772
rect 2006 1771 2012 1772
rect 2008 1751 2010 1771
rect 2048 1755 2050 1775
rect 2096 1755 2098 1776
rect 2232 1755 2234 1776
rect 2368 1755 2370 1776
rect 2512 1755 2514 1776
rect 2672 1755 2674 1776
rect 2856 1755 2858 1776
rect 3072 1755 3074 1776
rect 3304 1755 3306 1776
rect 3544 1755 3546 1776
rect 3792 1755 3794 1776
rect 3942 1775 3948 1776
rect 3944 1755 3946 1775
rect 2047 1754 2051 1755
rect 111 1750 115 1751
rect 111 1745 115 1746
rect 343 1750 347 1751
rect 343 1745 347 1746
rect 463 1750 467 1751
rect 463 1745 467 1746
rect 503 1750 507 1751
rect 503 1745 507 1746
rect 591 1750 595 1751
rect 591 1745 595 1746
rect 615 1750 619 1751
rect 615 1745 619 1746
rect 719 1750 723 1751
rect 719 1745 723 1746
rect 735 1750 739 1751
rect 735 1745 739 1746
rect 847 1750 851 1751
rect 847 1745 851 1746
rect 863 1750 867 1751
rect 863 1745 867 1746
rect 983 1750 987 1751
rect 983 1745 987 1746
rect 999 1750 1003 1751
rect 999 1745 1003 1746
rect 1127 1750 1131 1751
rect 1127 1745 1131 1746
rect 1151 1750 1155 1751
rect 1151 1745 1155 1746
rect 1279 1750 1283 1751
rect 1279 1745 1283 1746
rect 1319 1750 1323 1751
rect 1319 1745 1323 1746
rect 1439 1750 1443 1751
rect 1439 1745 1443 1746
rect 1487 1750 1491 1751
rect 1487 1745 1491 1746
rect 1599 1750 1603 1751
rect 1599 1745 1603 1746
rect 1663 1750 1667 1751
rect 1663 1745 1667 1746
rect 1847 1750 1851 1751
rect 1847 1745 1851 1746
rect 2007 1750 2011 1751
rect 2047 1749 2051 1750
rect 2095 1754 2099 1755
rect 2095 1749 2099 1750
rect 2183 1754 2187 1755
rect 2183 1749 2187 1750
rect 2231 1754 2235 1755
rect 2231 1749 2235 1750
rect 2287 1754 2291 1755
rect 2287 1749 2291 1750
rect 2367 1754 2371 1755
rect 2367 1749 2371 1750
rect 2391 1754 2395 1755
rect 2391 1749 2395 1750
rect 2495 1754 2499 1755
rect 2495 1749 2499 1750
rect 2511 1754 2515 1755
rect 2511 1749 2515 1750
rect 2599 1754 2603 1755
rect 2599 1749 2603 1750
rect 2671 1754 2675 1755
rect 2671 1749 2675 1750
rect 2703 1754 2707 1755
rect 2703 1749 2707 1750
rect 2807 1754 2811 1755
rect 2807 1749 2811 1750
rect 2855 1754 2859 1755
rect 2855 1749 2859 1750
rect 2911 1754 2915 1755
rect 2911 1749 2915 1750
rect 3015 1754 3019 1755
rect 3015 1749 3019 1750
rect 3071 1754 3075 1755
rect 3071 1749 3075 1750
rect 3127 1754 3131 1755
rect 3127 1749 3131 1750
rect 3303 1754 3307 1755
rect 3303 1749 3307 1750
rect 3543 1754 3547 1755
rect 3543 1749 3547 1750
rect 3791 1754 3795 1755
rect 3791 1749 3795 1750
rect 3943 1754 3947 1755
rect 3943 1749 3947 1750
rect 2007 1745 2011 1746
rect 112 1725 114 1745
rect 110 1724 116 1725
rect 344 1724 346 1745
rect 464 1724 466 1745
rect 592 1724 594 1745
rect 720 1724 722 1745
rect 848 1724 850 1745
rect 984 1724 986 1745
rect 1128 1724 1130 1745
rect 1280 1724 1282 1745
rect 1440 1724 1442 1745
rect 1600 1724 1602 1745
rect 2008 1725 2010 1745
rect 2048 1729 2050 1749
rect 2046 1728 2052 1729
rect 2184 1728 2186 1749
rect 2288 1728 2290 1749
rect 2392 1728 2394 1749
rect 2496 1728 2498 1749
rect 2600 1728 2602 1749
rect 2704 1728 2706 1749
rect 2808 1728 2810 1749
rect 2912 1728 2914 1749
rect 3016 1728 3018 1749
rect 3128 1728 3130 1749
rect 3944 1729 3946 1749
rect 3942 1728 3948 1729
rect 2006 1724 2012 1725
rect 110 1720 111 1724
rect 115 1720 116 1724
rect 110 1719 116 1720
rect 342 1723 348 1724
rect 342 1719 343 1723
rect 347 1719 348 1723
rect 342 1718 348 1719
rect 462 1723 468 1724
rect 462 1719 463 1723
rect 467 1719 468 1723
rect 462 1718 468 1719
rect 590 1723 596 1724
rect 590 1719 591 1723
rect 595 1719 596 1723
rect 590 1718 596 1719
rect 718 1723 724 1724
rect 718 1719 719 1723
rect 723 1719 724 1723
rect 718 1718 724 1719
rect 846 1723 852 1724
rect 846 1719 847 1723
rect 851 1719 852 1723
rect 846 1718 852 1719
rect 982 1723 988 1724
rect 982 1719 983 1723
rect 987 1719 988 1723
rect 982 1718 988 1719
rect 1126 1723 1132 1724
rect 1126 1719 1127 1723
rect 1131 1719 1132 1723
rect 1126 1718 1132 1719
rect 1278 1723 1284 1724
rect 1278 1719 1279 1723
rect 1283 1719 1284 1723
rect 1278 1718 1284 1719
rect 1438 1723 1444 1724
rect 1438 1719 1439 1723
rect 1443 1719 1444 1723
rect 1438 1718 1444 1719
rect 1598 1723 1604 1724
rect 1598 1719 1599 1723
rect 1603 1719 1604 1723
rect 2006 1720 2007 1724
rect 2011 1720 2012 1724
rect 2046 1724 2047 1728
rect 2051 1724 2052 1728
rect 2046 1723 2052 1724
rect 2182 1727 2188 1728
rect 2182 1723 2183 1727
rect 2187 1723 2188 1727
rect 2182 1722 2188 1723
rect 2286 1727 2292 1728
rect 2286 1723 2287 1727
rect 2291 1723 2292 1727
rect 2286 1722 2292 1723
rect 2390 1727 2396 1728
rect 2390 1723 2391 1727
rect 2395 1723 2396 1727
rect 2390 1722 2396 1723
rect 2494 1727 2500 1728
rect 2494 1723 2495 1727
rect 2499 1723 2500 1727
rect 2494 1722 2500 1723
rect 2598 1727 2604 1728
rect 2598 1723 2599 1727
rect 2603 1723 2604 1727
rect 2598 1722 2604 1723
rect 2702 1727 2708 1728
rect 2702 1723 2703 1727
rect 2707 1723 2708 1727
rect 2702 1722 2708 1723
rect 2806 1727 2812 1728
rect 2806 1723 2807 1727
rect 2811 1723 2812 1727
rect 2806 1722 2812 1723
rect 2910 1727 2916 1728
rect 2910 1723 2911 1727
rect 2915 1723 2916 1727
rect 2910 1722 2916 1723
rect 3014 1727 3020 1728
rect 3014 1723 3015 1727
rect 3019 1723 3020 1727
rect 3014 1722 3020 1723
rect 3126 1727 3132 1728
rect 3126 1723 3127 1727
rect 3131 1723 3132 1727
rect 3942 1724 3943 1728
rect 3947 1724 3948 1728
rect 3942 1723 3948 1724
rect 3126 1722 3132 1723
rect 2006 1719 2012 1720
rect 1598 1718 1604 1719
rect 2046 1711 2052 1712
rect 110 1707 116 1708
rect 110 1703 111 1707
rect 115 1703 116 1707
rect 2006 1707 2012 1708
rect 110 1702 116 1703
rect 342 1704 348 1705
rect 112 1671 114 1702
rect 342 1700 343 1704
rect 347 1700 348 1704
rect 342 1699 348 1700
rect 462 1704 468 1705
rect 462 1700 463 1704
rect 467 1700 468 1704
rect 462 1699 468 1700
rect 590 1704 596 1705
rect 590 1700 591 1704
rect 595 1700 596 1704
rect 590 1699 596 1700
rect 718 1704 724 1705
rect 718 1700 719 1704
rect 723 1700 724 1704
rect 718 1699 724 1700
rect 846 1704 852 1705
rect 846 1700 847 1704
rect 851 1700 852 1704
rect 846 1699 852 1700
rect 982 1704 988 1705
rect 982 1700 983 1704
rect 987 1700 988 1704
rect 982 1699 988 1700
rect 1126 1704 1132 1705
rect 1126 1700 1127 1704
rect 1131 1700 1132 1704
rect 1126 1699 1132 1700
rect 1278 1704 1284 1705
rect 1278 1700 1279 1704
rect 1283 1700 1284 1704
rect 1278 1699 1284 1700
rect 1438 1704 1444 1705
rect 1438 1700 1439 1704
rect 1443 1700 1444 1704
rect 1438 1699 1444 1700
rect 1598 1704 1604 1705
rect 1598 1700 1599 1704
rect 1603 1700 1604 1704
rect 2006 1703 2007 1707
rect 2011 1703 2012 1707
rect 2046 1707 2047 1711
rect 2051 1707 2052 1711
rect 3942 1711 3948 1712
rect 2046 1706 2052 1707
rect 2182 1708 2188 1709
rect 2006 1702 2012 1703
rect 1598 1699 1604 1700
rect 344 1671 346 1699
rect 464 1671 466 1699
rect 592 1671 594 1699
rect 720 1671 722 1699
rect 848 1671 850 1699
rect 984 1671 986 1699
rect 1128 1671 1130 1699
rect 1280 1671 1282 1699
rect 1440 1671 1442 1699
rect 1600 1671 1602 1699
rect 2008 1671 2010 1702
rect 2048 1679 2050 1706
rect 2182 1704 2183 1708
rect 2187 1704 2188 1708
rect 2182 1703 2188 1704
rect 2286 1708 2292 1709
rect 2286 1704 2287 1708
rect 2291 1704 2292 1708
rect 2286 1703 2292 1704
rect 2390 1708 2396 1709
rect 2390 1704 2391 1708
rect 2395 1704 2396 1708
rect 2390 1703 2396 1704
rect 2494 1708 2500 1709
rect 2494 1704 2495 1708
rect 2499 1704 2500 1708
rect 2494 1703 2500 1704
rect 2598 1708 2604 1709
rect 2598 1704 2599 1708
rect 2603 1704 2604 1708
rect 2598 1703 2604 1704
rect 2702 1708 2708 1709
rect 2702 1704 2703 1708
rect 2707 1704 2708 1708
rect 2702 1703 2708 1704
rect 2806 1708 2812 1709
rect 2806 1704 2807 1708
rect 2811 1704 2812 1708
rect 2806 1703 2812 1704
rect 2910 1708 2916 1709
rect 2910 1704 2911 1708
rect 2915 1704 2916 1708
rect 2910 1703 2916 1704
rect 3014 1708 3020 1709
rect 3014 1704 3015 1708
rect 3019 1704 3020 1708
rect 3014 1703 3020 1704
rect 3126 1708 3132 1709
rect 3126 1704 3127 1708
rect 3131 1704 3132 1708
rect 3942 1707 3943 1711
rect 3947 1707 3948 1711
rect 3942 1706 3948 1707
rect 3126 1703 3132 1704
rect 2184 1679 2186 1703
rect 2288 1679 2290 1703
rect 2392 1679 2394 1703
rect 2496 1679 2498 1703
rect 2600 1679 2602 1703
rect 2704 1679 2706 1703
rect 2808 1679 2810 1703
rect 2912 1679 2914 1703
rect 3016 1679 3018 1703
rect 3128 1679 3130 1703
rect 3944 1679 3946 1706
rect 2047 1678 2051 1679
rect 2047 1673 2051 1674
rect 2183 1678 2187 1679
rect 2183 1673 2187 1674
rect 2231 1678 2235 1679
rect 2231 1673 2235 1674
rect 2287 1678 2291 1679
rect 2287 1673 2291 1674
rect 2367 1678 2371 1679
rect 2367 1673 2371 1674
rect 2391 1678 2395 1679
rect 2391 1673 2395 1674
rect 2495 1678 2499 1679
rect 2495 1673 2499 1674
rect 2519 1678 2523 1679
rect 2519 1673 2523 1674
rect 2599 1678 2603 1679
rect 2599 1673 2603 1674
rect 2679 1678 2683 1679
rect 2679 1673 2683 1674
rect 2703 1678 2707 1679
rect 2703 1673 2707 1674
rect 2807 1678 2811 1679
rect 2807 1673 2811 1674
rect 2847 1678 2851 1679
rect 2847 1673 2851 1674
rect 2911 1678 2915 1679
rect 2911 1673 2915 1674
rect 3015 1678 3019 1679
rect 3015 1673 3019 1674
rect 3023 1678 3027 1679
rect 3023 1673 3027 1674
rect 3127 1678 3131 1679
rect 3127 1673 3131 1674
rect 3191 1678 3195 1679
rect 3191 1673 3195 1674
rect 3359 1678 3363 1679
rect 3359 1673 3363 1674
rect 3527 1678 3531 1679
rect 3527 1673 3531 1674
rect 3695 1678 3699 1679
rect 3695 1673 3699 1674
rect 3839 1678 3843 1679
rect 3839 1673 3843 1674
rect 3943 1678 3947 1679
rect 3943 1673 3947 1674
rect 111 1670 115 1671
rect 111 1665 115 1666
rect 159 1670 163 1671
rect 159 1665 163 1666
rect 295 1670 299 1671
rect 295 1665 299 1666
rect 343 1670 347 1671
rect 343 1665 347 1666
rect 455 1670 459 1671
rect 455 1665 459 1666
rect 463 1670 467 1671
rect 463 1665 467 1666
rect 591 1670 595 1671
rect 591 1665 595 1666
rect 623 1670 627 1671
rect 623 1665 627 1666
rect 719 1670 723 1671
rect 719 1665 723 1666
rect 799 1670 803 1671
rect 799 1665 803 1666
rect 847 1670 851 1671
rect 847 1665 851 1666
rect 983 1670 987 1671
rect 983 1665 987 1666
rect 1127 1670 1131 1671
rect 1127 1665 1131 1666
rect 1167 1670 1171 1671
rect 1167 1665 1171 1666
rect 1279 1670 1283 1671
rect 1279 1665 1283 1666
rect 1351 1670 1355 1671
rect 1351 1665 1355 1666
rect 1439 1670 1443 1671
rect 1439 1665 1443 1666
rect 1543 1670 1547 1671
rect 1543 1665 1547 1666
rect 1599 1670 1603 1671
rect 1599 1665 1603 1666
rect 1735 1670 1739 1671
rect 1735 1665 1739 1666
rect 2007 1670 2011 1671
rect 2007 1665 2011 1666
rect 112 1638 114 1665
rect 160 1641 162 1665
rect 296 1641 298 1665
rect 456 1641 458 1665
rect 624 1641 626 1665
rect 800 1641 802 1665
rect 984 1641 986 1665
rect 1168 1641 1170 1665
rect 1352 1641 1354 1665
rect 1544 1641 1546 1665
rect 1736 1641 1738 1665
rect 158 1640 164 1641
rect 110 1637 116 1638
rect 110 1633 111 1637
rect 115 1633 116 1637
rect 158 1636 159 1640
rect 163 1636 164 1640
rect 158 1635 164 1636
rect 294 1640 300 1641
rect 294 1636 295 1640
rect 299 1636 300 1640
rect 294 1635 300 1636
rect 454 1640 460 1641
rect 454 1636 455 1640
rect 459 1636 460 1640
rect 454 1635 460 1636
rect 622 1640 628 1641
rect 622 1636 623 1640
rect 627 1636 628 1640
rect 622 1635 628 1636
rect 798 1640 804 1641
rect 798 1636 799 1640
rect 803 1636 804 1640
rect 798 1635 804 1636
rect 982 1640 988 1641
rect 982 1636 983 1640
rect 987 1636 988 1640
rect 982 1635 988 1636
rect 1166 1640 1172 1641
rect 1166 1636 1167 1640
rect 1171 1636 1172 1640
rect 1166 1635 1172 1636
rect 1350 1640 1356 1641
rect 1350 1636 1351 1640
rect 1355 1636 1356 1640
rect 1350 1635 1356 1636
rect 1542 1640 1548 1641
rect 1542 1636 1543 1640
rect 1547 1636 1548 1640
rect 1542 1635 1548 1636
rect 1734 1640 1740 1641
rect 1734 1636 1735 1640
rect 1739 1636 1740 1640
rect 2008 1638 2010 1665
rect 2048 1646 2050 1673
rect 2232 1649 2234 1673
rect 2368 1649 2370 1673
rect 2520 1649 2522 1673
rect 2680 1649 2682 1673
rect 2848 1649 2850 1673
rect 3024 1649 3026 1673
rect 3192 1649 3194 1673
rect 3360 1649 3362 1673
rect 3528 1649 3530 1673
rect 3696 1649 3698 1673
rect 3840 1649 3842 1673
rect 2230 1648 2236 1649
rect 2046 1645 2052 1646
rect 2046 1641 2047 1645
rect 2051 1641 2052 1645
rect 2230 1644 2231 1648
rect 2235 1644 2236 1648
rect 2230 1643 2236 1644
rect 2366 1648 2372 1649
rect 2366 1644 2367 1648
rect 2371 1644 2372 1648
rect 2366 1643 2372 1644
rect 2518 1648 2524 1649
rect 2518 1644 2519 1648
rect 2523 1644 2524 1648
rect 2518 1643 2524 1644
rect 2678 1648 2684 1649
rect 2678 1644 2679 1648
rect 2683 1644 2684 1648
rect 2678 1643 2684 1644
rect 2846 1648 2852 1649
rect 2846 1644 2847 1648
rect 2851 1644 2852 1648
rect 2846 1643 2852 1644
rect 3022 1648 3028 1649
rect 3022 1644 3023 1648
rect 3027 1644 3028 1648
rect 3022 1643 3028 1644
rect 3190 1648 3196 1649
rect 3190 1644 3191 1648
rect 3195 1644 3196 1648
rect 3190 1643 3196 1644
rect 3358 1648 3364 1649
rect 3358 1644 3359 1648
rect 3363 1644 3364 1648
rect 3358 1643 3364 1644
rect 3526 1648 3532 1649
rect 3526 1644 3527 1648
rect 3531 1644 3532 1648
rect 3526 1643 3532 1644
rect 3694 1648 3700 1649
rect 3694 1644 3695 1648
rect 3699 1644 3700 1648
rect 3694 1643 3700 1644
rect 3838 1648 3844 1649
rect 3838 1644 3839 1648
rect 3843 1644 3844 1648
rect 3944 1646 3946 1673
rect 3838 1643 3844 1644
rect 3942 1645 3948 1646
rect 2046 1640 2052 1641
rect 3942 1641 3943 1645
rect 3947 1641 3948 1645
rect 3942 1640 3948 1641
rect 1734 1635 1740 1636
rect 2006 1637 2012 1638
rect 110 1632 116 1633
rect 2006 1633 2007 1637
rect 2011 1633 2012 1637
rect 2006 1632 2012 1633
rect 2230 1629 2236 1630
rect 2046 1628 2052 1629
rect 2046 1624 2047 1628
rect 2051 1624 2052 1628
rect 2230 1625 2231 1629
rect 2235 1625 2236 1629
rect 2230 1624 2236 1625
rect 2366 1629 2372 1630
rect 2366 1625 2367 1629
rect 2371 1625 2372 1629
rect 2366 1624 2372 1625
rect 2518 1629 2524 1630
rect 2518 1625 2519 1629
rect 2523 1625 2524 1629
rect 2518 1624 2524 1625
rect 2678 1629 2684 1630
rect 2678 1625 2679 1629
rect 2683 1625 2684 1629
rect 2678 1624 2684 1625
rect 2846 1629 2852 1630
rect 2846 1625 2847 1629
rect 2851 1625 2852 1629
rect 2846 1624 2852 1625
rect 3022 1629 3028 1630
rect 3022 1625 3023 1629
rect 3027 1625 3028 1629
rect 3022 1624 3028 1625
rect 3190 1629 3196 1630
rect 3190 1625 3191 1629
rect 3195 1625 3196 1629
rect 3190 1624 3196 1625
rect 3358 1629 3364 1630
rect 3358 1625 3359 1629
rect 3363 1625 3364 1629
rect 3358 1624 3364 1625
rect 3526 1629 3532 1630
rect 3526 1625 3527 1629
rect 3531 1625 3532 1629
rect 3526 1624 3532 1625
rect 3694 1629 3700 1630
rect 3694 1625 3695 1629
rect 3699 1625 3700 1629
rect 3694 1624 3700 1625
rect 3838 1629 3844 1630
rect 3838 1625 3839 1629
rect 3843 1625 3844 1629
rect 3838 1624 3844 1625
rect 3942 1628 3948 1629
rect 3942 1624 3943 1628
rect 3947 1624 3948 1628
rect 2046 1623 2052 1624
rect 158 1621 164 1622
rect 110 1620 116 1621
rect 110 1616 111 1620
rect 115 1616 116 1620
rect 158 1617 159 1621
rect 163 1617 164 1621
rect 158 1616 164 1617
rect 294 1621 300 1622
rect 294 1617 295 1621
rect 299 1617 300 1621
rect 294 1616 300 1617
rect 454 1621 460 1622
rect 454 1617 455 1621
rect 459 1617 460 1621
rect 454 1616 460 1617
rect 622 1621 628 1622
rect 622 1617 623 1621
rect 627 1617 628 1621
rect 622 1616 628 1617
rect 798 1621 804 1622
rect 798 1617 799 1621
rect 803 1617 804 1621
rect 798 1616 804 1617
rect 982 1621 988 1622
rect 982 1617 983 1621
rect 987 1617 988 1621
rect 982 1616 988 1617
rect 1166 1621 1172 1622
rect 1166 1617 1167 1621
rect 1171 1617 1172 1621
rect 1166 1616 1172 1617
rect 1350 1621 1356 1622
rect 1350 1617 1351 1621
rect 1355 1617 1356 1621
rect 1350 1616 1356 1617
rect 1542 1621 1548 1622
rect 1542 1617 1543 1621
rect 1547 1617 1548 1621
rect 1542 1616 1548 1617
rect 1734 1621 1740 1622
rect 1734 1617 1735 1621
rect 1739 1617 1740 1621
rect 1734 1616 1740 1617
rect 2006 1620 2012 1621
rect 2006 1616 2007 1620
rect 2011 1616 2012 1620
rect 110 1615 116 1616
rect 112 1595 114 1615
rect 160 1595 162 1616
rect 296 1595 298 1616
rect 456 1595 458 1616
rect 624 1595 626 1616
rect 800 1595 802 1616
rect 984 1595 986 1616
rect 1168 1595 1170 1616
rect 1352 1595 1354 1616
rect 1544 1595 1546 1616
rect 1736 1595 1738 1616
rect 2006 1615 2012 1616
rect 2008 1595 2010 1615
rect 2048 1595 2050 1623
rect 2232 1595 2234 1624
rect 2368 1595 2370 1624
rect 2520 1595 2522 1624
rect 2680 1595 2682 1624
rect 2848 1595 2850 1624
rect 3024 1595 3026 1624
rect 3192 1595 3194 1624
rect 3360 1595 3362 1624
rect 3528 1595 3530 1624
rect 3696 1595 3698 1624
rect 3840 1595 3842 1624
rect 3942 1623 3948 1624
rect 3944 1595 3946 1623
rect 111 1594 115 1595
rect 111 1589 115 1590
rect 135 1594 139 1595
rect 135 1589 139 1590
rect 159 1594 163 1595
rect 159 1589 163 1590
rect 255 1594 259 1595
rect 255 1589 259 1590
rect 295 1594 299 1595
rect 295 1589 299 1590
rect 423 1594 427 1595
rect 423 1589 427 1590
rect 455 1594 459 1595
rect 455 1589 459 1590
rect 607 1594 611 1595
rect 607 1589 611 1590
rect 623 1594 627 1595
rect 623 1589 627 1590
rect 799 1594 803 1595
rect 799 1589 803 1590
rect 983 1594 987 1595
rect 983 1589 987 1590
rect 991 1594 995 1595
rect 991 1589 995 1590
rect 1167 1594 1171 1595
rect 1167 1589 1171 1590
rect 1183 1594 1187 1595
rect 1183 1589 1187 1590
rect 1351 1594 1355 1595
rect 1351 1589 1355 1590
rect 1367 1594 1371 1595
rect 1367 1589 1371 1590
rect 1543 1594 1547 1595
rect 1543 1589 1547 1590
rect 1551 1594 1555 1595
rect 1551 1589 1555 1590
rect 1735 1594 1739 1595
rect 1735 1589 1739 1590
rect 1903 1594 1907 1595
rect 1903 1589 1907 1590
rect 2007 1594 2011 1595
rect 2007 1589 2011 1590
rect 2047 1594 2051 1595
rect 2047 1589 2051 1590
rect 2071 1594 2075 1595
rect 2071 1589 2075 1590
rect 2231 1594 2235 1595
rect 2231 1589 2235 1590
rect 2271 1594 2275 1595
rect 2271 1589 2275 1590
rect 2367 1594 2371 1595
rect 2367 1589 2371 1590
rect 2495 1594 2499 1595
rect 2495 1589 2499 1590
rect 2519 1594 2523 1595
rect 2519 1589 2523 1590
rect 2679 1594 2683 1595
rect 2679 1589 2683 1590
rect 2711 1594 2715 1595
rect 2711 1589 2715 1590
rect 2847 1594 2851 1595
rect 2847 1589 2851 1590
rect 2911 1594 2915 1595
rect 2911 1589 2915 1590
rect 3023 1594 3027 1595
rect 3023 1589 3027 1590
rect 3095 1594 3099 1595
rect 3095 1589 3099 1590
rect 3191 1594 3195 1595
rect 3191 1589 3195 1590
rect 3263 1594 3267 1595
rect 3263 1589 3267 1590
rect 3359 1594 3363 1595
rect 3359 1589 3363 1590
rect 3423 1594 3427 1595
rect 3423 1589 3427 1590
rect 3527 1594 3531 1595
rect 3527 1589 3531 1590
rect 3567 1594 3571 1595
rect 3567 1589 3571 1590
rect 3695 1594 3699 1595
rect 3695 1589 3699 1590
rect 3711 1594 3715 1595
rect 3711 1589 3715 1590
rect 3839 1594 3843 1595
rect 3839 1589 3843 1590
rect 3943 1594 3947 1595
rect 3943 1589 3947 1590
rect 112 1569 114 1589
rect 110 1568 116 1569
rect 136 1568 138 1589
rect 256 1568 258 1589
rect 424 1568 426 1589
rect 608 1568 610 1589
rect 800 1568 802 1589
rect 992 1568 994 1589
rect 1184 1568 1186 1589
rect 1368 1568 1370 1589
rect 1552 1568 1554 1589
rect 1736 1568 1738 1589
rect 1904 1568 1906 1589
rect 2008 1569 2010 1589
rect 2048 1569 2050 1589
rect 2006 1568 2012 1569
rect 110 1564 111 1568
rect 115 1564 116 1568
rect 110 1563 116 1564
rect 134 1567 140 1568
rect 134 1563 135 1567
rect 139 1563 140 1567
rect 134 1562 140 1563
rect 254 1567 260 1568
rect 254 1563 255 1567
rect 259 1563 260 1567
rect 254 1562 260 1563
rect 422 1567 428 1568
rect 422 1563 423 1567
rect 427 1563 428 1567
rect 422 1562 428 1563
rect 606 1567 612 1568
rect 606 1563 607 1567
rect 611 1563 612 1567
rect 606 1562 612 1563
rect 798 1567 804 1568
rect 798 1563 799 1567
rect 803 1563 804 1567
rect 798 1562 804 1563
rect 990 1567 996 1568
rect 990 1563 991 1567
rect 995 1563 996 1567
rect 990 1562 996 1563
rect 1182 1567 1188 1568
rect 1182 1563 1183 1567
rect 1187 1563 1188 1567
rect 1182 1562 1188 1563
rect 1366 1567 1372 1568
rect 1366 1563 1367 1567
rect 1371 1563 1372 1567
rect 1366 1562 1372 1563
rect 1550 1567 1556 1568
rect 1550 1563 1551 1567
rect 1555 1563 1556 1567
rect 1550 1562 1556 1563
rect 1734 1567 1740 1568
rect 1734 1563 1735 1567
rect 1739 1563 1740 1567
rect 1734 1562 1740 1563
rect 1902 1567 1908 1568
rect 1902 1563 1903 1567
rect 1907 1563 1908 1567
rect 2006 1564 2007 1568
rect 2011 1564 2012 1568
rect 2006 1563 2012 1564
rect 2046 1568 2052 1569
rect 2072 1568 2074 1589
rect 2272 1568 2274 1589
rect 2496 1568 2498 1589
rect 2712 1568 2714 1589
rect 2912 1568 2914 1589
rect 3096 1568 3098 1589
rect 3264 1568 3266 1589
rect 3424 1568 3426 1589
rect 3568 1568 3570 1589
rect 3712 1568 3714 1589
rect 3840 1568 3842 1589
rect 3944 1569 3946 1589
rect 3942 1568 3948 1569
rect 2046 1564 2047 1568
rect 2051 1564 2052 1568
rect 2046 1563 2052 1564
rect 2070 1567 2076 1568
rect 2070 1563 2071 1567
rect 2075 1563 2076 1567
rect 1902 1562 1908 1563
rect 2070 1562 2076 1563
rect 2270 1567 2276 1568
rect 2270 1563 2271 1567
rect 2275 1563 2276 1567
rect 2270 1562 2276 1563
rect 2494 1567 2500 1568
rect 2494 1563 2495 1567
rect 2499 1563 2500 1567
rect 2494 1562 2500 1563
rect 2710 1567 2716 1568
rect 2710 1563 2711 1567
rect 2715 1563 2716 1567
rect 2710 1562 2716 1563
rect 2910 1567 2916 1568
rect 2910 1563 2911 1567
rect 2915 1563 2916 1567
rect 2910 1562 2916 1563
rect 3094 1567 3100 1568
rect 3094 1563 3095 1567
rect 3099 1563 3100 1567
rect 3094 1562 3100 1563
rect 3262 1567 3268 1568
rect 3262 1563 3263 1567
rect 3267 1563 3268 1567
rect 3262 1562 3268 1563
rect 3422 1567 3428 1568
rect 3422 1563 3423 1567
rect 3427 1563 3428 1567
rect 3422 1562 3428 1563
rect 3566 1567 3572 1568
rect 3566 1563 3567 1567
rect 3571 1563 3572 1567
rect 3566 1562 3572 1563
rect 3710 1567 3716 1568
rect 3710 1563 3711 1567
rect 3715 1563 3716 1567
rect 3710 1562 3716 1563
rect 3838 1567 3844 1568
rect 3838 1563 3839 1567
rect 3843 1563 3844 1567
rect 3942 1564 3943 1568
rect 3947 1564 3948 1568
rect 3942 1563 3948 1564
rect 3838 1562 3844 1563
rect 110 1551 116 1552
rect 110 1547 111 1551
rect 115 1547 116 1551
rect 2006 1551 2012 1552
rect 110 1546 116 1547
rect 134 1548 140 1549
rect 112 1515 114 1546
rect 134 1544 135 1548
rect 139 1544 140 1548
rect 134 1543 140 1544
rect 254 1548 260 1549
rect 254 1544 255 1548
rect 259 1544 260 1548
rect 254 1543 260 1544
rect 422 1548 428 1549
rect 422 1544 423 1548
rect 427 1544 428 1548
rect 422 1543 428 1544
rect 606 1548 612 1549
rect 606 1544 607 1548
rect 611 1544 612 1548
rect 606 1543 612 1544
rect 798 1548 804 1549
rect 798 1544 799 1548
rect 803 1544 804 1548
rect 798 1543 804 1544
rect 990 1548 996 1549
rect 990 1544 991 1548
rect 995 1544 996 1548
rect 990 1543 996 1544
rect 1182 1548 1188 1549
rect 1182 1544 1183 1548
rect 1187 1544 1188 1548
rect 1182 1543 1188 1544
rect 1366 1548 1372 1549
rect 1366 1544 1367 1548
rect 1371 1544 1372 1548
rect 1366 1543 1372 1544
rect 1550 1548 1556 1549
rect 1550 1544 1551 1548
rect 1555 1544 1556 1548
rect 1550 1543 1556 1544
rect 1734 1548 1740 1549
rect 1734 1544 1735 1548
rect 1739 1544 1740 1548
rect 1734 1543 1740 1544
rect 1902 1548 1908 1549
rect 1902 1544 1903 1548
rect 1907 1544 1908 1548
rect 2006 1547 2007 1551
rect 2011 1547 2012 1551
rect 2006 1546 2012 1547
rect 2046 1551 2052 1552
rect 2046 1547 2047 1551
rect 2051 1547 2052 1551
rect 3942 1551 3948 1552
rect 2046 1546 2052 1547
rect 2070 1548 2076 1549
rect 1902 1543 1908 1544
rect 136 1515 138 1543
rect 256 1515 258 1543
rect 424 1515 426 1543
rect 608 1515 610 1543
rect 800 1515 802 1543
rect 992 1515 994 1543
rect 1184 1515 1186 1543
rect 1368 1515 1370 1543
rect 1552 1515 1554 1543
rect 1736 1515 1738 1543
rect 1904 1515 1906 1543
rect 2008 1515 2010 1546
rect 2048 1519 2050 1546
rect 2070 1544 2071 1548
rect 2075 1544 2076 1548
rect 2070 1543 2076 1544
rect 2270 1548 2276 1549
rect 2270 1544 2271 1548
rect 2275 1544 2276 1548
rect 2270 1543 2276 1544
rect 2494 1548 2500 1549
rect 2494 1544 2495 1548
rect 2499 1544 2500 1548
rect 2494 1543 2500 1544
rect 2710 1548 2716 1549
rect 2710 1544 2711 1548
rect 2715 1544 2716 1548
rect 2710 1543 2716 1544
rect 2910 1548 2916 1549
rect 2910 1544 2911 1548
rect 2915 1544 2916 1548
rect 2910 1543 2916 1544
rect 3094 1548 3100 1549
rect 3094 1544 3095 1548
rect 3099 1544 3100 1548
rect 3094 1543 3100 1544
rect 3262 1548 3268 1549
rect 3262 1544 3263 1548
rect 3267 1544 3268 1548
rect 3262 1543 3268 1544
rect 3422 1548 3428 1549
rect 3422 1544 3423 1548
rect 3427 1544 3428 1548
rect 3422 1543 3428 1544
rect 3566 1548 3572 1549
rect 3566 1544 3567 1548
rect 3571 1544 3572 1548
rect 3566 1543 3572 1544
rect 3710 1548 3716 1549
rect 3710 1544 3711 1548
rect 3715 1544 3716 1548
rect 3710 1543 3716 1544
rect 3838 1548 3844 1549
rect 3838 1544 3839 1548
rect 3843 1544 3844 1548
rect 3942 1547 3943 1551
rect 3947 1547 3948 1551
rect 3942 1546 3948 1547
rect 3838 1543 3844 1544
rect 2072 1519 2074 1543
rect 2272 1519 2274 1543
rect 2496 1519 2498 1543
rect 2712 1519 2714 1543
rect 2912 1519 2914 1543
rect 3096 1519 3098 1543
rect 3264 1519 3266 1543
rect 3424 1519 3426 1543
rect 3568 1519 3570 1543
rect 3712 1519 3714 1543
rect 3840 1519 3842 1543
rect 3944 1519 3946 1546
rect 2047 1518 2051 1519
rect 111 1514 115 1515
rect 111 1509 115 1510
rect 135 1514 139 1515
rect 135 1509 139 1510
rect 247 1514 251 1515
rect 247 1509 251 1510
rect 255 1514 259 1515
rect 255 1509 259 1510
rect 399 1514 403 1515
rect 399 1509 403 1510
rect 423 1514 427 1515
rect 423 1509 427 1510
rect 559 1514 563 1515
rect 559 1509 563 1510
rect 607 1514 611 1515
rect 607 1509 611 1510
rect 719 1514 723 1515
rect 719 1509 723 1510
rect 799 1514 803 1515
rect 799 1509 803 1510
rect 879 1514 883 1515
rect 879 1509 883 1510
rect 991 1514 995 1515
rect 991 1509 995 1510
rect 1039 1514 1043 1515
rect 1039 1509 1043 1510
rect 1183 1514 1187 1515
rect 1183 1509 1187 1510
rect 1319 1514 1323 1515
rect 1319 1509 1323 1510
rect 1367 1514 1371 1515
rect 1367 1509 1371 1510
rect 1447 1514 1451 1515
rect 1447 1509 1451 1510
rect 1551 1514 1555 1515
rect 1551 1509 1555 1510
rect 1567 1514 1571 1515
rect 1567 1509 1571 1510
rect 1687 1514 1691 1515
rect 1687 1509 1691 1510
rect 1735 1514 1739 1515
rect 1735 1509 1739 1510
rect 1807 1514 1811 1515
rect 1807 1509 1811 1510
rect 1903 1514 1907 1515
rect 1903 1509 1907 1510
rect 2007 1514 2011 1515
rect 2047 1513 2051 1514
rect 2071 1518 2075 1519
rect 2071 1513 2075 1514
rect 2271 1518 2275 1519
rect 2271 1513 2275 1514
rect 2431 1518 2435 1519
rect 2431 1513 2435 1514
rect 2495 1518 2499 1519
rect 2495 1513 2499 1514
rect 2711 1518 2715 1519
rect 2711 1513 2715 1514
rect 2791 1518 2795 1519
rect 2791 1513 2795 1514
rect 2911 1518 2915 1519
rect 2911 1513 2915 1514
rect 3095 1518 3099 1519
rect 3095 1513 3099 1514
rect 3127 1518 3131 1519
rect 3127 1513 3131 1514
rect 3263 1518 3267 1519
rect 3263 1513 3267 1514
rect 3423 1518 3427 1519
rect 3423 1513 3427 1514
rect 3463 1518 3467 1519
rect 3463 1513 3467 1514
rect 3567 1518 3571 1519
rect 3567 1513 3571 1514
rect 3711 1518 3715 1519
rect 3711 1513 3715 1514
rect 3799 1518 3803 1519
rect 3799 1513 3803 1514
rect 3839 1518 3843 1519
rect 3839 1513 3843 1514
rect 3943 1518 3947 1519
rect 3943 1513 3947 1514
rect 2007 1509 2011 1510
rect 112 1482 114 1509
rect 136 1485 138 1509
rect 248 1485 250 1509
rect 400 1485 402 1509
rect 560 1485 562 1509
rect 720 1485 722 1509
rect 880 1485 882 1509
rect 1040 1485 1042 1509
rect 1184 1485 1186 1509
rect 1320 1485 1322 1509
rect 1448 1485 1450 1509
rect 1568 1485 1570 1509
rect 1688 1485 1690 1509
rect 1808 1485 1810 1509
rect 1904 1485 1906 1509
rect 134 1484 140 1485
rect 110 1481 116 1482
rect 110 1477 111 1481
rect 115 1477 116 1481
rect 134 1480 135 1484
rect 139 1480 140 1484
rect 134 1479 140 1480
rect 246 1484 252 1485
rect 246 1480 247 1484
rect 251 1480 252 1484
rect 246 1479 252 1480
rect 398 1484 404 1485
rect 398 1480 399 1484
rect 403 1480 404 1484
rect 398 1479 404 1480
rect 558 1484 564 1485
rect 558 1480 559 1484
rect 563 1480 564 1484
rect 558 1479 564 1480
rect 718 1484 724 1485
rect 718 1480 719 1484
rect 723 1480 724 1484
rect 718 1479 724 1480
rect 878 1484 884 1485
rect 878 1480 879 1484
rect 883 1480 884 1484
rect 878 1479 884 1480
rect 1038 1484 1044 1485
rect 1038 1480 1039 1484
rect 1043 1480 1044 1484
rect 1038 1479 1044 1480
rect 1182 1484 1188 1485
rect 1182 1480 1183 1484
rect 1187 1480 1188 1484
rect 1182 1479 1188 1480
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1446 1484 1452 1485
rect 1446 1480 1447 1484
rect 1451 1480 1452 1484
rect 1446 1479 1452 1480
rect 1566 1484 1572 1485
rect 1566 1480 1567 1484
rect 1571 1480 1572 1484
rect 1566 1479 1572 1480
rect 1686 1484 1692 1485
rect 1686 1480 1687 1484
rect 1691 1480 1692 1484
rect 1686 1479 1692 1480
rect 1806 1484 1812 1485
rect 1806 1480 1807 1484
rect 1811 1480 1812 1484
rect 1806 1479 1812 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 2008 1482 2010 1509
rect 2048 1486 2050 1513
rect 2072 1489 2074 1513
rect 2432 1489 2434 1513
rect 2792 1489 2794 1513
rect 3128 1489 3130 1513
rect 3464 1489 3466 1513
rect 3800 1489 3802 1513
rect 2070 1488 2076 1489
rect 2046 1485 2052 1486
rect 1902 1479 1908 1480
rect 2006 1481 2012 1482
rect 110 1476 116 1477
rect 2006 1477 2007 1481
rect 2011 1477 2012 1481
rect 2046 1481 2047 1485
rect 2051 1481 2052 1485
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 2430 1488 2436 1489
rect 2430 1484 2431 1488
rect 2435 1484 2436 1488
rect 2430 1483 2436 1484
rect 2790 1488 2796 1489
rect 2790 1484 2791 1488
rect 2795 1484 2796 1488
rect 2790 1483 2796 1484
rect 3126 1488 3132 1489
rect 3126 1484 3127 1488
rect 3131 1484 3132 1488
rect 3126 1483 3132 1484
rect 3462 1488 3468 1489
rect 3462 1484 3463 1488
rect 3467 1484 3468 1488
rect 3462 1483 3468 1484
rect 3798 1488 3804 1489
rect 3798 1484 3799 1488
rect 3803 1484 3804 1488
rect 3944 1486 3946 1513
rect 3798 1483 3804 1484
rect 3942 1485 3948 1486
rect 2046 1480 2052 1481
rect 3942 1481 3943 1485
rect 3947 1481 3948 1485
rect 3942 1480 3948 1481
rect 2006 1476 2012 1477
rect 2070 1469 2076 1470
rect 2046 1468 2052 1469
rect 134 1465 140 1466
rect 110 1464 116 1465
rect 110 1460 111 1464
rect 115 1460 116 1464
rect 134 1461 135 1465
rect 139 1461 140 1465
rect 134 1460 140 1461
rect 246 1465 252 1466
rect 246 1461 247 1465
rect 251 1461 252 1465
rect 246 1460 252 1461
rect 398 1465 404 1466
rect 398 1461 399 1465
rect 403 1461 404 1465
rect 398 1460 404 1461
rect 558 1465 564 1466
rect 558 1461 559 1465
rect 563 1461 564 1465
rect 558 1460 564 1461
rect 718 1465 724 1466
rect 718 1461 719 1465
rect 723 1461 724 1465
rect 718 1460 724 1461
rect 878 1465 884 1466
rect 878 1461 879 1465
rect 883 1461 884 1465
rect 878 1460 884 1461
rect 1038 1465 1044 1466
rect 1038 1461 1039 1465
rect 1043 1461 1044 1465
rect 1038 1460 1044 1461
rect 1182 1465 1188 1466
rect 1182 1461 1183 1465
rect 1187 1461 1188 1465
rect 1182 1460 1188 1461
rect 1318 1465 1324 1466
rect 1318 1461 1319 1465
rect 1323 1461 1324 1465
rect 1318 1460 1324 1461
rect 1446 1465 1452 1466
rect 1446 1461 1447 1465
rect 1451 1461 1452 1465
rect 1446 1460 1452 1461
rect 1566 1465 1572 1466
rect 1566 1461 1567 1465
rect 1571 1461 1572 1465
rect 1566 1460 1572 1461
rect 1686 1465 1692 1466
rect 1686 1461 1687 1465
rect 1691 1461 1692 1465
rect 1686 1460 1692 1461
rect 1806 1465 1812 1466
rect 1806 1461 1807 1465
rect 1811 1461 1812 1465
rect 1806 1460 1812 1461
rect 1902 1465 1908 1466
rect 1902 1461 1903 1465
rect 1907 1461 1908 1465
rect 1902 1460 1908 1461
rect 2006 1464 2012 1465
rect 2006 1460 2007 1464
rect 2011 1460 2012 1464
rect 2046 1464 2047 1468
rect 2051 1464 2052 1468
rect 2070 1465 2071 1469
rect 2075 1465 2076 1469
rect 2070 1464 2076 1465
rect 2430 1469 2436 1470
rect 2430 1465 2431 1469
rect 2435 1465 2436 1469
rect 2430 1464 2436 1465
rect 2790 1469 2796 1470
rect 2790 1465 2791 1469
rect 2795 1465 2796 1469
rect 2790 1464 2796 1465
rect 3126 1469 3132 1470
rect 3126 1465 3127 1469
rect 3131 1465 3132 1469
rect 3126 1464 3132 1465
rect 3462 1469 3468 1470
rect 3462 1465 3463 1469
rect 3467 1465 3468 1469
rect 3462 1464 3468 1465
rect 3798 1469 3804 1470
rect 3798 1465 3799 1469
rect 3803 1465 3804 1469
rect 3798 1464 3804 1465
rect 3942 1468 3948 1469
rect 3942 1464 3943 1468
rect 3947 1464 3948 1468
rect 2046 1463 2052 1464
rect 110 1459 116 1460
rect 112 1439 114 1459
rect 136 1439 138 1460
rect 248 1439 250 1460
rect 400 1439 402 1460
rect 560 1439 562 1460
rect 720 1439 722 1460
rect 880 1439 882 1460
rect 1040 1439 1042 1460
rect 1184 1439 1186 1460
rect 1320 1439 1322 1460
rect 1448 1439 1450 1460
rect 1568 1439 1570 1460
rect 1688 1439 1690 1460
rect 1808 1439 1810 1460
rect 1904 1439 1906 1460
rect 2006 1459 2012 1460
rect 2008 1439 2010 1459
rect 111 1438 115 1439
rect 111 1433 115 1434
rect 135 1438 139 1439
rect 135 1433 139 1434
rect 247 1438 251 1439
rect 247 1433 251 1434
rect 263 1438 267 1439
rect 263 1433 267 1434
rect 399 1438 403 1439
rect 399 1433 403 1434
rect 431 1438 435 1439
rect 431 1433 435 1434
rect 559 1438 563 1439
rect 559 1433 563 1434
rect 607 1438 611 1439
rect 607 1433 611 1434
rect 719 1438 723 1439
rect 719 1433 723 1434
rect 791 1438 795 1439
rect 791 1433 795 1434
rect 879 1438 883 1439
rect 879 1433 883 1434
rect 975 1438 979 1439
rect 975 1433 979 1434
rect 1039 1438 1043 1439
rect 1039 1433 1043 1434
rect 1159 1438 1163 1439
rect 1159 1433 1163 1434
rect 1183 1438 1187 1439
rect 1183 1433 1187 1434
rect 1319 1438 1323 1439
rect 1319 1433 1323 1434
rect 1351 1438 1355 1439
rect 1351 1433 1355 1434
rect 1447 1438 1451 1439
rect 1447 1433 1451 1434
rect 1543 1438 1547 1439
rect 1543 1433 1547 1434
rect 1567 1438 1571 1439
rect 1567 1433 1571 1434
rect 1687 1438 1691 1439
rect 1687 1433 1691 1434
rect 1735 1438 1739 1439
rect 1735 1433 1739 1434
rect 1807 1438 1811 1439
rect 1807 1433 1811 1434
rect 1903 1438 1907 1439
rect 1903 1433 1907 1434
rect 2007 1438 2011 1439
rect 2048 1435 2050 1463
rect 2072 1435 2074 1464
rect 2432 1435 2434 1464
rect 2792 1435 2794 1464
rect 3128 1435 3130 1464
rect 3464 1435 3466 1464
rect 3800 1435 3802 1464
rect 3942 1463 3948 1464
rect 3944 1435 3946 1463
rect 2007 1433 2011 1434
rect 2047 1434 2051 1435
rect 112 1413 114 1433
rect 110 1412 116 1413
rect 136 1412 138 1433
rect 264 1412 266 1433
rect 432 1412 434 1433
rect 608 1412 610 1433
rect 792 1412 794 1433
rect 976 1412 978 1433
rect 1160 1412 1162 1433
rect 1352 1412 1354 1433
rect 1544 1412 1546 1433
rect 1736 1412 1738 1433
rect 1904 1412 1906 1433
rect 2008 1413 2010 1433
rect 2047 1429 2051 1430
rect 2071 1434 2075 1435
rect 2071 1429 2075 1430
rect 2271 1434 2275 1435
rect 2271 1429 2275 1430
rect 2431 1434 2435 1435
rect 2431 1429 2435 1430
rect 2495 1434 2499 1435
rect 2495 1429 2499 1430
rect 2711 1434 2715 1435
rect 2711 1429 2715 1430
rect 2791 1434 2795 1435
rect 2791 1429 2795 1430
rect 2911 1434 2915 1435
rect 2911 1429 2915 1430
rect 3095 1434 3099 1435
rect 3095 1429 3099 1430
rect 3127 1434 3131 1435
rect 3127 1429 3131 1430
rect 3271 1434 3275 1435
rect 3271 1429 3275 1430
rect 3439 1434 3443 1435
rect 3439 1429 3443 1430
rect 3463 1434 3467 1435
rect 3463 1429 3467 1430
rect 3607 1434 3611 1435
rect 3607 1429 3611 1430
rect 3783 1434 3787 1435
rect 3783 1429 3787 1430
rect 3799 1434 3803 1435
rect 3799 1429 3803 1430
rect 3943 1434 3947 1435
rect 3943 1429 3947 1430
rect 2006 1412 2012 1413
rect 110 1408 111 1412
rect 115 1408 116 1412
rect 110 1407 116 1408
rect 134 1411 140 1412
rect 134 1407 135 1411
rect 139 1407 140 1411
rect 134 1406 140 1407
rect 262 1411 268 1412
rect 262 1407 263 1411
rect 267 1407 268 1411
rect 262 1406 268 1407
rect 430 1411 436 1412
rect 430 1407 431 1411
rect 435 1407 436 1411
rect 430 1406 436 1407
rect 606 1411 612 1412
rect 606 1407 607 1411
rect 611 1407 612 1411
rect 606 1406 612 1407
rect 790 1411 796 1412
rect 790 1407 791 1411
rect 795 1407 796 1411
rect 790 1406 796 1407
rect 974 1411 980 1412
rect 974 1407 975 1411
rect 979 1407 980 1411
rect 974 1406 980 1407
rect 1158 1411 1164 1412
rect 1158 1407 1159 1411
rect 1163 1407 1164 1411
rect 1158 1406 1164 1407
rect 1350 1411 1356 1412
rect 1350 1407 1351 1411
rect 1355 1407 1356 1411
rect 1350 1406 1356 1407
rect 1542 1411 1548 1412
rect 1542 1407 1543 1411
rect 1547 1407 1548 1411
rect 1542 1406 1548 1407
rect 1734 1411 1740 1412
rect 1734 1407 1735 1411
rect 1739 1407 1740 1411
rect 1734 1406 1740 1407
rect 1902 1411 1908 1412
rect 1902 1407 1903 1411
rect 1907 1407 1908 1411
rect 2006 1408 2007 1412
rect 2011 1408 2012 1412
rect 2048 1409 2050 1429
rect 2006 1407 2012 1408
rect 2046 1408 2052 1409
rect 2072 1408 2074 1429
rect 2272 1408 2274 1429
rect 2496 1408 2498 1429
rect 2712 1408 2714 1429
rect 2912 1408 2914 1429
rect 3096 1408 3098 1429
rect 3272 1408 3274 1429
rect 3440 1408 3442 1429
rect 3608 1408 3610 1429
rect 3784 1408 3786 1429
rect 3944 1409 3946 1429
rect 3942 1408 3948 1409
rect 1902 1406 1908 1407
rect 2046 1404 2047 1408
rect 2051 1404 2052 1408
rect 2046 1403 2052 1404
rect 2070 1407 2076 1408
rect 2070 1403 2071 1407
rect 2075 1403 2076 1407
rect 2070 1402 2076 1403
rect 2270 1407 2276 1408
rect 2270 1403 2271 1407
rect 2275 1403 2276 1407
rect 2270 1402 2276 1403
rect 2494 1407 2500 1408
rect 2494 1403 2495 1407
rect 2499 1403 2500 1407
rect 2494 1402 2500 1403
rect 2710 1407 2716 1408
rect 2710 1403 2711 1407
rect 2715 1403 2716 1407
rect 2710 1402 2716 1403
rect 2910 1407 2916 1408
rect 2910 1403 2911 1407
rect 2915 1403 2916 1407
rect 2910 1402 2916 1403
rect 3094 1407 3100 1408
rect 3094 1403 3095 1407
rect 3099 1403 3100 1407
rect 3094 1402 3100 1403
rect 3270 1407 3276 1408
rect 3270 1403 3271 1407
rect 3275 1403 3276 1407
rect 3270 1402 3276 1403
rect 3438 1407 3444 1408
rect 3438 1403 3439 1407
rect 3443 1403 3444 1407
rect 3438 1402 3444 1403
rect 3606 1407 3612 1408
rect 3606 1403 3607 1407
rect 3611 1403 3612 1407
rect 3606 1402 3612 1403
rect 3782 1407 3788 1408
rect 3782 1403 3783 1407
rect 3787 1403 3788 1407
rect 3942 1404 3943 1408
rect 3947 1404 3948 1408
rect 3942 1403 3948 1404
rect 3782 1402 3788 1403
rect 110 1395 116 1396
rect 110 1391 111 1395
rect 115 1391 116 1395
rect 2006 1395 2012 1396
rect 110 1390 116 1391
rect 134 1392 140 1393
rect 112 1359 114 1390
rect 134 1388 135 1392
rect 139 1388 140 1392
rect 134 1387 140 1388
rect 262 1392 268 1393
rect 262 1388 263 1392
rect 267 1388 268 1392
rect 262 1387 268 1388
rect 430 1392 436 1393
rect 430 1388 431 1392
rect 435 1388 436 1392
rect 430 1387 436 1388
rect 606 1392 612 1393
rect 606 1388 607 1392
rect 611 1388 612 1392
rect 606 1387 612 1388
rect 790 1392 796 1393
rect 790 1388 791 1392
rect 795 1388 796 1392
rect 790 1387 796 1388
rect 974 1392 980 1393
rect 974 1388 975 1392
rect 979 1388 980 1392
rect 974 1387 980 1388
rect 1158 1392 1164 1393
rect 1158 1388 1159 1392
rect 1163 1388 1164 1392
rect 1158 1387 1164 1388
rect 1350 1392 1356 1393
rect 1350 1388 1351 1392
rect 1355 1388 1356 1392
rect 1350 1387 1356 1388
rect 1542 1392 1548 1393
rect 1542 1388 1543 1392
rect 1547 1388 1548 1392
rect 1542 1387 1548 1388
rect 1734 1392 1740 1393
rect 1734 1388 1735 1392
rect 1739 1388 1740 1392
rect 1734 1387 1740 1388
rect 1902 1392 1908 1393
rect 1902 1388 1903 1392
rect 1907 1388 1908 1392
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2006 1390 2012 1391
rect 2046 1391 2052 1392
rect 1902 1387 1908 1388
rect 136 1359 138 1387
rect 264 1359 266 1387
rect 432 1359 434 1387
rect 608 1359 610 1387
rect 792 1359 794 1387
rect 976 1359 978 1387
rect 1160 1359 1162 1387
rect 1352 1359 1354 1387
rect 1544 1359 1546 1387
rect 1736 1359 1738 1387
rect 1904 1359 1906 1387
rect 2008 1359 2010 1390
rect 2046 1387 2047 1391
rect 2051 1387 2052 1391
rect 3942 1391 3948 1392
rect 2046 1386 2052 1387
rect 2070 1388 2076 1389
rect 2048 1359 2050 1386
rect 2070 1384 2071 1388
rect 2075 1384 2076 1388
rect 2070 1383 2076 1384
rect 2270 1388 2276 1389
rect 2270 1384 2271 1388
rect 2275 1384 2276 1388
rect 2270 1383 2276 1384
rect 2494 1388 2500 1389
rect 2494 1384 2495 1388
rect 2499 1384 2500 1388
rect 2494 1383 2500 1384
rect 2710 1388 2716 1389
rect 2710 1384 2711 1388
rect 2715 1384 2716 1388
rect 2710 1383 2716 1384
rect 2910 1388 2916 1389
rect 2910 1384 2911 1388
rect 2915 1384 2916 1388
rect 2910 1383 2916 1384
rect 3094 1388 3100 1389
rect 3094 1384 3095 1388
rect 3099 1384 3100 1388
rect 3094 1383 3100 1384
rect 3270 1388 3276 1389
rect 3270 1384 3271 1388
rect 3275 1384 3276 1388
rect 3270 1383 3276 1384
rect 3438 1388 3444 1389
rect 3438 1384 3439 1388
rect 3443 1384 3444 1388
rect 3438 1383 3444 1384
rect 3606 1388 3612 1389
rect 3606 1384 3607 1388
rect 3611 1384 3612 1388
rect 3606 1383 3612 1384
rect 3782 1388 3788 1389
rect 3782 1384 3783 1388
rect 3787 1384 3788 1388
rect 3942 1387 3943 1391
rect 3947 1387 3948 1391
rect 3942 1386 3948 1387
rect 3782 1383 3788 1384
rect 2072 1359 2074 1383
rect 2272 1359 2274 1383
rect 2496 1359 2498 1383
rect 2712 1359 2714 1383
rect 2912 1359 2914 1383
rect 3096 1359 3098 1383
rect 3272 1359 3274 1383
rect 3440 1359 3442 1383
rect 3608 1359 3610 1383
rect 3784 1359 3786 1383
rect 3944 1359 3946 1386
rect 111 1358 115 1359
rect 111 1353 115 1354
rect 135 1358 139 1359
rect 135 1353 139 1354
rect 159 1358 163 1359
rect 159 1353 163 1354
rect 263 1358 267 1359
rect 263 1353 267 1354
rect 311 1358 315 1359
rect 311 1353 315 1354
rect 431 1358 435 1359
rect 431 1353 435 1354
rect 479 1358 483 1359
rect 479 1353 483 1354
rect 607 1358 611 1359
rect 607 1353 611 1354
rect 663 1358 667 1359
rect 663 1353 667 1354
rect 791 1358 795 1359
rect 791 1353 795 1354
rect 855 1358 859 1359
rect 855 1353 859 1354
rect 975 1358 979 1359
rect 975 1353 979 1354
rect 1047 1358 1051 1359
rect 1047 1353 1051 1354
rect 1159 1358 1163 1359
rect 1159 1353 1163 1354
rect 1247 1358 1251 1359
rect 1247 1353 1251 1354
rect 1351 1358 1355 1359
rect 1351 1353 1355 1354
rect 1447 1358 1451 1359
rect 1447 1353 1451 1354
rect 1543 1358 1547 1359
rect 1543 1353 1547 1354
rect 1655 1358 1659 1359
rect 1655 1353 1659 1354
rect 1735 1358 1739 1359
rect 1735 1353 1739 1354
rect 1863 1358 1867 1359
rect 1863 1353 1867 1354
rect 1903 1358 1907 1359
rect 1903 1353 1907 1354
rect 2007 1358 2011 1359
rect 2007 1353 2011 1354
rect 2047 1358 2051 1359
rect 2047 1353 2051 1354
rect 2071 1358 2075 1359
rect 2071 1353 2075 1354
rect 2207 1358 2211 1359
rect 2207 1353 2211 1354
rect 2271 1358 2275 1359
rect 2271 1353 2275 1354
rect 2383 1358 2387 1359
rect 2383 1353 2387 1354
rect 2495 1358 2499 1359
rect 2495 1353 2499 1354
rect 2567 1358 2571 1359
rect 2567 1353 2571 1354
rect 2711 1358 2715 1359
rect 2711 1353 2715 1354
rect 2751 1358 2755 1359
rect 2751 1353 2755 1354
rect 2911 1358 2915 1359
rect 2911 1353 2915 1354
rect 2935 1358 2939 1359
rect 2935 1353 2939 1354
rect 3095 1358 3099 1359
rect 3095 1353 3099 1354
rect 3111 1358 3115 1359
rect 3111 1353 3115 1354
rect 3271 1358 3275 1359
rect 3271 1353 3275 1354
rect 3279 1358 3283 1359
rect 3279 1353 3283 1354
rect 3439 1358 3443 1359
rect 3439 1353 3443 1354
rect 3447 1358 3451 1359
rect 3447 1353 3451 1354
rect 3607 1358 3611 1359
rect 3607 1353 3611 1354
rect 3623 1358 3627 1359
rect 3623 1353 3627 1354
rect 3783 1358 3787 1359
rect 3783 1353 3787 1354
rect 3943 1358 3947 1359
rect 3943 1353 3947 1354
rect 112 1326 114 1353
rect 160 1329 162 1353
rect 312 1329 314 1353
rect 480 1329 482 1353
rect 664 1329 666 1353
rect 856 1329 858 1353
rect 1048 1329 1050 1353
rect 1248 1329 1250 1353
rect 1448 1329 1450 1353
rect 1656 1329 1658 1353
rect 1864 1329 1866 1353
rect 158 1328 164 1329
rect 110 1325 116 1326
rect 110 1321 111 1325
rect 115 1321 116 1325
rect 158 1324 159 1328
rect 163 1324 164 1328
rect 158 1323 164 1324
rect 310 1328 316 1329
rect 310 1324 311 1328
rect 315 1324 316 1328
rect 310 1323 316 1324
rect 478 1328 484 1329
rect 478 1324 479 1328
rect 483 1324 484 1328
rect 478 1323 484 1324
rect 662 1328 668 1329
rect 662 1324 663 1328
rect 667 1324 668 1328
rect 662 1323 668 1324
rect 854 1328 860 1329
rect 854 1324 855 1328
rect 859 1324 860 1328
rect 854 1323 860 1324
rect 1046 1328 1052 1329
rect 1046 1324 1047 1328
rect 1051 1324 1052 1328
rect 1046 1323 1052 1324
rect 1246 1328 1252 1329
rect 1246 1324 1247 1328
rect 1251 1324 1252 1328
rect 1246 1323 1252 1324
rect 1446 1328 1452 1329
rect 1446 1324 1447 1328
rect 1451 1324 1452 1328
rect 1446 1323 1452 1324
rect 1654 1328 1660 1329
rect 1654 1324 1655 1328
rect 1659 1324 1660 1328
rect 1654 1323 1660 1324
rect 1862 1328 1868 1329
rect 1862 1324 1863 1328
rect 1867 1324 1868 1328
rect 2008 1326 2010 1353
rect 2048 1326 2050 1353
rect 2072 1329 2074 1353
rect 2208 1329 2210 1353
rect 2384 1329 2386 1353
rect 2568 1329 2570 1353
rect 2752 1329 2754 1353
rect 2936 1329 2938 1353
rect 3112 1329 3114 1353
rect 3280 1329 3282 1353
rect 3448 1329 3450 1353
rect 3624 1329 3626 1353
rect 2070 1328 2076 1329
rect 1862 1323 1868 1324
rect 2006 1325 2012 1326
rect 110 1320 116 1321
rect 2006 1321 2007 1325
rect 2011 1321 2012 1325
rect 2006 1320 2012 1321
rect 2046 1325 2052 1326
rect 2046 1321 2047 1325
rect 2051 1321 2052 1325
rect 2070 1324 2071 1328
rect 2075 1324 2076 1328
rect 2070 1323 2076 1324
rect 2206 1328 2212 1329
rect 2206 1324 2207 1328
rect 2211 1324 2212 1328
rect 2206 1323 2212 1324
rect 2382 1328 2388 1329
rect 2382 1324 2383 1328
rect 2387 1324 2388 1328
rect 2382 1323 2388 1324
rect 2566 1328 2572 1329
rect 2566 1324 2567 1328
rect 2571 1324 2572 1328
rect 2566 1323 2572 1324
rect 2750 1328 2756 1329
rect 2750 1324 2751 1328
rect 2755 1324 2756 1328
rect 2750 1323 2756 1324
rect 2934 1328 2940 1329
rect 2934 1324 2935 1328
rect 2939 1324 2940 1328
rect 2934 1323 2940 1324
rect 3110 1328 3116 1329
rect 3110 1324 3111 1328
rect 3115 1324 3116 1328
rect 3110 1323 3116 1324
rect 3278 1328 3284 1329
rect 3278 1324 3279 1328
rect 3283 1324 3284 1328
rect 3278 1323 3284 1324
rect 3446 1328 3452 1329
rect 3446 1324 3447 1328
rect 3451 1324 3452 1328
rect 3446 1323 3452 1324
rect 3622 1328 3628 1329
rect 3622 1324 3623 1328
rect 3627 1324 3628 1328
rect 3944 1326 3946 1353
rect 3622 1323 3628 1324
rect 3942 1325 3948 1326
rect 2046 1320 2052 1321
rect 3942 1321 3943 1325
rect 3947 1321 3948 1325
rect 3942 1320 3948 1321
rect 158 1309 164 1310
rect 110 1308 116 1309
rect 110 1304 111 1308
rect 115 1304 116 1308
rect 158 1305 159 1309
rect 163 1305 164 1309
rect 158 1304 164 1305
rect 310 1309 316 1310
rect 310 1305 311 1309
rect 315 1305 316 1309
rect 310 1304 316 1305
rect 478 1309 484 1310
rect 478 1305 479 1309
rect 483 1305 484 1309
rect 478 1304 484 1305
rect 662 1309 668 1310
rect 662 1305 663 1309
rect 667 1305 668 1309
rect 662 1304 668 1305
rect 854 1309 860 1310
rect 854 1305 855 1309
rect 859 1305 860 1309
rect 854 1304 860 1305
rect 1046 1309 1052 1310
rect 1046 1305 1047 1309
rect 1051 1305 1052 1309
rect 1046 1304 1052 1305
rect 1246 1309 1252 1310
rect 1246 1305 1247 1309
rect 1251 1305 1252 1309
rect 1246 1304 1252 1305
rect 1446 1309 1452 1310
rect 1446 1305 1447 1309
rect 1451 1305 1452 1309
rect 1446 1304 1452 1305
rect 1654 1309 1660 1310
rect 1654 1305 1655 1309
rect 1659 1305 1660 1309
rect 1654 1304 1660 1305
rect 1862 1309 1868 1310
rect 2070 1309 2076 1310
rect 1862 1305 1863 1309
rect 1867 1305 1868 1309
rect 1862 1304 1868 1305
rect 2006 1308 2012 1309
rect 2006 1304 2007 1308
rect 2011 1304 2012 1308
rect 110 1303 116 1304
rect 112 1279 114 1303
rect 160 1279 162 1304
rect 312 1279 314 1304
rect 480 1279 482 1304
rect 664 1279 666 1304
rect 856 1279 858 1304
rect 1048 1279 1050 1304
rect 1248 1279 1250 1304
rect 1448 1279 1450 1304
rect 1656 1279 1658 1304
rect 1864 1279 1866 1304
rect 2006 1303 2012 1304
rect 2046 1308 2052 1309
rect 2046 1304 2047 1308
rect 2051 1304 2052 1308
rect 2070 1305 2071 1309
rect 2075 1305 2076 1309
rect 2070 1304 2076 1305
rect 2206 1309 2212 1310
rect 2206 1305 2207 1309
rect 2211 1305 2212 1309
rect 2206 1304 2212 1305
rect 2382 1309 2388 1310
rect 2382 1305 2383 1309
rect 2387 1305 2388 1309
rect 2382 1304 2388 1305
rect 2566 1309 2572 1310
rect 2566 1305 2567 1309
rect 2571 1305 2572 1309
rect 2566 1304 2572 1305
rect 2750 1309 2756 1310
rect 2750 1305 2751 1309
rect 2755 1305 2756 1309
rect 2750 1304 2756 1305
rect 2934 1309 2940 1310
rect 2934 1305 2935 1309
rect 2939 1305 2940 1309
rect 2934 1304 2940 1305
rect 3110 1309 3116 1310
rect 3110 1305 3111 1309
rect 3115 1305 3116 1309
rect 3110 1304 3116 1305
rect 3278 1309 3284 1310
rect 3278 1305 3279 1309
rect 3283 1305 3284 1309
rect 3278 1304 3284 1305
rect 3446 1309 3452 1310
rect 3446 1305 3447 1309
rect 3451 1305 3452 1309
rect 3446 1304 3452 1305
rect 3622 1309 3628 1310
rect 3622 1305 3623 1309
rect 3627 1305 3628 1309
rect 3622 1304 3628 1305
rect 3942 1308 3948 1309
rect 3942 1304 3943 1308
rect 3947 1304 3948 1308
rect 2046 1303 2052 1304
rect 2008 1279 2010 1303
rect 2048 1283 2050 1303
rect 2072 1283 2074 1304
rect 2208 1283 2210 1304
rect 2384 1283 2386 1304
rect 2568 1283 2570 1304
rect 2752 1283 2754 1304
rect 2936 1283 2938 1304
rect 3112 1283 3114 1304
rect 3280 1283 3282 1304
rect 3448 1283 3450 1304
rect 3624 1283 3626 1304
rect 3942 1303 3948 1304
rect 3944 1283 3946 1303
rect 2047 1282 2051 1283
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 159 1278 163 1279
rect 159 1273 163 1274
rect 311 1278 315 1279
rect 311 1273 315 1274
rect 407 1278 411 1279
rect 407 1273 411 1274
rect 479 1278 483 1279
rect 479 1273 483 1274
rect 543 1278 547 1279
rect 543 1273 547 1274
rect 663 1278 667 1279
rect 663 1273 667 1274
rect 695 1278 699 1279
rect 695 1273 699 1274
rect 855 1278 859 1279
rect 855 1273 859 1274
rect 1023 1278 1027 1279
rect 1023 1273 1027 1274
rect 1047 1278 1051 1279
rect 1047 1273 1051 1274
rect 1191 1278 1195 1279
rect 1191 1273 1195 1274
rect 1247 1278 1251 1279
rect 1247 1273 1251 1274
rect 1367 1278 1371 1279
rect 1367 1273 1371 1274
rect 1447 1278 1451 1279
rect 1447 1273 1451 1274
rect 1543 1278 1547 1279
rect 1543 1273 1547 1274
rect 1655 1278 1659 1279
rect 1655 1273 1659 1274
rect 1719 1278 1723 1279
rect 1719 1273 1723 1274
rect 1863 1278 1867 1279
rect 1863 1273 1867 1274
rect 1895 1278 1899 1279
rect 1895 1273 1899 1274
rect 2007 1278 2011 1279
rect 2047 1277 2051 1278
rect 2071 1282 2075 1283
rect 2071 1277 2075 1278
rect 2151 1282 2155 1283
rect 2151 1277 2155 1278
rect 2207 1282 2211 1283
rect 2207 1277 2211 1278
rect 2287 1282 2291 1283
rect 2287 1277 2291 1278
rect 2383 1282 2387 1283
rect 2383 1277 2387 1278
rect 2431 1282 2435 1283
rect 2431 1277 2435 1278
rect 2567 1282 2571 1283
rect 2567 1277 2571 1278
rect 2583 1282 2587 1283
rect 2583 1277 2587 1278
rect 2743 1282 2747 1283
rect 2743 1277 2747 1278
rect 2751 1282 2755 1283
rect 2751 1277 2755 1278
rect 2903 1282 2907 1283
rect 2903 1277 2907 1278
rect 2935 1282 2939 1283
rect 2935 1277 2939 1278
rect 3071 1282 3075 1283
rect 3071 1277 3075 1278
rect 3111 1282 3115 1283
rect 3111 1277 3115 1278
rect 3247 1282 3251 1283
rect 3247 1277 3251 1278
rect 3279 1282 3283 1283
rect 3279 1277 3283 1278
rect 3431 1282 3435 1283
rect 3431 1277 3435 1278
rect 3447 1282 3451 1283
rect 3447 1277 3451 1278
rect 3615 1282 3619 1283
rect 3615 1277 3619 1278
rect 3623 1282 3627 1283
rect 3623 1277 3627 1278
rect 3807 1282 3811 1283
rect 3807 1277 3811 1278
rect 3943 1282 3947 1283
rect 3943 1277 3947 1278
rect 2007 1273 2011 1274
rect 112 1253 114 1273
rect 110 1252 116 1253
rect 408 1252 410 1273
rect 544 1252 546 1273
rect 696 1252 698 1273
rect 856 1252 858 1273
rect 1024 1252 1026 1273
rect 1192 1252 1194 1273
rect 1368 1252 1370 1273
rect 1544 1252 1546 1273
rect 1720 1252 1722 1273
rect 1896 1252 1898 1273
rect 2008 1253 2010 1273
rect 2048 1257 2050 1277
rect 2046 1256 2052 1257
rect 2152 1256 2154 1277
rect 2288 1256 2290 1277
rect 2432 1256 2434 1277
rect 2584 1256 2586 1277
rect 2744 1256 2746 1277
rect 2904 1256 2906 1277
rect 3072 1256 3074 1277
rect 3248 1256 3250 1277
rect 3432 1256 3434 1277
rect 3616 1256 3618 1277
rect 3808 1256 3810 1277
rect 3944 1257 3946 1277
rect 3942 1256 3948 1257
rect 2006 1252 2012 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 110 1247 116 1248
rect 406 1251 412 1252
rect 406 1247 407 1251
rect 411 1247 412 1251
rect 406 1246 412 1247
rect 542 1251 548 1252
rect 542 1247 543 1251
rect 547 1247 548 1251
rect 542 1246 548 1247
rect 694 1251 700 1252
rect 694 1247 695 1251
rect 699 1247 700 1251
rect 694 1246 700 1247
rect 854 1251 860 1252
rect 854 1247 855 1251
rect 859 1247 860 1251
rect 854 1246 860 1247
rect 1022 1251 1028 1252
rect 1022 1247 1023 1251
rect 1027 1247 1028 1251
rect 1022 1246 1028 1247
rect 1190 1251 1196 1252
rect 1190 1247 1191 1251
rect 1195 1247 1196 1251
rect 1190 1246 1196 1247
rect 1366 1251 1372 1252
rect 1366 1247 1367 1251
rect 1371 1247 1372 1251
rect 1366 1246 1372 1247
rect 1542 1251 1548 1252
rect 1542 1247 1543 1251
rect 1547 1247 1548 1251
rect 1542 1246 1548 1247
rect 1718 1251 1724 1252
rect 1718 1247 1719 1251
rect 1723 1247 1724 1251
rect 1718 1246 1724 1247
rect 1894 1251 1900 1252
rect 1894 1247 1895 1251
rect 1899 1247 1900 1251
rect 2006 1248 2007 1252
rect 2011 1248 2012 1252
rect 2046 1252 2047 1256
rect 2051 1252 2052 1256
rect 2046 1251 2052 1252
rect 2150 1255 2156 1256
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2286 1255 2292 1256
rect 2286 1251 2287 1255
rect 2291 1251 2292 1255
rect 2286 1250 2292 1251
rect 2430 1255 2436 1256
rect 2430 1251 2431 1255
rect 2435 1251 2436 1255
rect 2430 1250 2436 1251
rect 2582 1255 2588 1256
rect 2582 1251 2583 1255
rect 2587 1251 2588 1255
rect 2582 1250 2588 1251
rect 2742 1255 2748 1256
rect 2742 1251 2743 1255
rect 2747 1251 2748 1255
rect 2742 1250 2748 1251
rect 2902 1255 2908 1256
rect 2902 1251 2903 1255
rect 2907 1251 2908 1255
rect 2902 1250 2908 1251
rect 3070 1255 3076 1256
rect 3070 1251 3071 1255
rect 3075 1251 3076 1255
rect 3070 1250 3076 1251
rect 3246 1255 3252 1256
rect 3246 1251 3247 1255
rect 3251 1251 3252 1255
rect 3246 1250 3252 1251
rect 3430 1255 3436 1256
rect 3430 1251 3431 1255
rect 3435 1251 3436 1255
rect 3430 1250 3436 1251
rect 3614 1255 3620 1256
rect 3614 1251 3615 1255
rect 3619 1251 3620 1255
rect 3614 1250 3620 1251
rect 3806 1255 3812 1256
rect 3806 1251 3807 1255
rect 3811 1251 3812 1255
rect 3942 1252 3943 1256
rect 3947 1252 3948 1256
rect 3942 1251 3948 1252
rect 3806 1250 3812 1251
rect 2006 1247 2012 1248
rect 1894 1246 1900 1247
rect 2046 1239 2052 1240
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 2006 1235 2012 1236
rect 110 1230 116 1231
rect 406 1232 412 1233
rect 112 1203 114 1230
rect 406 1228 407 1232
rect 411 1228 412 1232
rect 406 1227 412 1228
rect 542 1232 548 1233
rect 542 1228 543 1232
rect 547 1228 548 1232
rect 542 1227 548 1228
rect 694 1232 700 1233
rect 694 1228 695 1232
rect 699 1228 700 1232
rect 694 1227 700 1228
rect 854 1232 860 1233
rect 854 1228 855 1232
rect 859 1228 860 1232
rect 854 1227 860 1228
rect 1022 1232 1028 1233
rect 1022 1228 1023 1232
rect 1027 1228 1028 1232
rect 1022 1227 1028 1228
rect 1190 1232 1196 1233
rect 1190 1228 1191 1232
rect 1195 1228 1196 1232
rect 1190 1227 1196 1228
rect 1366 1232 1372 1233
rect 1366 1228 1367 1232
rect 1371 1228 1372 1232
rect 1366 1227 1372 1228
rect 1542 1232 1548 1233
rect 1542 1228 1543 1232
rect 1547 1228 1548 1232
rect 1542 1227 1548 1228
rect 1718 1232 1724 1233
rect 1718 1228 1719 1232
rect 1723 1228 1724 1232
rect 1718 1227 1724 1228
rect 1894 1232 1900 1233
rect 1894 1228 1895 1232
rect 1899 1228 1900 1232
rect 2006 1231 2007 1235
rect 2011 1231 2012 1235
rect 2046 1235 2047 1239
rect 2051 1235 2052 1239
rect 3942 1239 3948 1240
rect 2046 1234 2052 1235
rect 2150 1236 2156 1237
rect 2006 1230 2012 1231
rect 1894 1227 1900 1228
rect 408 1203 410 1227
rect 544 1203 546 1227
rect 696 1203 698 1227
rect 856 1203 858 1227
rect 1024 1203 1026 1227
rect 1192 1203 1194 1227
rect 1368 1203 1370 1227
rect 1544 1203 1546 1227
rect 1720 1203 1722 1227
rect 1896 1203 1898 1227
rect 2008 1203 2010 1230
rect 2048 1207 2050 1234
rect 2150 1232 2151 1236
rect 2155 1232 2156 1236
rect 2150 1231 2156 1232
rect 2286 1236 2292 1237
rect 2286 1232 2287 1236
rect 2291 1232 2292 1236
rect 2286 1231 2292 1232
rect 2430 1236 2436 1237
rect 2430 1232 2431 1236
rect 2435 1232 2436 1236
rect 2430 1231 2436 1232
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 2582 1231 2588 1232
rect 2742 1236 2748 1237
rect 2742 1232 2743 1236
rect 2747 1232 2748 1236
rect 2742 1231 2748 1232
rect 2902 1236 2908 1237
rect 2902 1232 2903 1236
rect 2907 1232 2908 1236
rect 2902 1231 2908 1232
rect 3070 1236 3076 1237
rect 3070 1232 3071 1236
rect 3075 1232 3076 1236
rect 3070 1231 3076 1232
rect 3246 1236 3252 1237
rect 3246 1232 3247 1236
rect 3251 1232 3252 1236
rect 3246 1231 3252 1232
rect 3430 1236 3436 1237
rect 3430 1232 3431 1236
rect 3435 1232 3436 1236
rect 3430 1231 3436 1232
rect 3614 1236 3620 1237
rect 3614 1232 3615 1236
rect 3619 1232 3620 1236
rect 3614 1231 3620 1232
rect 3806 1236 3812 1237
rect 3806 1232 3807 1236
rect 3811 1232 3812 1236
rect 3942 1235 3943 1239
rect 3947 1235 3948 1239
rect 3942 1234 3948 1235
rect 3806 1231 3812 1232
rect 2152 1207 2154 1231
rect 2288 1207 2290 1231
rect 2432 1207 2434 1231
rect 2584 1207 2586 1231
rect 2744 1207 2746 1231
rect 2904 1207 2906 1231
rect 3072 1207 3074 1231
rect 3248 1207 3250 1231
rect 3432 1207 3434 1231
rect 3616 1207 3618 1231
rect 3808 1207 3810 1231
rect 3944 1207 3946 1234
rect 2047 1206 2051 1207
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 407 1202 411 1203
rect 407 1197 411 1198
rect 423 1202 427 1203
rect 423 1197 427 1198
rect 543 1202 547 1203
rect 543 1197 547 1198
rect 591 1202 595 1203
rect 591 1197 595 1198
rect 695 1202 699 1203
rect 695 1197 699 1198
rect 759 1202 763 1203
rect 759 1197 763 1198
rect 855 1202 859 1203
rect 855 1197 859 1198
rect 927 1202 931 1203
rect 927 1197 931 1198
rect 1023 1202 1027 1203
rect 1023 1197 1027 1198
rect 1095 1202 1099 1203
rect 1095 1197 1099 1198
rect 1191 1202 1195 1203
rect 1191 1197 1195 1198
rect 1247 1202 1251 1203
rect 1247 1197 1251 1198
rect 1367 1202 1371 1203
rect 1367 1197 1371 1198
rect 1399 1202 1403 1203
rect 1399 1197 1403 1198
rect 1543 1202 1547 1203
rect 1543 1197 1547 1198
rect 1687 1202 1691 1203
rect 1687 1197 1691 1198
rect 1719 1202 1723 1203
rect 1719 1197 1723 1198
rect 1839 1202 1843 1203
rect 1839 1197 1843 1198
rect 1895 1202 1899 1203
rect 1895 1197 1899 1198
rect 2007 1202 2011 1203
rect 2047 1201 2051 1202
rect 2151 1206 2155 1207
rect 2151 1201 2155 1202
rect 2287 1206 2291 1207
rect 2287 1201 2291 1202
rect 2311 1206 2315 1207
rect 2311 1201 2315 1202
rect 2415 1206 2419 1207
rect 2415 1201 2419 1202
rect 2431 1206 2435 1207
rect 2431 1201 2435 1202
rect 2527 1206 2531 1207
rect 2527 1201 2531 1202
rect 2583 1206 2587 1207
rect 2583 1201 2587 1202
rect 2639 1206 2643 1207
rect 2639 1201 2643 1202
rect 2743 1206 2747 1207
rect 2743 1201 2747 1202
rect 2767 1206 2771 1207
rect 2767 1201 2771 1202
rect 2903 1206 2907 1207
rect 2903 1201 2907 1202
rect 2911 1206 2915 1207
rect 2911 1201 2915 1202
rect 3071 1206 3075 1207
rect 3071 1201 3075 1202
rect 3247 1206 3251 1207
rect 3247 1201 3251 1202
rect 3431 1206 3435 1207
rect 3431 1201 3435 1202
rect 3439 1206 3443 1207
rect 3439 1201 3443 1202
rect 3615 1206 3619 1207
rect 3615 1201 3619 1202
rect 3631 1206 3635 1207
rect 3631 1201 3635 1202
rect 3807 1206 3811 1207
rect 3807 1201 3811 1202
rect 3831 1206 3835 1207
rect 3831 1201 3835 1202
rect 3943 1206 3947 1207
rect 3943 1201 3947 1202
rect 2007 1197 2011 1198
rect 112 1170 114 1197
rect 424 1173 426 1197
rect 592 1173 594 1197
rect 760 1173 762 1197
rect 928 1173 930 1197
rect 1096 1173 1098 1197
rect 1248 1173 1250 1197
rect 1400 1173 1402 1197
rect 1544 1173 1546 1197
rect 1688 1173 1690 1197
rect 1840 1173 1842 1197
rect 422 1172 428 1173
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 422 1168 423 1172
rect 427 1168 428 1172
rect 422 1167 428 1168
rect 590 1172 596 1173
rect 590 1168 591 1172
rect 595 1168 596 1172
rect 590 1167 596 1168
rect 758 1172 764 1173
rect 758 1168 759 1172
rect 763 1168 764 1172
rect 758 1167 764 1168
rect 926 1172 932 1173
rect 926 1168 927 1172
rect 931 1168 932 1172
rect 926 1167 932 1168
rect 1094 1172 1100 1173
rect 1094 1168 1095 1172
rect 1099 1168 1100 1172
rect 1094 1167 1100 1168
rect 1246 1172 1252 1173
rect 1246 1168 1247 1172
rect 1251 1168 1252 1172
rect 1246 1167 1252 1168
rect 1398 1172 1404 1173
rect 1398 1168 1399 1172
rect 1403 1168 1404 1172
rect 1398 1167 1404 1168
rect 1542 1172 1548 1173
rect 1542 1168 1543 1172
rect 1547 1168 1548 1172
rect 1542 1167 1548 1168
rect 1686 1172 1692 1173
rect 1686 1168 1687 1172
rect 1691 1168 1692 1172
rect 1686 1167 1692 1168
rect 1838 1172 1844 1173
rect 1838 1168 1839 1172
rect 1843 1168 1844 1172
rect 2008 1170 2010 1197
rect 2048 1174 2050 1201
rect 2312 1177 2314 1201
rect 2416 1177 2418 1201
rect 2528 1177 2530 1201
rect 2640 1177 2642 1201
rect 2768 1177 2770 1201
rect 2912 1177 2914 1201
rect 3072 1177 3074 1201
rect 3248 1177 3250 1201
rect 3440 1177 3442 1201
rect 3632 1177 3634 1201
rect 3832 1177 3834 1201
rect 2310 1176 2316 1177
rect 2046 1173 2052 1174
rect 1838 1167 1844 1168
rect 2006 1169 2012 1170
rect 110 1164 116 1165
rect 2006 1165 2007 1169
rect 2011 1165 2012 1169
rect 2046 1169 2047 1173
rect 2051 1169 2052 1173
rect 2310 1172 2311 1176
rect 2315 1172 2316 1176
rect 2310 1171 2316 1172
rect 2414 1176 2420 1177
rect 2414 1172 2415 1176
rect 2419 1172 2420 1176
rect 2414 1171 2420 1172
rect 2526 1176 2532 1177
rect 2526 1172 2527 1176
rect 2531 1172 2532 1176
rect 2526 1171 2532 1172
rect 2638 1176 2644 1177
rect 2638 1172 2639 1176
rect 2643 1172 2644 1176
rect 2638 1171 2644 1172
rect 2766 1176 2772 1177
rect 2766 1172 2767 1176
rect 2771 1172 2772 1176
rect 2766 1171 2772 1172
rect 2910 1176 2916 1177
rect 2910 1172 2911 1176
rect 2915 1172 2916 1176
rect 2910 1171 2916 1172
rect 3070 1176 3076 1177
rect 3070 1172 3071 1176
rect 3075 1172 3076 1176
rect 3070 1171 3076 1172
rect 3246 1176 3252 1177
rect 3246 1172 3247 1176
rect 3251 1172 3252 1176
rect 3246 1171 3252 1172
rect 3438 1176 3444 1177
rect 3438 1172 3439 1176
rect 3443 1172 3444 1176
rect 3438 1171 3444 1172
rect 3630 1176 3636 1177
rect 3630 1172 3631 1176
rect 3635 1172 3636 1176
rect 3630 1171 3636 1172
rect 3830 1176 3836 1177
rect 3830 1172 3831 1176
rect 3835 1172 3836 1176
rect 3944 1174 3946 1201
rect 3830 1171 3836 1172
rect 3942 1173 3948 1174
rect 2046 1168 2052 1169
rect 3942 1169 3943 1173
rect 3947 1169 3948 1173
rect 3942 1168 3948 1169
rect 2006 1164 2012 1165
rect 2310 1157 2316 1158
rect 2046 1156 2052 1157
rect 422 1153 428 1154
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 422 1149 423 1153
rect 427 1149 428 1153
rect 422 1148 428 1149
rect 590 1153 596 1154
rect 590 1149 591 1153
rect 595 1149 596 1153
rect 590 1148 596 1149
rect 758 1153 764 1154
rect 758 1149 759 1153
rect 763 1149 764 1153
rect 758 1148 764 1149
rect 926 1153 932 1154
rect 926 1149 927 1153
rect 931 1149 932 1153
rect 926 1148 932 1149
rect 1094 1153 1100 1154
rect 1094 1149 1095 1153
rect 1099 1149 1100 1153
rect 1094 1148 1100 1149
rect 1246 1153 1252 1154
rect 1246 1149 1247 1153
rect 1251 1149 1252 1153
rect 1246 1148 1252 1149
rect 1398 1153 1404 1154
rect 1398 1149 1399 1153
rect 1403 1149 1404 1153
rect 1398 1148 1404 1149
rect 1542 1153 1548 1154
rect 1542 1149 1543 1153
rect 1547 1149 1548 1153
rect 1542 1148 1548 1149
rect 1686 1153 1692 1154
rect 1686 1149 1687 1153
rect 1691 1149 1692 1153
rect 1686 1148 1692 1149
rect 1838 1153 1844 1154
rect 1838 1149 1839 1153
rect 1843 1149 1844 1153
rect 1838 1148 1844 1149
rect 2006 1152 2012 1153
rect 2006 1148 2007 1152
rect 2011 1148 2012 1152
rect 2046 1152 2047 1156
rect 2051 1152 2052 1156
rect 2310 1153 2311 1157
rect 2315 1153 2316 1157
rect 2310 1152 2316 1153
rect 2414 1157 2420 1158
rect 2414 1153 2415 1157
rect 2419 1153 2420 1157
rect 2414 1152 2420 1153
rect 2526 1157 2532 1158
rect 2526 1153 2527 1157
rect 2531 1153 2532 1157
rect 2526 1152 2532 1153
rect 2638 1157 2644 1158
rect 2638 1153 2639 1157
rect 2643 1153 2644 1157
rect 2638 1152 2644 1153
rect 2766 1157 2772 1158
rect 2766 1153 2767 1157
rect 2771 1153 2772 1157
rect 2766 1152 2772 1153
rect 2910 1157 2916 1158
rect 2910 1153 2911 1157
rect 2915 1153 2916 1157
rect 2910 1152 2916 1153
rect 3070 1157 3076 1158
rect 3070 1153 3071 1157
rect 3075 1153 3076 1157
rect 3070 1152 3076 1153
rect 3246 1157 3252 1158
rect 3246 1153 3247 1157
rect 3251 1153 3252 1157
rect 3246 1152 3252 1153
rect 3438 1157 3444 1158
rect 3438 1153 3439 1157
rect 3443 1153 3444 1157
rect 3438 1152 3444 1153
rect 3630 1157 3636 1158
rect 3630 1153 3631 1157
rect 3635 1153 3636 1157
rect 3630 1152 3636 1153
rect 3830 1157 3836 1158
rect 3830 1153 3831 1157
rect 3835 1153 3836 1157
rect 3830 1152 3836 1153
rect 3942 1156 3948 1157
rect 3942 1152 3943 1156
rect 3947 1152 3948 1156
rect 2046 1151 2052 1152
rect 110 1147 116 1148
rect 112 1123 114 1147
rect 424 1123 426 1148
rect 592 1123 594 1148
rect 760 1123 762 1148
rect 928 1123 930 1148
rect 1096 1123 1098 1148
rect 1248 1123 1250 1148
rect 1400 1123 1402 1148
rect 1544 1123 1546 1148
rect 1688 1123 1690 1148
rect 1840 1123 1842 1148
rect 2006 1147 2012 1148
rect 2008 1123 2010 1147
rect 2048 1127 2050 1151
rect 2312 1127 2314 1152
rect 2416 1127 2418 1152
rect 2528 1127 2530 1152
rect 2640 1127 2642 1152
rect 2768 1127 2770 1152
rect 2912 1127 2914 1152
rect 3072 1127 3074 1152
rect 3248 1127 3250 1152
rect 3440 1127 3442 1152
rect 3632 1127 3634 1152
rect 3832 1127 3834 1152
rect 3942 1151 3948 1152
rect 3944 1127 3946 1151
rect 2047 1126 2051 1127
rect 111 1122 115 1123
rect 111 1117 115 1118
rect 375 1122 379 1123
rect 375 1117 379 1118
rect 423 1122 427 1123
rect 423 1117 427 1118
rect 487 1122 491 1123
rect 487 1117 491 1118
rect 591 1122 595 1123
rect 591 1117 595 1118
rect 599 1122 603 1123
rect 599 1117 603 1118
rect 711 1122 715 1123
rect 711 1117 715 1118
rect 759 1122 763 1123
rect 759 1117 763 1118
rect 831 1122 835 1123
rect 831 1117 835 1118
rect 927 1122 931 1123
rect 927 1117 931 1118
rect 967 1122 971 1123
rect 967 1117 971 1118
rect 1095 1122 1099 1123
rect 1095 1117 1099 1118
rect 1119 1122 1123 1123
rect 1119 1117 1123 1118
rect 1247 1122 1251 1123
rect 1247 1117 1251 1118
rect 1279 1122 1283 1123
rect 1279 1117 1283 1118
rect 1399 1122 1403 1123
rect 1399 1117 1403 1118
rect 1447 1122 1451 1123
rect 1447 1117 1451 1118
rect 1543 1122 1547 1123
rect 1543 1117 1547 1118
rect 1623 1122 1627 1123
rect 1623 1117 1627 1118
rect 1687 1122 1691 1123
rect 1687 1117 1691 1118
rect 1839 1122 1843 1123
rect 1839 1117 1843 1118
rect 2007 1122 2011 1123
rect 2047 1121 2051 1122
rect 2311 1126 2315 1127
rect 2311 1121 2315 1122
rect 2407 1126 2411 1127
rect 2407 1121 2411 1122
rect 2415 1126 2419 1127
rect 2415 1121 2419 1122
rect 2503 1126 2507 1127
rect 2503 1121 2507 1122
rect 2527 1126 2531 1127
rect 2527 1121 2531 1122
rect 2599 1126 2603 1127
rect 2599 1121 2603 1122
rect 2639 1126 2643 1127
rect 2639 1121 2643 1122
rect 2695 1126 2699 1127
rect 2695 1121 2699 1122
rect 2767 1126 2771 1127
rect 2767 1121 2771 1122
rect 2807 1126 2811 1127
rect 2807 1121 2811 1122
rect 2911 1126 2915 1127
rect 2911 1121 2915 1122
rect 2943 1126 2947 1127
rect 2943 1121 2947 1122
rect 3071 1126 3075 1127
rect 3071 1121 3075 1122
rect 3095 1126 3099 1127
rect 3095 1121 3099 1122
rect 3247 1126 3251 1127
rect 3247 1121 3251 1122
rect 3263 1126 3267 1127
rect 3263 1121 3267 1122
rect 3439 1126 3443 1127
rect 3439 1121 3443 1122
rect 3447 1126 3451 1127
rect 3447 1121 3451 1122
rect 3631 1126 3635 1127
rect 3631 1121 3635 1122
rect 3639 1126 3643 1127
rect 3639 1121 3643 1122
rect 3831 1126 3835 1127
rect 3831 1121 3835 1122
rect 3839 1126 3843 1127
rect 3839 1121 3843 1122
rect 3943 1126 3947 1127
rect 3943 1121 3947 1122
rect 2007 1117 2011 1118
rect 112 1097 114 1117
rect 110 1096 116 1097
rect 376 1096 378 1117
rect 488 1096 490 1117
rect 600 1096 602 1117
rect 712 1096 714 1117
rect 832 1096 834 1117
rect 968 1096 970 1117
rect 1120 1096 1122 1117
rect 1280 1096 1282 1117
rect 1448 1096 1450 1117
rect 1624 1096 1626 1117
rect 2008 1097 2010 1117
rect 2048 1101 2050 1121
rect 2046 1100 2052 1101
rect 2408 1100 2410 1121
rect 2504 1100 2506 1121
rect 2600 1100 2602 1121
rect 2696 1100 2698 1121
rect 2808 1100 2810 1121
rect 2944 1100 2946 1121
rect 3096 1100 3098 1121
rect 3264 1100 3266 1121
rect 3448 1100 3450 1121
rect 3640 1100 3642 1121
rect 3840 1100 3842 1121
rect 3944 1101 3946 1121
rect 3942 1100 3948 1101
rect 2006 1096 2012 1097
rect 110 1092 111 1096
rect 115 1092 116 1096
rect 110 1091 116 1092
rect 374 1095 380 1096
rect 374 1091 375 1095
rect 379 1091 380 1095
rect 374 1090 380 1091
rect 486 1095 492 1096
rect 486 1091 487 1095
rect 491 1091 492 1095
rect 486 1090 492 1091
rect 598 1095 604 1096
rect 598 1091 599 1095
rect 603 1091 604 1095
rect 598 1090 604 1091
rect 710 1095 716 1096
rect 710 1091 711 1095
rect 715 1091 716 1095
rect 710 1090 716 1091
rect 830 1095 836 1096
rect 830 1091 831 1095
rect 835 1091 836 1095
rect 830 1090 836 1091
rect 966 1095 972 1096
rect 966 1091 967 1095
rect 971 1091 972 1095
rect 966 1090 972 1091
rect 1118 1095 1124 1096
rect 1118 1091 1119 1095
rect 1123 1091 1124 1095
rect 1118 1090 1124 1091
rect 1278 1095 1284 1096
rect 1278 1091 1279 1095
rect 1283 1091 1284 1095
rect 1278 1090 1284 1091
rect 1446 1095 1452 1096
rect 1446 1091 1447 1095
rect 1451 1091 1452 1095
rect 1446 1090 1452 1091
rect 1622 1095 1628 1096
rect 1622 1091 1623 1095
rect 1627 1091 1628 1095
rect 2006 1092 2007 1096
rect 2011 1092 2012 1096
rect 2046 1096 2047 1100
rect 2051 1096 2052 1100
rect 2046 1095 2052 1096
rect 2406 1099 2412 1100
rect 2406 1095 2407 1099
rect 2411 1095 2412 1099
rect 2406 1094 2412 1095
rect 2502 1099 2508 1100
rect 2502 1095 2503 1099
rect 2507 1095 2508 1099
rect 2502 1094 2508 1095
rect 2598 1099 2604 1100
rect 2598 1095 2599 1099
rect 2603 1095 2604 1099
rect 2598 1094 2604 1095
rect 2694 1099 2700 1100
rect 2694 1095 2695 1099
rect 2699 1095 2700 1099
rect 2694 1094 2700 1095
rect 2806 1099 2812 1100
rect 2806 1095 2807 1099
rect 2811 1095 2812 1099
rect 2806 1094 2812 1095
rect 2942 1099 2948 1100
rect 2942 1095 2943 1099
rect 2947 1095 2948 1099
rect 2942 1094 2948 1095
rect 3094 1099 3100 1100
rect 3094 1095 3095 1099
rect 3099 1095 3100 1099
rect 3094 1094 3100 1095
rect 3262 1099 3268 1100
rect 3262 1095 3263 1099
rect 3267 1095 3268 1099
rect 3262 1094 3268 1095
rect 3446 1099 3452 1100
rect 3446 1095 3447 1099
rect 3451 1095 3452 1099
rect 3446 1094 3452 1095
rect 3638 1099 3644 1100
rect 3638 1095 3639 1099
rect 3643 1095 3644 1099
rect 3638 1094 3644 1095
rect 3838 1099 3844 1100
rect 3838 1095 3839 1099
rect 3843 1095 3844 1099
rect 3942 1096 3943 1100
rect 3947 1096 3948 1100
rect 3942 1095 3948 1096
rect 3838 1094 3844 1095
rect 2006 1091 2012 1092
rect 1622 1090 1628 1091
rect 2046 1083 2052 1084
rect 110 1079 116 1080
rect 110 1075 111 1079
rect 115 1075 116 1079
rect 2006 1079 2012 1080
rect 110 1074 116 1075
rect 374 1076 380 1077
rect 112 1047 114 1074
rect 374 1072 375 1076
rect 379 1072 380 1076
rect 374 1071 380 1072
rect 486 1076 492 1077
rect 486 1072 487 1076
rect 491 1072 492 1076
rect 486 1071 492 1072
rect 598 1076 604 1077
rect 598 1072 599 1076
rect 603 1072 604 1076
rect 598 1071 604 1072
rect 710 1076 716 1077
rect 710 1072 711 1076
rect 715 1072 716 1076
rect 710 1071 716 1072
rect 830 1076 836 1077
rect 830 1072 831 1076
rect 835 1072 836 1076
rect 830 1071 836 1072
rect 966 1076 972 1077
rect 966 1072 967 1076
rect 971 1072 972 1076
rect 966 1071 972 1072
rect 1118 1076 1124 1077
rect 1118 1072 1119 1076
rect 1123 1072 1124 1076
rect 1118 1071 1124 1072
rect 1278 1076 1284 1077
rect 1278 1072 1279 1076
rect 1283 1072 1284 1076
rect 1278 1071 1284 1072
rect 1446 1076 1452 1077
rect 1446 1072 1447 1076
rect 1451 1072 1452 1076
rect 1446 1071 1452 1072
rect 1622 1076 1628 1077
rect 1622 1072 1623 1076
rect 1627 1072 1628 1076
rect 2006 1075 2007 1079
rect 2011 1075 2012 1079
rect 2046 1079 2047 1083
rect 2051 1079 2052 1083
rect 3942 1083 3948 1084
rect 2046 1078 2052 1079
rect 2406 1080 2412 1081
rect 2006 1074 2012 1075
rect 1622 1071 1628 1072
rect 376 1047 378 1071
rect 488 1047 490 1071
rect 600 1047 602 1071
rect 712 1047 714 1071
rect 832 1047 834 1071
rect 968 1047 970 1071
rect 1120 1047 1122 1071
rect 1280 1047 1282 1071
rect 1448 1047 1450 1071
rect 1624 1047 1626 1071
rect 2008 1047 2010 1074
rect 2048 1047 2050 1078
rect 2406 1076 2407 1080
rect 2411 1076 2412 1080
rect 2406 1075 2412 1076
rect 2502 1080 2508 1081
rect 2502 1076 2503 1080
rect 2507 1076 2508 1080
rect 2502 1075 2508 1076
rect 2598 1080 2604 1081
rect 2598 1076 2599 1080
rect 2603 1076 2604 1080
rect 2598 1075 2604 1076
rect 2694 1080 2700 1081
rect 2694 1076 2695 1080
rect 2699 1076 2700 1080
rect 2694 1075 2700 1076
rect 2806 1080 2812 1081
rect 2806 1076 2807 1080
rect 2811 1076 2812 1080
rect 2806 1075 2812 1076
rect 2942 1080 2948 1081
rect 2942 1076 2943 1080
rect 2947 1076 2948 1080
rect 2942 1075 2948 1076
rect 3094 1080 3100 1081
rect 3094 1076 3095 1080
rect 3099 1076 3100 1080
rect 3094 1075 3100 1076
rect 3262 1080 3268 1081
rect 3262 1076 3263 1080
rect 3267 1076 3268 1080
rect 3262 1075 3268 1076
rect 3446 1080 3452 1081
rect 3446 1076 3447 1080
rect 3451 1076 3452 1080
rect 3446 1075 3452 1076
rect 3638 1080 3644 1081
rect 3638 1076 3639 1080
rect 3643 1076 3644 1080
rect 3638 1075 3644 1076
rect 3838 1080 3844 1081
rect 3838 1076 3839 1080
rect 3843 1076 3844 1080
rect 3942 1079 3943 1083
rect 3947 1079 3948 1083
rect 3942 1078 3948 1079
rect 3838 1075 3844 1076
rect 2408 1047 2410 1075
rect 2504 1047 2506 1075
rect 2600 1047 2602 1075
rect 2696 1047 2698 1075
rect 2808 1047 2810 1075
rect 2944 1047 2946 1075
rect 3096 1047 3098 1075
rect 3264 1047 3266 1075
rect 3448 1047 3450 1075
rect 3640 1047 3642 1075
rect 3840 1047 3842 1075
rect 3944 1047 3946 1078
rect 111 1046 115 1047
rect 111 1041 115 1042
rect 303 1046 307 1047
rect 303 1041 307 1042
rect 375 1046 379 1047
rect 375 1041 379 1042
rect 447 1046 451 1047
rect 447 1041 451 1042
rect 487 1046 491 1047
rect 487 1041 491 1042
rect 591 1046 595 1047
rect 591 1041 595 1042
rect 599 1046 603 1047
rect 599 1041 603 1042
rect 711 1046 715 1047
rect 711 1041 715 1042
rect 727 1046 731 1047
rect 727 1041 731 1042
rect 831 1046 835 1047
rect 831 1041 835 1042
rect 855 1046 859 1047
rect 855 1041 859 1042
rect 967 1046 971 1047
rect 967 1041 971 1042
rect 975 1046 979 1047
rect 975 1041 979 1042
rect 1087 1046 1091 1047
rect 1087 1041 1091 1042
rect 1119 1046 1123 1047
rect 1119 1041 1123 1042
rect 1199 1046 1203 1047
rect 1199 1041 1203 1042
rect 1279 1046 1283 1047
rect 1279 1041 1283 1042
rect 1311 1046 1315 1047
rect 1311 1041 1315 1042
rect 1431 1046 1435 1047
rect 1431 1041 1435 1042
rect 1447 1046 1451 1047
rect 1447 1041 1451 1042
rect 1623 1046 1627 1047
rect 1623 1041 1627 1042
rect 2007 1046 2011 1047
rect 2007 1041 2011 1042
rect 2047 1046 2051 1047
rect 2047 1041 2051 1042
rect 2407 1046 2411 1047
rect 2407 1041 2411 1042
rect 2455 1046 2459 1047
rect 2455 1041 2459 1042
rect 2503 1046 2507 1047
rect 2503 1041 2507 1042
rect 2551 1046 2555 1047
rect 2551 1041 2555 1042
rect 2599 1046 2603 1047
rect 2599 1041 2603 1042
rect 2647 1046 2651 1047
rect 2647 1041 2651 1042
rect 2695 1046 2699 1047
rect 2695 1041 2699 1042
rect 2759 1046 2763 1047
rect 2759 1041 2763 1042
rect 2807 1046 2811 1047
rect 2807 1041 2811 1042
rect 2887 1046 2891 1047
rect 2887 1041 2891 1042
rect 2943 1046 2947 1047
rect 2943 1041 2947 1042
rect 3031 1046 3035 1047
rect 3031 1041 3035 1042
rect 3095 1046 3099 1047
rect 3095 1041 3099 1042
rect 3183 1046 3187 1047
rect 3183 1041 3187 1042
rect 3263 1046 3267 1047
rect 3263 1041 3267 1042
rect 3343 1046 3347 1047
rect 3343 1041 3347 1042
rect 3447 1046 3451 1047
rect 3447 1041 3451 1042
rect 3503 1046 3507 1047
rect 3503 1041 3507 1042
rect 3639 1046 3643 1047
rect 3639 1041 3643 1042
rect 3671 1046 3675 1047
rect 3671 1041 3675 1042
rect 3839 1046 3843 1047
rect 3839 1041 3843 1042
rect 3943 1046 3947 1047
rect 3943 1041 3947 1042
rect 112 1014 114 1041
rect 304 1017 306 1041
rect 448 1017 450 1041
rect 592 1017 594 1041
rect 728 1017 730 1041
rect 856 1017 858 1041
rect 976 1017 978 1041
rect 1088 1017 1090 1041
rect 1200 1017 1202 1041
rect 1312 1017 1314 1041
rect 1432 1017 1434 1041
rect 302 1016 308 1017
rect 110 1013 116 1014
rect 110 1009 111 1013
rect 115 1009 116 1013
rect 302 1012 303 1016
rect 307 1012 308 1016
rect 302 1011 308 1012
rect 446 1016 452 1017
rect 446 1012 447 1016
rect 451 1012 452 1016
rect 446 1011 452 1012
rect 590 1016 596 1017
rect 590 1012 591 1016
rect 595 1012 596 1016
rect 590 1011 596 1012
rect 726 1016 732 1017
rect 726 1012 727 1016
rect 731 1012 732 1016
rect 726 1011 732 1012
rect 854 1016 860 1017
rect 854 1012 855 1016
rect 859 1012 860 1016
rect 854 1011 860 1012
rect 974 1016 980 1017
rect 974 1012 975 1016
rect 979 1012 980 1016
rect 974 1011 980 1012
rect 1086 1016 1092 1017
rect 1086 1012 1087 1016
rect 1091 1012 1092 1016
rect 1086 1011 1092 1012
rect 1198 1016 1204 1017
rect 1198 1012 1199 1016
rect 1203 1012 1204 1016
rect 1198 1011 1204 1012
rect 1310 1016 1316 1017
rect 1310 1012 1311 1016
rect 1315 1012 1316 1016
rect 1310 1011 1316 1012
rect 1430 1016 1436 1017
rect 1430 1012 1431 1016
rect 1435 1012 1436 1016
rect 2008 1014 2010 1041
rect 2048 1014 2050 1041
rect 2456 1017 2458 1041
rect 2552 1017 2554 1041
rect 2648 1017 2650 1041
rect 2760 1017 2762 1041
rect 2888 1017 2890 1041
rect 3032 1017 3034 1041
rect 3184 1017 3186 1041
rect 3344 1017 3346 1041
rect 3504 1017 3506 1041
rect 3672 1017 3674 1041
rect 3840 1017 3842 1041
rect 2454 1016 2460 1017
rect 1430 1011 1436 1012
rect 2006 1013 2012 1014
rect 110 1008 116 1009
rect 2006 1009 2007 1013
rect 2011 1009 2012 1013
rect 2006 1008 2012 1009
rect 2046 1013 2052 1014
rect 2046 1009 2047 1013
rect 2051 1009 2052 1013
rect 2454 1012 2455 1016
rect 2459 1012 2460 1016
rect 2454 1011 2460 1012
rect 2550 1016 2556 1017
rect 2550 1012 2551 1016
rect 2555 1012 2556 1016
rect 2550 1011 2556 1012
rect 2646 1016 2652 1017
rect 2646 1012 2647 1016
rect 2651 1012 2652 1016
rect 2646 1011 2652 1012
rect 2758 1016 2764 1017
rect 2758 1012 2759 1016
rect 2763 1012 2764 1016
rect 2758 1011 2764 1012
rect 2886 1016 2892 1017
rect 2886 1012 2887 1016
rect 2891 1012 2892 1016
rect 2886 1011 2892 1012
rect 3030 1016 3036 1017
rect 3030 1012 3031 1016
rect 3035 1012 3036 1016
rect 3030 1011 3036 1012
rect 3182 1016 3188 1017
rect 3182 1012 3183 1016
rect 3187 1012 3188 1016
rect 3182 1011 3188 1012
rect 3342 1016 3348 1017
rect 3342 1012 3343 1016
rect 3347 1012 3348 1016
rect 3342 1011 3348 1012
rect 3502 1016 3508 1017
rect 3502 1012 3503 1016
rect 3507 1012 3508 1016
rect 3502 1011 3508 1012
rect 3670 1016 3676 1017
rect 3670 1012 3671 1016
rect 3675 1012 3676 1016
rect 3670 1011 3676 1012
rect 3838 1016 3844 1017
rect 3838 1012 3839 1016
rect 3843 1012 3844 1016
rect 3944 1014 3946 1041
rect 3838 1011 3844 1012
rect 3942 1013 3948 1014
rect 2046 1008 2052 1009
rect 3942 1009 3943 1013
rect 3947 1009 3948 1013
rect 3942 1008 3948 1009
rect 302 997 308 998
rect 110 996 116 997
rect 110 992 111 996
rect 115 992 116 996
rect 302 993 303 997
rect 307 993 308 997
rect 302 992 308 993
rect 446 997 452 998
rect 446 993 447 997
rect 451 993 452 997
rect 446 992 452 993
rect 590 997 596 998
rect 590 993 591 997
rect 595 993 596 997
rect 590 992 596 993
rect 726 997 732 998
rect 726 993 727 997
rect 731 993 732 997
rect 726 992 732 993
rect 854 997 860 998
rect 854 993 855 997
rect 859 993 860 997
rect 854 992 860 993
rect 974 997 980 998
rect 974 993 975 997
rect 979 993 980 997
rect 974 992 980 993
rect 1086 997 1092 998
rect 1086 993 1087 997
rect 1091 993 1092 997
rect 1086 992 1092 993
rect 1198 997 1204 998
rect 1198 993 1199 997
rect 1203 993 1204 997
rect 1198 992 1204 993
rect 1310 997 1316 998
rect 1310 993 1311 997
rect 1315 993 1316 997
rect 1310 992 1316 993
rect 1430 997 1436 998
rect 2454 997 2460 998
rect 1430 993 1431 997
rect 1435 993 1436 997
rect 1430 992 1436 993
rect 2006 996 2012 997
rect 2006 992 2007 996
rect 2011 992 2012 996
rect 110 991 116 992
rect 112 971 114 991
rect 304 971 306 992
rect 448 971 450 992
rect 592 971 594 992
rect 728 971 730 992
rect 856 971 858 992
rect 976 971 978 992
rect 1088 971 1090 992
rect 1200 971 1202 992
rect 1312 971 1314 992
rect 1432 971 1434 992
rect 2006 991 2012 992
rect 2046 996 2052 997
rect 2046 992 2047 996
rect 2051 992 2052 996
rect 2454 993 2455 997
rect 2459 993 2460 997
rect 2454 992 2460 993
rect 2550 997 2556 998
rect 2550 993 2551 997
rect 2555 993 2556 997
rect 2550 992 2556 993
rect 2646 997 2652 998
rect 2646 993 2647 997
rect 2651 993 2652 997
rect 2646 992 2652 993
rect 2758 997 2764 998
rect 2758 993 2759 997
rect 2763 993 2764 997
rect 2758 992 2764 993
rect 2886 997 2892 998
rect 2886 993 2887 997
rect 2891 993 2892 997
rect 2886 992 2892 993
rect 3030 997 3036 998
rect 3030 993 3031 997
rect 3035 993 3036 997
rect 3030 992 3036 993
rect 3182 997 3188 998
rect 3182 993 3183 997
rect 3187 993 3188 997
rect 3182 992 3188 993
rect 3342 997 3348 998
rect 3342 993 3343 997
rect 3347 993 3348 997
rect 3342 992 3348 993
rect 3502 997 3508 998
rect 3502 993 3503 997
rect 3507 993 3508 997
rect 3502 992 3508 993
rect 3670 997 3676 998
rect 3670 993 3671 997
rect 3675 993 3676 997
rect 3670 992 3676 993
rect 3838 997 3844 998
rect 3838 993 3839 997
rect 3843 993 3844 997
rect 3838 992 3844 993
rect 3942 996 3948 997
rect 3942 992 3943 996
rect 3947 992 3948 996
rect 2046 991 2052 992
rect 2008 971 2010 991
rect 111 970 115 971
rect 111 965 115 966
rect 255 970 259 971
rect 255 965 259 966
rect 303 970 307 971
rect 303 965 307 966
rect 447 970 451 971
rect 447 965 451 966
rect 591 970 595 971
rect 591 965 595 966
rect 631 970 635 971
rect 631 965 635 966
rect 727 970 731 971
rect 727 965 731 966
rect 807 970 811 971
rect 807 965 811 966
rect 855 970 859 971
rect 855 965 859 966
rect 975 970 979 971
rect 975 965 979 966
rect 1087 970 1091 971
rect 1087 965 1091 966
rect 1127 970 1131 971
rect 1127 965 1131 966
rect 1199 970 1203 971
rect 1199 965 1203 966
rect 1271 970 1275 971
rect 1271 965 1275 966
rect 1311 970 1315 971
rect 1311 965 1315 966
rect 1415 970 1419 971
rect 1415 965 1419 966
rect 1431 970 1435 971
rect 1431 965 1435 966
rect 1551 970 1555 971
rect 1551 965 1555 966
rect 1695 970 1699 971
rect 1695 965 1699 966
rect 2007 970 2011 971
rect 2048 967 2050 991
rect 2456 967 2458 992
rect 2552 967 2554 992
rect 2648 967 2650 992
rect 2760 967 2762 992
rect 2888 967 2890 992
rect 3032 967 3034 992
rect 3184 967 3186 992
rect 3344 967 3346 992
rect 3504 967 3506 992
rect 3672 967 3674 992
rect 3840 967 3842 992
rect 3942 991 3948 992
rect 3944 967 3946 991
rect 2007 965 2011 966
rect 2047 966 2051 967
rect 112 945 114 965
rect 110 944 116 945
rect 256 944 258 965
rect 448 944 450 965
rect 632 944 634 965
rect 808 944 810 965
rect 976 944 978 965
rect 1128 944 1130 965
rect 1272 944 1274 965
rect 1416 944 1418 965
rect 1552 944 1554 965
rect 1696 944 1698 965
rect 2008 945 2010 965
rect 2047 961 2051 962
rect 2423 966 2427 967
rect 2423 961 2427 962
rect 2455 966 2459 967
rect 2455 961 2459 962
rect 2519 966 2523 967
rect 2519 961 2523 962
rect 2551 966 2555 967
rect 2551 961 2555 962
rect 2615 966 2619 967
rect 2615 961 2619 962
rect 2647 966 2651 967
rect 2647 961 2651 962
rect 2711 966 2715 967
rect 2711 961 2715 962
rect 2759 966 2763 967
rect 2759 961 2763 962
rect 2823 966 2827 967
rect 2823 961 2827 962
rect 2887 966 2891 967
rect 2887 961 2891 962
rect 2951 966 2955 967
rect 2951 961 2955 962
rect 3031 966 3035 967
rect 3031 961 3035 962
rect 3103 966 3107 967
rect 3103 961 3107 962
rect 3183 966 3187 967
rect 3183 961 3187 962
rect 3271 966 3275 967
rect 3271 961 3275 962
rect 3343 966 3347 967
rect 3343 961 3347 962
rect 3455 966 3459 967
rect 3455 961 3459 962
rect 3503 966 3507 967
rect 3503 961 3507 962
rect 3647 966 3651 967
rect 3647 961 3651 962
rect 3671 966 3675 967
rect 3671 961 3675 962
rect 3839 966 3843 967
rect 3839 961 3843 962
rect 3943 966 3947 967
rect 3943 961 3947 962
rect 2006 944 2012 945
rect 110 940 111 944
rect 115 940 116 944
rect 110 939 116 940
rect 254 943 260 944
rect 254 939 255 943
rect 259 939 260 943
rect 254 938 260 939
rect 446 943 452 944
rect 446 939 447 943
rect 451 939 452 943
rect 446 938 452 939
rect 630 943 636 944
rect 630 939 631 943
rect 635 939 636 943
rect 630 938 636 939
rect 806 943 812 944
rect 806 939 807 943
rect 811 939 812 943
rect 806 938 812 939
rect 974 943 980 944
rect 974 939 975 943
rect 979 939 980 943
rect 974 938 980 939
rect 1126 943 1132 944
rect 1126 939 1127 943
rect 1131 939 1132 943
rect 1126 938 1132 939
rect 1270 943 1276 944
rect 1270 939 1271 943
rect 1275 939 1276 943
rect 1270 938 1276 939
rect 1414 943 1420 944
rect 1414 939 1415 943
rect 1419 939 1420 943
rect 1414 938 1420 939
rect 1550 943 1556 944
rect 1550 939 1551 943
rect 1555 939 1556 943
rect 1550 938 1556 939
rect 1694 943 1700 944
rect 1694 939 1695 943
rect 1699 939 1700 943
rect 2006 940 2007 944
rect 2011 940 2012 944
rect 2048 941 2050 961
rect 2006 939 2012 940
rect 2046 940 2052 941
rect 2424 940 2426 961
rect 2520 940 2522 961
rect 2616 940 2618 961
rect 2712 940 2714 961
rect 2824 940 2826 961
rect 2952 940 2954 961
rect 3104 940 3106 961
rect 3272 940 3274 961
rect 3456 940 3458 961
rect 3648 940 3650 961
rect 3840 940 3842 961
rect 3944 941 3946 961
rect 3942 940 3948 941
rect 1694 938 1700 939
rect 2046 936 2047 940
rect 2051 936 2052 940
rect 2046 935 2052 936
rect 2422 939 2428 940
rect 2422 935 2423 939
rect 2427 935 2428 939
rect 2422 934 2428 935
rect 2518 939 2524 940
rect 2518 935 2519 939
rect 2523 935 2524 939
rect 2518 934 2524 935
rect 2614 939 2620 940
rect 2614 935 2615 939
rect 2619 935 2620 939
rect 2614 934 2620 935
rect 2710 939 2716 940
rect 2710 935 2711 939
rect 2715 935 2716 939
rect 2710 934 2716 935
rect 2822 939 2828 940
rect 2822 935 2823 939
rect 2827 935 2828 939
rect 2822 934 2828 935
rect 2950 939 2956 940
rect 2950 935 2951 939
rect 2955 935 2956 939
rect 2950 934 2956 935
rect 3102 939 3108 940
rect 3102 935 3103 939
rect 3107 935 3108 939
rect 3102 934 3108 935
rect 3270 939 3276 940
rect 3270 935 3271 939
rect 3275 935 3276 939
rect 3270 934 3276 935
rect 3454 939 3460 940
rect 3454 935 3455 939
rect 3459 935 3460 939
rect 3454 934 3460 935
rect 3646 939 3652 940
rect 3646 935 3647 939
rect 3651 935 3652 939
rect 3646 934 3652 935
rect 3838 939 3844 940
rect 3838 935 3839 939
rect 3843 935 3844 939
rect 3942 936 3943 940
rect 3947 936 3948 940
rect 3942 935 3948 936
rect 3838 934 3844 935
rect 110 927 116 928
rect 110 923 111 927
rect 115 923 116 927
rect 2006 927 2012 928
rect 110 922 116 923
rect 254 924 260 925
rect 112 891 114 922
rect 254 920 255 924
rect 259 920 260 924
rect 254 919 260 920
rect 446 924 452 925
rect 446 920 447 924
rect 451 920 452 924
rect 446 919 452 920
rect 630 924 636 925
rect 630 920 631 924
rect 635 920 636 924
rect 630 919 636 920
rect 806 924 812 925
rect 806 920 807 924
rect 811 920 812 924
rect 806 919 812 920
rect 974 924 980 925
rect 974 920 975 924
rect 979 920 980 924
rect 974 919 980 920
rect 1126 924 1132 925
rect 1126 920 1127 924
rect 1131 920 1132 924
rect 1126 919 1132 920
rect 1270 924 1276 925
rect 1270 920 1271 924
rect 1275 920 1276 924
rect 1270 919 1276 920
rect 1414 924 1420 925
rect 1414 920 1415 924
rect 1419 920 1420 924
rect 1414 919 1420 920
rect 1550 924 1556 925
rect 1550 920 1551 924
rect 1555 920 1556 924
rect 1550 919 1556 920
rect 1694 924 1700 925
rect 1694 920 1695 924
rect 1699 920 1700 924
rect 2006 923 2007 927
rect 2011 923 2012 927
rect 2006 922 2012 923
rect 2046 923 2052 924
rect 1694 919 1700 920
rect 256 891 258 919
rect 448 891 450 919
rect 632 891 634 919
rect 808 891 810 919
rect 976 891 978 919
rect 1128 891 1130 919
rect 1272 891 1274 919
rect 1416 891 1418 919
rect 1552 891 1554 919
rect 1696 891 1698 919
rect 2008 891 2010 922
rect 2046 919 2047 923
rect 2051 919 2052 923
rect 3942 923 3948 924
rect 2046 918 2052 919
rect 2422 920 2428 921
rect 2048 891 2050 918
rect 2422 916 2423 920
rect 2427 916 2428 920
rect 2422 915 2428 916
rect 2518 920 2524 921
rect 2518 916 2519 920
rect 2523 916 2524 920
rect 2518 915 2524 916
rect 2614 920 2620 921
rect 2614 916 2615 920
rect 2619 916 2620 920
rect 2614 915 2620 916
rect 2710 920 2716 921
rect 2710 916 2711 920
rect 2715 916 2716 920
rect 2710 915 2716 916
rect 2822 920 2828 921
rect 2822 916 2823 920
rect 2827 916 2828 920
rect 2822 915 2828 916
rect 2950 920 2956 921
rect 2950 916 2951 920
rect 2955 916 2956 920
rect 2950 915 2956 916
rect 3102 920 3108 921
rect 3102 916 3103 920
rect 3107 916 3108 920
rect 3102 915 3108 916
rect 3270 920 3276 921
rect 3270 916 3271 920
rect 3275 916 3276 920
rect 3270 915 3276 916
rect 3454 920 3460 921
rect 3454 916 3455 920
rect 3459 916 3460 920
rect 3454 915 3460 916
rect 3646 920 3652 921
rect 3646 916 3647 920
rect 3651 916 3652 920
rect 3646 915 3652 916
rect 3838 920 3844 921
rect 3838 916 3839 920
rect 3843 916 3844 920
rect 3942 919 3943 923
rect 3947 919 3948 923
rect 3942 918 3948 919
rect 3838 915 3844 916
rect 2424 891 2426 915
rect 2520 891 2522 915
rect 2616 891 2618 915
rect 2712 891 2714 915
rect 2824 891 2826 915
rect 2952 891 2954 915
rect 3104 891 3106 915
rect 3272 891 3274 915
rect 3456 891 3458 915
rect 3648 891 3650 915
rect 3840 891 3842 915
rect 3944 891 3946 918
rect 111 890 115 891
rect 111 885 115 886
rect 255 890 259 891
rect 255 885 259 886
rect 447 890 451 891
rect 447 885 451 886
rect 631 890 635 891
rect 631 885 635 886
rect 639 890 643 891
rect 639 885 643 886
rect 807 890 811 891
rect 807 885 811 886
rect 823 890 827 891
rect 823 885 827 886
rect 975 890 979 891
rect 975 885 979 886
rect 999 890 1003 891
rect 999 885 1003 886
rect 1127 890 1131 891
rect 1127 885 1131 886
rect 1167 890 1171 891
rect 1167 885 1171 886
rect 1271 890 1275 891
rect 1271 885 1275 886
rect 1327 890 1331 891
rect 1327 885 1331 886
rect 1415 890 1419 891
rect 1415 885 1419 886
rect 1479 890 1483 891
rect 1479 885 1483 886
rect 1551 890 1555 891
rect 1551 885 1555 886
rect 1631 890 1635 891
rect 1631 885 1635 886
rect 1695 890 1699 891
rect 1695 885 1699 886
rect 1783 890 1787 891
rect 1783 885 1787 886
rect 2007 890 2011 891
rect 2007 885 2011 886
rect 2047 890 2051 891
rect 2047 885 2051 886
rect 2343 890 2347 891
rect 2343 885 2347 886
rect 2423 890 2427 891
rect 2423 885 2427 886
rect 2439 890 2443 891
rect 2439 885 2443 886
rect 2519 890 2523 891
rect 2519 885 2523 886
rect 2535 890 2539 891
rect 2535 885 2539 886
rect 2615 890 2619 891
rect 2615 885 2619 886
rect 2631 890 2635 891
rect 2631 885 2635 886
rect 2711 890 2715 891
rect 2711 885 2715 886
rect 2735 890 2739 891
rect 2735 885 2739 886
rect 2823 890 2827 891
rect 2823 885 2827 886
rect 2863 890 2867 891
rect 2863 885 2867 886
rect 2951 890 2955 891
rect 2951 885 2955 886
rect 3015 890 3019 891
rect 3015 885 3019 886
rect 3103 890 3107 891
rect 3103 885 3107 886
rect 3191 890 3195 891
rect 3191 885 3195 886
rect 3271 890 3275 891
rect 3271 885 3275 886
rect 3391 890 3395 891
rect 3391 885 3395 886
rect 3455 890 3459 891
rect 3455 885 3459 886
rect 3607 890 3611 891
rect 3607 885 3611 886
rect 3647 890 3651 891
rect 3647 885 3651 886
rect 3823 890 3827 891
rect 3823 885 3827 886
rect 3839 890 3843 891
rect 3839 885 3843 886
rect 3943 890 3947 891
rect 3943 885 3947 886
rect 112 858 114 885
rect 256 861 258 885
rect 448 861 450 885
rect 640 861 642 885
rect 824 861 826 885
rect 1000 861 1002 885
rect 1168 861 1170 885
rect 1328 861 1330 885
rect 1480 861 1482 885
rect 1632 861 1634 885
rect 1784 861 1786 885
rect 254 860 260 861
rect 110 857 116 858
rect 110 853 111 857
rect 115 853 116 857
rect 254 856 255 860
rect 259 856 260 860
rect 254 855 260 856
rect 446 860 452 861
rect 446 856 447 860
rect 451 856 452 860
rect 446 855 452 856
rect 638 860 644 861
rect 638 856 639 860
rect 643 856 644 860
rect 638 855 644 856
rect 822 860 828 861
rect 822 856 823 860
rect 827 856 828 860
rect 822 855 828 856
rect 998 860 1004 861
rect 998 856 999 860
rect 1003 856 1004 860
rect 998 855 1004 856
rect 1166 860 1172 861
rect 1166 856 1167 860
rect 1171 856 1172 860
rect 1166 855 1172 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1478 860 1484 861
rect 1478 856 1479 860
rect 1483 856 1484 860
rect 1478 855 1484 856
rect 1630 860 1636 861
rect 1630 856 1631 860
rect 1635 856 1636 860
rect 1630 855 1636 856
rect 1782 860 1788 861
rect 1782 856 1783 860
rect 1787 856 1788 860
rect 2008 858 2010 885
rect 2048 858 2050 885
rect 2344 861 2346 885
rect 2440 861 2442 885
rect 2536 861 2538 885
rect 2632 861 2634 885
rect 2736 861 2738 885
rect 2864 861 2866 885
rect 3016 861 3018 885
rect 3192 861 3194 885
rect 3392 861 3394 885
rect 3608 861 3610 885
rect 3824 861 3826 885
rect 2342 860 2348 861
rect 1782 855 1788 856
rect 2006 857 2012 858
rect 110 852 116 853
rect 2006 853 2007 857
rect 2011 853 2012 857
rect 2006 852 2012 853
rect 2046 857 2052 858
rect 2046 853 2047 857
rect 2051 853 2052 857
rect 2342 856 2343 860
rect 2347 856 2348 860
rect 2342 855 2348 856
rect 2438 860 2444 861
rect 2438 856 2439 860
rect 2443 856 2444 860
rect 2438 855 2444 856
rect 2534 860 2540 861
rect 2534 856 2535 860
rect 2539 856 2540 860
rect 2534 855 2540 856
rect 2630 860 2636 861
rect 2630 856 2631 860
rect 2635 856 2636 860
rect 2630 855 2636 856
rect 2734 860 2740 861
rect 2734 856 2735 860
rect 2739 856 2740 860
rect 2734 855 2740 856
rect 2862 860 2868 861
rect 2862 856 2863 860
rect 2867 856 2868 860
rect 2862 855 2868 856
rect 3014 860 3020 861
rect 3014 856 3015 860
rect 3019 856 3020 860
rect 3014 855 3020 856
rect 3190 860 3196 861
rect 3190 856 3191 860
rect 3195 856 3196 860
rect 3190 855 3196 856
rect 3390 860 3396 861
rect 3390 856 3391 860
rect 3395 856 3396 860
rect 3390 855 3396 856
rect 3606 860 3612 861
rect 3606 856 3607 860
rect 3611 856 3612 860
rect 3606 855 3612 856
rect 3822 860 3828 861
rect 3822 856 3823 860
rect 3827 856 3828 860
rect 3944 858 3946 885
rect 3822 855 3828 856
rect 3942 857 3948 858
rect 2046 852 2052 853
rect 3942 853 3943 857
rect 3947 853 3948 857
rect 3942 852 3948 853
rect 254 841 260 842
rect 110 840 116 841
rect 110 836 111 840
rect 115 836 116 840
rect 254 837 255 841
rect 259 837 260 841
rect 254 836 260 837
rect 446 841 452 842
rect 446 837 447 841
rect 451 837 452 841
rect 446 836 452 837
rect 638 841 644 842
rect 638 837 639 841
rect 643 837 644 841
rect 638 836 644 837
rect 822 841 828 842
rect 822 837 823 841
rect 827 837 828 841
rect 822 836 828 837
rect 998 841 1004 842
rect 998 837 999 841
rect 1003 837 1004 841
rect 998 836 1004 837
rect 1166 841 1172 842
rect 1166 837 1167 841
rect 1171 837 1172 841
rect 1166 836 1172 837
rect 1326 841 1332 842
rect 1326 837 1327 841
rect 1331 837 1332 841
rect 1326 836 1332 837
rect 1478 841 1484 842
rect 1478 837 1479 841
rect 1483 837 1484 841
rect 1478 836 1484 837
rect 1630 841 1636 842
rect 1630 837 1631 841
rect 1635 837 1636 841
rect 1630 836 1636 837
rect 1782 841 1788 842
rect 2342 841 2348 842
rect 1782 837 1783 841
rect 1787 837 1788 841
rect 1782 836 1788 837
rect 2006 840 2012 841
rect 2006 836 2007 840
rect 2011 836 2012 840
rect 110 835 116 836
rect 112 811 114 835
rect 256 811 258 836
rect 448 811 450 836
rect 640 811 642 836
rect 824 811 826 836
rect 1000 811 1002 836
rect 1168 811 1170 836
rect 1328 811 1330 836
rect 1480 811 1482 836
rect 1632 811 1634 836
rect 1784 811 1786 836
rect 2006 835 2012 836
rect 2046 840 2052 841
rect 2046 836 2047 840
rect 2051 836 2052 840
rect 2342 837 2343 841
rect 2347 837 2348 841
rect 2342 836 2348 837
rect 2438 841 2444 842
rect 2438 837 2439 841
rect 2443 837 2444 841
rect 2438 836 2444 837
rect 2534 841 2540 842
rect 2534 837 2535 841
rect 2539 837 2540 841
rect 2534 836 2540 837
rect 2630 841 2636 842
rect 2630 837 2631 841
rect 2635 837 2636 841
rect 2630 836 2636 837
rect 2734 841 2740 842
rect 2734 837 2735 841
rect 2739 837 2740 841
rect 2734 836 2740 837
rect 2862 841 2868 842
rect 2862 837 2863 841
rect 2867 837 2868 841
rect 2862 836 2868 837
rect 3014 841 3020 842
rect 3014 837 3015 841
rect 3019 837 3020 841
rect 3014 836 3020 837
rect 3190 841 3196 842
rect 3190 837 3191 841
rect 3195 837 3196 841
rect 3190 836 3196 837
rect 3390 841 3396 842
rect 3390 837 3391 841
rect 3395 837 3396 841
rect 3390 836 3396 837
rect 3606 841 3612 842
rect 3606 837 3607 841
rect 3611 837 3612 841
rect 3606 836 3612 837
rect 3822 841 3828 842
rect 3822 837 3823 841
rect 3827 837 3828 841
rect 3822 836 3828 837
rect 3942 840 3948 841
rect 3942 836 3943 840
rect 3947 836 3948 840
rect 2046 835 2052 836
rect 2008 811 2010 835
rect 2048 815 2050 835
rect 2344 815 2346 836
rect 2440 815 2442 836
rect 2536 815 2538 836
rect 2632 815 2634 836
rect 2736 815 2738 836
rect 2864 815 2866 836
rect 3016 815 3018 836
rect 3192 815 3194 836
rect 3392 815 3394 836
rect 3608 815 3610 836
rect 3824 815 3826 836
rect 3942 835 3948 836
rect 3944 815 3946 835
rect 2047 814 2051 815
rect 111 810 115 811
rect 111 805 115 806
rect 159 810 163 811
rect 159 805 163 806
rect 255 810 259 811
rect 255 805 259 806
rect 311 810 315 811
rect 311 805 315 806
rect 447 810 451 811
rect 447 805 451 806
rect 471 810 475 811
rect 471 805 475 806
rect 623 810 627 811
rect 623 805 627 806
rect 639 810 643 811
rect 639 805 643 806
rect 775 810 779 811
rect 775 805 779 806
rect 823 810 827 811
rect 823 805 827 806
rect 935 810 939 811
rect 935 805 939 806
rect 999 810 1003 811
rect 999 805 1003 806
rect 1095 810 1099 811
rect 1095 805 1099 806
rect 1167 810 1171 811
rect 1167 805 1171 806
rect 1255 810 1259 811
rect 1255 805 1259 806
rect 1327 810 1331 811
rect 1327 805 1331 806
rect 1415 810 1419 811
rect 1415 805 1419 806
rect 1479 810 1483 811
rect 1479 805 1483 806
rect 1583 810 1587 811
rect 1583 805 1587 806
rect 1631 810 1635 811
rect 1631 805 1635 806
rect 1751 810 1755 811
rect 1751 805 1755 806
rect 1783 810 1787 811
rect 1783 805 1787 806
rect 1903 810 1907 811
rect 1903 805 1907 806
rect 2007 810 2011 811
rect 2047 809 2051 810
rect 2311 814 2315 815
rect 2311 809 2315 810
rect 2343 814 2347 815
rect 2343 809 2347 810
rect 2439 814 2443 815
rect 2439 809 2443 810
rect 2495 814 2499 815
rect 2495 809 2499 810
rect 2535 814 2539 815
rect 2535 809 2539 810
rect 2631 814 2635 815
rect 2631 809 2635 810
rect 2687 814 2691 815
rect 2687 809 2691 810
rect 2735 814 2739 815
rect 2735 809 2739 810
rect 2863 814 2867 815
rect 2863 809 2867 810
rect 2879 814 2883 815
rect 2879 809 2883 810
rect 3015 814 3019 815
rect 3015 809 3019 810
rect 3079 814 3083 815
rect 3079 809 3083 810
rect 3191 814 3195 815
rect 3191 809 3195 810
rect 3287 814 3291 815
rect 3287 809 3291 810
rect 3391 814 3395 815
rect 3391 809 3395 810
rect 3503 814 3507 815
rect 3503 809 3507 810
rect 3607 814 3611 815
rect 3607 809 3611 810
rect 3719 814 3723 815
rect 3719 809 3723 810
rect 3823 814 3827 815
rect 3823 809 3827 810
rect 3943 814 3947 815
rect 3943 809 3947 810
rect 2007 805 2011 806
rect 112 785 114 805
rect 110 784 116 785
rect 160 784 162 805
rect 312 784 314 805
rect 472 784 474 805
rect 624 784 626 805
rect 776 784 778 805
rect 936 784 938 805
rect 1096 784 1098 805
rect 1256 784 1258 805
rect 1416 784 1418 805
rect 1584 784 1586 805
rect 1752 784 1754 805
rect 1904 784 1906 805
rect 2008 785 2010 805
rect 2048 789 2050 809
rect 2046 788 2052 789
rect 2312 788 2314 809
rect 2496 788 2498 809
rect 2688 788 2690 809
rect 2880 788 2882 809
rect 3080 788 3082 809
rect 3288 788 3290 809
rect 3504 788 3506 809
rect 3720 788 3722 809
rect 3944 789 3946 809
rect 3942 788 3948 789
rect 2006 784 2012 785
rect 110 780 111 784
rect 115 780 116 784
rect 110 779 116 780
rect 158 783 164 784
rect 158 779 159 783
rect 163 779 164 783
rect 158 778 164 779
rect 310 783 316 784
rect 310 779 311 783
rect 315 779 316 783
rect 310 778 316 779
rect 470 783 476 784
rect 470 779 471 783
rect 475 779 476 783
rect 470 778 476 779
rect 622 783 628 784
rect 622 779 623 783
rect 627 779 628 783
rect 622 778 628 779
rect 774 783 780 784
rect 774 779 775 783
rect 779 779 780 783
rect 774 778 780 779
rect 934 783 940 784
rect 934 779 935 783
rect 939 779 940 783
rect 934 778 940 779
rect 1094 783 1100 784
rect 1094 779 1095 783
rect 1099 779 1100 783
rect 1094 778 1100 779
rect 1254 783 1260 784
rect 1254 779 1255 783
rect 1259 779 1260 783
rect 1254 778 1260 779
rect 1414 783 1420 784
rect 1414 779 1415 783
rect 1419 779 1420 783
rect 1414 778 1420 779
rect 1582 783 1588 784
rect 1582 779 1583 783
rect 1587 779 1588 783
rect 1582 778 1588 779
rect 1750 783 1756 784
rect 1750 779 1751 783
rect 1755 779 1756 783
rect 1750 778 1756 779
rect 1902 783 1908 784
rect 1902 779 1903 783
rect 1907 779 1908 783
rect 2006 780 2007 784
rect 2011 780 2012 784
rect 2046 784 2047 788
rect 2051 784 2052 788
rect 2046 783 2052 784
rect 2310 787 2316 788
rect 2310 783 2311 787
rect 2315 783 2316 787
rect 2310 782 2316 783
rect 2494 787 2500 788
rect 2494 783 2495 787
rect 2499 783 2500 787
rect 2494 782 2500 783
rect 2686 787 2692 788
rect 2686 783 2687 787
rect 2691 783 2692 787
rect 2686 782 2692 783
rect 2878 787 2884 788
rect 2878 783 2879 787
rect 2883 783 2884 787
rect 2878 782 2884 783
rect 3078 787 3084 788
rect 3078 783 3079 787
rect 3083 783 3084 787
rect 3078 782 3084 783
rect 3286 787 3292 788
rect 3286 783 3287 787
rect 3291 783 3292 787
rect 3286 782 3292 783
rect 3502 787 3508 788
rect 3502 783 3503 787
rect 3507 783 3508 787
rect 3502 782 3508 783
rect 3718 787 3724 788
rect 3718 783 3719 787
rect 3723 783 3724 787
rect 3942 784 3943 788
rect 3947 784 3948 788
rect 3942 783 3948 784
rect 3718 782 3724 783
rect 2006 779 2012 780
rect 1902 778 1908 779
rect 2046 771 2052 772
rect 110 767 116 768
rect 110 763 111 767
rect 115 763 116 767
rect 2006 767 2012 768
rect 110 762 116 763
rect 158 764 164 765
rect 112 735 114 762
rect 158 760 159 764
rect 163 760 164 764
rect 158 759 164 760
rect 310 764 316 765
rect 310 760 311 764
rect 315 760 316 764
rect 310 759 316 760
rect 470 764 476 765
rect 470 760 471 764
rect 475 760 476 764
rect 470 759 476 760
rect 622 764 628 765
rect 622 760 623 764
rect 627 760 628 764
rect 622 759 628 760
rect 774 764 780 765
rect 774 760 775 764
rect 779 760 780 764
rect 774 759 780 760
rect 934 764 940 765
rect 934 760 935 764
rect 939 760 940 764
rect 934 759 940 760
rect 1094 764 1100 765
rect 1094 760 1095 764
rect 1099 760 1100 764
rect 1094 759 1100 760
rect 1254 764 1260 765
rect 1254 760 1255 764
rect 1259 760 1260 764
rect 1254 759 1260 760
rect 1414 764 1420 765
rect 1414 760 1415 764
rect 1419 760 1420 764
rect 1414 759 1420 760
rect 1582 764 1588 765
rect 1582 760 1583 764
rect 1587 760 1588 764
rect 1582 759 1588 760
rect 1750 764 1756 765
rect 1750 760 1751 764
rect 1755 760 1756 764
rect 1750 759 1756 760
rect 1902 764 1908 765
rect 1902 760 1903 764
rect 1907 760 1908 764
rect 2006 763 2007 767
rect 2011 763 2012 767
rect 2046 767 2047 771
rect 2051 767 2052 771
rect 3942 771 3948 772
rect 2046 766 2052 767
rect 2310 768 2316 769
rect 2006 762 2012 763
rect 1902 759 1908 760
rect 160 735 162 759
rect 312 735 314 759
rect 472 735 474 759
rect 624 735 626 759
rect 776 735 778 759
rect 936 735 938 759
rect 1096 735 1098 759
rect 1256 735 1258 759
rect 1416 735 1418 759
rect 1584 735 1586 759
rect 1752 735 1754 759
rect 1904 735 1906 759
rect 2008 735 2010 762
rect 2048 735 2050 766
rect 2310 764 2311 768
rect 2315 764 2316 768
rect 2310 763 2316 764
rect 2494 768 2500 769
rect 2494 764 2495 768
rect 2499 764 2500 768
rect 2494 763 2500 764
rect 2686 768 2692 769
rect 2686 764 2687 768
rect 2691 764 2692 768
rect 2686 763 2692 764
rect 2878 768 2884 769
rect 2878 764 2879 768
rect 2883 764 2884 768
rect 2878 763 2884 764
rect 3078 768 3084 769
rect 3078 764 3079 768
rect 3083 764 3084 768
rect 3078 763 3084 764
rect 3286 768 3292 769
rect 3286 764 3287 768
rect 3291 764 3292 768
rect 3286 763 3292 764
rect 3502 768 3508 769
rect 3502 764 3503 768
rect 3507 764 3508 768
rect 3502 763 3508 764
rect 3718 768 3724 769
rect 3718 764 3719 768
rect 3723 764 3724 768
rect 3942 767 3943 771
rect 3947 767 3948 771
rect 3942 766 3948 767
rect 3718 763 3724 764
rect 2312 735 2314 763
rect 2496 735 2498 763
rect 2688 735 2690 763
rect 2880 735 2882 763
rect 3080 735 3082 763
rect 3288 735 3290 763
rect 3504 735 3506 763
rect 3720 735 3722 763
rect 3944 735 3946 766
rect 111 734 115 735
rect 111 729 115 730
rect 135 734 139 735
rect 135 729 139 730
rect 159 734 163 735
rect 159 729 163 730
rect 263 734 267 735
rect 263 729 267 730
rect 311 734 315 735
rect 311 729 315 730
rect 431 734 435 735
rect 431 729 435 730
rect 471 734 475 735
rect 471 729 475 730
rect 623 734 627 735
rect 623 729 627 730
rect 775 734 779 735
rect 775 729 779 730
rect 823 734 827 735
rect 823 729 827 730
rect 935 734 939 735
rect 935 729 939 730
rect 1015 734 1019 735
rect 1015 729 1019 730
rect 1095 734 1099 735
rect 1095 729 1099 730
rect 1207 734 1211 735
rect 1207 729 1211 730
rect 1255 734 1259 735
rect 1255 729 1259 730
rect 1391 734 1395 735
rect 1391 729 1395 730
rect 1415 734 1419 735
rect 1415 729 1419 730
rect 1567 734 1571 735
rect 1567 729 1571 730
rect 1583 734 1587 735
rect 1583 729 1587 730
rect 1743 734 1747 735
rect 1743 729 1747 730
rect 1751 734 1755 735
rect 1751 729 1755 730
rect 1903 734 1907 735
rect 1903 729 1907 730
rect 2007 734 2011 735
rect 2007 729 2011 730
rect 2047 734 2051 735
rect 2047 729 2051 730
rect 2071 734 2075 735
rect 2071 729 2075 730
rect 2255 734 2259 735
rect 2255 729 2259 730
rect 2311 734 2315 735
rect 2311 729 2315 730
rect 2455 734 2459 735
rect 2455 729 2459 730
rect 2495 734 2499 735
rect 2495 729 2499 730
rect 2655 734 2659 735
rect 2655 729 2659 730
rect 2687 734 2691 735
rect 2687 729 2691 730
rect 2855 734 2859 735
rect 2855 729 2859 730
rect 2879 734 2883 735
rect 2879 729 2883 730
rect 3047 734 3051 735
rect 3047 729 3051 730
rect 3079 734 3083 735
rect 3079 729 3083 730
rect 3239 734 3243 735
rect 3239 729 3243 730
rect 3287 734 3291 735
rect 3287 729 3291 730
rect 3439 734 3443 735
rect 3439 729 3443 730
rect 3503 734 3507 735
rect 3503 729 3507 730
rect 3639 734 3643 735
rect 3639 729 3643 730
rect 3719 734 3723 735
rect 3719 729 3723 730
rect 3839 734 3843 735
rect 3839 729 3843 730
rect 3943 734 3947 735
rect 3943 729 3947 730
rect 112 702 114 729
rect 136 705 138 729
rect 264 705 266 729
rect 432 705 434 729
rect 624 705 626 729
rect 824 705 826 729
rect 1016 705 1018 729
rect 1208 705 1210 729
rect 1392 705 1394 729
rect 1568 705 1570 729
rect 1744 705 1746 729
rect 1904 705 1906 729
rect 134 704 140 705
rect 110 701 116 702
rect 110 697 111 701
rect 115 697 116 701
rect 134 700 135 704
rect 139 700 140 704
rect 134 699 140 700
rect 262 704 268 705
rect 262 700 263 704
rect 267 700 268 704
rect 262 699 268 700
rect 430 704 436 705
rect 430 700 431 704
rect 435 700 436 704
rect 430 699 436 700
rect 622 704 628 705
rect 622 700 623 704
rect 627 700 628 704
rect 622 699 628 700
rect 822 704 828 705
rect 822 700 823 704
rect 827 700 828 704
rect 822 699 828 700
rect 1014 704 1020 705
rect 1014 700 1015 704
rect 1019 700 1020 704
rect 1014 699 1020 700
rect 1206 704 1212 705
rect 1206 700 1207 704
rect 1211 700 1212 704
rect 1206 699 1212 700
rect 1390 704 1396 705
rect 1390 700 1391 704
rect 1395 700 1396 704
rect 1390 699 1396 700
rect 1566 704 1572 705
rect 1566 700 1567 704
rect 1571 700 1572 704
rect 1566 699 1572 700
rect 1742 704 1748 705
rect 1742 700 1743 704
rect 1747 700 1748 704
rect 1742 699 1748 700
rect 1902 704 1908 705
rect 1902 700 1903 704
rect 1907 700 1908 704
rect 2008 702 2010 729
rect 2048 702 2050 729
rect 2072 705 2074 729
rect 2256 705 2258 729
rect 2456 705 2458 729
rect 2656 705 2658 729
rect 2856 705 2858 729
rect 3048 705 3050 729
rect 3240 705 3242 729
rect 3440 705 3442 729
rect 3640 705 3642 729
rect 3840 705 3842 729
rect 2070 704 2076 705
rect 1902 699 1908 700
rect 2006 701 2012 702
rect 110 696 116 697
rect 2006 697 2007 701
rect 2011 697 2012 701
rect 2006 696 2012 697
rect 2046 701 2052 702
rect 2046 697 2047 701
rect 2051 697 2052 701
rect 2070 700 2071 704
rect 2075 700 2076 704
rect 2070 699 2076 700
rect 2254 704 2260 705
rect 2254 700 2255 704
rect 2259 700 2260 704
rect 2254 699 2260 700
rect 2454 704 2460 705
rect 2454 700 2455 704
rect 2459 700 2460 704
rect 2454 699 2460 700
rect 2654 704 2660 705
rect 2654 700 2655 704
rect 2659 700 2660 704
rect 2654 699 2660 700
rect 2854 704 2860 705
rect 2854 700 2855 704
rect 2859 700 2860 704
rect 2854 699 2860 700
rect 3046 704 3052 705
rect 3046 700 3047 704
rect 3051 700 3052 704
rect 3046 699 3052 700
rect 3238 704 3244 705
rect 3238 700 3239 704
rect 3243 700 3244 704
rect 3238 699 3244 700
rect 3438 704 3444 705
rect 3438 700 3439 704
rect 3443 700 3444 704
rect 3438 699 3444 700
rect 3638 704 3644 705
rect 3638 700 3639 704
rect 3643 700 3644 704
rect 3638 699 3644 700
rect 3838 704 3844 705
rect 3838 700 3839 704
rect 3843 700 3844 704
rect 3944 702 3946 729
rect 3838 699 3844 700
rect 3942 701 3948 702
rect 2046 696 2052 697
rect 3942 697 3943 701
rect 3947 697 3948 701
rect 3942 696 3948 697
rect 134 685 140 686
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 134 681 135 685
rect 139 681 140 685
rect 134 680 140 681
rect 262 685 268 686
rect 262 681 263 685
rect 267 681 268 685
rect 262 680 268 681
rect 430 685 436 686
rect 430 681 431 685
rect 435 681 436 685
rect 430 680 436 681
rect 622 685 628 686
rect 622 681 623 685
rect 627 681 628 685
rect 622 680 628 681
rect 822 685 828 686
rect 822 681 823 685
rect 827 681 828 685
rect 822 680 828 681
rect 1014 685 1020 686
rect 1014 681 1015 685
rect 1019 681 1020 685
rect 1014 680 1020 681
rect 1206 685 1212 686
rect 1206 681 1207 685
rect 1211 681 1212 685
rect 1206 680 1212 681
rect 1390 685 1396 686
rect 1390 681 1391 685
rect 1395 681 1396 685
rect 1390 680 1396 681
rect 1566 685 1572 686
rect 1566 681 1567 685
rect 1571 681 1572 685
rect 1566 680 1572 681
rect 1742 685 1748 686
rect 1742 681 1743 685
rect 1747 681 1748 685
rect 1742 680 1748 681
rect 1902 685 1908 686
rect 2070 685 2076 686
rect 1902 681 1903 685
rect 1907 681 1908 685
rect 1902 680 1908 681
rect 2006 684 2012 685
rect 2006 680 2007 684
rect 2011 680 2012 684
rect 110 679 116 680
rect 112 659 114 679
rect 136 659 138 680
rect 264 659 266 680
rect 432 659 434 680
rect 624 659 626 680
rect 824 659 826 680
rect 1016 659 1018 680
rect 1208 659 1210 680
rect 1392 659 1394 680
rect 1568 659 1570 680
rect 1744 659 1746 680
rect 1904 659 1906 680
rect 2006 679 2012 680
rect 2046 684 2052 685
rect 2046 680 2047 684
rect 2051 680 2052 684
rect 2070 681 2071 685
rect 2075 681 2076 685
rect 2070 680 2076 681
rect 2254 685 2260 686
rect 2254 681 2255 685
rect 2259 681 2260 685
rect 2254 680 2260 681
rect 2454 685 2460 686
rect 2454 681 2455 685
rect 2459 681 2460 685
rect 2454 680 2460 681
rect 2654 685 2660 686
rect 2654 681 2655 685
rect 2659 681 2660 685
rect 2654 680 2660 681
rect 2854 685 2860 686
rect 2854 681 2855 685
rect 2859 681 2860 685
rect 2854 680 2860 681
rect 3046 685 3052 686
rect 3046 681 3047 685
rect 3051 681 3052 685
rect 3046 680 3052 681
rect 3238 685 3244 686
rect 3238 681 3239 685
rect 3243 681 3244 685
rect 3238 680 3244 681
rect 3438 685 3444 686
rect 3438 681 3439 685
rect 3443 681 3444 685
rect 3438 680 3444 681
rect 3638 685 3644 686
rect 3638 681 3639 685
rect 3643 681 3644 685
rect 3638 680 3644 681
rect 3838 685 3844 686
rect 3838 681 3839 685
rect 3843 681 3844 685
rect 3838 680 3844 681
rect 3942 684 3948 685
rect 3942 680 3943 684
rect 3947 680 3948 684
rect 2046 679 2052 680
rect 2008 659 2010 679
rect 2048 659 2050 679
rect 2072 659 2074 680
rect 2256 659 2258 680
rect 2456 659 2458 680
rect 2656 659 2658 680
rect 2856 659 2858 680
rect 3048 659 3050 680
rect 3240 659 3242 680
rect 3440 659 3442 680
rect 3640 659 3642 680
rect 3840 659 3842 680
rect 3942 679 3948 680
rect 3944 659 3946 679
rect 111 658 115 659
rect 111 653 115 654
rect 135 658 139 659
rect 135 653 139 654
rect 247 658 251 659
rect 247 653 251 654
rect 263 658 267 659
rect 263 653 267 654
rect 383 658 387 659
rect 383 653 387 654
rect 431 658 435 659
rect 431 653 435 654
rect 527 658 531 659
rect 527 653 531 654
rect 623 658 627 659
rect 623 653 627 654
rect 687 658 691 659
rect 687 653 691 654
rect 823 658 827 659
rect 823 653 827 654
rect 871 658 875 659
rect 871 653 875 654
rect 1015 658 1019 659
rect 1015 653 1019 654
rect 1079 658 1083 659
rect 1079 653 1083 654
rect 1207 658 1211 659
rect 1207 653 1211 654
rect 1303 658 1307 659
rect 1303 653 1307 654
rect 1391 658 1395 659
rect 1391 653 1395 654
rect 1543 658 1547 659
rect 1543 653 1547 654
rect 1567 658 1571 659
rect 1567 653 1571 654
rect 1743 658 1747 659
rect 1743 653 1747 654
rect 1783 658 1787 659
rect 1783 653 1787 654
rect 1903 658 1907 659
rect 1903 653 1907 654
rect 2007 658 2011 659
rect 2007 653 2011 654
rect 2047 658 2051 659
rect 2047 653 2051 654
rect 2071 658 2075 659
rect 2071 653 2075 654
rect 2231 658 2235 659
rect 2231 653 2235 654
rect 2255 658 2259 659
rect 2255 653 2259 654
rect 2431 658 2435 659
rect 2431 653 2435 654
rect 2455 658 2459 659
rect 2455 653 2459 654
rect 2631 658 2635 659
rect 2631 653 2635 654
rect 2655 658 2659 659
rect 2655 653 2659 654
rect 2831 658 2835 659
rect 2831 653 2835 654
rect 2855 658 2859 659
rect 2855 653 2859 654
rect 3023 658 3027 659
rect 3023 653 3027 654
rect 3047 658 3051 659
rect 3047 653 3051 654
rect 3207 658 3211 659
rect 3207 653 3211 654
rect 3239 658 3243 659
rect 3239 653 3243 654
rect 3375 658 3379 659
rect 3375 653 3379 654
rect 3439 658 3443 659
rect 3439 653 3443 654
rect 3535 658 3539 659
rect 3535 653 3539 654
rect 3639 658 3643 659
rect 3639 653 3643 654
rect 3695 658 3699 659
rect 3695 653 3699 654
rect 3839 658 3843 659
rect 3839 653 3843 654
rect 3943 658 3947 659
rect 3943 653 3947 654
rect 112 633 114 653
rect 110 632 116 633
rect 136 632 138 653
rect 248 632 250 653
rect 384 632 386 653
rect 528 632 530 653
rect 688 632 690 653
rect 872 632 874 653
rect 1080 632 1082 653
rect 1304 632 1306 653
rect 1544 632 1546 653
rect 1784 632 1786 653
rect 2008 633 2010 653
rect 2048 633 2050 653
rect 2006 632 2012 633
rect 110 628 111 632
rect 115 628 116 632
rect 110 627 116 628
rect 134 631 140 632
rect 134 627 135 631
rect 139 627 140 631
rect 134 626 140 627
rect 246 631 252 632
rect 246 627 247 631
rect 251 627 252 631
rect 246 626 252 627
rect 382 631 388 632
rect 382 627 383 631
rect 387 627 388 631
rect 382 626 388 627
rect 526 631 532 632
rect 526 627 527 631
rect 531 627 532 631
rect 526 626 532 627
rect 686 631 692 632
rect 686 627 687 631
rect 691 627 692 631
rect 686 626 692 627
rect 870 631 876 632
rect 870 627 871 631
rect 875 627 876 631
rect 870 626 876 627
rect 1078 631 1084 632
rect 1078 627 1079 631
rect 1083 627 1084 631
rect 1078 626 1084 627
rect 1302 631 1308 632
rect 1302 627 1303 631
rect 1307 627 1308 631
rect 1302 626 1308 627
rect 1542 631 1548 632
rect 1542 627 1543 631
rect 1547 627 1548 631
rect 1542 626 1548 627
rect 1782 631 1788 632
rect 1782 627 1783 631
rect 1787 627 1788 631
rect 2006 628 2007 632
rect 2011 628 2012 632
rect 2006 627 2012 628
rect 2046 632 2052 633
rect 2072 632 2074 653
rect 2232 632 2234 653
rect 2432 632 2434 653
rect 2632 632 2634 653
rect 2832 632 2834 653
rect 3024 632 3026 653
rect 3208 632 3210 653
rect 3376 632 3378 653
rect 3536 632 3538 653
rect 3696 632 3698 653
rect 3840 632 3842 653
rect 3944 633 3946 653
rect 3942 632 3948 633
rect 2046 628 2047 632
rect 2051 628 2052 632
rect 2046 627 2052 628
rect 2070 631 2076 632
rect 2070 627 2071 631
rect 2075 627 2076 631
rect 1782 626 1788 627
rect 2070 626 2076 627
rect 2230 631 2236 632
rect 2230 627 2231 631
rect 2235 627 2236 631
rect 2230 626 2236 627
rect 2430 631 2436 632
rect 2430 627 2431 631
rect 2435 627 2436 631
rect 2430 626 2436 627
rect 2630 631 2636 632
rect 2630 627 2631 631
rect 2635 627 2636 631
rect 2630 626 2636 627
rect 2830 631 2836 632
rect 2830 627 2831 631
rect 2835 627 2836 631
rect 2830 626 2836 627
rect 3022 631 3028 632
rect 3022 627 3023 631
rect 3027 627 3028 631
rect 3022 626 3028 627
rect 3206 631 3212 632
rect 3206 627 3207 631
rect 3211 627 3212 631
rect 3206 626 3212 627
rect 3374 631 3380 632
rect 3374 627 3375 631
rect 3379 627 3380 631
rect 3374 626 3380 627
rect 3534 631 3540 632
rect 3534 627 3535 631
rect 3539 627 3540 631
rect 3534 626 3540 627
rect 3694 631 3700 632
rect 3694 627 3695 631
rect 3699 627 3700 631
rect 3694 626 3700 627
rect 3838 631 3844 632
rect 3838 627 3839 631
rect 3843 627 3844 631
rect 3942 628 3943 632
rect 3947 628 3948 632
rect 3942 627 3948 628
rect 3838 626 3844 627
rect 110 615 116 616
rect 110 611 111 615
rect 115 611 116 615
rect 2006 615 2012 616
rect 110 610 116 611
rect 134 612 140 613
rect 112 579 114 610
rect 134 608 135 612
rect 139 608 140 612
rect 134 607 140 608
rect 246 612 252 613
rect 246 608 247 612
rect 251 608 252 612
rect 246 607 252 608
rect 382 612 388 613
rect 382 608 383 612
rect 387 608 388 612
rect 382 607 388 608
rect 526 612 532 613
rect 526 608 527 612
rect 531 608 532 612
rect 526 607 532 608
rect 686 612 692 613
rect 686 608 687 612
rect 691 608 692 612
rect 686 607 692 608
rect 870 612 876 613
rect 870 608 871 612
rect 875 608 876 612
rect 870 607 876 608
rect 1078 612 1084 613
rect 1078 608 1079 612
rect 1083 608 1084 612
rect 1078 607 1084 608
rect 1302 612 1308 613
rect 1302 608 1303 612
rect 1307 608 1308 612
rect 1302 607 1308 608
rect 1542 612 1548 613
rect 1542 608 1543 612
rect 1547 608 1548 612
rect 1542 607 1548 608
rect 1782 612 1788 613
rect 1782 608 1783 612
rect 1787 608 1788 612
rect 2006 611 2007 615
rect 2011 611 2012 615
rect 2006 610 2012 611
rect 2046 615 2052 616
rect 2046 611 2047 615
rect 2051 611 2052 615
rect 3942 615 3948 616
rect 2046 610 2052 611
rect 2070 612 2076 613
rect 1782 607 1788 608
rect 136 579 138 607
rect 248 579 250 607
rect 384 579 386 607
rect 528 579 530 607
rect 688 579 690 607
rect 872 579 874 607
rect 1080 579 1082 607
rect 1304 579 1306 607
rect 1544 579 1546 607
rect 1784 579 1786 607
rect 2008 579 2010 610
rect 2048 579 2050 610
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 2230 612 2236 613
rect 2230 608 2231 612
rect 2235 608 2236 612
rect 2230 607 2236 608
rect 2430 612 2436 613
rect 2430 608 2431 612
rect 2435 608 2436 612
rect 2430 607 2436 608
rect 2630 612 2636 613
rect 2630 608 2631 612
rect 2635 608 2636 612
rect 2630 607 2636 608
rect 2830 612 2836 613
rect 2830 608 2831 612
rect 2835 608 2836 612
rect 2830 607 2836 608
rect 3022 612 3028 613
rect 3022 608 3023 612
rect 3027 608 3028 612
rect 3022 607 3028 608
rect 3206 612 3212 613
rect 3206 608 3207 612
rect 3211 608 3212 612
rect 3206 607 3212 608
rect 3374 612 3380 613
rect 3374 608 3375 612
rect 3379 608 3380 612
rect 3374 607 3380 608
rect 3534 612 3540 613
rect 3534 608 3535 612
rect 3539 608 3540 612
rect 3534 607 3540 608
rect 3694 612 3700 613
rect 3694 608 3695 612
rect 3699 608 3700 612
rect 3694 607 3700 608
rect 3838 612 3844 613
rect 3838 608 3839 612
rect 3843 608 3844 612
rect 3942 611 3943 615
rect 3947 611 3948 615
rect 3942 610 3948 611
rect 3838 607 3844 608
rect 2072 579 2074 607
rect 2232 579 2234 607
rect 2432 579 2434 607
rect 2632 579 2634 607
rect 2832 579 2834 607
rect 3024 579 3026 607
rect 3208 579 3210 607
rect 3376 579 3378 607
rect 3536 579 3538 607
rect 3696 579 3698 607
rect 3840 579 3842 607
rect 3944 579 3946 610
rect 111 578 115 579
rect 111 573 115 574
rect 135 578 139 579
rect 135 573 139 574
rect 247 578 251 579
rect 247 573 251 574
rect 295 578 299 579
rect 295 573 299 574
rect 383 578 387 579
rect 383 573 387 574
rect 479 578 483 579
rect 479 573 483 574
rect 527 578 531 579
rect 527 573 531 574
rect 663 578 667 579
rect 663 573 667 574
rect 687 578 691 579
rect 687 573 691 574
rect 847 578 851 579
rect 847 573 851 574
rect 871 578 875 579
rect 871 573 875 574
rect 1031 578 1035 579
rect 1031 573 1035 574
rect 1079 578 1083 579
rect 1079 573 1083 574
rect 1215 578 1219 579
rect 1215 573 1219 574
rect 1303 578 1307 579
rect 1303 573 1307 574
rect 1399 578 1403 579
rect 1399 573 1403 574
rect 1543 578 1547 579
rect 1543 573 1547 574
rect 1591 578 1595 579
rect 1591 573 1595 574
rect 1783 578 1787 579
rect 1783 573 1787 574
rect 2007 578 2011 579
rect 2007 573 2011 574
rect 2047 578 2051 579
rect 2047 573 2051 574
rect 2071 578 2075 579
rect 2071 573 2075 574
rect 2215 578 2219 579
rect 2215 573 2219 574
rect 2231 578 2235 579
rect 2231 573 2235 574
rect 2399 578 2403 579
rect 2399 573 2403 574
rect 2431 578 2435 579
rect 2431 573 2435 574
rect 2583 578 2587 579
rect 2583 573 2587 574
rect 2631 578 2635 579
rect 2631 573 2635 574
rect 2775 578 2779 579
rect 2775 573 2779 574
rect 2831 578 2835 579
rect 2831 573 2835 574
rect 2959 578 2963 579
rect 2959 573 2963 574
rect 3023 578 3027 579
rect 3023 573 3027 574
rect 3143 578 3147 579
rect 3143 573 3147 574
rect 3207 578 3211 579
rect 3207 573 3211 574
rect 3319 578 3323 579
rect 3319 573 3323 574
rect 3375 578 3379 579
rect 3375 573 3379 574
rect 3495 578 3499 579
rect 3495 573 3499 574
rect 3535 578 3539 579
rect 3535 573 3539 574
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3695 578 3699 579
rect 3695 573 3699 574
rect 3839 578 3843 579
rect 3839 573 3843 574
rect 3943 578 3947 579
rect 3943 573 3947 574
rect 112 546 114 573
rect 136 549 138 573
rect 296 549 298 573
rect 480 549 482 573
rect 664 549 666 573
rect 848 549 850 573
rect 1032 549 1034 573
rect 1216 549 1218 573
rect 1400 549 1402 573
rect 1592 549 1594 573
rect 1784 549 1786 573
rect 134 548 140 549
rect 110 545 116 546
rect 110 541 111 545
rect 115 541 116 545
rect 134 544 135 548
rect 139 544 140 548
rect 134 543 140 544
rect 294 548 300 549
rect 294 544 295 548
rect 299 544 300 548
rect 294 543 300 544
rect 478 548 484 549
rect 478 544 479 548
rect 483 544 484 548
rect 478 543 484 544
rect 662 548 668 549
rect 662 544 663 548
rect 667 544 668 548
rect 662 543 668 544
rect 846 548 852 549
rect 846 544 847 548
rect 851 544 852 548
rect 846 543 852 544
rect 1030 548 1036 549
rect 1030 544 1031 548
rect 1035 544 1036 548
rect 1030 543 1036 544
rect 1214 548 1220 549
rect 1214 544 1215 548
rect 1219 544 1220 548
rect 1214 543 1220 544
rect 1398 548 1404 549
rect 1398 544 1399 548
rect 1403 544 1404 548
rect 1398 543 1404 544
rect 1590 548 1596 549
rect 1590 544 1591 548
rect 1595 544 1596 548
rect 1590 543 1596 544
rect 1782 548 1788 549
rect 1782 544 1783 548
rect 1787 544 1788 548
rect 2008 546 2010 573
rect 2048 546 2050 573
rect 2072 549 2074 573
rect 2216 549 2218 573
rect 2400 549 2402 573
rect 2584 549 2586 573
rect 2776 549 2778 573
rect 2960 549 2962 573
rect 3144 549 3146 573
rect 3320 549 3322 573
rect 3496 549 3498 573
rect 3680 549 3682 573
rect 3840 549 3842 573
rect 2070 548 2076 549
rect 1782 543 1788 544
rect 2006 545 2012 546
rect 110 540 116 541
rect 2006 541 2007 545
rect 2011 541 2012 545
rect 2006 540 2012 541
rect 2046 545 2052 546
rect 2046 541 2047 545
rect 2051 541 2052 545
rect 2070 544 2071 548
rect 2075 544 2076 548
rect 2070 543 2076 544
rect 2214 548 2220 549
rect 2214 544 2215 548
rect 2219 544 2220 548
rect 2214 543 2220 544
rect 2398 548 2404 549
rect 2398 544 2399 548
rect 2403 544 2404 548
rect 2398 543 2404 544
rect 2582 548 2588 549
rect 2582 544 2583 548
rect 2587 544 2588 548
rect 2582 543 2588 544
rect 2774 548 2780 549
rect 2774 544 2775 548
rect 2779 544 2780 548
rect 2774 543 2780 544
rect 2958 548 2964 549
rect 2958 544 2959 548
rect 2963 544 2964 548
rect 2958 543 2964 544
rect 3142 548 3148 549
rect 3142 544 3143 548
rect 3147 544 3148 548
rect 3142 543 3148 544
rect 3318 548 3324 549
rect 3318 544 3319 548
rect 3323 544 3324 548
rect 3318 543 3324 544
rect 3494 548 3500 549
rect 3494 544 3495 548
rect 3499 544 3500 548
rect 3494 543 3500 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3678 543 3684 544
rect 3838 548 3844 549
rect 3838 544 3839 548
rect 3843 544 3844 548
rect 3944 546 3946 573
rect 3838 543 3844 544
rect 3942 545 3948 546
rect 2046 540 2052 541
rect 3942 541 3943 545
rect 3947 541 3948 545
rect 3942 540 3948 541
rect 134 529 140 530
rect 110 528 116 529
rect 110 524 111 528
rect 115 524 116 528
rect 134 525 135 529
rect 139 525 140 529
rect 134 524 140 525
rect 294 529 300 530
rect 294 525 295 529
rect 299 525 300 529
rect 294 524 300 525
rect 478 529 484 530
rect 478 525 479 529
rect 483 525 484 529
rect 478 524 484 525
rect 662 529 668 530
rect 662 525 663 529
rect 667 525 668 529
rect 662 524 668 525
rect 846 529 852 530
rect 846 525 847 529
rect 851 525 852 529
rect 846 524 852 525
rect 1030 529 1036 530
rect 1030 525 1031 529
rect 1035 525 1036 529
rect 1030 524 1036 525
rect 1214 529 1220 530
rect 1214 525 1215 529
rect 1219 525 1220 529
rect 1214 524 1220 525
rect 1398 529 1404 530
rect 1398 525 1399 529
rect 1403 525 1404 529
rect 1398 524 1404 525
rect 1590 529 1596 530
rect 1590 525 1591 529
rect 1595 525 1596 529
rect 1590 524 1596 525
rect 1782 529 1788 530
rect 2070 529 2076 530
rect 1782 525 1783 529
rect 1787 525 1788 529
rect 1782 524 1788 525
rect 2006 528 2012 529
rect 2006 524 2007 528
rect 2011 524 2012 528
rect 110 523 116 524
rect 112 503 114 523
rect 136 503 138 524
rect 296 503 298 524
rect 480 503 482 524
rect 664 503 666 524
rect 848 503 850 524
rect 1032 503 1034 524
rect 1216 503 1218 524
rect 1400 503 1402 524
rect 1592 503 1594 524
rect 1784 503 1786 524
rect 2006 523 2012 524
rect 2046 528 2052 529
rect 2046 524 2047 528
rect 2051 524 2052 528
rect 2070 525 2071 529
rect 2075 525 2076 529
rect 2070 524 2076 525
rect 2214 529 2220 530
rect 2214 525 2215 529
rect 2219 525 2220 529
rect 2214 524 2220 525
rect 2398 529 2404 530
rect 2398 525 2399 529
rect 2403 525 2404 529
rect 2398 524 2404 525
rect 2582 529 2588 530
rect 2582 525 2583 529
rect 2587 525 2588 529
rect 2582 524 2588 525
rect 2774 529 2780 530
rect 2774 525 2775 529
rect 2779 525 2780 529
rect 2774 524 2780 525
rect 2958 529 2964 530
rect 2958 525 2959 529
rect 2963 525 2964 529
rect 2958 524 2964 525
rect 3142 529 3148 530
rect 3142 525 3143 529
rect 3147 525 3148 529
rect 3142 524 3148 525
rect 3318 529 3324 530
rect 3318 525 3319 529
rect 3323 525 3324 529
rect 3318 524 3324 525
rect 3494 529 3500 530
rect 3494 525 3495 529
rect 3499 525 3500 529
rect 3494 524 3500 525
rect 3678 529 3684 530
rect 3678 525 3679 529
rect 3683 525 3684 529
rect 3678 524 3684 525
rect 3838 529 3844 530
rect 3838 525 3839 529
rect 3843 525 3844 529
rect 3838 524 3844 525
rect 3942 528 3948 529
rect 3942 524 3943 528
rect 3947 524 3948 528
rect 2046 523 2052 524
rect 2008 503 2010 523
rect 111 502 115 503
rect 111 497 115 498
rect 135 502 139 503
rect 135 497 139 498
rect 287 502 291 503
rect 287 497 291 498
rect 295 502 299 503
rect 295 497 299 498
rect 455 502 459 503
rect 455 497 459 498
rect 479 502 483 503
rect 479 497 483 498
rect 615 502 619 503
rect 615 497 619 498
rect 663 502 667 503
rect 663 497 667 498
rect 767 502 771 503
rect 767 497 771 498
rect 847 502 851 503
rect 847 497 851 498
rect 903 502 907 503
rect 903 497 907 498
rect 1031 502 1035 503
rect 1031 497 1035 498
rect 1159 502 1163 503
rect 1159 497 1163 498
rect 1215 502 1219 503
rect 1215 497 1219 498
rect 1287 502 1291 503
rect 1287 497 1291 498
rect 1399 502 1403 503
rect 1399 497 1403 498
rect 1415 502 1419 503
rect 1415 497 1419 498
rect 1591 502 1595 503
rect 1591 497 1595 498
rect 1783 502 1787 503
rect 1783 497 1787 498
rect 2007 502 2011 503
rect 2048 499 2050 523
rect 2072 499 2074 524
rect 2216 499 2218 524
rect 2400 499 2402 524
rect 2584 499 2586 524
rect 2776 499 2778 524
rect 2960 499 2962 524
rect 3144 499 3146 524
rect 3320 499 3322 524
rect 3496 499 3498 524
rect 3680 499 3682 524
rect 3840 499 3842 524
rect 3942 523 3948 524
rect 3944 499 3946 523
rect 2007 497 2011 498
rect 2047 498 2051 499
rect 112 477 114 497
rect 110 476 116 477
rect 136 476 138 497
rect 288 476 290 497
rect 456 476 458 497
rect 616 476 618 497
rect 768 476 770 497
rect 904 476 906 497
rect 1032 476 1034 497
rect 1160 476 1162 497
rect 1288 476 1290 497
rect 1416 476 1418 497
rect 2008 477 2010 497
rect 2047 493 2051 494
rect 2071 498 2075 499
rect 2071 493 2075 494
rect 2215 498 2219 499
rect 2215 493 2219 494
rect 2223 498 2227 499
rect 2223 493 2227 494
rect 2391 498 2395 499
rect 2391 493 2395 494
rect 2399 498 2403 499
rect 2399 493 2403 494
rect 2559 498 2563 499
rect 2559 493 2563 494
rect 2583 498 2587 499
rect 2583 493 2587 494
rect 2727 498 2731 499
rect 2727 493 2731 494
rect 2775 498 2779 499
rect 2775 493 2779 494
rect 2895 498 2899 499
rect 2895 493 2899 494
rect 2959 498 2963 499
rect 2959 493 2963 494
rect 3063 498 3067 499
rect 3063 493 3067 494
rect 3143 498 3147 499
rect 3143 493 3147 494
rect 3223 498 3227 499
rect 3223 493 3227 494
rect 3319 498 3323 499
rect 3319 493 3323 494
rect 3383 498 3387 499
rect 3383 493 3387 494
rect 3495 498 3499 499
rect 3495 493 3499 494
rect 3543 498 3547 499
rect 3543 493 3547 494
rect 3679 498 3683 499
rect 3679 493 3683 494
rect 3703 498 3707 499
rect 3703 493 3707 494
rect 3839 498 3843 499
rect 3839 493 3843 494
rect 3943 498 3947 499
rect 3943 493 3947 494
rect 2006 476 2012 477
rect 110 472 111 476
rect 115 472 116 476
rect 110 471 116 472
rect 134 475 140 476
rect 134 471 135 475
rect 139 471 140 475
rect 134 470 140 471
rect 286 475 292 476
rect 286 471 287 475
rect 291 471 292 475
rect 286 470 292 471
rect 454 475 460 476
rect 454 471 455 475
rect 459 471 460 475
rect 454 470 460 471
rect 614 475 620 476
rect 614 471 615 475
rect 619 471 620 475
rect 614 470 620 471
rect 766 475 772 476
rect 766 471 767 475
rect 771 471 772 475
rect 766 470 772 471
rect 902 475 908 476
rect 902 471 903 475
rect 907 471 908 475
rect 902 470 908 471
rect 1030 475 1036 476
rect 1030 471 1031 475
rect 1035 471 1036 475
rect 1030 470 1036 471
rect 1158 475 1164 476
rect 1158 471 1159 475
rect 1163 471 1164 475
rect 1158 470 1164 471
rect 1286 475 1292 476
rect 1286 471 1287 475
rect 1291 471 1292 475
rect 1286 470 1292 471
rect 1414 475 1420 476
rect 1414 471 1415 475
rect 1419 471 1420 475
rect 2006 472 2007 476
rect 2011 472 2012 476
rect 2048 473 2050 493
rect 2006 471 2012 472
rect 2046 472 2052 473
rect 2072 472 2074 493
rect 2224 472 2226 493
rect 2392 472 2394 493
rect 2560 472 2562 493
rect 2728 472 2730 493
rect 2896 472 2898 493
rect 3064 472 3066 493
rect 3224 472 3226 493
rect 3384 472 3386 493
rect 3544 472 3546 493
rect 3704 472 3706 493
rect 3840 472 3842 493
rect 3944 473 3946 493
rect 3942 472 3948 473
rect 1414 470 1420 471
rect 2046 468 2047 472
rect 2051 468 2052 472
rect 2046 467 2052 468
rect 2070 471 2076 472
rect 2070 467 2071 471
rect 2075 467 2076 471
rect 2070 466 2076 467
rect 2222 471 2228 472
rect 2222 467 2223 471
rect 2227 467 2228 471
rect 2222 466 2228 467
rect 2390 471 2396 472
rect 2390 467 2391 471
rect 2395 467 2396 471
rect 2390 466 2396 467
rect 2558 471 2564 472
rect 2558 467 2559 471
rect 2563 467 2564 471
rect 2558 466 2564 467
rect 2726 471 2732 472
rect 2726 467 2727 471
rect 2731 467 2732 471
rect 2726 466 2732 467
rect 2894 471 2900 472
rect 2894 467 2895 471
rect 2899 467 2900 471
rect 2894 466 2900 467
rect 3062 471 3068 472
rect 3062 467 3063 471
rect 3067 467 3068 471
rect 3062 466 3068 467
rect 3222 471 3228 472
rect 3222 467 3223 471
rect 3227 467 3228 471
rect 3222 466 3228 467
rect 3382 471 3388 472
rect 3382 467 3383 471
rect 3387 467 3388 471
rect 3382 466 3388 467
rect 3542 471 3548 472
rect 3542 467 3543 471
rect 3547 467 3548 471
rect 3542 466 3548 467
rect 3702 471 3708 472
rect 3702 467 3703 471
rect 3707 467 3708 471
rect 3702 466 3708 467
rect 3838 471 3844 472
rect 3838 467 3839 471
rect 3843 467 3844 471
rect 3942 468 3943 472
rect 3947 468 3948 472
rect 3942 467 3948 468
rect 3838 466 3844 467
rect 110 459 116 460
rect 110 455 111 459
rect 115 455 116 459
rect 2006 459 2012 460
rect 110 454 116 455
rect 134 456 140 457
rect 112 427 114 454
rect 134 452 135 456
rect 139 452 140 456
rect 134 451 140 452
rect 286 456 292 457
rect 286 452 287 456
rect 291 452 292 456
rect 286 451 292 452
rect 454 456 460 457
rect 454 452 455 456
rect 459 452 460 456
rect 454 451 460 452
rect 614 456 620 457
rect 614 452 615 456
rect 619 452 620 456
rect 614 451 620 452
rect 766 456 772 457
rect 766 452 767 456
rect 771 452 772 456
rect 766 451 772 452
rect 902 456 908 457
rect 902 452 903 456
rect 907 452 908 456
rect 902 451 908 452
rect 1030 456 1036 457
rect 1030 452 1031 456
rect 1035 452 1036 456
rect 1030 451 1036 452
rect 1158 456 1164 457
rect 1158 452 1159 456
rect 1163 452 1164 456
rect 1158 451 1164 452
rect 1286 456 1292 457
rect 1286 452 1287 456
rect 1291 452 1292 456
rect 1286 451 1292 452
rect 1414 456 1420 457
rect 1414 452 1415 456
rect 1419 452 1420 456
rect 2006 455 2007 459
rect 2011 455 2012 459
rect 2006 454 2012 455
rect 2046 455 2052 456
rect 1414 451 1420 452
rect 136 427 138 451
rect 288 427 290 451
rect 456 427 458 451
rect 616 427 618 451
rect 768 427 770 451
rect 904 427 906 451
rect 1032 427 1034 451
rect 1160 427 1162 451
rect 1288 427 1290 451
rect 1416 427 1418 451
rect 2008 427 2010 454
rect 2046 451 2047 455
rect 2051 451 2052 455
rect 3942 455 3948 456
rect 2046 450 2052 451
rect 2070 452 2076 453
rect 111 426 115 427
rect 111 421 115 422
rect 135 426 139 427
rect 135 421 139 422
rect 287 426 291 427
rect 287 421 291 422
rect 447 426 451 427
rect 447 421 451 422
rect 455 426 459 427
rect 455 421 459 422
rect 599 426 603 427
rect 599 421 603 422
rect 615 426 619 427
rect 615 421 619 422
rect 751 426 755 427
rect 751 421 755 422
rect 767 426 771 427
rect 767 421 771 422
rect 903 426 907 427
rect 903 421 907 422
rect 1031 426 1035 427
rect 1031 421 1035 422
rect 1079 426 1083 427
rect 1079 421 1083 422
rect 1159 426 1163 427
rect 1159 421 1163 422
rect 1271 426 1275 427
rect 1271 421 1275 422
rect 1287 426 1291 427
rect 1287 421 1291 422
rect 1415 426 1419 427
rect 1415 421 1419 422
rect 1479 426 1483 427
rect 1479 421 1483 422
rect 1703 426 1707 427
rect 1703 421 1707 422
rect 1903 426 1907 427
rect 1903 421 1907 422
rect 2007 426 2011 427
rect 2048 423 2050 450
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 2222 452 2228 453
rect 2222 448 2223 452
rect 2227 448 2228 452
rect 2222 447 2228 448
rect 2390 452 2396 453
rect 2390 448 2391 452
rect 2395 448 2396 452
rect 2390 447 2396 448
rect 2558 452 2564 453
rect 2558 448 2559 452
rect 2563 448 2564 452
rect 2558 447 2564 448
rect 2726 452 2732 453
rect 2726 448 2727 452
rect 2731 448 2732 452
rect 2726 447 2732 448
rect 2894 452 2900 453
rect 2894 448 2895 452
rect 2899 448 2900 452
rect 2894 447 2900 448
rect 3062 452 3068 453
rect 3062 448 3063 452
rect 3067 448 3068 452
rect 3062 447 3068 448
rect 3222 452 3228 453
rect 3222 448 3223 452
rect 3227 448 3228 452
rect 3222 447 3228 448
rect 3382 452 3388 453
rect 3382 448 3383 452
rect 3387 448 3388 452
rect 3382 447 3388 448
rect 3542 452 3548 453
rect 3542 448 3543 452
rect 3547 448 3548 452
rect 3542 447 3548 448
rect 3702 452 3708 453
rect 3702 448 3703 452
rect 3707 448 3708 452
rect 3702 447 3708 448
rect 3838 452 3844 453
rect 3838 448 3839 452
rect 3843 448 3844 452
rect 3942 451 3943 455
rect 3947 451 3948 455
rect 3942 450 3948 451
rect 3838 447 3844 448
rect 2072 423 2074 447
rect 2224 423 2226 447
rect 2392 423 2394 447
rect 2560 423 2562 447
rect 2728 423 2730 447
rect 2896 423 2898 447
rect 3064 423 3066 447
rect 3224 423 3226 447
rect 3384 423 3386 447
rect 3544 423 3546 447
rect 3704 423 3706 447
rect 3840 423 3842 447
rect 3944 423 3946 450
rect 2007 421 2011 422
rect 2047 422 2051 423
rect 112 394 114 421
rect 136 397 138 421
rect 288 397 290 421
rect 448 397 450 421
rect 600 397 602 421
rect 752 397 754 421
rect 904 397 906 421
rect 1080 397 1082 421
rect 1272 397 1274 421
rect 1480 397 1482 421
rect 1704 397 1706 421
rect 1904 397 1906 421
rect 134 396 140 397
rect 110 393 116 394
rect 110 389 111 393
rect 115 389 116 393
rect 134 392 135 396
rect 139 392 140 396
rect 134 391 140 392
rect 286 396 292 397
rect 286 392 287 396
rect 291 392 292 396
rect 286 391 292 392
rect 446 396 452 397
rect 446 392 447 396
rect 451 392 452 396
rect 446 391 452 392
rect 598 396 604 397
rect 598 392 599 396
rect 603 392 604 396
rect 598 391 604 392
rect 750 396 756 397
rect 750 392 751 396
rect 755 392 756 396
rect 750 391 756 392
rect 902 396 908 397
rect 902 392 903 396
rect 907 392 908 396
rect 902 391 908 392
rect 1078 396 1084 397
rect 1078 392 1079 396
rect 1083 392 1084 396
rect 1078 391 1084 392
rect 1270 396 1276 397
rect 1270 392 1271 396
rect 1275 392 1276 396
rect 1270 391 1276 392
rect 1478 396 1484 397
rect 1478 392 1479 396
rect 1483 392 1484 396
rect 1478 391 1484 392
rect 1702 396 1708 397
rect 1702 392 1703 396
rect 1707 392 1708 396
rect 1702 391 1708 392
rect 1902 396 1908 397
rect 1902 392 1903 396
rect 1907 392 1908 396
rect 2008 394 2010 421
rect 2047 417 2051 418
rect 2071 422 2075 423
rect 2071 417 2075 418
rect 2223 422 2227 423
rect 2223 417 2227 418
rect 2391 422 2395 423
rect 2391 417 2395 418
rect 2463 422 2467 423
rect 2463 417 2467 418
rect 2559 422 2563 423
rect 2559 417 2563 418
rect 2655 422 2659 423
rect 2655 417 2659 418
rect 2727 422 2731 423
rect 2727 417 2731 418
rect 2751 422 2755 423
rect 2751 417 2755 418
rect 2847 422 2851 423
rect 2847 417 2851 418
rect 2895 422 2899 423
rect 2895 417 2899 418
rect 2943 422 2947 423
rect 2943 417 2947 418
rect 3039 422 3043 423
rect 3039 417 3043 418
rect 3063 422 3067 423
rect 3063 417 3067 418
rect 3135 422 3139 423
rect 3135 417 3139 418
rect 3223 422 3227 423
rect 3223 417 3227 418
rect 3231 422 3235 423
rect 3231 417 3235 418
rect 3383 422 3387 423
rect 3383 417 3387 418
rect 3543 422 3547 423
rect 3543 417 3547 418
rect 3703 422 3707 423
rect 3703 417 3707 418
rect 3839 422 3843 423
rect 3839 417 3843 418
rect 3943 422 3947 423
rect 3943 417 3947 418
rect 1902 391 1908 392
rect 2006 393 2012 394
rect 110 388 116 389
rect 2006 389 2007 393
rect 2011 389 2012 393
rect 2048 390 2050 417
rect 2464 393 2466 417
rect 2560 393 2562 417
rect 2656 393 2658 417
rect 2752 393 2754 417
rect 2848 393 2850 417
rect 2944 393 2946 417
rect 3040 393 3042 417
rect 3136 393 3138 417
rect 3232 393 3234 417
rect 2462 392 2468 393
rect 2006 388 2012 389
rect 2046 389 2052 390
rect 2046 385 2047 389
rect 2051 385 2052 389
rect 2462 388 2463 392
rect 2467 388 2468 392
rect 2462 387 2468 388
rect 2558 392 2564 393
rect 2558 388 2559 392
rect 2563 388 2564 392
rect 2558 387 2564 388
rect 2654 392 2660 393
rect 2654 388 2655 392
rect 2659 388 2660 392
rect 2654 387 2660 388
rect 2750 392 2756 393
rect 2750 388 2751 392
rect 2755 388 2756 392
rect 2750 387 2756 388
rect 2846 392 2852 393
rect 2846 388 2847 392
rect 2851 388 2852 392
rect 2846 387 2852 388
rect 2942 392 2948 393
rect 2942 388 2943 392
rect 2947 388 2948 392
rect 2942 387 2948 388
rect 3038 392 3044 393
rect 3038 388 3039 392
rect 3043 388 3044 392
rect 3038 387 3044 388
rect 3134 392 3140 393
rect 3134 388 3135 392
rect 3139 388 3140 392
rect 3134 387 3140 388
rect 3230 392 3236 393
rect 3230 388 3231 392
rect 3235 388 3236 392
rect 3944 390 3946 417
rect 3230 387 3236 388
rect 3942 389 3948 390
rect 2046 384 2052 385
rect 3942 385 3943 389
rect 3947 385 3948 389
rect 3942 384 3948 385
rect 134 377 140 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 134 373 135 377
rect 139 373 140 377
rect 134 372 140 373
rect 286 377 292 378
rect 286 373 287 377
rect 291 373 292 377
rect 286 372 292 373
rect 446 377 452 378
rect 446 373 447 377
rect 451 373 452 377
rect 446 372 452 373
rect 598 377 604 378
rect 598 373 599 377
rect 603 373 604 377
rect 598 372 604 373
rect 750 377 756 378
rect 750 373 751 377
rect 755 373 756 377
rect 750 372 756 373
rect 902 377 908 378
rect 902 373 903 377
rect 907 373 908 377
rect 902 372 908 373
rect 1078 377 1084 378
rect 1078 373 1079 377
rect 1083 373 1084 377
rect 1078 372 1084 373
rect 1270 377 1276 378
rect 1270 373 1271 377
rect 1275 373 1276 377
rect 1270 372 1276 373
rect 1478 377 1484 378
rect 1478 373 1479 377
rect 1483 373 1484 377
rect 1478 372 1484 373
rect 1702 377 1708 378
rect 1702 373 1703 377
rect 1707 373 1708 377
rect 1702 372 1708 373
rect 1902 377 1908 378
rect 1902 373 1903 377
rect 1907 373 1908 377
rect 1902 372 1908 373
rect 2006 376 2012 377
rect 2006 372 2007 376
rect 2011 372 2012 376
rect 2462 373 2468 374
rect 110 371 116 372
rect 112 347 114 371
rect 136 347 138 372
rect 288 347 290 372
rect 448 347 450 372
rect 600 347 602 372
rect 752 347 754 372
rect 904 347 906 372
rect 1080 347 1082 372
rect 1272 347 1274 372
rect 1480 347 1482 372
rect 1704 347 1706 372
rect 1904 347 1906 372
rect 2006 371 2012 372
rect 2046 372 2052 373
rect 2008 347 2010 371
rect 2046 368 2047 372
rect 2051 368 2052 372
rect 2462 369 2463 373
rect 2467 369 2468 373
rect 2462 368 2468 369
rect 2558 373 2564 374
rect 2558 369 2559 373
rect 2563 369 2564 373
rect 2558 368 2564 369
rect 2654 373 2660 374
rect 2654 369 2655 373
rect 2659 369 2660 373
rect 2654 368 2660 369
rect 2750 373 2756 374
rect 2750 369 2751 373
rect 2755 369 2756 373
rect 2750 368 2756 369
rect 2846 373 2852 374
rect 2846 369 2847 373
rect 2851 369 2852 373
rect 2846 368 2852 369
rect 2942 373 2948 374
rect 2942 369 2943 373
rect 2947 369 2948 373
rect 2942 368 2948 369
rect 3038 373 3044 374
rect 3038 369 3039 373
rect 3043 369 3044 373
rect 3038 368 3044 369
rect 3134 373 3140 374
rect 3134 369 3135 373
rect 3139 369 3140 373
rect 3134 368 3140 369
rect 3230 373 3236 374
rect 3230 369 3231 373
rect 3235 369 3236 373
rect 3230 368 3236 369
rect 3942 372 3948 373
rect 3942 368 3943 372
rect 3947 368 3948 372
rect 2046 367 2052 368
rect 2048 347 2050 367
rect 2464 347 2466 368
rect 2560 347 2562 368
rect 2656 347 2658 368
rect 2752 347 2754 368
rect 2848 347 2850 368
rect 2944 347 2946 368
rect 3040 347 3042 368
rect 3136 347 3138 368
rect 3232 347 3234 368
rect 3942 367 3948 368
rect 3944 347 3946 367
rect 111 346 115 347
rect 111 341 115 342
rect 135 346 139 347
rect 135 341 139 342
rect 159 346 163 347
rect 159 341 163 342
rect 287 346 291 347
rect 287 341 291 342
rect 351 346 355 347
rect 351 341 355 342
rect 447 346 451 347
rect 447 341 451 342
rect 551 346 555 347
rect 551 341 555 342
rect 599 346 603 347
rect 599 341 603 342
rect 751 346 755 347
rect 751 341 755 342
rect 759 346 763 347
rect 759 341 763 342
rect 903 346 907 347
rect 903 341 907 342
rect 959 346 963 347
rect 959 341 963 342
rect 1079 346 1083 347
rect 1079 341 1083 342
rect 1159 346 1163 347
rect 1159 341 1163 342
rect 1271 346 1275 347
rect 1271 341 1275 342
rect 1343 346 1347 347
rect 1343 341 1347 342
rect 1479 346 1483 347
rect 1479 341 1483 342
rect 1527 346 1531 347
rect 1527 341 1531 342
rect 1703 346 1707 347
rect 1703 341 1707 342
rect 1711 346 1715 347
rect 1711 341 1715 342
rect 1895 346 1899 347
rect 1895 341 1899 342
rect 1903 346 1907 347
rect 1903 341 1907 342
rect 2007 346 2011 347
rect 2007 341 2011 342
rect 2047 346 2051 347
rect 2047 341 2051 342
rect 2399 346 2403 347
rect 2399 341 2403 342
rect 2463 346 2467 347
rect 2463 341 2467 342
rect 2503 346 2507 347
rect 2503 341 2507 342
rect 2559 346 2563 347
rect 2559 341 2563 342
rect 2623 346 2627 347
rect 2623 341 2627 342
rect 2655 346 2659 347
rect 2655 341 2659 342
rect 2751 346 2755 347
rect 2751 341 2755 342
rect 2759 346 2763 347
rect 2759 341 2763 342
rect 2847 346 2851 347
rect 2847 341 2851 342
rect 2911 346 2915 347
rect 2911 341 2915 342
rect 2943 346 2947 347
rect 2943 341 2947 342
rect 3039 346 3043 347
rect 3039 341 3043 342
rect 3071 346 3075 347
rect 3071 341 3075 342
rect 3135 346 3139 347
rect 3135 341 3139 342
rect 3231 346 3235 347
rect 3231 341 3235 342
rect 3247 346 3251 347
rect 3247 341 3251 342
rect 3423 346 3427 347
rect 3423 341 3427 342
rect 3607 346 3611 347
rect 3607 341 3611 342
rect 3791 346 3795 347
rect 3791 341 3795 342
rect 3943 346 3947 347
rect 3943 341 3947 342
rect 112 321 114 341
rect 110 320 116 321
rect 160 320 162 341
rect 352 320 354 341
rect 552 320 554 341
rect 760 320 762 341
rect 960 320 962 341
rect 1160 320 1162 341
rect 1344 320 1346 341
rect 1528 320 1530 341
rect 1712 320 1714 341
rect 1896 320 1898 341
rect 2008 321 2010 341
rect 2048 321 2050 341
rect 2006 320 2012 321
rect 110 316 111 320
rect 115 316 116 320
rect 110 315 116 316
rect 158 319 164 320
rect 158 315 159 319
rect 163 315 164 319
rect 158 314 164 315
rect 350 319 356 320
rect 350 315 351 319
rect 355 315 356 319
rect 350 314 356 315
rect 550 319 556 320
rect 550 315 551 319
rect 555 315 556 319
rect 550 314 556 315
rect 758 319 764 320
rect 758 315 759 319
rect 763 315 764 319
rect 758 314 764 315
rect 958 319 964 320
rect 958 315 959 319
rect 963 315 964 319
rect 958 314 964 315
rect 1158 319 1164 320
rect 1158 315 1159 319
rect 1163 315 1164 319
rect 1158 314 1164 315
rect 1342 319 1348 320
rect 1342 315 1343 319
rect 1347 315 1348 319
rect 1342 314 1348 315
rect 1526 319 1532 320
rect 1526 315 1527 319
rect 1531 315 1532 319
rect 1526 314 1532 315
rect 1710 319 1716 320
rect 1710 315 1711 319
rect 1715 315 1716 319
rect 1710 314 1716 315
rect 1894 319 1900 320
rect 1894 315 1895 319
rect 1899 315 1900 319
rect 2006 316 2007 320
rect 2011 316 2012 320
rect 2006 315 2012 316
rect 2046 320 2052 321
rect 2400 320 2402 341
rect 2504 320 2506 341
rect 2624 320 2626 341
rect 2760 320 2762 341
rect 2912 320 2914 341
rect 3072 320 3074 341
rect 3248 320 3250 341
rect 3424 320 3426 341
rect 3608 320 3610 341
rect 3792 320 3794 341
rect 3944 321 3946 341
rect 3942 320 3948 321
rect 2046 316 2047 320
rect 2051 316 2052 320
rect 2046 315 2052 316
rect 2398 319 2404 320
rect 2398 315 2399 319
rect 2403 315 2404 319
rect 1894 314 1900 315
rect 2398 314 2404 315
rect 2502 319 2508 320
rect 2502 315 2503 319
rect 2507 315 2508 319
rect 2502 314 2508 315
rect 2622 319 2628 320
rect 2622 315 2623 319
rect 2627 315 2628 319
rect 2622 314 2628 315
rect 2758 319 2764 320
rect 2758 315 2759 319
rect 2763 315 2764 319
rect 2758 314 2764 315
rect 2910 319 2916 320
rect 2910 315 2911 319
rect 2915 315 2916 319
rect 2910 314 2916 315
rect 3070 319 3076 320
rect 3070 315 3071 319
rect 3075 315 3076 319
rect 3070 314 3076 315
rect 3246 319 3252 320
rect 3246 315 3247 319
rect 3251 315 3252 319
rect 3246 314 3252 315
rect 3422 319 3428 320
rect 3422 315 3423 319
rect 3427 315 3428 319
rect 3422 314 3428 315
rect 3606 319 3612 320
rect 3606 315 3607 319
rect 3611 315 3612 319
rect 3606 314 3612 315
rect 3790 319 3796 320
rect 3790 315 3791 319
rect 3795 315 3796 319
rect 3942 316 3943 320
rect 3947 316 3948 320
rect 3942 315 3948 316
rect 3790 314 3796 315
rect 110 303 116 304
rect 110 299 111 303
rect 115 299 116 303
rect 2006 303 2012 304
rect 110 298 116 299
rect 158 300 164 301
rect 112 263 114 298
rect 158 296 159 300
rect 163 296 164 300
rect 158 295 164 296
rect 350 300 356 301
rect 350 296 351 300
rect 355 296 356 300
rect 350 295 356 296
rect 550 300 556 301
rect 550 296 551 300
rect 555 296 556 300
rect 550 295 556 296
rect 758 300 764 301
rect 758 296 759 300
rect 763 296 764 300
rect 758 295 764 296
rect 958 300 964 301
rect 958 296 959 300
rect 963 296 964 300
rect 958 295 964 296
rect 1158 300 1164 301
rect 1158 296 1159 300
rect 1163 296 1164 300
rect 1158 295 1164 296
rect 1342 300 1348 301
rect 1342 296 1343 300
rect 1347 296 1348 300
rect 1342 295 1348 296
rect 1526 300 1532 301
rect 1526 296 1527 300
rect 1531 296 1532 300
rect 1526 295 1532 296
rect 1710 300 1716 301
rect 1710 296 1711 300
rect 1715 296 1716 300
rect 1710 295 1716 296
rect 1894 300 1900 301
rect 1894 296 1895 300
rect 1899 296 1900 300
rect 2006 299 2007 303
rect 2011 299 2012 303
rect 2006 298 2012 299
rect 2046 303 2052 304
rect 2046 299 2047 303
rect 2051 299 2052 303
rect 3942 303 3948 304
rect 2046 298 2052 299
rect 2398 300 2404 301
rect 1894 295 1900 296
rect 160 263 162 295
rect 352 263 354 295
rect 552 263 554 295
rect 760 263 762 295
rect 960 263 962 295
rect 1160 263 1162 295
rect 1344 263 1346 295
rect 1528 263 1530 295
rect 1712 263 1714 295
rect 1896 263 1898 295
rect 2008 263 2010 298
rect 2048 271 2050 298
rect 2398 296 2399 300
rect 2403 296 2404 300
rect 2398 295 2404 296
rect 2502 300 2508 301
rect 2502 296 2503 300
rect 2507 296 2508 300
rect 2502 295 2508 296
rect 2622 300 2628 301
rect 2622 296 2623 300
rect 2627 296 2628 300
rect 2622 295 2628 296
rect 2758 300 2764 301
rect 2758 296 2759 300
rect 2763 296 2764 300
rect 2758 295 2764 296
rect 2910 300 2916 301
rect 2910 296 2911 300
rect 2915 296 2916 300
rect 2910 295 2916 296
rect 3070 300 3076 301
rect 3070 296 3071 300
rect 3075 296 3076 300
rect 3070 295 3076 296
rect 3246 300 3252 301
rect 3246 296 3247 300
rect 3251 296 3252 300
rect 3246 295 3252 296
rect 3422 300 3428 301
rect 3422 296 3423 300
rect 3427 296 3428 300
rect 3422 295 3428 296
rect 3606 300 3612 301
rect 3606 296 3607 300
rect 3611 296 3612 300
rect 3606 295 3612 296
rect 3790 300 3796 301
rect 3790 296 3791 300
rect 3795 296 3796 300
rect 3942 299 3943 303
rect 3947 299 3948 303
rect 3942 298 3948 299
rect 3790 295 3796 296
rect 2400 271 2402 295
rect 2504 271 2506 295
rect 2624 271 2626 295
rect 2760 271 2762 295
rect 2912 271 2914 295
rect 3072 271 3074 295
rect 3248 271 3250 295
rect 3424 271 3426 295
rect 3608 271 3610 295
rect 3792 271 3794 295
rect 3944 271 3946 298
rect 2047 270 2051 271
rect 2047 265 2051 266
rect 2191 270 2195 271
rect 2191 265 2195 266
rect 2351 270 2355 271
rect 2351 265 2355 266
rect 2399 270 2403 271
rect 2399 265 2403 266
rect 2503 270 2507 271
rect 2503 265 2507 266
rect 2519 270 2523 271
rect 2519 265 2523 266
rect 2623 270 2627 271
rect 2623 265 2627 266
rect 2687 270 2691 271
rect 2687 265 2691 266
rect 2759 270 2763 271
rect 2759 265 2763 266
rect 2855 270 2859 271
rect 2855 265 2859 266
rect 2911 270 2915 271
rect 2911 265 2915 266
rect 3031 270 3035 271
rect 3031 265 3035 266
rect 3071 270 3075 271
rect 3071 265 3075 266
rect 3215 270 3219 271
rect 3215 265 3219 266
rect 3247 270 3251 271
rect 3247 265 3251 266
rect 3407 270 3411 271
rect 3407 265 3411 266
rect 3423 270 3427 271
rect 3423 265 3427 266
rect 3607 270 3611 271
rect 3607 265 3611 266
rect 3791 270 3795 271
rect 3791 265 3795 266
rect 3807 270 3811 271
rect 3807 265 3811 266
rect 3943 270 3947 271
rect 3943 265 3947 266
rect 111 262 115 263
rect 111 257 115 258
rect 159 262 163 263
rect 159 257 163 258
rect 223 262 227 263
rect 223 257 227 258
rect 351 262 355 263
rect 351 257 355 258
rect 383 262 387 263
rect 383 257 387 258
rect 543 262 547 263
rect 543 257 547 258
rect 551 262 555 263
rect 551 257 555 258
rect 703 262 707 263
rect 703 257 707 258
rect 759 262 763 263
rect 759 257 763 258
rect 863 262 867 263
rect 863 257 867 258
rect 959 262 963 263
rect 959 257 963 258
rect 1031 262 1035 263
rect 1031 257 1035 258
rect 1159 262 1163 263
rect 1159 257 1163 258
rect 1199 262 1203 263
rect 1199 257 1203 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1367 262 1371 263
rect 1367 257 1371 258
rect 1527 262 1531 263
rect 1527 257 1531 258
rect 1543 262 1547 263
rect 1543 257 1547 258
rect 1711 262 1715 263
rect 1711 257 1715 258
rect 1727 262 1731 263
rect 1727 257 1731 258
rect 1895 262 1899 263
rect 1895 257 1899 258
rect 1903 262 1907 263
rect 1903 257 1907 258
rect 2007 262 2011 263
rect 2007 257 2011 258
rect 112 230 114 257
rect 224 233 226 257
rect 384 233 386 257
rect 544 233 546 257
rect 704 233 706 257
rect 864 233 866 257
rect 1032 233 1034 257
rect 1200 233 1202 257
rect 1368 233 1370 257
rect 1544 233 1546 257
rect 1728 233 1730 257
rect 1904 233 1906 257
rect 222 232 228 233
rect 110 229 116 230
rect 110 225 111 229
rect 115 225 116 229
rect 222 228 223 232
rect 227 228 228 232
rect 222 227 228 228
rect 382 232 388 233
rect 382 228 383 232
rect 387 228 388 232
rect 382 227 388 228
rect 542 232 548 233
rect 542 228 543 232
rect 547 228 548 232
rect 542 227 548 228
rect 702 232 708 233
rect 702 228 703 232
rect 707 228 708 232
rect 702 227 708 228
rect 862 232 868 233
rect 862 228 863 232
rect 867 228 868 232
rect 862 227 868 228
rect 1030 232 1036 233
rect 1030 228 1031 232
rect 1035 228 1036 232
rect 1030 227 1036 228
rect 1198 232 1204 233
rect 1198 228 1199 232
rect 1203 228 1204 232
rect 1198 227 1204 228
rect 1366 232 1372 233
rect 1366 228 1367 232
rect 1371 228 1372 232
rect 1366 227 1372 228
rect 1542 232 1548 233
rect 1542 228 1543 232
rect 1547 228 1548 232
rect 1542 227 1548 228
rect 1726 232 1732 233
rect 1726 228 1727 232
rect 1731 228 1732 232
rect 1726 227 1732 228
rect 1902 232 1908 233
rect 1902 228 1903 232
rect 1907 228 1908 232
rect 2008 230 2010 257
rect 2048 238 2050 265
rect 2192 241 2194 265
rect 2352 241 2354 265
rect 2520 241 2522 265
rect 2688 241 2690 265
rect 2856 241 2858 265
rect 3032 241 3034 265
rect 3216 241 3218 265
rect 3408 241 3410 265
rect 3608 241 3610 265
rect 3808 241 3810 265
rect 2190 240 2196 241
rect 2046 237 2052 238
rect 2046 233 2047 237
rect 2051 233 2052 237
rect 2190 236 2191 240
rect 2195 236 2196 240
rect 2190 235 2196 236
rect 2350 240 2356 241
rect 2350 236 2351 240
rect 2355 236 2356 240
rect 2350 235 2356 236
rect 2518 240 2524 241
rect 2518 236 2519 240
rect 2523 236 2524 240
rect 2518 235 2524 236
rect 2686 240 2692 241
rect 2686 236 2687 240
rect 2691 236 2692 240
rect 2686 235 2692 236
rect 2854 240 2860 241
rect 2854 236 2855 240
rect 2859 236 2860 240
rect 2854 235 2860 236
rect 3030 240 3036 241
rect 3030 236 3031 240
rect 3035 236 3036 240
rect 3030 235 3036 236
rect 3214 240 3220 241
rect 3214 236 3215 240
rect 3219 236 3220 240
rect 3214 235 3220 236
rect 3406 240 3412 241
rect 3406 236 3407 240
rect 3411 236 3412 240
rect 3406 235 3412 236
rect 3606 240 3612 241
rect 3606 236 3607 240
rect 3611 236 3612 240
rect 3606 235 3612 236
rect 3806 240 3812 241
rect 3806 236 3807 240
rect 3811 236 3812 240
rect 3944 238 3946 265
rect 3806 235 3812 236
rect 3942 237 3948 238
rect 2046 232 2052 233
rect 3942 233 3943 237
rect 3947 233 3948 237
rect 3942 232 3948 233
rect 1902 227 1908 228
rect 2006 229 2012 230
rect 110 224 116 225
rect 2006 225 2007 229
rect 2011 225 2012 229
rect 2006 224 2012 225
rect 2190 221 2196 222
rect 2046 220 2052 221
rect 2046 216 2047 220
rect 2051 216 2052 220
rect 2190 217 2191 221
rect 2195 217 2196 221
rect 2190 216 2196 217
rect 2350 221 2356 222
rect 2350 217 2351 221
rect 2355 217 2356 221
rect 2350 216 2356 217
rect 2518 221 2524 222
rect 2518 217 2519 221
rect 2523 217 2524 221
rect 2518 216 2524 217
rect 2686 221 2692 222
rect 2686 217 2687 221
rect 2691 217 2692 221
rect 2686 216 2692 217
rect 2854 221 2860 222
rect 2854 217 2855 221
rect 2859 217 2860 221
rect 2854 216 2860 217
rect 3030 221 3036 222
rect 3030 217 3031 221
rect 3035 217 3036 221
rect 3030 216 3036 217
rect 3214 221 3220 222
rect 3214 217 3215 221
rect 3219 217 3220 221
rect 3214 216 3220 217
rect 3406 221 3412 222
rect 3406 217 3407 221
rect 3411 217 3412 221
rect 3406 216 3412 217
rect 3606 221 3612 222
rect 3606 217 3607 221
rect 3611 217 3612 221
rect 3606 216 3612 217
rect 3806 221 3812 222
rect 3806 217 3807 221
rect 3811 217 3812 221
rect 3806 216 3812 217
rect 3942 220 3948 221
rect 3942 216 3943 220
rect 3947 216 3948 220
rect 2046 215 2052 216
rect 222 213 228 214
rect 110 212 116 213
rect 110 208 111 212
rect 115 208 116 212
rect 222 209 223 213
rect 227 209 228 213
rect 222 208 228 209
rect 382 213 388 214
rect 382 209 383 213
rect 387 209 388 213
rect 382 208 388 209
rect 542 213 548 214
rect 542 209 543 213
rect 547 209 548 213
rect 542 208 548 209
rect 702 213 708 214
rect 702 209 703 213
rect 707 209 708 213
rect 702 208 708 209
rect 862 213 868 214
rect 862 209 863 213
rect 867 209 868 213
rect 862 208 868 209
rect 1030 213 1036 214
rect 1030 209 1031 213
rect 1035 209 1036 213
rect 1030 208 1036 209
rect 1198 213 1204 214
rect 1198 209 1199 213
rect 1203 209 1204 213
rect 1198 208 1204 209
rect 1366 213 1372 214
rect 1366 209 1367 213
rect 1371 209 1372 213
rect 1366 208 1372 209
rect 1542 213 1548 214
rect 1542 209 1543 213
rect 1547 209 1548 213
rect 1542 208 1548 209
rect 1726 213 1732 214
rect 1726 209 1727 213
rect 1731 209 1732 213
rect 1726 208 1732 209
rect 1902 213 1908 214
rect 1902 209 1903 213
rect 1907 209 1908 213
rect 1902 208 1908 209
rect 2006 212 2012 213
rect 2006 208 2007 212
rect 2011 208 2012 212
rect 110 207 116 208
rect 112 167 114 207
rect 224 167 226 208
rect 384 167 386 208
rect 544 167 546 208
rect 704 167 706 208
rect 864 167 866 208
rect 1032 167 1034 208
rect 1200 167 1202 208
rect 1368 167 1370 208
rect 1544 167 1546 208
rect 1728 167 1730 208
rect 1904 167 1906 208
rect 2006 207 2012 208
rect 2008 167 2010 207
rect 111 166 115 167
rect 111 161 115 162
rect 135 166 139 167
rect 135 161 139 162
rect 223 166 227 167
rect 223 161 227 162
rect 231 166 235 167
rect 231 161 235 162
rect 327 166 331 167
rect 327 161 331 162
rect 383 166 387 167
rect 383 161 387 162
rect 423 166 427 167
rect 423 161 427 162
rect 527 166 531 167
rect 527 161 531 162
rect 543 166 547 167
rect 543 161 547 162
rect 647 166 651 167
rect 647 161 651 162
rect 703 166 707 167
rect 703 161 707 162
rect 775 166 779 167
rect 775 161 779 162
rect 863 166 867 167
rect 863 161 867 162
rect 903 166 907 167
rect 903 161 907 162
rect 1031 166 1035 167
rect 1031 161 1035 162
rect 1151 166 1155 167
rect 1151 161 1155 162
rect 1199 166 1203 167
rect 1199 161 1203 162
rect 1271 166 1275 167
rect 1271 161 1275 162
rect 1367 166 1371 167
rect 1367 161 1371 162
rect 1383 166 1387 167
rect 1383 161 1387 162
rect 1487 166 1491 167
rect 1487 161 1491 162
rect 1543 166 1547 167
rect 1543 161 1547 162
rect 1591 166 1595 167
rect 1591 161 1595 162
rect 1703 166 1707 167
rect 1703 161 1707 162
rect 1727 166 1731 167
rect 1727 161 1731 162
rect 1807 166 1811 167
rect 1807 161 1811 162
rect 1903 166 1907 167
rect 1903 161 1907 162
rect 2007 166 2011 167
rect 2048 163 2050 215
rect 2192 163 2194 216
rect 2352 163 2354 216
rect 2520 163 2522 216
rect 2688 163 2690 216
rect 2856 163 2858 216
rect 3032 163 3034 216
rect 3216 163 3218 216
rect 3408 163 3410 216
rect 3608 163 3610 216
rect 3808 163 3810 216
rect 3942 215 3948 216
rect 3944 163 3946 215
rect 2007 161 2011 162
rect 2047 162 2051 163
rect 112 141 114 161
rect 110 140 116 141
rect 136 140 138 161
rect 232 140 234 161
rect 328 140 330 161
rect 424 140 426 161
rect 528 140 530 161
rect 648 140 650 161
rect 776 140 778 161
rect 904 140 906 161
rect 1032 140 1034 161
rect 1152 140 1154 161
rect 1272 140 1274 161
rect 1384 140 1386 161
rect 1488 140 1490 161
rect 1592 140 1594 161
rect 1704 140 1706 161
rect 1808 140 1810 161
rect 1904 140 1906 161
rect 2008 141 2010 161
rect 2047 157 2051 158
rect 2071 162 2075 163
rect 2071 157 2075 158
rect 2167 162 2171 163
rect 2167 157 2171 158
rect 2191 162 2195 163
rect 2191 157 2195 158
rect 2263 162 2267 163
rect 2263 157 2267 158
rect 2351 162 2355 163
rect 2351 157 2355 158
rect 2367 162 2371 163
rect 2367 157 2371 158
rect 2487 162 2491 163
rect 2487 157 2491 158
rect 2519 162 2523 163
rect 2519 157 2523 158
rect 2615 162 2619 163
rect 2615 157 2619 158
rect 2687 162 2691 163
rect 2687 157 2691 158
rect 2743 162 2747 163
rect 2743 157 2747 158
rect 2855 162 2859 163
rect 2855 157 2859 158
rect 2871 162 2875 163
rect 2871 157 2875 158
rect 2991 162 2995 163
rect 2991 157 2995 158
rect 3031 162 3035 163
rect 3031 157 3035 158
rect 3111 162 3115 163
rect 3111 157 3115 158
rect 3215 162 3219 163
rect 3215 157 3219 158
rect 3223 162 3227 163
rect 3223 157 3227 158
rect 3327 162 3331 163
rect 3327 157 3331 158
rect 3407 162 3411 163
rect 3407 157 3411 158
rect 3431 162 3435 163
rect 3431 157 3435 158
rect 3535 162 3539 163
rect 3535 157 3539 158
rect 3607 162 3611 163
rect 3607 157 3611 158
rect 3639 162 3643 163
rect 3639 157 3643 158
rect 3743 162 3747 163
rect 3743 157 3747 158
rect 3807 162 3811 163
rect 3807 157 3811 158
rect 3839 162 3843 163
rect 3839 157 3843 158
rect 3943 162 3947 163
rect 3943 157 3947 158
rect 2006 140 2012 141
rect 110 136 111 140
rect 115 136 116 140
rect 110 135 116 136
rect 134 139 140 140
rect 134 135 135 139
rect 139 135 140 139
rect 134 134 140 135
rect 230 139 236 140
rect 230 135 231 139
rect 235 135 236 139
rect 230 134 236 135
rect 326 139 332 140
rect 326 135 327 139
rect 331 135 332 139
rect 326 134 332 135
rect 422 139 428 140
rect 422 135 423 139
rect 427 135 428 139
rect 422 134 428 135
rect 526 139 532 140
rect 526 135 527 139
rect 531 135 532 139
rect 526 134 532 135
rect 646 139 652 140
rect 646 135 647 139
rect 651 135 652 139
rect 646 134 652 135
rect 774 139 780 140
rect 774 135 775 139
rect 779 135 780 139
rect 774 134 780 135
rect 902 139 908 140
rect 902 135 903 139
rect 907 135 908 139
rect 902 134 908 135
rect 1030 139 1036 140
rect 1030 135 1031 139
rect 1035 135 1036 139
rect 1030 134 1036 135
rect 1150 139 1156 140
rect 1150 135 1151 139
rect 1155 135 1156 139
rect 1150 134 1156 135
rect 1270 139 1276 140
rect 1270 135 1271 139
rect 1275 135 1276 139
rect 1270 134 1276 135
rect 1382 139 1388 140
rect 1382 135 1383 139
rect 1387 135 1388 139
rect 1382 134 1388 135
rect 1486 139 1492 140
rect 1486 135 1487 139
rect 1491 135 1492 139
rect 1486 134 1492 135
rect 1590 139 1596 140
rect 1590 135 1591 139
rect 1595 135 1596 139
rect 1590 134 1596 135
rect 1702 139 1708 140
rect 1702 135 1703 139
rect 1707 135 1708 139
rect 1702 134 1708 135
rect 1806 139 1812 140
rect 1806 135 1807 139
rect 1811 135 1812 139
rect 1806 134 1812 135
rect 1902 139 1908 140
rect 1902 135 1903 139
rect 1907 135 1908 139
rect 2006 136 2007 140
rect 2011 136 2012 140
rect 2048 137 2050 157
rect 2006 135 2012 136
rect 2046 136 2052 137
rect 2072 136 2074 157
rect 2168 136 2170 157
rect 2264 136 2266 157
rect 2368 136 2370 157
rect 2488 136 2490 157
rect 2616 136 2618 157
rect 2744 136 2746 157
rect 2872 136 2874 157
rect 2992 136 2994 157
rect 3112 136 3114 157
rect 3224 136 3226 157
rect 3328 136 3330 157
rect 3432 136 3434 157
rect 3536 136 3538 157
rect 3640 136 3642 157
rect 3744 136 3746 157
rect 3840 136 3842 157
rect 3944 137 3946 157
rect 3942 136 3948 137
rect 1902 134 1908 135
rect 2046 132 2047 136
rect 2051 132 2052 136
rect 2046 131 2052 132
rect 2070 135 2076 136
rect 2070 131 2071 135
rect 2075 131 2076 135
rect 2070 130 2076 131
rect 2166 135 2172 136
rect 2166 131 2167 135
rect 2171 131 2172 135
rect 2166 130 2172 131
rect 2262 135 2268 136
rect 2262 131 2263 135
rect 2267 131 2268 135
rect 2262 130 2268 131
rect 2366 135 2372 136
rect 2366 131 2367 135
rect 2371 131 2372 135
rect 2366 130 2372 131
rect 2486 135 2492 136
rect 2486 131 2487 135
rect 2491 131 2492 135
rect 2486 130 2492 131
rect 2614 135 2620 136
rect 2614 131 2615 135
rect 2619 131 2620 135
rect 2614 130 2620 131
rect 2742 135 2748 136
rect 2742 131 2743 135
rect 2747 131 2748 135
rect 2742 130 2748 131
rect 2870 135 2876 136
rect 2870 131 2871 135
rect 2875 131 2876 135
rect 2870 130 2876 131
rect 2990 135 2996 136
rect 2990 131 2991 135
rect 2995 131 2996 135
rect 2990 130 2996 131
rect 3110 135 3116 136
rect 3110 131 3111 135
rect 3115 131 3116 135
rect 3110 130 3116 131
rect 3222 135 3228 136
rect 3222 131 3223 135
rect 3227 131 3228 135
rect 3222 130 3228 131
rect 3326 135 3332 136
rect 3326 131 3327 135
rect 3331 131 3332 135
rect 3326 130 3332 131
rect 3430 135 3436 136
rect 3430 131 3431 135
rect 3435 131 3436 135
rect 3430 130 3436 131
rect 3534 135 3540 136
rect 3534 131 3535 135
rect 3539 131 3540 135
rect 3534 130 3540 131
rect 3638 135 3644 136
rect 3638 131 3639 135
rect 3643 131 3644 135
rect 3638 130 3644 131
rect 3742 135 3748 136
rect 3742 131 3743 135
rect 3747 131 3748 135
rect 3742 130 3748 131
rect 3838 135 3844 136
rect 3838 131 3839 135
rect 3843 131 3844 135
rect 3942 132 3943 136
rect 3947 132 3948 136
rect 3942 131 3948 132
rect 3838 130 3844 131
rect 110 123 116 124
rect 110 119 111 123
rect 115 119 116 123
rect 2006 123 2012 124
rect 110 118 116 119
rect 134 120 140 121
rect 112 91 114 118
rect 134 116 135 120
rect 139 116 140 120
rect 134 115 140 116
rect 230 120 236 121
rect 230 116 231 120
rect 235 116 236 120
rect 230 115 236 116
rect 326 120 332 121
rect 326 116 327 120
rect 331 116 332 120
rect 326 115 332 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 526 120 532 121
rect 526 116 527 120
rect 531 116 532 120
rect 526 115 532 116
rect 646 120 652 121
rect 646 116 647 120
rect 651 116 652 120
rect 646 115 652 116
rect 774 120 780 121
rect 774 116 775 120
rect 779 116 780 120
rect 774 115 780 116
rect 902 120 908 121
rect 902 116 903 120
rect 907 116 908 120
rect 902 115 908 116
rect 1030 120 1036 121
rect 1030 116 1031 120
rect 1035 116 1036 120
rect 1030 115 1036 116
rect 1150 120 1156 121
rect 1150 116 1151 120
rect 1155 116 1156 120
rect 1150 115 1156 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1382 120 1388 121
rect 1382 116 1383 120
rect 1387 116 1388 120
rect 1382 115 1388 116
rect 1486 120 1492 121
rect 1486 116 1487 120
rect 1491 116 1492 120
rect 1486 115 1492 116
rect 1590 120 1596 121
rect 1590 116 1591 120
rect 1595 116 1596 120
rect 1590 115 1596 116
rect 1702 120 1708 121
rect 1702 116 1703 120
rect 1707 116 1708 120
rect 1702 115 1708 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 2006 119 2007 123
rect 2011 119 2012 123
rect 2006 118 2012 119
rect 2046 119 2052 120
rect 1902 115 1908 116
rect 136 91 138 115
rect 232 91 234 115
rect 328 91 330 115
rect 424 91 426 115
rect 528 91 530 115
rect 648 91 650 115
rect 776 91 778 115
rect 904 91 906 115
rect 1032 91 1034 115
rect 1152 91 1154 115
rect 1272 91 1274 115
rect 1384 91 1386 115
rect 1488 91 1490 115
rect 1592 91 1594 115
rect 1704 91 1706 115
rect 1808 91 1810 115
rect 1904 91 1906 115
rect 2008 91 2010 118
rect 2046 115 2047 119
rect 2051 115 2052 119
rect 3942 119 3948 120
rect 2046 114 2052 115
rect 2070 116 2076 117
rect 111 90 115 91
rect 111 85 115 86
rect 135 90 139 91
rect 135 85 139 86
rect 231 90 235 91
rect 231 85 235 86
rect 327 90 331 91
rect 327 85 331 86
rect 423 90 427 91
rect 423 85 427 86
rect 527 90 531 91
rect 527 85 531 86
rect 647 90 651 91
rect 647 85 651 86
rect 775 90 779 91
rect 775 85 779 86
rect 903 90 907 91
rect 903 85 907 86
rect 1031 90 1035 91
rect 1031 85 1035 86
rect 1151 90 1155 91
rect 1151 85 1155 86
rect 1271 90 1275 91
rect 1271 85 1275 86
rect 1383 90 1387 91
rect 1383 85 1387 86
rect 1487 90 1491 91
rect 1487 85 1491 86
rect 1591 90 1595 91
rect 1591 85 1595 86
rect 1703 90 1707 91
rect 1703 85 1707 86
rect 1807 90 1811 91
rect 1807 85 1811 86
rect 1903 90 1907 91
rect 1903 85 1907 86
rect 2007 90 2011 91
rect 2048 87 2050 114
rect 2070 112 2071 116
rect 2075 112 2076 116
rect 2070 111 2076 112
rect 2166 116 2172 117
rect 2166 112 2167 116
rect 2171 112 2172 116
rect 2166 111 2172 112
rect 2262 116 2268 117
rect 2262 112 2263 116
rect 2267 112 2268 116
rect 2262 111 2268 112
rect 2366 116 2372 117
rect 2366 112 2367 116
rect 2371 112 2372 116
rect 2366 111 2372 112
rect 2486 116 2492 117
rect 2486 112 2487 116
rect 2491 112 2492 116
rect 2486 111 2492 112
rect 2614 116 2620 117
rect 2614 112 2615 116
rect 2619 112 2620 116
rect 2614 111 2620 112
rect 2742 116 2748 117
rect 2742 112 2743 116
rect 2747 112 2748 116
rect 2742 111 2748 112
rect 2870 116 2876 117
rect 2870 112 2871 116
rect 2875 112 2876 116
rect 2870 111 2876 112
rect 2990 116 2996 117
rect 2990 112 2991 116
rect 2995 112 2996 116
rect 2990 111 2996 112
rect 3110 116 3116 117
rect 3110 112 3111 116
rect 3115 112 3116 116
rect 3110 111 3116 112
rect 3222 116 3228 117
rect 3222 112 3223 116
rect 3227 112 3228 116
rect 3222 111 3228 112
rect 3326 116 3332 117
rect 3326 112 3327 116
rect 3331 112 3332 116
rect 3326 111 3332 112
rect 3430 116 3436 117
rect 3430 112 3431 116
rect 3435 112 3436 116
rect 3430 111 3436 112
rect 3534 116 3540 117
rect 3534 112 3535 116
rect 3539 112 3540 116
rect 3534 111 3540 112
rect 3638 116 3644 117
rect 3638 112 3639 116
rect 3643 112 3644 116
rect 3638 111 3644 112
rect 3742 116 3748 117
rect 3742 112 3743 116
rect 3747 112 3748 116
rect 3742 111 3748 112
rect 3838 116 3844 117
rect 3838 112 3839 116
rect 3843 112 3844 116
rect 3942 115 3943 119
rect 3947 115 3948 119
rect 3942 114 3948 115
rect 3838 111 3844 112
rect 2072 87 2074 111
rect 2168 87 2170 111
rect 2264 87 2266 111
rect 2368 87 2370 111
rect 2488 87 2490 111
rect 2616 87 2618 111
rect 2744 87 2746 111
rect 2872 87 2874 111
rect 2992 87 2994 111
rect 3112 87 3114 111
rect 3224 87 3226 111
rect 3328 87 3330 111
rect 3432 87 3434 111
rect 3536 87 3538 111
rect 3640 87 3642 111
rect 3744 87 3746 111
rect 3840 87 3842 111
rect 3944 87 3946 114
rect 2007 85 2011 86
rect 2047 86 2051 87
rect 2047 81 2051 82
rect 2071 86 2075 87
rect 2071 81 2075 82
rect 2167 86 2171 87
rect 2167 81 2171 82
rect 2263 86 2267 87
rect 2263 81 2267 82
rect 2367 86 2371 87
rect 2367 81 2371 82
rect 2487 86 2491 87
rect 2487 81 2491 82
rect 2615 86 2619 87
rect 2615 81 2619 82
rect 2743 86 2747 87
rect 2743 81 2747 82
rect 2871 86 2875 87
rect 2871 81 2875 82
rect 2991 86 2995 87
rect 2991 81 2995 82
rect 3111 86 3115 87
rect 3111 81 3115 82
rect 3223 86 3227 87
rect 3223 81 3227 82
rect 3327 86 3331 87
rect 3327 81 3331 82
rect 3431 86 3435 87
rect 3431 81 3435 82
rect 3535 86 3539 87
rect 3535 81 3539 82
rect 3639 86 3643 87
rect 3639 81 3643 82
rect 3743 86 3747 87
rect 3743 81 3747 82
rect 3839 86 3843 87
rect 3839 81 3843 82
rect 3943 86 3947 87
rect 3943 81 3947 82
<< m4c >>
rect 2047 4026 2051 4030
rect 2071 4026 2075 4030
rect 3943 4026 3947 4030
rect 111 4006 115 4010
rect 151 4006 155 4010
rect 279 4006 283 4010
rect 431 4006 435 4010
rect 607 4006 611 4010
rect 791 4006 795 4010
rect 975 4006 979 4010
rect 1151 4006 1155 4010
rect 1311 4006 1315 4010
rect 1471 4006 1475 4010
rect 1623 4006 1627 4010
rect 1775 4006 1779 4010
rect 1903 4006 1907 4010
rect 2007 4006 2011 4010
rect 2047 3950 2051 3954
rect 2071 3950 2075 3954
rect 2079 3950 2083 3954
rect 2215 3950 2219 3954
rect 2359 3950 2363 3954
rect 2503 3950 2507 3954
rect 2647 3950 2651 3954
rect 2791 3950 2795 3954
rect 2927 3950 2931 3954
rect 3055 3950 3059 3954
rect 3175 3950 3179 3954
rect 3295 3950 3299 3954
rect 3415 3950 3419 3954
rect 3535 3950 3539 3954
rect 3943 3950 3947 3954
rect 111 3930 115 3934
rect 151 3930 155 3934
rect 279 3930 283 3934
rect 303 3930 307 3934
rect 423 3930 427 3934
rect 431 3930 435 3934
rect 551 3930 555 3934
rect 607 3930 611 3934
rect 687 3930 691 3934
rect 791 3930 795 3934
rect 815 3930 819 3934
rect 943 3930 947 3934
rect 975 3930 979 3934
rect 1071 3930 1075 3934
rect 1151 3930 1155 3934
rect 1199 3930 1203 3934
rect 1311 3930 1315 3934
rect 1327 3930 1331 3934
rect 1463 3930 1467 3934
rect 1471 3930 1475 3934
rect 1623 3930 1627 3934
rect 1775 3930 1779 3934
rect 1903 3930 1907 3934
rect 2007 3930 2011 3934
rect 2047 3874 2051 3878
rect 2079 3874 2083 3878
rect 2215 3874 2219 3878
rect 2255 3874 2259 3878
rect 2359 3874 2363 3878
rect 2383 3874 2387 3878
rect 2503 3874 2507 3878
rect 2519 3874 2523 3878
rect 2647 3874 2651 3878
rect 2671 3874 2675 3878
rect 2791 3874 2795 3878
rect 2831 3874 2835 3878
rect 2927 3874 2931 3878
rect 2991 3874 2995 3878
rect 3055 3874 3059 3878
rect 3159 3874 3163 3878
rect 3175 3874 3179 3878
rect 3295 3874 3299 3878
rect 3327 3874 3331 3878
rect 3415 3874 3419 3878
rect 3495 3874 3499 3878
rect 3535 3874 3539 3878
rect 3663 3874 3667 3878
rect 3943 3874 3947 3878
rect 111 3850 115 3854
rect 303 3850 307 3854
rect 415 3850 419 3854
rect 423 3850 427 3854
rect 551 3850 555 3854
rect 567 3850 571 3854
rect 687 3850 691 3854
rect 727 3850 731 3854
rect 815 3850 819 3854
rect 887 3850 891 3854
rect 943 3850 947 3854
rect 1039 3850 1043 3854
rect 1071 3850 1075 3854
rect 1191 3850 1195 3854
rect 1199 3850 1203 3854
rect 1327 3850 1331 3854
rect 1343 3850 1347 3854
rect 1463 3850 1467 3854
rect 1495 3850 1499 3854
rect 1647 3850 1651 3854
rect 2007 3850 2011 3854
rect 2047 3798 2051 3802
rect 2071 3798 2075 3802
rect 2199 3798 2203 3802
rect 2255 3798 2259 3802
rect 2375 3798 2379 3802
rect 2383 3798 2387 3802
rect 2519 3798 2523 3802
rect 2559 3798 2563 3802
rect 2671 3798 2675 3802
rect 2751 3798 2755 3802
rect 2831 3798 2835 3802
rect 2951 3798 2955 3802
rect 2991 3798 2995 3802
rect 3143 3798 3147 3802
rect 3159 3798 3163 3802
rect 3327 3798 3331 3802
rect 3335 3798 3339 3802
rect 3495 3798 3499 3802
rect 3535 3798 3539 3802
rect 3663 3798 3667 3802
rect 3735 3798 3739 3802
rect 3943 3798 3947 3802
rect 111 3770 115 3774
rect 399 3770 403 3774
rect 415 3770 419 3774
rect 567 3770 571 3774
rect 727 3770 731 3774
rect 751 3770 755 3774
rect 887 3770 891 3774
rect 935 3770 939 3774
rect 1039 3770 1043 3774
rect 1127 3770 1131 3774
rect 1191 3770 1195 3774
rect 1311 3770 1315 3774
rect 1343 3770 1347 3774
rect 1495 3770 1499 3774
rect 1503 3770 1507 3774
rect 1647 3770 1651 3774
rect 1695 3770 1699 3774
rect 1887 3770 1891 3774
rect 2007 3770 2011 3774
rect 2047 3710 2051 3714
rect 2071 3710 2075 3714
rect 2199 3710 2203 3714
rect 2263 3710 2267 3714
rect 2375 3710 2379 3714
rect 2479 3710 2483 3714
rect 2559 3710 2563 3714
rect 2695 3710 2699 3714
rect 2751 3710 2755 3714
rect 2911 3710 2915 3714
rect 2951 3710 2955 3714
rect 3119 3710 3123 3714
rect 3143 3710 3147 3714
rect 3319 3710 3323 3714
rect 3335 3710 3339 3714
rect 3519 3710 3523 3714
rect 3535 3710 3539 3714
rect 3727 3710 3731 3714
rect 3735 3710 3739 3714
rect 3943 3710 3947 3714
rect 111 3682 115 3686
rect 367 3682 371 3686
rect 399 3682 403 3686
rect 519 3682 523 3686
rect 567 3682 571 3686
rect 679 3682 683 3686
rect 751 3682 755 3686
rect 847 3682 851 3686
rect 935 3682 939 3686
rect 1015 3682 1019 3686
rect 1127 3682 1131 3686
rect 1175 3682 1179 3686
rect 1311 3682 1315 3686
rect 1327 3682 1331 3686
rect 1479 3682 1483 3686
rect 1503 3682 1507 3686
rect 1631 3682 1635 3686
rect 1695 3682 1699 3686
rect 1791 3682 1795 3686
rect 1887 3682 1891 3686
rect 2007 3682 2011 3686
rect 2047 3630 2051 3634
rect 2071 3630 2075 3634
rect 2111 3630 2115 3634
rect 2263 3630 2267 3634
rect 2271 3630 2275 3634
rect 2455 3630 2459 3634
rect 2479 3630 2483 3634
rect 2655 3630 2659 3634
rect 2695 3630 2699 3634
rect 2871 3630 2875 3634
rect 2911 3630 2915 3634
rect 3095 3630 3099 3634
rect 3119 3630 3123 3634
rect 3319 3630 3323 3634
rect 3327 3630 3331 3634
rect 3519 3630 3523 3634
rect 3567 3630 3571 3634
rect 3727 3630 3731 3634
rect 3943 3630 3947 3634
rect 111 3598 115 3602
rect 271 3598 275 3602
rect 367 3598 371 3602
rect 415 3598 419 3602
rect 519 3598 523 3602
rect 575 3598 579 3602
rect 679 3598 683 3602
rect 735 3598 739 3602
rect 847 3598 851 3602
rect 895 3598 899 3602
rect 1015 3598 1019 3602
rect 1055 3598 1059 3602
rect 1175 3598 1179 3602
rect 1215 3598 1219 3602
rect 1327 3598 1331 3602
rect 1375 3598 1379 3602
rect 1479 3598 1483 3602
rect 1543 3598 1547 3602
rect 1631 3598 1635 3602
rect 1791 3598 1795 3602
rect 2007 3598 2011 3602
rect 2047 3538 2051 3542
rect 2111 3538 2115 3542
rect 2271 3538 2275 3542
rect 2287 3538 2291 3542
rect 2383 3538 2387 3542
rect 2455 3538 2459 3542
rect 2479 3538 2483 3542
rect 2575 3538 2579 3542
rect 2655 3538 2659 3542
rect 2671 3538 2675 3542
rect 2767 3538 2771 3542
rect 2871 3538 2875 3542
rect 2983 3538 2987 3542
rect 3095 3538 3099 3542
rect 3103 3538 3107 3542
rect 3223 3538 3227 3542
rect 3327 3538 3331 3542
rect 3351 3538 3355 3542
rect 3487 3538 3491 3542
rect 3567 3538 3571 3542
rect 3943 3538 3947 3542
rect 111 3514 115 3518
rect 159 3514 163 3518
rect 271 3514 275 3518
rect 287 3514 291 3518
rect 415 3514 419 3518
rect 423 3514 427 3518
rect 559 3514 563 3518
rect 575 3514 579 3518
rect 695 3514 699 3518
rect 735 3514 739 3518
rect 831 3514 835 3518
rect 895 3514 899 3518
rect 967 3514 971 3518
rect 1055 3514 1059 3518
rect 1095 3514 1099 3518
rect 1215 3514 1219 3518
rect 1231 3514 1235 3518
rect 1367 3514 1371 3518
rect 1375 3514 1379 3518
rect 1543 3514 1547 3518
rect 2007 3514 2011 3518
rect 2047 3462 2051 3466
rect 2287 3462 2291 3466
rect 2383 3462 2387 3466
rect 2479 3462 2483 3466
rect 2487 3462 2491 3466
rect 2575 3462 2579 3466
rect 2583 3462 2587 3466
rect 2671 3462 2675 3466
rect 2679 3462 2683 3466
rect 2767 3462 2771 3466
rect 2783 3462 2787 3466
rect 2871 3462 2875 3466
rect 2895 3462 2899 3466
rect 2983 3462 2987 3466
rect 3015 3462 3019 3466
rect 3103 3462 3107 3466
rect 3143 3462 3147 3466
rect 3223 3462 3227 3466
rect 3271 3462 3275 3466
rect 3351 3462 3355 3466
rect 3407 3462 3411 3466
rect 3487 3462 3491 3466
rect 3943 3462 3947 3466
rect 111 3430 115 3434
rect 135 3430 139 3434
rect 159 3430 163 3434
rect 247 3430 251 3434
rect 287 3430 291 3434
rect 383 3430 387 3434
rect 423 3430 427 3434
rect 527 3430 531 3434
rect 559 3430 563 3434
rect 671 3430 675 3434
rect 695 3430 699 3434
rect 815 3430 819 3434
rect 831 3430 835 3434
rect 967 3430 971 3434
rect 1095 3430 1099 3434
rect 1119 3430 1123 3434
rect 1231 3430 1235 3434
rect 1271 3430 1275 3434
rect 1367 3430 1371 3434
rect 2007 3430 2011 3434
rect 2047 3378 2051 3382
rect 2351 3378 2355 3382
rect 2479 3378 2483 3382
rect 2487 3378 2491 3382
rect 2583 3378 2587 3382
rect 2615 3378 2619 3382
rect 2679 3378 2683 3382
rect 2751 3378 2755 3382
rect 2783 3378 2787 3382
rect 2887 3378 2891 3382
rect 2895 3378 2899 3382
rect 3015 3378 3019 3382
rect 3023 3378 3027 3382
rect 3143 3378 3147 3382
rect 3159 3378 3163 3382
rect 3271 3378 3275 3382
rect 3303 3378 3307 3382
rect 3407 3378 3411 3382
rect 3943 3378 3947 3382
rect 111 3346 115 3350
rect 135 3346 139 3350
rect 247 3346 251 3350
rect 263 3346 267 3350
rect 383 3346 387 3350
rect 431 3346 435 3350
rect 527 3346 531 3350
rect 599 3346 603 3350
rect 671 3346 675 3350
rect 767 3346 771 3350
rect 815 3346 819 3350
rect 927 3346 931 3350
rect 967 3346 971 3350
rect 1087 3346 1091 3350
rect 1119 3346 1123 3350
rect 1239 3346 1243 3350
rect 1271 3346 1275 3350
rect 1391 3346 1395 3350
rect 1551 3346 1555 3350
rect 2007 3346 2011 3350
rect 2047 3298 2051 3302
rect 2127 3298 2131 3302
rect 2295 3298 2299 3302
rect 2351 3298 2355 3302
rect 2455 3298 2459 3302
rect 2479 3298 2483 3302
rect 2615 3298 2619 3302
rect 2751 3298 2755 3302
rect 2775 3298 2779 3302
rect 2887 3298 2891 3302
rect 2935 3298 2939 3302
rect 3023 3298 3027 3302
rect 3095 3298 3099 3302
rect 3159 3298 3163 3302
rect 3263 3298 3267 3302
rect 3303 3298 3307 3302
rect 3943 3298 3947 3302
rect 111 3262 115 3266
rect 135 3262 139 3266
rect 143 3262 147 3266
rect 263 3262 267 3266
rect 295 3262 299 3266
rect 431 3262 435 3266
rect 455 3262 459 3266
rect 599 3262 603 3266
rect 623 3262 627 3266
rect 767 3262 771 3266
rect 791 3262 795 3266
rect 927 3262 931 3266
rect 959 3262 963 3266
rect 1087 3262 1091 3266
rect 1127 3262 1131 3266
rect 1239 3262 1243 3266
rect 1303 3262 1307 3266
rect 1391 3262 1395 3266
rect 1479 3262 1483 3266
rect 1551 3262 1555 3266
rect 2007 3262 2011 3266
rect 2047 3222 2051 3226
rect 2071 3222 2075 3226
rect 2127 3222 2131 3226
rect 2207 3222 2211 3226
rect 2295 3222 2299 3226
rect 2375 3222 2379 3226
rect 2455 3222 2459 3226
rect 2543 3222 2547 3226
rect 2615 3222 2619 3226
rect 2703 3222 2707 3226
rect 2775 3222 2779 3226
rect 2863 3222 2867 3226
rect 2935 3222 2939 3226
rect 3015 3222 3019 3226
rect 3095 3222 3099 3226
rect 3167 3222 3171 3226
rect 3263 3222 3267 3226
rect 3327 3222 3331 3226
rect 3943 3222 3947 3226
rect 111 3186 115 3190
rect 143 3186 147 3190
rect 295 3186 299 3190
rect 431 3186 435 3190
rect 455 3186 459 3190
rect 567 3186 571 3190
rect 623 3186 627 3190
rect 703 3186 707 3190
rect 791 3186 795 3190
rect 855 3186 859 3190
rect 959 3186 963 3190
rect 1031 3186 1035 3190
rect 1127 3186 1131 3190
rect 1231 3186 1235 3190
rect 1303 3186 1307 3190
rect 1455 3186 1459 3190
rect 1479 3186 1483 3190
rect 1687 3186 1691 3190
rect 1903 3186 1907 3190
rect 2007 3186 2011 3190
rect 2047 3142 2051 3146
rect 2071 3142 2075 3146
rect 2207 3142 2211 3146
rect 2343 3142 2347 3146
rect 2375 3142 2379 3146
rect 2543 3142 2547 3146
rect 2631 3142 2635 3146
rect 2703 3142 2707 3146
rect 2863 3142 2867 3146
rect 2903 3142 2907 3146
rect 3015 3142 3019 3146
rect 3167 3142 3171 3146
rect 3175 3142 3179 3146
rect 3327 3142 3331 3146
rect 3447 3142 3451 3146
rect 3943 3142 3947 3146
rect 111 3110 115 3114
rect 295 3110 299 3114
rect 311 3110 315 3114
rect 407 3110 411 3114
rect 431 3110 435 3114
rect 503 3110 507 3114
rect 567 3110 571 3114
rect 599 3110 603 3114
rect 695 3110 699 3114
rect 703 3110 707 3114
rect 807 3110 811 3114
rect 855 3110 859 3114
rect 943 3110 947 3114
rect 1031 3110 1035 3114
rect 1087 3110 1091 3114
rect 1231 3110 1235 3114
rect 1247 3110 1251 3114
rect 1407 3110 1411 3114
rect 1455 3110 1459 3114
rect 1575 3110 1579 3114
rect 1687 3110 1691 3114
rect 1751 3110 1755 3114
rect 1903 3110 1907 3114
rect 2007 3110 2011 3114
rect 2047 3062 2051 3066
rect 2071 3062 2075 3066
rect 2343 3062 2347 3066
rect 2487 3062 2491 3066
rect 2615 3062 2619 3066
rect 2631 3062 2635 3066
rect 2743 3062 2747 3066
rect 2863 3062 2867 3066
rect 2903 3062 2907 3066
rect 2983 3062 2987 3066
rect 3103 3062 3107 3066
rect 3175 3062 3179 3066
rect 3215 3062 3219 3066
rect 3327 3062 3331 3066
rect 3431 3062 3435 3066
rect 3447 3062 3451 3066
rect 3535 3062 3539 3066
rect 3639 3062 3643 3066
rect 3743 3062 3747 3066
rect 3839 3062 3843 3066
rect 3943 3062 3947 3066
rect 111 3034 115 3038
rect 311 3034 315 3038
rect 407 3034 411 3038
rect 423 3034 427 3038
rect 503 3034 507 3038
rect 519 3034 523 3038
rect 599 3034 603 3038
rect 615 3034 619 3038
rect 695 3034 699 3038
rect 711 3034 715 3038
rect 807 3034 811 3038
rect 815 3034 819 3038
rect 935 3034 939 3038
rect 943 3034 947 3038
rect 1055 3034 1059 3038
rect 1087 3034 1091 3038
rect 1183 3034 1187 3038
rect 1247 3034 1251 3038
rect 1311 3034 1315 3038
rect 1407 3034 1411 3038
rect 1431 3034 1435 3038
rect 1551 3034 1555 3038
rect 1575 3034 1579 3038
rect 1671 3034 1675 3038
rect 1751 3034 1755 3038
rect 1799 3034 1803 3038
rect 1903 3034 1907 3038
rect 2007 3034 2011 3038
rect 2047 2982 2051 2986
rect 2407 2982 2411 2986
rect 2487 2982 2491 2986
rect 2575 2982 2579 2986
rect 2615 2982 2619 2986
rect 2743 2982 2747 2986
rect 2767 2982 2771 2986
rect 2863 2982 2867 2986
rect 2967 2982 2971 2986
rect 2983 2982 2987 2986
rect 3103 2982 3107 2986
rect 3183 2982 3187 2986
rect 3215 2982 3219 2986
rect 3327 2982 3331 2986
rect 3399 2982 3403 2986
rect 3431 2982 3435 2986
rect 3535 2982 3539 2986
rect 3623 2982 3627 2986
rect 3639 2982 3643 2986
rect 3743 2982 3747 2986
rect 3839 2982 3843 2986
rect 3943 2982 3947 2986
rect 111 2934 115 2938
rect 423 2934 427 2938
rect 519 2934 523 2938
rect 615 2934 619 2938
rect 711 2934 715 2938
rect 815 2934 819 2938
rect 935 2934 939 2938
rect 1055 2934 1059 2938
rect 1183 2934 1187 2938
rect 1311 2934 1315 2938
rect 1431 2934 1435 2938
rect 1479 2934 1483 2938
rect 1551 2934 1555 2938
rect 1575 2934 1579 2938
rect 1671 2934 1675 2938
rect 1767 2934 1771 2938
rect 1799 2934 1803 2938
rect 1863 2934 1867 2938
rect 1903 2934 1907 2938
rect 2007 2934 2011 2938
rect 2047 2890 2051 2894
rect 2407 2890 2411 2894
rect 2551 2890 2555 2894
rect 2575 2890 2579 2894
rect 2671 2890 2675 2894
rect 2767 2890 2771 2894
rect 2799 2890 2803 2894
rect 2927 2890 2931 2894
rect 2967 2890 2971 2894
rect 3055 2890 3059 2894
rect 3183 2890 3187 2894
rect 3311 2890 3315 2894
rect 3399 2890 3403 2894
rect 3439 2890 3443 2894
rect 3575 2890 3579 2894
rect 3623 2890 3627 2894
rect 3839 2890 3843 2894
rect 3943 2890 3947 2894
rect 111 2850 115 2854
rect 279 2850 283 2854
rect 447 2850 451 2854
rect 631 2850 635 2854
rect 815 2850 819 2854
rect 999 2850 1003 2854
rect 1183 2850 1187 2854
rect 1359 2850 1363 2854
rect 1479 2850 1483 2854
rect 1527 2850 1531 2854
rect 1575 2850 1579 2854
rect 1671 2850 1675 2854
rect 1695 2850 1699 2854
rect 1767 2850 1771 2854
rect 1863 2850 1867 2854
rect 2007 2850 2011 2854
rect 2047 2814 2051 2818
rect 2439 2814 2443 2818
rect 2551 2814 2555 2818
rect 2567 2814 2571 2818
rect 2671 2814 2675 2818
rect 2695 2814 2699 2818
rect 2799 2814 2803 2818
rect 2831 2814 2835 2818
rect 2927 2814 2931 2818
rect 2967 2814 2971 2818
rect 3055 2814 3059 2818
rect 3103 2814 3107 2818
rect 3183 2814 3187 2818
rect 3247 2814 3251 2818
rect 3311 2814 3315 2818
rect 3391 2814 3395 2818
rect 3439 2814 3443 2818
rect 3543 2814 3547 2818
rect 3575 2814 3579 2818
rect 3703 2814 3707 2818
rect 3839 2814 3843 2818
rect 3943 2814 3947 2818
rect 111 2774 115 2778
rect 239 2774 243 2778
rect 279 2774 283 2778
rect 351 2774 355 2778
rect 447 2774 451 2778
rect 471 2774 475 2778
rect 607 2774 611 2778
rect 631 2774 635 2778
rect 743 2774 747 2778
rect 815 2774 819 2778
rect 879 2774 883 2778
rect 999 2774 1003 2778
rect 1015 2774 1019 2778
rect 1151 2774 1155 2778
rect 1183 2774 1187 2778
rect 1287 2774 1291 2778
rect 1359 2774 1363 2778
rect 1423 2774 1427 2778
rect 1527 2774 1531 2778
rect 1567 2774 1571 2778
rect 1695 2774 1699 2778
rect 1863 2774 1867 2778
rect 2007 2774 2011 2778
rect 2047 2730 2051 2734
rect 2335 2730 2339 2734
rect 2439 2730 2443 2734
rect 2495 2730 2499 2734
rect 2567 2730 2571 2734
rect 2663 2730 2667 2734
rect 2695 2730 2699 2734
rect 2831 2730 2835 2734
rect 2967 2730 2971 2734
rect 2999 2730 3003 2734
rect 3103 2730 3107 2734
rect 3167 2730 3171 2734
rect 3247 2730 3251 2734
rect 3335 2730 3339 2734
rect 3391 2730 3395 2734
rect 3511 2730 3515 2734
rect 3543 2730 3547 2734
rect 3687 2730 3691 2734
rect 3703 2730 3707 2734
rect 3839 2730 3843 2734
rect 3943 2730 3947 2734
rect 111 2698 115 2702
rect 223 2698 227 2702
rect 239 2698 243 2702
rect 351 2698 355 2702
rect 367 2698 371 2702
rect 471 2698 475 2702
rect 503 2698 507 2702
rect 607 2698 611 2702
rect 639 2698 643 2702
rect 743 2698 747 2702
rect 767 2698 771 2702
rect 879 2698 883 2702
rect 887 2698 891 2702
rect 999 2698 1003 2702
rect 1015 2698 1019 2702
rect 1111 2698 1115 2702
rect 1151 2698 1155 2702
rect 1231 2698 1235 2702
rect 1287 2698 1291 2702
rect 1351 2698 1355 2702
rect 1423 2698 1427 2702
rect 1567 2698 1571 2702
rect 2007 2698 2011 2702
rect 2047 2650 2051 2654
rect 2127 2650 2131 2654
rect 2279 2650 2283 2654
rect 2335 2650 2339 2654
rect 2447 2650 2451 2654
rect 2495 2650 2499 2654
rect 2623 2650 2627 2654
rect 2663 2650 2667 2654
rect 2807 2650 2811 2654
rect 2831 2650 2835 2654
rect 2991 2650 2995 2654
rect 2999 2650 3003 2654
rect 3167 2650 3171 2654
rect 3175 2650 3179 2654
rect 3335 2650 3339 2654
rect 3351 2650 3355 2654
rect 3511 2650 3515 2654
rect 3519 2650 3523 2654
rect 3687 2650 3691 2654
rect 3839 2650 3843 2654
rect 3943 2650 3947 2654
rect 111 2622 115 2626
rect 175 2622 179 2626
rect 223 2622 227 2626
rect 367 2622 371 2626
rect 503 2622 507 2626
rect 543 2622 547 2626
rect 639 2622 643 2626
rect 711 2622 715 2626
rect 767 2622 771 2626
rect 863 2622 867 2626
rect 887 2622 891 2626
rect 999 2622 1003 2626
rect 1007 2622 1011 2626
rect 1111 2622 1115 2626
rect 1143 2622 1147 2626
rect 1231 2622 1235 2626
rect 1279 2622 1283 2626
rect 1351 2622 1355 2626
rect 1423 2622 1427 2626
rect 2007 2622 2011 2626
rect 2047 2566 2051 2570
rect 2071 2566 2075 2570
rect 2127 2566 2131 2570
rect 2183 2566 2187 2570
rect 2279 2566 2283 2570
rect 2319 2566 2323 2570
rect 2447 2566 2451 2570
rect 2471 2566 2475 2570
rect 2623 2566 2627 2570
rect 2639 2566 2643 2570
rect 2807 2566 2811 2570
rect 2823 2566 2827 2570
rect 2991 2566 2995 2570
rect 3031 2566 3035 2570
rect 3175 2566 3179 2570
rect 3263 2566 3267 2570
rect 3351 2566 3355 2570
rect 3503 2566 3507 2570
rect 3519 2566 3523 2570
rect 3687 2566 3691 2570
rect 3743 2566 3747 2570
rect 3839 2566 3843 2570
rect 3943 2566 3947 2570
rect 111 2542 115 2546
rect 135 2542 139 2546
rect 175 2542 179 2546
rect 271 2542 275 2546
rect 367 2542 371 2546
rect 439 2542 443 2546
rect 543 2542 547 2546
rect 607 2542 611 2546
rect 711 2542 715 2546
rect 775 2542 779 2546
rect 863 2542 867 2546
rect 927 2542 931 2546
rect 1007 2542 1011 2546
rect 1079 2542 1083 2546
rect 1143 2542 1147 2546
rect 1223 2542 1227 2546
rect 1279 2542 1283 2546
rect 1359 2542 1363 2546
rect 1423 2542 1427 2546
rect 1495 2542 1499 2546
rect 1639 2542 1643 2546
rect 2007 2542 2011 2546
rect 2047 2486 2051 2490
rect 2071 2486 2075 2490
rect 2183 2486 2187 2490
rect 2215 2486 2219 2490
rect 2319 2486 2323 2490
rect 2383 2486 2387 2490
rect 2471 2486 2475 2490
rect 2559 2486 2563 2490
rect 2639 2486 2643 2490
rect 2751 2486 2755 2490
rect 2823 2486 2827 2490
rect 2951 2486 2955 2490
rect 3031 2486 3035 2490
rect 3167 2486 3171 2490
rect 3263 2486 3267 2490
rect 3391 2486 3395 2490
rect 3503 2486 3507 2490
rect 3623 2486 3627 2490
rect 3743 2486 3747 2490
rect 3839 2486 3843 2490
rect 3943 2486 3947 2490
rect 111 2462 115 2466
rect 135 2462 139 2466
rect 271 2462 275 2466
rect 311 2462 315 2466
rect 439 2462 443 2466
rect 511 2462 515 2466
rect 607 2462 611 2466
rect 711 2462 715 2466
rect 775 2462 779 2466
rect 903 2462 907 2466
rect 927 2462 931 2466
rect 1079 2462 1083 2466
rect 1223 2462 1227 2466
rect 1239 2462 1243 2466
rect 1359 2462 1363 2466
rect 1391 2462 1395 2466
rect 1495 2462 1499 2466
rect 1527 2462 1531 2466
rect 1639 2462 1643 2466
rect 1663 2462 1667 2466
rect 1791 2462 1795 2466
rect 1903 2462 1907 2466
rect 2007 2462 2011 2466
rect 2047 2394 2051 2398
rect 2071 2394 2075 2398
rect 2215 2394 2219 2398
rect 2247 2394 2251 2398
rect 2383 2394 2387 2398
rect 2431 2394 2435 2398
rect 2559 2394 2563 2398
rect 2607 2394 2611 2398
rect 2751 2394 2755 2398
rect 2775 2394 2779 2398
rect 2935 2394 2939 2398
rect 2951 2394 2955 2398
rect 3103 2394 3107 2398
rect 3167 2394 3171 2398
rect 3391 2394 3395 2398
rect 3623 2394 3627 2398
rect 3839 2394 3843 2398
rect 3943 2394 3947 2398
rect 111 2386 115 2390
rect 135 2386 139 2390
rect 311 2386 315 2390
rect 327 2386 331 2390
rect 511 2386 515 2390
rect 551 2386 555 2390
rect 711 2386 715 2390
rect 767 2386 771 2390
rect 903 2386 907 2390
rect 975 2386 979 2390
rect 1079 2386 1083 2390
rect 1175 2386 1179 2390
rect 1239 2386 1243 2390
rect 1367 2386 1371 2390
rect 1391 2386 1395 2390
rect 1527 2386 1531 2390
rect 1551 2386 1555 2390
rect 1663 2386 1667 2390
rect 1735 2386 1739 2390
rect 1791 2386 1795 2390
rect 1903 2386 1907 2390
rect 2007 2386 2011 2390
rect 2047 2318 2051 2322
rect 2071 2318 2075 2322
rect 2175 2318 2179 2322
rect 2247 2318 2251 2322
rect 2311 2318 2315 2322
rect 2431 2318 2435 2322
rect 2447 2318 2451 2322
rect 2591 2318 2595 2322
rect 2607 2318 2611 2322
rect 2751 2318 2755 2322
rect 2775 2318 2779 2322
rect 2935 2318 2939 2322
rect 3103 2318 3107 2322
rect 3143 2318 3147 2322
rect 3375 2318 3379 2322
rect 3615 2318 3619 2322
rect 3839 2318 3843 2322
rect 3943 2318 3947 2322
rect 111 2302 115 2306
rect 135 2302 139 2306
rect 271 2302 275 2306
rect 327 2302 331 2306
rect 431 2302 435 2306
rect 551 2302 555 2306
rect 591 2302 595 2306
rect 751 2302 755 2306
rect 767 2302 771 2306
rect 919 2302 923 2306
rect 975 2302 979 2306
rect 1087 2302 1091 2306
rect 1175 2302 1179 2306
rect 1263 2302 1267 2306
rect 1367 2302 1371 2306
rect 1447 2302 1451 2306
rect 1551 2302 1555 2306
rect 1631 2302 1635 2306
rect 1735 2302 1739 2306
rect 1815 2302 1819 2306
rect 1903 2302 1907 2306
rect 2007 2302 2011 2306
rect 2047 2234 2051 2238
rect 2071 2234 2075 2238
rect 2111 2234 2115 2238
rect 2175 2234 2179 2238
rect 2255 2234 2259 2238
rect 2311 2234 2315 2238
rect 2407 2234 2411 2238
rect 2447 2234 2451 2238
rect 2559 2234 2563 2238
rect 2591 2234 2595 2238
rect 2719 2234 2723 2238
rect 2751 2234 2755 2238
rect 2879 2234 2883 2238
rect 2935 2234 2939 2238
rect 3047 2234 3051 2238
rect 3143 2234 3147 2238
rect 3223 2234 3227 2238
rect 3375 2234 3379 2238
rect 3407 2234 3411 2238
rect 3591 2234 3595 2238
rect 3615 2234 3619 2238
rect 3783 2234 3787 2238
rect 3839 2234 3843 2238
rect 3943 2234 3947 2238
rect 111 2226 115 2230
rect 135 2226 139 2230
rect 159 2226 163 2230
rect 271 2226 275 2230
rect 327 2226 331 2230
rect 431 2226 435 2230
rect 495 2226 499 2230
rect 591 2226 595 2230
rect 679 2226 683 2230
rect 751 2226 755 2230
rect 879 2226 883 2230
rect 919 2226 923 2230
rect 1087 2226 1091 2230
rect 1095 2226 1099 2230
rect 1263 2226 1267 2230
rect 1327 2226 1331 2230
rect 1447 2226 1451 2230
rect 1567 2226 1571 2230
rect 1631 2226 1635 2230
rect 1815 2226 1819 2230
rect 2007 2226 2011 2230
rect 111 2150 115 2154
rect 159 2150 163 2154
rect 223 2150 227 2154
rect 327 2150 331 2154
rect 359 2150 363 2154
rect 495 2150 499 2154
rect 639 2150 643 2154
rect 679 2150 683 2154
rect 783 2150 787 2154
rect 879 2150 883 2154
rect 935 2150 939 2154
rect 1095 2150 1099 2154
rect 1263 2150 1267 2154
rect 1327 2150 1331 2154
rect 1447 2150 1451 2154
rect 1567 2150 1571 2154
rect 1631 2150 1635 2154
rect 1815 2150 1819 2154
rect 1823 2150 1827 2154
rect 2007 2150 2011 2154
rect 2047 2146 2051 2150
rect 2111 2146 2115 2150
rect 2255 2146 2259 2150
rect 2287 2146 2291 2150
rect 2407 2146 2411 2150
rect 2431 2146 2435 2150
rect 2559 2146 2563 2150
rect 2583 2146 2587 2150
rect 2719 2146 2723 2150
rect 2735 2146 2739 2150
rect 2879 2146 2883 2150
rect 2887 2146 2891 2150
rect 3047 2146 3051 2150
rect 3207 2146 3211 2150
rect 3223 2146 3227 2150
rect 3367 2146 3371 2150
rect 3407 2146 3411 2150
rect 3527 2146 3531 2150
rect 3591 2146 3595 2150
rect 3695 2146 3699 2150
rect 3783 2146 3787 2150
rect 3839 2146 3843 2150
rect 3943 2146 3947 2150
rect 111 2066 115 2070
rect 223 2066 227 2070
rect 359 2066 363 2070
rect 375 2066 379 2070
rect 495 2066 499 2070
rect 615 2066 619 2070
rect 639 2066 643 2070
rect 751 2066 755 2070
rect 783 2066 787 2070
rect 895 2066 899 2070
rect 935 2066 939 2070
rect 1047 2066 1051 2070
rect 1095 2066 1099 2070
rect 1215 2066 1219 2070
rect 1263 2066 1267 2070
rect 1399 2066 1403 2070
rect 1447 2066 1451 2070
rect 1583 2066 1587 2070
rect 1631 2066 1635 2070
rect 1775 2066 1779 2070
rect 1823 2066 1827 2070
rect 2007 2066 2011 2070
rect 2047 2062 2051 2066
rect 2287 2062 2291 2066
rect 2431 2062 2435 2066
rect 2503 2062 2507 2066
rect 2583 2062 2587 2066
rect 2671 2062 2675 2066
rect 2735 2062 2739 2066
rect 2839 2062 2843 2066
rect 2887 2062 2891 2066
rect 3007 2062 3011 2066
rect 3047 2062 3051 2066
rect 3167 2062 3171 2066
rect 3207 2062 3211 2066
rect 3311 2062 3315 2066
rect 3367 2062 3371 2066
rect 3455 2062 3459 2066
rect 3527 2062 3531 2066
rect 3591 2062 3595 2066
rect 3695 2062 3699 2066
rect 3727 2062 3731 2066
rect 3839 2062 3843 2066
rect 3943 2062 3947 2066
rect 111 1982 115 1986
rect 375 1982 379 1986
rect 495 1982 499 1986
rect 511 1982 515 1986
rect 615 1982 619 1986
rect 623 1982 627 1986
rect 743 1982 747 1986
rect 751 1982 755 1986
rect 871 1982 875 1986
rect 895 1982 899 1986
rect 1007 1982 1011 1986
rect 1047 1982 1051 1986
rect 1143 1982 1147 1986
rect 1215 1982 1219 1986
rect 1279 1982 1283 1986
rect 1399 1982 1403 1986
rect 1415 1982 1419 1986
rect 1559 1982 1563 1986
rect 1583 1982 1587 1986
rect 1703 1982 1707 1986
rect 1775 1982 1779 1986
rect 2007 1982 2011 1986
rect 2047 1982 2051 1986
rect 2495 1982 2499 1986
rect 2503 1982 2507 1986
rect 2591 1982 2595 1986
rect 2671 1982 2675 1986
rect 2695 1982 2699 1986
rect 2807 1982 2811 1986
rect 2839 1982 2843 1986
rect 2927 1982 2931 1986
rect 3007 1982 3011 1986
rect 3047 1982 3051 1986
rect 3167 1982 3171 1986
rect 3175 1982 3179 1986
rect 3295 1982 3299 1986
rect 3311 1982 3315 1986
rect 3415 1982 3419 1986
rect 3455 1982 3459 1986
rect 3543 1982 3547 1986
rect 3591 1982 3595 1986
rect 3671 1982 3675 1986
rect 3727 1982 3731 1986
rect 3799 1982 3803 1986
rect 3839 1982 3843 1986
rect 3943 1982 3947 1986
rect 111 1898 115 1902
rect 511 1898 515 1902
rect 551 1898 555 1902
rect 623 1898 627 1902
rect 663 1898 667 1902
rect 743 1898 747 1902
rect 783 1898 787 1902
rect 871 1898 875 1902
rect 911 1898 915 1902
rect 1007 1898 1011 1902
rect 1047 1898 1051 1902
rect 1143 1898 1147 1902
rect 1175 1898 1179 1902
rect 1279 1898 1283 1902
rect 1311 1898 1315 1902
rect 1415 1898 1419 1902
rect 1447 1898 1451 1902
rect 1559 1898 1563 1902
rect 1583 1898 1587 1902
rect 1703 1898 1707 1902
rect 1719 1898 1723 1902
rect 2007 1898 2011 1902
rect 2047 1902 2051 1906
rect 2071 1902 2075 1906
rect 2247 1902 2251 1906
rect 2439 1902 2443 1906
rect 2495 1902 2499 1906
rect 2591 1902 2595 1906
rect 2623 1902 2627 1906
rect 2695 1902 2699 1906
rect 2791 1902 2795 1906
rect 2807 1902 2811 1906
rect 2927 1902 2931 1906
rect 2959 1902 2963 1906
rect 3047 1902 3051 1906
rect 3127 1902 3131 1906
rect 3175 1902 3179 1906
rect 3295 1902 3299 1906
rect 3303 1902 3307 1906
rect 3415 1902 3419 1906
rect 3487 1902 3491 1906
rect 3543 1902 3547 1906
rect 3671 1902 3675 1906
rect 3799 1902 3803 1906
rect 3839 1902 3843 1906
rect 3943 1902 3947 1906
rect 111 1822 115 1826
rect 503 1822 507 1826
rect 551 1822 555 1826
rect 615 1822 619 1826
rect 663 1822 667 1826
rect 735 1822 739 1826
rect 783 1822 787 1826
rect 863 1822 867 1826
rect 911 1822 915 1826
rect 999 1822 1003 1826
rect 1047 1822 1051 1826
rect 1151 1822 1155 1826
rect 1175 1822 1179 1826
rect 1311 1822 1315 1826
rect 1319 1822 1323 1826
rect 1447 1822 1451 1826
rect 1487 1822 1491 1826
rect 1583 1822 1587 1826
rect 1663 1822 1667 1826
rect 1719 1822 1723 1826
rect 1847 1822 1851 1826
rect 2007 1822 2011 1826
rect 2047 1826 2051 1830
rect 2071 1826 2075 1830
rect 2095 1826 2099 1830
rect 2231 1826 2235 1830
rect 2247 1826 2251 1830
rect 2367 1826 2371 1830
rect 2439 1826 2443 1830
rect 2511 1826 2515 1830
rect 2623 1826 2627 1830
rect 2671 1826 2675 1830
rect 2791 1826 2795 1830
rect 2855 1826 2859 1830
rect 2959 1826 2963 1830
rect 3071 1826 3075 1830
rect 3127 1826 3131 1830
rect 3303 1826 3307 1830
rect 3487 1826 3491 1830
rect 3543 1826 3547 1830
rect 3671 1826 3675 1830
rect 3791 1826 3795 1830
rect 3839 1826 3843 1830
rect 3943 1826 3947 1830
rect 111 1746 115 1750
rect 343 1746 347 1750
rect 463 1746 467 1750
rect 503 1746 507 1750
rect 591 1746 595 1750
rect 615 1746 619 1750
rect 719 1746 723 1750
rect 735 1746 739 1750
rect 847 1746 851 1750
rect 863 1746 867 1750
rect 983 1746 987 1750
rect 999 1746 1003 1750
rect 1127 1746 1131 1750
rect 1151 1746 1155 1750
rect 1279 1746 1283 1750
rect 1319 1746 1323 1750
rect 1439 1746 1443 1750
rect 1487 1746 1491 1750
rect 1599 1746 1603 1750
rect 1663 1746 1667 1750
rect 1847 1746 1851 1750
rect 2007 1746 2011 1750
rect 2047 1750 2051 1754
rect 2095 1750 2099 1754
rect 2183 1750 2187 1754
rect 2231 1750 2235 1754
rect 2287 1750 2291 1754
rect 2367 1750 2371 1754
rect 2391 1750 2395 1754
rect 2495 1750 2499 1754
rect 2511 1750 2515 1754
rect 2599 1750 2603 1754
rect 2671 1750 2675 1754
rect 2703 1750 2707 1754
rect 2807 1750 2811 1754
rect 2855 1750 2859 1754
rect 2911 1750 2915 1754
rect 3015 1750 3019 1754
rect 3071 1750 3075 1754
rect 3127 1750 3131 1754
rect 3303 1750 3307 1754
rect 3543 1750 3547 1754
rect 3791 1750 3795 1754
rect 3943 1750 3947 1754
rect 2047 1674 2051 1678
rect 2183 1674 2187 1678
rect 2231 1674 2235 1678
rect 2287 1674 2291 1678
rect 2367 1674 2371 1678
rect 2391 1674 2395 1678
rect 2495 1674 2499 1678
rect 2519 1674 2523 1678
rect 2599 1674 2603 1678
rect 2679 1674 2683 1678
rect 2703 1674 2707 1678
rect 2807 1674 2811 1678
rect 2847 1674 2851 1678
rect 2911 1674 2915 1678
rect 3015 1674 3019 1678
rect 3023 1674 3027 1678
rect 3127 1674 3131 1678
rect 3191 1674 3195 1678
rect 3359 1674 3363 1678
rect 3527 1674 3531 1678
rect 3695 1674 3699 1678
rect 3839 1674 3843 1678
rect 3943 1674 3947 1678
rect 111 1666 115 1670
rect 159 1666 163 1670
rect 295 1666 299 1670
rect 343 1666 347 1670
rect 455 1666 459 1670
rect 463 1666 467 1670
rect 591 1666 595 1670
rect 623 1666 627 1670
rect 719 1666 723 1670
rect 799 1666 803 1670
rect 847 1666 851 1670
rect 983 1666 987 1670
rect 1127 1666 1131 1670
rect 1167 1666 1171 1670
rect 1279 1666 1283 1670
rect 1351 1666 1355 1670
rect 1439 1666 1443 1670
rect 1543 1666 1547 1670
rect 1599 1666 1603 1670
rect 1735 1666 1739 1670
rect 2007 1666 2011 1670
rect 111 1590 115 1594
rect 135 1590 139 1594
rect 159 1590 163 1594
rect 255 1590 259 1594
rect 295 1590 299 1594
rect 423 1590 427 1594
rect 455 1590 459 1594
rect 607 1590 611 1594
rect 623 1590 627 1594
rect 799 1590 803 1594
rect 983 1590 987 1594
rect 991 1590 995 1594
rect 1167 1590 1171 1594
rect 1183 1590 1187 1594
rect 1351 1590 1355 1594
rect 1367 1590 1371 1594
rect 1543 1590 1547 1594
rect 1551 1590 1555 1594
rect 1735 1590 1739 1594
rect 1903 1590 1907 1594
rect 2007 1590 2011 1594
rect 2047 1590 2051 1594
rect 2071 1590 2075 1594
rect 2231 1590 2235 1594
rect 2271 1590 2275 1594
rect 2367 1590 2371 1594
rect 2495 1590 2499 1594
rect 2519 1590 2523 1594
rect 2679 1590 2683 1594
rect 2711 1590 2715 1594
rect 2847 1590 2851 1594
rect 2911 1590 2915 1594
rect 3023 1590 3027 1594
rect 3095 1590 3099 1594
rect 3191 1590 3195 1594
rect 3263 1590 3267 1594
rect 3359 1590 3363 1594
rect 3423 1590 3427 1594
rect 3527 1590 3531 1594
rect 3567 1590 3571 1594
rect 3695 1590 3699 1594
rect 3711 1590 3715 1594
rect 3839 1590 3843 1594
rect 3943 1590 3947 1594
rect 111 1510 115 1514
rect 135 1510 139 1514
rect 247 1510 251 1514
rect 255 1510 259 1514
rect 399 1510 403 1514
rect 423 1510 427 1514
rect 559 1510 563 1514
rect 607 1510 611 1514
rect 719 1510 723 1514
rect 799 1510 803 1514
rect 879 1510 883 1514
rect 991 1510 995 1514
rect 1039 1510 1043 1514
rect 1183 1510 1187 1514
rect 1319 1510 1323 1514
rect 1367 1510 1371 1514
rect 1447 1510 1451 1514
rect 1551 1510 1555 1514
rect 1567 1510 1571 1514
rect 1687 1510 1691 1514
rect 1735 1510 1739 1514
rect 1807 1510 1811 1514
rect 1903 1510 1907 1514
rect 2007 1510 2011 1514
rect 2047 1514 2051 1518
rect 2071 1514 2075 1518
rect 2271 1514 2275 1518
rect 2431 1514 2435 1518
rect 2495 1514 2499 1518
rect 2711 1514 2715 1518
rect 2791 1514 2795 1518
rect 2911 1514 2915 1518
rect 3095 1514 3099 1518
rect 3127 1514 3131 1518
rect 3263 1514 3267 1518
rect 3423 1514 3427 1518
rect 3463 1514 3467 1518
rect 3567 1514 3571 1518
rect 3711 1514 3715 1518
rect 3799 1514 3803 1518
rect 3839 1514 3843 1518
rect 3943 1514 3947 1518
rect 111 1434 115 1438
rect 135 1434 139 1438
rect 247 1434 251 1438
rect 263 1434 267 1438
rect 399 1434 403 1438
rect 431 1434 435 1438
rect 559 1434 563 1438
rect 607 1434 611 1438
rect 719 1434 723 1438
rect 791 1434 795 1438
rect 879 1434 883 1438
rect 975 1434 979 1438
rect 1039 1434 1043 1438
rect 1159 1434 1163 1438
rect 1183 1434 1187 1438
rect 1319 1434 1323 1438
rect 1351 1434 1355 1438
rect 1447 1434 1451 1438
rect 1543 1434 1547 1438
rect 1567 1434 1571 1438
rect 1687 1434 1691 1438
rect 1735 1434 1739 1438
rect 1807 1434 1811 1438
rect 1903 1434 1907 1438
rect 2007 1434 2011 1438
rect 2047 1430 2051 1434
rect 2071 1430 2075 1434
rect 2271 1430 2275 1434
rect 2431 1430 2435 1434
rect 2495 1430 2499 1434
rect 2711 1430 2715 1434
rect 2791 1430 2795 1434
rect 2911 1430 2915 1434
rect 3095 1430 3099 1434
rect 3127 1430 3131 1434
rect 3271 1430 3275 1434
rect 3439 1430 3443 1434
rect 3463 1430 3467 1434
rect 3607 1430 3611 1434
rect 3783 1430 3787 1434
rect 3799 1430 3803 1434
rect 3943 1430 3947 1434
rect 111 1354 115 1358
rect 135 1354 139 1358
rect 159 1354 163 1358
rect 263 1354 267 1358
rect 311 1354 315 1358
rect 431 1354 435 1358
rect 479 1354 483 1358
rect 607 1354 611 1358
rect 663 1354 667 1358
rect 791 1354 795 1358
rect 855 1354 859 1358
rect 975 1354 979 1358
rect 1047 1354 1051 1358
rect 1159 1354 1163 1358
rect 1247 1354 1251 1358
rect 1351 1354 1355 1358
rect 1447 1354 1451 1358
rect 1543 1354 1547 1358
rect 1655 1354 1659 1358
rect 1735 1354 1739 1358
rect 1863 1354 1867 1358
rect 1903 1354 1907 1358
rect 2007 1354 2011 1358
rect 2047 1354 2051 1358
rect 2071 1354 2075 1358
rect 2207 1354 2211 1358
rect 2271 1354 2275 1358
rect 2383 1354 2387 1358
rect 2495 1354 2499 1358
rect 2567 1354 2571 1358
rect 2711 1354 2715 1358
rect 2751 1354 2755 1358
rect 2911 1354 2915 1358
rect 2935 1354 2939 1358
rect 3095 1354 3099 1358
rect 3111 1354 3115 1358
rect 3271 1354 3275 1358
rect 3279 1354 3283 1358
rect 3439 1354 3443 1358
rect 3447 1354 3451 1358
rect 3607 1354 3611 1358
rect 3623 1354 3627 1358
rect 3783 1354 3787 1358
rect 3943 1354 3947 1358
rect 111 1274 115 1278
rect 159 1274 163 1278
rect 311 1274 315 1278
rect 407 1274 411 1278
rect 479 1274 483 1278
rect 543 1274 547 1278
rect 663 1274 667 1278
rect 695 1274 699 1278
rect 855 1274 859 1278
rect 1023 1274 1027 1278
rect 1047 1274 1051 1278
rect 1191 1274 1195 1278
rect 1247 1274 1251 1278
rect 1367 1274 1371 1278
rect 1447 1274 1451 1278
rect 1543 1274 1547 1278
rect 1655 1274 1659 1278
rect 1719 1274 1723 1278
rect 1863 1274 1867 1278
rect 1895 1274 1899 1278
rect 2007 1274 2011 1278
rect 2047 1278 2051 1282
rect 2071 1278 2075 1282
rect 2151 1278 2155 1282
rect 2207 1278 2211 1282
rect 2287 1278 2291 1282
rect 2383 1278 2387 1282
rect 2431 1278 2435 1282
rect 2567 1278 2571 1282
rect 2583 1278 2587 1282
rect 2743 1278 2747 1282
rect 2751 1278 2755 1282
rect 2903 1278 2907 1282
rect 2935 1278 2939 1282
rect 3071 1278 3075 1282
rect 3111 1278 3115 1282
rect 3247 1278 3251 1282
rect 3279 1278 3283 1282
rect 3431 1278 3435 1282
rect 3447 1278 3451 1282
rect 3615 1278 3619 1282
rect 3623 1278 3627 1282
rect 3807 1278 3811 1282
rect 3943 1278 3947 1282
rect 111 1198 115 1202
rect 407 1198 411 1202
rect 423 1198 427 1202
rect 543 1198 547 1202
rect 591 1198 595 1202
rect 695 1198 699 1202
rect 759 1198 763 1202
rect 855 1198 859 1202
rect 927 1198 931 1202
rect 1023 1198 1027 1202
rect 1095 1198 1099 1202
rect 1191 1198 1195 1202
rect 1247 1198 1251 1202
rect 1367 1198 1371 1202
rect 1399 1198 1403 1202
rect 1543 1198 1547 1202
rect 1687 1198 1691 1202
rect 1719 1198 1723 1202
rect 1839 1198 1843 1202
rect 1895 1198 1899 1202
rect 2007 1198 2011 1202
rect 2047 1202 2051 1206
rect 2151 1202 2155 1206
rect 2287 1202 2291 1206
rect 2311 1202 2315 1206
rect 2415 1202 2419 1206
rect 2431 1202 2435 1206
rect 2527 1202 2531 1206
rect 2583 1202 2587 1206
rect 2639 1202 2643 1206
rect 2743 1202 2747 1206
rect 2767 1202 2771 1206
rect 2903 1202 2907 1206
rect 2911 1202 2915 1206
rect 3071 1202 3075 1206
rect 3247 1202 3251 1206
rect 3431 1202 3435 1206
rect 3439 1202 3443 1206
rect 3615 1202 3619 1206
rect 3631 1202 3635 1206
rect 3807 1202 3811 1206
rect 3831 1202 3835 1206
rect 3943 1202 3947 1206
rect 111 1118 115 1122
rect 375 1118 379 1122
rect 423 1118 427 1122
rect 487 1118 491 1122
rect 591 1118 595 1122
rect 599 1118 603 1122
rect 711 1118 715 1122
rect 759 1118 763 1122
rect 831 1118 835 1122
rect 927 1118 931 1122
rect 967 1118 971 1122
rect 1095 1118 1099 1122
rect 1119 1118 1123 1122
rect 1247 1118 1251 1122
rect 1279 1118 1283 1122
rect 1399 1118 1403 1122
rect 1447 1118 1451 1122
rect 1543 1118 1547 1122
rect 1623 1118 1627 1122
rect 1687 1118 1691 1122
rect 1839 1118 1843 1122
rect 2007 1118 2011 1122
rect 2047 1122 2051 1126
rect 2311 1122 2315 1126
rect 2407 1122 2411 1126
rect 2415 1122 2419 1126
rect 2503 1122 2507 1126
rect 2527 1122 2531 1126
rect 2599 1122 2603 1126
rect 2639 1122 2643 1126
rect 2695 1122 2699 1126
rect 2767 1122 2771 1126
rect 2807 1122 2811 1126
rect 2911 1122 2915 1126
rect 2943 1122 2947 1126
rect 3071 1122 3075 1126
rect 3095 1122 3099 1126
rect 3247 1122 3251 1126
rect 3263 1122 3267 1126
rect 3439 1122 3443 1126
rect 3447 1122 3451 1126
rect 3631 1122 3635 1126
rect 3639 1122 3643 1126
rect 3831 1122 3835 1126
rect 3839 1122 3843 1126
rect 3943 1122 3947 1126
rect 111 1042 115 1046
rect 303 1042 307 1046
rect 375 1042 379 1046
rect 447 1042 451 1046
rect 487 1042 491 1046
rect 591 1042 595 1046
rect 599 1042 603 1046
rect 711 1042 715 1046
rect 727 1042 731 1046
rect 831 1042 835 1046
rect 855 1042 859 1046
rect 967 1042 971 1046
rect 975 1042 979 1046
rect 1087 1042 1091 1046
rect 1119 1042 1123 1046
rect 1199 1042 1203 1046
rect 1279 1042 1283 1046
rect 1311 1042 1315 1046
rect 1431 1042 1435 1046
rect 1447 1042 1451 1046
rect 1623 1042 1627 1046
rect 2007 1042 2011 1046
rect 2047 1042 2051 1046
rect 2407 1042 2411 1046
rect 2455 1042 2459 1046
rect 2503 1042 2507 1046
rect 2551 1042 2555 1046
rect 2599 1042 2603 1046
rect 2647 1042 2651 1046
rect 2695 1042 2699 1046
rect 2759 1042 2763 1046
rect 2807 1042 2811 1046
rect 2887 1042 2891 1046
rect 2943 1042 2947 1046
rect 3031 1042 3035 1046
rect 3095 1042 3099 1046
rect 3183 1042 3187 1046
rect 3263 1042 3267 1046
rect 3343 1042 3347 1046
rect 3447 1042 3451 1046
rect 3503 1042 3507 1046
rect 3639 1042 3643 1046
rect 3671 1042 3675 1046
rect 3839 1042 3843 1046
rect 3943 1042 3947 1046
rect 111 966 115 970
rect 255 966 259 970
rect 303 966 307 970
rect 447 966 451 970
rect 591 966 595 970
rect 631 966 635 970
rect 727 966 731 970
rect 807 966 811 970
rect 855 966 859 970
rect 975 966 979 970
rect 1087 966 1091 970
rect 1127 966 1131 970
rect 1199 966 1203 970
rect 1271 966 1275 970
rect 1311 966 1315 970
rect 1415 966 1419 970
rect 1431 966 1435 970
rect 1551 966 1555 970
rect 1695 966 1699 970
rect 2007 966 2011 970
rect 2047 962 2051 966
rect 2423 962 2427 966
rect 2455 962 2459 966
rect 2519 962 2523 966
rect 2551 962 2555 966
rect 2615 962 2619 966
rect 2647 962 2651 966
rect 2711 962 2715 966
rect 2759 962 2763 966
rect 2823 962 2827 966
rect 2887 962 2891 966
rect 2951 962 2955 966
rect 3031 962 3035 966
rect 3103 962 3107 966
rect 3183 962 3187 966
rect 3271 962 3275 966
rect 3343 962 3347 966
rect 3455 962 3459 966
rect 3503 962 3507 966
rect 3647 962 3651 966
rect 3671 962 3675 966
rect 3839 962 3843 966
rect 3943 962 3947 966
rect 111 886 115 890
rect 255 886 259 890
rect 447 886 451 890
rect 631 886 635 890
rect 639 886 643 890
rect 807 886 811 890
rect 823 886 827 890
rect 975 886 979 890
rect 999 886 1003 890
rect 1127 886 1131 890
rect 1167 886 1171 890
rect 1271 886 1275 890
rect 1327 886 1331 890
rect 1415 886 1419 890
rect 1479 886 1483 890
rect 1551 886 1555 890
rect 1631 886 1635 890
rect 1695 886 1699 890
rect 1783 886 1787 890
rect 2007 886 2011 890
rect 2047 886 2051 890
rect 2343 886 2347 890
rect 2423 886 2427 890
rect 2439 886 2443 890
rect 2519 886 2523 890
rect 2535 886 2539 890
rect 2615 886 2619 890
rect 2631 886 2635 890
rect 2711 886 2715 890
rect 2735 886 2739 890
rect 2823 886 2827 890
rect 2863 886 2867 890
rect 2951 886 2955 890
rect 3015 886 3019 890
rect 3103 886 3107 890
rect 3191 886 3195 890
rect 3271 886 3275 890
rect 3391 886 3395 890
rect 3455 886 3459 890
rect 3607 886 3611 890
rect 3647 886 3651 890
rect 3823 886 3827 890
rect 3839 886 3843 890
rect 3943 886 3947 890
rect 111 806 115 810
rect 159 806 163 810
rect 255 806 259 810
rect 311 806 315 810
rect 447 806 451 810
rect 471 806 475 810
rect 623 806 627 810
rect 639 806 643 810
rect 775 806 779 810
rect 823 806 827 810
rect 935 806 939 810
rect 999 806 1003 810
rect 1095 806 1099 810
rect 1167 806 1171 810
rect 1255 806 1259 810
rect 1327 806 1331 810
rect 1415 806 1419 810
rect 1479 806 1483 810
rect 1583 806 1587 810
rect 1631 806 1635 810
rect 1751 806 1755 810
rect 1783 806 1787 810
rect 1903 806 1907 810
rect 2007 806 2011 810
rect 2047 810 2051 814
rect 2311 810 2315 814
rect 2343 810 2347 814
rect 2439 810 2443 814
rect 2495 810 2499 814
rect 2535 810 2539 814
rect 2631 810 2635 814
rect 2687 810 2691 814
rect 2735 810 2739 814
rect 2863 810 2867 814
rect 2879 810 2883 814
rect 3015 810 3019 814
rect 3079 810 3083 814
rect 3191 810 3195 814
rect 3287 810 3291 814
rect 3391 810 3395 814
rect 3503 810 3507 814
rect 3607 810 3611 814
rect 3719 810 3723 814
rect 3823 810 3827 814
rect 3943 810 3947 814
rect 111 730 115 734
rect 135 730 139 734
rect 159 730 163 734
rect 263 730 267 734
rect 311 730 315 734
rect 431 730 435 734
rect 471 730 475 734
rect 623 730 627 734
rect 775 730 779 734
rect 823 730 827 734
rect 935 730 939 734
rect 1015 730 1019 734
rect 1095 730 1099 734
rect 1207 730 1211 734
rect 1255 730 1259 734
rect 1391 730 1395 734
rect 1415 730 1419 734
rect 1567 730 1571 734
rect 1583 730 1587 734
rect 1743 730 1747 734
rect 1751 730 1755 734
rect 1903 730 1907 734
rect 2007 730 2011 734
rect 2047 730 2051 734
rect 2071 730 2075 734
rect 2255 730 2259 734
rect 2311 730 2315 734
rect 2455 730 2459 734
rect 2495 730 2499 734
rect 2655 730 2659 734
rect 2687 730 2691 734
rect 2855 730 2859 734
rect 2879 730 2883 734
rect 3047 730 3051 734
rect 3079 730 3083 734
rect 3239 730 3243 734
rect 3287 730 3291 734
rect 3439 730 3443 734
rect 3503 730 3507 734
rect 3639 730 3643 734
rect 3719 730 3723 734
rect 3839 730 3843 734
rect 3943 730 3947 734
rect 111 654 115 658
rect 135 654 139 658
rect 247 654 251 658
rect 263 654 267 658
rect 383 654 387 658
rect 431 654 435 658
rect 527 654 531 658
rect 623 654 627 658
rect 687 654 691 658
rect 823 654 827 658
rect 871 654 875 658
rect 1015 654 1019 658
rect 1079 654 1083 658
rect 1207 654 1211 658
rect 1303 654 1307 658
rect 1391 654 1395 658
rect 1543 654 1547 658
rect 1567 654 1571 658
rect 1743 654 1747 658
rect 1783 654 1787 658
rect 1903 654 1907 658
rect 2007 654 2011 658
rect 2047 654 2051 658
rect 2071 654 2075 658
rect 2231 654 2235 658
rect 2255 654 2259 658
rect 2431 654 2435 658
rect 2455 654 2459 658
rect 2631 654 2635 658
rect 2655 654 2659 658
rect 2831 654 2835 658
rect 2855 654 2859 658
rect 3023 654 3027 658
rect 3047 654 3051 658
rect 3207 654 3211 658
rect 3239 654 3243 658
rect 3375 654 3379 658
rect 3439 654 3443 658
rect 3535 654 3539 658
rect 3639 654 3643 658
rect 3695 654 3699 658
rect 3839 654 3843 658
rect 3943 654 3947 658
rect 111 574 115 578
rect 135 574 139 578
rect 247 574 251 578
rect 295 574 299 578
rect 383 574 387 578
rect 479 574 483 578
rect 527 574 531 578
rect 663 574 667 578
rect 687 574 691 578
rect 847 574 851 578
rect 871 574 875 578
rect 1031 574 1035 578
rect 1079 574 1083 578
rect 1215 574 1219 578
rect 1303 574 1307 578
rect 1399 574 1403 578
rect 1543 574 1547 578
rect 1591 574 1595 578
rect 1783 574 1787 578
rect 2007 574 2011 578
rect 2047 574 2051 578
rect 2071 574 2075 578
rect 2215 574 2219 578
rect 2231 574 2235 578
rect 2399 574 2403 578
rect 2431 574 2435 578
rect 2583 574 2587 578
rect 2631 574 2635 578
rect 2775 574 2779 578
rect 2831 574 2835 578
rect 2959 574 2963 578
rect 3023 574 3027 578
rect 3143 574 3147 578
rect 3207 574 3211 578
rect 3319 574 3323 578
rect 3375 574 3379 578
rect 3495 574 3499 578
rect 3535 574 3539 578
rect 3679 574 3683 578
rect 3695 574 3699 578
rect 3839 574 3843 578
rect 3943 574 3947 578
rect 111 498 115 502
rect 135 498 139 502
rect 287 498 291 502
rect 295 498 299 502
rect 455 498 459 502
rect 479 498 483 502
rect 615 498 619 502
rect 663 498 667 502
rect 767 498 771 502
rect 847 498 851 502
rect 903 498 907 502
rect 1031 498 1035 502
rect 1159 498 1163 502
rect 1215 498 1219 502
rect 1287 498 1291 502
rect 1399 498 1403 502
rect 1415 498 1419 502
rect 1591 498 1595 502
rect 1783 498 1787 502
rect 2007 498 2011 502
rect 2047 494 2051 498
rect 2071 494 2075 498
rect 2215 494 2219 498
rect 2223 494 2227 498
rect 2391 494 2395 498
rect 2399 494 2403 498
rect 2559 494 2563 498
rect 2583 494 2587 498
rect 2727 494 2731 498
rect 2775 494 2779 498
rect 2895 494 2899 498
rect 2959 494 2963 498
rect 3063 494 3067 498
rect 3143 494 3147 498
rect 3223 494 3227 498
rect 3319 494 3323 498
rect 3383 494 3387 498
rect 3495 494 3499 498
rect 3543 494 3547 498
rect 3679 494 3683 498
rect 3703 494 3707 498
rect 3839 494 3843 498
rect 3943 494 3947 498
rect 111 422 115 426
rect 135 422 139 426
rect 287 422 291 426
rect 447 422 451 426
rect 455 422 459 426
rect 599 422 603 426
rect 615 422 619 426
rect 751 422 755 426
rect 767 422 771 426
rect 903 422 907 426
rect 1031 422 1035 426
rect 1079 422 1083 426
rect 1159 422 1163 426
rect 1271 422 1275 426
rect 1287 422 1291 426
rect 1415 422 1419 426
rect 1479 422 1483 426
rect 1703 422 1707 426
rect 1903 422 1907 426
rect 2007 422 2011 426
rect 2047 418 2051 422
rect 2071 418 2075 422
rect 2223 418 2227 422
rect 2391 418 2395 422
rect 2463 418 2467 422
rect 2559 418 2563 422
rect 2655 418 2659 422
rect 2727 418 2731 422
rect 2751 418 2755 422
rect 2847 418 2851 422
rect 2895 418 2899 422
rect 2943 418 2947 422
rect 3039 418 3043 422
rect 3063 418 3067 422
rect 3135 418 3139 422
rect 3223 418 3227 422
rect 3231 418 3235 422
rect 3383 418 3387 422
rect 3543 418 3547 422
rect 3703 418 3707 422
rect 3839 418 3843 422
rect 3943 418 3947 422
rect 111 342 115 346
rect 135 342 139 346
rect 159 342 163 346
rect 287 342 291 346
rect 351 342 355 346
rect 447 342 451 346
rect 551 342 555 346
rect 599 342 603 346
rect 751 342 755 346
rect 759 342 763 346
rect 903 342 907 346
rect 959 342 963 346
rect 1079 342 1083 346
rect 1159 342 1163 346
rect 1271 342 1275 346
rect 1343 342 1347 346
rect 1479 342 1483 346
rect 1527 342 1531 346
rect 1703 342 1707 346
rect 1711 342 1715 346
rect 1895 342 1899 346
rect 1903 342 1907 346
rect 2007 342 2011 346
rect 2047 342 2051 346
rect 2399 342 2403 346
rect 2463 342 2467 346
rect 2503 342 2507 346
rect 2559 342 2563 346
rect 2623 342 2627 346
rect 2655 342 2659 346
rect 2751 342 2755 346
rect 2759 342 2763 346
rect 2847 342 2851 346
rect 2911 342 2915 346
rect 2943 342 2947 346
rect 3039 342 3043 346
rect 3071 342 3075 346
rect 3135 342 3139 346
rect 3231 342 3235 346
rect 3247 342 3251 346
rect 3423 342 3427 346
rect 3607 342 3611 346
rect 3791 342 3795 346
rect 3943 342 3947 346
rect 2047 266 2051 270
rect 2191 266 2195 270
rect 2351 266 2355 270
rect 2399 266 2403 270
rect 2503 266 2507 270
rect 2519 266 2523 270
rect 2623 266 2627 270
rect 2687 266 2691 270
rect 2759 266 2763 270
rect 2855 266 2859 270
rect 2911 266 2915 270
rect 3031 266 3035 270
rect 3071 266 3075 270
rect 3215 266 3219 270
rect 3247 266 3251 270
rect 3407 266 3411 270
rect 3423 266 3427 270
rect 3607 266 3611 270
rect 3791 266 3795 270
rect 3807 266 3811 270
rect 3943 266 3947 270
rect 111 258 115 262
rect 159 258 163 262
rect 223 258 227 262
rect 351 258 355 262
rect 383 258 387 262
rect 543 258 547 262
rect 551 258 555 262
rect 703 258 707 262
rect 759 258 763 262
rect 863 258 867 262
rect 959 258 963 262
rect 1031 258 1035 262
rect 1159 258 1163 262
rect 1199 258 1203 262
rect 1343 258 1347 262
rect 1367 258 1371 262
rect 1527 258 1531 262
rect 1543 258 1547 262
rect 1711 258 1715 262
rect 1727 258 1731 262
rect 1895 258 1899 262
rect 1903 258 1907 262
rect 2007 258 2011 262
rect 111 162 115 166
rect 135 162 139 166
rect 223 162 227 166
rect 231 162 235 166
rect 327 162 331 166
rect 383 162 387 166
rect 423 162 427 166
rect 527 162 531 166
rect 543 162 547 166
rect 647 162 651 166
rect 703 162 707 166
rect 775 162 779 166
rect 863 162 867 166
rect 903 162 907 166
rect 1031 162 1035 166
rect 1151 162 1155 166
rect 1199 162 1203 166
rect 1271 162 1275 166
rect 1367 162 1371 166
rect 1383 162 1387 166
rect 1487 162 1491 166
rect 1543 162 1547 166
rect 1591 162 1595 166
rect 1703 162 1707 166
rect 1727 162 1731 166
rect 1807 162 1811 166
rect 1903 162 1907 166
rect 2007 162 2011 166
rect 2047 158 2051 162
rect 2071 158 2075 162
rect 2167 158 2171 162
rect 2191 158 2195 162
rect 2263 158 2267 162
rect 2351 158 2355 162
rect 2367 158 2371 162
rect 2487 158 2491 162
rect 2519 158 2523 162
rect 2615 158 2619 162
rect 2687 158 2691 162
rect 2743 158 2747 162
rect 2855 158 2859 162
rect 2871 158 2875 162
rect 2991 158 2995 162
rect 3031 158 3035 162
rect 3111 158 3115 162
rect 3215 158 3219 162
rect 3223 158 3227 162
rect 3327 158 3331 162
rect 3407 158 3411 162
rect 3431 158 3435 162
rect 3535 158 3539 162
rect 3607 158 3611 162
rect 3639 158 3643 162
rect 3743 158 3747 162
rect 3807 158 3811 162
rect 3839 158 3843 162
rect 3943 158 3947 162
rect 111 86 115 90
rect 135 86 139 90
rect 231 86 235 90
rect 327 86 331 90
rect 423 86 427 90
rect 527 86 531 90
rect 647 86 651 90
rect 775 86 779 90
rect 903 86 907 90
rect 1031 86 1035 90
rect 1151 86 1155 90
rect 1271 86 1275 90
rect 1383 86 1387 90
rect 1487 86 1491 90
rect 1591 86 1595 90
rect 1703 86 1707 90
rect 1807 86 1811 90
rect 1903 86 1907 90
rect 2007 86 2011 90
rect 2047 82 2051 86
rect 2071 82 2075 86
rect 2167 82 2171 86
rect 2263 82 2267 86
rect 2367 82 2371 86
rect 2487 82 2491 86
rect 2615 82 2619 86
rect 2743 82 2747 86
rect 2871 82 2875 86
rect 2991 82 2995 86
rect 3111 82 3115 86
rect 3223 82 3227 86
rect 3327 82 3331 86
rect 3431 82 3435 86
rect 3535 82 3539 86
rect 3639 82 3643 86
rect 3743 82 3747 86
rect 3839 82 3843 86
rect 3943 82 3947 86
<< m4 >>
rect 2030 4025 2031 4031
rect 2037 4030 3979 4031
rect 2037 4026 2047 4030
rect 2051 4026 2071 4030
rect 2075 4026 3943 4030
rect 3947 4026 3979 4030
rect 2037 4025 3979 4026
rect 3985 4025 3986 4031
rect 96 4005 97 4011
rect 103 4010 2031 4011
rect 103 4006 111 4010
rect 115 4006 151 4010
rect 155 4006 279 4010
rect 283 4006 431 4010
rect 435 4006 607 4010
rect 611 4006 791 4010
rect 795 4006 975 4010
rect 979 4006 1151 4010
rect 1155 4006 1311 4010
rect 1315 4006 1471 4010
rect 1475 4006 1623 4010
rect 1627 4006 1775 4010
rect 1779 4006 1903 4010
rect 1907 4006 2007 4010
rect 2011 4006 2031 4010
rect 103 4005 2031 4006
rect 2037 4005 2038 4011
rect 2018 3949 2019 3955
rect 2025 3954 3967 3955
rect 2025 3950 2047 3954
rect 2051 3950 2071 3954
rect 2075 3950 2079 3954
rect 2083 3950 2215 3954
rect 2219 3950 2359 3954
rect 2363 3950 2503 3954
rect 2507 3950 2647 3954
rect 2651 3950 2791 3954
rect 2795 3950 2927 3954
rect 2931 3950 3055 3954
rect 3059 3950 3175 3954
rect 3179 3950 3295 3954
rect 3299 3950 3415 3954
rect 3419 3950 3535 3954
rect 3539 3950 3943 3954
rect 3947 3950 3967 3954
rect 2025 3949 3967 3950
rect 3973 3949 3974 3955
rect 84 3929 85 3935
rect 91 3934 2019 3935
rect 91 3930 111 3934
rect 115 3930 151 3934
rect 155 3930 279 3934
rect 283 3930 303 3934
rect 307 3930 423 3934
rect 427 3930 431 3934
rect 435 3930 551 3934
rect 555 3930 607 3934
rect 611 3930 687 3934
rect 691 3930 791 3934
rect 795 3930 815 3934
rect 819 3930 943 3934
rect 947 3930 975 3934
rect 979 3930 1071 3934
rect 1075 3930 1151 3934
rect 1155 3930 1199 3934
rect 1203 3930 1311 3934
rect 1315 3930 1327 3934
rect 1331 3930 1463 3934
rect 1467 3930 1471 3934
rect 1475 3930 1623 3934
rect 1627 3930 1775 3934
rect 1779 3930 1903 3934
rect 1907 3930 2007 3934
rect 2011 3930 2019 3934
rect 91 3929 2019 3930
rect 2025 3929 2026 3935
rect 2030 3873 2031 3879
rect 2037 3878 3979 3879
rect 2037 3874 2047 3878
rect 2051 3874 2079 3878
rect 2083 3874 2215 3878
rect 2219 3874 2255 3878
rect 2259 3874 2359 3878
rect 2363 3874 2383 3878
rect 2387 3874 2503 3878
rect 2507 3874 2519 3878
rect 2523 3874 2647 3878
rect 2651 3874 2671 3878
rect 2675 3874 2791 3878
rect 2795 3874 2831 3878
rect 2835 3874 2927 3878
rect 2931 3874 2991 3878
rect 2995 3874 3055 3878
rect 3059 3874 3159 3878
rect 3163 3874 3175 3878
rect 3179 3874 3295 3878
rect 3299 3874 3327 3878
rect 3331 3874 3415 3878
rect 3419 3874 3495 3878
rect 3499 3874 3535 3878
rect 3539 3874 3663 3878
rect 3667 3874 3943 3878
rect 3947 3874 3979 3878
rect 2037 3873 3979 3874
rect 3985 3873 3986 3879
rect 96 3849 97 3855
rect 103 3854 2031 3855
rect 103 3850 111 3854
rect 115 3850 303 3854
rect 307 3850 415 3854
rect 419 3850 423 3854
rect 427 3850 551 3854
rect 555 3850 567 3854
rect 571 3850 687 3854
rect 691 3850 727 3854
rect 731 3850 815 3854
rect 819 3850 887 3854
rect 891 3850 943 3854
rect 947 3850 1039 3854
rect 1043 3850 1071 3854
rect 1075 3850 1191 3854
rect 1195 3850 1199 3854
rect 1203 3850 1327 3854
rect 1331 3850 1343 3854
rect 1347 3850 1463 3854
rect 1467 3850 1495 3854
rect 1499 3850 1647 3854
rect 1651 3850 2007 3854
rect 2011 3850 2031 3854
rect 103 3849 2031 3850
rect 2037 3849 2038 3855
rect 2018 3797 2019 3803
rect 2025 3802 3967 3803
rect 2025 3798 2047 3802
rect 2051 3798 2071 3802
rect 2075 3798 2199 3802
rect 2203 3798 2255 3802
rect 2259 3798 2375 3802
rect 2379 3798 2383 3802
rect 2387 3798 2519 3802
rect 2523 3798 2559 3802
rect 2563 3798 2671 3802
rect 2675 3798 2751 3802
rect 2755 3798 2831 3802
rect 2835 3798 2951 3802
rect 2955 3798 2991 3802
rect 2995 3798 3143 3802
rect 3147 3798 3159 3802
rect 3163 3798 3327 3802
rect 3331 3798 3335 3802
rect 3339 3798 3495 3802
rect 3499 3798 3535 3802
rect 3539 3798 3663 3802
rect 3667 3798 3735 3802
rect 3739 3798 3943 3802
rect 3947 3798 3967 3802
rect 2025 3797 3967 3798
rect 3973 3797 3974 3803
rect 84 3769 85 3775
rect 91 3774 2019 3775
rect 91 3770 111 3774
rect 115 3770 399 3774
rect 403 3770 415 3774
rect 419 3770 567 3774
rect 571 3770 727 3774
rect 731 3770 751 3774
rect 755 3770 887 3774
rect 891 3770 935 3774
rect 939 3770 1039 3774
rect 1043 3770 1127 3774
rect 1131 3770 1191 3774
rect 1195 3770 1311 3774
rect 1315 3770 1343 3774
rect 1347 3770 1495 3774
rect 1499 3770 1503 3774
rect 1507 3770 1647 3774
rect 1651 3770 1695 3774
rect 1699 3770 1887 3774
rect 1891 3770 2007 3774
rect 2011 3770 2019 3774
rect 91 3769 2019 3770
rect 2025 3769 2026 3775
rect 2030 3709 2031 3715
rect 2037 3714 3979 3715
rect 2037 3710 2047 3714
rect 2051 3710 2071 3714
rect 2075 3710 2199 3714
rect 2203 3710 2263 3714
rect 2267 3710 2375 3714
rect 2379 3710 2479 3714
rect 2483 3710 2559 3714
rect 2563 3710 2695 3714
rect 2699 3710 2751 3714
rect 2755 3710 2911 3714
rect 2915 3710 2951 3714
rect 2955 3710 3119 3714
rect 3123 3710 3143 3714
rect 3147 3710 3319 3714
rect 3323 3710 3335 3714
rect 3339 3710 3519 3714
rect 3523 3710 3535 3714
rect 3539 3710 3727 3714
rect 3731 3710 3735 3714
rect 3739 3710 3943 3714
rect 3947 3710 3979 3714
rect 2037 3709 3979 3710
rect 3985 3709 3986 3715
rect 96 3681 97 3687
rect 103 3686 2031 3687
rect 103 3682 111 3686
rect 115 3682 367 3686
rect 371 3682 399 3686
rect 403 3682 519 3686
rect 523 3682 567 3686
rect 571 3682 679 3686
rect 683 3682 751 3686
rect 755 3682 847 3686
rect 851 3682 935 3686
rect 939 3682 1015 3686
rect 1019 3682 1127 3686
rect 1131 3682 1175 3686
rect 1179 3682 1311 3686
rect 1315 3682 1327 3686
rect 1331 3682 1479 3686
rect 1483 3682 1503 3686
rect 1507 3682 1631 3686
rect 1635 3682 1695 3686
rect 1699 3682 1791 3686
rect 1795 3682 1887 3686
rect 1891 3682 2007 3686
rect 2011 3682 2031 3686
rect 103 3681 2031 3682
rect 2037 3681 2038 3687
rect 2018 3629 2019 3635
rect 2025 3634 3967 3635
rect 2025 3630 2047 3634
rect 2051 3630 2071 3634
rect 2075 3630 2111 3634
rect 2115 3630 2263 3634
rect 2267 3630 2271 3634
rect 2275 3630 2455 3634
rect 2459 3630 2479 3634
rect 2483 3630 2655 3634
rect 2659 3630 2695 3634
rect 2699 3630 2871 3634
rect 2875 3630 2911 3634
rect 2915 3630 3095 3634
rect 3099 3630 3119 3634
rect 3123 3630 3319 3634
rect 3323 3630 3327 3634
rect 3331 3630 3519 3634
rect 3523 3630 3567 3634
rect 3571 3630 3727 3634
rect 3731 3630 3943 3634
rect 3947 3630 3967 3634
rect 2025 3629 3967 3630
rect 3973 3629 3974 3635
rect 84 3597 85 3603
rect 91 3602 2019 3603
rect 91 3598 111 3602
rect 115 3598 271 3602
rect 275 3598 367 3602
rect 371 3598 415 3602
rect 419 3598 519 3602
rect 523 3598 575 3602
rect 579 3598 679 3602
rect 683 3598 735 3602
rect 739 3598 847 3602
rect 851 3598 895 3602
rect 899 3598 1015 3602
rect 1019 3598 1055 3602
rect 1059 3598 1175 3602
rect 1179 3598 1215 3602
rect 1219 3598 1327 3602
rect 1331 3598 1375 3602
rect 1379 3598 1479 3602
rect 1483 3598 1543 3602
rect 1547 3598 1631 3602
rect 1635 3598 1791 3602
rect 1795 3598 2007 3602
rect 2011 3598 2019 3602
rect 91 3597 2019 3598
rect 2025 3597 2026 3603
rect 2030 3537 2031 3543
rect 2037 3542 3979 3543
rect 2037 3538 2047 3542
rect 2051 3538 2111 3542
rect 2115 3538 2271 3542
rect 2275 3538 2287 3542
rect 2291 3538 2383 3542
rect 2387 3538 2455 3542
rect 2459 3538 2479 3542
rect 2483 3538 2575 3542
rect 2579 3538 2655 3542
rect 2659 3538 2671 3542
rect 2675 3538 2767 3542
rect 2771 3538 2871 3542
rect 2875 3538 2983 3542
rect 2987 3538 3095 3542
rect 3099 3538 3103 3542
rect 3107 3538 3223 3542
rect 3227 3538 3327 3542
rect 3331 3538 3351 3542
rect 3355 3538 3487 3542
rect 3491 3538 3567 3542
rect 3571 3538 3943 3542
rect 3947 3538 3979 3542
rect 2037 3537 3979 3538
rect 3985 3537 3986 3543
rect 96 3513 97 3519
rect 103 3518 2031 3519
rect 103 3514 111 3518
rect 115 3514 159 3518
rect 163 3514 271 3518
rect 275 3514 287 3518
rect 291 3514 415 3518
rect 419 3514 423 3518
rect 427 3514 559 3518
rect 563 3514 575 3518
rect 579 3514 695 3518
rect 699 3514 735 3518
rect 739 3514 831 3518
rect 835 3514 895 3518
rect 899 3514 967 3518
rect 971 3514 1055 3518
rect 1059 3514 1095 3518
rect 1099 3514 1215 3518
rect 1219 3514 1231 3518
rect 1235 3514 1367 3518
rect 1371 3514 1375 3518
rect 1379 3514 1543 3518
rect 1547 3514 2007 3518
rect 2011 3514 2031 3518
rect 103 3513 2031 3514
rect 2037 3513 2038 3519
rect 2018 3461 2019 3467
rect 2025 3466 3967 3467
rect 2025 3462 2047 3466
rect 2051 3462 2287 3466
rect 2291 3462 2383 3466
rect 2387 3462 2479 3466
rect 2483 3462 2487 3466
rect 2491 3462 2575 3466
rect 2579 3462 2583 3466
rect 2587 3462 2671 3466
rect 2675 3462 2679 3466
rect 2683 3462 2767 3466
rect 2771 3462 2783 3466
rect 2787 3462 2871 3466
rect 2875 3462 2895 3466
rect 2899 3462 2983 3466
rect 2987 3462 3015 3466
rect 3019 3462 3103 3466
rect 3107 3462 3143 3466
rect 3147 3462 3223 3466
rect 3227 3462 3271 3466
rect 3275 3462 3351 3466
rect 3355 3462 3407 3466
rect 3411 3462 3487 3466
rect 3491 3462 3943 3466
rect 3947 3462 3967 3466
rect 2025 3461 3967 3462
rect 3973 3461 3974 3467
rect 84 3429 85 3435
rect 91 3434 2019 3435
rect 91 3430 111 3434
rect 115 3430 135 3434
rect 139 3430 159 3434
rect 163 3430 247 3434
rect 251 3430 287 3434
rect 291 3430 383 3434
rect 387 3430 423 3434
rect 427 3430 527 3434
rect 531 3430 559 3434
rect 563 3430 671 3434
rect 675 3430 695 3434
rect 699 3430 815 3434
rect 819 3430 831 3434
rect 835 3430 967 3434
rect 971 3430 1095 3434
rect 1099 3430 1119 3434
rect 1123 3430 1231 3434
rect 1235 3430 1271 3434
rect 1275 3430 1367 3434
rect 1371 3430 2007 3434
rect 2011 3430 2019 3434
rect 91 3429 2019 3430
rect 2025 3429 2026 3435
rect 2030 3377 2031 3383
rect 2037 3382 3979 3383
rect 2037 3378 2047 3382
rect 2051 3378 2351 3382
rect 2355 3378 2479 3382
rect 2483 3378 2487 3382
rect 2491 3378 2583 3382
rect 2587 3378 2615 3382
rect 2619 3378 2679 3382
rect 2683 3378 2751 3382
rect 2755 3378 2783 3382
rect 2787 3378 2887 3382
rect 2891 3378 2895 3382
rect 2899 3378 3015 3382
rect 3019 3378 3023 3382
rect 3027 3378 3143 3382
rect 3147 3378 3159 3382
rect 3163 3378 3271 3382
rect 3275 3378 3303 3382
rect 3307 3378 3407 3382
rect 3411 3378 3943 3382
rect 3947 3378 3979 3382
rect 2037 3377 3979 3378
rect 3985 3377 3986 3383
rect 96 3345 97 3351
rect 103 3350 2031 3351
rect 103 3346 111 3350
rect 115 3346 135 3350
rect 139 3346 247 3350
rect 251 3346 263 3350
rect 267 3346 383 3350
rect 387 3346 431 3350
rect 435 3346 527 3350
rect 531 3346 599 3350
rect 603 3346 671 3350
rect 675 3346 767 3350
rect 771 3346 815 3350
rect 819 3346 927 3350
rect 931 3346 967 3350
rect 971 3346 1087 3350
rect 1091 3346 1119 3350
rect 1123 3346 1239 3350
rect 1243 3346 1271 3350
rect 1275 3346 1391 3350
rect 1395 3346 1551 3350
rect 1555 3346 2007 3350
rect 2011 3346 2031 3350
rect 103 3345 2031 3346
rect 2037 3345 2038 3351
rect 2018 3297 2019 3303
rect 2025 3302 3967 3303
rect 2025 3298 2047 3302
rect 2051 3298 2127 3302
rect 2131 3298 2295 3302
rect 2299 3298 2351 3302
rect 2355 3298 2455 3302
rect 2459 3298 2479 3302
rect 2483 3298 2615 3302
rect 2619 3298 2751 3302
rect 2755 3298 2775 3302
rect 2779 3298 2887 3302
rect 2891 3298 2935 3302
rect 2939 3298 3023 3302
rect 3027 3298 3095 3302
rect 3099 3298 3159 3302
rect 3163 3298 3263 3302
rect 3267 3298 3303 3302
rect 3307 3298 3943 3302
rect 3947 3298 3967 3302
rect 2025 3297 3967 3298
rect 3973 3297 3974 3303
rect 84 3261 85 3267
rect 91 3266 2019 3267
rect 91 3262 111 3266
rect 115 3262 135 3266
rect 139 3262 143 3266
rect 147 3262 263 3266
rect 267 3262 295 3266
rect 299 3262 431 3266
rect 435 3262 455 3266
rect 459 3262 599 3266
rect 603 3262 623 3266
rect 627 3262 767 3266
rect 771 3262 791 3266
rect 795 3262 927 3266
rect 931 3262 959 3266
rect 963 3262 1087 3266
rect 1091 3262 1127 3266
rect 1131 3262 1239 3266
rect 1243 3262 1303 3266
rect 1307 3262 1391 3266
rect 1395 3262 1479 3266
rect 1483 3262 1551 3266
rect 1555 3262 2007 3266
rect 2011 3262 2019 3266
rect 91 3261 2019 3262
rect 2025 3261 2026 3267
rect 2030 3221 2031 3227
rect 2037 3226 3979 3227
rect 2037 3222 2047 3226
rect 2051 3222 2071 3226
rect 2075 3222 2127 3226
rect 2131 3222 2207 3226
rect 2211 3222 2295 3226
rect 2299 3222 2375 3226
rect 2379 3222 2455 3226
rect 2459 3222 2543 3226
rect 2547 3222 2615 3226
rect 2619 3222 2703 3226
rect 2707 3222 2775 3226
rect 2779 3222 2863 3226
rect 2867 3222 2935 3226
rect 2939 3222 3015 3226
rect 3019 3222 3095 3226
rect 3099 3222 3167 3226
rect 3171 3222 3263 3226
rect 3267 3222 3327 3226
rect 3331 3222 3943 3226
rect 3947 3222 3979 3226
rect 2037 3221 3979 3222
rect 3985 3221 3986 3227
rect 96 3185 97 3191
rect 103 3190 2031 3191
rect 103 3186 111 3190
rect 115 3186 143 3190
rect 147 3186 295 3190
rect 299 3186 431 3190
rect 435 3186 455 3190
rect 459 3186 567 3190
rect 571 3186 623 3190
rect 627 3186 703 3190
rect 707 3186 791 3190
rect 795 3186 855 3190
rect 859 3186 959 3190
rect 963 3186 1031 3190
rect 1035 3186 1127 3190
rect 1131 3186 1231 3190
rect 1235 3186 1303 3190
rect 1307 3186 1455 3190
rect 1459 3186 1479 3190
rect 1483 3186 1687 3190
rect 1691 3186 1903 3190
rect 1907 3186 2007 3190
rect 2011 3186 2031 3190
rect 103 3185 2031 3186
rect 2037 3185 2038 3191
rect 2018 3141 2019 3147
rect 2025 3146 3967 3147
rect 2025 3142 2047 3146
rect 2051 3142 2071 3146
rect 2075 3142 2207 3146
rect 2211 3142 2343 3146
rect 2347 3142 2375 3146
rect 2379 3142 2543 3146
rect 2547 3142 2631 3146
rect 2635 3142 2703 3146
rect 2707 3142 2863 3146
rect 2867 3142 2903 3146
rect 2907 3142 3015 3146
rect 3019 3142 3167 3146
rect 3171 3142 3175 3146
rect 3179 3142 3327 3146
rect 3331 3142 3447 3146
rect 3451 3142 3943 3146
rect 3947 3142 3967 3146
rect 2025 3141 3967 3142
rect 3973 3141 3974 3147
rect 84 3109 85 3115
rect 91 3114 2019 3115
rect 91 3110 111 3114
rect 115 3110 295 3114
rect 299 3110 311 3114
rect 315 3110 407 3114
rect 411 3110 431 3114
rect 435 3110 503 3114
rect 507 3110 567 3114
rect 571 3110 599 3114
rect 603 3110 695 3114
rect 699 3110 703 3114
rect 707 3110 807 3114
rect 811 3110 855 3114
rect 859 3110 943 3114
rect 947 3110 1031 3114
rect 1035 3110 1087 3114
rect 1091 3110 1231 3114
rect 1235 3110 1247 3114
rect 1251 3110 1407 3114
rect 1411 3110 1455 3114
rect 1459 3110 1575 3114
rect 1579 3110 1687 3114
rect 1691 3110 1751 3114
rect 1755 3110 1903 3114
rect 1907 3110 2007 3114
rect 2011 3110 2019 3114
rect 91 3109 2019 3110
rect 2025 3109 2026 3115
rect 2030 3061 2031 3067
rect 2037 3066 3979 3067
rect 2037 3062 2047 3066
rect 2051 3062 2071 3066
rect 2075 3062 2343 3066
rect 2347 3062 2487 3066
rect 2491 3062 2615 3066
rect 2619 3062 2631 3066
rect 2635 3062 2743 3066
rect 2747 3062 2863 3066
rect 2867 3062 2903 3066
rect 2907 3062 2983 3066
rect 2987 3062 3103 3066
rect 3107 3062 3175 3066
rect 3179 3062 3215 3066
rect 3219 3062 3327 3066
rect 3331 3062 3431 3066
rect 3435 3062 3447 3066
rect 3451 3062 3535 3066
rect 3539 3062 3639 3066
rect 3643 3062 3743 3066
rect 3747 3062 3839 3066
rect 3843 3062 3943 3066
rect 3947 3062 3979 3066
rect 2037 3061 3979 3062
rect 3985 3061 3986 3067
rect 96 3033 97 3039
rect 103 3038 2031 3039
rect 103 3034 111 3038
rect 115 3034 311 3038
rect 315 3034 407 3038
rect 411 3034 423 3038
rect 427 3034 503 3038
rect 507 3034 519 3038
rect 523 3034 599 3038
rect 603 3034 615 3038
rect 619 3034 695 3038
rect 699 3034 711 3038
rect 715 3034 807 3038
rect 811 3034 815 3038
rect 819 3034 935 3038
rect 939 3034 943 3038
rect 947 3034 1055 3038
rect 1059 3034 1087 3038
rect 1091 3034 1183 3038
rect 1187 3034 1247 3038
rect 1251 3034 1311 3038
rect 1315 3034 1407 3038
rect 1411 3034 1431 3038
rect 1435 3034 1551 3038
rect 1555 3034 1575 3038
rect 1579 3034 1671 3038
rect 1675 3034 1751 3038
rect 1755 3034 1799 3038
rect 1803 3034 1903 3038
rect 1907 3034 2007 3038
rect 2011 3034 2031 3038
rect 103 3033 2031 3034
rect 2037 3033 2038 3039
rect 2018 2981 2019 2987
rect 2025 2986 3967 2987
rect 2025 2982 2047 2986
rect 2051 2982 2407 2986
rect 2411 2982 2487 2986
rect 2491 2982 2575 2986
rect 2579 2982 2615 2986
rect 2619 2982 2743 2986
rect 2747 2982 2767 2986
rect 2771 2982 2863 2986
rect 2867 2982 2967 2986
rect 2971 2982 2983 2986
rect 2987 2982 3103 2986
rect 3107 2982 3183 2986
rect 3187 2982 3215 2986
rect 3219 2982 3327 2986
rect 3331 2982 3399 2986
rect 3403 2982 3431 2986
rect 3435 2982 3535 2986
rect 3539 2982 3623 2986
rect 3627 2982 3639 2986
rect 3643 2982 3743 2986
rect 3747 2982 3839 2986
rect 3843 2982 3943 2986
rect 3947 2982 3967 2986
rect 2025 2981 3967 2982
rect 3973 2981 3974 2987
rect 84 2933 85 2939
rect 91 2938 2019 2939
rect 91 2934 111 2938
rect 115 2934 423 2938
rect 427 2934 519 2938
rect 523 2934 615 2938
rect 619 2934 711 2938
rect 715 2934 815 2938
rect 819 2934 935 2938
rect 939 2934 1055 2938
rect 1059 2934 1183 2938
rect 1187 2934 1311 2938
rect 1315 2934 1431 2938
rect 1435 2934 1479 2938
rect 1483 2934 1551 2938
rect 1555 2934 1575 2938
rect 1579 2934 1671 2938
rect 1675 2934 1767 2938
rect 1771 2934 1799 2938
rect 1803 2934 1863 2938
rect 1867 2934 1903 2938
rect 1907 2934 2007 2938
rect 2011 2934 2019 2938
rect 91 2933 2019 2934
rect 2025 2933 2026 2939
rect 2030 2889 2031 2895
rect 2037 2894 3979 2895
rect 2037 2890 2047 2894
rect 2051 2890 2407 2894
rect 2411 2890 2551 2894
rect 2555 2890 2575 2894
rect 2579 2890 2671 2894
rect 2675 2890 2767 2894
rect 2771 2890 2799 2894
rect 2803 2890 2927 2894
rect 2931 2890 2967 2894
rect 2971 2890 3055 2894
rect 3059 2890 3183 2894
rect 3187 2890 3311 2894
rect 3315 2890 3399 2894
rect 3403 2890 3439 2894
rect 3443 2890 3575 2894
rect 3579 2890 3623 2894
rect 3627 2890 3839 2894
rect 3843 2890 3943 2894
rect 3947 2890 3979 2894
rect 2037 2889 3979 2890
rect 3985 2889 3986 2895
rect 96 2849 97 2855
rect 103 2854 2031 2855
rect 103 2850 111 2854
rect 115 2850 279 2854
rect 283 2850 447 2854
rect 451 2850 631 2854
rect 635 2850 815 2854
rect 819 2850 999 2854
rect 1003 2850 1183 2854
rect 1187 2850 1359 2854
rect 1363 2850 1479 2854
rect 1483 2850 1527 2854
rect 1531 2850 1575 2854
rect 1579 2850 1671 2854
rect 1675 2850 1695 2854
rect 1699 2850 1767 2854
rect 1771 2850 1863 2854
rect 1867 2850 2007 2854
rect 2011 2850 2031 2854
rect 103 2849 2031 2850
rect 2037 2849 2038 2855
rect 2018 2813 2019 2819
rect 2025 2818 3967 2819
rect 2025 2814 2047 2818
rect 2051 2814 2439 2818
rect 2443 2814 2551 2818
rect 2555 2814 2567 2818
rect 2571 2814 2671 2818
rect 2675 2814 2695 2818
rect 2699 2814 2799 2818
rect 2803 2814 2831 2818
rect 2835 2814 2927 2818
rect 2931 2814 2967 2818
rect 2971 2814 3055 2818
rect 3059 2814 3103 2818
rect 3107 2814 3183 2818
rect 3187 2814 3247 2818
rect 3251 2814 3311 2818
rect 3315 2814 3391 2818
rect 3395 2814 3439 2818
rect 3443 2814 3543 2818
rect 3547 2814 3575 2818
rect 3579 2814 3703 2818
rect 3707 2814 3839 2818
rect 3843 2814 3943 2818
rect 3947 2814 3967 2818
rect 2025 2813 3967 2814
rect 3973 2813 3974 2819
rect 84 2773 85 2779
rect 91 2778 2019 2779
rect 91 2774 111 2778
rect 115 2774 239 2778
rect 243 2774 279 2778
rect 283 2774 351 2778
rect 355 2774 447 2778
rect 451 2774 471 2778
rect 475 2774 607 2778
rect 611 2774 631 2778
rect 635 2774 743 2778
rect 747 2774 815 2778
rect 819 2774 879 2778
rect 883 2774 999 2778
rect 1003 2774 1015 2778
rect 1019 2774 1151 2778
rect 1155 2774 1183 2778
rect 1187 2774 1287 2778
rect 1291 2774 1359 2778
rect 1363 2774 1423 2778
rect 1427 2774 1527 2778
rect 1531 2774 1567 2778
rect 1571 2774 1695 2778
rect 1699 2774 1863 2778
rect 1867 2774 2007 2778
rect 2011 2774 2019 2778
rect 91 2773 2019 2774
rect 2025 2773 2026 2779
rect 2030 2729 2031 2735
rect 2037 2734 3979 2735
rect 2037 2730 2047 2734
rect 2051 2730 2335 2734
rect 2339 2730 2439 2734
rect 2443 2730 2495 2734
rect 2499 2730 2567 2734
rect 2571 2730 2663 2734
rect 2667 2730 2695 2734
rect 2699 2730 2831 2734
rect 2835 2730 2967 2734
rect 2971 2730 2999 2734
rect 3003 2730 3103 2734
rect 3107 2730 3167 2734
rect 3171 2730 3247 2734
rect 3251 2730 3335 2734
rect 3339 2730 3391 2734
rect 3395 2730 3511 2734
rect 3515 2730 3543 2734
rect 3547 2730 3687 2734
rect 3691 2730 3703 2734
rect 3707 2730 3839 2734
rect 3843 2730 3943 2734
rect 3947 2730 3979 2734
rect 2037 2729 3979 2730
rect 3985 2729 3986 2735
rect 96 2697 97 2703
rect 103 2702 2031 2703
rect 103 2698 111 2702
rect 115 2698 223 2702
rect 227 2698 239 2702
rect 243 2698 351 2702
rect 355 2698 367 2702
rect 371 2698 471 2702
rect 475 2698 503 2702
rect 507 2698 607 2702
rect 611 2698 639 2702
rect 643 2698 743 2702
rect 747 2698 767 2702
rect 771 2698 879 2702
rect 883 2698 887 2702
rect 891 2698 999 2702
rect 1003 2698 1015 2702
rect 1019 2698 1111 2702
rect 1115 2698 1151 2702
rect 1155 2698 1231 2702
rect 1235 2698 1287 2702
rect 1291 2698 1351 2702
rect 1355 2698 1423 2702
rect 1427 2698 1567 2702
rect 1571 2698 2007 2702
rect 2011 2698 2031 2702
rect 103 2697 2031 2698
rect 2037 2697 2038 2703
rect 2018 2649 2019 2655
rect 2025 2654 3967 2655
rect 2025 2650 2047 2654
rect 2051 2650 2127 2654
rect 2131 2650 2279 2654
rect 2283 2650 2335 2654
rect 2339 2650 2447 2654
rect 2451 2650 2495 2654
rect 2499 2650 2623 2654
rect 2627 2650 2663 2654
rect 2667 2650 2807 2654
rect 2811 2650 2831 2654
rect 2835 2650 2991 2654
rect 2995 2650 2999 2654
rect 3003 2650 3167 2654
rect 3171 2650 3175 2654
rect 3179 2650 3335 2654
rect 3339 2650 3351 2654
rect 3355 2650 3511 2654
rect 3515 2650 3519 2654
rect 3523 2650 3687 2654
rect 3691 2650 3839 2654
rect 3843 2650 3943 2654
rect 3947 2650 3967 2654
rect 2025 2649 3967 2650
rect 3973 2649 3974 2655
rect 84 2621 85 2627
rect 91 2626 2019 2627
rect 91 2622 111 2626
rect 115 2622 175 2626
rect 179 2622 223 2626
rect 227 2622 367 2626
rect 371 2622 503 2626
rect 507 2622 543 2626
rect 547 2622 639 2626
rect 643 2622 711 2626
rect 715 2622 767 2626
rect 771 2622 863 2626
rect 867 2622 887 2626
rect 891 2622 999 2626
rect 1003 2622 1007 2626
rect 1011 2622 1111 2626
rect 1115 2622 1143 2626
rect 1147 2622 1231 2626
rect 1235 2622 1279 2626
rect 1283 2622 1351 2626
rect 1355 2622 1423 2626
rect 1427 2622 2007 2626
rect 2011 2622 2019 2626
rect 91 2621 2019 2622
rect 2025 2621 2026 2627
rect 2030 2565 2031 2571
rect 2037 2570 3979 2571
rect 2037 2566 2047 2570
rect 2051 2566 2071 2570
rect 2075 2566 2127 2570
rect 2131 2566 2183 2570
rect 2187 2566 2279 2570
rect 2283 2566 2319 2570
rect 2323 2566 2447 2570
rect 2451 2566 2471 2570
rect 2475 2566 2623 2570
rect 2627 2566 2639 2570
rect 2643 2566 2807 2570
rect 2811 2566 2823 2570
rect 2827 2566 2991 2570
rect 2995 2566 3031 2570
rect 3035 2566 3175 2570
rect 3179 2566 3263 2570
rect 3267 2566 3351 2570
rect 3355 2566 3503 2570
rect 3507 2566 3519 2570
rect 3523 2566 3687 2570
rect 3691 2566 3743 2570
rect 3747 2566 3839 2570
rect 3843 2566 3943 2570
rect 3947 2566 3979 2570
rect 2037 2565 3979 2566
rect 3985 2565 3986 2571
rect 96 2541 97 2547
rect 103 2546 2031 2547
rect 103 2542 111 2546
rect 115 2542 135 2546
rect 139 2542 175 2546
rect 179 2542 271 2546
rect 275 2542 367 2546
rect 371 2542 439 2546
rect 443 2542 543 2546
rect 547 2542 607 2546
rect 611 2542 711 2546
rect 715 2542 775 2546
rect 779 2542 863 2546
rect 867 2542 927 2546
rect 931 2542 1007 2546
rect 1011 2542 1079 2546
rect 1083 2542 1143 2546
rect 1147 2542 1223 2546
rect 1227 2542 1279 2546
rect 1283 2542 1359 2546
rect 1363 2542 1423 2546
rect 1427 2542 1495 2546
rect 1499 2542 1639 2546
rect 1643 2542 2007 2546
rect 2011 2542 2031 2546
rect 103 2541 2031 2542
rect 2037 2541 2038 2547
rect 2018 2485 2019 2491
rect 2025 2490 3967 2491
rect 2025 2486 2047 2490
rect 2051 2486 2071 2490
rect 2075 2486 2183 2490
rect 2187 2486 2215 2490
rect 2219 2486 2319 2490
rect 2323 2486 2383 2490
rect 2387 2486 2471 2490
rect 2475 2486 2559 2490
rect 2563 2486 2639 2490
rect 2643 2486 2751 2490
rect 2755 2486 2823 2490
rect 2827 2486 2951 2490
rect 2955 2486 3031 2490
rect 3035 2486 3167 2490
rect 3171 2486 3263 2490
rect 3267 2486 3391 2490
rect 3395 2486 3503 2490
rect 3507 2486 3623 2490
rect 3627 2486 3743 2490
rect 3747 2486 3839 2490
rect 3843 2486 3943 2490
rect 3947 2486 3967 2490
rect 2025 2485 3967 2486
rect 3973 2485 3974 2491
rect 84 2461 85 2467
rect 91 2466 2019 2467
rect 91 2462 111 2466
rect 115 2462 135 2466
rect 139 2462 271 2466
rect 275 2462 311 2466
rect 315 2462 439 2466
rect 443 2462 511 2466
rect 515 2462 607 2466
rect 611 2462 711 2466
rect 715 2462 775 2466
rect 779 2462 903 2466
rect 907 2462 927 2466
rect 931 2462 1079 2466
rect 1083 2462 1223 2466
rect 1227 2462 1239 2466
rect 1243 2462 1359 2466
rect 1363 2462 1391 2466
rect 1395 2462 1495 2466
rect 1499 2462 1527 2466
rect 1531 2462 1639 2466
rect 1643 2462 1663 2466
rect 1667 2462 1791 2466
rect 1795 2462 1903 2466
rect 1907 2462 2007 2466
rect 2011 2462 2019 2466
rect 91 2461 2019 2462
rect 2025 2461 2026 2467
rect 2030 2393 2031 2399
rect 2037 2398 3979 2399
rect 2037 2394 2047 2398
rect 2051 2394 2071 2398
rect 2075 2394 2215 2398
rect 2219 2394 2247 2398
rect 2251 2394 2383 2398
rect 2387 2394 2431 2398
rect 2435 2394 2559 2398
rect 2563 2394 2607 2398
rect 2611 2394 2751 2398
rect 2755 2394 2775 2398
rect 2779 2394 2935 2398
rect 2939 2394 2951 2398
rect 2955 2394 3103 2398
rect 3107 2394 3167 2398
rect 3171 2394 3391 2398
rect 3395 2394 3623 2398
rect 3627 2394 3839 2398
rect 3843 2394 3943 2398
rect 3947 2394 3979 2398
rect 2037 2393 3979 2394
rect 3985 2393 3986 2399
rect 2030 2391 2038 2393
rect 96 2385 97 2391
rect 103 2390 2031 2391
rect 103 2386 111 2390
rect 115 2386 135 2390
rect 139 2386 311 2390
rect 315 2386 327 2390
rect 331 2386 511 2390
rect 515 2386 551 2390
rect 555 2386 711 2390
rect 715 2386 767 2390
rect 771 2386 903 2390
rect 907 2386 975 2390
rect 979 2386 1079 2390
rect 1083 2386 1175 2390
rect 1179 2386 1239 2390
rect 1243 2386 1367 2390
rect 1371 2386 1391 2390
rect 1395 2386 1527 2390
rect 1531 2386 1551 2390
rect 1555 2386 1663 2390
rect 1667 2386 1735 2390
rect 1739 2386 1791 2390
rect 1795 2386 1903 2390
rect 1907 2386 2007 2390
rect 2011 2386 2031 2390
rect 103 2385 2031 2386
rect 2037 2385 2038 2391
rect 2018 2317 2019 2323
rect 2025 2322 3967 2323
rect 2025 2318 2047 2322
rect 2051 2318 2071 2322
rect 2075 2318 2175 2322
rect 2179 2318 2247 2322
rect 2251 2318 2311 2322
rect 2315 2318 2431 2322
rect 2435 2318 2447 2322
rect 2451 2318 2591 2322
rect 2595 2318 2607 2322
rect 2611 2318 2751 2322
rect 2755 2318 2775 2322
rect 2779 2318 2935 2322
rect 2939 2318 3103 2322
rect 3107 2318 3143 2322
rect 3147 2318 3375 2322
rect 3379 2318 3615 2322
rect 3619 2318 3839 2322
rect 3843 2318 3943 2322
rect 3947 2318 3967 2322
rect 2025 2317 3967 2318
rect 3973 2317 3974 2323
rect 84 2301 85 2307
rect 91 2306 2019 2307
rect 91 2302 111 2306
rect 115 2302 135 2306
rect 139 2302 271 2306
rect 275 2302 327 2306
rect 331 2302 431 2306
rect 435 2302 551 2306
rect 555 2302 591 2306
rect 595 2302 751 2306
rect 755 2302 767 2306
rect 771 2302 919 2306
rect 923 2302 975 2306
rect 979 2302 1087 2306
rect 1091 2302 1175 2306
rect 1179 2302 1263 2306
rect 1267 2302 1367 2306
rect 1371 2302 1447 2306
rect 1451 2302 1551 2306
rect 1555 2302 1631 2306
rect 1635 2302 1735 2306
rect 1739 2302 1815 2306
rect 1819 2302 1903 2306
rect 1907 2302 2007 2306
rect 2011 2302 2019 2306
rect 91 2301 2019 2302
rect 2025 2301 2026 2307
rect 2030 2233 2031 2239
rect 2037 2238 3979 2239
rect 2037 2234 2047 2238
rect 2051 2234 2071 2238
rect 2075 2234 2111 2238
rect 2115 2234 2175 2238
rect 2179 2234 2255 2238
rect 2259 2234 2311 2238
rect 2315 2234 2407 2238
rect 2411 2234 2447 2238
rect 2451 2234 2559 2238
rect 2563 2234 2591 2238
rect 2595 2234 2719 2238
rect 2723 2234 2751 2238
rect 2755 2234 2879 2238
rect 2883 2234 2935 2238
rect 2939 2234 3047 2238
rect 3051 2234 3143 2238
rect 3147 2234 3223 2238
rect 3227 2234 3375 2238
rect 3379 2234 3407 2238
rect 3411 2234 3591 2238
rect 3595 2234 3615 2238
rect 3619 2234 3783 2238
rect 3787 2234 3839 2238
rect 3843 2234 3943 2238
rect 3947 2234 3979 2238
rect 2037 2233 3979 2234
rect 3985 2233 3986 2239
rect 2030 2231 2038 2233
rect 96 2225 97 2231
rect 103 2230 2031 2231
rect 103 2226 111 2230
rect 115 2226 135 2230
rect 139 2226 159 2230
rect 163 2226 271 2230
rect 275 2226 327 2230
rect 331 2226 431 2230
rect 435 2226 495 2230
rect 499 2226 591 2230
rect 595 2226 679 2230
rect 683 2226 751 2230
rect 755 2226 879 2230
rect 883 2226 919 2230
rect 923 2226 1087 2230
rect 1091 2226 1095 2230
rect 1099 2226 1263 2230
rect 1267 2226 1327 2230
rect 1331 2226 1447 2230
rect 1451 2226 1567 2230
rect 1571 2226 1631 2230
rect 1635 2226 1815 2230
rect 1819 2226 2007 2230
rect 2011 2226 2031 2230
rect 103 2225 2031 2226
rect 2037 2225 2038 2231
rect 84 2149 85 2155
rect 91 2154 2019 2155
rect 91 2150 111 2154
rect 115 2150 159 2154
rect 163 2150 223 2154
rect 227 2150 327 2154
rect 331 2150 359 2154
rect 363 2150 495 2154
rect 499 2150 639 2154
rect 643 2150 679 2154
rect 683 2150 783 2154
rect 787 2150 879 2154
rect 883 2150 935 2154
rect 939 2150 1095 2154
rect 1099 2150 1263 2154
rect 1267 2150 1327 2154
rect 1331 2150 1447 2154
rect 1451 2150 1567 2154
rect 1571 2150 1631 2154
rect 1635 2150 1815 2154
rect 1819 2150 1823 2154
rect 1827 2150 2007 2154
rect 2011 2150 2019 2154
rect 91 2149 2019 2150
rect 2025 2151 2026 2155
rect 2025 2150 3974 2151
rect 2025 2149 2047 2150
rect 2018 2146 2047 2149
rect 2051 2146 2111 2150
rect 2115 2146 2255 2150
rect 2259 2146 2287 2150
rect 2291 2146 2407 2150
rect 2411 2146 2431 2150
rect 2435 2146 2559 2150
rect 2563 2146 2583 2150
rect 2587 2146 2719 2150
rect 2723 2146 2735 2150
rect 2739 2146 2879 2150
rect 2883 2146 2887 2150
rect 2891 2146 3047 2150
rect 3051 2146 3207 2150
rect 3211 2146 3223 2150
rect 3227 2146 3367 2150
rect 3371 2146 3407 2150
rect 3411 2146 3527 2150
rect 3531 2146 3591 2150
rect 3595 2146 3695 2150
rect 3699 2146 3783 2150
rect 3787 2146 3839 2150
rect 3843 2146 3943 2150
rect 3947 2146 3974 2150
rect 2018 2145 3974 2146
rect 96 2065 97 2071
rect 103 2070 2031 2071
rect 103 2066 111 2070
rect 115 2066 223 2070
rect 227 2066 359 2070
rect 363 2066 375 2070
rect 379 2066 495 2070
rect 499 2066 615 2070
rect 619 2066 639 2070
rect 643 2066 751 2070
rect 755 2066 783 2070
rect 787 2066 895 2070
rect 899 2066 935 2070
rect 939 2066 1047 2070
rect 1051 2066 1095 2070
rect 1099 2066 1215 2070
rect 1219 2066 1263 2070
rect 1267 2066 1399 2070
rect 1403 2066 1447 2070
rect 1451 2066 1583 2070
rect 1587 2066 1631 2070
rect 1635 2066 1775 2070
rect 1779 2066 1823 2070
rect 1827 2066 2007 2070
rect 2011 2066 2031 2070
rect 103 2065 2031 2066
rect 2037 2067 2038 2071
rect 2037 2066 3986 2067
rect 2037 2065 2047 2066
rect 2030 2062 2047 2065
rect 2051 2062 2287 2066
rect 2291 2062 2431 2066
rect 2435 2062 2503 2066
rect 2507 2062 2583 2066
rect 2587 2062 2671 2066
rect 2675 2062 2735 2066
rect 2739 2062 2839 2066
rect 2843 2062 2887 2066
rect 2891 2062 3007 2066
rect 3011 2062 3047 2066
rect 3051 2062 3167 2066
rect 3171 2062 3207 2066
rect 3211 2062 3311 2066
rect 3315 2062 3367 2066
rect 3371 2062 3455 2066
rect 3459 2062 3527 2066
rect 3531 2062 3591 2066
rect 3595 2062 3695 2066
rect 3699 2062 3727 2066
rect 3731 2062 3839 2066
rect 3843 2062 3943 2066
rect 3947 2062 3986 2066
rect 2030 2061 3986 2062
rect 84 1981 85 1987
rect 91 1986 2019 1987
rect 91 1982 111 1986
rect 115 1982 375 1986
rect 379 1982 495 1986
rect 499 1982 511 1986
rect 515 1982 615 1986
rect 619 1982 623 1986
rect 627 1982 743 1986
rect 747 1982 751 1986
rect 755 1982 871 1986
rect 875 1982 895 1986
rect 899 1982 1007 1986
rect 1011 1982 1047 1986
rect 1051 1982 1143 1986
rect 1147 1982 1215 1986
rect 1219 1982 1279 1986
rect 1283 1982 1399 1986
rect 1403 1982 1415 1986
rect 1419 1982 1559 1986
rect 1563 1982 1583 1986
rect 1587 1982 1703 1986
rect 1707 1982 1775 1986
rect 1779 1982 2007 1986
rect 2011 1982 2019 1986
rect 91 1981 2019 1982
rect 2025 1986 3974 1987
rect 2025 1982 2047 1986
rect 2051 1982 2495 1986
rect 2499 1982 2503 1986
rect 2507 1982 2591 1986
rect 2595 1982 2671 1986
rect 2675 1982 2695 1986
rect 2699 1982 2807 1986
rect 2811 1982 2839 1986
rect 2843 1982 2927 1986
rect 2931 1982 3007 1986
rect 3011 1982 3047 1986
rect 3051 1982 3167 1986
rect 3171 1982 3175 1986
rect 3179 1982 3295 1986
rect 3299 1982 3311 1986
rect 3315 1982 3415 1986
rect 3419 1982 3455 1986
rect 3459 1982 3543 1986
rect 3547 1982 3591 1986
rect 3595 1982 3671 1986
rect 3675 1982 3727 1986
rect 3731 1982 3799 1986
rect 3803 1982 3839 1986
rect 3843 1982 3943 1986
rect 3947 1982 3974 1986
rect 2025 1981 3974 1982
rect 2030 1906 3986 1907
rect 2030 1903 2047 1906
rect 96 1897 97 1903
rect 103 1902 2031 1903
rect 103 1898 111 1902
rect 115 1898 511 1902
rect 515 1898 551 1902
rect 555 1898 623 1902
rect 627 1898 663 1902
rect 667 1898 743 1902
rect 747 1898 783 1902
rect 787 1898 871 1902
rect 875 1898 911 1902
rect 915 1898 1007 1902
rect 1011 1898 1047 1902
rect 1051 1898 1143 1902
rect 1147 1898 1175 1902
rect 1179 1898 1279 1902
rect 1283 1898 1311 1902
rect 1315 1898 1415 1902
rect 1419 1898 1447 1902
rect 1451 1898 1559 1902
rect 1563 1898 1583 1902
rect 1587 1898 1703 1902
rect 1707 1898 1719 1902
rect 1723 1898 2007 1902
rect 2011 1898 2031 1902
rect 103 1897 2031 1898
rect 2037 1902 2047 1903
rect 2051 1902 2071 1906
rect 2075 1902 2247 1906
rect 2251 1902 2439 1906
rect 2443 1902 2495 1906
rect 2499 1902 2591 1906
rect 2595 1902 2623 1906
rect 2627 1902 2695 1906
rect 2699 1902 2791 1906
rect 2795 1902 2807 1906
rect 2811 1902 2927 1906
rect 2931 1902 2959 1906
rect 2963 1902 3047 1906
rect 3051 1902 3127 1906
rect 3131 1902 3175 1906
rect 3179 1902 3295 1906
rect 3299 1902 3303 1906
rect 3307 1902 3415 1906
rect 3419 1902 3487 1906
rect 3491 1902 3543 1906
rect 3547 1902 3671 1906
rect 3675 1902 3799 1906
rect 3803 1902 3839 1906
rect 3843 1902 3943 1906
rect 3947 1902 3986 1906
rect 2037 1901 3986 1902
rect 2037 1897 2038 1901
rect 2018 1830 3974 1831
rect 2018 1827 2047 1830
rect 84 1821 85 1827
rect 91 1826 2019 1827
rect 91 1822 111 1826
rect 115 1822 503 1826
rect 507 1822 551 1826
rect 555 1822 615 1826
rect 619 1822 663 1826
rect 667 1822 735 1826
rect 739 1822 783 1826
rect 787 1822 863 1826
rect 867 1822 911 1826
rect 915 1822 999 1826
rect 1003 1822 1047 1826
rect 1051 1822 1151 1826
rect 1155 1822 1175 1826
rect 1179 1822 1311 1826
rect 1315 1822 1319 1826
rect 1323 1822 1447 1826
rect 1451 1822 1487 1826
rect 1491 1822 1583 1826
rect 1587 1822 1663 1826
rect 1667 1822 1719 1826
rect 1723 1822 1847 1826
rect 1851 1822 2007 1826
rect 2011 1822 2019 1826
rect 91 1821 2019 1822
rect 2025 1826 2047 1827
rect 2051 1826 2071 1830
rect 2075 1826 2095 1830
rect 2099 1826 2231 1830
rect 2235 1826 2247 1830
rect 2251 1826 2367 1830
rect 2371 1826 2439 1830
rect 2443 1826 2511 1830
rect 2515 1826 2623 1830
rect 2627 1826 2671 1830
rect 2675 1826 2791 1830
rect 2795 1826 2855 1830
rect 2859 1826 2959 1830
rect 2963 1826 3071 1830
rect 3075 1826 3127 1830
rect 3131 1826 3303 1830
rect 3307 1826 3487 1830
rect 3491 1826 3543 1830
rect 3547 1826 3671 1830
rect 3675 1826 3791 1830
rect 3795 1826 3839 1830
rect 3843 1826 3943 1830
rect 3947 1826 3974 1830
rect 2025 1825 3974 1826
rect 2025 1821 2026 1825
rect 2030 1754 3986 1755
rect 2030 1751 2047 1754
rect 96 1745 97 1751
rect 103 1750 2031 1751
rect 103 1746 111 1750
rect 115 1746 343 1750
rect 347 1746 463 1750
rect 467 1746 503 1750
rect 507 1746 591 1750
rect 595 1746 615 1750
rect 619 1746 719 1750
rect 723 1746 735 1750
rect 739 1746 847 1750
rect 851 1746 863 1750
rect 867 1746 983 1750
rect 987 1746 999 1750
rect 1003 1746 1127 1750
rect 1131 1746 1151 1750
rect 1155 1746 1279 1750
rect 1283 1746 1319 1750
rect 1323 1746 1439 1750
rect 1443 1746 1487 1750
rect 1491 1746 1599 1750
rect 1603 1746 1663 1750
rect 1667 1746 1847 1750
rect 1851 1746 2007 1750
rect 2011 1746 2031 1750
rect 103 1745 2031 1746
rect 2037 1750 2047 1751
rect 2051 1750 2095 1754
rect 2099 1750 2183 1754
rect 2187 1750 2231 1754
rect 2235 1750 2287 1754
rect 2291 1750 2367 1754
rect 2371 1750 2391 1754
rect 2395 1750 2495 1754
rect 2499 1750 2511 1754
rect 2515 1750 2599 1754
rect 2603 1750 2671 1754
rect 2675 1750 2703 1754
rect 2707 1750 2807 1754
rect 2811 1750 2855 1754
rect 2859 1750 2911 1754
rect 2915 1750 3015 1754
rect 3019 1750 3071 1754
rect 3075 1750 3127 1754
rect 3131 1750 3303 1754
rect 3307 1750 3543 1754
rect 3547 1750 3791 1754
rect 3795 1750 3943 1754
rect 3947 1750 3986 1754
rect 2037 1749 3986 1750
rect 2037 1745 2038 1749
rect 2018 1673 2019 1679
rect 2025 1678 3967 1679
rect 2025 1674 2047 1678
rect 2051 1674 2183 1678
rect 2187 1674 2231 1678
rect 2235 1674 2287 1678
rect 2291 1674 2367 1678
rect 2371 1674 2391 1678
rect 2395 1674 2495 1678
rect 2499 1674 2519 1678
rect 2523 1674 2599 1678
rect 2603 1674 2679 1678
rect 2683 1674 2703 1678
rect 2707 1674 2807 1678
rect 2811 1674 2847 1678
rect 2851 1674 2911 1678
rect 2915 1674 3015 1678
rect 3019 1674 3023 1678
rect 3027 1674 3127 1678
rect 3131 1674 3191 1678
rect 3195 1674 3359 1678
rect 3363 1674 3527 1678
rect 3531 1674 3695 1678
rect 3699 1674 3839 1678
rect 3843 1674 3943 1678
rect 3947 1674 3967 1678
rect 2025 1673 3967 1674
rect 3973 1673 3974 1679
rect 2018 1671 2026 1673
rect 84 1665 85 1671
rect 91 1670 2019 1671
rect 91 1666 111 1670
rect 115 1666 159 1670
rect 163 1666 295 1670
rect 299 1666 343 1670
rect 347 1666 455 1670
rect 459 1666 463 1670
rect 467 1666 591 1670
rect 595 1666 623 1670
rect 627 1666 719 1670
rect 723 1666 799 1670
rect 803 1666 847 1670
rect 851 1666 983 1670
rect 987 1666 1127 1670
rect 1131 1666 1167 1670
rect 1171 1666 1279 1670
rect 1283 1666 1351 1670
rect 1355 1666 1439 1670
rect 1443 1666 1543 1670
rect 1547 1666 1599 1670
rect 1603 1666 1735 1670
rect 1739 1666 2007 1670
rect 2011 1666 2019 1670
rect 91 1665 2019 1666
rect 2025 1665 2026 1671
rect 96 1589 97 1595
rect 103 1594 2031 1595
rect 103 1590 111 1594
rect 115 1590 135 1594
rect 139 1590 159 1594
rect 163 1590 255 1594
rect 259 1590 295 1594
rect 299 1590 423 1594
rect 427 1590 455 1594
rect 459 1590 607 1594
rect 611 1590 623 1594
rect 627 1590 799 1594
rect 803 1590 983 1594
rect 987 1590 991 1594
rect 995 1590 1167 1594
rect 1171 1590 1183 1594
rect 1187 1590 1351 1594
rect 1355 1590 1367 1594
rect 1371 1590 1543 1594
rect 1547 1590 1551 1594
rect 1555 1590 1735 1594
rect 1739 1590 1903 1594
rect 1907 1590 2007 1594
rect 2011 1590 2031 1594
rect 103 1589 2031 1590
rect 2037 1594 3986 1595
rect 2037 1590 2047 1594
rect 2051 1590 2071 1594
rect 2075 1590 2231 1594
rect 2235 1590 2271 1594
rect 2275 1590 2367 1594
rect 2371 1590 2495 1594
rect 2499 1590 2519 1594
rect 2523 1590 2679 1594
rect 2683 1590 2711 1594
rect 2715 1590 2847 1594
rect 2851 1590 2911 1594
rect 2915 1590 3023 1594
rect 3027 1590 3095 1594
rect 3099 1590 3191 1594
rect 3195 1590 3263 1594
rect 3267 1590 3359 1594
rect 3363 1590 3423 1594
rect 3427 1590 3527 1594
rect 3531 1590 3567 1594
rect 3571 1590 3695 1594
rect 3699 1590 3711 1594
rect 3715 1590 3839 1594
rect 3843 1590 3943 1594
rect 3947 1590 3986 1594
rect 2037 1589 3986 1590
rect 2018 1518 3974 1519
rect 2018 1515 2047 1518
rect 84 1509 85 1515
rect 91 1514 2019 1515
rect 91 1510 111 1514
rect 115 1510 135 1514
rect 139 1510 247 1514
rect 251 1510 255 1514
rect 259 1510 399 1514
rect 403 1510 423 1514
rect 427 1510 559 1514
rect 563 1510 607 1514
rect 611 1510 719 1514
rect 723 1510 799 1514
rect 803 1510 879 1514
rect 883 1510 991 1514
rect 995 1510 1039 1514
rect 1043 1510 1183 1514
rect 1187 1510 1319 1514
rect 1323 1510 1367 1514
rect 1371 1510 1447 1514
rect 1451 1510 1551 1514
rect 1555 1510 1567 1514
rect 1571 1510 1687 1514
rect 1691 1510 1735 1514
rect 1739 1510 1807 1514
rect 1811 1510 1903 1514
rect 1907 1510 2007 1514
rect 2011 1510 2019 1514
rect 91 1509 2019 1510
rect 2025 1514 2047 1515
rect 2051 1514 2071 1518
rect 2075 1514 2271 1518
rect 2275 1514 2431 1518
rect 2435 1514 2495 1518
rect 2499 1514 2711 1518
rect 2715 1514 2791 1518
rect 2795 1514 2911 1518
rect 2915 1514 3095 1518
rect 3099 1514 3127 1518
rect 3131 1514 3263 1518
rect 3267 1514 3423 1518
rect 3427 1514 3463 1518
rect 3467 1514 3567 1518
rect 3571 1514 3711 1518
rect 3715 1514 3799 1518
rect 3803 1514 3839 1518
rect 3843 1514 3943 1518
rect 3947 1514 3974 1518
rect 2025 1513 3974 1514
rect 2025 1509 2026 1513
rect 96 1433 97 1439
rect 103 1438 2031 1439
rect 103 1434 111 1438
rect 115 1434 135 1438
rect 139 1434 247 1438
rect 251 1434 263 1438
rect 267 1434 399 1438
rect 403 1434 431 1438
rect 435 1434 559 1438
rect 563 1434 607 1438
rect 611 1434 719 1438
rect 723 1434 791 1438
rect 795 1434 879 1438
rect 883 1434 975 1438
rect 979 1434 1039 1438
rect 1043 1434 1159 1438
rect 1163 1434 1183 1438
rect 1187 1434 1319 1438
rect 1323 1434 1351 1438
rect 1355 1434 1447 1438
rect 1451 1434 1543 1438
rect 1547 1434 1567 1438
rect 1571 1434 1687 1438
rect 1691 1434 1735 1438
rect 1739 1434 1807 1438
rect 1811 1434 1903 1438
rect 1907 1434 2007 1438
rect 2011 1434 2031 1438
rect 103 1433 2031 1434
rect 2037 1435 2038 1439
rect 2037 1434 3986 1435
rect 2037 1433 2047 1434
rect 2030 1430 2047 1433
rect 2051 1430 2071 1434
rect 2075 1430 2271 1434
rect 2275 1430 2431 1434
rect 2435 1430 2495 1434
rect 2499 1430 2711 1434
rect 2715 1430 2791 1434
rect 2795 1430 2911 1434
rect 2915 1430 3095 1434
rect 3099 1430 3127 1434
rect 3131 1430 3271 1434
rect 3275 1430 3439 1434
rect 3443 1430 3463 1434
rect 3467 1430 3607 1434
rect 3611 1430 3783 1434
rect 3787 1430 3799 1434
rect 3803 1430 3943 1434
rect 3947 1430 3986 1434
rect 2030 1429 3986 1430
rect 84 1353 85 1359
rect 91 1358 2019 1359
rect 91 1354 111 1358
rect 115 1354 135 1358
rect 139 1354 159 1358
rect 163 1354 263 1358
rect 267 1354 311 1358
rect 315 1354 431 1358
rect 435 1354 479 1358
rect 483 1354 607 1358
rect 611 1354 663 1358
rect 667 1354 791 1358
rect 795 1354 855 1358
rect 859 1354 975 1358
rect 979 1354 1047 1358
rect 1051 1354 1159 1358
rect 1163 1354 1247 1358
rect 1251 1354 1351 1358
rect 1355 1354 1447 1358
rect 1451 1354 1543 1358
rect 1547 1354 1655 1358
rect 1659 1354 1735 1358
rect 1739 1354 1863 1358
rect 1867 1354 1903 1358
rect 1907 1354 2007 1358
rect 2011 1354 2019 1358
rect 91 1353 2019 1354
rect 2025 1358 3974 1359
rect 2025 1354 2047 1358
rect 2051 1354 2071 1358
rect 2075 1354 2207 1358
rect 2211 1354 2271 1358
rect 2275 1354 2383 1358
rect 2387 1354 2495 1358
rect 2499 1354 2567 1358
rect 2571 1354 2711 1358
rect 2715 1354 2751 1358
rect 2755 1354 2911 1358
rect 2915 1354 2935 1358
rect 2939 1354 3095 1358
rect 3099 1354 3111 1358
rect 3115 1354 3271 1358
rect 3275 1354 3279 1358
rect 3283 1354 3439 1358
rect 3443 1354 3447 1358
rect 3451 1354 3607 1358
rect 3611 1354 3623 1358
rect 3627 1354 3783 1358
rect 3787 1354 3943 1358
rect 3947 1354 3974 1358
rect 2025 1353 3974 1354
rect 2030 1282 3986 1283
rect 2030 1279 2047 1282
rect 96 1273 97 1279
rect 103 1278 2031 1279
rect 103 1274 111 1278
rect 115 1274 159 1278
rect 163 1274 311 1278
rect 315 1274 407 1278
rect 411 1274 479 1278
rect 483 1274 543 1278
rect 547 1274 663 1278
rect 667 1274 695 1278
rect 699 1274 855 1278
rect 859 1274 1023 1278
rect 1027 1274 1047 1278
rect 1051 1274 1191 1278
rect 1195 1274 1247 1278
rect 1251 1274 1367 1278
rect 1371 1274 1447 1278
rect 1451 1274 1543 1278
rect 1547 1274 1655 1278
rect 1659 1274 1719 1278
rect 1723 1274 1863 1278
rect 1867 1274 1895 1278
rect 1899 1274 2007 1278
rect 2011 1274 2031 1278
rect 103 1273 2031 1274
rect 2037 1278 2047 1279
rect 2051 1278 2071 1282
rect 2075 1278 2151 1282
rect 2155 1278 2207 1282
rect 2211 1278 2287 1282
rect 2291 1278 2383 1282
rect 2387 1278 2431 1282
rect 2435 1278 2567 1282
rect 2571 1278 2583 1282
rect 2587 1278 2743 1282
rect 2747 1278 2751 1282
rect 2755 1278 2903 1282
rect 2907 1278 2935 1282
rect 2939 1278 3071 1282
rect 3075 1278 3111 1282
rect 3115 1278 3247 1282
rect 3251 1278 3279 1282
rect 3283 1278 3431 1282
rect 3435 1278 3447 1282
rect 3451 1278 3615 1282
rect 3619 1278 3623 1282
rect 3627 1278 3807 1282
rect 3811 1278 3943 1282
rect 3947 1278 3986 1282
rect 2037 1277 3986 1278
rect 2037 1273 2038 1277
rect 2018 1206 3974 1207
rect 2018 1203 2047 1206
rect 84 1197 85 1203
rect 91 1202 2019 1203
rect 91 1198 111 1202
rect 115 1198 407 1202
rect 411 1198 423 1202
rect 427 1198 543 1202
rect 547 1198 591 1202
rect 595 1198 695 1202
rect 699 1198 759 1202
rect 763 1198 855 1202
rect 859 1198 927 1202
rect 931 1198 1023 1202
rect 1027 1198 1095 1202
rect 1099 1198 1191 1202
rect 1195 1198 1247 1202
rect 1251 1198 1367 1202
rect 1371 1198 1399 1202
rect 1403 1198 1543 1202
rect 1547 1198 1687 1202
rect 1691 1198 1719 1202
rect 1723 1198 1839 1202
rect 1843 1198 1895 1202
rect 1899 1198 2007 1202
rect 2011 1198 2019 1202
rect 91 1197 2019 1198
rect 2025 1202 2047 1203
rect 2051 1202 2151 1206
rect 2155 1202 2287 1206
rect 2291 1202 2311 1206
rect 2315 1202 2415 1206
rect 2419 1202 2431 1206
rect 2435 1202 2527 1206
rect 2531 1202 2583 1206
rect 2587 1202 2639 1206
rect 2643 1202 2743 1206
rect 2747 1202 2767 1206
rect 2771 1202 2903 1206
rect 2907 1202 2911 1206
rect 2915 1202 3071 1206
rect 3075 1202 3247 1206
rect 3251 1202 3431 1206
rect 3435 1202 3439 1206
rect 3443 1202 3615 1206
rect 3619 1202 3631 1206
rect 3635 1202 3807 1206
rect 3811 1202 3831 1206
rect 3835 1202 3943 1206
rect 3947 1202 3974 1206
rect 2025 1201 3974 1202
rect 2025 1197 2026 1201
rect 2030 1126 3986 1127
rect 2030 1123 2047 1126
rect 96 1117 97 1123
rect 103 1122 2031 1123
rect 103 1118 111 1122
rect 115 1118 375 1122
rect 379 1118 423 1122
rect 427 1118 487 1122
rect 491 1118 591 1122
rect 595 1118 599 1122
rect 603 1118 711 1122
rect 715 1118 759 1122
rect 763 1118 831 1122
rect 835 1118 927 1122
rect 931 1118 967 1122
rect 971 1118 1095 1122
rect 1099 1118 1119 1122
rect 1123 1118 1247 1122
rect 1251 1118 1279 1122
rect 1283 1118 1399 1122
rect 1403 1118 1447 1122
rect 1451 1118 1543 1122
rect 1547 1118 1623 1122
rect 1627 1118 1687 1122
rect 1691 1118 1839 1122
rect 1843 1118 2007 1122
rect 2011 1118 2031 1122
rect 103 1117 2031 1118
rect 2037 1122 2047 1123
rect 2051 1122 2311 1126
rect 2315 1122 2407 1126
rect 2411 1122 2415 1126
rect 2419 1122 2503 1126
rect 2507 1122 2527 1126
rect 2531 1122 2599 1126
rect 2603 1122 2639 1126
rect 2643 1122 2695 1126
rect 2699 1122 2767 1126
rect 2771 1122 2807 1126
rect 2811 1122 2911 1126
rect 2915 1122 2943 1126
rect 2947 1122 3071 1126
rect 3075 1122 3095 1126
rect 3099 1122 3247 1126
rect 3251 1122 3263 1126
rect 3267 1122 3439 1126
rect 3443 1122 3447 1126
rect 3451 1122 3631 1126
rect 3635 1122 3639 1126
rect 3643 1122 3831 1126
rect 3835 1122 3839 1126
rect 3843 1122 3943 1126
rect 3947 1122 3986 1126
rect 2037 1121 3986 1122
rect 2037 1117 2038 1121
rect 84 1041 85 1047
rect 91 1046 2019 1047
rect 91 1042 111 1046
rect 115 1042 303 1046
rect 307 1042 375 1046
rect 379 1042 447 1046
rect 451 1042 487 1046
rect 491 1042 591 1046
rect 595 1042 599 1046
rect 603 1042 711 1046
rect 715 1042 727 1046
rect 731 1042 831 1046
rect 835 1042 855 1046
rect 859 1042 967 1046
rect 971 1042 975 1046
rect 979 1042 1087 1046
rect 1091 1042 1119 1046
rect 1123 1042 1199 1046
rect 1203 1042 1279 1046
rect 1283 1042 1311 1046
rect 1315 1042 1431 1046
rect 1435 1042 1447 1046
rect 1451 1042 1623 1046
rect 1627 1042 2007 1046
rect 2011 1042 2019 1046
rect 91 1041 2019 1042
rect 2025 1046 3974 1047
rect 2025 1042 2047 1046
rect 2051 1042 2407 1046
rect 2411 1042 2455 1046
rect 2459 1042 2503 1046
rect 2507 1042 2551 1046
rect 2555 1042 2599 1046
rect 2603 1042 2647 1046
rect 2651 1042 2695 1046
rect 2699 1042 2759 1046
rect 2763 1042 2807 1046
rect 2811 1042 2887 1046
rect 2891 1042 2943 1046
rect 2947 1042 3031 1046
rect 3035 1042 3095 1046
rect 3099 1042 3183 1046
rect 3187 1042 3263 1046
rect 3267 1042 3343 1046
rect 3347 1042 3447 1046
rect 3451 1042 3503 1046
rect 3507 1042 3639 1046
rect 3643 1042 3671 1046
rect 3675 1042 3839 1046
rect 3843 1042 3943 1046
rect 3947 1042 3974 1046
rect 2025 1041 3974 1042
rect 96 965 97 971
rect 103 970 2031 971
rect 103 966 111 970
rect 115 966 255 970
rect 259 966 303 970
rect 307 966 447 970
rect 451 966 591 970
rect 595 966 631 970
rect 635 966 727 970
rect 731 966 807 970
rect 811 966 855 970
rect 859 966 975 970
rect 979 966 1087 970
rect 1091 966 1127 970
rect 1131 966 1199 970
rect 1203 966 1271 970
rect 1275 966 1311 970
rect 1315 966 1415 970
rect 1419 966 1431 970
rect 1435 966 1551 970
rect 1555 966 1695 970
rect 1699 966 2007 970
rect 2011 966 2031 970
rect 103 965 2031 966
rect 2037 967 2038 971
rect 2037 966 3986 967
rect 2037 965 2047 966
rect 2030 962 2047 965
rect 2051 962 2423 966
rect 2427 962 2455 966
rect 2459 962 2519 966
rect 2523 962 2551 966
rect 2555 962 2615 966
rect 2619 962 2647 966
rect 2651 962 2711 966
rect 2715 962 2759 966
rect 2763 962 2823 966
rect 2827 962 2887 966
rect 2891 962 2951 966
rect 2955 962 3031 966
rect 3035 962 3103 966
rect 3107 962 3183 966
rect 3187 962 3271 966
rect 3275 962 3343 966
rect 3347 962 3455 966
rect 3459 962 3503 966
rect 3507 962 3647 966
rect 3651 962 3671 966
rect 3675 962 3839 966
rect 3843 962 3943 966
rect 3947 962 3986 966
rect 2030 961 3986 962
rect 84 885 85 891
rect 91 890 2019 891
rect 91 886 111 890
rect 115 886 255 890
rect 259 886 447 890
rect 451 886 631 890
rect 635 886 639 890
rect 643 886 807 890
rect 811 886 823 890
rect 827 886 975 890
rect 979 886 999 890
rect 1003 886 1127 890
rect 1131 886 1167 890
rect 1171 886 1271 890
rect 1275 886 1327 890
rect 1331 886 1415 890
rect 1419 886 1479 890
rect 1483 886 1551 890
rect 1555 886 1631 890
rect 1635 886 1695 890
rect 1699 886 1783 890
rect 1787 886 2007 890
rect 2011 886 2019 890
rect 91 885 2019 886
rect 2025 890 3974 891
rect 2025 886 2047 890
rect 2051 886 2343 890
rect 2347 886 2423 890
rect 2427 886 2439 890
rect 2443 886 2519 890
rect 2523 886 2535 890
rect 2539 886 2615 890
rect 2619 886 2631 890
rect 2635 886 2711 890
rect 2715 886 2735 890
rect 2739 886 2823 890
rect 2827 886 2863 890
rect 2867 886 2951 890
rect 2955 886 3015 890
rect 3019 886 3103 890
rect 3107 886 3191 890
rect 3195 886 3271 890
rect 3275 886 3391 890
rect 3395 886 3455 890
rect 3459 886 3607 890
rect 3611 886 3647 890
rect 3651 886 3823 890
rect 3827 886 3839 890
rect 3843 886 3943 890
rect 3947 886 3974 890
rect 2025 885 3974 886
rect 2030 814 3986 815
rect 2030 811 2047 814
rect 96 805 97 811
rect 103 810 2031 811
rect 103 806 111 810
rect 115 806 159 810
rect 163 806 255 810
rect 259 806 311 810
rect 315 806 447 810
rect 451 806 471 810
rect 475 806 623 810
rect 627 806 639 810
rect 643 806 775 810
rect 779 806 823 810
rect 827 806 935 810
rect 939 806 999 810
rect 1003 806 1095 810
rect 1099 806 1167 810
rect 1171 806 1255 810
rect 1259 806 1327 810
rect 1331 806 1415 810
rect 1419 806 1479 810
rect 1483 806 1583 810
rect 1587 806 1631 810
rect 1635 806 1751 810
rect 1755 806 1783 810
rect 1787 806 1903 810
rect 1907 806 2007 810
rect 2011 806 2031 810
rect 103 805 2031 806
rect 2037 810 2047 811
rect 2051 810 2311 814
rect 2315 810 2343 814
rect 2347 810 2439 814
rect 2443 810 2495 814
rect 2499 810 2535 814
rect 2539 810 2631 814
rect 2635 810 2687 814
rect 2691 810 2735 814
rect 2739 810 2863 814
rect 2867 810 2879 814
rect 2883 810 3015 814
rect 3019 810 3079 814
rect 3083 810 3191 814
rect 3195 810 3287 814
rect 3291 810 3391 814
rect 3395 810 3503 814
rect 3507 810 3607 814
rect 3611 810 3719 814
rect 3723 810 3823 814
rect 3827 810 3943 814
rect 3947 810 3986 814
rect 2037 809 3986 810
rect 2037 805 2038 809
rect 84 729 85 735
rect 91 734 2019 735
rect 91 730 111 734
rect 115 730 135 734
rect 139 730 159 734
rect 163 730 263 734
rect 267 730 311 734
rect 315 730 431 734
rect 435 730 471 734
rect 475 730 623 734
rect 627 730 775 734
rect 779 730 823 734
rect 827 730 935 734
rect 939 730 1015 734
rect 1019 730 1095 734
rect 1099 730 1207 734
rect 1211 730 1255 734
rect 1259 730 1391 734
rect 1395 730 1415 734
rect 1419 730 1567 734
rect 1571 730 1583 734
rect 1587 730 1743 734
rect 1747 730 1751 734
rect 1755 730 1903 734
rect 1907 730 2007 734
rect 2011 730 2019 734
rect 91 729 2019 730
rect 2025 734 3974 735
rect 2025 730 2047 734
rect 2051 730 2071 734
rect 2075 730 2255 734
rect 2259 730 2311 734
rect 2315 730 2455 734
rect 2459 730 2495 734
rect 2499 730 2655 734
rect 2659 730 2687 734
rect 2691 730 2855 734
rect 2859 730 2879 734
rect 2883 730 3047 734
rect 3051 730 3079 734
rect 3083 730 3239 734
rect 3243 730 3287 734
rect 3291 730 3439 734
rect 3443 730 3503 734
rect 3507 730 3639 734
rect 3643 730 3719 734
rect 3723 730 3839 734
rect 3843 730 3943 734
rect 3947 730 3974 734
rect 2025 729 3974 730
rect 96 653 97 659
rect 103 658 2031 659
rect 103 654 111 658
rect 115 654 135 658
rect 139 654 247 658
rect 251 654 263 658
rect 267 654 383 658
rect 387 654 431 658
rect 435 654 527 658
rect 531 654 623 658
rect 627 654 687 658
rect 691 654 823 658
rect 827 654 871 658
rect 875 654 1015 658
rect 1019 654 1079 658
rect 1083 654 1207 658
rect 1211 654 1303 658
rect 1307 654 1391 658
rect 1395 654 1543 658
rect 1547 654 1567 658
rect 1571 654 1743 658
rect 1747 654 1783 658
rect 1787 654 1903 658
rect 1907 654 2007 658
rect 2011 654 2031 658
rect 103 653 2031 654
rect 2037 658 3986 659
rect 2037 654 2047 658
rect 2051 654 2071 658
rect 2075 654 2231 658
rect 2235 654 2255 658
rect 2259 654 2431 658
rect 2435 654 2455 658
rect 2459 654 2631 658
rect 2635 654 2655 658
rect 2659 654 2831 658
rect 2835 654 2855 658
rect 2859 654 3023 658
rect 3027 654 3047 658
rect 3051 654 3207 658
rect 3211 654 3239 658
rect 3243 654 3375 658
rect 3379 654 3439 658
rect 3443 654 3535 658
rect 3539 654 3639 658
rect 3643 654 3695 658
rect 3699 654 3839 658
rect 3843 654 3943 658
rect 3947 654 3986 658
rect 2037 653 3986 654
rect 84 573 85 579
rect 91 578 2019 579
rect 91 574 111 578
rect 115 574 135 578
rect 139 574 247 578
rect 251 574 295 578
rect 299 574 383 578
rect 387 574 479 578
rect 483 574 527 578
rect 531 574 663 578
rect 667 574 687 578
rect 691 574 847 578
rect 851 574 871 578
rect 875 574 1031 578
rect 1035 574 1079 578
rect 1083 574 1215 578
rect 1219 574 1303 578
rect 1307 574 1399 578
rect 1403 574 1543 578
rect 1547 574 1591 578
rect 1595 574 1783 578
rect 1787 574 2007 578
rect 2011 574 2019 578
rect 91 573 2019 574
rect 2025 578 3974 579
rect 2025 574 2047 578
rect 2051 574 2071 578
rect 2075 574 2215 578
rect 2219 574 2231 578
rect 2235 574 2399 578
rect 2403 574 2431 578
rect 2435 574 2583 578
rect 2587 574 2631 578
rect 2635 574 2775 578
rect 2779 574 2831 578
rect 2835 574 2959 578
rect 2963 574 3023 578
rect 3027 574 3143 578
rect 3147 574 3207 578
rect 3211 574 3319 578
rect 3323 574 3375 578
rect 3379 574 3495 578
rect 3499 574 3535 578
rect 3539 574 3679 578
rect 3683 574 3695 578
rect 3699 574 3839 578
rect 3843 574 3943 578
rect 3947 574 3974 578
rect 2025 573 3974 574
rect 96 497 97 503
rect 103 502 2031 503
rect 103 498 111 502
rect 115 498 135 502
rect 139 498 287 502
rect 291 498 295 502
rect 299 498 455 502
rect 459 498 479 502
rect 483 498 615 502
rect 619 498 663 502
rect 667 498 767 502
rect 771 498 847 502
rect 851 498 903 502
rect 907 498 1031 502
rect 1035 498 1159 502
rect 1163 498 1215 502
rect 1219 498 1287 502
rect 1291 498 1399 502
rect 1403 498 1415 502
rect 1419 498 1591 502
rect 1595 498 1783 502
rect 1787 498 2007 502
rect 2011 498 2031 502
rect 103 497 2031 498
rect 2037 499 2038 503
rect 2037 498 3986 499
rect 2037 497 2047 498
rect 2030 494 2047 497
rect 2051 494 2071 498
rect 2075 494 2215 498
rect 2219 494 2223 498
rect 2227 494 2391 498
rect 2395 494 2399 498
rect 2403 494 2559 498
rect 2563 494 2583 498
rect 2587 494 2727 498
rect 2731 494 2775 498
rect 2779 494 2895 498
rect 2899 494 2959 498
rect 2963 494 3063 498
rect 3067 494 3143 498
rect 3147 494 3223 498
rect 3227 494 3319 498
rect 3323 494 3383 498
rect 3387 494 3495 498
rect 3499 494 3543 498
rect 3547 494 3679 498
rect 3683 494 3703 498
rect 3707 494 3839 498
rect 3843 494 3943 498
rect 3947 494 3986 498
rect 2030 493 3986 494
rect 84 421 85 427
rect 91 426 2019 427
rect 91 422 111 426
rect 115 422 135 426
rect 139 422 287 426
rect 291 422 447 426
rect 451 422 455 426
rect 459 422 599 426
rect 603 422 615 426
rect 619 422 751 426
rect 755 422 767 426
rect 771 422 903 426
rect 907 422 1031 426
rect 1035 422 1079 426
rect 1083 422 1159 426
rect 1163 422 1271 426
rect 1275 422 1287 426
rect 1291 422 1415 426
rect 1419 422 1479 426
rect 1483 422 1703 426
rect 1707 422 1903 426
rect 1907 422 2007 426
rect 2011 422 2019 426
rect 91 421 2019 422
rect 2025 423 2026 427
rect 2025 422 3974 423
rect 2025 421 2047 422
rect 2018 418 2047 421
rect 2051 418 2071 422
rect 2075 418 2223 422
rect 2227 418 2391 422
rect 2395 418 2463 422
rect 2467 418 2559 422
rect 2563 418 2655 422
rect 2659 418 2727 422
rect 2731 418 2751 422
rect 2755 418 2847 422
rect 2851 418 2895 422
rect 2899 418 2943 422
rect 2947 418 3039 422
rect 3043 418 3063 422
rect 3067 418 3135 422
rect 3139 418 3223 422
rect 3227 418 3231 422
rect 3235 418 3383 422
rect 3387 418 3543 422
rect 3547 418 3703 422
rect 3707 418 3839 422
rect 3843 418 3943 422
rect 3947 418 3974 422
rect 2018 417 3974 418
rect 96 341 97 347
rect 103 346 2031 347
rect 103 342 111 346
rect 115 342 135 346
rect 139 342 159 346
rect 163 342 287 346
rect 291 342 351 346
rect 355 342 447 346
rect 451 342 551 346
rect 555 342 599 346
rect 603 342 751 346
rect 755 342 759 346
rect 763 342 903 346
rect 907 342 959 346
rect 963 342 1079 346
rect 1083 342 1159 346
rect 1163 342 1271 346
rect 1275 342 1343 346
rect 1347 342 1479 346
rect 1483 342 1527 346
rect 1531 342 1703 346
rect 1707 342 1711 346
rect 1715 342 1895 346
rect 1899 342 1903 346
rect 1907 342 2007 346
rect 2011 342 2031 346
rect 103 341 2031 342
rect 2037 346 3986 347
rect 2037 342 2047 346
rect 2051 342 2399 346
rect 2403 342 2463 346
rect 2467 342 2503 346
rect 2507 342 2559 346
rect 2563 342 2623 346
rect 2627 342 2655 346
rect 2659 342 2751 346
rect 2755 342 2759 346
rect 2763 342 2847 346
rect 2851 342 2911 346
rect 2915 342 2943 346
rect 2947 342 3039 346
rect 3043 342 3071 346
rect 3075 342 3135 346
rect 3139 342 3231 346
rect 3235 342 3247 346
rect 3251 342 3423 346
rect 3427 342 3607 346
rect 3611 342 3791 346
rect 3795 342 3943 346
rect 3947 342 3986 346
rect 2037 341 3986 342
rect 2018 265 2019 271
rect 2025 270 3967 271
rect 2025 266 2047 270
rect 2051 266 2191 270
rect 2195 266 2351 270
rect 2355 266 2399 270
rect 2403 266 2503 270
rect 2507 266 2519 270
rect 2523 266 2623 270
rect 2627 266 2687 270
rect 2691 266 2759 270
rect 2763 266 2855 270
rect 2859 266 2911 270
rect 2915 266 3031 270
rect 3035 266 3071 270
rect 3075 266 3215 270
rect 3219 266 3247 270
rect 3251 266 3407 270
rect 3411 266 3423 270
rect 3427 266 3607 270
rect 3611 266 3791 270
rect 3795 266 3807 270
rect 3811 266 3943 270
rect 3947 266 3967 270
rect 2025 265 3967 266
rect 3973 265 3974 271
rect 2018 263 2026 265
rect 84 257 85 263
rect 91 262 2019 263
rect 91 258 111 262
rect 115 258 159 262
rect 163 258 223 262
rect 227 258 351 262
rect 355 258 383 262
rect 387 258 543 262
rect 547 258 551 262
rect 555 258 703 262
rect 707 258 759 262
rect 763 258 863 262
rect 867 258 959 262
rect 963 258 1031 262
rect 1035 258 1159 262
rect 1163 258 1199 262
rect 1203 258 1343 262
rect 1347 258 1367 262
rect 1371 258 1527 262
rect 1531 258 1543 262
rect 1547 258 1711 262
rect 1715 258 1727 262
rect 1731 258 1895 262
rect 1899 258 1903 262
rect 1907 258 2007 262
rect 2011 258 2019 262
rect 91 257 2019 258
rect 2025 257 2026 263
rect 96 161 97 167
rect 103 166 2031 167
rect 103 162 111 166
rect 115 162 135 166
rect 139 162 223 166
rect 227 162 231 166
rect 235 162 327 166
rect 331 162 383 166
rect 387 162 423 166
rect 427 162 527 166
rect 531 162 543 166
rect 547 162 647 166
rect 651 162 703 166
rect 707 162 775 166
rect 779 162 863 166
rect 867 162 903 166
rect 907 162 1031 166
rect 1035 162 1151 166
rect 1155 162 1199 166
rect 1203 162 1271 166
rect 1275 162 1367 166
rect 1371 162 1383 166
rect 1387 162 1487 166
rect 1491 162 1543 166
rect 1547 162 1591 166
rect 1595 162 1703 166
rect 1707 162 1727 166
rect 1731 162 1807 166
rect 1811 162 1903 166
rect 1907 162 2007 166
rect 2011 162 2031 166
rect 103 161 2031 162
rect 2037 163 2038 167
rect 2037 162 3986 163
rect 2037 161 2047 162
rect 2030 158 2047 161
rect 2051 158 2071 162
rect 2075 158 2167 162
rect 2171 158 2191 162
rect 2195 158 2263 162
rect 2267 158 2351 162
rect 2355 158 2367 162
rect 2371 158 2487 162
rect 2491 158 2519 162
rect 2523 158 2615 162
rect 2619 158 2687 162
rect 2691 158 2743 162
rect 2747 158 2855 162
rect 2859 158 2871 162
rect 2875 158 2991 162
rect 2995 158 3031 162
rect 3035 158 3111 162
rect 3115 158 3215 162
rect 3219 158 3223 162
rect 3227 158 3327 162
rect 3331 158 3407 162
rect 3411 158 3431 162
rect 3435 158 3535 162
rect 3539 158 3607 162
rect 3611 158 3639 162
rect 3643 158 3743 162
rect 3747 158 3807 162
rect 3811 158 3839 162
rect 3843 158 3943 162
rect 3947 158 3986 162
rect 2030 157 3986 158
rect 84 85 85 91
rect 91 90 2019 91
rect 91 86 111 90
rect 115 86 135 90
rect 139 86 231 90
rect 235 86 327 90
rect 331 86 423 90
rect 427 86 527 90
rect 531 86 647 90
rect 651 86 775 90
rect 779 86 903 90
rect 907 86 1031 90
rect 1035 86 1151 90
rect 1155 86 1271 90
rect 1275 86 1383 90
rect 1387 86 1487 90
rect 1491 86 1591 90
rect 1595 86 1703 90
rect 1707 86 1807 90
rect 1811 86 1903 90
rect 1907 86 2007 90
rect 2011 86 2019 90
rect 91 85 2019 86
rect 2025 87 2026 91
rect 2025 86 3974 87
rect 2025 85 2047 86
rect 2018 82 2047 85
rect 2051 82 2071 86
rect 2075 82 2167 86
rect 2171 82 2263 86
rect 2267 82 2367 86
rect 2371 82 2487 86
rect 2491 82 2615 86
rect 2619 82 2743 86
rect 2747 82 2871 86
rect 2875 82 2991 86
rect 2995 82 3111 86
rect 3115 82 3223 86
rect 3227 82 3327 86
rect 3331 82 3431 86
rect 3435 82 3535 86
rect 3539 82 3639 86
rect 3643 82 3743 86
rect 3747 82 3839 86
rect 3843 82 3943 86
rect 3947 82 3974 86
rect 2018 81 3974 82
<< m5c >>
rect 2031 4025 2037 4031
rect 3979 4025 3985 4031
rect 97 4005 103 4011
rect 2031 4005 2037 4011
rect 2019 3949 2025 3955
rect 3967 3949 3973 3955
rect 85 3929 91 3935
rect 2019 3929 2025 3935
rect 2031 3873 2037 3879
rect 3979 3873 3985 3879
rect 97 3849 103 3855
rect 2031 3849 2037 3855
rect 2019 3797 2025 3803
rect 3967 3797 3973 3803
rect 85 3769 91 3775
rect 2019 3769 2025 3775
rect 2031 3709 2037 3715
rect 3979 3709 3985 3715
rect 97 3681 103 3687
rect 2031 3681 2037 3687
rect 2019 3629 2025 3635
rect 3967 3629 3973 3635
rect 85 3597 91 3603
rect 2019 3597 2025 3603
rect 2031 3537 2037 3543
rect 3979 3537 3985 3543
rect 97 3513 103 3519
rect 2031 3513 2037 3519
rect 2019 3461 2025 3467
rect 3967 3461 3973 3467
rect 85 3429 91 3435
rect 2019 3429 2025 3435
rect 2031 3377 2037 3383
rect 3979 3377 3985 3383
rect 97 3345 103 3351
rect 2031 3345 2037 3351
rect 2019 3297 2025 3303
rect 3967 3297 3973 3303
rect 85 3261 91 3267
rect 2019 3261 2025 3267
rect 2031 3221 2037 3227
rect 3979 3221 3985 3227
rect 97 3185 103 3191
rect 2031 3185 2037 3191
rect 2019 3141 2025 3147
rect 3967 3141 3973 3147
rect 85 3109 91 3115
rect 2019 3109 2025 3115
rect 2031 3061 2037 3067
rect 3979 3061 3985 3067
rect 97 3033 103 3039
rect 2031 3033 2037 3039
rect 2019 2981 2025 2987
rect 3967 2981 3973 2987
rect 85 2933 91 2939
rect 2019 2933 2025 2939
rect 2031 2889 2037 2895
rect 3979 2889 3985 2895
rect 97 2849 103 2855
rect 2031 2849 2037 2855
rect 2019 2813 2025 2819
rect 3967 2813 3973 2819
rect 85 2773 91 2779
rect 2019 2773 2025 2779
rect 2031 2729 2037 2735
rect 3979 2729 3985 2735
rect 97 2697 103 2703
rect 2031 2697 2037 2703
rect 2019 2649 2025 2655
rect 3967 2649 3973 2655
rect 85 2621 91 2627
rect 2019 2621 2025 2627
rect 2031 2565 2037 2571
rect 3979 2565 3985 2571
rect 97 2541 103 2547
rect 2031 2541 2037 2547
rect 2019 2485 2025 2491
rect 3967 2485 3973 2491
rect 85 2461 91 2467
rect 2019 2461 2025 2467
rect 2031 2393 2037 2399
rect 3979 2393 3985 2399
rect 97 2385 103 2391
rect 2031 2385 2037 2391
rect 2019 2317 2025 2323
rect 3967 2317 3973 2323
rect 85 2301 91 2307
rect 2019 2301 2025 2307
rect 2031 2233 2037 2239
rect 3979 2233 3985 2239
rect 97 2225 103 2231
rect 2031 2225 2037 2231
rect 85 2149 91 2155
rect 2019 2149 2025 2155
rect 97 2065 103 2071
rect 2031 2065 2037 2071
rect 85 1981 91 1987
rect 2019 1981 2025 1987
rect 97 1897 103 1903
rect 2031 1897 2037 1903
rect 85 1821 91 1827
rect 2019 1821 2025 1827
rect 97 1745 103 1751
rect 2031 1745 2037 1751
rect 2019 1673 2025 1679
rect 3967 1673 3973 1679
rect 85 1665 91 1671
rect 2019 1665 2025 1671
rect 97 1589 103 1595
rect 2031 1589 2037 1595
rect 85 1509 91 1515
rect 2019 1509 2025 1515
rect 97 1433 103 1439
rect 2031 1433 2037 1439
rect 85 1353 91 1359
rect 2019 1353 2025 1359
rect 97 1273 103 1279
rect 2031 1273 2037 1279
rect 85 1197 91 1203
rect 2019 1197 2025 1203
rect 97 1117 103 1123
rect 2031 1117 2037 1123
rect 85 1041 91 1047
rect 2019 1041 2025 1047
rect 97 965 103 971
rect 2031 965 2037 971
rect 85 885 91 891
rect 2019 885 2025 891
rect 97 805 103 811
rect 2031 805 2037 811
rect 85 729 91 735
rect 2019 729 2025 735
rect 97 653 103 659
rect 2031 653 2037 659
rect 85 573 91 579
rect 2019 573 2025 579
rect 97 497 103 503
rect 2031 497 2037 503
rect 85 421 91 427
rect 2019 421 2025 427
rect 97 341 103 347
rect 2031 341 2037 347
rect 2019 265 2025 271
rect 3967 265 3973 271
rect 85 257 91 263
rect 2019 257 2025 263
rect 97 161 103 167
rect 2031 161 2037 167
rect 85 85 91 91
rect 2019 85 2025 91
<< m5 >>
rect 84 3935 92 4032
rect 84 3929 85 3935
rect 91 3929 92 3935
rect 84 3775 92 3929
rect 84 3769 85 3775
rect 91 3769 92 3775
rect 84 3603 92 3769
rect 84 3597 85 3603
rect 91 3597 92 3603
rect 84 3435 92 3597
rect 84 3429 85 3435
rect 91 3429 92 3435
rect 84 3267 92 3429
rect 84 3261 85 3267
rect 91 3261 92 3267
rect 84 3115 92 3261
rect 84 3109 85 3115
rect 91 3109 92 3115
rect 84 2939 92 3109
rect 84 2933 85 2939
rect 91 2933 92 2939
rect 84 2779 92 2933
rect 84 2773 85 2779
rect 91 2773 92 2779
rect 84 2627 92 2773
rect 84 2621 85 2627
rect 91 2621 92 2627
rect 84 2467 92 2621
rect 84 2461 85 2467
rect 91 2461 92 2467
rect 84 2307 92 2461
rect 84 2301 85 2307
rect 91 2301 92 2307
rect 84 2155 92 2301
rect 84 2149 85 2155
rect 91 2149 92 2155
rect 84 1987 92 2149
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1827 92 1981
rect 84 1821 85 1827
rect 91 1821 92 1827
rect 84 1671 92 1821
rect 84 1665 85 1671
rect 91 1665 92 1671
rect 84 1515 92 1665
rect 84 1509 85 1515
rect 91 1509 92 1515
rect 84 1359 92 1509
rect 84 1353 85 1359
rect 91 1353 92 1359
rect 84 1203 92 1353
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1047 92 1197
rect 84 1041 85 1047
rect 91 1041 92 1047
rect 84 891 92 1041
rect 84 885 85 891
rect 91 885 92 891
rect 84 735 92 885
rect 84 729 85 735
rect 91 729 92 735
rect 84 579 92 729
rect 84 573 85 579
rect 91 573 92 579
rect 84 427 92 573
rect 84 421 85 427
rect 91 421 92 427
rect 84 263 92 421
rect 84 257 85 263
rect 91 257 92 263
rect 84 91 92 257
rect 84 85 85 91
rect 91 85 92 91
rect 84 72 92 85
rect 96 4011 104 4032
rect 96 4005 97 4011
rect 103 4005 104 4011
rect 96 3855 104 4005
rect 96 3849 97 3855
rect 103 3849 104 3855
rect 96 3687 104 3849
rect 96 3681 97 3687
rect 103 3681 104 3687
rect 96 3519 104 3681
rect 96 3513 97 3519
rect 103 3513 104 3519
rect 96 3351 104 3513
rect 96 3345 97 3351
rect 103 3345 104 3351
rect 96 3191 104 3345
rect 96 3185 97 3191
rect 103 3185 104 3191
rect 96 3039 104 3185
rect 96 3033 97 3039
rect 103 3033 104 3039
rect 96 2855 104 3033
rect 96 2849 97 2855
rect 103 2849 104 2855
rect 96 2703 104 2849
rect 96 2697 97 2703
rect 103 2697 104 2703
rect 96 2547 104 2697
rect 96 2541 97 2547
rect 103 2541 104 2547
rect 96 2391 104 2541
rect 96 2385 97 2391
rect 103 2385 104 2391
rect 96 2231 104 2385
rect 96 2225 97 2231
rect 103 2225 104 2231
rect 96 2071 104 2225
rect 96 2065 97 2071
rect 103 2065 104 2071
rect 96 1903 104 2065
rect 96 1897 97 1903
rect 103 1897 104 1903
rect 96 1751 104 1897
rect 96 1745 97 1751
rect 103 1745 104 1751
rect 96 1595 104 1745
rect 96 1589 97 1595
rect 103 1589 104 1595
rect 96 1439 104 1589
rect 96 1433 97 1439
rect 103 1433 104 1439
rect 96 1279 104 1433
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1123 104 1273
rect 96 1117 97 1123
rect 103 1117 104 1123
rect 96 971 104 1117
rect 96 965 97 971
rect 103 965 104 971
rect 96 811 104 965
rect 96 805 97 811
rect 103 805 104 811
rect 96 659 104 805
rect 96 653 97 659
rect 103 653 104 659
rect 96 503 104 653
rect 96 497 97 503
rect 103 497 104 503
rect 96 347 104 497
rect 96 341 97 347
rect 103 341 104 347
rect 96 167 104 341
rect 96 161 97 167
rect 103 161 104 167
rect 96 72 104 161
rect 2018 3955 2026 4032
rect 2018 3949 2019 3955
rect 2025 3949 2026 3955
rect 2018 3935 2026 3949
rect 2018 3929 2019 3935
rect 2025 3929 2026 3935
rect 2018 3803 2026 3929
rect 2018 3797 2019 3803
rect 2025 3797 2026 3803
rect 2018 3775 2026 3797
rect 2018 3769 2019 3775
rect 2025 3769 2026 3775
rect 2018 3635 2026 3769
rect 2018 3629 2019 3635
rect 2025 3629 2026 3635
rect 2018 3603 2026 3629
rect 2018 3597 2019 3603
rect 2025 3597 2026 3603
rect 2018 3467 2026 3597
rect 2018 3461 2019 3467
rect 2025 3461 2026 3467
rect 2018 3435 2026 3461
rect 2018 3429 2019 3435
rect 2025 3429 2026 3435
rect 2018 3303 2026 3429
rect 2018 3297 2019 3303
rect 2025 3297 2026 3303
rect 2018 3267 2026 3297
rect 2018 3261 2019 3267
rect 2025 3261 2026 3267
rect 2018 3147 2026 3261
rect 2018 3141 2019 3147
rect 2025 3141 2026 3147
rect 2018 3115 2026 3141
rect 2018 3109 2019 3115
rect 2025 3109 2026 3115
rect 2018 2987 2026 3109
rect 2018 2981 2019 2987
rect 2025 2981 2026 2987
rect 2018 2939 2026 2981
rect 2018 2933 2019 2939
rect 2025 2933 2026 2939
rect 2018 2819 2026 2933
rect 2018 2813 2019 2819
rect 2025 2813 2026 2819
rect 2018 2779 2026 2813
rect 2018 2773 2019 2779
rect 2025 2773 2026 2779
rect 2018 2655 2026 2773
rect 2018 2649 2019 2655
rect 2025 2649 2026 2655
rect 2018 2627 2026 2649
rect 2018 2621 2019 2627
rect 2025 2621 2026 2627
rect 2018 2491 2026 2621
rect 2018 2485 2019 2491
rect 2025 2485 2026 2491
rect 2018 2467 2026 2485
rect 2018 2461 2019 2467
rect 2025 2461 2026 2467
rect 2018 2323 2026 2461
rect 2018 2317 2019 2323
rect 2025 2317 2026 2323
rect 2018 2307 2026 2317
rect 2018 2301 2019 2307
rect 2025 2301 2026 2307
rect 2018 2155 2026 2301
rect 2018 2149 2019 2155
rect 2025 2149 2026 2155
rect 2018 1987 2026 2149
rect 2018 1981 2019 1987
rect 2025 1981 2026 1987
rect 2018 1827 2026 1981
rect 2018 1821 2019 1827
rect 2025 1821 2026 1827
rect 2018 1679 2026 1821
rect 2018 1673 2019 1679
rect 2025 1673 2026 1679
rect 2018 1671 2026 1673
rect 2018 1665 2019 1671
rect 2025 1665 2026 1671
rect 2018 1515 2026 1665
rect 2018 1509 2019 1515
rect 2025 1509 2026 1515
rect 2018 1359 2026 1509
rect 2018 1353 2019 1359
rect 2025 1353 2026 1359
rect 2018 1203 2026 1353
rect 2018 1197 2019 1203
rect 2025 1197 2026 1203
rect 2018 1047 2026 1197
rect 2018 1041 2019 1047
rect 2025 1041 2026 1047
rect 2018 891 2026 1041
rect 2018 885 2019 891
rect 2025 885 2026 891
rect 2018 735 2026 885
rect 2018 729 2019 735
rect 2025 729 2026 735
rect 2018 579 2026 729
rect 2018 573 2019 579
rect 2025 573 2026 579
rect 2018 427 2026 573
rect 2018 421 2019 427
rect 2025 421 2026 427
rect 2018 271 2026 421
rect 2018 265 2019 271
rect 2025 265 2026 271
rect 2018 263 2026 265
rect 2018 257 2019 263
rect 2025 257 2026 263
rect 2018 91 2026 257
rect 2018 85 2019 91
rect 2025 85 2026 91
rect 2018 72 2026 85
rect 2030 4031 2038 4032
rect 2030 4025 2031 4031
rect 2037 4025 2038 4031
rect 2030 4011 2038 4025
rect 2030 4005 2031 4011
rect 2037 4005 2038 4011
rect 2030 3879 2038 4005
rect 2030 3873 2031 3879
rect 2037 3873 2038 3879
rect 2030 3855 2038 3873
rect 2030 3849 2031 3855
rect 2037 3849 2038 3855
rect 2030 3715 2038 3849
rect 2030 3709 2031 3715
rect 2037 3709 2038 3715
rect 2030 3687 2038 3709
rect 2030 3681 2031 3687
rect 2037 3681 2038 3687
rect 2030 3543 2038 3681
rect 2030 3537 2031 3543
rect 2037 3537 2038 3543
rect 2030 3519 2038 3537
rect 2030 3513 2031 3519
rect 2037 3513 2038 3519
rect 2030 3383 2038 3513
rect 2030 3377 2031 3383
rect 2037 3377 2038 3383
rect 2030 3351 2038 3377
rect 2030 3345 2031 3351
rect 2037 3345 2038 3351
rect 2030 3227 2038 3345
rect 2030 3221 2031 3227
rect 2037 3221 2038 3227
rect 2030 3191 2038 3221
rect 2030 3185 2031 3191
rect 2037 3185 2038 3191
rect 2030 3067 2038 3185
rect 2030 3061 2031 3067
rect 2037 3061 2038 3067
rect 2030 3039 2038 3061
rect 2030 3033 2031 3039
rect 2037 3033 2038 3039
rect 2030 2895 2038 3033
rect 2030 2889 2031 2895
rect 2037 2889 2038 2895
rect 2030 2855 2038 2889
rect 2030 2849 2031 2855
rect 2037 2849 2038 2855
rect 2030 2735 2038 2849
rect 2030 2729 2031 2735
rect 2037 2729 2038 2735
rect 2030 2703 2038 2729
rect 2030 2697 2031 2703
rect 2037 2697 2038 2703
rect 2030 2571 2038 2697
rect 2030 2565 2031 2571
rect 2037 2565 2038 2571
rect 2030 2547 2038 2565
rect 2030 2541 2031 2547
rect 2037 2541 2038 2547
rect 2030 2399 2038 2541
rect 2030 2393 2031 2399
rect 2037 2393 2038 2399
rect 2030 2391 2038 2393
rect 2030 2385 2031 2391
rect 2037 2385 2038 2391
rect 2030 2239 2038 2385
rect 2030 2233 2031 2239
rect 2037 2233 2038 2239
rect 2030 2231 2038 2233
rect 2030 2225 2031 2231
rect 2037 2225 2038 2231
rect 2030 2071 2038 2225
rect 2030 2065 2031 2071
rect 2037 2065 2038 2071
rect 2030 1903 2038 2065
rect 2030 1897 2031 1903
rect 2037 1897 2038 1903
rect 2030 1751 2038 1897
rect 2030 1745 2031 1751
rect 2037 1745 2038 1751
rect 2030 1595 2038 1745
rect 2030 1589 2031 1595
rect 2037 1589 2038 1595
rect 2030 1439 2038 1589
rect 2030 1433 2031 1439
rect 2037 1433 2038 1439
rect 2030 1279 2038 1433
rect 2030 1273 2031 1279
rect 2037 1273 2038 1279
rect 2030 1123 2038 1273
rect 2030 1117 2031 1123
rect 2037 1117 2038 1123
rect 2030 971 2038 1117
rect 2030 965 2031 971
rect 2037 965 2038 971
rect 2030 811 2038 965
rect 2030 805 2031 811
rect 2037 805 2038 811
rect 2030 659 2038 805
rect 2030 653 2031 659
rect 2037 653 2038 659
rect 2030 503 2038 653
rect 2030 497 2031 503
rect 2037 497 2038 503
rect 2030 347 2038 497
rect 2030 341 2031 347
rect 2037 341 2038 347
rect 2030 167 2038 341
rect 2030 161 2031 167
rect 2037 161 2038 167
rect 2030 72 2038 161
rect 3966 3955 3974 4032
rect 3966 3949 3967 3955
rect 3973 3949 3974 3955
rect 3966 3803 3974 3949
rect 3966 3797 3967 3803
rect 3973 3797 3974 3803
rect 3966 3635 3974 3797
rect 3966 3629 3967 3635
rect 3973 3629 3974 3635
rect 3966 3467 3974 3629
rect 3966 3461 3967 3467
rect 3973 3461 3974 3467
rect 3966 3303 3974 3461
rect 3966 3297 3967 3303
rect 3973 3297 3974 3303
rect 3966 3147 3974 3297
rect 3966 3141 3967 3147
rect 3973 3141 3974 3147
rect 3966 2987 3974 3141
rect 3966 2981 3967 2987
rect 3973 2981 3974 2987
rect 3966 2819 3974 2981
rect 3966 2813 3967 2819
rect 3973 2813 3974 2819
rect 3966 2655 3974 2813
rect 3966 2649 3967 2655
rect 3973 2649 3974 2655
rect 3966 2491 3974 2649
rect 3966 2485 3967 2491
rect 3973 2485 3974 2491
rect 3966 2323 3974 2485
rect 3966 2317 3967 2323
rect 3973 2317 3974 2323
rect 3966 1679 3974 2317
rect 3966 1673 3967 1679
rect 3973 1673 3974 1679
rect 3966 271 3974 1673
rect 3966 265 3967 271
rect 3973 265 3974 271
rect 3966 72 3974 265
rect 3978 4031 3986 4032
rect 3978 4025 3979 4031
rect 3985 4025 3986 4031
rect 3978 3879 3986 4025
rect 3978 3873 3979 3879
rect 3985 3873 3986 3879
rect 3978 3715 3986 3873
rect 3978 3709 3979 3715
rect 3985 3709 3986 3715
rect 3978 3543 3986 3709
rect 3978 3537 3979 3543
rect 3985 3537 3986 3543
rect 3978 3383 3986 3537
rect 3978 3377 3979 3383
rect 3985 3377 3986 3383
rect 3978 3227 3986 3377
rect 3978 3221 3979 3227
rect 3985 3221 3986 3227
rect 3978 3067 3986 3221
rect 3978 3061 3979 3067
rect 3985 3061 3986 3067
rect 3978 2895 3986 3061
rect 3978 2889 3979 2895
rect 3985 2889 3986 2895
rect 3978 2735 3986 2889
rect 3978 2729 3979 2735
rect 3985 2729 3986 2735
rect 3978 2571 3986 2729
rect 3978 2565 3979 2571
rect 3985 2565 3986 2571
rect 3978 2399 3986 2565
rect 3978 2393 3979 2399
rect 3985 2393 3986 2399
rect 3978 2239 3986 2393
rect 3978 2233 3979 2239
rect 3985 2233 3986 2239
rect 3978 72 3986 2233
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__195
timestamp 1731220342
transform 1 0 3936 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220342
transform 1 0 2040 0 1 3980
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220342
transform 1 0 3936 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220342
transform 1 0 2040 0 -1 3924
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220342
transform 1 0 3936 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220342
transform 1 0 2040 0 1 3828
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220342
transform 1 0 3936 0 -1 3772
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220342
transform 1 0 2040 0 -1 3772
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220342
transform 1 0 3936 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220342
transform 1 0 2040 0 1 3664
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220342
transform 1 0 3936 0 -1 3604
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220342
transform 1 0 2040 0 -1 3604
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220342
transform 1 0 3936 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220342
transform 1 0 2040 0 1 3492
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220342
transform 1 0 3936 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220342
transform 1 0 2040 0 -1 3436
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220342
transform 1 0 3936 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220342
transform 1 0 2040 0 1 3332
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220342
transform 1 0 3936 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220342
transform 1 0 2040 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220342
transform 1 0 3936 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220342
transform 1 0 2040 0 1 3176
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220342
transform 1 0 3936 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220342
transform 1 0 2040 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220342
transform 1 0 3936 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220342
transform 1 0 2040 0 1 3016
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220342
transform 1 0 3936 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220342
transform 1 0 2040 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220342
transform 1 0 3936 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220342
transform 1 0 2040 0 1 2844
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220342
transform 1 0 3936 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220342
transform 1 0 2040 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220342
transform 1 0 3936 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220342
transform 1 0 2040 0 1 2684
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220342
transform 1 0 3936 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220342
transform 1 0 2040 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220342
transform 1 0 3936 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220342
transform 1 0 2040 0 1 2520
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220342
transform 1 0 3936 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220342
transform 1 0 2040 0 -1 2460
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220342
transform 1 0 3936 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220342
transform 1 0 2040 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220342
transform 1 0 3936 0 -1 2292
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220342
transform 1 0 2040 0 -1 2292
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220342
transform 1 0 3936 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220342
transform 1 0 2040 0 1 2188
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220342
transform 1 0 3936 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220342
transform 1 0 2040 0 -1 2120
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220342
transform 1 0 3936 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220342
transform 1 0 2040 0 1 2016
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220342
transform 1 0 3936 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220342
transform 1 0 2040 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220342
transform 1 0 3936 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220342
transform 1 0 2040 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220342
transform 1 0 3936 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220342
transform 1 0 2040 0 -1 1800
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220342
transform 1 0 3936 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220342
transform 1 0 2040 0 1 1704
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220342
transform 1 0 3936 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220342
transform 1 0 2040 0 -1 1648
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220342
transform 1 0 3936 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220342
transform 1 0 2040 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220342
transform 1 0 3936 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220342
transform 1 0 2040 0 -1 1488
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220342
transform 1 0 3936 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220342
transform 1 0 2040 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220342
transform 1 0 3936 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220342
transform 1 0 2040 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220342
transform 1 0 3936 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220342
transform 1 0 2040 0 1 1232
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220342
transform 1 0 3936 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220342
transform 1 0 2040 0 -1 1176
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220342
transform 1 0 3936 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220342
transform 1 0 2040 0 1 1076
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220342
transform 1 0 3936 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220342
transform 1 0 2040 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220342
transform 1 0 3936 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220342
transform 1 0 2040 0 1 916
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220342
transform 1 0 3936 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220342
transform 1 0 2040 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220342
transform 1 0 3936 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220342
transform 1 0 2040 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220342
transform 1 0 3936 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220342
transform 1 0 2040 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220342
transform 1 0 3936 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220342
transform 1 0 2040 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220342
transform 1 0 3936 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220342
transform 1 0 2040 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220342
transform 1 0 3936 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220342
transform 1 0 2040 0 1 448
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220342
transform 1 0 3936 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220342
transform 1 0 2040 0 -1 392
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220342
transform 1 0 3936 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220342
transform 1 0 2040 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220342
transform 1 0 3936 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220342
transform 1 0 2040 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220342
transform 1 0 3936 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220342
transform 1 0 2040 0 1 112
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220342
transform 1 0 2000 0 1 3960
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220342
transform 1 0 104 0 1 3960
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220342
transform 1 0 2000 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220342
transform 1 0 104 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220342
transform 1 0 2000 0 1 3804
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220342
transform 1 0 104 0 1 3804
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220342
transform 1 0 2000 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220342
transform 1 0 104 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220342
transform 1 0 2000 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220342
transform 1 0 104 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220342
transform 1 0 2000 0 -1 3572
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220342
transform 1 0 104 0 -1 3572
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220342
transform 1 0 2000 0 1 3468
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220342
transform 1 0 104 0 1 3468
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220342
transform 1 0 2000 0 -1 3404
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220342
transform 1 0 104 0 -1 3404
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220342
transform 1 0 2000 0 1 3300
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220342
transform 1 0 104 0 1 3300
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220342
transform 1 0 2000 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220342
transform 1 0 104 0 -1 3236
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220342
transform 1 0 2000 0 1 3140
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220342
transform 1 0 104 0 1 3140
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220342
transform 1 0 2000 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220342
transform 1 0 104 0 -1 3084
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220342
transform 1 0 2000 0 1 2988
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220342
transform 1 0 104 0 1 2988
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220342
transform 1 0 2000 0 -1 2908
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220342
transform 1 0 104 0 -1 2908
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220342
transform 1 0 2000 0 1 2804
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220342
transform 1 0 104 0 1 2804
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220342
transform 1 0 2000 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220342
transform 1 0 104 0 -1 2748
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220342
transform 1 0 2000 0 1 2652
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220342
transform 1 0 104 0 1 2652
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220342
transform 1 0 2000 0 -1 2596
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220342
transform 1 0 104 0 -1 2596
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220342
transform 1 0 2000 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220342
transform 1 0 104 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220342
transform 1 0 2000 0 -1 2436
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220342
transform 1 0 104 0 -1 2436
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220342
transform 1 0 2000 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220342
transform 1 0 104 0 1 2340
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220342
transform 1 0 2000 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220342
transform 1 0 104 0 -1 2276
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220342
transform 1 0 2000 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220342
transform 1 0 104 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220342
transform 1 0 2000 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220342
transform 1 0 104 0 -1 2124
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220342
transform 1 0 2000 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220342
transform 1 0 104 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220342
transform 1 0 2000 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220342
transform 1 0 104 0 -1 1956
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220342
transform 1 0 2000 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220342
transform 1 0 104 0 1 1852
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220342
transform 1 0 2000 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220342
transform 1 0 104 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220342
transform 1 0 2000 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220342
transform 1 0 104 0 1 1700
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220342
transform 1 0 2000 0 -1 1640
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220342
transform 1 0 104 0 -1 1640
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220342
transform 1 0 2000 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220342
transform 1 0 104 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220342
transform 1 0 2000 0 -1 1484
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220342
transform 1 0 104 0 -1 1484
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220342
transform 1 0 2000 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220342
transform 1 0 104 0 1 1388
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220342
transform 1 0 2000 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220342
transform 1 0 104 0 -1 1328
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220342
transform 1 0 2000 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220342
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220342
transform 1 0 2000 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220342
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220342
transform 1 0 2000 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220342
transform 1 0 104 0 1 1072
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220342
transform 1 0 2000 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220342
transform 1 0 104 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220342
transform 1 0 2000 0 1 920
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220342
transform 1 0 104 0 1 920
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220342
transform 1 0 2000 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220342
transform 1 0 104 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220342
transform 1 0 2000 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220342
transform 1 0 104 0 1 760
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220342
transform 1 0 2000 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220342
transform 1 0 104 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220342
transform 1 0 2000 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220342
transform 1 0 104 0 1 608
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220342
transform 1 0 2000 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220342
transform 1 0 104 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220342
transform 1 0 2000 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220342
transform 1 0 104 0 1 452
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220342
transform 1 0 2000 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220342
transform 1 0 104 0 -1 396
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220342
transform 1 0 2000 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220342
transform 1 0 104 0 1 296
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220342
transform 1 0 2000 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220342
transform 1 0 104 0 -1 232
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220342
transform 1 0 2000 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220342
transform 1 0 104 0 1 116
box 7 3 12 24
use _0_0cell_0_0gcelem3x0  tst_5999_6
timestamp 1731220342
transform 1 0 3832 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5998_6
timestamp 1731220342
transform 1 0 3736 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5997_6
timestamp 1731220342
transform 1 0 3800 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5996_6
timestamp 1731220342
transform 1 0 3784 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5995_6
timestamp 1731220342
transform 1 0 3600 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5994_6
timestamp 1731220342
transform 1 0 3416 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5993_6
timestamp 1731220342
transform 1 0 3600 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5992_6
timestamp 1731220342
transform 1 0 3632 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5991_6
timestamp 1731220342
transform 1 0 3528 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5990_6
timestamp 1731220342
transform 1 0 3424 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5989_6
timestamp 1731220342
transform 1 0 3320 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5988_6
timestamp 1731220342
transform 1 0 3216 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5987_6
timestamp 1731220342
transform 1 0 3104 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5986_6
timestamp 1731220342
transform 1 0 2984 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5985_6
timestamp 1731220342
transform 1 0 2864 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5984_6
timestamp 1731220342
transform 1 0 3400 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5983_6
timestamp 1731220342
transform 1 0 3208 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5982_6
timestamp 1731220342
transform 1 0 3024 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5981_6
timestamp 1731220342
transform 1 0 2848 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5980_6
timestamp 1731220342
transform 1 0 3064 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5979_6
timestamp 1731220342
transform 1 0 3240 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5978_6
timestamp 1731220342
transform 1 0 3224 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5977_6
timestamp 1731220342
transform 1 0 3128 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5976_6
timestamp 1731220342
transform 1 0 3032 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5975_6
timestamp 1731220342
transform 1 0 2936 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5974_6
timestamp 1731220342
transform 1 0 2840 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5973_6
timestamp 1731220342
transform 1 0 2888 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5972_6
timestamp 1731220342
transform 1 0 3056 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5971_6
timestamp 1731220342
transform 1 0 3376 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5970_6
timestamp 1731220342
transform 1 0 3216 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5969_6
timestamp 1731220342
transform 1 0 3136 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5968_6
timestamp 1731220342
transform 1 0 2952 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5967_6
timestamp 1731220342
transform 1 0 3312 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5966_6
timestamp 1731220342
transform 1 0 3488 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5965_6
timestamp 1731220342
transform 1 0 3672 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5964_6
timestamp 1731220342
transform 1 0 3528 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5963_6
timestamp 1731220342
transform 1 0 3368 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5962_6
timestamp 1731220342
transform 1 0 3200 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5961_6
timestamp 1731220342
transform 1 0 3016 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5960_6
timestamp 1731220342
transform 1 0 3632 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5959_6
timestamp 1731220342
transform 1 0 3432 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5958_6
timestamp 1731220342
transform 1 0 3232 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5957_6
timestamp 1731220342
transform 1 0 3040 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5956_6
timestamp 1731220342
transform 1 0 2848 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5955_6
timestamp 1731220342
transform 1 0 3496 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5954_6
timestamp 1731220342
transform 1 0 3280 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5953_6
timestamp 1731220342
transform 1 0 3072 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5952_6
timestamp 1731220342
transform 1 0 2872 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5951_6
timestamp 1731220342
transform 1 0 3600 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5950_6
timestamp 1731220342
transform 1 0 3384 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5949_6
timestamp 1731220342
transform 1 0 3184 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5948_6
timestamp 1731220342
transform 1 0 3008 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5947_6
timestamp 1731220342
transform 1 0 2856 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5946_6
timestamp 1731220342
transform 1 0 3448 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5945_6
timestamp 1731220342
transform 1 0 3264 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5944_6
timestamp 1731220342
transform 1 0 3096 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5943_6
timestamp 1731220342
transform 1 0 2944 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5942_6
timestamp 1731220342
transform 1 0 3024 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5941_6
timestamp 1731220342
transform 1 0 2816 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5940_6
timestamp 1731220342
transform 1 0 2752 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5939_6
timestamp 1731220342
transform 1 0 2704 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5938_6
timestamp 1731220342
transform 1 0 2640 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5937_6
timestamp 1731220342
transform 1 0 2880 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5936_6
timestamp 1731220342
transform 1 0 2800 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5935_6
timestamp 1731220342
transform 1 0 2936 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5934_6
timestamp 1731220342
transform 1 0 3176 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5933_6
timestamp 1731220342
transform 1 0 3336 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5932_6
timestamp 1731220342
transform 1 0 3440 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5931_6
timestamp 1731220342
transform 1 0 3256 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5930_6
timestamp 1731220342
transform 1 0 3088 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5929_6
timestamp 1731220342
transform 1 0 3064 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5928_6
timestamp 1731220342
transform 1 0 2904 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5927_6
timestamp 1731220342
transform 1 0 3432 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5926_6
timestamp 1731220342
transform 1 0 3240 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5925_6
timestamp 1731220342
transform 1 0 3064 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5924_6
timestamp 1731220342
transform 1 0 2896 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5923_6
timestamp 1731220342
transform 1 0 3240 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5922_6
timestamp 1731220342
transform 1 0 3424 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5921_6
timestamp 1731220342
transform 1 0 3272 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5920_6
timestamp 1731220342
transform 1 0 3104 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5919_6
timestamp 1731220342
transform 1 0 2928 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5918_6
timestamp 1731220342
transform 1 0 3264 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5917_6
timestamp 1731220342
transform 1 0 3432 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5916_6
timestamp 1731220342
transform 1 0 3600 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5915_6
timestamp 1731220342
transform 1 0 3440 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5914_6
timestamp 1731220342
transform 1 0 3616 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5913_6
timestamp 1731220342
transform 1 0 3608 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5912_6
timestamp 1731220342
transform 1 0 3624 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5911_6
timestamp 1731220342
transform 1 0 3632 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5910_6
timestamp 1731220342
transform 1 0 3496 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5909_6
timestamp 1731220342
transform 1 0 3664 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5908_6
timestamp 1731220342
transform 1 0 3640 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5907_6
timestamp 1731220342
transform 1 0 3712 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5906_6
timestamp 1731220342
transform 1 0 3688 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5905_6
timestamp 1731220342
transform 1 0 3696 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5904_6
timestamp 1731220342
transform 1 0 3536 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5903_6
timestamp 1731220342
transform 1 0 3832 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5902_6
timestamp 1731220342
transform 1 0 3832 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5901_6
timestamp 1731220342
transform 1 0 3832 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5900_6
timestamp 1731220342
transform 1 0 3832 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5899_6
timestamp 1731220342
transform 1 0 3816 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5898_6
timestamp 1731220342
transform 1 0 3832 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5897_6
timestamp 1731220342
transform 1 0 3832 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5896_6
timestamp 1731220342
transform 1 0 3832 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5895_6
timestamp 1731220342
transform 1 0 3824 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5894_6
timestamp 1731220342
transform 1 0 3800 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5893_6
timestamp 1731220342
transform 1 0 3776 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5892_6
timestamp 1731220342
transform 1 0 3792 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5891_6
timestamp 1731220342
transform 1 0 3456 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5890_6
timestamp 1731220342
transform 1 0 3560 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5889_6
timestamp 1731220342
transform 1 0 3688 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5888_6
timestamp 1731220342
transform 1 0 3520 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5887_6
timestamp 1731220342
transform 1 0 3352 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5886_6
timestamp 1731220342
transform 1 0 3416 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5885_6
timestamp 1731220342
transform 1 0 3256 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5884_6
timestamp 1731220342
transform 1 0 3120 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5883_6
timestamp 1731220342
transform 1 0 3088 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5882_6
timestamp 1731220342
transform 1 0 2904 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5881_6
timestamp 1731220342
transform 1 0 2784 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5880_6
timestamp 1731220342
transform 1 0 2424 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5879_6
timestamp 1731220342
transform 1 0 2904 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5878_6
timestamp 1731220342
transform 1 0 3088 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5877_6
timestamp 1731220342
transform 1 0 3016 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5876_6
timestamp 1731220342
transform 1 0 3184 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5875_6
timestamp 1731220342
transform 1 0 3120 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5874_6
timestamp 1731220342
transform 1 0 3008 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5873_6
timestamp 1731220342
transform 1 0 2904 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5872_6
timestamp 1731220342
transform 1 0 2800 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5871_6
timestamp 1731220342
transform 1 0 2696 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5870_6
timestamp 1731220342
transform 1 0 2848 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5869_6
timestamp 1731220342
transform 1 0 3064 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5868_6
timestamp 1731220342
transform 1 0 3296 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5867_6
timestamp 1731220342
transform 1 0 3536 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5866_6
timestamp 1731220342
transform 1 0 3664 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5865_6
timestamp 1731220342
transform 1 0 3480 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5864_6
timestamp 1731220342
transform 1 0 3296 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5863_6
timestamp 1731220342
transform 1 0 3120 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5862_6
timestamp 1731220342
transform 1 0 2952 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5861_6
timestamp 1731220342
transform 1 0 3288 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5860_6
timestamp 1731220342
transform 1 0 3408 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5859_6
timestamp 1731220342
transform 1 0 3536 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5858_6
timestamp 1731220342
transform 1 0 3664 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5857_6
timestamp 1731220342
transform 1 0 3720 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5856_6
timestamp 1731220342
transform 1 0 3584 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5855_6
timestamp 1731220342
transform 1 0 3448 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5854_6
timestamp 1731220342
transform 1 0 3304 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5853_6
timestamp 1731220342
transform 1 0 3160 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5852_6
timestamp 1731220342
transform 1 0 3688 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5851_6
timestamp 1731220342
transform 1 0 3520 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5850_6
timestamp 1731220342
transform 1 0 3360 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5849_6
timestamp 1731220342
transform 1 0 3200 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5848_6
timestamp 1731220342
transform 1 0 3040 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5847_6
timestamp 1731220342
transform 1 0 3584 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5846_6
timestamp 1731220342
transform 1 0 3400 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5845_6
timestamp 1731220342
transform 1 0 3216 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5844_6
timestamp 1731220342
transform 1 0 3040 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5843_6
timestamp 1731220342
transform 1 0 2872 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5842_6
timestamp 1731220342
transform 1 0 3608 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5841_6
timestamp 1731220342
transform 1 0 3368 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5840_6
timestamp 1731220342
transform 1 0 3136 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5839_6
timestamp 1731220342
transform 1 0 2928 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5838_6
timestamp 1731220342
transform 1 0 2744 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5837_6
timestamp 1731220342
transform 1 0 3096 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5836_6
timestamp 1731220342
transform 1 0 2928 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5835_6
timestamp 1731220342
transform 1 0 2768 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5834_6
timestamp 1731220342
transform 1 0 2600 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5833_6
timestamp 1731220342
transform 1 0 2424 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5832_6
timestamp 1731220342
transform 1 0 2552 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5831_6
timestamp 1731220342
transform 1 0 2744 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5830_6
timestamp 1731220342
transform 1 0 2944 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5829_6
timestamp 1731220342
transform 1 0 3160 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5828_6
timestamp 1731220342
transform 1 0 3384 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5827_6
timestamp 1731220342
transform 1 0 3496 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5826_6
timestamp 1731220342
transform 1 0 3256 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5825_6
timestamp 1731220342
transform 1 0 3024 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5824_6
timestamp 1731220342
transform 1 0 2816 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5823_6
timestamp 1731220342
transform 1 0 2984 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5822_6
timestamp 1731220342
transform 1 0 3168 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5821_6
timestamp 1731220342
transform 1 0 3160 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5820_6
timestamp 1731220342
transform 1 0 2992 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5819_6
timestamp 1731220342
transform 1 0 3328 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5818_6
timestamp 1731220342
transform 1 0 3240 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5817_6
timestamp 1731220342
transform 1 0 3096 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5816_6
timestamp 1731220342
transform 1 0 3176 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5815_6
timestamp 1731220342
transform 1 0 3304 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5814_6
timestamp 1731220342
transform 1 0 3568 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5813_6
timestamp 1731220342
transform 1 0 3432 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5812_6
timestamp 1731220342
transform 1 0 3384 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5811_6
timestamp 1731220342
transform 1 0 3536 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5810_6
timestamp 1731220342
transform 1 0 3696 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5809_6
timestamp 1731220342
transform 1 0 3680 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5808_6
timestamp 1731220342
transform 1 0 3504 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5807_6
timestamp 1731220342
transform 1 0 3512 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5806_6
timestamp 1731220342
transform 1 0 3344 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5805_6
timestamp 1731220342
transform 1 0 3680 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5804_6
timestamp 1731220342
transform 1 0 3736 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5803_6
timestamp 1731220342
transform 1 0 3616 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5802_6
timestamp 1731220342
transform 1 0 3776 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5801_6
timestamp 1731220342
transform 1 0 3792 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5800_6
timestamp 1731220342
transform 1 0 3784 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5799_6
timestamp 1731220342
transform 1 0 3704 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5798_6
timestamp 1731220342
transform 1 0 3832 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5797_6
timestamp 1731220342
transform 1 0 3832 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5796_6
timestamp 1731220342
transform 1 0 3832 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5795_6
timestamp 1731220342
transform 1 0 3832 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5794_6
timestamp 1731220342
transform 1 0 3832 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5793_6
timestamp 1731220342
transform 1 0 3832 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5792_6
timestamp 1731220342
transform 1 0 3832 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5791_6
timestamp 1731220342
transform 1 0 3832 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5790_6
timestamp 1731220342
transform 1 0 3832 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5789_6
timestamp 1731220342
transform 1 0 3832 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5788_6
timestamp 1731220342
transform 1 0 3832 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5787_6
timestamp 1731220342
transform 1 0 3832 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5786_6
timestamp 1731220342
transform 1 0 3736 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5785_6
timestamp 1731220342
transform 1 0 3632 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5784_6
timestamp 1731220342
transform 1 0 3528 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5783_6
timestamp 1731220342
transform 1 0 3616 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5782_6
timestamp 1731220342
transform 1 0 3392 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5781_6
timestamp 1731220342
transform 1 0 3424 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5780_6
timestamp 1731220342
transform 1 0 3320 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5779_6
timestamp 1731220342
transform 1 0 3208 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5778_6
timestamp 1731220342
transform 1 0 3096 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5777_6
timestamp 1731220342
transform 1 0 2976 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5776_6
timestamp 1731220342
transform 1 0 2896 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5775_6
timestamp 1731220342
transform 1 0 3168 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5774_6
timestamp 1731220342
transform 1 0 3440 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5773_6
timestamp 1731220342
transform 1 0 3320 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5772_6
timestamp 1731220342
transform 1 0 3160 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5771_6
timestamp 1731220342
transform 1 0 3008 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5770_6
timestamp 1731220342
transform 1 0 2928 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5769_6
timestamp 1731220342
transform 1 0 3088 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5768_6
timestamp 1731220342
transform 1 0 3256 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5767_6
timestamp 1731220342
transform 1 0 3152 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5766_6
timestamp 1731220342
transform 1 0 3296 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5765_6
timestamp 1731220342
transform 1 0 3264 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5764_6
timestamp 1731220342
transform 1 0 3400 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5763_6
timestamp 1731220342
transform 1 0 3480 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5762_6
timestamp 1731220342
transform 1 0 3344 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5761_6
timestamp 1731220342
transform 1 0 3320 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5760_6
timestamp 1731220342
transform 1 0 3560 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5759_6
timestamp 1731220342
transform 1 0 3512 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5758_6
timestamp 1731220342
transform 1 0 3312 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5757_6
timestamp 1731220342
transform 1 0 3720 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5756_6
timestamp 1731220342
transform 1 0 3728 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5755_6
timestamp 1731220342
transform 1 0 3528 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5754_6
timestamp 1731220342
transform 1 0 3328 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5753_6
timestamp 1731220342
transform 1 0 3320 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5752_6
timestamp 1731220342
transform 1 0 3488 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5751_6
timestamp 1731220342
transform 1 0 3656 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5750_6
timestamp 1731220342
transform 1 0 3528 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5749_6
timestamp 1731220342
transform 1 0 3408 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5748_6
timestamp 1731220342
transform 1 0 3288 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5747_6
timestamp 1731220342
transform 1 0 3168 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5746_6
timestamp 1731220342
transform 1 0 3048 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5745_6
timestamp 1731220342
transform 1 0 2920 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5744_6
timestamp 1731220342
transform 1 0 2784 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5743_6
timestamp 1731220342
transform 1 0 3152 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5742_6
timestamp 1731220342
transform 1 0 2984 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5741_6
timestamp 1731220342
transform 1 0 2944 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5740_6
timestamp 1731220342
transform 1 0 3136 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5739_6
timestamp 1731220342
transform 1 0 3112 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5738_6
timestamp 1731220342
transform 1 0 2904 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5737_6
timestamp 1731220342
transform 1 0 3088 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5736_6
timestamp 1731220342
transform 1 0 3216 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5735_6
timestamp 1731220342
transform 1 0 3136 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5734_6
timestamp 1731220342
transform 1 0 3016 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5733_6
timestamp 1731220342
transform 1 0 2880 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5732_6
timestamp 1731220342
transform 1 0 2768 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5731_6
timestamp 1731220342
transform 1 0 2856 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5730_6
timestamp 1731220342
transform 1 0 2696 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5729_6
timestamp 1731220342
transform 1 0 2624 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5728_6
timestamp 1731220342
transform 1 0 2336 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5727_6
timestamp 1731220342
transform 1 0 2856 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5726_6
timestamp 1731220342
transform 1 0 2736 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5725_6
timestamp 1731220342
transform 1 0 2608 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5724_6
timestamp 1731220342
transform 1 0 2480 0 1 2988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5723_6
timestamp 1731220342
transform 1 0 2400 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5722_6
timestamp 1731220342
transform 1 0 2568 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5721_6
timestamp 1731220342
transform 1 0 2760 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5720_6
timestamp 1731220342
transform 1 0 2960 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5719_6
timestamp 1731220342
transform 1 0 3176 0 -1 2984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5718_6
timestamp 1731220342
transform 1 0 3048 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5717_6
timestamp 1731220342
transform 1 0 2920 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5716_6
timestamp 1731220342
transform 1 0 2792 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5715_6
timestamp 1731220342
transform 1 0 2664 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5714_6
timestamp 1731220342
transform 1 0 2544 0 1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5713_6
timestamp 1731220342
transform 1 0 2960 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5712_6
timestamp 1731220342
transform 1 0 2824 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5711_6
timestamp 1731220342
transform 1 0 2688 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5710_6
timestamp 1731220342
transform 1 0 2560 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5709_6
timestamp 1731220342
transform 1 0 2432 0 -1 2816
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5708_6
timestamp 1731220342
transform 1 0 2824 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5707_6
timestamp 1731220342
transform 1 0 2656 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5706_6
timestamp 1731220342
transform 1 0 2488 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5705_6
timestamp 1731220342
transform 1 0 2328 0 1 2656
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5704_6
timestamp 1731220342
transform 1 0 2800 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5703_6
timestamp 1731220342
transform 1 0 2616 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5702_6
timestamp 1731220342
transform 1 0 2440 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5701_6
timestamp 1731220342
transform 1 0 2272 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5700_6
timestamp 1731220342
transform 1 0 2120 0 -1 2652
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5699_6
timestamp 1731220342
transform 1 0 2632 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5698_6
timestamp 1731220342
transform 1 0 2464 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5697_6
timestamp 1731220342
transform 1 0 2312 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5696_6
timestamp 1731220342
transform 1 0 2176 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5695_6
timestamp 1731220342
transform 1 0 2064 0 1 2492
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5694_6
timestamp 1731220342
transform 1 0 2376 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5693_6
timestamp 1731220342
transform 1 0 2208 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5692_6
timestamp 1731220342
transform 1 0 2064 0 -1 2488
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5691_6
timestamp 1731220342
transform 1 0 1896 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5690_6
timestamp 1731220342
transform 1 0 1784 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5689_6
timestamp 1731220342
transform 1 0 1656 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5688_6
timestamp 1731220342
transform 1 0 1896 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5687_6
timestamp 1731220342
transform 1 0 2064 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5686_6
timestamp 1731220342
transform 1 0 2240 0 1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5685_6
timestamp 1731220342
transform 1 0 2168 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5684_6
timestamp 1731220342
transform 1 0 2064 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5683_6
timestamp 1731220342
transform 1 0 2304 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5682_6
timestamp 1731220342
transform 1 0 2584 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5681_6
timestamp 1731220342
transform 1 0 2440 0 -1 2320
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5680_6
timestamp 1731220342
transform 1 0 2400 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5679_6
timestamp 1731220342
transform 1 0 2248 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5678_6
timestamp 1731220342
transform 1 0 2104 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5677_6
timestamp 1731220342
transform 1 0 2552 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5676_6
timestamp 1731220342
transform 1 0 2712 0 1 2160
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5675_6
timestamp 1731220342
transform 1 0 2576 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5674_6
timestamp 1731220342
transform 1 0 2424 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5673_6
timestamp 1731220342
transform 1 0 2280 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5672_6
timestamp 1731220342
transform 1 0 2728 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5671_6
timestamp 1731220342
transform 1 0 2880 0 -1 2148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5670_6
timestamp 1731220342
transform 1 0 3000 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5669_6
timestamp 1731220342
transform 1 0 2832 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5668_6
timestamp 1731220342
transform 1 0 2664 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5667_6
timestamp 1731220342
transform 1 0 2496 0 1 1988
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5666_6
timestamp 1731220342
transform 1 0 2488 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5665_6
timestamp 1731220342
transform 1 0 2584 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5664_6
timestamp 1731220342
transform 1 0 2688 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5663_6
timestamp 1731220342
transform 1 0 2800 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5662_6
timestamp 1731220342
transform 1 0 3168 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5661_6
timestamp 1731220342
transform 1 0 3040 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5660_6
timestamp 1731220342
transform 1 0 2920 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5659_6
timestamp 1731220342
transform 1 0 2784 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5658_6
timestamp 1731220342
transform 1 0 2616 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5657_6
timestamp 1731220342
transform 1 0 2432 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5656_6
timestamp 1731220342
transform 1 0 2240 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5655_6
timestamp 1731220342
transform 1 0 2504 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5654_6
timestamp 1731220342
transform 1 0 2664 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5653_6
timestamp 1731220342
transform 1 0 2592 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5652_6
timestamp 1731220342
transform 1 0 2488 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5651_6
timestamp 1731220342
transform 1 0 2672 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5650_6
timestamp 1731220342
transform 1 0 2840 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5649_6
timestamp 1731220342
transform 1 0 2704 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5648_6
timestamp 1731220342
transform 1 0 2512 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5647_6
timestamp 1731220342
transform 1 0 2360 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5646_6
timestamp 1731220342
transform 1 0 2224 0 -1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5645_6
timestamp 1731220342
transform 1 0 2176 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5644_6
timestamp 1731220342
transform 1 0 2280 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5643_6
timestamp 1731220342
transform 1 0 2384 0 1 1676
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5642_6
timestamp 1731220342
transform 1 0 2360 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5641_6
timestamp 1731220342
transform 1 0 2224 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5640_6
timestamp 1731220342
transform 1 0 2088 0 -1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5639_6
timestamp 1731220342
transform 1 0 2064 0 1 1828
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5638_6
timestamp 1731220342
transform 1 0 1840 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5637_6
timestamp 1731220342
transform 1 0 1576 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5636_6
timestamp 1731220342
transform 1 0 1440 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5635_6
timestamp 1731220342
transform 1 0 1304 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5634_6
timestamp 1731220342
transform 1 0 1272 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5633_6
timestamp 1731220342
transform 1 0 1552 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5632_6
timestamp 1731220342
transform 1 0 1408 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5631_6
timestamp 1731220342
transform 1 0 1392 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5630_6
timestamp 1731220342
transform 1 0 1576 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5629_6
timestamp 1731220342
transform 1 0 1624 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5628_6
timestamp 1731220342
transform 1 0 1440 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5627_6
timestamp 1731220342
transform 1 0 1256 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5626_6
timestamp 1731220342
transform 1 0 1320 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5625_6
timestamp 1731220342
transform 1 0 1560 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5624_6
timestamp 1731220342
transform 1 0 1440 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5623_6
timestamp 1731220342
transform 1 0 1256 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5622_6
timestamp 1731220342
transform 1 0 1080 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5621_6
timestamp 1731220342
transform 1 0 912 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5620_6
timestamp 1731220342
transform 1 0 1088 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5619_6
timestamp 1731220342
transform 1 0 1088 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5618_6
timestamp 1731220342
transform 1 0 928 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5617_6
timestamp 1731220342
transform 1 0 1040 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5616_6
timestamp 1731220342
transform 1 0 1208 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5615_6
timestamp 1731220342
transform 1 0 1136 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5614_6
timestamp 1731220342
transform 1 0 1168 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5613_6
timestamp 1731220342
transform 1 0 1144 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5612_6
timestamp 1731220342
transform 1 0 1312 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5611_6
timestamp 1731220342
transform 1 0 1432 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5610_6
timestamp 1731220342
transform 1 0 1272 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5609_6
timestamp 1731220342
transform 1 0 1120 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5608_6
timestamp 1731220342
transform 1 0 1160 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5607_6
timestamp 1731220342
transform 1 0 1344 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5606_6
timestamp 1731220342
transform 1 0 1360 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5605_6
timestamp 1731220342
transform 1 0 1176 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5604_6
timestamp 1731220342
transform 1 0 1176 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5603_6
timestamp 1731220342
transform 1 0 1344 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5602_6
timestamp 1731220342
transform 1 0 1536 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5601_6
timestamp 1731220342
transform 1 0 1728 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5600_6
timestamp 1731220342
transform 1 0 1648 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5599_6
timestamp 1731220342
transform 1 0 1856 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5598_6
timestamp 1731220342
transform 1 0 1888 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5597_6
timestamp 1731220342
transform 1 0 1712 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5596_6
timestamp 1731220342
transform 1 0 1832 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5595_6
timestamp 1731220342
transform 1 0 1680 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5594_6
timestamp 1731220342
transform 1 0 1536 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5593_6
timestamp 1731220342
transform 1 0 1616 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5592_6
timestamp 1731220342
transform 1 0 1392 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5591_6
timestamp 1731220342
transform 1 0 1240 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5590_6
timestamp 1731220342
transform 1 0 1184 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5589_6
timestamp 1731220342
transform 1 0 1360 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5588_6
timestamp 1731220342
transform 1 0 1536 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5587_6
timestamp 1731220342
transform 1 0 1440 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5586_6
timestamp 1731220342
transform 1 0 1240 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5585_6
timestamp 1731220342
transform 1 0 1040 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5584_6
timestamp 1731220342
transform 1 0 1152 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5583_6
timestamp 1731220342
transform 1 0 968 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5582_6
timestamp 1731220342
transform 1 0 872 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5581_6
timestamp 1731220342
transform 1 0 1032 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5580_6
timestamp 1731220342
transform 1 0 984 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5579_6
timestamp 1731220342
transform 1 0 976 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5578_6
timestamp 1731220342
transform 1 0 976 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5577_6
timestamp 1731220342
transform 1 0 840 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5576_6
timestamp 1731220342
transform 1 0 856 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5575_6
timestamp 1731220342
transform 1 0 992 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5574_6
timestamp 1731220342
transform 1 0 1040 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5573_6
timestamp 1731220342
transform 1 0 1000 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5572_6
timestamp 1731220342
transform 1 0 864 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5571_6
timestamp 1731220342
transform 1 0 888 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5570_6
timestamp 1731220342
transform 1 0 744 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5569_6
timestamp 1731220342
transform 1 0 776 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5568_6
timestamp 1731220342
transform 1 0 872 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5567_6
timestamp 1731220342
transform 1 0 672 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5566_6
timestamp 1731220342
transform 1 0 584 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5565_6
timestamp 1731220342
transform 1 0 744 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5564_6
timestamp 1731220342
transform 1 0 968 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5563_6
timestamp 1731220342
transform 1 0 760 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5562_6
timestamp 1731220342
transform 1 0 544 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5561_6
timestamp 1731220342
transform 1 0 704 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5560_6
timestamp 1731220342
transform 1 0 896 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5559_6
timestamp 1731220342
transform 1 0 920 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5558_6
timestamp 1731220342
transform 1 0 768 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5557_6
timestamp 1731220342
transform 1 0 600 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5556_6
timestamp 1731220342
transform 1 0 536 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5555_6
timestamp 1731220342
transform 1 0 704 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5554_6
timestamp 1731220342
transform 1 0 760 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5553_6
timestamp 1731220342
transform 1 0 632 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5552_6
timestamp 1731220342
transform 1 0 496 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5551_6
timestamp 1731220342
transform 1 0 600 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5550_6
timestamp 1731220342
transform 1 0 736 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5549_6
timestamp 1731220342
transform 1 0 872 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5548_6
timestamp 1731220342
transform 1 0 992 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5547_6
timestamp 1731220342
transform 1 0 808 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5546_6
timestamp 1731220342
transform 1 0 624 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5545_6
timestamp 1731220342
transform 1 0 440 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5544_6
timestamp 1731220342
transform 1 0 272 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5543_6
timestamp 1731220342
transform 1 0 464 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5542_6
timestamp 1731220342
transform 1 0 344 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5541_6
timestamp 1731220342
transform 1 0 232 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5540_6
timestamp 1731220342
transform 1 0 216 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5539_6
timestamp 1731220342
transform 1 0 360 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5538_6
timestamp 1731220342
transform 1 0 360 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5537_6
timestamp 1731220342
transform 1 0 168 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5536_6
timestamp 1731220342
transform 1 0 128 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5535_6
timestamp 1731220342
transform 1 0 264 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5534_6
timestamp 1731220342
transform 1 0 432 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5533_6
timestamp 1731220342
transform 1 0 504 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5532_6
timestamp 1731220342
transform 1 0 304 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5531_6
timestamp 1731220342
transform 1 0 128 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5530_6
timestamp 1731220342
transform 1 0 128 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5529_6
timestamp 1731220342
transform 1 0 320 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5528_6
timestamp 1731220342
transform 1 0 264 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5527_6
timestamp 1731220342
transform 1 0 128 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5526_6
timestamp 1731220342
transform 1 0 424 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5525_6
timestamp 1731220342
transform 1 0 320 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5524_6
timestamp 1731220342
transform 1 0 152 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5523_6
timestamp 1731220342
transform 1 0 488 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5522_6
timestamp 1731220342
transform 1 0 488 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5521_6
timestamp 1731220342
transform 1 0 352 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5520_6
timestamp 1731220342
transform 1 0 216 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5519_6
timestamp 1731220342
transform 1 0 632 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5518_6
timestamp 1731220342
transform 1 0 608 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5517_6
timestamp 1731220342
transform 1 0 488 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5516_6
timestamp 1731220342
transform 1 0 368 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5515_6
timestamp 1731220342
transform 1 0 504 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5514_6
timestamp 1731220342
transform 1 0 616 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5513_6
timestamp 1731220342
transform 1 0 736 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5512_6
timestamp 1731220342
transform 1 0 904 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5511_6
timestamp 1731220342
transform 1 0 776 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5510_6
timestamp 1731220342
transform 1 0 656 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5509_6
timestamp 1731220342
transform 1 0 544 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5508_6
timestamp 1731220342
transform 1 0 496 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5507_6
timestamp 1731220342
transform 1 0 608 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5506_6
timestamp 1731220342
transform 1 0 728 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5505_6
timestamp 1731220342
transform 1 0 712 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5504_6
timestamp 1731220342
transform 1 0 584 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5503_6
timestamp 1731220342
transform 1 0 456 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5502_6
timestamp 1731220342
transform 1 0 336 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5501_6
timestamp 1731220342
transform 1 0 792 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5500_6
timestamp 1731220342
transform 1 0 616 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5499_6
timestamp 1731220342
transform 1 0 448 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5498_6
timestamp 1731220342
transform 1 0 288 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5497_6
timestamp 1731220342
transform 1 0 152 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5496_6
timestamp 1731220342
transform 1 0 792 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5495_6
timestamp 1731220342
transform 1 0 600 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5494_6
timestamp 1731220342
transform 1 0 416 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5493_6
timestamp 1731220342
transform 1 0 248 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5492_6
timestamp 1731220342
transform 1 0 128 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5491_6
timestamp 1731220342
transform 1 0 712 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5490_6
timestamp 1731220342
transform 1 0 552 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5489_6
timestamp 1731220342
transform 1 0 392 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5488_6
timestamp 1731220342
transform 1 0 240 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5487_6
timestamp 1731220342
transform 1 0 128 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5486_6
timestamp 1731220342
transform 1 0 128 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5485_6
timestamp 1731220342
transform 1 0 256 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5484_6
timestamp 1731220342
transform 1 0 424 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5483_6
timestamp 1731220342
transform 1 0 784 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5482_6
timestamp 1731220342
transform 1 0 600 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5481_6
timestamp 1731220342
transform 1 0 472 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5480_6
timestamp 1731220342
transform 1 0 304 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5479_6
timestamp 1731220342
transform 1 0 152 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5478_6
timestamp 1731220342
transform 1 0 848 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5477_6
timestamp 1731220342
transform 1 0 656 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5476_6
timestamp 1731220342
transform 1 0 536 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5475_6
timestamp 1731220342
transform 1 0 400 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5474_6
timestamp 1731220342
transform 1 0 1016 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5473_6
timestamp 1731220342
transform 1 0 848 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5472_6
timestamp 1731220342
transform 1 0 688 0 1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5471_6
timestamp 1731220342
transform 1 0 584 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5470_6
timestamp 1731220342
transform 1 0 416 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5469_6
timestamp 1731220342
transform 1 0 368 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5468_6
timestamp 1731220342
transform 1 0 296 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5467_6
timestamp 1731220342
transform 1 0 440 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5466_6
timestamp 1731220342
transform 1 0 440 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5465_6
timestamp 1731220342
transform 1 0 248 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5464_6
timestamp 1731220342
transform 1 0 248 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5463_6
timestamp 1731220342
transform 1 0 152 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5462_6
timestamp 1731220342
transform 1 0 304 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5461_6
timestamp 1731220342
transform 1 0 256 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5460_6
timestamp 1731220342
transform 1 0 128 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5459_6
timestamp 1731220342
transform 1 0 128 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5458_6
timestamp 1731220342
transform 1 0 240 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5457_6
timestamp 1731220342
transform 1 0 288 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5456_6
timestamp 1731220342
transform 1 0 128 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5455_6
timestamp 1731220342
transform 1 0 128 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5454_6
timestamp 1731220342
transform 1 0 280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5453_6
timestamp 1731220342
transform 1 0 280 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5452_6
timestamp 1731220342
transform 1 0 128 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5451_6
timestamp 1731220342
transform 1 0 152 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5450_6
timestamp 1731220342
transform 1 0 344 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5449_6
timestamp 1731220342
transform 1 0 376 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5448_6
timestamp 1731220342
transform 1 0 216 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5447_6
timestamp 1731220342
transform 1 0 224 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5446_6
timestamp 1731220342
transform 1 0 128 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5445_6
timestamp 1731220342
transform 1 0 320 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5444_6
timestamp 1731220342
transform 1 0 416 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5443_6
timestamp 1731220342
transform 1 0 520 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5442_6
timestamp 1731220342
transform 1 0 896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5441_6
timestamp 1731220342
transform 1 0 768 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5440_6
timestamp 1731220342
transform 1 0 640 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5439_6
timestamp 1731220342
transform 1 0 536 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5438_6
timestamp 1731220342
transform 1 0 696 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5437_6
timestamp 1731220342
transform 1 0 856 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5436_6
timestamp 1731220342
transform 1 0 952 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5435_6
timestamp 1731220342
transform 1 0 752 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5434_6
timestamp 1731220342
transform 1 0 544 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5433_6
timestamp 1731220342
transform 1 0 440 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5432_6
timestamp 1731220342
transform 1 0 592 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5431_6
timestamp 1731220342
transform 1 0 744 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5430_6
timestamp 1731220342
transform 1 0 760 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5429_6
timestamp 1731220342
transform 1 0 608 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5428_6
timestamp 1731220342
transform 1 0 448 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5427_6
timestamp 1731220342
transform 1 0 472 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5426_6
timestamp 1731220342
transform 1 0 656 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5425_6
timestamp 1731220342
transform 1 0 680 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5424_6
timestamp 1731220342
transform 1 0 520 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5423_6
timestamp 1731220342
transform 1 0 376 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5422_6
timestamp 1731220342
transform 1 0 424 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5421_6
timestamp 1731220342
transform 1 0 616 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5420_6
timestamp 1731220342
transform 1 0 816 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5419_6
timestamp 1731220342
transform 1 0 768 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5418_6
timestamp 1731220342
transform 1 0 616 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5417_6
timestamp 1731220342
transform 1 0 464 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5416_6
timestamp 1731220342
transform 1 0 440 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5415_6
timestamp 1731220342
transform 1 0 632 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5414_6
timestamp 1731220342
transform 1 0 816 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5413_6
timestamp 1731220342
transform 1 0 992 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5412_6
timestamp 1731220342
transform 1 0 968 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5411_6
timestamp 1731220342
transform 1 0 800 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5410_6
timestamp 1731220342
transform 1 0 624 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5409_6
timestamp 1731220342
transform 1 0 584 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5408_6
timestamp 1731220342
transform 1 0 848 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5407_6
timestamp 1731220342
transform 1 0 720 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5406_6
timestamp 1731220342
transform 1 0 704 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5405_6
timestamp 1731220342
transform 1 0 592 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5404_6
timestamp 1731220342
transform 1 0 480 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5403_6
timestamp 1731220342
transform 1 0 752 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5402_6
timestamp 1731220342
transform 1 0 920 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5401_6
timestamp 1731220342
transform 1 0 1088 0 -1 1200
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5400_6
timestamp 1731220342
transform 1 0 1112 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5399_6
timestamp 1731220342
transform 1 0 960 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5398_6
timestamp 1731220342
transform 1 0 824 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5397_6
timestamp 1731220342
transform 1 0 1272 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5396_6
timestamp 1731220342
transform 1 0 1440 0 1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5395_6
timestamp 1731220342
transform 1 0 1424 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5394_6
timestamp 1731220342
transform 1 0 1304 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5393_6
timestamp 1731220342
transform 1 0 1192 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5392_6
timestamp 1731220342
transform 1 0 1080 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5391_6
timestamp 1731220342
transform 1 0 968 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5390_6
timestamp 1731220342
transform 1 0 1120 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5389_6
timestamp 1731220342
transform 1 0 1264 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5388_6
timestamp 1731220342
transform 1 0 1408 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5387_6
timestamp 1731220342
transform 1 0 1544 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5386_6
timestamp 1731220342
transform 1 0 1688 0 1 892
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5385_6
timestamp 1731220342
transform 1 0 1776 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5384_6
timestamp 1731220342
transform 1 0 1624 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5383_6
timestamp 1731220342
transform 1 0 1472 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5382_6
timestamp 1731220342
transform 1 0 1320 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5381_6
timestamp 1731220342
transform 1 0 1160 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5380_6
timestamp 1731220342
transform 1 0 1576 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5379_6
timestamp 1731220342
transform 1 0 1408 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5378_6
timestamp 1731220342
transform 1 0 1248 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5377_6
timestamp 1731220342
transform 1 0 1088 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5376_6
timestamp 1731220342
transform 1 0 928 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5375_6
timestamp 1731220342
transform 1 0 1008 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5374_6
timestamp 1731220342
transform 1 0 1200 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5373_6
timestamp 1731220342
transform 1 0 1536 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5372_6
timestamp 1731220342
transform 1 0 1296 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5371_6
timestamp 1731220342
transform 1 0 1072 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5370_6
timestamp 1731220342
transform 1 0 864 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5369_6
timestamp 1731220342
transform 1 0 840 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5368_6
timestamp 1731220342
transform 1 0 1208 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5367_6
timestamp 1731220342
transform 1 0 1024 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5366_6
timestamp 1731220342
transform 1 0 896 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5365_6
timestamp 1731220342
transform 1 0 896 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5364_6
timestamp 1731220342
transform 1 0 1072 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5363_6
timestamp 1731220342
transform 1 0 1264 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5362_6
timestamp 1731220342
transform 1 0 1152 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5361_6
timestamp 1731220342
transform 1 0 1696 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5360_6
timestamp 1731220342
transform 1 0 1472 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5359_6
timestamp 1731220342
transform 1 0 1280 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5358_6
timestamp 1731220342
transform 1 0 1152 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5357_6
timestamp 1731220342
transform 1 0 1024 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5356_6
timestamp 1731220342
transform 1 0 1408 0 1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5355_6
timestamp 1731220342
transform 1 0 1392 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5354_6
timestamp 1731220342
transform 1 0 1584 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5353_6
timestamp 1731220342
transform 1 0 1776 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5352_6
timestamp 1731220342
transform 1 0 1776 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5351_6
timestamp 1731220342
transform 1 0 1560 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5350_6
timestamp 1731220342
transform 1 0 1384 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5349_6
timestamp 1731220342
transform 1 0 1736 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5348_6
timestamp 1731220342
transform 1 0 1896 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5347_6
timestamp 1731220342
transform 1 0 1744 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5346_6
timestamp 1731220342
transform 1 0 1896 0 1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5345_6
timestamp 1731220342
transform 1 0 2064 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5344_6
timestamp 1731220342
transform 1 0 2248 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5343_6
timestamp 1731220342
transform 1 0 2448 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5342_6
timestamp 1731220342
transform 1 0 2424 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5341_6
timestamp 1731220342
transform 1 0 2224 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5340_6
timestamp 1731220342
transform 1 0 2064 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5339_6
timestamp 1731220342
transform 1 0 2392 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5338_6
timestamp 1731220342
transform 1 0 2576 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5337_6
timestamp 1731220342
transform 1 0 2768 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5336_6
timestamp 1731220342
transform 1 0 2720 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5335_6
timestamp 1731220342
transform 1 0 2552 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5334_6
timestamp 1731220342
transform 1 0 2384 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5333_6
timestamp 1731220342
transform 1 0 2216 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5332_6
timestamp 1731220342
transform 1 0 2456 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5331_6
timestamp 1731220342
transform 1 0 2552 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5330_6
timestamp 1731220342
transform 1 0 2648 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5329_6
timestamp 1731220342
transform 1 0 2744 0 -1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5328_6
timestamp 1731220342
transform 1 0 2904 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5327_6
timestamp 1731220342
transform 1 0 2752 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5326_6
timestamp 1731220342
transform 1 0 2616 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5325_6
timestamp 1731220342
transform 1 0 2496 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5324_6
timestamp 1731220342
transform 1 0 2392 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5323_6
timestamp 1731220342
transform 1 0 2680 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5322_6
timestamp 1731220342
transform 1 0 2512 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5321_6
timestamp 1731220342
transform 1 0 2344 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5320_6
timestamp 1731220342
transform 1 0 2184 0 -1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5319_6
timestamp 1731220342
transform 1 0 2736 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5318_6
timestamp 1731220342
transform 1 0 2608 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5317_6
timestamp 1731220342
transform 1 0 2480 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5316_6
timestamp 1731220342
transform 1 0 2360 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5315_6
timestamp 1731220342
transform 1 0 2256 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5314_6
timestamp 1731220342
transform 1 0 2160 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5313_6
timestamp 1731220342
transform 1 0 2064 0 1 84
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5312_6
timestamp 1731220342
transform 1 0 1896 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5311_6
timestamp 1731220342
transform 1 0 1896 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5310_6
timestamp 1731220342
transform 1 0 1800 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5309_6
timestamp 1731220342
transform 1 0 1696 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5308_6
timestamp 1731220342
transform 1 0 1584 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5307_6
timestamp 1731220342
transform 1 0 1480 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5306_6
timestamp 1731220342
transform 1 0 1376 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5305_6
timestamp 1731220342
transform 1 0 1264 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5304_6
timestamp 1731220342
transform 1 0 1144 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5303_6
timestamp 1731220342
transform 1 0 1024 0 1 88
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5302_6
timestamp 1731220342
transform 1 0 1024 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5301_6
timestamp 1731220342
transform 1 0 1192 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5300_6
timestamp 1731220342
transform 1 0 1360 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5299_6
timestamp 1731220342
transform 1 0 1536 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5298_6
timestamp 1731220342
transform 1 0 1720 0 -1 260
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5297_6
timestamp 1731220342
transform 1 0 1704 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5296_6
timestamp 1731220342
transform 1 0 1520 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5295_6
timestamp 1731220342
transform 1 0 1336 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5294_6
timestamp 1731220342
transform 1 0 1888 0 1 268
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5293_6
timestamp 1731220342
transform 1 0 1896 0 -1 424
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5292_6
timestamp 1731220342
transform 1 0 2064 0 1 420
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5291_6
timestamp 1731220342
transform 1 0 2064 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5290_6
timestamp 1731220342
transform 1 0 2208 0 -1 576
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5289_6
timestamp 1731220342
transform 1 0 2624 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5288_6
timestamp 1731220342
transform 1 0 2824 0 1 580
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5287_6
timestamp 1731220342
transform 1 0 2648 0 -1 732
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5286_6
timestamp 1731220342
transform 1 0 2680 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5285_6
timestamp 1731220342
transform 1 0 2488 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5284_6
timestamp 1731220342
transform 1 0 2304 0 1 736
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5283_6
timestamp 1731220342
transform 1 0 2336 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5282_6
timestamp 1731220342
transform 1 0 2432 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5281_6
timestamp 1731220342
transform 1 0 2528 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5280_6
timestamp 1731220342
transform 1 0 2728 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5279_6
timestamp 1731220342
transform 1 0 2624 0 -1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5278_6
timestamp 1731220342
transform 1 0 2608 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5277_6
timestamp 1731220342
transform 1 0 2512 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5276_6
timestamp 1731220342
transform 1 0 2416 0 1 888
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5275_6
timestamp 1731220342
transform 1 0 2448 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5274_6
timestamp 1731220342
transform 1 0 2544 0 -1 1044
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5273_6
timestamp 1731220342
transform 1 0 2688 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5272_6
timestamp 1731220342
transform 1 0 2592 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5271_6
timestamp 1731220342
transform 1 0 2496 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5270_6
timestamp 1731220342
transform 1 0 2400 0 1 1048
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5269_6
timestamp 1731220342
transform 1 0 2760 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5268_6
timestamp 1731220342
transform 1 0 2632 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5267_6
timestamp 1731220342
transform 1 0 2520 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5266_6
timestamp 1731220342
transform 1 0 2408 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5265_6
timestamp 1731220342
transform 1 0 2304 0 -1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5264_6
timestamp 1731220342
transform 1 0 2736 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5263_6
timestamp 1731220342
transform 1 0 2576 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5262_6
timestamp 1731220342
transform 1 0 2424 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5261_6
timestamp 1731220342
transform 1 0 2280 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5260_6
timestamp 1731220342
transform 1 0 2144 0 1 1204
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5259_6
timestamp 1731220342
transform 1 0 2744 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5258_6
timestamp 1731220342
transform 1 0 2560 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5257_6
timestamp 1731220342
transform 1 0 2376 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5256_6
timestamp 1731220342
transform 1 0 2200 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5255_6
timestamp 1731220342
transform 1 0 2064 0 -1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5254_6
timestamp 1731220342
transform 1 0 2704 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5253_6
timestamp 1731220342
transform 1 0 2488 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5252_6
timestamp 1731220342
transform 1 0 2264 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5251_6
timestamp 1731220342
transform 1 0 2064 0 1 1356
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5250_6
timestamp 1731220342
transform 1 0 1896 0 1 1360
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5249_6
timestamp 1731220342
transform 1 0 1800 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5248_6
timestamp 1731220342
transform 1 0 1896 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5247_6
timestamp 1731220342
transform 1 0 2064 0 -1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5246_6
timestamp 1731220342
transform 1 0 2488 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5245_6
timestamp 1731220342
transform 1 0 2264 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5244_6
timestamp 1731220342
transform 1 0 2064 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5243_6
timestamp 1731220342
transform 1 0 1896 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5242_6
timestamp 1731220342
transform 1 0 1680 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5241_6
timestamp 1731220342
transform 1 0 1560 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5240_6
timestamp 1731220342
transform 1 0 1440 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5239_6
timestamp 1731220342
transform 1 0 1312 0 -1 1512
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5238_6
timestamp 1731220342
transform 1 0 1544 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5237_6
timestamp 1731220342
transform 1 0 1728 0 1 1516
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5236_6
timestamp 1731220342
transform 1 0 1728 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5235_6
timestamp 1731220342
transform 1 0 1536 0 -1 1668
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5234_6
timestamp 1731220342
transform 1 0 1592 0 1 1672
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5233_6
timestamp 1731220342
transform 1 0 1480 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5232_6
timestamp 1731220342
transform 1 0 1656 0 -1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5231_6
timestamp 1731220342
transform 1 0 1712 0 1 1824
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5230_6
timestamp 1731220342
transform 1 0 1696 0 -1 1984
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5229_6
timestamp 1731220342
transform 1 0 1768 0 1 1992
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5228_6
timestamp 1731220342
transform 1 0 1816 0 -1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5227_6
timestamp 1731220342
transform 1 0 1808 0 1 2152
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5226_6
timestamp 1731220342
transform 1 0 1808 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5225_6
timestamp 1731220342
transform 1 0 1624 0 -1 2304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5224_6
timestamp 1731220342
transform 1 0 1728 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5223_6
timestamp 1731220342
transform 1 0 1544 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5222_6
timestamp 1731220342
transform 1 0 1360 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5221_6
timestamp 1731220342
transform 1 0 1168 0 1 2312
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5220_6
timestamp 1731220342
transform 1 0 1520 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5219_6
timestamp 1731220342
transform 1 0 1384 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5218_6
timestamp 1731220342
transform 1 0 1232 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5217_6
timestamp 1731220342
transform 1 0 1072 0 -1 2464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5216_6
timestamp 1731220342
transform 1 0 1632 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5215_6
timestamp 1731220342
transform 1 0 1488 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5214_6
timestamp 1731220342
transform 1 0 1352 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5213_6
timestamp 1731220342
transform 1 0 1216 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5212_6
timestamp 1731220342
transform 1 0 1072 0 1 2468
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5211_6
timestamp 1731220342
transform 1 0 1416 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5210_6
timestamp 1731220342
transform 1 0 1272 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5209_6
timestamp 1731220342
transform 1 0 1136 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5208_6
timestamp 1731220342
transform 1 0 1000 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5207_6
timestamp 1731220342
transform 1 0 856 0 -1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5206_6
timestamp 1731220342
transform 1 0 880 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5205_6
timestamp 1731220342
transform 1 0 992 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5204_6
timestamp 1731220342
transform 1 0 1104 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5203_6
timestamp 1731220342
transform 1 0 1344 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5202_6
timestamp 1731220342
transform 1 0 1224 0 1 2624
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5201_6
timestamp 1731220342
transform 1 0 1144 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5200_6
timestamp 1731220342
transform 1 0 1008 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5199_6
timestamp 1731220342
transform 1 0 1280 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5198_6
timestamp 1731220342
transform 1 0 1560 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5197_6
timestamp 1731220342
transform 1 0 1416 0 -1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5196_6
timestamp 1731220342
transform 1 0 1352 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5195_6
timestamp 1731220342
transform 1 0 1176 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5194_6
timestamp 1731220342
transform 1 0 1520 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5193_6
timestamp 1731220342
transform 1 0 1688 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5192_6
timestamp 1731220342
transform 1 0 1856 0 1 2776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5191_6
timestamp 1731220342
transform 1 0 1856 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5190_6
timestamp 1731220342
transform 1 0 1760 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5189_6
timestamp 1731220342
transform 1 0 1664 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5188_6
timestamp 1731220342
transform 1 0 1568 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5187_6
timestamp 1731220342
transform 1 0 1472 0 -1 2936
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5186_6
timestamp 1731220342
transform 1 0 1424 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5185_6
timestamp 1731220342
transform 1 0 1544 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5184_6
timestamp 1731220342
transform 1 0 1664 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5183_6
timestamp 1731220342
transform 1 0 1896 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5182_6
timestamp 1731220342
transform 1 0 1792 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5181_6
timestamp 1731220342
transform 1 0 1744 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5180_6
timestamp 1731220342
transform 1 0 1568 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5179_6
timestamp 1731220342
transform 1 0 1896 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5178_6
timestamp 1731220342
transform 1 0 1896 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5177_6
timestamp 1731220342
transform 1 0 2064 0 -1 3144
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5176_6
timestamp 1731220342
transform 1 0 2064 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5175_6
timestamp 1731220342
transform 1 0 2536 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5174_6
timestamp 1731220342
transform 1 0 2368 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5173_6
timestamp 1731220342
transform 1 0 2200 0 1 3148
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5172_6
timestamp 1731220342
transform 1 0 2120 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5171_6
timestamp 1731220342
transform 1 0 2288 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5170_6
timestamp 1731220342
transform 1 0 2448 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5169_6
timestamp 1731220342
transform 1 0 2608 0 -1 3300
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5168_6
timestamp 1731220342
transform 1 0 2608 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5167_6
timestamp 1731220342
transform 1 0 2472 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5166_6
timestamp 1731220342
transform 1 0 2344 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5165_6
timestamp 1731220342
transform 1 0 2744 0 1 3304
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5164_6
timestamp 1731220342
transform 1 0 2776 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5163_6
timestamp 1731220342
transform 1 0 2888 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5162_6
timestamp 1731220342
transform 1 0 3008 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5161_6
timestamp 1731220342
transform 1 0 3096 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5160_6
timestamp 1731220342
transform 1 0 2976 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5159_6
timestamp 1731220342
transform 1 0 2864 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5158_6
timestamp 1731220342
transform 1 0 2760 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5157_6
timestamp 1731220342
transform 1 0 2664 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5156_6
timestamp 1731220342
transform 1 0 2672 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5155_6
timestamp 1731220342
transform 1 0 2576 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5154_6
timestamp 1731220342
transform 1 0 2480 0 -1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5153_6
timestamp 1731220342
transform 1 0 2568 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5152_6
timestamp 1731220342
transform 1 0 2472 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5151_6
timestamp 1731220342
transform 1 0 2376 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5150_6
timestamp 1731220342
transform 1 0 2280 0 1 3464
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5149_6
timestamp 1731220342
transform 1 0 2864 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5148_6
timestamp 1731220342
transform 1 0 2648 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5147_6
timestamp 1731220342
transform 1 0 2448 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5146_6
timestamp 1731220342
transform 1 0 2264 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5145_6
timestamp 1731220342
transform 1 0 2104 0 -1 3632
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5144_6
timestamp 1731220342
transform 1 0 2688 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5143_6
timestamp 1731220342
transform 1 0 2472 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5142_6
timestamp 1731220342
transform 1 0 2256 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5141_6
timestamp 1731220342
transform 1 0 2064 0 1 3636
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5140_6
timestamp 1731220342
transform 1 0 2064 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5139_6
timestamp 1731220342
transform 1 0 2192 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5138_6
timestamp 1731220342
transform 1 0 2368 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5137_6
timestamp 1731220342
transform 1 0 2744 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5136_6
timestamp 1731220342
transform 1 0 2552 0 -1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5135_6
timestamp 1731220342
transform 1 0 2512 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5134_6
timestamp 1731220342
transform 1 0 2376 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5133_6
timestamp 1731220342
transform 1 0 2248 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5132_6
timestamp 1731220342
transform 1 0 2824 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5131_6
timestamp 1731220342
transform 1 0 2664 0 1 3800
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5130_6
timestamp 1731220342
transform 1 0 2640 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5129_6
timestamp 1731220342
transform 1 0 2496 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5128_6
timestamp 1731220342
transform 1 0 2352 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5127_6
timestamp 1731220342
transform 1 0 2208 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5126_6
timestamp 1731220342
transform 1 0 2072 0 -1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5125_6
timestamp 1731220342
transform 1 0 2064 0 1 3952
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5124_6
timestamp 1731220342
transform 1 0 1896 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5123_6
timestamp 1731220342
transform 1 0 1768 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5122_6
timestamp 1731220342
transform 1 0 1616 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5121_6
timestamp 1731220342
transform 1 0 1464 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5120_6
timestamp 1731220342
transform 1 0 1304 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5119_6
timestamp 1731220342
transform 1 0 1144 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5118_6
timestamp 1731220342
transform 1 0 1456 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5117_6
timestamp 1731220342
transform 1 0 1320 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5116_6
timestamp 1731220342
transform 1 0 1192 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5115_6
timestamp 1731220342
transform 1 0 1064 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5114_6
timestamp 1731220342
transform 1 0 936 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5113_6
timestamp 1731220342
transform 1 0 1032 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5112_6
timestamp 1731220342
transform 1 0 1184 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5111_6
timestamp 1731220342
transform 1 0 1336 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5110_6
timestamp 1731220342
transform 1 0 1488 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5109_6
timestamp 1731220342
transform 1 0 1640 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5108_6
timestamp 1731220342
transform 1 0 1496 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5107_6
timestamp 1731220342
transform 1 0 1304 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5106_6
timestamp 1731220342
transform 1 0 1688 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5105_6
timestamp 1731220342
transform 1 0 1880 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5104_6
timestamp 1731220342
transform 1 0 1784 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5103_6
timestamp 1731220342
transform 1 0 1624 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5102_6
timestamp 1731220342
transform 1 0 1472 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5101_6
timestamp 1731220342
transform 1 0 1320 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_5100_6
timestamp 1731220342
transform 1 0 1168 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_599_6
timestamp 1731220342
transform 1 0 1536 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_598_6
timestamp 1731220342
transform 1 0 1368 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_597_6
timestamp 1731220342
transform 1 0 1208 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_596_6
timestamp 1731220342
transform 1 0 1048 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_595_6
timestamp 1731220342
transform 1 0 1360 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_594_6
timestamp 1731220342
transform 1 0 1224 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_593_6
timestamp 1731220342
transform 1 0 1088 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_592_6
timestamp 1731220342
transform 1 0 960 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_591_6
timestamp 1731220342
transform 1 0 824 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_590_6
timestamp 1731220342
transform 1 0 808 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_589_6
timestamp 1731220342
transform 1 0 960 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_588_6
timestamp 1731220342
transform 1 0 1264 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_587_6
timestamp 1731220342
transform 1 0 1112 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_586_6
timestamp 1731220342
transform 1 0 1080 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_585_6
timestamp 1731220342
transform 1 0 920 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_584_6
timestamp 1731220342
transform 1 0 1232 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_583_6
timestamp 1731220342
transform 1 0 1384 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_582_6
timestamp 1731220342
transform 1 0 1544 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_581_6
timestamp 1731220342
transform 1 0 1472 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_580_6
timestamp 1731220342
transform 1 0 1296 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_579_6
timestamp 1731220342
transform 1 0 1120 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_578_6
timestamp 1731220342
transform 1 0 952 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_577_6
timestamp 1731220342
transform 1 0 1680 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_576_6
timestamp 1731220342
transform 1 0 1448 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_575_6
timestamp 1731220342
transform 1 0 1224 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_574_6
timestamp 1731220342
transform 1 0 1024 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_573_6
timestamp 1731220342
transform 1 0 848 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_572_6
timestamp 1731220342
transform 1 0 1400 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_571_6
timestamp 1731220342
transform 1 0 1240 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_570_6
timestamp 1731220342
transform 1 0 1080 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_569_6
timestamp 1731220342
transform 1 0 936 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_568_6
timestamp 1731220342
transform 1 0 1304 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_567_6
timestamp 1731220342
transform 1 0 1176 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_566_6
timestamp 1731220342
transform 1 0 1048 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_565_6
timestamp 1731220342
transform 1 0 928 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_564_6
timestamp 1731220342
transform 1 0 808 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_563_6
timestamp 1731220342
transform 1 0 704 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_562_6
timestamp 1731220342
transform 1 0 608 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_561_6
timestamp 1731220342
transform 1 0 512 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_560_6
timestamp 1731220342
transform 1 0 416 0 1 2960
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_559_6
timestamp 1731220342
transform 1 0 800 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_558_6
timestamp 1731220342
transform 1 0 688 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_557_6
timestamp 1731220342
transform 1 0 592 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_556_6
timestamp 1731220342
transform 1 0 496 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_555_6
timestamp 1731220342
transform 1 0 400 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_554_6
timestamp 1731220342
transform 1 0 304 0 -1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_553_6
timestamp 1731220342
transform 1 0 696 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_552_6
timestamp 1731220342
transform 1 0 560 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_551_6
timestamp 1731220342
transform 1 0 424 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_550_6
timestamp 1731220342
transform 1 0 288 0 1 3112
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_549_6
timestamp 1731220342
transform 1 0 784 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_548_6
timestamp 1731220342
transform 1 0 616 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_547_6
timestamp 1731220342
transform 1 0 448 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_546_6
timestamp 1731220342
transform 1 0 288 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_545_6
timestamp 1731220342
transform 1 0 136 0 -1 3264
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_544_6
timestamp 1731220342
transform 1 0 760 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_543_6
timestamp 1731220342
transform 1 0 592 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_542_6
timestamp 1731220342
transform 1 0 424 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_541_6
timestamp 1731220342
transform 1 0 256 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_540_6
timestamp 1731220342
transform 1 0 128 0 1 3272
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_539_6
timestamp 1731220342
transform 1 0 128 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_538_6
timestamp 1731220342
transform 1 0 240 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_537_6
timestamp 1731220342
transform 1 0 664 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_536_6
timestamp 1731220342
transform 1 0 520 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_535_6
timestamp 1731220342
transform 1 0 376 0 -1 3432
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_534_6
timestamp 1731220342
transform 1 0 280 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_533_6
timestamp 1731220342
transform 1 0 152 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_532_6
timestamp 1731220342
transform 1 0 688 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_531_6
timestamp 1731220342
transform 1 0 552 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_530_6
timestamp 1731220342
transform 1 0 416 0 1 3440
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_529_6
timestamp 1731220342
transform 1 0 408 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_528_6
timestamp 1731220342
transform 1 0 264 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_527_6
timestamp 1731220342
transform 1 0 888 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_526_6
timestamp 1731220342
transform 1 0 728 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_525_6
timestamp 1731220342
transform 1 0 568 0 -1 3600
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_524_6
timestamp 1731220342
transform 1 0 512 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_523_6
timestamp 1731220342
transform 1 0 360 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_522_6
timestamp 1731220342
transform 1 0 672 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_521_6
timestamp 1731220342
transform 1 0 840 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_520_6
timestamp 1731220342
transform 1 0 1008 0 1 3608
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_519_6
timestamp 1731220342
transform 1 0 1120 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_518_6
timestamp 1731220342
transform 1 0 928 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_517_6
timestamp 1731220342
transform 1 0 744 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_516_6
timestamp 1731220342
transform 1 0 560 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_515_6
timestamp 1731220342
transform 1 0 392 0 -1 3772
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_514_6
timestamp 1731220342
transform 1 0 880 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_513_6
timestamp 1731220342
transform 1 0 720 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_512_6
timestamp 1731220342
transform 1 0 560 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_511_6
timestamp 1731220342
transform 1 0 408 0 1 3776
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_510_6
timestamp 1731220342
transform 1 0 808 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_59_6
timestamp 1731220342
transform 1 0 680 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_58_6
timestamp 1731220342
transform 1 0 544 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_57_6
timestamp 1731220342
transform 1 0 416 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_56_6
timestamp 1731220342
transform 1 0 296 0 -1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_55_6
timestamp 1731220342
transform 1 0 968 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_54_6
timestamp 1731220342
transform 1 0 784 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_53_6
timestamp 1731220342
transform 1 0 600 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_52_6
timestamp 1731220342
transform 1 0 424 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_51_6
timestamp 1731220342
transform 1 0 272 0 1 3932
box 8 5 92 72
use _0_0cell_0_0gcelem3x0  tst_50_6
timestamp 1731220342
transform 1 0 144 0 1 3932
box 8 5 92 72
<< end >>
