magic
tech sky130l
timestamp 1731220628
<< m1 >>
rect 456 2123 460 2143
rect 544 2123 548 2163
rect 624 2123 628 2143
rect 688 2123 692 2143
rect 736 2051 740 2071
rect 896 2051 900 2071
rect 984 2051 988 2071
rect 1192 2027 1196 2047
rect 1248 2027 1252 2047
rect 1432 2027 1436 2047
rect 1792 2027 1796 2047
rect 1864 2027 1868 2047
rect 1488 1991 1492 2011
rect 2008 1991 2012 2023
rect 792 1943 796 1963
rect 280 1855 284 1915
rect 1520 1911 1524 1931
rect 1664 1911 1668 1931
rect 1736 1911 1740 1931
rect 1808 1911 1812 1931
rect 1880 1911 1884 1931
rect 1360 1875 1364 1895
rect 640 1791 644 1811
rect 2048 1803 2052 1871
rect 1584 1759 1588 1779
rect 808 1707 812 1735
rect 856 1715 860 1735
rect 496 1675 500 1695
rect 720 1675 724 1695
rect 1864 1687 1868 1707
rect 1928 1687 1932 1707
rect 1992 1687 1996 1707
rect 1456 1651 1460 1671
rect 1960 1651 1964 1671
rect 1232 1579 1236 1599
rect 216 1559 220 1579
rect 400 1559 404 1579
rect 1608 1547 1612 1563
rect 1800 1471 1804 1491
rect 1888 1471 1892 1491
rect 736 1439 740 1459
rect 728 1367 732 1387
rect 792 1367 796 1387
rect 712 1331 716 1351
rect 2016 1323 2020 1343
rect 800 1255 804 1283
rect 936 1263 940 1283
rect 1232 1251 1236 1271
rect 1912 1251 1916 1271
rect 392 1223 396 1243
rect 640 1223 644 1243
rect 1312 1211 1316 1231
rect 1408 1215 1412 1231
rect 1648 1215 1652 1231
rect 1664 1191 1668 1207
rect 344 1119 348 1139
rect 1400 1135 1404 1163
rect 232 1043 236 1063
rect 280 1043 284 1063
rect 400 1043 404 1063
rect 1880 1031 1884 1051
rect 1960 1031 1964 1051
rect 304 1003 308 1023
rect 2048 927 2052 947
rect 448 895 452 915
rect 384 823 388 843
rect 808 823 812 843
rect 204 791 212 795
rect 208 787 212 791
rect 208 783 216 787
rect 248 719 252 783
rect 616 743 620 807
rect 1536 775 1540 795
rect 480 719 484 739
rect 1840 707 1844 727
rect 1936 707 1940 727
rect 744 679 748 699
rect 856 679 860 699
rect 1424 667 1428 687
rect 1808 667 1812 687
rect 488 603 492 623
rect 1032 563 1036 583
rect 200 487 204 507
rect 464 487 468 507
rect 792 487 796 507
rect 1376 491 1380 511
rect 272 451 276 471
rect 784 455 788 483
rect 264 383 268 403
rect 400 383 404 403
rect 456 383 460 403
rect 1856 387 1860 407
rect 256 323 260 379
rect 616 351 620 367
rect 1952 347 1956 367
rect 192 275 196 295
rect 504 275 508 295
rect 656 275 660 295
rect 784 275 788 295
rect 840 275 844 295
rect 1280 275 1284 295
rect 1656 263 1660 295
rect 2048 275 2052 295
rect 472 239 476 259
rect 680 239 684 259
rect 360 167 364 187
rect 1232 163 1236 183
rect 1640 163 1644 183
rect 1704 163 1708 183
rect 912 107 916 127
rect 1888 107 1892 127
<< m2c >>
rect 1684 2219 1688 2223
rect 1724 2219 1728 2223
rect 1764 2219 1768 2223
rect 1804 2219 1808 2223
rect 1712 2195 1716 2199
rect 1752 2195 1756 2199
rect 1792 2195 1796 2199
rect 1832 2195 1836 2199
rect 160 2187 164 2191
rect 200 2187 204 2191
rect 240 2187 244 2191
rect 280 2187 284 2191
rect 344 2187 348 2191
rect 408 2187 412 2191
rect 472 2187 476 2191
rect 536 2187 540 2191
rect 600 2187 604 2191
rect 656 2187 660 2191
rect 712 2187 716 2191
rect 760 2187 764 2191
rect 816 2187 820 2191
rect 872 2187 876 2191
rect 928 2187 932 2191
rect 172 2163 176 2167
rect 212 2163 216 2167
rect 252 2163 256 2167
rect 316 2163 320 2167
rect 380 2163 384 2167
rect 444 2163 448 2167
rect 508 2163 512 2167
rect 544 2163 548 2167
rect 572 2163 576 2167
rect 628 2163 632 2167
rect 684 2163 688 2167
rect 732 2163 736 2167
rect 788 2163 792 2167
rect 844 2163 848 2167
rect 900 2163 904 2167
rect 228 2145 232 2149
rect 268 2143 272 2147
rect 308 2143 312 2147
rect 356 2143 360 2147
rect 420 2143 424 2147
rect 456 2143 460 2147
rect 484 2143 488 2147
rect 256 2121 260 2125
rect 1184 2151 1188 2155
rect 1224 2151 1228 2155
rect 1264 2151 1268 2155
rect 1304 2151 1308 2155
rect 1360 2151 1364 2155
rect 1416 2151 1420 2155
rect 1480 2151 1484 2155
rect 1552 2151 1556 2155
rect 1616 2151 1620 2155
rect 1688 2151 1692 2155
rect 1760 2151 1764 2155
rect 1832 2151 1836 2155
rect 1904 2151 1908 2155
rect 556 2143 560 2147
rect 624 2143 628 2147
rect 636 2143 640 2147
rect 688 2143 692 2147
rect 716 2143 720 2147
rect 796 2145 800 2149
rect 876 2143 880 2147
rect 964 2143 968 2147
rect 1156 2127 1160 2131
rect 1196 2127 1200 2131
rect 1236 2127 1240 2131
rect 1276 2127 1280 2131
rect 1332 2127 1336 2131
rect 1388 2127 1392 2131
rect 1452 2127 1456 2131
rect 1524 2127 1528 2131
rect 1588 2127 1592 2131
rect 1660 2127 1664 2131
rect 1732 2127 1736 2131
rect 1804 2127 1808 2131
rect 1876 2127 1880 2131
rect 296 2119 300 2123
rect 336 2119 340 2123
rect 384 2119 388 2123
rect 448 2119 452 2123
rect 456 2119 460 2123
rect 512 2119 516 2123
rect 544 2119 548 2123
rect 584 2119 588 2123
rect 624 2119 628 2123
rect 664 2119 668 2123
rect 688 2119 692 2123
rect 744 2119 748 2123
rect 824 2119 828 2123
rect 904 2121 908 2125
rect 992 2119 996 2123
rect 1156 2115 1160 2119
rect 1196 2115 1200 2119
rect 1236 2115 1240 2119
rect 1292 2115 1296 2119
rect 1364 2115 1368 2119
rect 1436 2115 1440 2119
rect 1516 2115 1520 2119
rect 1596 2115 1600 2119
rect 1676 2115 1680 2119
rect 1748 2115 1752 2119
rect 1820 2115 1824 2119
rect 1884 2115 1888 2119
rect 1948 2115 1952 2119
rect 2020 2115 2024 2119
rect 2068 2115 2072 2119
rect 1184 2091 1188 2095
rect 1224 2091 1228 2095
rect 1264 2091 1268 2095
rect 1320 2091 1324 2095
rect 1392 2091 1396 2095
rect 1464 2091 1468 2095
rect 1544 2091 1548 2095
rect 1624 2091 1628 2095
rect 1704 2091 1708 2095
rect 1776 2091 1780 2095
rect 1848 2091 1852 2095
rect 1912 2091 1916 2095
rect 1976 2091 1980 2095
rect 2048 2091 2052 2095
rect 2096 2091 2100 2095
rect 328 2071 332 2075
rect 376 2071 380 2075
rect 432 2071 436 2075
rect 496 2071 500 2075
rect 568 2071 572 2075
rect 648 2071 652 2075
rect 728 2071 732 2075
rect 736 2071 740 2075
rect 808 2071 812 2075
rect 888 2071 892 2075
rect 896 2071 900 2075
rect 976 2071 980 2075
rect 984 2071 988 2075
rect 1064 2071 1068 2075
rect 300 2047 304 2051
rect 348 2047 352 2051
rect 404 2047 408 2051
rect 468 2047 472 2051
rect 540 2047 544 2051
rect 620 2047 624 2051
rect 700 2047 704 2051
rect 736 2047 740 2051
rect 780 2047 784 2051
rect 860 2047 864 2051
rect 896 2047 900 2051
rect 948 2047 952 2051
rect 984 2047 988 2051
rect 1036 2047 1040 2051
rect 1184 2047 1188 2051
rect 1192 2047 1196 2051
rect 1240 2047 1244 2051
rect 1248 2047 1252 2051
rect 1328 2047 1332 2051
rect 1424 2047 1428 2051
rect 1432 2047 1436 2051
rect 1520 2047 1524 2051
rect 1616 2047 1620 2051
rect 1704 2047 1708 2051
rect 1784 2047 1788 2051
rect 1792 2047 1796 2051
rect 1856 2047 1860 2051
rect 1864 2047 1868 2051
rect 1920 2047 1924 2051
rect 1984 2047 1988 2051
rect 2048 2047 2052 2051
rect 2096 2047 2100 2051
rect 180 2031 184 2035
rect 276 2031 280 2035
rect 372 2031 376 2035
rect 460 2031 464 2035
rect 540 2033 544 2037
rect 620 2031 624 2035
rect 692 2031 696 2035
rect 756 2031 760 2035
rect 812 2031 816 2035
rect 860 2031 864 2035
rect 908 2031 912 2035
rect 956 2031 960 2035
rect 1004 2031 1008 2035
rect 1044 2031 1048 2035
rect 1156 2023 1160 2027
rect 1192 2023 1196 2027
rect 1212 2023 1216 2027
rect 1248 2023 1252 2027
rect 1300 2023 1304 2027
rect 1396 2023 1400 2027
rect 1432 2023 1436 2027
rect 1492 2023 1496 2027
rect 1588 2023 1592 2027
rect 1676 2023 1680 2027
rect 1756 2023 1760 2027
rect 1792 2023 1796 2027
rect 1828 2023 1832 2027
rect 1864 2023 1868 2027
rect 1892 2023 1896 2027
rect 1956 2023 1960 2027
rect 2008 2023 2012 2027
rect 2020 2023 2024 2027
rect 2068 2023 2072 2027
rect 1156 2011 1160 2015
rect 1236 2011 1240 2015
rect 1348 2011 1352 2015
rect 1452 2011 1456 2015
rect 1488 2011 1492 2015
rect 1556 2011 1560 2015
rect 1652 2011 1656 2015
rect 1740 2011 1744 2015
rect 1820 2011 1824 2015
rect 1892 2011 1896 2015
rect 1956 2011 1960 2015
rect 208 2007 212 2011
rect 304 2007 308 2011
rect 400 2007 404 2011
rect 488 2007 492 2011
rect 568 2007 572 2011
rect 648 2007 652 2011
rect 720 2007 724 2011
rect 784 2007 788 2011
rect 840 2007 844 2011
rect 888 2007 892 2011
rect 936 2007 940 2011
rect 984 2007 988 2011
rect 1032 2007 1036 2011
rect 1072 2007 1076 2011
rect 2020 2011 2024 2015
rect 2068 2011 2072 2015
rect 1184 1987 1188 1991
rect 1264 1987 1268 1991
rect 1376 1987 1380 1991
rect 1480 1987 1484 1991
rect 1488 1987 1492 1991
rect 1584 1987 1588 1991
rect 1680 1987 1684 1991
rect 1768 1987 1772 1991
rect 1848 1987 1852 1991
rect 1920 1987 1924 1991
rect 1984 1987 1988 1991
rect 2008 1987 2012 1991
rect 2048 1987 2052 1991
rect 2096 1987 2100 1991
rect 184 1963 188 1967
rect 256 1963 260 1967
rect 328 1963 332 1967
rect 400 1963 404 1967
rect 472 1963 476 1967
rect 552 1963 556 1967
rect 632 1963 636 1967
rect 712 1963 716 1967
rect 784 1963 788 1967
rect 792 1963 796 1967
rect 856 1963 860 1967
rect 936 1963 940 1967
rect 1016 1963 1020 1967
rect 156 1939 160 1943
rect 228 1939 232 1943
rect 300 1939 304 1943
rect 372 1939 376 1943
rect 444 1939 448 1943
rect 524 1939 528 1943
rect 604 1939 608 1943
rect 684 1939 688 1943
rect 756 1939 760 1943
rect 792 1939 796 1943
rect 828 1939 832 1943
rect 908 1939 912 1943
rect 988 1939 992 1943
rect 1384 1931 1388 1935
rect 1448 1931 1452 1935
rect 1512 1931 1516 1935
rect 1520 1931 1524 1935
rect 1584 1931 1588 1935
rect 1656 1931 1660 1935
rect 1664 1931 1668 1935
rect 1728 1931 1732 1935
rect 1736 1931 1740 1935
rect 1800 1931 1804 1935
rect 1808 1931 1812 1935
rect 1872 1931 1876 1935
rect 1880 1931 1884 1935
rect 1952 1931 1956 1935
rect 2032 1931 2036 1935
rect 2096 1931 2100 1935
rect 132 1925 136 1929
rect 172 1923 176 1927
rect 228 1923 232 1927
rect 292 1923 296 1927
rect 364 1923 368 1927
rect 444 1923 448 1927
rect 524 1925 528 1929
rect 612 1923 616 1927
rect 700 1923 704 1927
rect 788 1923 792 1927
rect 876 1923 880 1927
rect 280 1915 284 1919
rect 160 1899 164 1903
rect 200 1899 204 1903
rect 256 1899 260 1903
rect 1356 1907 1360 1911
rect 1420 1907 1424 1911
rect 1484 1907 1488 1911
rect 1520 1907 1524 1911
rect 1556 1907 1560 1911
rect 1628 1907 1632 1911
rect 1664 1907 1668 1911
rect 1700 1907 1704 1911
rect 1736 1907 1740 1911
rect 1772 1907 1776 1911
rect 1808 1907 1812 1911
rect 1844 1907 1848 1911
rect 1880 1907 1884 1911
rect 1924 1907 1928 1911
rect 2004 1907 2008 1911
rect 2068 1907 2072 1911
rect 320 1899 324 1903
rect 392 1899 396 1903
rect 472 1899 476 1903
rect 552 1899 556 1903
rect 640 1899 644 1903
rect 728 1899 732 1903
rect 816 1899 820 1903
rect 904 1899 908 1903
rect 1228 1897 1232 1901
rect 1268 1895 1272 1899
rect 1316 1895 1320 1899
rect 1360 1895 1364 1899
rect 1372 1897 1376 1901
rect 1436 1895 1440 1899
rect 1500 1895 1504 1899
rect 1572 1895 1576 1899
rect 1652 1895 1656 1899
rect 1748 1895 1752 1899
rect 1860 1895 1864 1899
rect 1972 1895 1976 1899
rect 2068 1895 2072 1899
rect 1256 1871 1260 1875
rect 1296 1871 1300 1875
rect 1344 1871 1348 1875
rect 1360 1871 1364 1875
rect 1400 1871 1404 1875
rect 1464 1871 1468 1875
rect 1528 1871 1532 1875
rect 1600 1871 1604 1875
rect 1680 1871 1684 1875
rect 1776 1871 1780 1875
rect 1888 1871 1892 1875
rect 2000 1871 2004 1875
rect 2048 1871 2052 1875
rect 2096 1871 2100 1875
rect 160 1851 164 1855
rect 200 1851 204 1855
rect 248 1851 252 1855
rect 280 1851 284 1855
rect 312 1851 316 1855
rect 384 1851 388 1855
rect 456 1851 460 1855
rect 528 1851 532 1855
rect 592 1851 596 1855
rect 656 1851 660 1855
rect 720 1851 724 1855
rect 784 1851 788 1855
rect 856 1851 860 1855
rect 132 1827 136 1831
rect 172 1827 176 1831
rect 220 1827 224 1831
rect 284 1827 288 1831
rect 356 1827 360 1831
rect 428 1827 432 1831
rect 500 1827 504 1831
rect 564 1827 568 1831
rect 628 1827 632 1831
rect 692 1827 696 1831
rect 756 1827 760 1831
rect 828 1827 832 1831
rect 1184 1823 1188 1827
rect 1224 1823 1228 1827
rect 1264 1823 1268 1827
rect 1328 1823 1332 1827
rect 1392 1823 1396 1827
rect 1456 1823 1460 1827
rect 1528 1823 1532 1827
rect 1608 1823 1612 1827
rect 1696 1823 1700 1827
rect 1792 1823 1796 1827
rect 1896 1823 1900 1827
rect 2008 1823 2012 1827
rect 132 1811 136 1815
rect 180 1811 184 1815
rect 260 1813 264 1817
rect 348 1811 352 1815
rect 436 1811 440 1815
rect 524 1811 528 1815
rect 604 1811 608 1815
rect 640 1811 644 1815
rect 684 1811 688 1815
rect 764 1811 768 1815
rect 836 1813 840 1817
rect 908 1811 912 1815
rect 988 1811 992 1815
rect 1044 1811 1048 1815
rect 1156 1801 1160 1805
rect 1196 1801 1200 1805
rect 2096 1823 2100 1827
rect 1236 1799 1240 1803
rect 1300 1799 1304 1803
rect 1364 1799 1368 1803
rect 1428 1799 1432 1803
rect 1500 1799 1504 1803
rect 1580 1799 1584 1803
rect 1668 1799 1672 1803
rect 1764 1799 1768 1803
rect 1868 1799 1872 1803
rect 1980 1799 1984 1803
rect 2048 1799 2052 1803
rect 2068 1799 2072 1803
rect 160 1787 164 1791
rect 208 1787 212 1791
rect 288 1787 292 1791
rect 376 1787 380 1791
rect 464 1787 468 1791
rect 552 1787 556 1791
rect 632 1787 636 1791
rect 640 1787 644 1791
rect 712 1787 716 1791
rect 792 1787 796 1791
rect 864 1787 868 1791
rect 936 1787 940 1791
rect 1016 1787 1020 1791
rect 1072 1787 1076 1791
rect 1308 1779 1312 1783
rect 1348 1779 1352 1783
rect 1388 1779 1392 1783
rect 1428 1779 1432 1783
rect 1468 1779 1472 1783
rect 1508 1779 1512 1783
rect 1548 1779 1552 1783
rect 1584 1779 1588 1783
rect 1604 1779 1608 1783
rect 1676 1779 1680 1783
rect 1764 1779 1768 1783
rect 1868 1779 1872 1783
rect 1980 1779 1984 1783
rect 2068 1779 2072 1783
rect 1336 1755 1340 1759
rect 1376 1755 1380 1759
rect 1416 1755 1420 1759
rect 1456 1755 1460 1759
rect 1496 1755 1500 1759
rect 1536 1755 1540 1759
rect 1576 1755 1580 1759
rect 1584 1755 1588 1759
rect 1632 1755 1636 1759
rect 1704 1755 1708 1759
rect 1792 1755 1796 1759
rect 1896 1755 1900 1759
rect 2008 1755 2012 1759
rect 2096 1755 2100 1759
rect 160 1735 164 1739
rect 224 1735 228 1739
rect 320 1735 324 1739
rect 424 1735 428 1739
rect 520 1735 524 1739
rect 616 1735 620 1739
rect 696 1735 700 1739
rect 776 1735 780 1739
rect 808 1735 812 1739
rect 848 1735 852 1739
rect 856 1735 860 1739
rect 912 1735 916 1739
rect 984 1735 988 1739
rect 1056 1735 1060 1739
rect 132 1711 136 1715
rect 196 1711 200 1715
rect 292 1711 296 1715
rect 396 1711 400 1715
rect 492 1711 496 1715
rect 588 1711 592 1715
rect 668 1711 672 1715
rect 748 1711 752 1715
rect 820 1711 824 1715
rect 856 1711 860 1715
rect 884 1711 888 1715
rect 956 1711 960 1715
rect 1028 1711 1032 1715
rect 1288 1707 1292 1711
rect 1344 1707 1348 1711
rect 1408 1707 1412 1711
rect 1480 1707 1484 1711
rect 1560 1707 1564 1711
rect 1640 1707 1644 1711
rect 1712 1707 1716 1711
rect 1784 1707 1788 1711
rect 1856 1707 1860 1711
rect 1864 1707 1868 1711
rect 1920 1707 1924 1711
rect 1928 1707 1932 1711
rect 1984 1707 1988 1711
rect 1992 1707 1996 1711
rect 2048 1707 2052 1711
rect 2096 1707 2100 1711
rect 808 1703 812 1707
rect 148 1695 152 1699
rect 220 1697 224 1701
rect 300 1695 304 1699
rect 380 1695 384 1699
rect 460 1695 464 1699
rect 496 1695 500 1699
rect 532 1695 536 1699
rect 604 1695 608 1699
rect 668 1695 672 1699
rect 720 1695 724 1699
rect 732 1695 736 1699
rect 804 1695 808 1699
rect 876 1695 880 1699
rect 1260 1683 1264 1687
rect 1316 1683 1320 1687
rect 1380 1683 1384 1687
rect 1452 1683 1456 1687
rect 1532 1683 1536 1687
rect 1612 1683 1616 1687
rect 1684 1683 1688 1687
rect 1756 1683 1760 1687
rect 1828 1683 1832 1687
rect 1864 1683 1868 1687
rect 1892 1683 1896 1687
rect 1928 1683 1932 1687
rect 1956 1683 1960 1687
rect 1992 1683 1996 1687
rect 2020 1683 2024 1687
rect 2068 1683 2072 1687
rect 176 1671 180 1675
rect 248 1671 252 1675
rect 328 1671 332 1675
rect 408 1671 412 1675
rect 488 1671 492 1675
rect 496 1671 500 1675
rect 560 1671 564 1675
rect 632 1671 636 1675
rect 696 1671 700 1675
rect 720 1671 724 1675
rect 760 1671 764 1675
rect 832 1671 836 1675
rect 904 1671 908 1675
rect 1164 1671 1168 1675
rect 1244 1671 1248 1675
rect 1332 1671 1336 1675
rect 1420 1671 1424 1675
rect 1456 1671 1460 1675
rect 1508 1671 1512 1675
rect 1596 1671 1600 1675
rect 1676 1671 1680 1675
rect 1748 1671 1752 1675
rect 1812 1671 1816 1675
rect 1868 1671 1872 1675
rect 1924 1671 1928 1675
rect 1960 1671 1964 1675
rect 1980 1671 1984 1675
rect 2028 1671 2032 1675
rect 2068 1671 2072 1675
rect 1192 1647 1196 1651
rect 1272 1647 1276 1651
rect 1360 1647 1364 1651
rect 1448 1647 1452 1651
rect 1456 1647 1460 1651
rect 1536 1647 1540 1651
rect 1624 1647 1628 1651
rect 1704 1647 1708 1651
rect 1776 1647 1780 1651
rect 1840 1647 1844 1651
rect 1896 1647 1900 1651
rect 1952 1647 1956 1651
rect 1960 1647 1964 1651
rect 2008 1647 2012 1651
rect 2056 1647 2060 1651
rect 2096 1647 2100 1651
rect 200 1623 204 1627
rect 240 1623 244 1627
rect 280 1623 284 1627
rect 328 1623 332 1627
rect 384 1623 388 1627
rect 432 1623 436 1627
rect 480 1623 484 1627
rect 528 1623 532 1627
rect 576 1623 580 1627
rect 632 1623 636 1627
rect 688 1623 692 1627
rect 744 1623 748 1627
rect 172 1599 176 1603
rect 212 1599 216 1603
rect 252 1599 256 1603
rect 300 1599 304 1603
rect 356 1599 360 1603
rect 404 1599 408 1603
rect 452 1599 456 1603
rect 500 1599 504 1603
rect 548 1599 552 1603
rect 604 1599 608 1603
rect 660 1599 664 1603
rect 716 1599 720 1603
rect 1184 1599 1188 1603
rect 1224 1599 1228 1603
rect 1232 1599 1236 1603
rect 1272 1599 1276 1603
rect 1344 1599 1348 1603
rect 1416 1599 1420 1603
rect 1488 1599 1492 1603
rect 1560 1599 1564 1603
rect 1632 1599 1636 1603
rect 1704 1599 1708 1603
rect 1776 1599 1780 1603
rect 1856 1599 1860 1603
rect 140 1579 144 1583
rect 180 1579 184 1583
rect 216 1579 220 1583
rect 228 1579 232 1583
rect 284 1579 288 1583
rect 348 1579 352 1583
rect 400 1579 404 1583
rect 412 1579 416 1583
rect 476 1581 480 1585
rect 540 1579 544 1583
rect 604 1579 608 1583
rect 660 1579 664 1583
rect 724 1579 728 1583
rect 788 1579 792 1583
rect 852 1579 856 1583
rect 1156 1575 1160 1579
rect 1196 1575 1200 1579
rect 1232 1575 1236 1579
rect 1244 1575 1248 1579
rect 1316 1575 1320 1579
rect 1388 1575 1392 1579
rect 1460 1575 1464 1579
rect 1532 1575 1536 1579
rect 1604 1575 1608 1579
rect 1676 1575 1680 1579
rect 1748 1575 1752 1579
rect 1828 1575 1832 1579
rect 1236 1563 1240 1567
rect 1276 1563 1280 1567
rect 1324 1563 1328 1567
rect 1372 1563 1376 1567
rect 1420 1563 1424 1567
rect 1468 1565 1472 1569
rect 1516 1563 1520 1567
rect 1564 1563 1568 1567
rect 1608 1563 1612 1567
rect 1620 1563 1624 1567
rect 1676 1563 1680 1567
rect 1732 1563 1736 1567
rect 168 1555 172 1559
rect 208 1555 212 1559
rect 216 1555 220 1559
rect 256 1555 260 1559
rect 312 1555 316 1559
rect 376 1555 380 1559
rect 400 1555 404 1559
rect 440 1555 444 1559
rect 504 1555 508 1559
rect 568 1555 572 1559
rect 632 1555 636 1559
rect 688 1555 692 1559
rect 752 1555 756 1559
rect 816 1555 820 1559
rect 880 1555 884 1559
rect 1608 1543 1612 1547
rect 1264 1539 1268 1543
rect 1304 1539 1308 1543
rect 1352 1539 1356 1543
rect 1400 1539 1404 1543
rect 1448 1539 1452 1543
rect 1496 1539 1500 1543
rect 1544 1539 1548 1543
rect 1592 1539 1596 1543
rect 1648 1539 1652 1543
rect 1704 1539 1708 1543
rect 1760 1539 1764 1543
rect 160 1503 164 1507
rect 200 1503 204 1507
rect 240 1503 244 1507
rect 280 1503 284 1507
rect 320 1503 324 1507
rect 360 1503 364 1507
rect 400 1503 404 1507
rect 440 1503 444 1507
rect 480 1503 484 1507
rect 520 1503 524 1507
rect 560 1503 564 1507
rect 600 1503 604 1507
rect 640 1503 644 1507
rect 680 1503 684 1507
rect 720 1503 724 1507
rect 760 1503 764 1507
rect 800 1503 804 1507
rect 856 1503 860 1507
rect 912 1503 916 1507
rect 1344 1491 1348 1495
rect 1384 1491 1388 1495
rect 1424 1491 1428 1495
rect 1464 1491 1468 1495
rect 1504 1491 1508 1495
rect 1544 1491 1548 1495
rect 1584 1491 1588 1495
rect 1632 1491 1636 1495
rect 1688 1491 1692 1495
rect 1760 1491 1764 1495
rect 1800 1491 1804 1495
rect 1840 1491 1844 1495
rect 1888 1491 1892 1495
rect 1928 1491 1932 1495
rect 2016 1491 2020 1495
rect 2096 1491 2100 1495
rect 132 1479 136 1483
rect 172 1479 176 1483
rect 212 1479 216 1483
rect 252 1479 256 1483
rect 292 1479 296 1483
rect 332 1479 336 1483
rect 372 1479 376 1483
rect 412 1479 416 1483
rect 452 1479 456 1483
rect 492 1479 496 1483
rect 532 1479 536 1483
rect 572 1479 576 1483
rect 612 1479 616 1483
rect 652 1479 656 1483
rect 692 1479 696 1483
rect 732 1479 736 1483
rect 772 1479 776 1483
rect 828 1479 832 1483
rect 884 1479 888 1483
rect 1316 1467 1320 1471
rect 1356 1467 1360 1471
rect 1396 1467 1400 1471
rect 1436 1467 1440 1471
rect 1476 1467 1480 1471
rect 1516 1467 1520 1471
rect 1556 1467 1560 1471
rect 1604 1467 1608 1471
rect 1660 1467 1664 1471
rect 1732 1467 1736 1471
rect 1800 1467 1804 1471
rect 1812 1467 1816 1471
rect 1888 1467 1892 1471
rect 1900 1467 1904 1471
rect 1988 1467 1992 1471
rect 2068 1467 2072 1471
rect 516 1461 520 1465
rect 556 1459 560 1463
rect 596 1459 600 1463
rect 644 1461 648 1465
rect 692 1459 696 1463
rect 736 1459 740 1463
rect 748 1459 752 1463
rect 804 1459 808 1463
rect 868 1459 872 1463
rect 932 1459 936 1463
rect 1228 1455 1232 1459
rect 1276 1455 1280 1459
rect 1332 1455 1336 1459
rect 1388 1455 1392 1459
rect 1452 1455 1456 1459
rect 1516 1455 1520 1459
rect 1580 1455 1584 1459
rect 1644 1455 1648 1459
rect 1716 1455 1720 1459
rect 1804 1455 1808 1459
rect 1892 1455 1896 1459
rect 1988 1455 1992 1459
rect 2068 1455 2072 1459
rect 544 1435 548 1439
rect 584 1435 588 1439
rect 624 1435 628 1439
rect 672 1435 676 1439
rect 720 1435 724 1439
rect 736 1435 740 1439
rect 776 1437 780 1441
rect 832 1435 836 1439
rect 896 1435 900 1439
rect 960 1435 964 1439
rect 1256 1431 1260 1435
rect 1304 1431 1308 1435
rect 1360 1431 1364 1435
rect 1416 1431 1420 1435
rect 1480 1431 1484 1435
rect 1544 1431 1548 1435
rect 1608 1431 1612 1435
rect 1672 1431 1676 1435
rect 1744 1431 1748 1435
rect 1832 1431 1836 1435
rect 1920 1431 1924 1435
rect 2016 1431 2020 1435
rect 2096 1431 2100 1435
rect 456 1387 460 1391
rect 496 1387 500 1391
rect 544 1387 548 1391
rect 600 1387 604 1391
rect 656 1387 660 1391
rect 720 1387 724 1391
rect 728 1387 732 1391
rect 784 1387 788 1391
rect 792 1387 796 1391
rect 848 1387 852 1391
rect 920 1387 924 1391
rect 992 1387 996 1391
rect 1184 1383 1188 1387
rect 1224 1383 1228 1387
rect 1288 1383 1292 1387
rect 1376 1383 1380 1387
rect 1472 1383 1476 1387
rect 1568 1383 1572 1387
rect 1656 1383 1660 1387
rect 1744 1383 1748 1387
rect 1824 1383 1828 1387
rect 1896 1383 1900 1387
rect 1968 1383 1972 1387
rect 2040 1383 2044 1387
rect 2096 1383 2100 1387
rect 428 1363 432 1367
rect 468 1363 472 1367
rect 516 1363 520 1367
rect 572 1363 576 1367
rect 628 1363 632 1367
rect 692 1363 696 1367
rect 728 1363 732 1367
rect 756 1363 760 1367
rect 792 1363 796 1367
rect 820 1363 824 1367
rect 892 1363 896 1367
rect 964 1363 968 1367
rect 1156 1359 1160 1363
rect 1196 1359 1200 1363
rect 1260 1359 1264 1363
rect 1348 1359 1352 1363
rect 1444 1359 1448 1363
rect 1540 1359 1544 1363
rect 1628 1359 1632 1363
rect 1716 1359 1720 1363
rect 1796 1359 1800 1363
rect 1868 1359 1872 1363
rect 1940 1359 1944 1363
rect 2012 1359 2016 1363
rect 2068 1359 2072 1363
rect 372 1351 376 1355
rect 420 1351 424 1355
rect 476 1351 480 1355
rect 540 1351 544 1355
rect 604 1351 608 1355
rect 668 1351 672 1355
rect 712 1351 716 1355
rect 732 1351 736 1355
rect 796 1351 800 1355
rect 860 1351 864 1355
rect 924 1351 928 1355
rect 996 1351 1000 1355
rect 1044 1351 1048 1355
rect 1156 1343 1160 1347
rect 1252 1343 1256 1347
rect 1372 1343 1376 1347
rect 1484 1343 1488 1347
rect 1588 1345 1592 1349
rect 1676 1343 1680 1347
rect 1756 1343 1760 1347
rect 1828 1343 1832 1347
rect 1900 1345 1904 1349
rect 1964 1343 1968 1347
rect 2016 1343 2020 1347
rect 2028 1343 2032 1347
rect 2068 1343 2072 1347
rect 400 1327 404 1331
rect 448 1327 452 1331
rect 504 1327 508 1331
rect 568 1327 572 1331
rect 632 1327 636 1331
rect 696 1327 700 1331
rect 712 1327 716 1331
rect 760 1327 764 1331
rect 824 1327 828 1331
rect 888 1327 892 1331
rect 952 1327 956 1331
rect 1024 1327 1028 1331
rect 1072 1327 1076 1331
rect 1184 1319 1188 1323
rect 1280 1319 1284 1323
rect 1400 1319 1404 1323
rect 1512 1319 1516 1323
rect 1616 1319 1620 1323
rect 1704 1319 1708 1323
rect 1784 1319 1788 1323
rect 1856 1319 1860 1323
rect 1928 1319 1932 1323
rect 1992 1319 1996 1323
rect 2016 1319 2020 1323
rect 2056 1319 2060 1323
rect 2096 1319 2100 1323
rect 360 1283 364 1287
rect 416 1283 420 1287
rect 480 1283 484 1287
rect 552 1283 556 1287
rect 624 1283 628 1287
rect 696 1283 700 1287
rect 768 1283 772 1287
rect 800 1283 804 1287
rect 848 1283 852 1287
rect 928 1283 932 1287
rect 936 1283 940 1287
rect 1008 1283 1012 1287
rect 1072 1283 1076 1287
rect 332 1259 336 1263
rect 388 1259 392 1263
rect 452 1259 456 1263
rect 524 1259 528 1263
rect 596 1259 600 1263
rect 668 1259 672 1263
rect 740 1259 744 1263
rect 1184 1271 1188 1275
rect 1224 1271 1228 1275
rect 1232 1271 1236 1275
rect 1272 1271 1276 1275
rect 1344 1271 1348 1275
rect 1424 1271 1428 1275
rect 1504 1271 1508 1275
rect 1584 1271 1588 1275
rect 1664 1271 1668 1275
rect 1744 1271 1748 1275
rect 1824 1271 1828 1275
rect 1904 1271 1908 1275
rect 1912 1271 1916 1275
rect 1992 1271 1996 1275
rect 2080 1271 2084 1275
rect 820 1259 824 1263
rect 900 1259 904 1263
rect 936 1259 940 1263
rect 980 1259 984 1263
rect 1044 1259 1048 1263
rect 800 1251 804 1255
rect 1156 1249 1160 1253
rect 1196 1247 1200 1251
rect 1232 1247 1236 1251
rect 1244 1249 1248 1253
rect 1316 1247 1320 1251
rect 1396 1247 1400 1251
rect 1476 1247 1480 1251
rect 1556 1247 1560 1251
rect 1636 1247 1640 1251
rect 1716 1247 1720 1251
rect 1796 1247 1800 1251
rect 1876 1247 1880 1251
rect 1912 1247 1916 1251
rect 1964 1247 1968 1251
rect 2052 1247 2056 1251
rect 260 1243 264 1247
rect 308 1243 312 1247
rect 356 1243 360 1247
rect 392 1243 396 1247
rect 412 1243 416 1247
rect 476 1243 480 1247
rect 540 1243 544 1247
rect 604 1243 608 1247
rect 640 1243 644 1247
rect 668 1243 672 1247
rect 732 1243 736 1247
rect 796 1243 800 1247
rect 860 1243 864 1247
rect 924 1243 928 1247
rect 288 1219 292 1223
rect 336 1221 340 1225
rect 1156 1233 1160 1237
rect 1196 1231 1200 1235
rect 1236 1231 1240 1235
rect 1276 1231 1280 1235
rect 1312 1231 1316 1235
rect 1324 1233 1328 1237
rect 1372 1231 1376 1235
rect 1408 1231 1412 1235
rect 1420 1231 1424 1235
rect 1468 1233 1472 1237
rect 1532 1231 1536 1235
rect 1612 1231 1616 1235
rect 1648 1231 1652 1235
rect 1716 1231 1720 1235
rect 1836 1231 1840 1235
rect 1964 1231 1968 1235
rect 2068 1231 2072 1235
rect 384 1219 388 1223
rect 392 1219 396 1223
rect 440 1219 444 1223
rect 504 1219 508 1223
rect 568 1219 572 1223
rect 632 1219 636 1223
rect 640 1219 644 1223
rect 696 1219 700 1223
rect 760 1219 764 1223
rect 824 1219 828 1223
rect 888 1219 892 1223
rect 952 1219 956 1223
rect 1408 1211 1412 1215
rect 1648 1211 1652 1215
rect 1184 1207 1188 1211
rect 1224 1207 1228 1211
rect 1264 1207 1268 1211
rect 1304 1207 1308 1211
rect 1312 1207 1316 1211
rect 1352 1207 1356 1211
rect 1400 1207 1404 1211
rect 1448 1207 1452 1211
rect 1496 1207 1500 1211
rect 1560 1207 1564 1211
rect 1640 1207 1644 1211
rect 1664 1207 1668 1211
rect 1744 1207 1748 1211
rect 1864 1207 1868 1211
rect 1992 1207 1996 1211
rect 2096 1207 2100 1211
rect 1664 1187 1668 1191
rect 248 1175 252 1179
rect 304 1175 308 1179
rect 368 1175 372 1179
rect 432 1175 436 1179
rect 504 1175 508 1179
rect 576 1175 580 1179
rect 656 1175 660 1179
rect 736 1175 740 1179
rect 816 1175 820 1179
rect 896 1175 900 1179
rect 984 1175 988 1179
rect 1312 1163 1316 1167
rect 1352 1163 1356 1167
rect 1392 1163 1396 1167
rect 1400 1163 1404 1167
rect 1440 1163 1444 1167
rect 1496 1163 1500 1167
rect 1552 1163 1556 1167
rect 1608 1163 1612 1167
rect 1664 1163 1668 1167
rect 1728 1163 1732 1167
rect 1792 1163 1796 1167
rect 1864 1163 1868 1167
rect 1944 1163 1948 1167
rect 2032 1163 2036 1167
rect 2096 1163 2100 1167
rect 220 1151 224 1155
rect 276 1151 280 1155
rect 340 1151 344 1155
rect 404 1151 408 1155
rect 476 1151 480 1155
rect 548 1151 552 1155
rect 628 1151 632 1155
rect 708 1151 712 1155
rect 788 1151 792 1155
rect 868 1151 872 1155
rect 956 1151 960 1155
rect 156 1139 160 1143
rect 196 1139 200 1143
rect 244 1139 248 1143
rect 300 1139 304 1143
rect 344 1139 348 1143
rect 364 1139 368 1143
rect 436 1139 440 1143
rect 508 1139 512 1143
rect 588 1139 592 1143
rect 676 1139 680 1143
rect 772 1139 776 1143
rect 876 1139 880 1143
rect 988 1139 992 1143
rect 1284 1139 1288 1143
rect 1324 1139 1328 1143
rect 1364 1139 1368 1143
rect 1412 1139 1416 1143
rect 1468 1139 1472 1143
rect 1524 1139 1528 1143
rect 1580 1139 1584 1143
rect 1636 1139 1640 1143
rect 1700 1139 1704 1143
rect 1764 1139 1768 1143
rect 1836 1139 1840 1143
rect 1916 1139 1920 1143
rect 2004 1139 2008 1143
rect 2068 1139 2072 1143
rect 1400 1131 1404 1135
rect 1380 1119 1384 1123
rect 1420 1119 1424 1123
rect 1468 1119 1472 1123
rect 1524 1121 1528 1125
rect 1588 1119 1592 1123
rect 1652 1119 1656 1123
rect 1708 1121 1712 1125
rect 1764 1119 1768 1123
rect 1820 1119 1824 1123
rect 1868 1119 1872 1123
rect 1924 1119 1928 1123
rect 1980 1119 1984 1123
rect 2028 1119 2032 1123
rect 2068 1119 2072 1123
rect 184 1115 188 1119
rect 224 1115 228 1119
rect 272 1115 276 1119
rect 328 1115 332 1119
rect 344 1115 348 1119
rect 392 1115 396 1119
rect 464 1115 468 1119
rect 536 1115 540 1119
rect 616 1115 620 1119
rect 704 1115 708 1119
rect 800 1115 804 1119
rect 904 1115 908 1119
rect 1016 1115 1020 1119
rect 1408 1095 1412 1099
rect 1448 1095 1452 1099
rect 1496 1095 1500 1099
rect 1552 1095 1556 1099
rect 1616 1095 1620 1099
rect 1680 1095 1684 1099
rect 1736 1095 1740 1099
rect 1792 1095 1796 1099
rect 1848 1095 1852 1099
rect 1896 1095 1900 1099
rect 1952 1095 1956 1099
rect 2008 1095 2012 1099
rect 2056 1095 2060 1099
rect 2096 1095 2100 1099
rect 224 1063 228 1067
rect 232 1063 236 1067
rect 272 1063 276 1067
rect 280 1063 284 1067
rect 328 1063 332 1067
rect 392 1063 396 1067
rect 400 1063 404 1067
rect 456 1063 460 1067
rect 528 1063 532 1067
rect 600 1063 604 1067
rect 672 1063 676 1067
rect 744 1063 748 1067
rect 808 1063 812 1067
rect 864 1063 868 1067
rect 920 1063 924 1067
rect 976 1063 980 1067
rect 1032 1063 1036 1067
rect 1072 1063 1076 1067
rect 1184 1051 1188 1055
rect 1272 1051 1276 1055
rect 1384 1051 1388 1055
rect 1496 1051 1500 1055
rect 1600 1051 1604 1055
rect 1696 1051 1700 1055
rect 1784 1051 1788 1055
rect 1872 1051 1876 1055
rect 1880 1051 1884 1055
rect 1952 1051 1956 1055
rect 1960 1051 1964 1055
rect 2032 1051 2036 1055
rect 2096 1051 2100 1055
rect 196 1039 200 1043
rect 232 1039 236 1043
rect 244 1039 248 1043
rect 280 1039 284 1043
rect 300 1039 304 1043
rect 364 1039 368 1043
rect 400 1039 404 1043
rect 428 1039 432 1043
rect 500 1039 504 1043
rect 572 1039 576 1043
rect 644 1039 648 1043
rect 716 1039 720 1043
rect 780 1039 784 1043
rect 836 1039 840 1043
rect 892 1039 896 1043
rect 948 1039 952 1043
rect 1004 1039 1008 1043
rect 1044 1039 1048 1043
rect 1156 1027 1160 1031
rect 1244 1027 1248 1031
rect 1356 1027 1360 1031
rect 1468 1027 1472 1031
rect 1572 1027 1576 1031
rect 1668 1027 1672 1031
rect 1756 1027 1760 1031
rect 1844 1027 1848 1031
rect 1880 1027 1884 1031
rect 1924 1027 1928 1031
rect 1960 1027 1964 1031
rect 2004 1027 2008 1031
rect 2068 1027 2072 1031
rect 220 1023 224 1027
rect 268 1023 272 1027
rect 304 1023 308 1027
rect 332 1023 336 1027
rect 404 1023 408 1027
rect 476 1023 480 1027
rect 556 1023 560 1027
rect 628 1023 632 1027
rect 700 1023 704 1027
rect 772 1023 776 1027
rect 836 1023 840 1027
rect 900 1023 904 1027
rect 964 1023 968 1027
rect 1036 1023 1040 1027
rect 1156 1015 1160 1019
rect 1228 1015 1232 1019
rect 1300 1015 1304 1019
rect 1380 1015 1384 1019
rect 1460 1015 1464 1019
rect 1540 1015 1544 1019
rect 1620 1015 1624 1019
rect 1692 1015 1696 1019
rect 1756 1015 1760 1019
rect 1820 1015 1824 1019
rect 1884 1015 1888 1019
rect 1948 1015 1952 1019
rect 248 999 252 1003
rect 296 999 300 1003
rect 304 999 308 1003
rect 360 999 364 1003
rect 432 999 436 1003
rect 504 999 508 1003
rect 584 999 588 1003
rect 656 999 660 1003
rect 728 999 732 1003
rect 800 999 804 1003
rect 864 999 868 1003
rect 928 999 932 1003
rect 992 999 996 1003
rect 1064 999 1068 1003
rect 1184 991 1188 995
rect 1256 991 1260 995
rect 1328 991 1332 995
rect 1408 991 1412 995
rect 1488 991 1492 995
rect 1568 991 1572 995
rect 1648 991 1652 995
rect 1720 991 1724 995
rect 1784 991 1788 995
rect 1848 991 1852 995
rect 1912 991 1916 995
rect 1976 991 1980 995
rect 176 951 180 955
rect 240 951 244 955
rect 312 951 316 955
rect 392 951 396 955
rect 472 951 476 955
rect 552 951 556 955
rect 624 951 628 955
rect 696 951 700 955
rect 760 951 764 955
rect 824 951 828 955
rect 888 951 892 955
rect 952 951 956 955
rect 1016 951 1020 955
rect 1072 951 1076 955
rect 1264 947 1268 951
rect 1328 947 1332 951
rect 1400 947 1404 951
rect 1464 947 1468 951
rect 1536 947 1540 951
rect 1608 947 1612 951
rect 1680 947 1684 951
rect 1752 947 1756 951
rect 1824 947 1828 951
rect 1896 947 1900 951
rect 1968 947 1972 951
rect 2040 947 2044 951
rect 2048 947 2052 951
rect 2096 947 2100 951
rect 148 927 152 931
rect 212 927 216 931
rect 284 927 288 931
rect 364 927 368 931
rect 444 927 448 931
rect 524 927 528 931
rect 596 927 600 931
rect 668 927 672 931
rect 732 927 736 931
rect 796 927 800 931
rect 860 927 864 931
rect 924 927 928 931
rect 988 927 992 931
rect 1044 927 1048 931
rect 1236 923 1240 927
rect 1300 923 1304 927
rect 1372 923 1376 927
rect 1436 923 1440 927
rect 1508 923 1512 927
rect 1580 923 1584 927
rect 1652 923 1656 927
rect 1724 923 1728 927
rect 1796 923 1800 927
rect 1868 923 1872 927
rect 1940 923 1944 927
rect 2012 923 2016 927
rect 2048 923 2052 927
rect 2068 923 2072 927
rect 132 915 136 919
rect 180 915 184 919
rect 252 915 256 919
rect 324 915 328 919
rect 396 915 400 919
rect 448 915 452 919
rect 460 915 464 919
rect 524 915 528 919
rect 596 915 600 919
rect 668 915 672 919
rect 740 915 744 919
rect 812 915 816 919
rect 892 915 896 919
rect 980 915 984 919
rect 1044 915 1048 919
rect 1284 907 1288 911
rect 1324 907 1328 911
rect 1372 907 1376 911
rect 1420 907 1424 911
rect 1476 907 1480 911
rect 1548 907 1552 911
rect 1620 907 1624 911
rect 1700 907 1704 911
rect 1788 907 1792 911
rect 1876 907 1880 911
rect 1964 907 1968 911
rect 2060 907 2064 911
rect 160 891 164 895
rect 208 891 212 895
rect 280 891 284 895
rect 352 891 356 895
rect 424 891 428 895
rect 448 891 452 895
rect 488 891 492 895
rect 552 891 556 895
rect 624 891 628 895
rect 696 891 700 895
rect 768 891 772 895
rect 840 891 844 895
rect 920 891 924 895
rect 1008 891 1012 895
rect 1072 891 1076 895
rect 1312 883 1316 887
rect 1352 883 1356 887
rect 1400 883 1404 887
rect 1448 883 1452 887
rect 1504 883 1508 887
rect 1576 883 1580 887
rect 1648 883 1652 887
rect 1728 883 1732 887
rect 1816 883 1820 887
rect 1904 883 1908 887
rect 1992 883 1996 887
rect 2088 883 2092 887
rect 160 843 164 847
rect 200 843 204 847
rect 240 843 244 847
rect 304 843 308 847
rect 368 843 372 847
rect 384 843 388 847
rect 424 843 428 847
rect 488 843 492 847
rect 560 843 564 847
rect 640 843 644 847
rect 736 843 740 847
rect 808 843 812 847
rect 848 843 852 847
rect 968 843 972 847
rect 1072 843 1076 847
rect 1184 839 1188 843
rect 1224 839 1228 843
rect 1288 839 1292 843
rect 1352 839 1356 843
rect 1424 839 1428 843
rect 1496 839 1500 843
rect 1568 839 1572 843
rect 1648 839 1652 843
rect 1728 839 1732 843
rect 1800 839 1804 843
rect 1880 839 1884 843
rect 1960 839 1964 843
rect 2040 839 2044 843
rect 2096 839 2100 843
rect 132 819 136 823
rect 172 819 176 823
rect 212 819 216 823
rect 276 819 280 823
rect 340 819 344 823
rect 384 819 388 823
rect 396 819 400 823
rect 460 819 464 823
rect 532 819 536 823
rect 612 819 616 823
rect 708 819 712 823
rect 808 819 812 823
rect 820 819 824 823
rect 940 819 944 823
rect 1044 819 1048 823
rect 1156 817 1160 821
rect 1196 815 1200 819
rect 1260 815 1264 819
rect 1324 815 1328 819
rect 1396 815 1400 819
rect 1468 815 1472 819
rect 1540 815 1544 819
rect 1620 815 1624 819
rect 1700 815 1704 819
rect 1772 815 1776 819
rect 1852 815 1856 819
rect 1932 815 1936 819
rect 2012 815 2016 819
rect 2068 815 2072 819
rect 132 807 136 811
rect 172 807 176 811
rect 212 807 216 811
rect 276 807 280 811
rect 332 807 336 811
rect 388 807 392 811
rect 452 807 456 811
rect 516 807 520 811
rect 580 807 584 811
rect 616 807 620 811
rect 652 807 656 811
rect 732 807 736 811
rect 812 807 816 811
rect 892 807 896 811
rect 980 807 984 811
rect 1044 807 1048 811
rect 200 791 204 795
rect 160 783 164 787
rect 200 783 204 787
rect 216 783 220 787
rect 240 783 244 787
rect 248 783 252 787
rect 304 783 308 787
rect 360 783 364 787
rect 416 783 420 787
rect 480 783 484 787
rect 544 783 548 787
rect 608 783 612 787
rect 160 739 164 743
rect 232 739 236 743
rect 1156 795 1160 799
rect 1236 795 1240 799
rect 1340 795 1344 799
rect 1444 795 1448 799
rect 1536 795 1540 799
rect 1548 795 1552 799
rect 1652 795 1656 799
rect 1748 795 1752 799
rect 1836 795 1840 799
rect 1916 795 1920 799
rect 2004 795 2008 799
rect 2068 795 2072 799
rect 680 783 684 787
rect 760 783 764 787
rect 840 783 844 787
rect 920 783 924 787
rect 1008 783 1012 787
rect 1072 783 1076 787
rect 1184 771 1188 775
rect 1264 771 1268 775
rect 1368 771 1372 775
rect 1472 771 1476 775
rect 1536 771 1540 775
rect 1576 771 1580 775
rect 1680 771 1684 775
rect 1776 771 1780 775
rect 1864 771 1868 775
rect 1944 771 1948 775
rect 2032 771 2036 775
rect 2096 771 2100 775
rect 320 739 324 743
rect 400 739 404 743
rect 472 739 476 743
rect 480 739 484 743
rect 544 739 548 743
rect 608 739 612 743
rect 616 739 620 743
rect 664 739 668 743
rect 712 739 716 743
rect 768 739 772 743
rect 824 739 828 743
rect 880 739 884 743
rect 1184 727 1188 731
rect 1224 727 1228 731
rect 1264 727 1268 731
rect 1312 727 1316 731
rect 1384 727 1388 731
rect 1464 727 1468 731
rect 1552 727 1556 731
rect 1640 727 1644 731
rect 1736 727 1740 731
rect 1832 727 1836 731
rect 1840 727 1844 731
rect 1928 727 1932 731
rect 1936 727 1940 731
rect 2024 727 2028 731
rect 2096 727 2100 731
rect 132 715 136 719
rect 204 715 208 719
rect 248 715 252 719
rect 292 715 296 719
rect 372 715 376 719
rect 444 715 448 719
rect 480 715 484 719
rect 516 715 520 719
rect 580 715 584 719
rect 636 715 640 719
rect 684 715 688 719
rect 740 715 744 719
rect 796 715 800 719
rect 852 715 856 719
rect 1156 703 1160 707
rect 1196 703 1200 707
rect 1236 703 1240 707
rect 1284 703 1288 707
rect 1356 703 1360 707
rect 1436 703 1440 707
rect 1524 703 1528 707
rect 1612 703 1616 707
rect 1708 703 1712 707
rect 1804 703 1808 707
rect 1840 703 1844 707
rect 1900 703 1904 707
rect 1936 703 1940 707
rect 1996 703 2000 707
rect 2068 703 2072 707
rect 132 699 136 703
rect 180 699 184 703
rect 244 699 248 703
rect 308 699 312 703
rect 380 699 384 703
rect 452 699 456 703
rect 516 699 520 703
rect 580 699 584 703
rect 644 699 648 703
rect 708 699 712 703
rect 744 699 748 703
rect 764 699 768 703
rect 820 699 824 703
rect 856 699 860 703
rect 876 699 880 703
rect 940 699 944 703
rect 1236 687 1240 691
rect 1284 687 1288 691
rect 1332 687 1336 691
rect 1388 689 1392 693
rect 1424 687 1428 691
rect 1444 687 1448 691
rect 1508 687 1512 691
rect 1572 687 1576 691
rect 1636 689 1640 693
rect 1700 687 1704 691
rect 1764 687 1768 691
rect 1808 687 1812 691
rect 1828 687 1832 691
rect 1892 687 1896 691
rect 1956 687 1960 691
rect 2020 687 2024 691
rect 2068 687 2072 691
rect 160 675 164 679
rect 208 675 212 679
rect 272 675 276 679
rect 336 675 340 679
rect 408 675 412 679
rect 480 675 484 679
rect 544 675 548 679
rect 608 675 612 679
rect 672 675 676 679
rect 736 675 740 679
rect 744 675 748 679
rect 792 675 796 679
rect 848 675 852 679
rect 856 675 860 679
rect 904 675 908 679
rect 968 675 972 679
rect 1264 663 1268 667
rect 1312 663 1316 667
rect 1360 663 1364 667
rect 1416 663 1420 667
rect 1424 663 1428 667
rect 1472 663 1476 667
rect 1536 663 1540 667
rect 1600 663 1604 667
rect 1664 663 1668 667
rect 1728 663 1732 667
rect 1792 663 1796 667
rect 1808 663 1812 667
rect 1856 663 1860 667
rect 1920 663 1924 667
rect 1984 663 1988 667
rect 2048 663 2052 667
rect 2096 663 2100 667
rect 184 623 188 627
rect 240 623 244 627
rect 312 623 316 627
rect 392 623 396 627
rect 480 623 484 627
rect 488 623 492 627
rect 568 623 572 627
rect 656 623 660 627
rect 744 623 748 627
rect 824 623 828 627
rect 896 623 900 627
rect 976 623 980 627
rect 1056 623 1060 627
rect 1304 619 1308 623
rect 1344 619 1348 623
rect 1392 619 1396 623
rect 1448 619 1452 623
rect 1504 619 1508 623
rect 1560 619 1564 623
rect 1616 619 1620 623
rect 1672 619 1676 623
rect 1744 619 1748 623
rect 1824 619 1828 623
rect 1904 619 1908 623
rect 1992 619 1996 623
rect 2088 619 2092 623
rect 156 599 160 603
rect 212 599 216 603
rect 284 599 288 603
rect 364 599 368 603
rect 452 599 456 603
rect 488 599 492 603
rect 540 599 544 603
rect 628 599 632 603
rect 716 599 720 603
rect 796 599 800 603
rect 868 599 872 603
rect 948 599 952 603
rect 1028 599 1032 603
rect 1276 595 1280 599
rect 1316 595 1320 599
rect 1364 595 1368 599
rect 1420 595 1424 599
rect 1476 595 1480 599
rect 1532 595 1536 599
rect 1588 595 1592 599
rect 1644 595 1648 599
rect 1716 595 1720 599
rect 1796 595 1800 599
rect 1876 595 1880 599
rect 1964 595 1968 599
rect 2060 595 2064 599
rect 156 585 160 589
rect 204 583 208 587
rect 252 583 256 587
rect 308 583 312 587
rect 380 583 384 587
rect 460 583 464 587
rect 540 583 544 587
rect 620 583 624 587
rect 700 583 704 587
rect 780 585 784 589
rect 852 583 856 587
rect 924 583 928 587
rect 996 583 1000 587
rect 1032 583 1036 587
rect 1044 583 1048 587
rect 1332 583 1336 587
rect 1372 583 1376 587
rect 1412 583 1416 587
rect 1460 583 1464 587
rect 1516 583 1520 587
rect 1580 583 1584 587
rect 1652 583 1656 587
rect 1724 583 1728 587
rect 1804 583 1808 587
rect 1884 583 1888 587
rect 1972 583 1976 587
rect 2060 583 2064 587
rect 184 559 188 563
rect 232 559 236 563
rect 280 559 284 563
rect 336 559 340 563
rect 408 559 412 563
rect 488 559 492 563
rect 568 559 572 563
rect 648 559 652 563
rect 728 559 732 563
rect 808 559 812 563
rect 880 559 884 563
rect 952 559 956 563
rect 1024 559 1028 563
rect 1032 559 1036 563
rect 1072 559 1076 563
rect 1360 559 1364 563
rect 1400 559 1404 563
rect 1440 559 1444 563
rect 1488 559 1492 563
rect 1544 559 1548 563
rect 1608 559 1612 563
rect 1680 559 1684 563
rect 1752 559 1756 563
rect 1832 559 1836 563
rect 1912 559 1916 563
rect 2000 559 2004 563
rect 2088 559 2092 563
rect 1216 511 1220 515
rect 1264 511 1268 515
rect 1312 511 1316 515
rect 1368 511 1372 515
rect 1376 511 1380 515
rect 1432 511 1436 515
rect 1504 511 1508 515
rect 1568 511 1572 515
rect 1632 511 1636 515
rect 1696 511 1700 515
rect 1760 511 1764 515
rect 1824 511 1828 515
rect 1888 512 1892 516
rect 1960 511 1964 515
rect 2032 511 2036 515
rect 2096 511 2100 515
rect 192 507 196 511
rect 200 507 204 511
rect 248 507 252 511
rect 312 507 316 511
rect 384 507 388 511
rect 456 507 460 511
rect 464 507 468 511
rect 536 507 540 511
rect 616 507 620 511
rect 688 507 692 511
rect 760 507 764 511
rect 792 507 796 511
rect 832 507 836 511
rect 896 507 900 511
rect 960 507 964 511
rect 1024 507 1028 511
rect 1072 507 1076 511
rect 164 483 168 487
rect 200 483 204 487
rect 220 485 224 489
rect 1188 487 1192 491
rect 1236 487 1240 491
rect 1284 487 1288 491
rect 1340 487 1344 491
rect 1376 487 1380 491
rect 1404 487 1408 491
rect 1476 487 1480 491
rect 1540 487 1544 491
rect 1604 487 1608 491
rect 1668 487 1672 491
rect 1732 487 1736 491
rect 1796 487 1800 491
rect 1860 487 1864 491
rect 1932 487 1936 491
rect 2004 487 2008 491
rect 2068 487 2072 491
rect 284 483 288 487
rect 356 483 360 487
rect 428 483 432 487
rect 464 483 468 487
rect 508 483 512 487
rect 588 483 592 487
rect 660 483 664 487
rect 732 483 736 487
rect 784 483 788 487
rect 792 483 796 487
rect 804 483 808 487
rect 868 483 872 487
rect 932 483 936 487
rect 996 483 1000 487
rect 1044 483 1048 487
rect 164 471 168 475
rect 228 471 232 475
rect 272 471 276 475
rect 300 471 304 475
rect 372 471 376 475
rect 452 471 456 475
rect 532 471 536 475
rect 604 471 608 475
rect 676 471 680 475
rect 740 471 744 475
rect 1156 475 1160 479
rect 1260 475 1264 479
rect 1380 475 1384 479
rect 1492 475 1496 479
rect 1596 475 1600 479
rect 1700 475 1704 479
rect 1796 475 1800 479
rect 1884 475 1888 479
rect 1980 475 1984 479
rect 2068 475 2072 479
rect 796 471 800 475
rect 852 471 856 475
rect 900 471 904 475
rect 956 471 960 475
rect 1004 471 1008 475
rect 1044 471 1048 475
rect 784 451 788 455
rect 1184 451 1188 455
rect 1288 451 1292 455
rect 1408 451 1412 455
rect 1520 451 1524 455
rect 1624 451 1628 455
rect 1728 451 1732 455
rect 1824 451 1828 455
rect 1912 451 1916 455
rect 2008 451 2012 455
rect 2096 451 2100 455
rect 192 447 196 451
rect 256 447 260 451
rect 272 447 276 451
rect 328 447 332 451
rect 400 447 404 451
rect 480 447 484 451
rect 560 447 564 451
rect 632 447 636 451
rect 704 447 708 451
rect 768 447 772 451
rect 824 447 828 451
rect 880 447 884 451
rect 928 447 932 451
rect 984 447 988 451
rect 1032 447 1036 451
rect 1072 447 1076 451
rect 1184 407 1188 411
rect 1224 407 1228 411
rect 1280 407 1284 411
rect 1360 407 1364 411
rect 1440 407 1444 411
rect 1528 407 1532 411
rect 1616 407 1620 411
rect 1696 407 1700 411
rect 1776 407 1780 411
rect 1848 407 1852 411
rect 1856 407 1860 411
rect 1912 407 1916 411
rect 1976 407 1980 411
rect 2048 407 2052 411
rect 2096 407 2100 411
rect 176 403 180 407
rect 240 403 244 407
rect 264 403 268 407
rect 304 403 308 407
rect 376 403 380 407
rect 400 403 404 407
rect 448 403 452 407
rect 456 403 460 407
rect 512 403 516 407
rect 576 403 580 407
rect 640 403 644 407
rect 696 403 700 407
rect 752 403 756 407
rect 816 403 820 407
rect 880 403 884 407
rect 1156 383 1160 387
rect 1196 383 1200 387
rect 1252 383 1256 387
rect 1332 383 1336 387
rect 1412 383 1416 387
rect 1500 383 1504 387
rect 1588 383 1592 387
rect 1668 383 1672 387
rect 1748 383 1752 387
rect 1820 383 1824 387
rect 1856 383 1860 387
rect 1884 383 1888 387
rect 1948 383 1952 387
rect 2020 383 2024 387
rect 2068 383 2072 387
rect 148 379 152 383
rect 212 379 216 383
rect 256 379 260 383
rect 264 379 268 383
rect 276 379 280 383
rect 348 379 352 383
rect 400 379 404 383
rect 420 379 424 383
rect 456 379 460 383
rect 484 379 488 383
rect 548 379 552 383
rect 612 379 616 383
rect 668 379 672 383
rect 724 379 728 383
rect 788 379 792 383
rect 852 379 856 383
rect 132 367 136 371
rect 172 367 176 371
rect 212 367 216 371
rect 160 343 164 347
rect 200 343 204 347
rect 240 343 244 347
rect 268 367 272 371
rect 332 367 336 371
rect 396 367 400 371
rect 460 367 464 371
rect 516 367 520 371
rect 572 367 576 371
rect 616 367 620 371
rect 628 367 632 371
rect 684 367 688 371
rect 748 367 752 371
rect 1300 369 1304 373
rect 1340 367 1344 371
rect 1380 367 1384 371
rect 1420 367 1424 371
rect 1460 367 1464 371
rect 1500 367 1504 371
rect 1548 367 1552 371
rect 1612 367 1616 371
rect 1676 367 1680 371
rect 1748 367 1752 371
rect 1828 367 1832 371
rect 1916 367 1920 371
rect 1952 367 1956 371
rect 2004 367 2008 371
rect 2068 367 2072 371
rect 616 347 620 351
rect 296 343 300 347
rect 360 343 364 347
rect 424 343 428 347
rect 488 343 492 347
rect 544 343 548 347
rect 600 343 604 347
rect 656 343 660 347
rect 712 343 716 347
rect 776 343 780 347
rect 1328 343 1332 347
rect 1368 343 1372 347
rect 1408 343 1412 347
rect 1448 343 1452 347
rect 1488 343 1492 347
rect 1528 343 1532 347
rect 1576 343 1580 347
rect 1640 343 1644 347
rect 1704 343 1708 347
rect 1776 343 1780 347
rect 1856 343 1860 347
rect 1944 343 1948 347
rect 1952 343 1956 347
rect 2032 343 2036 347
rect 2096 343 2100 347
rect 256 319 260 323
rect 160 295 164 299
rect 192 295 196 299
rect 232 295 236 299
rect 320 295 324 299
rect 408 295 412 299
rect 496 295 500 299
rect 504 295 508 299
rect 576 295 580 299
rect 648 295 652 299
rect 656 295 660 299
rect 712 295 716 299
rect 776 295 780 299
rect 784 295 788 299
rect 832 295 836 299
rect 840 295 844 299
rect 896 295 900 299
rect 960 295 964 299
rect 1192 295 1196 299
rect 1232 295 1236 299
rect 1272 295 1276 299
rect 1280 295 1284 299
rect 1320 295 1324 299
rect 1368 295 1372 299
rect 1416 295 1420 299
rect 1464 295 1468 299
rect 1520 295 1524 299
rect 1584 295 1588 299
rect 1648 295 1652 299
rect 1656 295 1660 299
rect 1720 295 1724 299
rect 1800 295 1804 299
rect 1880 295 1884 299
rect 1960 295 1964 299
rect 2040 295 2044 299
rect 2048 295 2052 299
rect 2096 295 2100 299
rect 132 271 136 275
rect 192 271 196 275
rect 204 271 208 275
rect 292 271 296 275
rect 380 271 384 275
rect 468 271 472 275
rect 504 271 508 275
rect 548 271 552 275
rect 620 271 624 275
rect 656 271 660 275
rect 684 271 688 275
rect 748 271 752 275
rect 784 271 788 275
rect 804 271 808 275
rect 840 271 844 275
rect 868 273 872 277
rect 932 271 936 275
rect 1164 273 1168 277
rect 1204 273 1208 277
rect 1244 271 1248 275
rect 1280 271 1284 275
rect 1292 271 1296 275
rect 1340 271 1344 275
rect 1388 271 1392 275
rect 1436 271 1440 275
rect 1492 271 1496 275
rect 1556 271 1560 275
rect 1620 271 1624 275
rect 1692 271 1696 275
rect 1772 271 1776 275
rect 1852 271 1856 275
rect 1932 271 1936 275
rect 2012 271 2016 275
rect 2048 271 2052 275
rect 2068 271 2072 275
rect 132 259 136 263
rect 196 259 200 263
rect 276 259 280 263
rect 356 259 360 263
rect 436 259 440 263
rect 472 259 476 263
rect 508 259 512 263
rect 580 259 584 263
rect 644 259 648 263
rect 680 259 684 263
rect 700 259 704 263
rect 756 259 760 263
rect 812 259 816 263
rect 876 259 880 263
rect 1656 259 1660 263
rect 1156 251 1160 255
rect 1204 251 1208 255
rect 1268 251 1272 255
rect 1324 251 1328 255
rect 1388 251 1392 255
rect 1452 251 1456 255
rect 1524 251 1528 255
rect 1604 253 1608 257
rect 1684 251 1688 255
rect 1764 251 1768 255
rect 1836 251 1840 255
rect 1916 251 1920 255
rect 1996 251 2000 255
rect 2068 251 2072 255
rect 160 235 164 239
rect 224 235 228 239
rect 304 235 308 239
rect 384 235 388 239
rect 464 235 468 239
rect 472 235 476 239
rect 536 235 540 239
rect 608 235 612 239
rect 672 235 676 239
rect 680 235 684 239
rect 728 235 732 239
rect 784 235 788 239
rect 840 235 844 239
rect 904 235 908 239
rect 1184 227 1188 231
rect 1232 227 1236 231
rect 1296 227 1300 231
rect 1352 227 1356 231
rect 1416 227 1420 231
rect 1480 227 1484 231
rect 1552 227 1556 231
rect 1632 227 1636 231
rect 1712 227 1716 231
rect 1792 227 1796 231
rect 1864 227 1868 231
rect 1944 227 1948 231
rect 2024 227 2028 231
rect 2096 227 2100 231
rect 160 187 164 191
rect 208 187 212 191
rect 256 187 260 191
rect 304 187 308 191
rect 352 187 356 191
rect 360 187 364 191
rect 400 187 404 191
rect 440 187 444 191
rect 480 187 484 191
rect 528 187 532 191
rect 576 187 580 191
rect 624 187 628 191
rect 672 187 676 191
rect 720 187 724 191
rect 768 187 772 191
rect 1184 183 1188 187
rect 1224 183 1228 187
rect 1232 183 1236 187
rect 1288 183 1292 187
rect 1352 183 1356 187
rect 1424 183 1428 187
rect 1496 183 1500 187
rect 1568 183 1572 187
rect 1632 183 1636 187
rect 1640 183 1644 187
rect 1696 183 1700 187
rect 1704 183 1708 187
rect 1760 183 1764 187
rect 1832 183 1836 187
rect 1904 183 1908 187
rect 1976 183 1980 187
rect 2048 183 2052 187
rect 2096 183 2100 187
rect 132 163 136 167
rect 180 163 184 167
rect 228 163 232 167
rect 276 163 280 167
rect 324 163 328 167
rect 360 163 364 167
rect 372 165 376 169
rect 412 163 416 167
rect 452 163 456 167
rect 500 163 504 167
rect 548 163 552 167
rect 596 163 600 167
rect 644 163 648 167
rect 692 163 696 167
rect 740 163 744 167
rect 1156 161 1160 165
rect 1196 159 1200 163
rect 1232 159 1236 163
rect 1260 159 1264 163
rect 1324 159 1328 163
rect 1396 159 1400 163
rect 1468 159 1472 163
rect 1540 159 1544 163
rect 1604 159 1608 163
rect 1640 159 1644 163
rect 1668 159 1672 163
rect 1704 159 1708 163
rect 1732 159 1736 163
rect 1804 159 1808 163
rect 1876 159 1880 163
rect 1948 159 1952 163
rect 2020 159 2024 163
rect 2068 159 2072 163
rect 140 129 144 133
rect 180 127 184 131
rect 220 127 224 131
rect 260 127 264 131
rect 300 127 304 131
rect 340 127 344 131
rect 380 127 384 131
rect 420 127 424 131
rect 460 127 464 131
rect 500 127 504 131
rect 540 127 544 131
rect 580 127 584 131
rect 620 127 624 131
rect 660 127 664 131
rect 700 127 704 131
rect 740 127 744 131
rect 780 127 784 131
rect 828 127 832 131
rect 876 127 880 131
rect 912 127 916 131
rect 924 127 928 131
rect 964 127 968 131
rect 1004 127 1008 131
rect 1044 127 1048 131
rect 1156 127 1160 131
rect 1204 129 1208 133
rect 1268 127 1272 131
rect 1332 127 1336 131
rect 1396 127 1400 131
rect 1452 127 1456 131
rect 1508 129 1512 133
rect 1556 127 1560 131
rect 1604 127 1608 131
rect 1644 127 1648 131
rect 1684 127 1688 131
rect 1724 127 1728 131
rect 1764 127 1768 131
rect 1804 127 1808 131
rect 1852 127 1856 131
rect 1888 127 1892 131
rect 1900 127 1904 131
rect 1948 127 1952 131
rect 1988 127 1992 131
rect 2028 127 2032 131
rect 2068 127 2072 131
rect 168 103 172 107
rect 208 103 212 107
rect 248 103 252 107
rect 288 103 292 107
rect 328 103 332 107
rect 368 103 372 107
rect 408 103 412 107
rect 448 103 452 107
rect 488 103 492 107
rect 528 103 532 107
rect 568 103 572 107
rect 608 103 612 107
rect 648 103 652 107
rect 688 103 692 107
rect 728 103 732 107
rect 768 103 772 107
rect 808 103 812 107
rect 856 103 860 107
rect 904 103 908 107
rect 912 103 916 107
rect 952 103 956 107
rect 992 103 996 107
rect 1032 103 1036 107
rect 1072 103 1076 107
rect 1184 103 1188 107
rect 1232 103 1236 107
rect 1296 103 1300 107
rect 1360 103 1364 107
rect 1424 103 1428 107
rect 1480 103 1484 107
rect 1536 103 1540 107
rect 1584 103 1588 107
rect 1632 103 1636 107
rect 1672 103 1676 107
rect 1712 103 1716 107
rect 1752 103 1756 107
rect 1792 103 1796 107
rect 1832 103 1836 107
rect 1880 103 1884 107
rect 1888 103 1892 107
rect 1928 103 1932 107
rect 1976 103 1980 107
rect 2056 103 2060 107
rect 2096 103 2100 107
<< m2 >>
rect 1678 2223 1689 2224
rect 1678 2219 1679 2223
rect 1683 2219 1684 2223
rect 1688 2219 1689 2223
rect 1678 2218 1689 2219
rect 1714 2223 1720 2224
rect 1714 2219 1715 2223
rect 1719 2222 1720 2223
rect 1723 2223 1729 2224
rect 1723 2222 1724 2223
rect 1719 2220 1724 2222
rect 1719 2219 1720 2220
rect 1714 2218 1720 2219
rect 1723 2219 1724 2220
rect 1728 2219 1729 2223
rect 1723 2218 1729 2219
rect 1750 2223 1756 2224
rect 1750 2219 1751 2223
rect 1755 2222 1756 2223
rect 1763 2223 1769 2224
rect 1763 2222 1764 2223
rect 1755 2220 1764 2222
rect 1755 2219 1756 2220
rect 1750 2218 1756 2219
rect 1763 2219 1764 2220
rect 1768 2219 1769 2223
rect 1763 2218 1769 2219
rect 1794 2223 1800 2224
rect 1794 2219 1795 2223
rect 1799 2222 1800 2223
rect 1803 2223 1809 2224
rect 1803 2222 1804 2223
rect 1799 2220 1804 2222
rect 1799 2219 1800 2220
rect 1794 2218 1800 2219
rect 1803 2219 1804 2220
rect 1808 2219 1809 2223
rect 1803 2218 1809 2219
rect 1686 2212 1692 2213
rect 134 2208 140 2209
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 134 2204 135 2208
rect 139 2204 140 2208
rect 134 2203 140 2204
rect 174 2208 180 2209
rect 174 2204 175 2208
rect 179 2204 180 2208
rect 174 2203 180 2204
rect 214 2208 220 2209
rect 214 2204 215 2208
rect 219 2204 220 2208
rect 214 2203 220 2204
rect 254 2208 260 2209
rect 254 2204 255 2208
rect 259 2204 260 2208
rect 254 2203 260 2204
rect 318 2208 324 2209
rect 318 2204 319 2208
rect 323 2204 324 2208
rect 318 2203 324 2204
rect 382 2208 388 2209
rect 382 2204 383 2208
rect 387 2204 388 2208
rect 382 2203 388 2204
rect 446 2208 452 2209
rect 446 2204 447 2208
rect 451 2204 452 2208
rect 446 2203 452 2204
rect 510 2208 516 2209
rect 510 2204 511 2208
rect 515 2204 516 2208
rect 510 2203 516 2204
rect 574 2208 580 2209
rect 574 2204 575 2208
rect 579 2204 580 2208
rect 574 2203 580 2204
rect 630 2208 636 2209
rect 630 2204 631 2208
rect 635 2204 636 2208
rect 630 2203 636 2204
rect 686 2208 692 2209
rect 686 2204 687 2208
rect 691 2204 692 2208
rect 686 2203 692 2204
rect 734 2208 740 2209
rect 734 2204 735 2208
rect 739 2204 740 2208
rect 734 2203 740 2204
rect 790 2208 796 2209
rect 790 2204 791 2208
rect 795 2204 796 2208
rect 790 2203 796 2204
rect 846 2208 852 2209
rect 846 2204 847 2208
rect 851 2204 852 2208
rect 846 2203 852 2204
rect 902 2208 908 2209
rect 902 2204 903 2208
rect 907 2204 908 2208
rect 1686 2208 1687 2212
rect 1691 2208 1692 2212
rect 1686 2207 1692 2208
rect 1726 2212 1732 2213
rect 1726 2208 1727 2212
rect 1731 2208 1732 2212
rect 1726 2207 1732 2208
rect 1766 2212 1772 2213
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1766 2207 1772 2208
rect 1806 2212 1812 2213
rect 1806 2208 1807 2212
rect 1811 2208 1812 2212
rect 1806 2207 1812 2208
rect 902 2203 908 2204
rect 1094 2205 1100 2206
rect 110 2200 116 2201
rect 1094 2201 1095 2205
rect 1099 2201 1100 2205
rect 1094 2200 1100 2201
rect 1134 2204 1140 2205
rect 1134 2200 1135 2204
rect 1139 2200 1140 2204
rect 2118 2204 2124 2205
rect 2118 2200 2119 2204
rect 2123 2200 2124 2204
rect 1134 2199 1140 2200
rect 1711 2199 1720 2200
rect 1711 2195 1712 2199
rect 1719 2195 1720 2199
rect 1711 2194 1720 2195
rect 1750 2199 1757 2200
rect 1750 2195 1751 2199
rect 1756 2195 1757 2199
rect 1750 2194 1757 2195
rect 1791 2199 1800 2200
rect 1791 2195 1792 2199
rect 1799 2195 1800 2199
rect 1791 2194 1800 2195
rect 1814 2199 1820 2200
rect 1814 2195 1815 2199
rect 1819 2198 1820 2199
rect 1831 2199 1837 2200
rect 2118 2199 2124 2200
rect 1831 2198 1832 2199
rect 1819 2196 1832 2198
rect 1819 2195 1820 2196
rect 1814 2194 1820 2195
rect 1831 2195 1832 2196
rect 1836 2195 1837 2199
rect 1831 2194 1837 2195
rect 159 2191 168 2192
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 159 2187 160 2191
rect 167 2187 168 2191
rect 159 2186 168 2187
rect 199 2191 208 2192
rect 199 2187 200 2191
rect 207 2187 208 2191
rect 199 2186 208 2187
rect 239 2191 248 2192
rect 239 2187 240 2191
rect 247 2187 248 2191
rect 239 2186 248 2187
rect 279 2191 285 2192
rect 279 2187 280 2191
rect 284 2190 285 2191
rect 310 2191 316 2192
rect 310 2190 311 2191
rect 284 2188 311 2190
rect 284 2187 285 2188
rect 279 2186 285 2187
rect 310 2187 311 2188
rect 315 2187 316 2191
rect 310 2186 316 2187
rect 343 2191 349 2192
rect 343 2187 344 2191
rect 348 2190 349 2191
rect 374 2191 380 2192
rect 374 2190 375 2191
rect 348 2188 375 2190
rect 348 2187 349 2188
rect 343 2186 349 2187
rect 374 2187 375 2188
rect 379 2187 380 2191
rect 374 2186 380 2187
rect 407 2191 413 2192
rect 407 2187 408 2191
rect 412 2190 413 2191
rect 438 2191 444 2192
rect 438 2190 439 2191
rect 412 2188 439 2190
rect 412 2187 413 2188
rect 407 2186 413 2187
rect 438 2187 439 2188
rect 443 2187 444 2191
rect 438 2186 444 2187
rect 454 2191 460 2192
rect 454 2187 455 2191
rect 459 2190 460 2191
rect 471 2191 477 2192
rect 471 2190 472 2191
rect 459 2188 472 2190
rect 459 2187 460 2188
rect 454 2186 460 2187
rect 471 2187 472 2188
rect 476 2187 477 2191
rect 471 2186 477 2187
rect 535 2191 541 2192
rect 535 2187 536 2191
rect 540 2190 541 2191
rect 566 2191 572 2192
rect 566 2190 567 2191
rect 540 2188 567 2190
rect 540 2187 541 2188
rect 535 2186 541 2187
rect 566 2187 567 2188
rect 571 2187 572 2191
rect 566 2186 572 2187
rect 599 2191 605 2192
rect 599 2187 600 2191
rect 604 2190 605 2191
rect 622 2191 628 2192
rect 622 2190 623 2191
rect 604 2188 623 2190
rect 604 2187 605 2188
rect 599 2186 605 2187
rect 622 2187 623 2188
rect 627 2187 628 2191
rect 622 2186 628 2187
rect 655 2191 661 2192
rect 655 2187 656 2191
rect 660 2190 661 2191
rect 678 2191 684 2192
rect 678 2190 679 2191
rect 660 2188 679 2190
rect 660 2187 661 2188
rect 655 2186 661 2187
rect 678 2187 679 2188
rect 683 2187 684 2191
rect 678 2186 684 2187
rect 711 2191 717 2192
rect 711 2187 712 2191
rect 716 2190 717 2191
rect 726 2191 732 2192
rect 726 2190 727 2191
rect 716 2188 727 2190
rect 716 2187 717 2188
rect 711 2186 717 2187
rect 726 2187 727 2188
rect 731 2187 732 2191
rect 726 2186 732 2187
rect 759 2191 765 2192
rect 759 2187 760 2191
rect 764 2190 765 2191
rect 782 2191 788 2192
rect 782 2190 783 2191
rect 764 2188 783 2190
rect 764 2187 765 2188
rect 759 2186 765 2187
rect 782 2187 783 2188
rect 787 2187 788 2191
rect 782 2186 788 2187
rect 815 2191 821 2192
rect 815 2187 816 2191
rect 820 2190 821 2191
rect 838 2191 844 2192
rect 838 2190 839 2191
rect 820 2188 839 2190
rect 820 2187 821 2188
rect 815 2186 821 2187
rect 838 2187 839 2188
rect 843 2187 844 2191
rect 838 2186 844 2187
rect 871 2191 877 2192
rect 871 2187 872 2191
rect 876 2190 877 2191
rect 894 2191 900 2192
rect 894 2190 895 2191
rect 876 2188 895 2190
rect 876 2187 877 2188
rect 871 2186 877 2187
rect 894 2187 895 2188
rect 899 2187 900 2191
rect 894 2186 900 2187
rect 910 2191 916 2192
rect 910 2187 911 2191
rect 915 2190 916 2191
rect 927 2191 933 2192
rect 927 2190 928 2191
rect 915 2188 928 2190
rect 915 2187 916 2188
rect 910 2186 916 2187
rect 927 2187 928 2188
rect 932 2187 933 2191
rect 927 2186 933 2187
rect 1094 2188 1100 2189
rect 110 2183 116 2184
rect 1094 2184 1095 2188
rect 1099 2184 1100 2188
rect 1094 2183 1100 2184
rect 1134 2187 1140 2188
rect 1134 2183 1135 2187
rect 1139 2183 1140 2187
rect 2118 2187 2124 2188
rect 1134 2182 1140 2183
rect 1686 2184 1692 2185
rect 134 2180 140 2181
rect 134 2176 135 2180
rect 139 2176 140 2180
rect 134 2175 140 2176
rect 174 2180 180 2181
rect 174 2176 175 2180
rect 179 2176 180 2180
rect 174 2175 180 2176
rect 214 2180 220 2181
rect 214 2176 215 2180
rect 219 2176 220 2180
rect 214 2175 220 2176
rect 254 2180 260 2181
rect 254 2176 255 2180
rect 259 2176 260 2180
rect 254 2175 260 2176
rect 318 2180 324 2181
rect 318 2176 319 2180
rect 323 2176 324 2180
rect 318 2175 324 2176
rect 382 2180 388 2181
rect 382 2176 383 2180
rect 387 2176 388 2180
rect 382 2175 388 2176
rect 446 2180 452 2181
rect 446 2176 447 2180
rect 451 2176 452 2180
rect 446 2175 452 2176
rect 510 2180 516 2181
rect 510 2176 511 2180
rect 515 2176 516 2180
rect 510 2175 516 2176
rect 574 2180 580 2181
rect 574 2176 575 2180
rect 579 2176 580 2180
rect 574 2175 580 2176
rect 630 2180 636 2181
rect 630 2176 631 2180
rect 635 2176 636 2180
rect 630 2175 636 2176
rect 686 2180 692 2181
rect 686 2176 687 2180
rect 691 2176 692 2180
rect 686 2175 692 2176
rect 734 2180 740 2181
rect 734 2176 735 2180
rect 739 2176 740 2180
rect 734 2175 740 2176
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 846 2180 852 2181
rect 846 2176 847 2180
rect 851 2176 852 2180
rect 846 2175 852 2176
rect 902 2180 908 2181
rect 902 2176 903 2180
rect 907 2176 908 2180
rect 1686 2180 1687 2184
rect 1691 2180 1692 2184
rect 1686 2179 1692 2180
rect 1726 2184 1732 2185
rect 1726 2180 1727 2184
rect 1731 2180 1732 2184
rect 1726 2179 1732 2180
rect 1766 2184 1772 2185
rect 1766 2180 1767 2184
rect 1771 2180 1772 2184
rect 1766 2179 1772 2180
rect 1806 2184 1812 2185
rect 1806 2180 1807 2184
rect 1811 2180 1812 2184
rect 2118 2183 2119 2187
rect 2123 2183 2124 2187
rect 2118 2182 2124 2183
rect 1806 2179 1812 2180
rect 902 2175 908 2176
rect 1158 2172 1164 2173
rect 1134 2169 1140 2170
rect 162 2167 168 2168
rect 162 2163 163 2167
rect 167 2166 168 2167
rect 171 2167 177 2168
rect 171 2166 172 2167
rect 167 2164 172 2166
rect 167 2163 168 2164
rect 162 2162 168 2163
rect 171 2163 172 2164
rect 176 2163 177 2167
rect 171 2162 177 2163
rect 202 2167 208 2168
rect 202 2163 203 2167
rect 207 2166 208 2167
rect 211 2167 217 2168
rect 211 2166 212 2167
rect 207 2164 212 2166
rect 207 2163 208 2164
rect 202 2162 208 2163
rect 211 2163 212 2164
rect 216 2163 217 2167
rect 211 2162 217 2163
rect 242 2167 248 2168
rect 242 2163 243 2167
rect 247 2166 248 2167
rect 251 2167 257 2168
rect 251 2166 252 2167
rect 247 2164 252 2166
rect 247 2163 248 2164
rect 242 2162 248 2163
rect 251 2163 252 2164
rect 256 2163 257 2167
rect 251 2162 257 2163
rect 310 2167 321 2168
rect 310 2163 311 2167
rect 315 2163 316 2167
rect 320 2163 321 2167
rect 310 2162 321 2163
rect 374 2167 385 2168
rect 374 2163 375 2167
rect 379 2163 380 2167
rect 384 2163 385 2167
rect 374 2162 385 2163
rect 438 2167 449 2168
rect 438 2163 439 2167
rect 443 2163 444 2167
rect 448 2163 449 2167
rect 438 2162 449 2163
rect 507 2167 513 2168
rect 507 2163 508 2167
rect 512 2166 513 2167
rect 543 2167 549 2168
rect 543 2166 544 2167
rect 512 2164 544 2166
rect 512 2163 513 2164
rect 507 2162 513 2163
rect 543 2163 544 2164
rect 548 2163 549 2167
rect 543 2162 549 2163
rect 566 2167 577 2168
rect 566 2163 567 2167
rect 571 2163 572 2167
rect 576 2163 577 2167
rect 566 2162 577 2163
rect 622 2167 633 2168
rect 622 2163 623 2167
rect 627 2163 628 2167
rect 632 2163 633 2167
rect 622 2162 633 2163
rect 678 2167 689 2168
rect 678 2163 679 2167
rect 683 2163 684 2167
rect 688 2163 689 2167
rect 678 2162 689 2163
rect 726 2167 737 2168
rect 726 2163 727 2167
rect 731 2163 732 2167
rect 736 2163 737 2167
rect 726 2162 737 2163
rect 782 2167 793 2168
rect 782 2163 783 2167
rect 787 2163 788 2167
rect 792 2163 793 2167
rect 782 2162 793 2163
rect 838 2167 849 2168
rect 838 2163 839 2167
rect 843 2163 844 2167
rect 848 2163 849 2167
rect 838 2162 849 2163
rect 894 2167 905 2168
rect 894 2163 895 2167
rect 899 2163 900 2167
rect 904 2163 905 2167
rect 1134 2165 1135 2169
rect 1139 2165 1140 2169
rect 1158 2168 1159 2172
rect 1163 2168 1164 2172
rect 1158 2167 1164 2168
rect 1198 2172 1204 2173
rect 1198 2168 1199 2172
rect 1203 2168 1204 2172
rect 1198 2167 1204 2168
rect 1238 2172 1244 2173
rect 1238 2168 1239 2172
rect 1243 2168 1244 2172
rect 1238 2167 1244 2168
rect 1278 2172 1284 2173
rect 1278 2168 1279 2172
rect 1283 2168 1284 2172
rect 1278 2167 1284 2168
rect 1334 2172 1340 2173
rect 1334 2168 1335 2172
rect 1339 2168 1340 2172
rect 1334 2167 1340 2168
rect 1390 2172 1396 2173
rect 1390 2168 1391 2172
rect 1395 2168 1396 2172
rect 1390 2167 1396 2168
rect 1454 2172 1460 2173
rect 1454 2168 1455 2172
rect 1459 2168 1460 2172
rect 1454 2167 1460 2168
rect 1526 2172 1532 2173
rect 1526 2168 1527 2172
rect 1531 2168 1532 2172
rect 1526 2167 1532 2168
rect 1590 2172 1596 2173
rect 1590 2168 1591 2172
rect 1595 2168 1596 2172
rect 1590 2167 1596 2168
rect 1662 2172 1668 2173
rect 1662 2168 1663 2172
rect 1667 2168 1668 2172
rect 1662 2167 1668 2168
rect 1734 2172 1740 2173
rect 1734 2168 1735 2172
rect 1739 2168 1740 2172
rect 1734 2167 1740 2168
rect 1806 2172 1812 2173
rect 1806 2168 1807 2172
rect 1811 2168 1812 2172
rect 1806 2167 1812 2168
rect 1878 2172 1884 2173
rect 1878 2168 1879 2172
rect 1883 2168 1884 2172
rect 1878 2167 1884 2168
rect 2118 2169 2124 2170
rect 1134 2164 1140 2165
rect 2118 2165 2119 2169
rect 2123 2165 2124 2169
rect 2118 2164 2124 2165
rect 894 2162 905 2163
rect 1318 2163 1324 2164
rect 1318 2162 1319 2163
rect 1176 2160 1319 2162
rect 1174 2159 1180 2160
rect 454 2155 460 2156
rect 454 2154 455 2155
rect 228 2152 455 2154
rect 228 2150 230 2152
rect 454 2151 455 2152
rect 459 2151 460 2155
rect 910 2155 916 2156
rect 910 2154 911 2155
rect 454 2150 460 2151
rect 796 2152 911 2154
rect 796 2150 798 2152
rect 910 2151 911 2152
rect 915 2151 916 2155
rect 1174 2155 1175 2159
rect 1179 2155 1180 2159
rect 1318 2159 1319 2160
rect 1323 2159 1324 2163
rect 1318 2158 1324 2159
rect 1766 2163 1772 2164
rect 1766 2159 1767 2163
rect 1771 2162 1772 2163
rect 1771 2160 1882 2162
rect 1771 2159 1772 2160
rect 1766 2158 1772 2159
rect 1174 2154 1180 2155
rect 1183 2155 1192 2156
rect 910 2150 916 2151
rect 1134 2152 1140 2153
rect 227 2149 233 2150
rect 227 2145 228 2149
rect 232 2145 233 2149
rect 795 2149 801 2150
rect 227 2144 233 2145
rect 267 2147 273 2148
rect 267 2143 268 2147
rect 272 2143 273 2147
rect 267 2142 273 2143
rect 298 2147 304 2148
rect 298 2143 299 2147
rect 303 2146 304 2147
rect 307 2147 313 2148
rect 307 2146 308 2147
rect 303 2144 308 2146
rect 303 2143 304 2144
rect 298 2142 304 2143
rect 307 2143 308 2144
rect 312 2143 313 2147
rect 307 2142 313 2143
rect 338 2147 344 2148
rect 338 2143 339 2147
rect 343 2146 344 2147
rect 355 2147 361 2148
rect 355 2146 356 2147
rect 343 2144 356 2146
rect 343 2143 344 2144
rect 338 2142 344 2143
rect 355 2143 356 2144
rect 360 2143 361 2147
rect 419 2147 425 2148
rect 419 2146 420 2147
rect 384 2144 420 2146
rect 355 2142 361 2143
rect 382 2143 388 2144
rect 257 2140 271 2142
rect 230 2136 236 2137
rect 230 2132 231 2136
rect 235 2132 236 2136
rect 230 2131 236 2132
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 257 2126 259 2140
rect 382 2139 383 2143
rect 387 2139 388 2143
rect 419 2143 420 2144
rect 424 2143 425 2147
rect 419 2142 425 2143
rect 455 2147 461 2148
rect 455 2143 456 2147
rect 460 2146 461 2147
rect 483 2147 489 2148
rect 483 2146 484 2147
rect 460 2144 484 2146
rect 460 2143 461 2144
rect 455 2142 461 2143
rect 483 2143 484 2144
rect 488 2143 489 2147
rect 483 2142 489 2143
rect 555 2147 561 2148
rect 555 2143 556 2147
rect 560 2146 561 2147
rect 623 2147 629 2148
rect 623 2146 624 2147
rect 560 2144 624 2146
rect 560 2143 561 2144
rect 555 2142 561 2143
rect 623 2143 624 2144
rect 628 2143 629 2147
rect 623 2142 629 2143
rect 635 2147 641 2148
rect 635 2143 636 2147
rect 640 2146 641 2147
rect 687 2147 693 2148
rect 687 2146 688 2147
rect 640 2144 688 2146
rect 640 2143 641 2144
rect 635 2142 641 2143
rect 687 2143 688 2144
rect 692 2143 693 2147
rect 687 2142 693 2143
rect 715 2147 721 2148
rect 715 2143 716 2147
rect 720 2146 721 2147
rect 726 2147 732 2148
rect 726 2146 727 2147
rect 720 2144 727 2146
rect 720 2143 721 2144
rect 715 2142 721 2143
rect 726 2143 727 2144
rect 731 2143 732 2147
rect 795 2145 796 2149
rect 800 2145 801 2149
rect 1134 2148 1135 2152
rect 1139 2148 1140 2152
rect 1183 2151 1184 2155
rect 1191 2151 1192 2155
rect 1183 2150 1192 2151
rect 1223 2155 1232 2156
rect 1223 2151 1224 2155
rect 1231 2151 1232 2155
rect 1223 2150 1232 2151
rect 1263 2155 1272 2156
rect 1263 2151 1264 2155
rect 1271 2151 1272 2155
rect 1263 2150 1272 2151
rect 1303 2155 1309 2156
rect 1303 2151 1304 2155
rect 1308 2154 1309 2155
rect 1326 2155 1332 2156
rect 1326 2154 1327 2155
rect 1308 2152 1327 2154
rect 1308 2151 1309 2152
rect 1303 2150 1309 2151
rect 1326 2151 1327 2152
rect 1331 2151 1332 2155
rect 1326 2150 1332 2151
rect 1359 2155 1365 2156
rect 1359 2151 1360 2155
rect 1364 2154 1365 2155
rect 1382 2155 1388 2156
rect 1382 2154 1383 2155
rect 1364 2152 1383 2154
rect 1364 2151 1365 2152
rect 1359 2150 1365 2151
rect 1382 2151 1383 2152
rect 1387 2151 1388 2155
rect 1382 2150 1388 2151
rect 1415 2155 1421 2156
rect 1415 2151 1416 2155
rect 1420 2154 1421 2155
rect 1446 2155 1452 2156
rect 1446 2154 1447 2155
rect 1420 2152 1447 2154
rect 1420 2151 1421 2152
rect 1415 2150 1421 2151
rect 1446 2151 1447 2152
rect 1451 2151 1452 2155
rect 1446 2150 1452 2151
rect 1479 2155 1485 2156
rect 1479 2151 1480 2155
rect 1484 2154 1485 2155
rect 1498 2155 1504 2156
rect 1498 2154 1499 2155
rect 1484 2152 1499 2154
rect 1484 2151 1485 2152
rect 1479 2150 1485 2151
rect 1498 2151 1499 2152
rect 1503 2151 1504 2155
rect 1498 2150 1504 2151
rect 1534 2155 1540 2156
rect 1534 2151 1535 2155
rect 1539 2154 1540 2155
rect 1551 2155 1557 2156
rect 1551 2154 1552 2155
rect 1539 2152 1552 2154
rect 1539 2151 1540 2152
rect 1534 2150 1540 2151
rect 1551 2151 1552 2152
rect 1556 2151 1557 2155
rect 1551 2150 1557 2151
rect 1615 2155 1621 2156
rect 1615 2151 1616 2155
rect 1620 2154 1621 2155
rect 1654 2155 1660 2156
rect 1654 2154 1655 2155
rect 1620 2152 1655 2154
rect 1620 2151 1621 2152
rect 1615 2150 1621 2151
rect 1654 2151 1655 2152
rect 1659 2151 1660 2155
rect 1654 2150 1660 2151
rect 1678 2155 1684 2156
rect 1678 2151 1679 2155
rect 1683 2154 1684 2155
rect 1687 2155 1693 2156
rect 1687 2154 1688 2155
rect 1683 2152 1688 2154
rect 1683 2151 1684 2152
rect 1678 2150 1684 2151
rect 1687 2151 1688 2152
rect 1692 2151 1693 2155
rect 1687 2150 1693 2151
rect 1758 2155 1765 2156
rect 1758 2151 1759 2155
rect 1764 2151 1765 2155
rect 1758 2150 1765 2151
rect 1831 2155 1837 2156
rect 1831 2151 1832 2155
rect 1836 2154 1837 2155
rect 1870 2155 1876 2156
rect 1870 2154 1871 2155
rect 1836 2152 1871 2154
rect 1836 2151 1837 2152
rect 1831 2150 1837 2151
rect 1870 2151 1871 2152
rect 1875 2151 1876 2155
rect 1880 2154 1882 2160
rect 1903 2155 1909 2156
rect 1903 2154 1904 2155
rect 1880 2152 1904 2154
rect 1870 2150 1876 2151
rect 1903 2151 1904 2152
rect 1908 2151 1909 2155
rect 1903 2150 1909 2151
rect 2118 2152 2124 2153
rect 795 2144 801 2145
rect 826 2147 832 2148
rect 726 2142 732 2143
rect 826 2143 827 2147
rect 831 2146 832 2147
rect 875 2147 881 2148
rect 875 2146 876 2147
rect 831 2144 876 2146
rect 831 2143 832 2144
rect 826 2142 832 2143
rect 875 2143 876 2144
rect 880 2143 881 2147
rect 963 2147 969 2148
rect 1134 2147 1140 2148
rect 2118 2148 2119 2152
rect 2123 2148 2124 2152
rect 2118 2147 2124 2148
rect 963 2146 964 2147
rect 875 2142 881 2143
rect 919 2144 964 2146
rect 382 2138 388 2139
rect 270 2136 276 2137
rect 270 2132 271 2136
rect 275 2132 276 2136
rect 270 2131 276 2132
rect 310 2136 316 2137
rect 310 2132 311 2136
rect 315 2132 316 2136
rect 310 2131 316 2132
rect 358 2136 364 2137
rect 358 2132 359 2136
rect 363 2132 364 2136
rect 358 2131 364 2132
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 486 2136 492 2137
rect 486 2132 487 2136
rect 491 2132 492 2136
rect 486 2131 492 2132
rect 558 2136 564 2137
rect 558 2132 559 2136
rect 563 2132 564 2136
rect 558 2131 564 2132
rect 638 2136 644 2137
rect 638 2132 639 2136
rect 643 2132 644 2136
rect 638 2131 644 2132
rect 718 2136 724 2137
rect 718 2132 719 2136
rect 723 2132 724 2136
rect 718 2131 724 2132
rect 798 2136 804 2137
rect 798 2132 799 2136
rect 803 2132 804 2136
rect 798 2131 804 2132
rect 878 2136 884 2137
rect 878 2132 879 2136
rect 883 2132 884 2136
rect 878 2131 884 2132
rect 919 2130 921 2144
rect 963 2143 964 2144
rect 968 2143 969 2147
rect 963 2142 969 2143
rect 1158 2144 1164 2145
rect 1158 2140 1159 2144
rect 1163 2140 1164 2144
rect 1158 2139 1164 2140
rect 1198 2144 1204 2145
rect 1198 2140 1199 2144
rect 1203 2140 1204 2144
rect 1198 2139 1204 2140
rect 1238 2144 1244 2145
rect 1238 2140 1239 2144
rect 1243 2140 1244 2144
rect 1238 2139 1244 2140
rect 1278 2144 1284 2145
rect 1278 2140 1279 2144
rect 1283 2140 1284 2144
rect 1278 2139 1284 2140
rect 1334 2144 1340 2145
rect 1334 2140 1335 2144
rect 1339 2140 1340 2144
rect 1334 2139 1340 2140
rect 1390 2144 1396 2145
rect 1390 2140 1391 2144
rect 1395 2140 1396 2144
rect 1390 2139 1396 2140
rect 1454 2144 1460 2145
rect 1454 2140 1455 2144
rect 1459 2140 1460 2144
rect 1454 2139 1460 2140
rect 1526 2144 1532 2145
rect 1526 2140 1527 2144
rect 1531 2140 1532 2144
rect 1526 2139 1532 2140
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1662 2144 1668 2145
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1734 2144 1740 2145
rect 1734 2140 1735 2144
rect 1739 2140 1740 2144
rect 1734 2139 1740 2140
rect 1806 2144 1812 2145
rect 1806 2140 1807 2144
rect 1811 2140 1812 2144
rect 1806 2139 1812 2140
rect 1878 2144 1884 2145
rect 1878 2140 1879 2144
rect 1883 2140 1884 2144
rect 1878 2139 1884 2140
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1155 2131 1161 2132
rect 905 2128 921 2130
rect 1094 2128 1100 2129
rect 905 2126 907 2128
rect 110 2123 116 2124
rect 255 2125 261 2126
rect 255 2121 256 2125
rect 260 2121 261 2125
rect 903 2125 909 2126
rect 255 2120 261 2121
rect 295 2123 304 2124
rect 295 2119 296 2123
rect 303 2119 304 2123
rect 295 2118 304 2119
rect 335 2123 344 2124
rect 335 2119 336 2123
rect 343 2119 344 2123
rect 335 2118 344 2119
rect 382 2123 389 2124
rect 382 2119 383 2123
rect 388 2119 389 2123
rect 382 2118 389 2119
rect 447 2123 453 2124
rect 447 2119 448 2123
rect 452 2122 453 2123
rect 455 2123 461 2124
rect 455 2122 456 2123
rect 452 2120 456 2122
rect 452 2119 453 2120
rect 447 2118 453 2119
rect 455 2119 456 2120
rect 460 2119 461 2123
rect 455 2118 461 2119
rect 478 2123 484 2124
rect 478 2119 479 2123
rect 483 2122 484 2123
rect 511 2123 517 2124
rect 511 2122 512 2123
rect 483 2120 512 2122
rect 483 2119 484 2120
rect 478 2118 484 2119
rect 511 2119 512 2120
rect 516 2119 517 2123
rect 511 2118 517 2119
rect 543 2123 549 2124
rect 543 2119 544 2123
rect 548 2122 549 2123
rect 583 2123 589 2124
rect 583 2122 584 2123
rect 548 2120 584 2122
rect 548 2119 549 2120
rect 543 2118 549 2119
rect 583 2119 584 2120
rect 588 2119 589 2123
rect 583 2118 589 2119
rect 623 2123 629 2124
rect 623 2119 624 2123
rect 628 2122 629 2123
rect 663 2123 669 2124
rect 663 2122 664 2123
rect 628 2120 664 2122
rect 628 2119 629 2120
rect 623 2118 629 2119
rect 663 2119 664 2120
rect 668 2119 669 2123
rect 663 2118 669 2119
rect 687 2123 693 2124
rect 687 2119 688 2123
rect 692 2122 693 2123
rect 743 2123 749 2124
rect 743 2122 744 2123
rect 692 2120 744 2122
rect 692 2119 693 2120
rect 687 2118 693 2119
rect 743 2119 744 2120
rect 748 2119 749 2123
rect 743 2118 749 2119
rect 823 2123 832 2124
rect 823 2119 824 2123
rect 831 2119 832 2123
rect 903 2121 904 2125
rect 908 2121 909 2125
rect 1094 2124 1095 2128
rect 1099 2124 1100 2128
rect 1155 2127 1156 2131
rect 1160 2130 1161 2131
rect 1174 2131 1180 2132
rect 1174 2130 1175 2131
rect 1160 2128 1175 2130
rect 1160 2127 1161 2128
rect 1155 2126 1161 2127
rect 1174 2127 1175 2128
rect 1179 2127 1180 2131
rect 1174 2126 1180 2127
rect 1186 2131 1192 2132
rect 1186 2127 1187 2131
rect 1191 2130 1192 2131
rect 1195 2131 1201 2132
rect 1195 2130 1196 2131
rect 1191 2128 1196 2130
rect 1191 2127 1192 2128
rect 1186 2126 1192 2127
rect 1195 2127 1196 2128
rect 1200 2127 1201 2131
rect 1195 2126 1201 2127
rect 1226 2131 1232 2132
rect 1226 2127 1227 2131
rect 1231 2130 1232 2131
rect 1235 2131 1241 2132
rect 1235 2130 1236 2131
rect 1231 2128 1236 2130
rect 1231 2127 1232 2128
rect 1226 2126 1232 2127
rect 1235 2127 1236 2128
rect 1240 2127 1241 2131
rect 1235 2126 1241 2127
rect 1266 2131 1272 2132
rect 1266 2127 1267 2131
rect 1271 2130 1272 2131
rect 1275 2131 1281 2132
rect 1275 2130 1276 2131
rect 1271 2128 1276 2130
rect 1271 2127 1272 2128
rect 1266 2126 1272 2127
rect 1275 2127 1276 2128
rect 1280 2127 1281 2131
rect 1275 2126 1281 2127
rect 1326 2131 1337 2132
rect 1326 2127 1327 2131
rect 1331 2127 1332 2131
rect 1336 2127 1337 2131
rect 1326 2126 1337 2127
rect 1382 2131 1393 2132
rect 1382 2127 1383 2131
rect 1387 2127 1388 2131
rect 1392 2127 1393 2131
rect 1382 2126 1393 2127
rect 1446 2131 1457 2132
rect 1446 2127 1447 2131
rect 1451 2127 1452 2131
rect 1456 2127 1457 2131
rect 1446 2126 1457 2127
rect 1498 2131 1504 2132
rect 1498 2127 1499 2131
rect 1503 2130 1504 2131
rect 1523 2131 1529 2132
rect 1523 2130 1524 2131
rect 1503 2128 1524 2130
rect 1503 2127 1504 2128
rect 1498 2126 1504 2127
rect 1523 2127 1524 2128
rect 1528 2127 1529 2131
rect 1523 2126 1529 2127
rect 1587 2131 1593 2132
rect 1587 2127 1588 2131
rect 1592 2130 1593 2131
rect 1646 2131 1652 2132
rect 1646 2130 1647 2131
rect 1592 2128 1647 2130
rect 1592 2127 1593 2128
rect 1587 2126 1593 2127
rect 1646 2127 1647 2128
rect 1651 2127 1652 2131
rect 1646 2126 1652 2127
rect 1654 2131 1665 2132
rect 1654 2127 1655 2131
rect 1659 2127 1660 2131
rect 1664 2127 1665 2131
rect 1654 2126 1665 2127
rect 1731 2131 1737 2132
rect 1731 2127 1732 2131
rect 1736 2130 1737 2131
rect 1766 2131 1772 2132
rect 1766 2130 1767 2131
rect 1736 2128 1767 2130
rect 1736 2127 1737 2128
rect 1731 2126 1737 2127
rect 1766 2127 1767 2128
rect 1771 2127 1772 2131
rect 1766 2126 1772 2127
rect 1803 2131 1809 2132
rect 1803 2127 1804 2131
rect 1808 2130 1809 2131
rect 1814 2131 1820 2132
rect 1814 2130 1815 2131
rect 1808 2128 1815 2130
rect 1808 2127 1809 2128
rect 1803 2126 1809 2127
rect 1814 2127 1815 2128
rect 1819 2127 1820 2131
rect 1814 2126 1820 2127
rect 1870 2131 1881 2132
rect 1870 2127 1871 2131
rect 1875 2127 1876 2131
rect 1880 2127 1881 2131
rect 1870 2126 1881 2127
rect 903 2120 909 2121
rect 991 2123 997 2124
rect 823 2118 832 2119
rect 991 2119 992 2123
rect 996 2122 997 2123
rect 1030 2123 1036 2124
rect 1094 2123 1100 2124
rect 1030 2122 1031 2123
rect 996 2120 1031 2122
rect 996 2119 997 2120
rect 991 2118 997 2119
rect 1030 2119 1031 2120
rect 1035 2119 1036 2123
rect 1030 2118 1036 2119
rect 1155 2119 1161 2120
rect 1155 2115 1156 2119
rect 1160 2118 1161 2119
rect 1178 2119 1184 2120
rect 1178 2118 1179 2119
rect 1160 2116 1179 2118
rect 1160 2115 1161 2116
rect 1155 2114 1161 2115
rect 1178 2115 1179 2116
rect 1183 2115 1184 2119
rect 1178 2114 1184 2115
rect 1186 2119 1192 2120
rect 1186 2115 1187 2119
rect 1191 2118 1192 2119
rect 1195 2119 1201 2120
rect 1195 2118 1196 2119
rect 1191 2116 1196 2118
rect 1191 2115 1192 2116
rect 1186 2114 1192 2115
rect 1195 2115 1196 2116
rect 1200 2115 1201 2119
rect 1195 2114 1201 2115
rect 1226 2119 1232 2120
rect 1226 2115 1227 2119
rect 1231 2118 1232 2119
rect 1235 2119 1241 2120
rect 1235 2118 1236 2119
rect 1231 2116 1236 2118
rect 1231 2115 1232 2116
rect 1226 2114 1232 2115
rect 1235 2115 1236 2116
rect 1240 2115 1241 2119
rect 1235 2114 1241 2115
rect 1266 2119 1272 2120
rect 1266 2115 1267 2119
rect 1271 2118 1272 2119
rect 1291 2119 1297 2120
rect 1291 2118 1292 2119
rect 1271 2116 1292 2118
rect 1271 2115 1272 2116
rect 1266 2114 1272 2115
rect 1291 2115 1292 2116
rect 1296 2115 1297 2119
rect 1291 2114 1297 2115
rect 1363 2119 1369 2120
rect 1363 2115 1364 2119
rect 1368 2118 1369 2119
rect 1402 2119 1408 2120
rect 1368 2116 1394 2118
rect 1368 2115 1369 2116
rect 1363 2114 1369 2115
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 1094 2111 1100 2112
rect 110 2106 116 2107
rect 230 2108 236 2109
rect 230 2104 231 2108
rect 235 2104 236 2108
rect 230 2103 236 2104
rect 270 2108 276 2109
rect 270 2104 271 2108
rect 275 2104 276 2108
rect 270 2103 276 2104
rect 310 2108 316 2109
rect 310 2104 311 2108
rect 315 2104 316 2108
rect 310 2103 316 2104
rect 358 2108 364 2109
rect 358 2104 359 2108
rect 363 2104 364 2108
rect 358 2103 364 2104
rect 422 2108 428 2109
rect 422 2104 423 2108
rect 427 2104 428 2108
rect 422 2103 428 2104
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 558 2108 564 2109
rect 558 2104 559 2108
rect 563 2104 564 2108
rect 558 2103 564 2104
rect 638 2108 644 2109
rect 638 2104 639 2108
rect 643 2104 644 2108
rect 638 2103 644 2104
rect 718 2108 724 2109
rect 718 2104 719 2108
rect 723 2104 724 2108
rect 718 2103 724 2104
rect 798 2108 804 2109
rect 798 2104 799 2108
rect 803 2104 804 2108
rect 798 2103 804 2104
rect 878 2108 884 2109
rect 878 2104 879 2108
rect 883 2104 884 2108
rect 878 2103 884 2104
rect 966 2108 972 2109
rect 966 2104 967 2108
rect 971 2104 972 2108
rect 1094 2107 1095 2111
rect 1099 2107 1100 2111
rect 1094 2106 1100 2107
rect 1158 2108 1164 2109
rect 966 2103 972 2104
rect 1158 2104 1159 2108
rect 1163 2104 1164 2108
rect 1158 2103 1164 2104
rect 1198 2108 1204 2109
rect 1198 2104 1199 2108
rect 1203 2104 1204 2108
rect 1198 2103 1204 2104
rect 1238 2108 1244 2109
rect 1238 2104 1239 2108
rect 1243 2104 1244 2108
rect 1238 2103 1244 2104
rect 1294 2108 1300 2109
rect 1294 2104 1295 2108
rect 1299 2104 1300 2108
rect 1294 2103 1300 2104
rect 1366 2108 1372 2109
rect 1366 2104 1367 2108
rect 1371 2104 1372 2108
rect 1392 2106 1394 2116
rect 1402 2115 1403 2119
rect 1407 2118 1408 2119
rect 1435 2119 1441 2120
rect 1435 2118 1436 2119
rect 1407 2116 1436 2118
rect 1407 2115 1408 2116
rect 1402 2114 1408 2115
rect 1435 2115 1436 2116
rect 1440 2115 1441 2119
rect 1435 2114 1441 2115
rect 1515 2119 1521 2120
rect 1515 2115 1516 2119
rect 1520 2118 1521 2119
rect 1534 2119 1540 2120
rect 1534 2118 1535 2119
rect 1520 2116 1535 2118
rect 1520 2115 1521 2116
rect 1515 2114 1521 2115
rect 1534 2115 1535 2116
rect 1539 2115 1540 2119
rect 1534 2114 1540 2115
rect 1595 2119 1601 2120
rect 1595 2115 1596 2119
rect 1600 2118 1601 2119
rect 1614 2119 1620 2120
rect 1614 2118 1615 2119
rect 1600 2116 1615 2118
rect 1600 2115 1601 2116
rect 1595 2114 1601 2115
rect 1614 2115 1615 2116
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1626 2119 1632 2120
rect 1626 2115 1627 2119
rect 1631 2118 1632 2119
rect 1675 2119 1681 2120
rect 1675 2118 1676 2119
rect 1631 2116 1676 2118
rect 1631 2115 1632 2116
rect 1626 2114 1632 2115
rect 1675 2115 1676 2116
rect 1680 2115 1681 2119
rect 1675 2114 1681 2115
rect 1747 2119 1753 2120
rect 1747 2115 1748 2119
rect 1752 2118 1753 2119
rect 1758 2119 1764 2120
rect 1758 2118 1759 2119
rect 1752 2116 1759 2118
rect 1752 2115 1753 2116
rect 1747 2114 1753 2115
rect 1758 2115 1759 2116
rect 1763 2115 1764 2119
rect 1758 2114 1764 2115
rect 1798 2119 1804 2120
rect 1798 2115 1799 2119
rect 1803 2118 1804 2119
rect 1819 2119 1825 2120
rect 1819 2118 1820 2119
rect 1803 2116 1820 2118
rect 1803 2115 1804 2116
rect 1798 2114 1804 2115
rect 1819 2115 1820 2116
rect 1824 2115 1825 2119
rect 1819 2114 1825 2115
rect 1866 2119 1872 2120
rect 1866 2115 1867 2119
rect 1871 2118 1872 2119
rect 1883 2119 1889 2120
rect 1883 2118 1884 2119
rect 1871 2116 1884 2118
rect 1871 2115 1872 2116
rect 1866 2114 1872 2115
rect 1883 2115 1884 2116
rect 1888 2115 1889 2119
rect 1883 2114 1889 2115
rect 1947 2119 1953 2120
rect 1947 2115 1948 2119
rect 1952 2118 1953 2119
rect 1982 2119 1988 2120
rect 1982 2118 1983 2119
rect 1952 2116 1983 2118
rect 1952 2115 1953 2116
rect 1947 2114 1953 2115
rect 1982 2115 1983 2116
rect 1987 2115 1988 2119
rect 1982 2114 1988 2115
rect 1994 2119 2000 2120
rect 1994 2115 1995 2119
rect 1999 2118 2000 2119
rect 2019 2119 2025 2120
rect 2019 2118 2020 2119
rect 1999 2116 2020 2118
rect 1999 2115 2000 2116
rect 1994 2114 2000 2115
rect 2019 2115 2020 2116
rect 2024 2115 2025 2119
rect 2019 2114 2025 2115
rect 2050 2119 2056 2120
rect 2050 2115 2051 2119
rect 2055 2118 2056 2119
rect 2067 2119 2073 2120
rect 2067 2118 2068 2119
rect 2055 2116 2068 2118
rect 2055 2115 2056 2116
rect 2050 2114 2056 2115
rect 2067 2115 2068 2116
rect 2072 2115 2073 2119
rect 2067 2114 2073 2115
rect 1438 2108 1444 2109
rect 1392 2104 1434 2106
rect 1366 2103 1372 2104
rect 1134 2100 1140 2101
rect 1134 2096 1135 2100
rect 1139 2096 1140 2100
rect 1432 2098 1434 2104
rect 1438 2104 1439 2108
rect 1443 2104 1444 2108
rect 1438 2103 1444 2104
rect 1518 2108 1524 2109
rect 1518 2104 1519 2108
rect 1523 2104 1524 2108
rect 1518 2103 1524 2104
rect 1598 2108 1604 2109
rect 1598 2104 1599 2108
rect 1603 2104 1604 2108
rect 1598 2103 1604 2104
rect 1678 2108 1684 2109
rect 1678 2104 1679 2108
rect 1683 2104 1684 2108
rect 1678 2103 1684 2104
rect 1750 2108 1756 2109
rect 1750 2104 1751 2108
rect 1755 2104 1756 2108
rect 1750 2103 1756 2104
rect 1822 2108 1828 2109
rect 1822 2104 1823 2108
rect 1827 2104 1828 2108
rect 1822 2103 1828 2104
rect 1886 2108 1892 2109
rect 1886 2104 1887 2108
rect 1891 2104 1892 2108
rect 1886 2103 1892 2104
rect 1950 2108 1956 2109
rect 1950 2104 1951 2108
rect 1955 2104 1956 2108
rect 1950 2103 1956 2104
rect 2022 2108 2028 2109
rect 2022 2104 2023 2108
rect 2027 2104 2028 2108
rect 2022 2103 2028 2104
rect 2070 2108 2076 2109
rect 2070 2104 2071 2108
rect 2075 2104 2076 2108
rect 2070 2103 2076 2104
rect 1456 2100 1498 2102
rect 1456 2098 1458 2100
rect 1432 2096 1458 2098
rect 1134 2095 1140 2096
rect 1183 2095 1192 2096
rect 302 2092 308 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 302 2088 303 2092
rect 307 2088 308 2092
rect 302 2087 308 2088
rect 350 2092 356 2093
rect 350 2088 351 2092
rect 355 2088 356 2092
rect 350 2087 356 2088
rect 406 2092 412 2093
rect 406 2088 407 2092
rect 411 2088 412 2092
rect 406 2087 412 2088
rect 470 2092 476 2093
rect 470 2088 471 2092
rect 475 2088 476 2092
rect 470 2087 476 2088
rect 542 2092 548 2093
rect 542 2088 543 2092
rect 547 2088 548 2092
rect 542 2087 548 2088
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 702 2092 708 2093
rect 702 2088 703 2092
rect 707 2088 708 2092
rect 702 2087 708 2088
rect 782 2092 788 2093
rect 782 2088 783 2092
rect 787 2088 788 2092
rect 782 2087 788 2088
rect 862 2092 868 2093
rect 862 2088 863 2092
rect 867 2088 868 2092
rect 862 2087 868 2088
rect 950 2092 956 2093
rect 950 2088 951 2092
rect 955 2088 956 2092
rect 950 2087 956 2088
rect 1038 2092 1044 2093
rect 1038 2088 1039 2092
rect 1043 2088 1044 2092
rect 1183 2091 1184 2095
rect 1191 2091 1192 2095
rect 1183 2090 1192 2091
rect 1223 2095 1232 2096
rect 1223 2091 1224 2095
rect 1231 2091 1232 2095
rect 1223 2090 1232 2091
rect 1263 2095 1272 2096
rect 1263 2091 1264 2095
rect 1271 2091 1272 2095
rect 1263 2090 1272 2091
rect 1318 2095 1325 2096
rect 1318 2091 1319 2095
rect 1324 2091 1325 2095
rect 1318 2090 1325 2091
rect 1391 2095 1397 2096
rect 1391 2091 1392 2095
rect 1396 2094 1397 2095
rect 1402 2095 1408 2096
rect 1402 2094 1403 2095
rect 1396 2092 1403 2094
rect 1396 2091 1397 2092
rect 1391 2090 1397 2091
rect 1402 2091 1403 2092
rect 1407 2091 1408 2095
rect 1402 2090 1408 2091
rect 1463 2095 1469 2096
rect 1463 2091 1464 2095
rect 1468 2094 1469 2095
rect 1486 2095 1492 2096
rect 1486 2094 1487 2095
rect 1468 2092 1487 2094
rect 1468 2091 1469 2092
rect 1463 2090 1469 2091
rect 1486 2091 1487 2092
rect 1491 2091 1492 2095
rect 1496 2094 1498 2100
rect 2118 2100 2124 2101
rect 2118 2096 2119 2100
rect 2123 2096 2124 2100
rect 1543 2095 1549 2096
rect 1543 2094 1544 2095
rect 1496 2092 1544 2094
rect 1486 2090 1492 2091
rect 1543 2091 1544 2092
rect 1548 2091 1549 2095
rect 1543 2090 1549 2091
rect 1623 2095 1632 2096
rect 1623 2091 1624 2095
rect 1631 2091 1632 2095
rect 1623 2090 1632 2091
rect 1646 2095 1652 2096
rect 1646 2091 1647 2095
rect 1651 2094 1652 2095
rect 1703 2095 1709 2096
rect 1703 2094 1704 2095
rect 1651 2092 1704 2094
rect 1651 2091 1652 2092
rect 1646 2090 1652 2091
rect 1703 2091 1704 2092
rect 1708 2091 1709 2095
rect 1703 2090 1709 2091
rect 1775 2095 1781 2096
rect 1775 2091 1776 2095
rect 1780 2094 1781 2095
rect 1798 2095 1804 2096
rect 1798 2094 1799 2095
rect 1780 2092 1799 2094
rect 1780 2091 1781 2092
rect 1775 2090 1781 2091
rect 1798 2091 1799 2092
rect 1803 2091 1804 2095
rect 1798 2090 1804 2091
rect 1847 2095 1853 2096
rect 1847 2091 1848 2095
rect 1852 2094 1853 2095
rect 1866 2095 1872 2096
rect 1866 2094 1867 2095
rect 1852 2092 1867 2094
rect 1852 2091 1853 2092
rect 1847 2090 1853 2091
rect 1866 2091 1867 2092
rect 1871 2091 1872 2095
rect 1866 2090 1872 2091
rect 1902 2095 1908 2096
rect 1902 2091 1903 2095
rect 1907 2094 1908 2095
rect 1911 2095 1917 2096
rect 1911 2094 1912 2095
rect 1907 2092 1912 2094
rect 1907 2091 1908 2092
rect 1902 2090 1908 2091
rect 1911 2091 1912 2092
rect 1916 2091 1917 2095
rect 1911 2090 1917 2091
rect 1975 2095 1981 2096
rect 1975 2091 1976 2095
rect 1980 2094 1981 2095
rect 1994 2095 2000 2096
rect 1994 2094 1995 2095
rect 1980 2092 1995 2094
rect 1980 2091 1981 2092
rect 1975 2090 1981 2091
rect 1994 2091 1995 2092
rect 1999 2091 2000 2095
rect 1994 2090 2000 2091
rect 2047 2095 2056 2096
rect 2047 2091 2048 2095
rect 2055 2091 2056 2095
rect 2047 2090 2056 2091
rect 2058 2095 2064 2096
rect 2058 2091 2059 2095
rect 2063 2094 2064 2095
rect 2095 2095 2101 2096
rect 2118 2095 2124 2096
rect 2095 2094 2096 2095
rect 2063 2092 2096 2094
rect 2063 2091 2064 2092
rect 2058 2090 2064 2091
rect 2095 2091 2096 2092
rect 2100 2091 2101 2095
rect 2095 2090 2101 2091
rect 1038 2087 1044 2088
rect 1094 2089 1100 2090
rect 110 2084 116 2085
rect 1094 2085 1095 2089
rect 1099 2085 1100 2089
rect 1094 2084 1100 2085
rect 1134 2083 1140 2084
rect 1134 2079 1135 2083
rect 1139 2079 1140 2083
rect 2118 2083 2124 2084
rect 1134 2078 1140 2079
rect 1158 2080 1164 2081
rect 1158 2076 1159 2080
rect 1163 2076 1164 2080
rect 286 2075 292 2076
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 286 2071 287 2075
rect 291 2074 292 2075
rect 327 2075 333 2076
rect 327 2074 328 2075
rect 291 2072 328 2074
rect 291 2071 292 2072
rect 286 2070 292 2071
rect 327 2071 328 2072
rect 332 2071 333 2075
rect 327 2070 333 2071
rect 375 2075 381 2076
rect 375 2071 376 2075
rect 380 2074 381 2075
rect 398 2075 404 2076
rect 398 2074 399 2075
rect 380 2072 399 2074
rect 380 2071 381 2072
rect 375 2070 381 2071
rect 398 2071 399 2072
rect 403 2071 404 2075
rect 398 2070 404 2071
rect 431 2075 437 2076
rect 431 2071 432 2075
rect 436 2074 437 2075
rect 462 2075 468 2076
rect 462 2074 463 2075
rect 436 2072 463 2074
rect 436 2071 437 2072
rect 431 2070 437 2071
rect 462 2071 463 2072
rect 467 2071 468 2075
rect 462 2070 468 2071
rect 495 2075 501 2076
rect 495 2071 496 2075
rect 500 2074 501 2075
rect 534 2075 540 2076
rect 534 2074 535 2075
rect 500 2072 535 2074
rect 500 2071 501 2072
rect 495 2070 501 2071
rect 534 2071 535 2072
rect 539 2071 540 2075
rect 534 2070 540 2071
rect 567 2075 573 2076
rect 567 2071 568 2075
rect 572 2074 573 2075
rect 614 2075 620 2076
rect 614 2074 615 2075
rect 572 2072 615 2074
rect 572 2071 573 2072
rect 567 2070 573 2071
rect 614 2071 615 2072
rect 619 2071 620 2075
rect 614 2070 620 2071
rect 630 2075 636 2076
rect 630 2071 631 2075
rect 635 2074 636 2075
rect 647 2075 653 2076
rect 647 2074 648 2075
rect 635 2072 648 2074
rect 635 2071 636 2072
rect 630 2070 636 2071
rect 647 2071 648 2072
rect 652 2071 653 2075
rect 647 2070 653 2071
rect 726 2075 733 2076
rect 726 2071 727 2075
rect 732 2071 733 2075
rect 726 2070 733 2071
rect 735 2075 741 2076
rect 735 2071 736 2075
rect 740 2074 741 2075
rect 807 2075 813 2076
rect 807 2074 808 2075
rect 740 2072 808 2074
rect 740 2071 741 2072
rect 735 2070 741 2071
rect 807 2071 808 2072
rect 812 2071 813 2075
rect 807 2070 813 2071
rect 822 2075 828 2076
rect 822 2071 823 2075
rect 827 2074 828 2075
rect 887 2075 893 2076
rect 887 2074 888 2075
rect 827 2072 888 2074
rect 827 2071 828 2072
rect 822 2070 828 2071
rect 887 2071 888 2072
rect 892 2071 893 2075
rect 887 2070 893 2071
rect 895 2075 901 2076
rect 895 2071 896 2075
rect 900 2074 901 2075
rect 975 2075 981 2076
rect 975 2074 976 2075
rect 900 2072 976 2074
rect 900 2071 901 2072
rect 895 2070 901 2071
rect 975 2071 976 2072
rect 980 2071 981 2075
rect 975 2070 981 2071
rect 983 2075 989 2076
rect 983 2071 984 2075
rect 988 2074 989 2075
rect 1063 2075 1069 2076
rect 1158 2075 1164 2076
rect 1198 2080 1204 2081
rect 1198 2076 1199 2080
rect 1203 2076 1204 2080
rect 1198 2075 1204 2076
rect 1238 2080 1244 2081
rect 1238 2076 1239 2080
rect 1243 2076 1244 2080
rect 1238 2075 1244 2076
rect 1294 2080 1300 2081
rect 1294 2076 1295 2080
rect 1299 2076 1300 2080
rect 1294 2075 1300 2076
rect 1366 2080 1372 2081
rect 1366 2076 1367 2080
rect 1371 2076 1372 2080
rect 1366 2075 1372 2076
rect 1438 2080 1444 2081
rect 1438 2076 1439 2080
rect 1443 2076 1444 2080
rect 1438 2075 1444 2076
rect 1518 2080 1524 2081
rect 1518 2076 1519 2080
rect 1523 2076 1524 2080
rect 1518 2075 1524 2076
rect 1598 2080 1604 2081
rect 1598 2076 1599 2080
rect 1603 2076 1604 2080
rect 1598 2075 1604 2076
rect 1678 2080 1684 2081
rect 1678 2076 1679 2080
rect 1683 2076 1684 2080
rect 1678 2075 1684 2076
rect 1750 2080 1756 2081
rect 1750 2076 1751 2080
rect 1755 2076 1756 2080
rect 1750 2075 1756 2076
rect 1822 2080 1828 2081
rect 1822 2076 1823 2080
rect 1827 2076 1828 2080
rect 1822 2075 1828 2076
rect 1886 2080 1892 2081
rect 1886 2076 1887 2080
rect 1891 2076 1892 2080
rect 1886 2075 1892 2076
rect 1950 2080 1956 2081
rect 1950 2076 1951 2080
rect 1955 2076 1956 2080
rect 1950 2075 1956 2076
rect 2022 2080 2028 2081
rect 2022 2076 2023 2080
rect 2027 2076 2028 2080
rect 2022 2075 2028 2076
rect 2070 2080 2076 2081
rect 2070 2076 2071 2080
rect 2075 2076 2076 2080
rect 2118 2079 2119 2083
rect 2123 2079 2124 2083
rect 2118 2078 2124 2079
rect 2070 2075 2076 2076
rect 1063 2074 1064 2075
rect 988 2072 1064 2074
rect 988 2071 989 2072
rect 983 2070 989 2071
rect 1063 2071 1064 2072
rect 1068 2071 1069 2075
rect 1063 2070 1069 2071
rect 1094 2072 1100 2073
rect 110 2067 116 2068
rect 1094 2068 1095 2072
rect 1099 2068 1100 2072
rect 1094 2067 1100 2068
rect 1158 2068 1164 2069
rect 1134 2065 1140 2066
rect 302 2064 308 2065
rect 302 2060 303 2064
rect 307 2060 308 2064
rect 302 2059 308 2060
rect 350 2064 356 2065
rect 350 2060 351 2064
rect 355 2060 356 2064
rect 350 2059 356 2060
rect 406 2064 412 2065
rect 406 2060 407 2064
rect 411 2060 412 2064
rect 406 2059 412 2060
rect 470 2064 476 2065
rect 470 2060 471 2064
rect 475 2060 476 2064
rect 470 2059 476 2060
rect 542 2064 548 2065
rect 542 2060 543 2064
rect 547 2060 548 2064
rect 542 2059 548 2060
rect 622 2064 628 2065
rect 622 2060 623 2064
rect 627 2060 628 2064
rect 622 2059 628 2060
rect 702 2064 708 2065
rect 702 2060 703 2064
rect 707 2060 708 2064
rect 702 2059 708 2060
rect 782 2064 788 2065
rect 782 2060 783 2064
rect 787 2060 788 2064
rect 782 2059 788 2060
rect 862 2064 868 2065
rect 862 2060 863 2064
rect 867 2060 868 2064
rect 862 2059 868 2060
rect 950 2064 956 2065
rect 950 2060 951 2064
rect 955 2060 956 2064
rect 950 2059 956 2060
rect 1038 2064 1044 2065
rect 1038 2060 1039 2064
rect 1043 2060 1044 2064
rect 1134 2061 1135 2065
rect 1139 2061 1140 2065
rect 1158 2064 1159 2068
rect 1163 2064 1164 2068
rect 1158 2063 1164 2064
rect 1214 2068 1220 2069
rect 1214 2064 1215 2068
rect 1219 2064 1220 2068
rect 1214 2063 1220 2064
rect 1302 2068 1308 2069
rect 1302 2064 1303 2068
rect 1307 2064 1308 2068
rect 1302 2063 1308 2064
rect 1398 2068 1404 2069
rect 1398 2064 1399 2068
rect 1403 2064 1404 2068
rect 1398 2063 1404 2064
rect 1494 2068 1500 2069
rect 1494 2064 1495 2068
rect 1499 2064 1500 2068
rect 1494 2063 1500 2064
rect 1590 2068 1596 2069
rect 1590 2064 1591 2068
rect 1595 2064 1596 2068
rect 1590 2063 1596 2064
rect 1678 2068 1684 2069
rect 1678 2064 1679 2068
rect 1683 2064 1684 2068
rect 1678 2063 1684 2064
rect 1758 2068 1764 2069
rect 1758 2064 1759 2068
rect 1763 2064 1764 2068
rect 1758 2063 1764 2064
rect 1830 2068 1836 2069
rect 1830 2064 1831 2068
rect 1835 2064 1836 2068
rect 1830 2063 1836 2064
rect 1894 2068 1900 2069
rect 1894 2064 1895 2068
rect 1899 2064 1900 2068
rect 1894 2063 1900 2064
rect 1958 2068 1964 2069
rect 1958 2064 1959 2068
rect 1963 2064 1964 2068
rect 1958 2063 1964 2064
rect 2022 2068 2028 2069
rect 2022 2064 2023 2068
rect 2027 2064 2028 2068
rect 2022 2063 2028 2064
rect 2070 2068 2076 2069
rect 2070 2064 2071 2068
rect 2075 2064 2076 2068
rect 2070 2063 2076 2064
rect 2118 2065 2124 2066
rect 1134 2060 1140 2061
rect 2118 2061 2119 2065
rect 2123 2061 2124 2065
rect 2118 2060 2124 2061
rect 1038 2059 1044 2060
rect 299 2051 305 2052
rect 299 2047 300 2051
rect 304 2050 305 2051
rect 347 2051 353 2052
rect 304 2048 321 2050
rect 304 2047 305 2048
rect 299 2046 305 2047
rect 319 2042 321 2048
rect 347 2047 348 2051
rect 352 2050 353 2051
rect 390 2051 396 2052
rect 390 2050 391 2051
rect 352 2048 391 2050
rect 352 2047 353 2048
rect 347 2046 353 2047
rect 390 2047 391 2048
rect 395 2047 396 2051
rect 390 2046 396 2047
rect 398 2051 409 2052
rect 398 2047 399 2051
rect 403 2047 404 2051
rect 408 2047 409 2051
rect 398 2046 409 2047
rect 462 2051 473 2052
rect 462 2047 463 2051
rect 467 2047 468 2051
rect 472 2047 473 2051
rect 462 2046 473 2047
rect 534 2051 545 2052
rect 534 2047 535 2051
rect 539 2047 540 2051
rect 544 2047 545 2051
rect 534 2046 545 2047
rect 614 2051 625 2052
rect 614 2047 615 2051
rect 619 2047 620 2051
rect 624 2047 625 2051
rect 614 2046 625 2047
rect 699 2051 705 2052
rect 699 2047 700 2051
rect 704 2050 705 2051
rect 735 2051 741 2052
rect 735 2050 736 2051
rect 704 2048 736 2050
rect 704 2047 705 2048
rect 699 2046 705 2047
rect 735 2047 736 2048
rect 740 2047 741 2051
rect 735 2046 741 2047
rect 774 2051 785 2052
rect 774 2047 775 2051
rect 779 2047 780 2051
rect 784 2047 785 2051
rect 774 2046 785 2047
rect 859 2051 865 2052
rect 859 2047 860 2051
rect 864 2050 865 2051
rect 895 2051 901 2052
rect 895 2050 896 2051
rect 864 2048 896 2050
rect 864 2047 865 2048
rect 859 2046 865 2047
rect 895 2047 896 2048
rect 900 2047 901 2051
rect 895 2046 901 2047
rect 947 2051 953 2052
rect 947 2047 948 2051
rect 952 2050 953 2051
rect 983 2051 989 2052
rect 983 2050 984 2051
rect 952 2048 984 2050
rect 952 2047 953 2048
rect 947 2046 953 2047
rect 983 2047 984 2048
rect 988 2047 989 2051
rect 983 2046 989 2047
rect 1030 2051 1041 2052
rect 1030 2047 1031 2051
rect 1035 2047 1036 2051
rect 1040 2047 1041 2051
rect 1178 2051 1189 2052
rect 1030 2046 1041 2047
rect 1134 2048 1140 2049
rect 1134 2044 1135 2048
rect 1139 2044 1140 2048
rect 1178 2047 1179 2051
rect 1183 2047 1184 2051
rect 1188 2047 1189 2051
rect 1178 2046 1189 2047
rect 1191 2051 1197 2052
rect 1191 2047 1192 2051
rect 1196 2050 1197 2051
rect 1239 2051 1245 2052
rect 1239 2050 1240 2051
rect 1196 2048 1240 2050
rect 1196 2047 1197 2048
rect 1191 2046 1197 2047
rect 1239 2047 1240 2048
rect 1244 2047 1245 2051
rect 1239 2046 1245 2047
rect 1247 2051 1253 2052
rect 1247 2047 1248 2051
rect 1252 2050 1253 2051
rect 1327 2051 1333 2052
rect 1327 2050 1328 2051
rect 1252 2048 1328 2050
rect 1252 2047 1253 2048
rect 1247 2046 1253 2047
rect 1327 2047 1328 2048
rect 1332 2047 1333 2051
rect 1327 2046 1333 2047
rect 1358 2051 1364 2052
rect 1358 2047 1359 2051
rect 1363 2050 1364 2051
rect 1423 2051 1429 2052
rect 1423 2050 1424 2051
rect 1363 2048 1424 2050
rect 1363 2047 1364 2048
rect 1358 2046 1364 2047
rect 1423 2047 1424 2048
rect 1428 2047 1429 2051
rect 1423 2046 1429 2047
rect 1431 2051 1437 2052
rect 1431 2047 1432 2051
rect 1436 2050 1437 2051
rect 1519 2051 1525 2052
rect 1519 2050 1520 2051
rect 1436 2048 1520 2050
rect 1436 2047 1437 2048
rect 1431 2046 1437 2047
rect 1519 2047 1520 2048
rect 1524 2047 1525 2051
rect 1519 2046 1525 2047
rect 1614 2051 1621 2052
rect 1614 2047 1615 2051
rect 1620 2047 1621 2051
rect 1614 2046 1621 2047
rect 1646 2051 1652 2052
rect 1646 2047 1647 2051
rect 1651 2050 1652 2051
rect 1703 2051 1709 2052
rect 1703 2050 1704 2051
rect 1651 2048 1704 2050
rect 1651 2047 1652 2048
rect 1646 2046 1652 2047
rect 1703 2047 1704 2048
rect 1708 2047 1709 2051
rect 1703 2046 1709 2047
rect 1750 2051 1756 2052
rect 1750 2047 1751 2051
rect 1755 2050 1756 2051
rect 1783 2051 1789 2052
rect 1783 2050 1784 2051
rect 1755 2048 1784 2050
rect 1755 2047 1756 2048
rect 1750 2046 1756 2047
rect 1783 2047 1784 2048
rect 1788 2047 1789 2051
rect 1783 2046 1789 2047
rect 1791 2051 1797 2052
rect 1791 2047 1792 2051
rect 1796 2050 1797 2051
rect 1855 2051 1861 2052
rect 1855 2050 1856 2051
rect 1796 2048 1856 2050
rect 1796 2047 1797 2048
rect 1791 2046 1797 2047
rect 1855 2047 1856 2048
rect 1860 2047 1861 2051
rect 1855 2046 1861 2047
rect 1863 2051 1869 2052
rect 1863 2047 1864 2051
rect 1868 2050 1869 2051
rect 1919 2051 1925 2052
rect 1919 2050 1920 2051
rect 1868 2048 1920 2050
rect 1868 2047 1869 2048
rect 1863 2046 1869 2047
rect 1919 2047 1920 2048
rect 1924 2047 1925 2051
rect 1919 2046 1925 2047
rect 1982 2051 1989 2052
rect 1982 2047 1983 2051
rect 1988 2047 1989 2051
rect 1982 2046 1989 2047
rect 2047 2051 2053 2052
rect 2047 2047 2048 2051
rect 2052 2050 2053 2051
rect 2062 2051 2068 2052
rect 2062 2050 2063 2051
rect 2052 2048 2063 2050
rect 2052 2047 2053 2048
rect 2047 2046 2053 2047
rect 2062 2047 2063 2048
rect 2067 2047 2068 2051
rect 2062 2046 2068 2047
rect 2078 2051 2084 2052
rect 2078 2047 2079 2051
rect 2083 2050 2084 2051
rect 2095 2051 2101 2052
rect 2095 2050 2096 2051
rect 2083 2048 2096 2050
rect 2083 2047 2084 2048
rect 2078 2046 2084 2047
rect 2095 2047 2096 2048
rect 2100 2047 2101 2051
rect 2095 2046 2101 2047
rect 2118 2048 2124 2049
rect 478 2043 484 2044
rect 478 2042 479 2043
rect 319 2040 479 2042
rect 478 2039 479 2040
rect 483 2039 484 2043
rect 630 2043 636 2044
rect 1134 2043 1140 2044
rect 2118 2044 2119 2048
rect 2123 2044 2124 2048
rect 2118 2043 2124 2044
rect 630 2042 631 2043
rect 478 2038 484 2039
rect 540 2040 631 2042
rect 540 2038 542 2040
rect 630 2039 631 2040
rect 635 2039 636 2043
rect 630 2038 636 2039
rect 1158 2040 1164 2041
rect 539 2037 545 2038
rect 179 2035 185 2036
rect 179 2031 180 2035
rect 184 2034 185 2035
rect 254 2035 260 2036
rect 254 2034 255 2035
rect 184 2032 255 2034
rect 184 2031 185 2032
rect 179 2030 185 2031
rect 254 2031 255 2032
rect 259 2031 260 2035
rect 254 2030 260 2031
rect 275 2035 281 2036
rect 275 2031 276 2035
rect 280 2034 281 2035
rect 286 2035 292 2036
rect 286 2034 287 2035
rect 280 2032 287 2034
rect 280 2031 281 2032
rect 275 2030 281 2031
rect 286 2031 287 2032
rect 291 2031 292 2035
rect 286 2030 292 2031
rect 371 2035 377 2036
rect 371 2031 372 2035
rect 376 2034 377 2035
rect 398 2035 404 2036
rect 398 2034 399 2035
rect 376 2032 399 2034
rect 376 2031 377 2032
rect 371 2030 377 2031
rect 398 2031 399 2032
rect 403 2031 404 2035
rect 398 2030 404 2031
rect 459 2035 465 2036
rect 459 2031 460 2035
rect 464 2034 465 2035
rect 530 2035 536 2036
rect 530 2034 531 2035
rect 464 2032 531 2034
rect 464 2031 465 2032
rect 459 2030 465 2031
rect 530 2031 531 2032
rect 535 2031 536 2035
rect 539 2033 540 2037
rect 544 2033 545 2037
rect 1158 2036 1159 2040
rect 1163 2036 1164 2040
rect 539 2032 545 2033
rect 619 2035 625 2036
rect 530 2030 536 2031
rect 619 2031 620 2035
rect 624 2034 625 2035
rect 642 2035 648 2036
rect 642 2034 643 2035
rect 624 2032 643 2034
rect 624 2031 625 2032
rect 619 2030 625 2031
rect 642 2031 643 2032
rect 647 2031 648 2035
rect 642 2030 648 2031
rect 650 2035 656 2036
rect 650 2031 651 2035
rect 655 2034 656 2035
rect 691 2035 697 2036
rect 691 2034 692 2035
rect 655 2032 692 2034
rect 655 2031 656 2032
rect 650 2030 656 2031
rect 691 2031 692 2032
rect 696 2031 697 2035
rect 691 2030 697 2031
rect 722 2035 728 2036
rect 722 2031 723 2035
rect 727 2034 728 2035
rect 755 2035 761 2036
rect 755 2034 756 2035
rect 727 2032 756 2034
rect 727 2031 728 2032
rect 722 2030 728 2031
rect 755 2031 756 2032
rect 760 2031 761 2035
rect 755 2030 761 2031
rect 811 2035 817 2036
rect 811 2031 812 2035
rect 816 2034 817 2035
rect 822 2035 828 2036
rect 822 2034 823 2035
rect 816 2032 823 2034
rect 816 2031 817 2032
rect 811 2030 817 2031
rect 822 2031 823 2032
rect 827 2031 828 2035
rect 822 2030 828 2031
rect 842 2035 848 2036
rect 842 2031 843 2035
rect 847 2034 848 2035
rect 859 2035 865 2036
rect 859 2034 860 2035
rect 847 2032 860 2034
rect 847 2031 848 2032
rect 842 2030 848 2031
rect 859 2031 860 2032
rect 864 2031 865 2035
rect 859 2030 865 2031
rect 890 2035 896 2036
rect 890 2031 891 2035
rect 895 2034 896 2035
rect 907 2035 913 2036
rect 907 2034 908 2035
rect 895 2032 908 2034
rect 895 2031 896 2032
rect 890 2030 896 2031
rect 907 2031 908 2032
rect 912 2031 913 2035
rect 907 2030 913 2031
rect 938 2035 944 2036
rect 938 2031 939 2035
rect 943 2034 944 2035
rect 955 2035 961 2036
rect 955 2034 956 2035
rect 943 2032 956 2034
rect 943 2031 944 2032
rect 938 2030 944 2031
rect 955 2031 956 2032
rect 960 2031 961 2035
rect 955 2030 961 2031
rect 986 2035 992 2036
rect 986 2031 987 2035
rect 991 2034 992 2035
rect 1003 2035 1009 2036
rect 1003 2034 1004 2035
rect 991 2032 1004 2034
rect 991 2031 992 2032
rect 986 2030 992 2031
rect 1003 2031 1004 2032
rect 1008 2031 1009 2035
rect 1003 2030 1009 2031
rect 1030 2035 1036 2036
rect 1030 2031 1031 2035
rect 1035 2034 1036 2035
rect 1043 2035 1049 2036
rect 1158 2035 1164 2036
rect 1214 2040 1220 2041
rect 1214 2036 1215 2040
rect 1219 2036 1220 2040
rect 1214 2035 1220 2036
rect 1302 2040 1308 2041
rect 1302 2036 1303 2040
rect 1307 2036 1308 2040
rect 1302 2035 1308 2036
rect 1398 2040 1404 2041
rect 1398 2036 1399 2040
rect 1403 2036 1404 2040
rect 1398 2035 1404 2036
rect 1494 2040 1500 2041
rect 1494 2036 1495 2040
rect 1499 2036 1500 2040
rect 1494 2035 1500 2036
rect 1590 2040 1596 2041
rect 1590 2036 1591 2040
rect 1595 2036 1596 2040
rect 1590 2035 1596 2036
rect 1678 2040 1684 2041
rect 1678 2036 1679 2040
rect 1683 2036 1684 2040
rect 1678 2035 1684 2036
rect 1758 2040 1764 2041
rect 1758 2036 1759 2040
rect 1763 2036 1764 2040
rect 1758 2035 1764 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1894 2040 1900 2041
rect 1894 2036 1895 2040
rect 1899 2036 1900 2040
rect 1894 2035 1900 2036
rect 1958 2040 1964 2041
rect 1958 2036 1959 2040
rect 1963 2036 1964 2040
rect 1958 2035 1964 2036
rect 2022 2040 2028 2041
rect 2022 2036 2023 2040
rect 2027 2036 2028 2040
rect 2022 2035 2028 2036
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 1043 2034 1044 2035
rect 1035 2032 1044 2034
rect 1035 2031 1036 2032
rect 1030 2030 1036 2031
rect 1043 2031 1044 2032
rect 1048 2031 1049 2035
rect 1043 2030 1049 2031
rect 1155 2027 1161 2028
rect 182 2024 188 2025
rect 182 2020 183 2024
rect 187 2020 188 2024
rect 182 2019 188 2020
rect 278 2024 284 2025
rect 278 2020 279 2024
rect 283 2020 284 2024
rect 278 2019 284 2020
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 462 2024 468 2025
rect 462 2020 463 2024
rect 467 2020 468 2024
rect 462 2019 468 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 622 2024 628 2025
rect 622 2020 623 2024
rect 627 2020 628 2024
rect 622 2019 628 2020
rect 694 2024 700 2025
rect 694 2020 695 2024
rect 699 2020 700 2024
rect 694 2019 700 2020
rect 758 2024 764 2025
rect 758 2020 759 2024
rect 763 2020 764 2024
rect 758 2019 764 2020
rect 814 2024 820 2025
rect 814 2020 815 2024
rect 819 2020 820 2024
rect 814 2019 820 2020
rect 862 2024 868 2025
rect 862 2020 863 2024
rect 867 2020 868 2024
rect 862 2019 868 2020
rect 910 2024 916 2025
rect 910 2020 911 2024
rect 915 2020 916 2024
rect 910 2019 916 2020
rect 958 2024 964 2025
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 1006 2024 1012 2025
rect 1006 2020 1007 2024
rect 1011 2020 1012 2024
rect 1006 2019 1012 2020
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1155 2023 1156 2027
rect 1160 2026 1161 2027
rect 1191 2027 1197 2028
rect 1191 2026 1192 2027
rect 1160 2024 1192 2026
rect 1160 2023 1161 2024
rect 1155 2022 1161 2023
rect 1191 2023 1192 2024
rect 1196 2023 1197 2027
rect 1191 2022 1197 2023
rect 1211 2027 1217 2028
rect 1211 2023 1212 2027
rect 1216 2026 1217 2027
rect 1247 2027 1253 2028
rect 1247 2026 1248 2027
rect 1216 2024 1248 2026
rect 1216 2023 1217 2024
rect 1211 2022 1217 2023
rect 1247 2023 1248 2024
rect 1252 2023 1253 2027
rect 1247 2022 1253 2023
rect 1266 2027 1272 2028
rect 1266 2023 1267 2027
rect 1271 2026 1272 2027
rect 1299 2027 1305 2028
rect 1299 2026 1300 2027
rect 1271 2024 1300 2026
rect 1271 2023 1272 2024
rect 1266 2022 1272 2023
rect 1299 2023 1300 2024
rect 1304 2023 1305 2027
rect 1299 2022 1305 2023
rect 1395 2027 1401 2028
rect 1395 2023 1396 2027
rect 1400 2026 1401 2027
rect 1431 2027 1437 2028
rect 1431 2026 1432 2027
rect 1400 2024 1432 2026
rect 1400 2023 1401 2024
rect 1395 2022 1401 2023
rect 1431 2023 1432 2024
rect 1436 2023 1437 2027
rect 1431 2022 1437 2023
rect 1486 2027 1497 2028
rect 1486 2023 1487 2027
rect 1491 2023 1492 2027
rect 1496 2023 1497 2027
rect 1486 2022 1497 2023
rect 1587 2027 1593 2028
rect 1587 2023 1588 2027
rect 1592 2026 1593 2027
rect 1646 2027 1652 2028
rect 1646 2026 1647 2027
rect 1592 2024 1647 2026
rect 1592 2023 1593 2024
rect 1587 2022 1593 2023
rect 1646 2023 1647 2024
rect 1651 2023 1652 2027
rect 1646 2022 1652 2023
rect 1670 2027 1681 2028
rect 1670 2023 1671 2027
rect 1675 2023 1676 2027
rect 1680 2023 1681 2027
rect 1670 2022 1681 2023
rect 1755 2027 1761 2028
rect 1755 2023 1756 2027
rect 1760 2026 1761 2027
rect 1791 2027 1797 2028
rect 1791 2026 1792 2027
rect 1760 2024 1792 2026
rect 1760 2023 1761 2024
rect 1755 2022 1761 2023
rect 1791 2023 1792 2024
rect 1796 2023 1797 2027
rect 1791 2022 1797 2023
rect 1827 2027 1833 2028
rect 1827 2023 1828 2027
rect 1832 2026 1833 2027
rect 1863 2027 1869 2028
rect 1863 2026 1864 2027
rect 1832 2024 1864 2026
rect 1832 2023 1833 2024
rect 1827 2022 1833 2023
rect 1863 2023 1864 2024
rect 1868 2023 1869 2027
rect 1863 2022 1869 2023
rect 1891 2027 1897 2028
rect 1891 2023 1892 2027
rect 1896 2026 1897 2027
rect 1902 2027 1908 2028
rect 1902 2026 1903 2027
rect 1896 2024 1903 2026
rect 1896 2023 1897 2024
rect 1891 2022 1897 2023
rect 1902 2023 1903 2024
rect 1907 2023 1908 2027
rect 1902 2022 1908 2023
rect 1955 2027 1961 2028
rect 1955 2023 1956 2027
rect 1960 2026 1961 2027
rect 2007 2027 2013 2028
rect 2007 2026 2008 2027
rect 1960 2024 2008 2026
rect 1960 2023 1961 2024
rect 1955 2022 1961 2023
rect 2007 2023 2008 2024
rect 2012 2023 2013 2027
rect 2007 2022 2013 2023
rect 2019 2027 2025 2028
rect 2019 2023 2020 2027
rect 2024 2026 2025 2027
rect 2054 2027 2060 2028
rect 2054 2026 2055 2027
rect 2024 2024 2055 2026
rect 2024 2023 2025 2024
rect 2019 2022 2025 2023
rect 2054 2023 2055 2024
rect 2059 2023 2060 2027
rect 2054 2022 2060 2023
rect 2062 2027 2073 2028
rect 2062 2023 2063 2027
rect 2067 2023 2068 2027
rect 2072 2023 2073 2027
rect 2062 2022 2073 2023
rect 1046 2019 1052 2020
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 1155 2015 1161 2016
rect 1155 2014 1156 2015
rect 110 2011 116 2012
rect 166 2011 172 2012
rect 166 2007 167 2011
rect 171 2010 172 2011
rect 207 2011 213 2012
rect 207 2010 208 2011
rect 171 2008 208 2010
rect 171 2007 172 2008
rect 166 2006 172 2007
rect 207 2007 208 2008
rect 212 2007 213 2011
rect 207 2006 213 2007
rect 254 2011 260 2012
rect 254 2007 255 2011
rect 259 2010 260 2011
rect 303 2011 309 2012
rect 303 2010 304 2011
rect 259 2008 304 2010
rect 259 2007 260 2008
rect 254 2006 260 2007
rect 303 2007 304 2008
rect 308 2007 309 2011
rect 303 2006 309 2007
rect 390 2011 396 2012
rect 390 2007 391 2011
rect 395 2010 396 2011
rect 399 2011 405 2012
rect 399 2010 400 2011
rect 395 2008 400 2010
rect 395 2007 396 2008
rect 390 2006 396 2007
rect 399 2007 400 2008
rect 404 2007 405 2011
rect 399 2006 405 2007
rect 454 2011 460 2012
rect 454 2007 455 2011
rect 459 2010 460 2011
rect 487 2011 493 2012
rect 487 2010 488 2011
rect 459 2008 488 2010
rect 459 2007 460 2008
rect 454 2006 460 2007
rect 487 2007 488 2008
rect 492 2007 493 2011
rect 487 2006 493 2007
rect 530 2011 536 2012
rect 530 2007 531 2011
rect 535 2010 536 2011
rect 567 2011 573 2012
rect 567 2010 568 2011
rect 535 2008 568 2010
rect 535 2007 536 2008
rect 530 2006 536 2007
rect 567 2007 568 2008
rect 572 2007 573 2011
rect 567 2006 573 2007
rect 647 2011 656 2012
rect 647 2007 648 2011
rect 655 2007 656 2011
rect 647 2006 656 2007
rect 719 2011 728 2012
rect 719 2007 720 2011
rect 727 2007 728 2011
rect 719 2006 728 2007
rect 774 2011 780 2012
rect 774 2007 775 2011
rect 779 2010 780 2011
rect 783 2011 789 2012
rect 783 2010 784 2011
rect 779 2008 784 2010
rect 779 2007 780 2008
rect 774 2006 780 2007
rect 783 2007 784 2008
rect 788 2007 789 2011
rect 783 2006 789 2007
rect 839 2011 848 2012
rect 839 2007 840 2011
rect 847 2007 848 2011
rect 839 2006 848 2007
rect 887 2011 896 2012
rect 887 2007 888 2011
rect 895 2007 896 2011
rect 887 2006 896 2007
rect 935 2011 944 2012
rect 935 2007 936 2011
rect 943 2007 944 2011
rect 935 2006 944 2007
rect 983 2011 992 2012
rect 983 2007 984 2011
rect 991 2007 992 2011
rect 983 2006 992 2007
rect 1030 2011 1037 2012
rect 1030 2007 1031 2011
rect 1036 2007 1037 2011
rect 1030 2006 1037 2007
rect 1071 2011 1077 2012
rect 1094 2011 1100 2012
rect 1116 2012 1156 2014
rect 1071 2007 1072 2011
rect 1076 2010 1077 2011
rect 1076 2008 1090 2010
rect 1076 2007 1077 2008
rect 1071 2006 1077 2007
rect 1088 2006 1090 2008
rect 1116 2006 1118 2012
rect 1155 2011 1156 2012
rect 1160 2011 1161 2015
rect 1155 2010 1161 2011
rect 1186 2015 1192 2016
rect 1186 2011 1187 2015
rect 1191 2014 1192 2015
rect 1235 2015 1241 2016
rect 1235 2014 1236 2015
rect 1191 2012 1236 2014
rect 1191 2011 1192 2012
rect 1186 2010 1192 2011
rect 1235 2011 1236 2012
rect 1240 2011 1241 2015
rect 1235 2010 1241 2011
rect 1347 2015 1353 2016
rect 1347 2011 1348 2015
rect 1352 2014 1353 2015
rect 1358 2015 1364 2016
rect 1358 2014 1359 2015
rect 1352 2012 1359 2014
rect 1352 2011 1353 2012
rect 1347 2010 1353 2011
rect 1358 2011 1359 2012
rect 1363 2011 1364 2015
rect 1358 2010 1364 2011
rect 1378 2015 1384 2016
rect 1378 2011 1379 2015
rect 1383 2014 1384 2015
rect 1451 2015 1457 2016
rect 1451 2014 1452 2015
rect 1383 2012 1452 2014
rect 1383 2011 1384 2012
rect 1378 2010 1384 2011
rect 1451 2011 1452 2012
rect 1456 2011 1457 2015
rect 1451 2010 1457 2011
rect 1487 2015 1493 2016
rect 1487 2011 1488 2015
rect 1492 2014 1493 2015
rect 1555 2015 1561 2016
rect 1555 2014 1556 2015
rect 1492 2012 1556 2014
rect 1492 2011 1493 2012
rect 1487 2010 1493 2011
rect 1555 2011 1556 2012
rect 1560 2011 1561 2015
rect 1555 2010 1561 2011
rect 1646 2015 1657 2016
rect 1646 2011 1647 2015
rect 1651 2011 1652 2015
rect 1656 2011 1657 2015
rect 1646 2010 1657 2011
rect 1739 2015 1745 2016
rect 1739 2011 1740 2015
rect 1744 2014 1745 2015
rect 1750 2015 1756 2016
rect 1750 2014 1751 2015
rect 1744 2012 1751 2014
rect 1744 2011 1745 2012
rect 1739 2010 1745 2011
rect 1750 2011 1751 2012
rect 1755 2011 1756 2015
rect 1750 2010 1756 2011
rect 1770 2015 1776 2016
rect 1770 2011 1771 2015
rect 1775 2014 1776 2015
rect 1819 2015 1825 2016
rect 1819 2014 1820 2015
rect 1775 2012 1820 2014
rect 1775 2011 1776 2012
rect 1770 2010 1776 2011
rect 1819 2011 1820 2012
rect 1824 2011 1825 2015
rect 1819 2010 1825 2011
rect 1850 2015 1856 2016
rect 1850 2011 1851 2015
rect 1855 2014 1856 2015
rect 1891 2015 1897 2016
rect 1891 2014 1892 2015
rect 1855 2012 1892 2014
rect 1855 2011 1856 2012
rect 1850 2010 1856 2011
rect 1891 2011 1892 2012
rect 1896 2011 1897 2015
rect 1891 2010 1897 2011
rect 1938 2015 1944 2016
rect 1938 2011 1939 2015
rect 1943 2014 1944 2015
rect 1955 2015 1961 2016
rect 1955 2014 1956 2015
rect 1943 2012 1956 2014
rect 1943 2011 1944 2012
rect 1938 2010 1944 2011
rect 1955 2011 1956 2012
rect 1960 2011 1961 2015
rect 1955 2010 1961 2011
rect 1986 2015 1992 2016
rect 1986 2011 1987 2015
rect 1991 2014 1992 2015
rect 2019 2015 2025 2016
rect 2019 2014 2020 2015
rect 1991 2012 2020 2014
rect 1991 2011 1992 2012
rect 1986 2010 1992 2011
rect 2019 2011 2020 2012
rect 2024 2011 2025 2015
rect 2019 2010 2025 2011
rect 2067 2015 2073 2016
rect 2067 2011 2068 2015
rect 2072 2014 2073 2015
rect 2078 2015 2084 2016
rect 2078 2014 2079 2015
rect 2072 2012 2079 2014
rect 2072 2011 2073 2012
rect 2067 2010 2073 2011
rect 2078 2011 2079 2012
rect 2083 2011 2084 2015
rect 2078 2010 2084 2011
rect 1088 2004 1118 2006
rect 1158 2004 1164 2005
rect 1158 2000 1159 2004
rect 1163 2000 1164 2004
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1094 1999 1100 2000
rect 1158 1999 1164 2000
rect 1238 2004 1244 2005
rect 1238 2000 1239 2004
rect 1243 2000 1244 2004
rect 1238 1999 1244 2000
rect 1350 2004 1356 2005
rect 1350 2000 1351 2004
rect 1355 2000 1356 2004
rect 1350 1999 1356 2000
rect 1454 2004 1460 2005
rect 1454 2000 1455 2004
rect 1459 2000 1460 2004
rect 1454 1999 1460 2000
rect 1558 2004 1564 2005
rect 1558 2000 1559 2004
rect 1563 2000 1564 2004
rect 1558 1999 1564 2000
rect 1654 2004 1660 2005
rect 1654 2000 1655 2004
rect 1659 2000 1660 2004
rect 1654 1999 1660 2000
rect 1742 2004 1748 2005
rect 1742 2000 1743 2004
rect 1747 2000 1748 2004
rect 1742 1999 1748 2000
rect 1822 2004 1828 2005
rect 1822 2000 1823 2004
rect 1827 2000 1828 2004
rect 1822 1999 1828 2000
rect 1894 2004 1900 2005
rect 1894 2000 1895 2004
rect 1899 2000 1900 2004
rect 1894 1999 1900 2000
rect 1958 2004 1964 2005
rect 1958 2000 1959 2004
rect 1963 2000 1964 2004
rect 1958 1999 1964 2000
rect 2022 2004 2028 2005
rect 2022 2000 2023 2004
rect 2027 2000 2028 2004
rect 2022 1999 2028 2000
rect 2070 2004 2076 2005
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 110 1994 116 1995
rect 182 1996 188 1997
rect 182 1992 183 1996
rect 187 1992 188 1996
rect 182 1991 188 1992
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 374 1996 380 1997
rect 374 1992 375 1996
rect 379 1992 380 1996
rect 374 1991 380 1992
rect 462 1996 468 1997
rect 462 1992 463 1996
rect 467 1992 468 1996
rect 462 1991 468 1992
rect 542 1996 548 1997
rect 542 1992 543 1996
rect 547 1992 548 1996
rect 542 1991 548 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 694 1996 700 1997
rect 694 1992 695 1996
rect 699 1992 700 1996
rect 694 1991 700 1992
rect 758 1996 764 1997
rect 758 1992 759 1996
rect 763 1992 764 1996
rect 758 1991 764 1992
rect 814 1996 820 1997
rect 814 1992 815 1996
rect 819 1992 820 1996
rect 814 1991 820 1992
rect 862 1996 868 1997
rect 862 1992 863 1996
rect 867 1992 868 1996
rect 862 1991 868 1992
rect 910 1996 916 1997
rect 910 1992 911 1996
rect 915 1992 916 1996
rect 910 1991 916 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1006 1996 1012 1997
rect 1006 1992 1007 1996
rect 1011 1992 1012 1996
rect 1006 1991 1012 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1094 1995 1095 1999
rect 1099 1995 1100 1999
rect 1094 1994 1100 1995
rect 1134 1996 1140 1997
rect 1046 1991 1052 1992
rect 1134 1992 1135 1996
rect 1139 1992 1140 1996
rect 2118 1996 2124 1997
rect 2118 1992 2119 1996
rect 2123 1992 2124 1996
rect 1134 1991 1140 1992
rect 1183 1991 1192 1992
rect 1183 1987 1184 1991
rect 1191 1987 1192 1991
rect 1183 1986 1192 1987
rect 1263 1991 1272 1992
rect 1263 1987 1264 1991
rect 1271 1987 1272 1991
rect 1263 1986 1272 1987
rect 1375 1991 1384 1992
rect 1375 1987 1376 1991
rect 1383 1987 1384 1991
rect 1375 1986 1384 1987
rect 1479 1991 1485 1992
rect 1479 1987 1480 1991
rect 1484 1990 1485 1991
rect 1487 1991 1493 1992
rect 1487 1990 1488 1991
rect 1484 1988 1488 1990
rect 1484 1987 1485 1988
rect 1479 1986 1485 1987
rect 1487 1987 1488 1988
rect 1492 1987 1493 1991
rect 1487 1986 1493 1987
rect 1566 1991 1572 1992
rect 1566 1987 1567 1991
rect 1571 1990 1572 1991
rect 1583 1991 1589 1992
rect 1583 1990 1584 1991
rect 1571 1988 1584 1990
rect 1571 1987 1572 1988
rect 1566 1986 1572 1987
rect 1583 1987 1584 1988
rect 1588 1987 1589 1991
rect 1583 1986 1589 1987
rect 1670 1991 1676 1992
rect 1670 1987 1671 1991
rect 1675 1990 1676 1991
rect 1679 1991 1685 1992
rect 1679 1990 1680 1991
rect 1675 1988 1680 1990
rect 1675 1987 1676 1988
rect 1670 1986 1676 1987
rect 1679 1987 1680 1988
rect 1684 1987 1685 1991
rect 1679 1986 1685 1987
rect 1767 1991 1776 1992
rect 1767 1987 1768 1991
rect 1775 1987 1776 1991
rect 1767 1986 1776 1987
rect 1847 1991 1856 1992
rect 1847 1987 1848 1991
rect 1855 1987 1856 1991
rect 1847 1986 1856 1987
rect 1919 1991 1925 1992
rect 1919 1987 1920 1991
rect 1924 1990 1925 1991
rect 1938 1991 1944 1992
rect 1938 1990 1939 1991
rect 1924 1988 1939 1990
rect 1924 1987 1925 1988
rect 1919 1986 1925 1987
rect 1938 1987 1939 1988
rect 1943 1987 1944 1991
rect 1938 1986 1944 1987
rect 1983 1991 1992 1992
rect 1983 1987 1984 1991
rect 1991 1987 1992 1991
rect 1983 1986 1992 1987
rect 2007 1991 2013 1992
rect 2007 1987 2008 1991
rect 2012 1990 2013 1991
rect 2047 1991 2053 1992
rect 2047 1990 2048 1991
rect 2012 1988 2048 1990
rect 2012 1987 2013 1988
rect 2007 1986 2013 1987
rect 2047 1987 2048 1988
rect 2052 1987 2053 1991
rect 2047 1986 2053 1987
rect 2058 1991 2064 1992
rect 2058 1987 2059 1991
rect 2063 1990 2064 1991
rect 2095 1991 2101 1992
rect 2118 1991 2124 1992
rect 2095 1990 2096 1991
rect 2063 1988 2096 1990
rect 2063 1987 2064 1988
rect 2058 1986 2064 1987
rect 2095 1987 2096 1988
rect 2100 1987 2101 1991
rect 2095 1986 2101 1987
rect 158 1984 164 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 158 1980 159 1984
rect 163 1980 164 1984
rect 158 1979 164 1980
rect 230 1984 236 1985
rect 230 1980 231 1984
rect 235 1980 236 1984
rect 230 1979 236 1980
rect 302 1984 308 1985
rect 302 1980 303 1984
rect 307 1980 308 1984
rect 302 1979 308 1980
rect 374 1984 380 1985
rect 374 1980 375 1984
rect 379 1980 380 1984
rect 374 1979 380 1980
rect 446 1984 452 1985
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 526 1984 532 1985
rect 526 1980 527 1984
rect 531 1980 532 1984
rect 526 1979 532 1980
rect 606 1984 612 1985
rect 606 1980 607 1984
rect 611 1980 612 1984
rect 606 1979 612 1980
rect 686 1984 692 1985
rect 686 1980 687 1984
rect 691 1980 692 1984
rect 686 1979 692 1980
rect 758 1984 764 1985
rect 758 1980 759 1984
rect 763 1980 764 1984
rect 758 1979 764 1980
rect 830 1984 836 1985
rect 830 1980 831 1984
rect 835 1980 836 1984
rect 830 1979 836 1980
rect 910 1984 916 1985
rect 910 1980 911 1984
rect 915 1980 916 1984
rect 910 1979 916 1980
rect 990 1984 996 1985
rect 990 1980 991 1984
rect 995 1980 996 1984
rect 990 1979 996 1980
rect 1094 1981 1100 1982
rect 110 1976 116 1977
rect 1094 1977 1095 1981
rect 1099 1977 1100 1981
rect 1094 1976 1100 1977
rect 1134 1979 1140 1980
rect 642 1975 648 1976
rect 642 1971 643 1975
rect 647 1974 648 1975
rect 858 1975 864 1976
rect 647 1972 734 1974
rect 647 1971 648 1972
rect 642 1970 648 1971
rect 182 1967 189 1968
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 182 1963 183 1967
rect 188 1963 189 1967
rect 182 1962 189 1963
rect 255 1967 261 1968
rect 255 1963 256 1967
rect 260 1966 261 1967
rect 294 1967 300 1968
rect 294 1966 295 1967
rect 260 1964 295 1966
rect 260 1963 261 1964
rect 255 1962 261 1963
rect 294 1963 295 1964
rect 299 1963 300 1967
rect 294 1962 300 1963
rect 327 1967 333 1968
rect 327 1963 328 1967
rect 332 1966 333 1967
rect 366 1967 372 1968
rect 366 1966 367 1967
rect 332 1964 367 1966
rect 332 1963 333 1964
rect 327 1962 333 1963
rect 366 1963 367 1964
rect 371 1963 372 1967
rect 366 1962 372 1963
rect 398 1967 405 1968
rect 398 1963 399 1967
rect 404 1963 405 1967
rect 398 1962 405 1963
rect 471 1967 477 1968
rect 471 1963 472 1967
rect 476 1966 477 1967
rect 518 1967 524 1968
rect 518 1966 519 1967
rect 476 1964 519 1966
rect 476 1963 477 1964
rect 471 1962 477 1963
rect 518 1963 519 1964
rect 523 1963 524 1967
rect 518 1962 524 1963
rect 551 1967 557 1968
rect 551 1963 552 1967
rect 556 1966 557 1967
rect 598 1967 604 1968
rect 598 1966 599 1967
rect 556 1964 599 1966
rect 556 1963 557 1964
rect 551 1962 557 1963
rect 598 1963 599 1964
rect 603 1963 604 1967
rect 598 1962 604 1963
rect 631 1967 637 1968
rect 631 1963 632 1967
rect 636 1966 637 1967
rect 678 1967 684 1968
rect 678 1966 679 1967
rect 636 1964 679 1966
rect 636 1963 637 1964
rect 631 1962 637 1963
rect 678 1963 679 1964
rect 683 1963 684 1967
rect 678 1962 684 1963
rect 710 1967 717 1968
rect 710 1963 711 1967
rect 716 1963 717 1967
rect 732 1966 734 1972
rect 858 1971 859 1975
rect 863 1974 864 1975
rect 1134 1975 1135 1979
rect 1139 1975 1140 1979
rect 2118 1979 2124 1980
rect 1134 1974 1140 1975
rect 1158 1976 1164 1977
rect 863 1972 994 1974
rect 863 1971 864 1972
rect 858 1970 864 1971
rect 783 1967 789 1968
rect 783 1966 784 1967
rect 732 1964 784 1966
rect 710 1962 717 1963
rect 783 1963 784 1964
rect 788 1963 789 1967
rect 783 1962 789 1963
rect 791 1967 797 1968
rect 791 1963 792 1967
rect 796 1966 797 1967
rect 855 1967 861 1968
rect 855 1966 856 1967
rect 796 1964 856 1966
rect 796 1963 797 1964
rect 791 1962 797 1963
rect 855 1963 856 1964
rect 860 1963 861 1967
rect 855 1962 861 1963
rect 935 1967 941 1968
rect 935 1963 936 1967
rect 940 1966 941 1967
rect 982 1967 988 1968
rect 982 1966 983 1967
rect 940 1964 983 1966
rect 940 1963 941 1964
rect 935 1962 941 1963
rect 982 1963 983 1964
rect 987 1963 988 1967
rect 992 1966 994 1972
rect 1158 1972 1159 1976
rect 1163 1972 1164 1976
rect 1158 1971 1164 1972
rect 1238 1976 1244 1977
rect 1238 1972 1239 1976
rect 1243 1972 1244 1976
rect 1238 1971 1244 1972
rect 1350 1976 1356 1977
rect 1350 1972 1351 1976
rect 1355 1972 1356 1976
rect 1350 1971 1356 1972
rect 1454 1976 1460 1977
rect 1454 1972 1455 1976
rect 1459 1972 1460 1976
rect 1454 1971 1460 1972
rect 1558 1976 1564 1977
rect 1558 1972 1559 1976
rect 1563 1972 1564 1976
rect 1558 1971 1564 1972
rect 1654 1976 1660 1977
rect 1654 1972 1655 1976
rect 1659 1972 1660 1976
rect 1654 1971 1660 1972
rect 1742 1976 1748 1977
rect 1742 1972 1743 1976
rect 1747 1972 1748 1976
rect 1742 1971 1748 1972
rect 1822 1976 1828 1977
rect 1822 1972 1823 1976
rect 1827 1972 1828 1976
rect 1822 1971 1828 1972
rect 1894 1976 1900 1977
rect 1894 1972 1895 1976
rect 1899 1972 1900 1976
rect 1894 1971 1900 1972
rect 1958 1976 1964 1977
rect 1958 1972 1959 1976
rect 1963 1972 1964 1976
rect 1958 1971 1964 1972
rect 2022 1976 2028 1977
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 2070 1976 2076 1977
rect 2070 1972 2071 1976
rect 2075 1972 2076 1976
rect 2118 1975 2119 1979
rect 2123 1975 2124 1979
rect 2118 1974 2124 1975
rect 2070 1971 2076 1972
rect 1015 1967 1021 1968
rect 1015 1966 1016 1967
rect 992 1964 1016 1966
rect 982 1962 988 1963
rect 1015 1963 1016 1964
rect 1020 1963 1021 1967
rect 1015 1962 1021 1963
rect 1094 1964 1100 1965
rect 110 1959 116 1960
rect 1094 1960 1095 1964
rect 1099 1960 1100 1964
rect 1094 1959 1100 1960
rect 158 1956 164 1957
rect 158 1952 159 1956
rect 163 1952 164 1956
rect 158 1951 164 1952
rect 230 1956 236 1957
rect 230 1952 231 1956
rect 235 1952 236 1956
rect 230 1951 236 1952
rect 302 1956 308 1957
rect 302 1952 303 1956
rect 307 1952 308 1956
rect 302 1951 308 1952
rect 374 1956 380 1957
rect 374 1952 375 1956
rect 379 1952 380 1956
rect 374 1951 380 1952
rect 446 1956 452 1957
rect 446 1952 447 1956
rect 451 1952 452 1956
rect 446 1951 452 1952
rect 526 1956 532 1957
rect 526 1952 527 1956
rect 531 1952 532 1956
rect 526 1951 532 1952
rect 606 1956 612 1957
rect 606 1952 607 1956
rect 611 1952 612 1956
rect 606 1951 612 1952
rect 686 1956 692 1957
rect 686 1952 687 1956
rect 691 1952 692 1956
rect 686 1951 692 1952
rect 758 1956 764 1957
rect 758 1952 759 1956
rect 763 1952 764 1956
rect 758 1951 764 1952
rect 830 1956 836 1957
rect 830 1952 831 1956
rect 835 1952 836 1956
rect 830 1951 836 1952
rect 910 1956 916 1957
rect 910 1952 911 1956
rect 915 1952 916 1956
rect 910 1951 916 1952
rect 990 1956 996 1957
rect 990 1952 991 1956
rect 995 1952 996 1956
rect 990 1951 996 1952
rect 1358 1952 1364 1953
rect 1134 1949 1140 1950
rect 1134 1945 1135 1949
rect 1139 1945 1140 1949
rect 1358 1948 1359 1952
rect 1363 1948 1364 1952
rect 1358 1947 1364 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1486 1952 1492 1953
rect 1486 1948 1487 1952
rect 1491 1948 1492 1952
rect 1486 1947 1492 1948
rect 1558 1952 1564 1953
rect 1558 1948 1559 1952
rect 1563 1948 1564 1952
rect 1558 1947 1564 1948
rect 1630 1952 1636 1953
rect 1630 1948 1631 1952
rect 1635 1948 1636 1952
rect 1630 1947 1636 1948
rect 1702 1952 1708 1953
rect 1702 1948 1703 1952
rect 1707 1948 1708 1952
rect 1702 1947 1708 1948
rect 1774 1952 1780 1953
rect 1774 1948 1775 1952
rect 1779 1948 1780 1952
rect 1774 1947 1780 1948
rect 1846 1952 1852 1953
rect 1846 1948 1847 1952
rect 1851 1948 1852 1952
rect 1846 1947 1852 1948
rect 1926 1952 1932 1953
rect 1926 1948 1927 1952
rect 1931 1948 1932 1952
rect 1926 1947 1932 1948
rect 2006 1952 2012 1953
rect 2006 1948 2007 1952
rect 2011 1948 2012 1952
rect 2006 1947 2012 1948
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2070 1947 2076 1948
rect 2118 1949 2124 1950
rect 1134 1944 1140 1945
rect 2118 1945 2119 1949
rect 2123 1945 2124 1949
rect 2118 1944 2124 1945
rect 155 1943 161 1944
rect 155 1939 156 1943
rect 160 1942 161 1943
rect 166 1943 172 1944
rect 166 1942 167 1943
rect 160 1940 167 1942
rect 160 1939 161 1940
rect 155 1938 161 1939
rect 166 1939 167 1940
rect 171 1939 172 1943
rect 166 1938 172 1939
rect 227 1943 233 1944
rect 227 1939 228 1943
rect 232 1942 233 1943
rect 294 1943 305 1944
rect 232 1940 278 1942
rect 232 1939 233 1940
rect 227 1938 233 1939
rect 198 1935 204 1936
rect 198 1934 199 1935
rect 132 1932 199 1934
rect 132 1930 134 1932
rect 198 1931 199 1932
rect 203 1931 204 1935
rect 276 1934 278 1940
rect 294 1939 295 1943
rect 299 1939 300 1943
rect 304 1939 305 1943
rect 294 1938 305 1939
rect 366 1943 377 1944
rect 366 1939 367 1943
rect 371 1939 372 1943
rect 376 1939 377 1943
rect 366 1938 377 1939
rect 443 1943 449 1944
rect 443 1939 444 1943
rect 448 1942 449 1943
rect 454 1943 460 1944
rect 454 1942 455 1943
rect 448 1940 455 1942
rect 448 1939 449 1940
rect 443 1938 449 1939
rect 454 1939 455 1940
rect 459 1939 460 1943
rect 454 1938 460 1939
rect 518 1943 529 1944
rect 518 1939 519 1943
rect 523 1939 524 1943
rect 528 1939 529 1943
rect 518 1938 529 1939
rect 598 1943 609 1944
rect 598 1939 599 1943
rect 603 1939 604 1943
rect 608 1939 609 1943
rect 598 1938 609 1939
rect 678 1943 689 1944
rect 678 1939 679 1943
rect 683 1939 684 1943
rect 688 1939 689 1943
rect 678 1938 689 1939
rect 755 1943 761 1944
rect 755 1939 756 1943
rect 760 1942 761 1943
rect 791 1943 797 1944
rect 791 1942 792 1943
rect 760 1940 792 1942
rect 760 1939 761 1940
rect 755 1938 761 1939
rect 791 1939 792 1940
rect 796 1939 797 1943
rect 791 1938 797 1939
rect 827 1943 833 1944
rect 827 1939 828 1943
rect 832 1942 833 1943
rect 858 1943 864 1944
rect 858 1942 859 1943
rect 832 1940 859 1942
rect 832 1939 833 1940
rect 827 1938 833 1939
rect 858 1939 859 1940
rect 863 1939 864 1943
rect 858 1938 864 1939
rect 902 1943 913 1944
rect 902 1939 903 1943
rect 907 1939 908 1943
rect 912 1939 913 1943
rect 902 1938 913 1939
rect 982 1943 993 1944
rect 982 1939 983 1943
rect 987 1939 988 1943
rect 992 1939 993 1943
rect 982 1938 993 1939
rect 1382 1943 1388 1944
rect 1382 1939 1383 1943
rect 1387 1942 1388 1943
rect 1387 1940 1458 1942
rect 1387 1939 1388 1940
rect 1382 1938 1388 1939
rect 470 1935 476 1936
rect 470 1934 471 1935
rect 276 1932 471 1934
rect 198 1930 204 1931
rect 470 1931 471 1932
rect 475 1931 476 1935
rect 726 1935 732 1936
rect 726 1934 727 1935
rect 470 1930 476 1931
rect 524 1932 727 1934
rect 524 1930 526 1932
rect 726 1931 727 1932
rect 731 1931 732 1935
rect 1383 1935 1389 1936
rect 726 1930 732 1931
rect 1134 1932 1140 1933
rect 131 1929 137 1930
rect 131 1925 132 1929
rect 136 1925 137 1929
rect 523 1929 529 1930
rect 131 1924 137 1925
rect 171 1927 177 1928
rect 171 1923 172 1927
rect 176 1926 177 1927
rect 182 1927 188 1928
rect 182 1926 183 1927
rect 176 1924 183 1926
rect 176 1923 177 1924
rect 171 1922 177 1923
rect 182 1923 183 1924
rect 187 1923 188 1927
rect 182 1922 188 1923
rect 227 1927 233 1928
rect 227 1923 228 1927
rect 232 1926 233 1927
rect 258 1927 264 1928
rect 232 1924 254 1926
rect 232 1923 233 1924
rect 227 1922 233 1923
rect 252 1918 254 1924
rect 258 1923 259 1927
rect 263 1926 264 1927
rect 291 1927 297 1928
rect 291 1926 292 1927
rect 263 1924 292 1926
rect 263 1923 264 1924
rect 258 1922 264 1923
rect 291 1923 292 1924
rect 296 1923 297 1927
rect 291 1922 297 1923
rect 322 1927 328 1928
rect 322 1923 323 1927
rect 327 1926 328 1927
rect 363 1927 369 1928
rect 363 1926 364 1927
rect 327 1924 364 1926
rect 327 1923 328 1924
rect 322 1922 328 1923
rect 363 1923 364 1924
rect 368 1923 369 1927
rect 363 1922 369 1923
rect 394 1927 400 1928
rect 394 1923 395 1927
rect 399 1926 400 1927
rect 443 1927 449 1928
rect 443 1926 444 1927
rect 399 1924 444 1926
rect 399 1923 400 1924
rect 394 1922 400 1923
rect 443 1923 444 1924
rect 448 1923 449 1927
rect 523 1925 524 1929
rect 528 1925 529 1929
rect 1134 1928 1135 1932
rect 1139 1928 1140 1932
rect 1383 1931 1384 1935
rect 1388 1934 1389 1935
rect 1414 1935 1420 1936
rect 1414 1934 1415 1935
rect 1388 1932 1415 1934
rect 1388 1931 1389 1932
rect 1383 1930 1389 1931
rect 1414 1931 1415 1932
rect 1419 1931 1420 1935
rect 1414 1930 1420 1931
rect 1446 1935 1453 1936
rect 1446 1931 1447 1935
rect 1452 1931 1453 1935
rect 1456 1934 1458 1940
rect 1511 1935 1517 1936
rect 1511 1934 1512 1935
rect 1456 1932 1512 1934
rect 1446 1930 1453 1931
rect 1511 1931 1512 1932
rect 1516 1931 1517 1935
rect 1511 1930 1517 1931
rect 1519 1935 1525 1936
rect 1519 1931 1520 1935
rect 1524 1934 1525 1935
rect 1583 1935 1589 1936
rect 1583 1934 1584 1935
rect 1524 1932 1584 1934
rect 1524 1931 1525 1932
rect 1519 1930 1525 1931
rect 1583 1931 1584 1932
rect 1588 1931 1589 1935
rect 1583 1930 1589 1931
rect 1646 1935 1652 1936
rect 1646 1931 1647 1935
rect 1651 1934 1652 1935
rect 1655 1935 1661 1936
rect 1655 1934 1656 1935
rect 1651 1932 1656 1934
rect 1651 1931 1652 1932
rect 1646 1930 1652 1931
rect 1655 1931 1656 1932
rect 1660 1931 1661 1935
rect 1655 1930 1661 1931
rect 1663 1935 1669 1936
rect 1663 1931 1664 1935
rect 1668 1934 1669 1935
rect 1727 1935 1733 1936
rect 1727 1934 1728 1935
rect 1668 1932 1728 1934
rect 1668 1931 1669 1932
rect 1663 1930 1669 1931
rect 1727 1931 1728 1932
rect 1732 1931 1733 1935
rect 1727 1930 1733 1931
rect 1735 1935 1741 1936
rect 1735 1931 1736 1935
rect 1740 1934 1741 1935
rect 1799 1935 1805 1936
rect 1799 1934 1800 1935
rect 1740 1932 1800 1934
rect 1740 1931 1741 1932
rect 1735 1930 1741 1931
rect 1799 1931 1800 1932
rect 1804 1931 1805 1935
rect 1799 1930 1805 1931
rect 1807 1935 1813 1936
rect 1807 1931 1808 1935
rect 1812 1934 1813 1935
rect 1871 1935 1877 1936
rect 1871 1934 1872 1935
rect 1812 1932 1872 1934
rect 1812 1931 1813 1932
rect 1807 1930 1813 1931
rect 1871 1931 1872 1932
rect 1876 1931 1877 1935
rect 1871 1930 1877 1931
rect 1879 1935 1885 1936
rect 1879 1931 1880 1935
rect 1884 1934 1885 1935
rect 1951 1935 1957 1936
rect 1951 1934 1952 1935
rect 1884 1932 1952 1934
rect 1884 1931 1885 1932
rect 1879 1930 1885 1931
rect 1951 1931 1952 1932
rect 1956 1931 1957 1935
rect 1951 1930 1957 1931
rect 2031 1935 2037 1936
rect 2031 1931 2032 1935
rect 2036 1934 2037 1935
rect 2062 1935 2068 1936
rect 2062 1934 2063 1935
rect 2036 1932 2063 1934
rect 2036 1931 2037 1932
rect 2031 1930 2037 1931
rect 2062 1931 2063 1932
rect 2067 1931 2068 1935
rect 2062 1930 2068 1931
rect 2078 1935 2084 1936
rect 2078 1931 2079 1935
rect 2083 1934 2084 1935
rect 2095 1935 2101 1936
rect 2095 1934 2096 1935
rect 2083 1932 2096 1934
rect 2083 1931 2084 1932
rect 2078 1930 2084 1931
rect 2095 1931 2096 1932
rect 2100 1931 2101 1935
rect 2095 1930 2101 1931
rect 2118 1932 2124 1933
rect 523 1924 529 1925
rect 554 1927 560 1928
rect 443 1922 449 1923
rect 554 1923 555 1927
rect 559 1926 560 1927
rect 611 1927 617 1928
rect 611 1926 612 1927
rect 559 1924 612 1926
rect 559 1923 560 1924
rect 554 1922 560 1923
rect 611 1923 612 1924
rect 616 1923 617 1927
rect 611 1922 617 1923
rect 699 1927 705 1928
rect 699 1923 700 1927
rect 704 1926 705 1927
rect 710 1927 716 1928
rect 710 1926 711 1927
rect 704 1924 711 1926
rect 704 1923 705 1924
rect 699 1922 705 1923
rect 710 1923 711 1924
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 787 1927 793 1928
rect 787 1923 788 1927
rect 792 1926 793 1927
rect 810 1927 816 1928
rect 810 1926 811 1927
rect 792 1924 811 1926
rect 792 1923 793 1924
rect 787 1922 793 1923
rect 810 1923 811 1924
rect 815 1923 816 1927
rect 810 1922 816 1923
rect 818 1927 824 1928
rect 818 1923 819 1927
rect 823 1926 824 1927
rect 875 1927 881 1928
rect 1134 1927 1140 1928
rect 2118 1928 2119 1932
rect 2123 1928 2124 1932
rect 2118 1927 2124 1928
rect 875 1926 876 1927
rect 823 1924 876 1926
rect 823 1923 824 1924
rect 818 1922 824 1923
rect 875 1923 876 1924
rect 880 1923 881 1927
rect 875 1922 881 1923
rect 1358 1924 1364 1925
rect 1358 1920 1359 1924
rect 1363 1920 1364 1924
rect 279 1919 285 1920
rect 1358 1919 1364 1920
rect 1422 1924 1428 1925
rect 1422 1920 1423 1924
rect 1427 1920 1428 1924
rect 1422 1919 1428 1920
rect 1486 1924 1492 1925
rect 1486 1920 1487 1924
rect 1491 1920 1492 1924
rect 1486 1919 1492 1920
rect 1558 1924 1564 1925
rect 1558 1920 1559 1924
rect 1563 1920 1564 1924
rect 1558 1919 1564 1920
rect 1630 1924 1636 1925
rect 1630 1920 1631 1924
rect 1635 1920 1636 1924
rect 1630 1919 1636 1920
rect 1702 1924 1708 1925
rect 1702 1920 1703 1924
rect 1707 1920 1708 1924
rect 1702 1919 1708 1920
rect 1774 1924 1780 1925
rect 1774 1920 1775 1924
rect 1779 1920 1780 1924
rect 1774 1919 1780 1920
rect 1846 1924 1852 1925
rect 1846 1920 1847 1924
rect 1851 1920 1852 1924
rect 1846 1919 1852 1920
rect 1926 1924 1932 1925
rect 1926 1920 1927 1924
rect 1931 1920 1932 1924
rect 1926 1919 1932 1920
rect 2006 1924 2012 1925
rect 2006 1920 2007 1924
rect 2011 1920 2012 1924
rect 2006 1919 2012 1920
rect 2070 1924 2076 1925
rect 2070 1920 2071 1924
rect 2075 1920 2076 1924
rect 2070 1919 2076 1920
rect 279 1918 280 1919
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 174 1916 180 1917
rect 174 1912 175 1916
rect 179 1912 180 1916
rect 174 1911 180 1912
rect 230 1916 236 1917
rect 252 1916 280 1918
rect 230 1912 231 1916
rect 235 1912 236 1916
rect 279 1915 280 1916
rect 284 1915 285 1919
rect 279 1914 285 1915
rect 294 1916 300 1917
rect 230 1911 236 1912
rect 294 1912 295 1916
rect 299 1912 300 1916
rect 294 1911 300 1912
rect 366 1916 372 1917
rect 366 1912 367 1916
rect 371 1912 372 1916
rect 366 1911 372 1912
rect 446 1916 452 1917
rect 446 1912 447 1916
rect 451 1912 452 1916
rect 446 1911 452 1912
rect 526 1916 532 1917
rect 526 1912 527 1916
rect 531 1912 532 1916
rect 526 1911 532 1912
rect 614 1916 620 1917
rect 614 1912 615 1916
rect 619 1912 620 1916
rect 614 1911 620 1912
rect 702 1916 708 1917
rect 702 1912 703 1916
rect 707 1912 708 1916
rect 702 1911 708 1912
rect 790 1916 796 1917
rect 790 1912 791 1916
rect 795 1912 796 1916
rect 790 1911 796 1912
rect 878 1916 884 1917
rect 878 1912 879 1916
rect 883 1912 884 1916
rect 878 1911 884 1912
rect 1355 1911 1361 1912
rect 110 1908 116 1909
rect 110 1904 111 1908
rect 115 1904 116 1908
rect 1094 1908 1100 1909
rect 1094 1904 1095 1908
rect 1099 1904 1100 1908
rect 1342 1907 1348 1908
rect 1342 1906 1343 1907
rect 110 1903 116 1904
rect 159 1903 168 1904
rect 159 1899 160 1903
rect 167 1899 168 1903
rect 159 1898 168 1899
rect 198 1903 205 1904
rect 198 1899 199 1903
rect 204 1899 205 1903
rect 198 1898 205 1899
rect 255 1903 264 1904
rect 255 1899 256 1903
rect 263 1899 264 1903
rect 255 1898 264 1899
rect 319 1903 328 1904
rect 319 1899 320 1903
rect 327 1899 328 1903
rect 319 1898 328 1899
rect 391 1903 400 1904
rect 391 1899 392 1903
rect 399 1899 400 1903
rect 391 1898 400 1899
rect 470 1903 477 1904
rect 470 1899 471 1903
rect 476 1899 477 1903
rect 470 1898 477 1899
rect 551 1903 560 1904
rect 551 1899 552 1903
rect 559 1899 560 1903
rect 551 1898 560 1899
rect 638 1903 645 1904
rect 638 1899 639 1903
rect 644 1899 645 1903
rect 638 1898 645 1899
rect 726 1903 733 1904
rect 726 1899 727 1903
rect 732 1899 733 1903
rect 726 1898 733 1899
rect 815 1903 824 1904
rect 815 1899 816 1903
rect 823 1899 824 1903
rect 815 1898 824 1899
rect 902 1903 909 1904
rect 1094 1903 1100 1904
rect 1228 1904 1343 1906
rect 902 1899 903 1903
rect 908 1899 909 1903
rect 1228 1902 1230 1904
rect 1342 1903 1343 1904
rect 1347 1903 1348 1907
rect 1355 1907 1356 1911
rect 1360 1910 1361 1911
rect 1382 1911 1388 1912
rect 1382 1910 1383 1911
rect 1360 1908 1383 1910
rect 1360 1907 1361 1908
rect 1355 1906 1361 1907
rect 1382 1907 1383 1908
rect 1387 1907 1388 1911
rect 1382 1906 1388 1907
rect 1414 1911 1425 1912
rect 1414 1907 1415 1911
rect 1419 1907 1420 1911
rect 1424 1907 1425 1911
rect 1483 1911 1489 1912
rect 1414 1906 1425 1907
rect 1474 1907 1480 1908
rect 1474 1906 1475 1907
rect 1342 1902 1348 1903
rect 1428 1904 1475 1906
rect 1428 1902 1430 1904
rect 1474 1903 1475 1904
rect 1479 1903 1480 1907
rect 1483 1907 1484 1911
rect 1488 1910 1489 1911
rect 1519 1911 1525 1912
rect 1519 1910 1520 1911
rect 1488 1908 1520 1910
rect 1488 1907 1489 1908
rect 1483 1906 1489 1907
rect 1519 1907 1520 1908
rect 1524 1907 1525 1911
rect 1519 1906 1525 1907
rect 1555 1911 1561 1912
rect 1555 1907 1556 1911
rect 1560 1910 1561 1911
rect 1566 1911 1572 1912
rect 1566 1910 1567 1911
rect 1560 1908 1567 1910
rect 1560 1907 1561 1908
rect 1555 1906 1561 1907
rect 1566 1907 1567 1908
rect 1571 1907 1572 1911
rect 1566 1906 1572 1907
rect 1627 1911 1633 1912
rect 1627 1907 1628 1911
rect 1632 1910 1633 1911
rect 1663 1911 1669 1912
rect 1663 1910 1664 1911
rect 1632 1908 1664 1910
rect 1632 1907 1633 1908
rect 1627 1906 1633 1907
rect 1663 1907 1664 1908
rect 1668 1907 1669 1911
rect 1663 1906 1669 1907
rect 1699 1911 1705 1912
rect 1699 1907 1700 1911
rect 1704 1910 1705 1911
rect 1735 1911 1741 1912
rect 1735 1910 1736 1911
rect 1704 1908 1736 1910
rect 1704 1907 1705 1908
rect 1699 1906 1705 1907
rect 1735 1907 1736 1908
rect 1740 1907 1741 1911
rect 1735 1906 1741 1907
rect 1771 1911 1777 1912
rect 1771 1907 1772 1911
rect 1776 1910 1777 1911
rect 1807 1911 1813 1912
rect 1807 1910 1808 1911
rect 1776 1908 1808 1910
rect 1776 1907 1777 1908
rect 1771 1906 1777 1907
rect 1807 1907 1808 1908
rect 1812 1907 1813 1911
rect 1807 1906 1813 1907
rect 1843 1911 1849 1912
rect 1843 1907 1844 1911
rect 1848 1910 1849 1911
rect 1879 1911 1885 1912
rect 1879 1910 1880 1911
rect 1848 1908 1880 1910
rect 1848 1907 1849 1908
rect 1843 1906 1849 1907
rect 1879 1907 1880 1908
rect 1884 1907 1885 1911
rect 1879 1906 1885 1907
rect 1923 1911 1929 1912
rect 1923 1907 1924 1911
rect 1928 1910 1929 1911
rect 1986 1911 1992 1912
rect 1986 1910 1987 1911
rect 1928 1908 1987 1910
rect 1928 1907 1929 1908
rect 1923 1906 1929 1907
rect 1986 1907 1987 1908
rect 1991 1907 1992 1911
rect 1986 1906 1992 1907
rect 2003 1911 2009 1912
rect 2003 1907 2004 1911
rect 2008 1910 2009 1911
rect 2054 1911 2060 1912
rect 2054 1910 2055 1911
rect 2008 1908 2055 1910
rect 2008 1907 2009 1908
rect 2003 1906 2009 1907
rect 2054 1907 2055 1908
rect 2059 1907 2060 1911
rect 2054 1906 2060 1907
rect 2062 1911 2073 1912
rect 2062 1907 2063 1911
rect 2067 1907 2068 1911
rect 2072 1907 2073 1911
rect 2062 1906 2073 1907
rect 1474 1902 1480 1903
rect 902 1898 909 1899
rect 1227 1901 1233 1902
rect 1227 1897 1228 1901
rect 1232 1897 1233 1901
rect 1371 1901 1430 1902
rect 1227 1896 1233 1897
rect 1258 1899 1264 1900
rect 1258 1895 1259 1899
rect 1263 1898 1264 1899
rect 1267 1899 1273 1900
rect 1267 1898 1268 1899
rect 1263 1896 1268 1898
rect 1263 1895 1264 1896
rect 1258 1894 1264 1895
rect 1267 1895 1268 1896
rect 1272 1895 1273 1899
rect 1267 1894 1273 1895
rect 1315 1899 1321 1900
rect 1315 1895 1316 1899
rect 1320 1898 1321 1899
rect 1359 1899 1365 1900
rect 1359 1898 1360 1899
rect 1320 1896 1360 1898
rect 1320 1895 1321 1896
rect 1315 1894 1321 1895
rect 1359 1895 1360 1896
rect 1364 1895 1365 1899
rect 1371 1897 1372 1901
rect 1376 1900 1430 1901
rect 1376 1897 1377 1900
rect 1371 1896 1377 1897
rect 1435 1899 1441 1900
rect 1359 1894 1365 1895
rect 1435 1895 1436 1899
rect 1440 1898 1441 1899
rect 1446 1899 1452 1900
rect 1446 1898 1447 1899
rect 1440 1896 1447 1898
rect 1440 1895 1441 1896
rect 1435 1894 1441 1895
rect 1446 1895 1447 1896
rect 1451 1895 1452 1899
rect 1446 1894 1452 1895
rect 1466 1899 1472 1900
rect 1466 1895 1467 1899
rect 1471 1898 1472 1899
rect 1499 1899 1505 1900
rect 1499 1898 1500 1899
rect 1471 1896 1500 1898
rect 1471 1895 1472 1896
rect 1466 1894 1472 1895
rect 1499 1895 1500 1896
rect 1504 1895 1505 1899
rect 1499 1894 1505 1895
rect 1566 1899 1577 1900
rect 1566 1895 1567 1899
rect 1571 1895 1572 1899
rect 1576 1895 1577 1899
rect 1566 1894 1577 1895
rect 1602 1899 1608 1900
rect 1602 1895 1603 1899
rect 1607 1898 1608 1899
rect 1651 1899 1657 1900
rect 1651 1898 1652 1899
rect 1607 1896 1652 1898
rect 1607 1895 1608 1896
rect 1602 1894 1608 1895
rect 1651 1895 1652 1896
rect 1656 1895 1657 1899
rect 1651 1894 1657 1895
rect 1682 1899 1688 1900
rect 1682 1895 1683 1899
rect 1687 1898 1688 1899
rect 1747 1899 1753 1900
rect 1747 1898 1748 1899
rect 1687 1896 1748 1898
rect 1687 1895 1688 1896
rect 1682 1894 1688 1895
rect 1747 1895 1748 1896
rect 1752 1895 1753 1899
rect 1859 1899 1865 1900
rect 1859 1898 1860 1899
rect 1776 1896 1860 1898
rect 1747 1894 1753 1895
rect 1774 1895 1780 1896
rect 110 1891 116 1892
rect 110 1887 111 1891
rect 115 1887 116 1891
rect 1094 1891 1100 1892
rect 110 1886 116 1887
rect 134 1888 140 1889
rect 134 1884 135 1888
rect 139 1884 140 1888
rect 134 1883 140 1884
rect 174 1888 180 1889
rect 174 1884 175 1888
rect 179 1884 180 1888
rect 174 1883 180 1884
rect 230 1888 236 1889
rect 230 1884 231 1888
rect 235 1884 236 1888
rect 230 1883 236 1884
rect 294 1888 300 1889
rect 294 1884 295 1888
rect 299 1884 300 1888
rect 294 1883 300 1884
rect 366 1888 372 1889
rect 366 1884 367 1888
rect 371 1884 372 1888
rect 366 1883 372 1884
rect 446 1888 452 1889
rect 446 1884 447 1888
rect 451 1884 452 1888
rect 446 1883 452 1884
rect 526 1888 532 1889
rect 526 1884 527 1888
rect 531 1884 532 1888
rect 526 1883 532 1884
rect 614 1888 620 1889
rect 614 1884 615 1888
rect 619 1884 620 1888
rect 614 1883 620 1884
rect 702 1888 708 1889
rect 702 1884 703 1888
rect 707 1884 708 1888
rect 702 1883 708 1884
rect 790 1888 796 1889
rect 790 1884 791 1888
rect 795 1884 796 1888
rect 790 1883 796 1884
rect 878 1888 884 1889
rect 878 1884 879 1888
rect 883 1884 884 1888
rect 1094 1887 1095 1891
rect 1099 1887 1100 1891
rect 1774 1891 1775 1895
rect 1779 1891 1780 1895
rect 1859 1895 1860 1896
rect 1864 1895 1865 1899
rect 1859 1894 1865 1895
rect 1890 1899 1896 1900
rect 1890 1895 1891 1899
rect 1895 1898 1896 1899
rect 1971 1899 1977 1900
rect 1971 1898 1972 1899
rect 1895 1896 1972 1898
rect 1895 1895 1896 1896
rect 1890 1894 1896 1895
rect 1971 1895 1972 1896
rect 1976 1895 1977 1899
rect 1971 1894 1977 1895
rect 2067 1899 2073 1900
rect 2067 1895 2068 1899
rect 2072 1898 2073 1899
rect 2078 1899 2084 1900
rect 2078 1898 2079 1899
rect 2072 1896 2079 1898
rect 2072 1895 2073 1896
rect 2067 1894 2073 1895
rect 2078 1895 2079 1896
rect 2083 1895 2084 1899
rect 2078 1894 2084 1895
rect 1774 1890 1780 1891
rect 1094 1886 1100 1887
rect 1230 1888 1236 1889
rect 878 1883 884 1884
rect 1230 1884 1231 1888
rect 1235 1884 1236 1888
rect 1230 1883 1236 1884
rect 1270 1888 1276 1889
rect 1270 1884 1271 1888
rect 1275 1884 1276 1888
rect 1270 1883 1276 1884
rect 1318 1888 1324 1889
rect 1318 1884 1319 1888
rect 1323 1884 1324 1888
rect 1318 1883 1324 1884
rect 1374 1888 1380 1889
rect 1374 1884 1375 1888
rect 1379 1884 1380 1888
rect 1374 1883 1380 1884
rect 1438 1888 1444 1889
rect 1438 1884 1439 1888
rect 1443 1884 1444 1888
rect 1438 1883 1444 1884
rect 1502 1888 1508 1889
rect 1502 1884 1503 1888
rect 1507 1884 1508 1888
rect 1502 1883 1508 1884
rect 1574 1888 1580 1889
rect 1574 1884 1575 1888
rect 1579 1884 1580 1888
rect 1574 1883 1580 1884
rect 1654 1888 1660 1889
rect 1654 1884 1655 1888
rect 1659 1884 1660 1888
rect 1654 1883 1660 1884
rect 1750 1888 1756 1889
rect 1750 1884 1751 1888
rect 1755 1884 1756 1888
rect 1750 1883 1756 1884
rect 1862 1888 1868 1889
rect 1862 1884 1863 1888
rect 1867 1884 1868 1888
rect 1862 1883 1868 1884
rect 1974 1888 1980 1889
rect 1974 1884 1975 1888
rect 1979 1884 1980 1888
rect 1974 1883 1980 1884
rect 2070 1888 2076 1889
rect 2070 1884 2071 1888
rect 2075 1884 2076 1888
rect 2070 1883 2076 1884
rect 1134 1880 1140 1881
rect 1134 1876 1135 1880
rect 1139 1876 1140 1880
rect 2118 1880 2124 1881
rect 2118 1876 2119 1880
rect 2123 1876 2124 1880
rect 1134 1875 1140 1876
rect 1255 1875 1264 1876
rect 134 1872 140 1873
rect 110 1869 116 1870
rect 110 1865 111 1869
rect 115 1865 116 1869
rect 134 1868 135 1872
rect 139 1868 140 1872
rect 134 1867 140 1868
rect 174 1872 180 1873
rect 174 1868 175 1872
rect 179 1868 180 1872
rect 174 1867 180 1868
rect 222 1872 228 1873
rect 222 1868 223 1872
rect 227 1868 228 1872
rect 222 1867 228 1868
rect 286 1872 292 1873
rect 286 1868 287 1872
rect 291 1868 292 1872
rect 286 1867 292 1868
rect 358 1872 364 1873
rect 358 1868 359 1872
rect 363 1868 364 1872
rect 358 1867 364 1868
rect 430 1872 436 1873
rect 430 1868 431 1872
rect 435 1868 436 1872
rect 430 1867 436 1868
rect 502 1872 508 1873
rect 502 1868 503 1872
rect 507 1868 508 1872
rect 502 1867 508 1868
rect 566 1872 572 1873
rect 566 1868 567 1872
rect 571 1868 572 1872
rect 566 1867 572 1868
rect 630 1872 636 1873
rect 630 1868 631 1872
rect 635 1868 636 1872
rect 630 1867 636 1868
rect 694 1872 700 1873
rect 694 1868 695 1872
rect 699 1868 700 1872
rect 694 1867 700 1868
rect 758 1872 764 1873
rect 758 1868 759 1872
rect 763 1868 764 1872
rect 758 1867 764 1868
rect 830 1872 836 1873
rect 830 1868 831 1872
rect 835 1868 836 1872
rect 1255 1871 1256 1875
rect 1263 1871 1264 1875
rect 1255 1870 1264 1871
rect 1294 1875 1301 1876
rect 1294 1871 1295 1875
rect 1300 1871 1301 1875
rect 1294 1870 1301 1871
rect 1342 1875 1349 1876
rect 1342 1871 1343 1875
rect 1348 1871 1349 1875
rect 1342 1870 1349 1871
rect 1359 1875 1365 1876
rect 1359 1871 1360 1875
rect 1364 1874 1365 1875
rect 1399 1875 1405 1876
rect 1399 1874 1400 1875
rect 1364 1872 1400 1874
rect 1364 1871 1365 1872
rect 1359 1870 1365 1871
rect 1399 1871 1400 1872
rect 1404 1871 1405 1875
rect 1399 1870 1405 1871
rect 1463 1875 1472 1876
rect 1463 1871 1464 1875
rect 1471 1871 1472 1875
rect 1463 1870 1472 1871
rect 1474 1875 1480 1876
rect 1474 1871 1475 1875
rect 1479 1874 1480 1875
rect 1527 1875 1533 1876
rect 1527 1874 1528 1875
rect 1479 1872 1528 1874
rect 1479 1871 1480 1872
rect 1474 1870 1480 1871
rect 1527 1871 1528 1872
rect 1532 1871 1533 1875
rect 1527 1870 1533 1871
rect 1599 1875 1608 1876
rect 1599 1871 1600 1875
rect 1607 1871 1608 1875
rect 1599 1870 1608 1871
rect 1679 1875 1688 1876
rect 1679 1871 1680 1875
rect 1687 1871 1688 1875
rect 1679 1870 1688 1871
rect 1774 1875 1781 1876
rect 1774 1871 1775 1875
rect 1780 1871 1781 1875
rect 1774 1870 1781 1871
rect 1887 1875 1896 1876
rect 1887 1871 1888 1875
rect 1895 1871 1896 1875
rect 1887 1870 1896 1871
rect 1986 1875 1992 1876
rect 1986 1871 1987 1875
rect 1991 1874 1992 1875
rect 1999 1875 2005 1876
rect 1999 1874 2000 1875
rect 1991 1872 2000 1874
rect 1991 1871 1992 1872
rect 1986 1870 1992 1871
rect 1999 1871 2000 1872
rect 2004 1871 2005 1875
rect 1999 1870 2005 1871
rect 2047 1875 2053 1876
rect 2047 1871 2048 1875
rect 2052 1874 2053 1875
rect 2095 1875 2101 1876
rect 2118 1875 2124 1876
rect 2095 1874 2096 1875
rect 2052 1872 2096 1874
rect 2052 1871 2053 1872
rect 2047 1870 2053 1871
rect 2095 1871 2096 1872
rect 2100 1871 2101 1875
rect 2095 1870 2101 1871
rect 830 1867 836 1868
rect 1094 1869 1100 1870
rect 110 1864 116 1865
rect 1094 1865 1095 1869
rect 1099 1865 1100 1869
rect 1094 1864 1100 1865
rect 310 1863 316 1864
rect 310 1859 311 1863
rect 315 1862 316 1863
rect 526 1863 532 1864
rect 315 1860 434 1862
rect 315 1859 316 1860
rect 310 1858 316 1859
rect 142 1855 148 1856
rect 110 1852 116 1853
rect 110 1848 111 1852
rect 115 1848 116 1852
rect 142 1851 143 1855
rect 147 1854 148 1855
rect 159 1855 165 1856
rect 159 1854 160 1855
rect 147 1852 160 1854
rect 147 1851 148 1852
rect 142 1850 148 1851
rect 159 1851 160 1852
rect 164 1851 165 1855
rect 159 1850 165 1851
rect 199 1855 205 1856
rect 199 1851 200 1855
rect 204 1854 205 1855
rect 214 1855 220 1856
rect 214 1854 215 1855
rect 204 1852 215 1854
rect 204 1851 205 1852
rect 199 1850 205 1851
rect 214 1851 215 1852
rect 219 1851 220 1855
rect 214 1850 220 1851
rect 230 1855 236 1856
rect 230 1851 231 1855
rect 235 1854 236 1855
rect 247 1855 253 1856
rect 247 1854 248 1855
rect 235 1852 248 1854
rect 235 1851 236 1852
rect 230 1850 236 1851
rect 247 1851 248 1852
rect 252 1851 253 1855
rect 247 1850 253 1851
rect 279 1855 285 1856
rect 279 1851 280 1855
rect 284 1854 285 1855
rect 311 1855 317 1856
rect 311 1854 312 1855
rect 284 1852 312 1854
rect 284 1851 285 1852
rect 279 1850 285 1851
rect 311 1851 312 1852
rect 316 1851 317 1855
rect 311 1850 317 1851
rect 383 1855 389 1856
rect 383 1851 384 1855
rect 388 1854 389 1855
rect 422 1855 428 1856
rect 422 1854 423 1855
rect 388 1852 423 1854
rect 388 1851 389 1852
rect 383 1850 389 1851
rect 422 1851 423 1852
rect 427 1851 428 1855
rect 432 1854 434 1860
rect 526 1859 527 1863
rect 531 1862 532 1863
rect 810 1863 816 1864
rect 531 1860 606 1862
rect 531 1859 532 1860
rect 526 1858 532 1859
rect 455 1855 461 1856
rect 455 1854 456 1855
rect 432 1852 456 1854
rect 422 1850 428 1851
rect 455 1851 456 1852
rect 460 1851 461 1855
rect 455 1850 461 1851
rect 527 1855 533 1856
rect 527 1851 528 1855
rect 532 1854 533 1855
rect 558 1855 564 1856
rect 558 1854 559 1855
rect 532 1852 559 1854
rect 532 1851 533 1852
rect 527 1850 533 1851
rect 558 1851 559 1852
rect 563 1851 564 1855
rect 558 1850 564 1851
rect 591 1855 600 1856
rect 591 1851 592 1855
rect 599 1851 600 1855
rect 604 1854 606 1860
rect 810 1859 811 1863
rect 815 1862 816 1863
rect 1134 1863 1140 1864
rect 815 1860 859 1862
rect 815 1859 816 1860
rect 810 1858 816 1859
rect 857 1856 859 1860
rect 1134 1859 1135 1863
rect 1139 1859 1140 1863
rect 2118 1863 2124 1864
rect 1134 1858 1140 1859
rect 1230 1860 1236 1861
rect 1230 1856 1231 1860
rect 1235 1856 1236 1860
rect 655 1855 661 1856
rect 655 1854 656 1855
rect 604 1852 656 1854
rect 591 1850 600 1851
rect 655 1851 656 1852
rect 660 1851 661 1855
rect 655 1850 661 1851
rect 719 1855 725 1856
rect 719 1851 720 1855
rect 724 1854 725 1855
rect 750 1855 756 1856
rect 750 1854 751 1855
rect 724 1852 751 1854
rect 724 1851 725 1852
rect 719 1850 725 1851
rect 750 1851 751 1852
rect 755 1851 756 1855
rect 750 1850 756 1851
rect 783 1855 789 1856
rect 783 1851 784 1855
rect 788 1854 789 1855
rect 822 1855 828 1856
rect 822 1854 823 1855
rect 788 1852 823 1854
rect 788 1851 789 1852
rect 783 1850 789 1851
rect 822 1851 823 1852
rect 827 1851 828 1855
rect 822 1850 828 1851
rect 855 1855 861 1856
rect 1230 1855 1236 1856
rect 1270 1860 1276 1861
rect 1270 1856 1271 1860
rect 1275 1856 1276 1860
rect 1270 1855 1276 1856
rect 1318 1860 1324 1861
rect 1318 1856 1319 1860
rect 1323 1856 1324 1860
rect 1318 1855 1324 1856
rect 1374 1860 1380 1861
rect 1374 1856 1375 1860
rect 1379 1856 1380 1860
rect 1374 1855 1380 1856
rect 1438 1860 1444 1861
rect 1438 1856 1439 1860
rect 1443 1856 1444 1860
rect 1438 1855 1444 1856
rect 1502 1860 1508 1861
rect 1502 1856 1503 1860
rect 1507 1856 1508 1860
rect 1502 1855 1508 1856
rect 1574 1860 1580 1861
rect 1574 1856 1575 1860
rect 1579 1856 1580 1860
rect 1574 1855 1580 1856
rect 1654 1860 1660 1861
rect 1654 1856 1655 1860
rect 1659 1856 1660 1860
rect 1654 1855 1660 1856
rect 1750 1860 1756 1861
rect 1750 1856 1751 1860
rect 1755 1856 1756 1860
rect 1750 1855 1756 1856
rect 1862 1860 1868 1861
rect 1862 1856 1863 1860
rect 1867 1856 1868 1860
rect 1862 1855 1868 1856
rect 1974 1860 1980 1861
rect 1974 1856 1975 1860
rect 1979 1856 1980 1860
rect 1974 1855 1980 1856
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2118 1859 2119 1863
rect 2123 1859 2124 1863
rect 2118 1858 2124 1859
rect 2070 1855 2076 1856
rect 855 1851 856 1855
rect 860 1851 861 1855
rect 855 1850 861 1851
rect 1094 1852 1100 1853
rect 110 1847 116 1848
rect 1094 1848 1095 1852
rect 1099 1848 1100 1852
rect 1094 1847 1100 1848
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 222 1844 228 1845
rect 222 1840 223 1844
rect 227 1840 228 1844
rect 222 1839 228 1840
rect 286 1844 292 1845
rect 286 1840 287 1844
rect 291 1840 292 1844
rect 286 1839 292 1840
rect 358 1844 364 1845
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 430 1844 436 1845
rect 430 1840 431 1844
rect 435 1840 436 1844
rect 430 1839 436 1840
rect 502 1844 508 1845
rect 502 1840 503 1844
rect 507 1840 508 1844
rect 502 1839 508 1840
rect 566 1844 572 1845
rect 566 1840 567 1844
rect 571 1840 572 1844
rect 566 1839 572 1840
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 758 1844 764 1845
rect 758 1840 759 1844
rect 763 1840 764 1844
rect 758 1839 764 1840
rect 830 1844 836 1845
rect 830 1840 831 1844
rect 835 1840 836 1844
rect 1158 1844 1164 1845
rect 830 1839 836 1840
rect 1134 1841 1140 1842
rect 1134 1837 1135 1841
rect 1139 1837 1140 1841
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1238 1844 1244 1845
rect 1238 1840 1239 1844
rect 1243 1840 1244 1844
rect 1238 1839 1244 1840
rect 1302 1844 1308 1845
rect 1302 1840 1303 1844
rect 1307 1840 1308 1844
rect 1302 1839 1308 1840
rect 1366 1844 1372 1845
rect 1366 1840 1367 1844
rect 1371 1840 1372 1844
rect 1366 1839 1372 1840
rect 1430 1844 1436 1845
rect 1430 1840 1431 1844
rect 1435 1840 1436 1844
rect 1430 1839 1436 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1582 1844 1588 1845
rect 1582 1840 1583 1844
rect 1587 1840 1588 1844
rect 1582 1839 1588 1840
rect 1670 1844 1676 1845
rect 1670 1840 1671 1844
rect 1675 1840 1676 1844
rect 1670 1839 1676 1840
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1766 1839 1772 1840
rect 1870 1844 1876 1845
rect 1870 1840 1871 1844
rect 1875 1840 1876 1844
rect 1870 1839 1876 1840
rect 1982 1844 1988 1845
rect 1982 1840 1983 1844
rect 1987 1840 1988 1844
rect 1982 1839 1988 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2070 1839 2076 1840
rect 2118 1841 2124 1842
rect 1134 1836 1140 1837
rect 2118 1837 2119 1841
rect 2123 1837 2124 1841
rect 2118 1836 2124 1837
rect 1566 1835 1572 1836
rect 131 1831 137 1832
rect 131 1827 132 1831
rect 136 1830 137 1831
rect 162 1831 168 1832
rect 136 1828 159 1830
rect 136 1827 137 1828
rect 131 1826 137 1827
rect 157 1822 159 1828
rect 162 1827 163 1831
rect 167 1830 168 1831
rect 171 1831 177 1832
rect 171 1830 172 1831
rect 167 1828 172 1830
rect 167 1827 168 1828
rect 162 1826 168 1827
rect 171 1827 172 1828
rect 176 1827 177 1831
rect 171 1826 177 1827
rect 214 1831 225 1832
rect 214 1827 215 1831
rect 219 1827 220 1831
rect 224 1827 225 1831
rect 214 1826 225 1827
rect 283 1831 289 1832
rect 283 1827 284 1831
rect 288 1830 289 1831
rect 310 1831 316 1832
rect 310 1830 311 1831
rect 288 1828 311 1830
rect 288 1827 289 1828
rect 283 1826 289 1827
rect 310 1827 311 1828
rect 315 1827 316 1831
rect 310 1826 316 1827
rect 355 1831 361 1832
rect 355 1827 356 1831
rect 360 1830 361 1831
rect 374 1831 380 1832
rect 374 1830 375 1831
rect 360 1828 375 1830
rect 360 1827 361 1828
rect 355 1826 361 1827
rect 374 1827 375 1828
rect 379 1827 380 1831
rect 374 1826 380 1827
rect 422 1831 433 1832
rect 422 1827 423 1831
rect 427 1827 428 1831
rect 432 1827 433 1831
rect 422 1826 433 1827
rect 499 1831 505 1832
rect 499 1827 500 1831
rect 504 1830 505 1831
rect 526 1831 532 1832
rect 526 1830 527 1831
rect 504 1828 527 1830
rect 504 1827 505 1828
rect 499 1826 505 1827
rect 526 1827 527 1828
rect 531 1827 532 1831
rect 526 1826 532 1827
rect 558 1831 569 1832
rect 558 1827 559 1831
rect 563 1827 564 1831
rect 568 1827 569 1831
rect 558 1826 569 1827
rect 627 1831 633 1832
rect 627 1827 628 1831
rect 632 1830 633 1831
rect 638 1831 644 1832
rect 638 1830 639 1831
rect 632 1828 639 1830
rect 632 1827 633 1828
rect 627 1826 633 1827
rect 638 1827 639 1828
rect 643 1827 644 1831
rect 638 1826 644 1827
rect 691 1831 697 1832
rect 691 1827 692 1831
rect 696 1830 697 1831
rect 742 1831 748 1832
rect 742 1830 743 1831
rect 696 1828 743 1830
rect 696 1827 697 1828
rect 691 1826 697 1827
rect 742 1827 743 1828
rect 747 1827 748 1831
rect 742 1826 748 1827
rect 750 1831 761 1832
rect 750 1827 751 1831
rect 755 1827 756 1831
rect 760 1827 761 1831
rect 750 1826 761 1827
rect 822 1831 833 1832
rect 822 1827 823 1831
rect 827 1827 828 1831
rect 832 1827 833 1831
rect 1566 1831 1567 1835
rect 1571 1834 1572 1835
rect 1571 1832 1874 1834
rect 1571 1831 1572 1832
rect 1566 1830 1572 1831
rect 822 1826 833 1827
rect 1183 1827 1189 1828
rect 1183 1826 1184 1827
rect 1134 1824 1140 1825
rect 230 1823 236 1824
rect 230 1822 231 1823
rect 157 1820 231 1822
rect 230 1819 231 1820
rect 235 1819 236 1823
rect 462 1823 468 1824
rect 462 1822 463 1823
rect 230 1818 236 1819
rect 260 1820 463 1822
rect 260 1818 262 1820
rect 462 1819 463 1820
rect 467 1819 468 1823
rect 1014 1823 1020 1824
rect 1014 1822 1015 1823
rect 462 1818 468 1819
rect 836 1820 1015 1822
rect 836 1818 838 1820
rect 1014 1819 1015 1820
rect 1019 1819 1020 1823
rect 1134 1820 1135 1824
rect 1139 1820 1140 1824
rect 1134 1819 1140 1820
rect 1144 1824 1184 1826
rect 1014 1818 1020 1819
rect 259 1817 265 1818
rect 131 1815 137 1816
rect 131 1811 132 1815
rect 136 1814 137 1815
rect 142 1815 148 1816
rect 142 1814 143 1815
rect 136 1812 143 1814
rect 136 1811 137 1812
rect 131 1810 137 1811
rect 142 1811 143 1812
rect 147 1811 148 1815
rect 142 1810 148 1811
rect 162 1815 168 1816
rect 162 1811 163 1815
rect 167 1814 168 1815
rect 179 1815 185 1816
rect 179 1814 180 1815
rect 167 1812 180 1814
rect 167 1811 168 1812
rect 162 1810 168 1811
rect 179 1811 180 1812
rect 184 1811 185 1815
rect 259 1813 260 1817
rect 264 1813 265 1817
rect 835 1817 841 1818
rect 259 1812 265 1813
rect 298 1815 304 1816
rect 179 1810 185 1811
rect 298 1811 299 1815
rect 303 1814 304 1815
rect 347 1815 353 1816
rect 347 1814 348 1815
rect 303 1812 348 1814
rect 303 1811 304 1812
rect 298 1810 304 1811
rect 347 1811 348 1812
rect 352 1811 353 1815
rect 347 1810 353 1811
rect 435 1815 441 1816
rect 435 1811 436 1815
rect 440 1814 441 1815
rect 510 1815 516 1816
rect 510 1814 511 1815
rect 440 1812 511 1814
rect 440 1811 441 1812
rect 435 1810 441 1811
rect 510 1811 511 1812
rect 515 1811 516 1815
rect 510 1810 516 1811
rect 518 1815 529 1816
rect 518 1811 519 1815
rect 523 1811 524 1815
rect 528 1811 529 1815
rect 518 1810 529 1811
rect 594 1815 600 1816
rect 594 1811 595 1815
rect 599 1814 600 1815
rect 603 1815 609 1816
rect 603 1814 604 1815
rect 599 1812 604 1814
rect 599 1811 600 1812
rect 594 1810 600 1811
rect 603 1811 604 1812
rect 608 1811 609 1815
rect 603 1810 609 1811
rect 639 1815 645 1816
rect 639 1811 640 1815
rect 644 1814 645 1815
rect 683 1815 689 1816
rect 683 1814 684 1815
rect 644 1812 684 1814
rect 644 1811 645 1812
rect 639 1810 645 1811
rect 683 1811 684 1812
rect 688 1811 689 1815
rect 683 1810 689 1811
rect 714 1815 720 1816
rect 714 1811 715 1815
rect 719 1814 720 1815
rect 763 1815 769 1816
rect 763 1814 764 1815
rect 719 1812 764 1814
rect 719 1811 720 1812
rect 714 1810 720 1811
rect 763 1811 764 1812
rect 768 1811 769 1815
rect 835 1813 836 1817
rect 840 1813 841 1817
rect 835 1812 841 1813
rect 866 1815 872 1816
rect 763 1810 769 1811
rect 866 1811 867 1815
rect 871 1814 872 1815
rect 907 1815 913 1816
rect 907 1814 908 1815
rect 871 1812 908 1814
rect 871 1811 872 1812
rect 866 1810 872 1811
rect 907 1811 908 1812
rect 912 1811 913 1815
rect 907 1810 913 1811
rect 987 1815 993 1816
rect 987 1811 988 1815
rect 992 1814 993 1815
rect 1034 1815 1040 1816
rect 1034 1814 1035 1815
rect 992 1812 1035 1814
rect 992 1811 993 1812
rect 987 1810 993 1811
rect 1034 1811 1035 1812
rect 1039 1811 1040 1815
rect 1034 1810 1040 1811
rect 1043 1815 1049 1816
rect 1043 1811 1044 1815
rect 1048 1814 1049 1815
rect 1144 1814 1146 1824
rect 1183 1823 1184 1824
rect 1188 1823 1189 1827
rect 1223 1827 1229 1828
rect 1223 1826 1224 1827
rect 1183 1822 1189 1823
rect 1192 1824 1224 1826
rect 1048 1812 1146 1814
rect 1158 1816 1164 1817
rect 1158 1812 1159 1816
rect 1163 1812 1164 1816
rect 1048 1811 1049 1812
rect 1158 1811 1164 1812
rect 1043 1810 1049 1811
rect 1192 1810 1194 1824
rect 1223 1823 1224 1824
rect 1228 1823 1229 1827
rect 1263 1827 1269 1828
rect 1263 1826 1264 1827
rect 1223 1822 1229 1823
rect 1232 1824 1264 1826
rect 1198 1816 1204 1817
rect 1198 1812 1199 1816
rect 1203 1812 1204 1816
rect 1232 1814 1234 1824
rect 1263 1823 1264 1824
rect 1268 1823 1269 1827
rect 1263 1822 1269 1823
rect 1327 1827 1333 1828
rect 1327 1823 1328 1827
rect 1332 1826 1333 1827
rect 1358 1827 1364 1828
rect 1358 1826 1359 1827
rect 1332 1824 1359 1826
rect 1332 1823 1333 1824
rect 1327 1822 1333 1823
rect 1358 1823 1359 1824
rect 1363 1823 1364 1827
rect 1358 1822 1364 1823
rect 1374 1827 1380 1828
rect 1374 1823 1375 1827
rect 1379 1826 1380 1827
rect 1391 1827 1397 1828
rect 1391 1826 1392 1827
rect 1379 1824 1392 1826
rect 1379 1823 1380 1824
rect 1374 1822 1380 1823
rect 1391 1823 1392 1824
rect 1396 1823 1397 1827
rect 1391 1822 1397 1823
rect 1455 1827 1461 1828
rect 1455 1823 1456 1827
rect 1460 1826 1461 1827
rect 1494 1827 1500 1828
rect 1494 1826 1495 1827
rect 1460 1824 1495 1826
rect 1460 1823 1461 1824
rect 1455 1822 1461 1823
rect 1494 1823 1495 1824
rect 1499 1823 1500 1827
rect 1494 1822 1500 1823
rect 1527 1827 1533 1828
rect 1527 1823 1528 1827
rect 1532 1826 1533 1827
rect 1574 1827 1580 1828
rect 1574 1826 1575 1827
rect 1532 1824 1575 1826
rect 1532 1823 1533 1824
rect 1527 1822 1533 1823
rect 1574 1823 1575 1824
rect 1579 1823 1580 1827
rect 1574 1822 1580 1823
rect 1607 1827 1613 1828
rect 1607 1823 1608 1827
rect 1612 1826 1613 1827
rect 1662 1827 1668 1828
rect 1662 1826 1663 1827
rect 1612 1824 1663 1826
rect 1612 1823 1613 1824
rect 1607 1822 1613 1823
rect 1662 1823 1663 1824
rect 1667 1823 1668 1827
rect 1662 1822 1668 1823
rect 1695 1827 1701 1828
rect 1695 1823 1696 1827
rect 1700 1826 1701 1827
rect 1758 1827 1764 1828
rect 1758 1826 1759 1827
rect 1700 1824 1759 1826
rect 1700 1823 1701 1824
rect 1695 1822 1701 1823
rect 1758 1823 1759 1824
rect 1763 1823 1764 1827
rect 1758 1822 1764 1823
rect 1791 1827 1797 1828
rect 1791 1823 1792 1827
rect 1796 1826 1797 1827
rect 1862 1827 1868 1828
rect 1862 1826 1863 1827
rect 1796 1824 1863 1826
rect 1796 1823 1797 1824
rect 1791 1822 1797 1823
rect 1862 1823 1863 1824
rect 1867 1823 1868 1827
rect 1872 1826 1874 1832
rect 1895 1827 1901 1828
rect 1895 1826 1896 1827
rect 1872 1824 1896 1826
rect 1862 1822 1868 1823
rect 1895 1823 1896 1824
rect 1900 1823 1901 1827
rect 1895 1822 1901 1823
rect 2007 1827 2013 1828
rect 2007 1823 2008 1827
rect 2012 1826 2013 1827
rect 2062 1827 2068 1828
rect 2062 1826 2063 1827
rect 2012 1824 2063 1826
rect 2012 1823 2013 1824
rect 2007 1822 2013 1823
rect 2062 1823 2063 1824
rect 2067 1823 2068 1827
rect 2062 1822 2068 1823
rect 2078 1827 2084 1828
rect 2078 1823 2079 1827
rect 2083 1826 2084 1827
rect 2095 1827 2101 1828
rect 2095 1826 2096 1827
rect 2083 1824 2096 1826
rect 2083 1823 2084 1824
rect 2078 1822 2084 1823
rect 2095 1823 2096 1824
rect 2100 1823 2101 1827
rect 2095 1822 2101 1823
rect 2118 1824 2124 1825
rect 2118 1820 2119 1824
rect 2123 1820 2124 1824
rect 2118 1819 2124 1820
rect 1198 1811 1204 1812
rect 1208 1812 1234 1814
rect 1238 1816 1244 1817
rect 1238 1812 1239 1816
rect 1243 1812 1244 1816
rect 1188 1808 1194 1810
rect 1188 1806 1190 1808
rect 1208 1806 1210 1812
rect 1238 1811 1244 1812
rect 1302 1816 1308 1817
rect 1302 1812 1303 1816
rect 1307 1812 1308 1816
rect 1302 1811 1308 1812
rect 1366 1816 1372 1817
rect 1366 1812 1367 1816
rect 1371 1812 1372 1816
rect 1366 1811 1372 1812
rect 1430 1816 1436 1817
rect 1430 1812 1431 1816
rect 1435 1812 1436 1816
rect 1430 1811 1436 1812
rect 1502 1816 1508 1817
rect 1502 1812 1503 1816
rect 1507 1812 1508 1816
rect 1502 1811 1508 1812
rect 1582 1816 1588 1817
rect 1582 1812 1583 1816
rect 1587 1812 1588 1816
rect 1582 1811 1588 1812
rect 1670 1816 1676 1817
rect 1670 1812 1671 1816
rect 1675 1812 1676 1816
rect 1670 1811 1676 1812
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1870 1816 1876 1817
rect 1870 1812 1871 1816
rect 1875 1812 1876 1816
rect 1870 1811 1876 1812
rect 1982 1816 1988 1817
rect 1982 1812 1983 1816
rect 1987 1812 1988 1816
rect 1982 1811 1988 1812
rect 2070 1816 2076 1817
rect 2070 1812 2071 1816
rect 2075 1812 2076 1816
rect 2070 1811 2076 1812
rect 1155 1805 1190 1806
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 182 1804 188 1805
rect 182 1800 183 1804
rect 187 1800 188 1804
rect 182 1799 188 1800
rect 262 1804 268 1805
rect 262 1800 263 1804
rect 267 1800 268 1804
rect 262 1799 268 1800
rect 350 1804 356 1805
rect 350 1800 351 1804
rect 355 1800 356 1804
rect 350 1799 356 1800
rect 438 1804 444 1805
rect 438 1800 439 1804
rect 443 1800 444 1804
rect 438 1799 444 1800
rect 526 1804 532 1805
rect 526 1800 527 1804
rect 531 1800 532 1804
rect 526 1799 532 1800
rect 606 1804 612 1805
rect 606 1800 607 1804
rect 611 1800 612 1804
rect 606 1799 612 1800
rect 686 1804 692 1805
rect 686 1800 687 1804
rect 691 1800 692 1804
rect 686 1799 692 1800
rect 766 1804 772 1805
rect 766 1800 767 1804
rect 771 1800 772 1804
rect 766 1799 772 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 990 1804 996 1805
rect 990 1800 991 1804
rect 995 1800 996 1804
rect 990 1799 996 1800
rect 1046 1804 1052 1805
rect 1046 1800 1047 1804
rect 1051 1800 1052 1804
rect 1155 1801 1156 1805
rect 1160 1804 1190 1805
rect 1195 1805 1210 1806
rect 1160 1801 1161 1804
rect 1155 1800 1161 1801
rect 1195 1801 1196 1805
rect 1200 1804 1210 1805
rect 1200 1801 1201 1804
rect 1195 1800 1201 1801
rect 1235 1803 1241 1804
rect 1046 1799 1052 1800
rect 1235 1799 1236 1803
rect 1240 1799 1241 1803
rect 1235 1798 1241 1799
rect 1294 1803 1305 1804
rect 1294 1799 1295 1803
rect 1299 1799 1300 1803
rect 1304 1799 1305 1803
rect 1294 1798 1305 1799
rect 1358 1803 1369 1804
rect 1358 1799 1359 1803
rect 1363 1799 1364 1803
rect 1368 1799 1369 1803
rect 1358 1798 1369 1799
rect 1427 1803 1433 1804
rect 1427 1799 1428 1803
rect 1432 1802 1433 1803
rect 1438 1803 1444 1804
rect 1438 1802 1439 1803
rect 1432 1800 1439 1802
rect 1432 1799 1433 1800
rect 1427 1798 1433 1799
rect 1438 1799 1439 1800
rect 1443 1799 1444 1803
rect 1438 1798 1444 1799
rect 1494 1803 1505 1804
rect 1494 1799 1495 1803
rect 1499 1799 1500 1803
rect 1504 1799 1505 1803
rect 1494 1798 1505 1799
rect 1574 1803 1585 1804
rect 1574 1799 1575 1803
rect 1579 1799 1580 1803
rect 1584 1799 1585 1803
rect 1574 1798 1585 1799
rect 1662 1803 1673 1804
rect 1662 1799 1663 1803
rect 1667 1799 1668 1803
rect 1672 1799 1673 1803
rect 1662 1798 1673 1799
rect 1758 1803 1769 1804
rect 1758 1799 1759 1803
rect 1763 1799 1764 1803
rect 1768 1799 1769 1803
rect 1758 1798 1769 1799
rect 1862 1803 1873 1804
rect 1862 1799 1863 1803
rect 1867 1799 1868 1803
rect 1872 1799 1873 1803
rect 1862 1798 1873 1799
rect 1979 1803 1985 1804
rect 1979 1799 1980 1803
rect 1984 1802 1985 1803
rect 2047 1803 2053 1804
rect 2047 1802 2048 1803
rect 1984 1800 2048 1802
rect 1984 1799 1985 1800
rect 1979 1798 1985 1799
rect 2047 1799 2048 1800
rect 2052 1799 2053 1803
rect 2047 1798 2053 1799
rect 2062 1803 2073 1804
rect 2062 1799 2063 1803
rect 2067 1799 2068 1803
rect 2072 1799 2073 1803
rect 2062 1798 2073 1799
rect 110 1796 116 1797
rect 110 1792 111 1796
rect 115 1792 116 1796
rect 1094 1796 1100 1797
rect 1094 1792 1095 1796
rect 1099 1792 1100 1796
rect 1237 1794 1239 1798
rect 1374 1795 1380 1796
rect 1374 1794 1375 1795
rect 1237 1792 1375 1794
rect 110 1791 116 1792
rect 159 1791 168 1792
rect 159 1787 160 1791
rect 167 1787 168 1791
rect 159 1786 168 1787
rect 170 1791 176 1792
rect 170 1787 171 1791
rect 175 1790 176 1791
rect 207 1791 213 1792
rect 207 1790 208 1791
rect 175 1788 208 1790
rect 175 1787 176 1788
rect 170 1786 176 1787
rect 207 1787 208 1788
rect 212 1787 213 1791
rect 207 1786 213 1787
rect 287 1791 293 1792
rect 287 1787 288 1791
rect 292 1790 293 1791
rect 298 1791 304 1792
rect 298 1790 299 1791
rect 292 1788 299 1790
rect 292 1787 293 1788
rect 287 1786 293 1787
rect 298 1787 299 1788
rect 303 1787 304 1791
rect 298 1786 304 1787
rect 374 1791 381 1792
rect 374 1787 375 1791
rect 380 1787 381 1791
rect 374 1786 381 1787
rect 462 1791 469 1792
rect 462 1787 463 1791
rect 468 1787 469 1791
rect 462 1786 469 1787
rect 510 1791 516 1792
rect 510 1787 511 1791
rect 515 1790 516 1791
rect 551 1791 557 1792
rect 551 1790 552 1791
rect 515 1788 552 1790
rect 515 1787 516 1788
rect 510 1786 516 1787
rect 551 1787 552 1788
rect 556 1787 557 1791
rect 551 1786 557 1787
rect 631 1791 637 1792
rect 631 1787 632 1791
rect 636 1790 637 1791
rect 639 1791 645 1792
rect 639 1790 640 1791
rect 636 1788 640 1790
rect 636 1787 637 1788
rect 631 1786 637 1787
rect 639 1787 640 1788
rect 644 1787 645 1791
rect 639 1786 645 1787
rect 711 1791 720 1792
rect 711 1787 712 1791
rect 719 1787 720 1791
rect 711 1786 720 1787
rect 742 1791 748 1792
rect 742 1787 743 1791
rect 747 1790 748 1791
rect 791 1791 797 1792
rect 791 1790 792 1791
rect 747 1788 792 1790
rect 747 1787 748 1788
rect 742 1786 748 1787
rect 791 1787 792 1788
rect 796 1787 797 1791
rect 791 1786 797 1787
rect 863 1791 872 1792
rect 863 1787 864 1791
rect 871 1787 872 1791
rect 863 1786 872 1787
rect 935 1791 941 1792
rect 935 1787 936 1791
rect 940 1790 941 1791
rect 950 1791 956 1792
rect 950 1790 951 1791
rect 940 1788 951 1790
rect 940 1787 941 1788
rect 935 1786 941 1787
rect 950 1787 951 1788
rect 955 1787 956 1791
rect 950 1786 956 1787
rect 1014 1791 1021 1792
rect 1014 1787 1015 1791
rect 1020 1787 1021 1791
rect 1014 1786 1021 1787
rect 1034 1791 1040 1792
rect 1034 1787 1035 1791
rect 1039 1790 1040 1791
rect 1071 1791 1077 1792
rect 1094 1791 1100 1792
rect 1374 1791 1375 1792
rect 1379 1791 1380 1795
rect 1071 1790 1072 1791
rect 1039 1788 1072 1790
rect 1039 1787 1040 1788
rect 1034 1786 1040 1787
rect 1071 1787 1072 1788
rect 1076 1787 1077 1791
rect 1374 1790 1380 1791
rect 1071 1786 1077 1787
rect 1307 1783 1313 1784
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 1094 1779 1100 1780
rect 110 1774 116 1775
rect 134 1776 140 1777
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 182 1776 188 1777
rect 182 1772 183 1776
rect 187 1772 188 1776
rect 182 1771 188 1772
rect 262 1776 268 1777
rect 262 1772 263 1776
rect 267 1772 268 1776
rect 262 1771 268 1772
rect 350 1776 356 1777
rect 350 1772 351 1776
rect 355 1772 356 1776
rect 350 1771 356 1772
rect 438 1776 444 1777
rect 438 1772 439 1776
rect 443 1772 444 1776
rect 438 1771 444 1772
rect 526 1776 532 1777
rect 526 1772 527 1776
rect 531 1772 532 1776
rect 526 1771 532 1772
rect 606 1776 612 1777
rect 606 1772 607 1776
rect 611 1772 612 1776
rect 606 1771 612 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 766 1776 772 1777
rect 766 1772 767 1776
rect 771 1772 772 1776
rect 766 1771 772 1772
rect 838 1776 844 1777
rect 838 1772 839 1776
rect 843 1772 844 1776
rect 838 1771 844 1772
rect 910 1776 916 1777
rect 910 1772 911 1776
rect 915 1772 916 1776
rect 910 1771 916 1772
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1046 1776 1052 1777
rect 1046 1772 1047 1776
rect 1051 1772 1052 1776
rect 1094 1775 1095 1779
rect 1099 1775 1100 1779
rect 1307 1779 1308 1783
rect 1312 1782 1313 1783
rect 1330 1783 1336 1784
rect 1330 1782 1331 1783
rect 1312 1780 1331 1782
rect 1312 1779 1313 1780
rect 1307 1778 1313 1779
rect 1330 1779 1331 1780
rect 1335 1779 1336 1783
rect 1330 1778 1336 1779
rect 1338 1783 1344 1784
rect 1338 1779 1339 1783
rect 1343 1782 1344 1783
rect 1347 1783 1353 1784
rect 1347 1782 1348 1783
rect 1343 1780 1348 1782
rect 1343 1779 1344 1780
rect 1338 1778 1344 1779
rect 1347 1779 1348 1780
rect 1352 1779 1353 1783
rect 1347 1778 1353 1779
rect 1378 1783 1384 1784
rect 1378 1779 1379 1783
rect 1383 1782 1384 1783
rect 1387 1783 1393 1784
rect 1387 1782 1388 1783
rect 1383 1780 1388 1782
rect 1383 1779 1384 1780
rect 1378 1778 1384 1779
rect 1387 1779 1388 1780
rect 1392 1779 1393 1783
rect 1387 1778 1393 1779
rect 1418 1783 1424 1784
rect 1418 1779 1419 1783
rect 1423 1782 1424 1783
rect 1427 1783 1433 1784
rect 1427 1782 1428 1783
rect 1423 1780 1428 1782
rect 1423 1779 1424 1780
rect 1418 1778 1424 1779
rect 1427 1779 1428 1780
rect 1432 1779 1433 1783
rect 1427 1778 1433 1779
rect 1454 1783 1460 1784
rect 1454 1779 1455 1783
rect 1459 1782 1460 1783
rect 1467 1783 1473 1784
rect 1467 1782 1468 1783
rect 1459 1780 1468 1782
rect 1459 1779 1460 1780
rect 1454 1778 1460 1779
rect 1467 1779 1468 1780
rect 1472 1779 1473 1783
rect 1467 1778 1473 1779
rect 1494 1783 1500 1784
rect 1494 1779 1495 1783
rect 1499 1782 1500 1783
rect 1507 1783 1513 1784
rect 1507 1782 1508 1783
rect 1499 1780 1508 1782
rect 1499 1779 1500 1780
rect 1494 1778 1500 1779
rect 1507 1779 1508 1780
rect 1512 1779 1513 1783
rect 1507 1778 1513 1779
rect 1538 1783 1544 1784
rect 1538 1779 1539 1783
rect 1543 1782 1544 1783
rect 1547 1783 1553 1784
rect 1547 1782 1548 1783
rect 1543 1780 1548 1782
rect 1543 1779 1544 1780
rect 1538 1778 1544 1779
rect 1547 1779 1548 1780
rect 1552 1779 1553 1783
rect 1547 1778 1553 1779
rect 1583 1783 1589 1784
rect 1583 1779 1584 1783
rect 1588 1782 1589 1783
rect 1603 1783 1609 1784
rect 1603 1782 1604 1783
rect 1588 1780 1604 1782
rect 1588 1779 1589 1780
rect 1583 1778 1589 1779
rect 1603 1779 1604 1780
rect 1608 1779 1609 1783
rect 1603 1778 1609 1779
rect 1634 1783 1640 1784
rect 1634 1779 1635 1783
rect 1639 1782 1640 1783
rect 1675 1783 1681 1784
rect 1675 1782 1676 1783
rect 1639 1780 1676 1782
rect 1639 1779 1640 1780
rect 1634 1778 1640 1779
rect 1675 1779 1676 1780
rect 1680 1779 1681 1783
rect 1675 1778 1681 1779
rect 1706 1783 1712 1784
rect 1706 1779 1707 1783
rect 1711 1782 1712 1783
rect 1763 1783 1769 1784
rect 1763 1782 1764 1783
rect 1711 1780 1764 1782
rect 1711 1779 1712 1780
rect 1706 1778 1712 1779
rect 1763 1779 1764 1780
rect 1768 1779 1769 1783
rect 1763 1778 1769 1779
rect 1794 1783 1800 1784
rect 1794 1779 1795 1783
rect 1799 1782 1800 1783
rect 1867 1783 1873 1784
rect 1867 1782 1868 1783
rect 1799 1780 1868 1782
rect 1799 1779 1800 1780
rect 1794 1778 1800 1779
rect 1867 1779 1868 1780
rect 1872 1779 1873 1783
rect 1867 1778 1873 1779
rect 1898 1783 1904 1784
rect 1898 1779 1899 1783
rect 1903 1782 1904 1783
rect 1979 1783 1985 1784
rect 1979 1782 1980 1783
rect 1903 1780 1980 1782
rect 1903 1779 1904 1780
rect 1898 1778 1904 1779
rect 1979 1779 1980 1780
rect 1984 1779 1985 1783
rect 1979 1778 1985 1779
rect 2067 1783 2073 1784
rect 2067 1779 2068 1783
rect 2072 1782 2073 1783
rect 2078 1783 2084 1784
rect 2078 1782 2079 1783
rect 2072 1780 2079 1782
rect 2072 1779 2073 1780
rect 2067 1778 2073 1779
rect 2078 1779 2079 1780
rect 2083 1779 2084 1783
rect 2078 1778 2084 1779
rect 1094 1774 1100 1775
rect 1046 1771 1052 1772
rect 1310 1772 1316 1773
rect 1310 1768 1311 1772
rect 1315 1768 1316 1772
rect 1310 1767 1316 1768
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1430 1772 1436 1773
rect 1430 1768 1431 1772
rect 1435 1768 1436 1772
rect 1430 1767 1436 1768
rect 1470 1772 1476 1773
rect 1470 1768 1471 1772
rect 1475 1768 1476 1772
rect 1470 1767 1476 1768
rect 1510 1772 1516 1773
rect 1510 1768 1511 1772
rect 1515 1768 1516 1772
rect 1510 1767 1516 1768
rect 1550 1772 1556 1773
rect 1550 1768 1551 1772
rect 1555 1768 1556 1772
rect 1550 1767 1556 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1678 1772 1684 1773
rect 1678 1768 1679 1772
rect 1683 1768 1684 1772
rect 1678 1767 1684 1768
rect 1766 1772 1772 1773
rect 1766 1768 1767 1772
rect 1771 1768 1772 1772
rect 1766 1767 1772 1768
rect 1870 1772 1876 1773
rect 1870 1768 1871 1772
rect 1875 1768 1876 1772
rect 1870 1767 1876 1768
rect 1982 1772 1988 1773
rect 1982 1768 1983 1772
rect 1987 1768 1988 1772
rect 1982 1767 1988 1768
rect 2070 1772 2076 1773
rect 2070 1768 2071 1772
rect 2075 1768 2076 1772
rect 2070 1767 2076 1768
rect 1134 1764 1140 1765
rect 1134 1760 1135 1764
rect 1139 1760 1140 1764
rect 2118 1764 2124 1765
rect 2118 1760 2119 1764
rect 2123 1760 2124 1764
rect 1134 1759 1140 1760
rect 1335 1759 1344 1760
rect 134 1756 140 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 134 1752 135 1756
rect 139 1752 140 1756
rect 134 1751 140 1752
rect 198 1756 204 1757
rect 198 1752 199 1756
rect 203 1752 204 1756
rect 198 1751 204 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 398 1756 404 1757
rect 398 1752 399 1756
rect 403 1752 404 1756
rect 398 1751 404 1752
rect 494 1756 500 1757
rect 494 1752 495 1756
rect 499 1752 500 1756
rect 494 1751 500 1752
rect 590 1756 596 1757
rect 590 1752 591 1756
rect 595 1752 596 1756
rect 590 1751 596 1752
rect 670 1756 676 1757
rect 670 1752 671 1756
rect 675 1752 676 1756
rect 670 1751 676 1752
rect 750 1756 756 1757
rect 750 1752 751 1756
rect 755 1752 756 1756
rect 750 1751 756 1752
rect 822 1756 828 1757
rect 822 1752 823 1756
rect 827 1752 828 1756
rect 822 1751 828 1752
rect 886 1756 892 1757
rect 886 1752 887 1756
rect 891 1752 892 1756
rect 886 1751 892 1752
rect 958 1756 964 1757
rect 958 1752 959 1756
rect 963 1752 964 1756
rect 958 1751 964 1752
rect 1030 1756 1036 1757
rect 1030 1752 1031 1756
rect 1035 1752 1036 1756
rect 1335 1755 1336 1759
rect 1343 1755 1344 1759
rect 1335 1754 1344 1755
rect 1375 1759 1384 1760
rect 1375 1755 1376 1759
rect 1383 1755 1384 1759
rect 1375 1754 1384 1755
rect 1415 1759 1424 1760
rect 1415 1755 1416 1759
rect 1423 1755 1424 1759
rect 1415 1754 1424 1755
rect 1454 1759 1461 1760
rect 1454 1755 1455 1759
rect 1460 1755 1461 1759
rect 1454 1754 1461 1755
rect 1494 1759 1501 1760
rect 1494 1755 1495 1759
rect 1500 1755 1501 1759
rect 1494 1754 1501 1755
rect 1535 1759 1544 1760
rect 1535 1755 1536 1759
rect 1543 1755 1544 1759
rect 1535 1754 1544 1755
rect 1575 1759 1581 1760
rect 1575 1755 1576 1759
rect 1580 1758 1581 1759
rect 1583 1759 1589 1760
rect 1583 1758 1584 1759
rect 1580 1756 1584 1758
rect 1580 1755 1581 1756
rect 1575 1754 1581 1755
rect 1583 1755 1584 1756
rect 1588 1755 1589 1759
rect 1583 1754 1589 1755
rect 1631 1759 1640 1760
rect 1631 1755 1632 1759
rect 1639 1755 1640 1759
rect 1631 1754 1640 1755
rect 1703 1759 1712 1760
rect 1703 1755 1704 1759
rect 1711 1755 1712 1759
rect 1703 1754 1712 1755
rect 1791 1759 1800 1760
rect 1791 1755 1792 1759
rect 1799 1755 1800 1759
rect 1791 1754 1800 1755
rect 1895 1759 1904 1760
rect 1895 1755 1896 1759
rect 1903 1755 1904 1759
rect 1895 1754 1904 1755
rect 2006 1759 2013 1760
rect 2006 1755 2007 1759
rect 2012 1755 2013 1759
rect 2006 1754 2013 1755
rect 2090 1759 2101 1760
rect 2118 1759 2124 1760
rect 2090 1755 2091 1759
rect 2095 1755 2096 1759
rect 2100 1755 2101 1759
rect 2090 1754 2101 1755
rect 1030 1751 1036 1752
rect 1094 1753 1100 1754
rect 110 1748 116 1749
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 430 1747 436 1748
rect 430 1743 431 1747
rect 435 1746 436 1747
rect 910 1747 916 1748
rect 435 1744 530 1746
rect 435 1743 436 1744
rect 430 1742 436 1743
rect 159 1739 165 1740
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 159 1735 160 1739
rect 164 1738 165 1739
rect 182 1739 188 1740
rect 182 1738 183 1739
rect 164 1736 183 1738
rect 164 1735 165 1736
rect 159 1734 165 1735
rect 182 1735 183 1736
rect 187 1735 188 1739
rect 182 1734 188 1735
rect 223 1739 229 1740
rect 223 1735 224 1739
rect 228 1738 229 1739
rect 286 1739 292 1740
rect 286 1738 287 1739
rect 228 1736 287 1738
rect 228 1735 229 1736
rect 223 1734 229 1735
rect 286 1735 287 1736
rect 291 1735 292 1739
rect 286 1734 292 1735
rect 310 1739 316 1740
rect 310 1735 311 1739
rect 315 1738 316 1739
rect 319 1739 325 1740
rect 319 1738 320 1739
rect 315 1736 320 1738
rect 315 1735 316 1736
rect 310 1734 316 1735
rect 319 1735 320 1736
rect 324 1735 325 1739
rect 319 1734 325 1735
rect 423 1739 429 1740
rect 423 1735 424 1739
rect 428 1738 429 1739
rect 486 1739 492 1740
rect 486 1738 487 1739
rect 428 1736 487 1738
rect 428 1735 429 1736
rect 423 1734 429 1735
rect 486 1735 487 1736
rect 491 1735 492 1739
rect 486 1734 492 1735
rect 518 1739 525 1740
rect 518 1735 519 1739
rect 524 1735 525 1739
rect 528 1738 530 1744
rect 910 1743 911 1747
rect 915 1746 916 1747
rect 1134 1747 1140 1748
rect 915 1744 1034 1746
rect 915 1743 916 1744
rect 910 1742 916 1743
rect 615 1739 621 1740
rect 615 1738 616 1739
rect 528 1736 616 1738
rect 518 1734 525 1735
rect 615 1735 616 1736
rect 620 1735 621 1739
rect 615 1734 621 1735
rect 695 1739 701 1740
rect 695 1735 696 1739
rect 700 1738 701 1739
rect 742 1739 748 1740
rect 742 1738 743 1739
rect 700 1736 743 1738
rect 700 1735 701 1736
rect 695 1734 701 1735
rect 742 1735 743 1736
rect 747 1735 748 1739
rect 742 1734 748 1735
rect 775 1739 781 1740
rect 775 1735 776 1739
rect 780 1738 781 1739
rect 798 1739 804 1740
rect 798 1738 799 1739
rect 780 1736 799 1738
rect 780 1735 781 1736
rect 775 1734 781 1735
rect 798 1735 799 1736
rect 803 1735 804 1739
rect 798 1734 804 1735
rect 807 1739 813 1740
rect 807 1735 808 1739
rect 812 1738 813 1739
rect 847 1739 853 1740
rect 847 1738 848 1739
rect 812 1736 848 1738
rect 812 1735 813 1736
rect 807 1734 813 1735
rect 847 1735 848 1736
rect 852 1735 853 1739
rect 847 1734 853 1735
rect 855 1739 861 1740
rect 855 1735 856 1739
rect 860 1738 861 1739
rect 911 1739 917 1740
rect 911 1738 912 1739
rect 860 1736 912 1738
rect 860 1735 861 1736
rect 855 1734 861 1735
rect 911 1735 912 1736
rect 916 1735 917 1739
rect 911 1734 917 1735
rect 983 1739 989 1740
rect 983 1735 984 1739
rect 988 1738 989 1739
rect 1022 1739 1028 1740
rect 1022 1738 1023 1739
rect 988 1736 1023 1738
rect 988 1735 989 1736
rect 983 1734 989 1735
rect 1022 1735 1023 1736
rect 1027 1735 1028 1739
rect 1032 1738 1034 1744
rect 1134 1743 1135 1747
rect 1139 1743 1140 1747
rect 2118 1747 2124 1748
rect 1134 1742 1140 1743
rect 1310 1744 1316 1745
rect 1310 1740 1311 1744
rect 1315 1740 1316 1744
rect 1055 1739 1061 1740
rect 1310 1739 1316 1740
rect 1350 1744 1356 1745
rect 1350 1740 1351 1744
rect 1355 1740 1356 1744
rect 1350 1739 1356 1740
rect 1390 1744 1396 1745
rect 1390 1740 1391 1744
rect 1395 1740 1396 1744
rect 1390 1739 1396 1740
rect 1430 1744 1436 1745
rect 1430 1740 1431 1744
rect 1435 1740 1436 1744
rect 1430 1739 1436 1740
rect 1470 1744 1476 1745
rect 1470 1740 1471 1744
rect 1475 1740 1476 1744
rect 1470 1739 1476 1740
rect 1510 1744 1516 1745
rect 1510 1740 1511 1744
rect 1515 1740 1516 1744
rect 1510 1739 1516 1740
rect 1550 1744 1556 1745
rect 1550 1740 1551 1744
rect 1555 1740 1556 1744
rect 1550 1739 1556 1740
rect 1606 1744 1612 1745
rect 1606 1740 1607 1744
rect 1611 1740 1612 1744
rect 1606 1739 1612 1740
rect 1678 1744 1684 1745
rect 1678 1740 1679 1744
rect 1683 1740 1684 1744
rect 1678 1739 1684 1740
rect 1766 1744 1772 1745
rect 1766 1740 1767 1744
rect 1771 1740 1772 1744
rect 1766 1739 1772 1740
rect 1870 1744 1876 1745
rect 1870 1740 1871 1744
rect 1875 1740 1876 1744
rect 1870 1739 1876 1740
rect 1982 1744 1988 1745
rect 1982 1740 1983 1744
rect 1987 1740 1988 1744
rect 1982 1739 1988 1740
rect 2070 1744 2076 1745
rect 2070 1740 2071 1744
rect 2075 1740 2076 1744
rect 2118 1743 2119 1747
rect 2123 1743 2124 1747
rect 2118 1742 2124 1743
rect 2070 1739 2076 1740
rect 1055 1738 1056 1739
rect 1032 1736 1056 1738
rect 1022 1734 1028 1735
rect 1055 1735 1056 1736
rect 1060 1735 1061 1739
rect 1055 1734 1061 1735
rect 1094 1736 1100 1737
rect 110 1731 116 1732
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1094 1731 1100 1732
rect 134 1728 140 1729
rect 134 1724 135 1728
rect 139 1724 140 1728
rect 134 1723 140 1724
rect 198 1728 204 1729
rect 198 1724 199 1728
rect 203 1724 204 1728
rect 198 1723 204 1724
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 398 1728 404 1729
rect 398 1724 399 1728
rect 403 1724 404 1728
rect 398 1723 404 1724
rect 494 1728 500 1729
rect 494 1724 495 1728
rect 499 1724 500 1728
rect 494 1723 500 1724
rect 590 1728 596 1729
rect 590 1724 591 1728
rect 595 1724 596 1728
rect 590 1723 596 1724
rect 670 1728 676 1729
rect 670 1724 671 1728
rect 675 1724 676 1728
rect 670 1723 676 1724
rect 750 1728 756 1729
rect 750 1724 751 1728
rect 755 1724 756 1728
rect 750 1723 756 1724
rect 822 1728 828 1729
rect 822 1724 823 1728
rect 827 1724 828 1728
rect 822 1723 828 1724
rect 886 1728 892 1729
rect 886 1724 887 1728
rect 891 1724 892 1728
rect 886 1723 892 1724
rect 958 1728 964 1729
rect 958 1724 959 1728
rect 963 1724 964 1728
rect 958 1723 964 1724
rect 1030 1728 1036 1729
rect 1030 1724 1031 1728
rect 1035 1724 1036 1728
rect 1262 1728 1268 1729
rect 1030 1723 1036 1724
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1262 1724 1263 1728
rect 1267 1724 1268 1728
rect 1262 1723 1268 1724
rect 1318 1728 1324 1729
rect 1318 1724 1319 1728
rect 1323 1724 1324 1728
rect 1318 1723 1324 1724
rect 1382 1728 1388 1729
rect 1382 1724 1383 1728
rect 1387 1724 1388 1728
rect 1382 1723 1388 1724
rect 1454 1728 1460 1729
rect 1454 1724 1455 1728
rect 1459 1724 1460 1728
rect 1454 1723 1460 1724
rect 1534 1728 1540 1729
rect 1534 1724 1535 1728
rect 1539 1724 1540 1728
rect 1534 1723 1540 1724
rect 1614 1728 1620 1729
rect 1614 1724 1615 1728
rect 1619 1724 1620 1728
rect 1614 1723 1620 1724
rect 1686 1728 1692 1729
rect 1686 1724 1687 1728
rect 1691 1724 1692 1728
rect 1686 1723 1692 1724
rect 1758 1728 1764 1729
rect 1758 1724 1759 1728
rect 1763 1724 1764 1728
rect 1758 1723 1764 1724
rect 1830 1728 1836 1729
rect 1830 1724 1831 1728
rect 1835 1724 1836 1728
rect 1830 1723 1836 1724
rect 1894 1728 1900 1729
rect 1894 1724 1895 1728
rect 1899 1724 1900 1728
rect 1894 1723 1900 1724
rect 1958 1728 1964 1729
rect 1958 1724 1959 1728
rect 1963 1724 1964 1728
rect 1958 1723 1964 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 2118 1725 2124 1726
rect 1134 1720 1140 1721
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 1710 1719 1716 1720
rect 1332 1716 1618 1718
rect 131 1715 137 1716
rect 131 1711 132 1715
rect 136 1714 137 1715
rect 170 1715 176 1716
rect 170 1714 171 1715
rect 136 1712 171 1714
rect 136 1711 137 1712
rect 131 1710 137 1711
rect 170 1711 171 1712
rect 175 1711 176 1715
rect 170 1710 176 1711
rect 182 1715 188 1716
rect 182 1711 183 1715
rect 187 1714 188 1715
rect 195 1715 201 1716
rect 195 1714 196 1715
rect 187 1712 196 1714
rect 187 1711 188 1712
rect 182 1710 188 1711
rect 195 1711 196 1712
rect 200 1711 201 1715
rect 195 1710 201 1711
rect 286 1715 297 1716
rect 286 1711 287 1715
rect 291 1711 292 1715
rect 296 1711 297 1715
rect 286 1710 297 1711
rect 395 1715 401 1716
rect 395 1711 396 1715
rect 400 1714 401 1715
rect 430 1715 436 1716
rect 430 1714 431 1715
rect 400 1712 431 1714
rect 400 1711 401 1712
rect 395 1710 401 1711
rect 430 1711 431 1712
rect 435 1711 436 1715
rect 430 1710 436 1711
rect 486 1715 497 1716
rect 486 1711 487 1715
rect 491 1711 492 1715
rect 496 1711 497 1715
rect 486 1710 497 1711
rect 562 1715 568 1716
rect 562 1711 563 1715
rect 567 1714 568 1715
rect 587 1715 593 1716
rect 587 1714 588 1715
rect 567 1712 588 1714
rect 567 1711 568 1712
rect 562 1710 568 1711
rect 587 1711 588 1712
rect 592 1711 593 1715
rect 587 1710 593 1711
rect 667 1715 673 1716
rect 667 1711 668 1715
rect 672 1714 673 1715
rect 742 1715 753 1716
rect 672 1712 681 1714
rect 672 1711 673 1712
rect 667 1710 673 1711
rect 310 1707 316 1708
rect 310 1706 311 1707
rect 220 1704 311 1706
rect 220 1702 222 1704
rect 310 1703 311 1704
rect 315 1703 316 1707
rect 679 1706 681 1712
rect 742 1711 743 1715
rect 747 1711 748 1715
rect 752 1711 753 1715
rect 742 1710 753 1711
rect 819 1715 825 1716
rect 819 1711 820 1715
rect 824 1714 825 1715
rect 855 1715 861 1716
rect 855 1714 856 1715
rect 824 1712 856 1714
rect 824 1711 825 1712
rect 819 1710 825 1711
rect 855 1711 856 1712
rect 860 1711 861 1715
rect 855 1710 861 1711
rect 883 1715 889 1716
rect 883 1711 884 1715
rect 888 1714 889 1715
rect 910 1715 916 1716
rect 910 1714 911 1715
rect 888 1712 911 1714
rect 888 1711 889 1712
rect 883 1710 889 1711
rect 910 1711 911 1712
rect 915 1711 916 1715
rect 910 1710 916 1711
rect 950 1715 961 1716
rect 950 1711 951 1715
rect 955 1711 956 1715
rect 960 1711 961 1715
rect 950 1710 961 1711
rect 1022 1715 1033 1716
rect 1022 1711 1023 1715
rect 1027 1711 1028 1715
rect 1032 1711 1033 1715
rect 1330 1715 1336 1716
rect 1022 1710 1033 1711
rect 1287 1711 1293 1712
rect 1134 1708 1140 1709
rect 807 1707 813 1708
rect 807 1706 808 1707
rect 679 1704 808 1706
rect 310 1702 316 1703
rect 807 1703 808 1704
rect 812 1703 813 1707
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1287 1707 1288 1711
rect 1292 1710 1293 1711
rect 1310 1711 1316 1712
rect 1310 1710 1311 1711
rect 1292 1708 1311 1710
rect 1292 1707 1293 1708
rect 1287 1706 1293 1707
rect 1310 1707 1311 1708
rect 1315 1707 1316 1711
rect 1330 1711 1331 1715
rect 1335 1711 1336 1715
rect 1330 1710 1336 1711
rect 1343 1711 1349 1712
rect 1310 1706 1316 1707
rect 1343 1707 1344 1711
rect 1348 1710 1349 1711
rect 1374 1711 1380 1712
rect 1374 1710 1375 1711
rect 1348 1708 1375 1710
rect 1348 1707 1349 1708
rect 1343 1706 1349 1707
rect 1374 1707 1375 1708
rect 1379 1707 1380 1711
rect 1374 1706 1380 1707
rect 1407 1711 1413 1712
rect 1407 1707 1408 1711
rect 1412 1710 1413 1711
rect 1446 1711 1452 1712
rect 1446 1710 1447 1711
rect 1412 1708 1447 1710
rect 1412 1707 1413 1708
rect 1407 1706 1413 1707
rect 1446 1707 1447 1708
rect 1451 1707 1452 1711
rect 1446 1706 1452 1707
rect 1479 1711 1485 1712
rect 1479 1707 1480 1711
rect 1484 1710 1485 1711
rect 1526 1711 1532 1712
rect 1526 1710 1527 1711
rect 1484 1708 1527 1710
rect 1484 1707 1485 1708
rect 1479 1706 1485 1707
rect 1526 1707 1527 1708
rect 1531 1707 1532 1711
rect 1526 1706 1532 1707
rect 1559 1711 1565 1712
rect 1559 1707 1560 1711
rect 1564 1710 1565 1711
rect 1606 1711 1612 1712
rect 1606 1710 1607 1711
rect 1564 1708 1607 1710
rect 1564 1707 1565 1708
rect 1559 1706 1565 1707
rect 1606 1707 1607 1708
rect 1611 1707 1612 1711
rect 1616 1710 1618 1716
rect 1710 1715 1711 1719
rect 1715 1718 1716 1719
rect 1715 1716 1818 1718
rect 1715 1715 1716 1716
rect 1710 1714 1716 1715
rect 1639 1711 1645 1712
rect 1639 1710 1640 1711
rect 1616 1708 1640 1710
rect 1606 1706 1612 1707
rect 1639 1707 1640 1708
rect 1644 1707 1645 1711
rect 1639 1706 1645 1707
rect 1711 1711 1717 1712
rect 1711 1707 1712 1711
rect 1716 1710 1717 1711
rect 1742 1711 1748 1712
rect 1742 1710 1743 1711
rect 1716 1708 1743 1710
rect 1716 1707 1717 1708
rect 1711 1706 1717 1707
rect 1742 1707 1743 1708
rect 1747 1707 1748 1711
rect 1742 1706 1748 1707
rect 1783 1711 1789 1712
rect 1783 1707 1784 1711
rect 1788 1710 1789 1711
rect 1806 1711 1812 1712
rect 1806 1710 1807 1711
rect 1788 1708 1807 1710
rect 1788 1707 1789 1708
rect 1783 1706 1789 1707
rect 1806 1707 1807 1708
rect 1811 1707 1812 1711
rect 1816 1710 1818 1716
rect 1855 1711 1861 1712
rect 1855 1710 1856 1711
rect 1816 1708 1856 1710
rect 1806 1706 1812 1707
rect 1855 1707 1856 1708
rect 1860 1707 1861 1711
rect 1855 1706 1861 1707
rect 1863 1711 1869 1712
rect 1863 1707 1864 1711
rect 1868 1710 1869 1711
rect 1919 1711 1925 1712
rect 1919 1710 1920 1711
rect 1868 1708 1920 1710
rect 1868 1707 1869 1708
rect 1863 1706 1869 1707
rect 1919 1707 1920 1708
rect 1924 1707 1925 1711
rect 1919 1706 1925 1707
rect 1927 1711 1933 1712
rect 1927 1707 1928 1711
rect 1932 1710 1933 1711
rect 1983 1711 1989 1712
rect 1983 1710 1984 1711
rect 1932 1708 1984 1710
rect 1932 1707 1933 1708
rect 1927 1706 1933 1707
rect 1983 1707 1984 1708
rect 1988 1707 1989 1711
rect 1983 1706 1989 1707
rect 1991 1711 1997 1712
rect 1991 1707 1992 1711
rect 1996 1710 1997 1711
rect 2047 1711 2053 1712
rect 2047 1710 2048 1711
rect 1996 1708 2048 1710
rect 1996 1707 1997 1708
rect 1991 1706 1997 1707
rect 2047 1707 2048 1708
rect 2052 1707 2053 1711
rect 2047 1706 2053 1707
rect 2082 1711 2088 1712
rect 2082 1707 2083 1711
rect 2087 1710 2088 1711
rect 2095 1711 2101 1712
rect 2095 1710 2096 1711
rect 2087 1708 2096 1710
rect 2087 1707 2088 1708
rect 2082 1706 2088 1707
rect 2095 1707 2096 1708
rect 2100 1707 2101 1711
rect 2095 1706 2101 1707
rect 2118 1708 2124 1709
rect 1134 1703 1140 1704
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 807 1702 813 1703
rect 219 1701 225 1702
rect 147 1699 153 1700
rect 147 1695 148 1699
rect 152 1698 153 1699
rect 210 1699 216 1700
rect 210 1698 211 1699
rect 152 1696 211 1698
rect 152 1695 153 1696
rect 147 1694 153 1695
rect 210 1695 211 1696
rect 215 1695 216 1699
rect 219 1697 220 1701
rect 224 1697 225 1701
rect 1262 1700 1268 1701
rect 219 1696 225 1697
rect 299 1699 305 1700
rect 210 1694 216 1695
rect 299 1695 300 1699
rect 304 1698 305 1699
rect 322 1699 328 1700
rect 322 1698 323 1699
rect 304 1696 323 1698
rect 304 1695 305 1696
rect 299 1694 305 1695
rect 322 1695 323 1696
rect 327 1695 328 1699
rect 322 1694 328 1695
rect 330 1699 336 1700
rect 330 1695 331 1699
rect 335 1698 336 1699
rect 379 1699 385 1700
rect 379 1698 380 1699
rect 335 1696 380 1698
rect 335 1695 336 1696
rect 330 1694 336 1695
rect 379 1695 380 1696
rect 384 1695 385 1699
rect 379 1694 385 1695
rect 410 1699 416 1700
rect 410 1695 411 1699
rect 415 1698 416 1699
rect 459 1699 465 1700
rect 459 1698 460 1699
rect 415 1696 460 1698
rect 415 1695 416 1696
rect 410 1694 416 1695
rect 459 1695 460 1696
rect 464 1695 465 1699
rect 459 1694 465 1695
rect 495 1699 501 1700
rect 495 1695 496 1699
rect 500 1698 501 1699
rect 531 1699 537 1700
rect 531 1698 532 1699
rect 500 1696 532 1698
rect 500 1695 501 1696
rect 495 1694 501 1695
rect 531 1695 532 1696
rect 536 1695 537 1699
rect 531 1694 537 1695
rect 603 1699 609 1700
rect 603 1695 604 1699
rect 608 1698 609 1699
rect 658 1699 664 1700
rect 658 1698 659 1699
rect 608 1696 659 1698
rect 608 1695 609 1696
rect 603 1694 609 1695
rect 658 1695 659 1696
rect 663 1695 664 1699
rect 658 1694 664 1695
rect 667 1699 673 1700
rect 667 1695 668 1699
rect 672 1698 673 1699
rect 719 1699 725 1700
rect 719 1698 720 1699
rect 672 1696 720 1698
rect 672 1695 673 1696
rect 667 1694 673 1695
rect 719 1695 720 1696
rect 724 1695 725 1699
rect 719 1694 725 1695
rect 731 1699 737 1700
rect 731 1695 732 1699
rect 736 1698 737 1699
rect 790 1699 796 1700
rect 790 1698 791 1699
rect 736 1696 791 1698
rect 736 1695 737 1696
rect 731 1694 737 1695
rect 790 1695 791 1696
rect 795 1695 796 1699
rect 790 1694 796 1695
rect 798 1699 809 1700
rect 798 1695 799 1699
rect 803 1695 804 1699
rect 808 1695 809 1699
rect 798 1694 809 1695
rect 834 1699 840 1700
rect 834 1695 835 1699
rect 839 1698 840 1699
rect 875 1699 881 1700
rect 875 1698 876 1699
rect 839 1696 876 1698
rect 839 1695 840 1696
rect 834 1694 840 1695
rect 875 1695 876 1696
rect 880 1695 881 1699
rect 1262 1696 1263 1700
rect 1267 1696 1268 1700
rect 1262 1695 1268 1696
rect 1318 1700 1324 1701
rect 1318 1696 1319 1700
rect 1323 1696 1324 1700
rect 1318 1695 1324 1696
rect 1382 1700 1388 1701
rect 1382 1696 1383 1700
rect 1387 1696 1388 1700
rect 1382 1695 1388 1696
rect 1454 1700 1460 1701
rect 1454 1696 1455 1700
rect 1459 1696 1460 1700
rect 1454 1695 1460 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1614 1700 1620 1701
rect 1614 1696 1615 1700
rect 1619 1696 1620 1700
rect 1614 1695 1620 1696
rect 1686 1700 1692 1701
rect 1686 1696 1687 1700
rect 1691 1696 1692 1700
rect 1686 1695 1692 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1830 1700 1836 1701
rect 1830 1696 1831 1700
rect 1835 1696 1836 1700
rect 1830 1695 1836 1696
rect 1894 1700 1900 1701
rect 1894 1696 1895 1700
rect 1899 1696 1900 1700
rect 1894 1695 1900 1696
rect 1958 1700 1964 1701
rect 1958 1696 1959 1700
rect 1963 1696 1964 1700
rect 1958 1695 1964 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 875 1694 881 1695
rect 150 1688 156 1689
rect 150 1684 151 1688
rect 155 1684 156 1688
rect 150 1683 156 1684
rect 222 1688 228 1689
rect 222 1684 223 1688
rect 227 1684 228 1688
rect 222 1683 228 1684
rect 302 1688 308 1689
rect 302 1684 303 1688
rect 307 1684 308 1688
rect 302 1683 308 1684
rect 382 1688 388 1689
rect 382 1684 383 1688
rect 387 1684 388 1688
rect 382 1683 388 1684
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 534 1688 540 1689
rect 534 1684 535 1688
rect 539 1684 540 1688
rect 534 1683 540 1684
rect 606 1688 612 1689
rect 606 1684 607 1688
rect 611 1684 612 1688
rect 606 1683 612 1684
rect 670 1688 676 1689
rect 670 1684 671 1688
rect 675 1684 676 1688
rect 670 1683 676 1684
rect 734 1688 740 1689
rect 734 1684 735 1688
rect 739 1684 740 1688
rect 734 1683 740 1684
rect 806 1688 812 1689
rect 806 1684 807 1688
rect 811 1684 812 1688
rect 806 1683 812 1684
rect 878 1688 884 1689
rect 878 1684 879 1688
rect 883 1684 884 1688
rect 878 1683 884 1684
rect 1259 1687 1265 1688
rect 1259 1683 1260 1687
rect 1264 1686 1265 1687
rect 1302 1687 1308 1688
rect 1302 1686 1303 1687
rect 1264 1684 1303 1686
rect 1264 1683 1265 1684
rect 1259 1682 1265 1683
rect 1302 1683 1303 1684
rect 1307 1683 1308 1687
rect 1302 1682 1308 1683
rect 1310 1687 1321 1688
rect 1310 1683 1311 1687
rect 1315 1683 1316 1687
rect 1320 1683 1321 1687
rect 1310 1682 1321 1683
rect 1374 1687 1385 1688
rect 1374 1683 1375 1687
rect 1379 1683 1380 1687
rect 1384 1683 1385 1687
rect 1374 1682 1385 1683
rect 1446 1687 1457 1688
rect 1446 1683 1447 1687
rect 1451 1683 1452 1687
rect 1456 1683 1457 1687
rect 1446 1682 1457 1683
rect 1526 1687 1537 1688
rect 1526 1683 1527 1687
rect 1531 1683 1532 1687
rect 1536 1683 1537 1687
rect 1526 1682 1537 1683
rect 1606 1687 1617 1688
rect 1606 1683 1607 1687
rect 1611 1683 1612 1687
rect 1616 1683 1617 1687
rect 1606 1682 1617 1683
rect 1683 1687 1689 1688
rect 1683 1683 1684 1687
rect 1688 1686 1689 1687
rect 1710 1687 1716 1688
rect 1710 1686 1711 1687
rect 1688 1684 1711 1686
rect 1688 1683 1689 1684
rect 1683 1682 1689 1683
rect 1710 1683 1711 1684
rect 1715 1683 1716 1687
rect 1710 1682 1716 1683
rect 1742 1687 1748 1688
rect 1742 1683 1743 1687
rect 1747 1686 1748 1687
rect 1755 1687 1761 1688
rect 1755 1686 1756 1687
rect 1747 1684 1756 1686
rect 1747 1683 1748 1684
rect 1742 1682 1748 1683
rect 1755 1683 1756 1684
rect 1760 1683 1761 1687
rect 1755 1682 1761 1683
rect 1827 1687 1833 1688
rect 1827 1683 1828 1687
rect 1832 1686 1833 1687
rect 1863 1687 1869 1688
rect 1863 1686 1864 1687
rect 1832 1684 1864 1686
rect 1832 1683 1833 1684
rect 1827 1682 1833 1683
rect 1863 1683 1864 1684
rect 1868 1683 1869 1687
rect 1863 1682 1869 1683
rect 1891 1687 1897 1688
rect 1891 1683 1892 1687
rect 1896 1686 1897 1687
rect 1927 1687 1933 1688
rect 1927 1686 1928 1687
rect 1896 1684 1928 1686
rect 1896 1683 1897 1684
rect 1891 1682 1897 1683
rect 1927 1683 1928 1684
rect 1932 1683 1933 1687
rect 1927 1682 1933 1683
rect 1955 1687 1961 1688
rect 1955 1683 1956 1687
rect 1960 1686 1961 1687
rect 1991 1687 1997 1688
rect 1991 1686 1992 1687
rect 1960 1684 1992 1686
rect 1960 1683 1961 1684
rect 1955 1682 1961 1683
rect 1991 1683 1992 1684
rect 1996 1683 1997 1687
rect 1991 1682 1997 1683
rect 2010 1687 2016 1688
rect 2010 1683 2011 1687
rect 2015 1686 2016 1687
rect 2019 1687 2025 1688
rect 2019 1686 2020 1687
rect 2015 1684 2020 1686
rect 2015 1683 2016 1684
rect 2010 1682 2016 1683
rect 2019 1683 2020 1684
rect 2024 1683 2025 1687
rect 2019 1682 2025 1683
rect 2067 1687 2073 1688
rect 2067 1683 2068 1687
rect 2072 1686 2073 1687
rect 2090 1687 2096 1688
rect 2090 1686 2091 1687
rect 2072 1684 2091 1686
rect 2072 1683 2073 1684
rect 2067 1682 2073 1683
rect 2090 1683 2091 1684
rect 2095 1683 2096 1687
rect 2090 1682 2096 1683
rect 110 1680 116 1681
rect 824 1680 846 1682
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 790 1679 796 1680
rect 110 1675 116 1676
rect 166 1675 172 1676
rect 166 1671 167 1675
rect 171 1674 172 1675
rect 175 1675 181 1676
rect 175 1674 176 1675
rect 171 1672 176 1674
rect 171 1671 172 1672
rect 166 1670 172 1671
rect 175 1671 176 1672
rect 180 1671 181 1675
rect 175 1670 181 1671
rect 210 1675 216 1676
rect 210 1671 211 1675
rect 215 1674 216 1675
rect 247 1675 253 1676
rect 247 1674 248 1675
rect 215 1672 248 1674
rect 215 1671 216 1672
rect 210 1670 216 1671
rect 247 1671 248 1672
rect 252 1671 253 1675
rect 247 1670 253 1671
rect 327 1675 336 1676
rect 327 1671 328 1675
rect 335 1671 336 1675
rect 327 1670 336 1671
rect 407 1675 416 1676
rect 407 1671 408 1675
rect 415 1671 416 1675
rect 407 1670 416 1671
rect 487 1675 493 1676
rect 487 1671 488 1675
rect 492 1674 493 1675
rect 495 1675 501 1676
rect 495 1674 496 1675
rect 492 1672 496 1674
rect 492 1671 493 1672
rect 487 1670 493 1671
rect 495 1671 496 1672
rect 500 1671 501 1675
rect 495 1670 501 1671
rect 559 1675 568 1676
rect 559 1671 560 1675
rect 567 1671 568 1675
rect 559 1670 568 1671
rect 631 1675 637 1676
rect 631 1671 632 1675
rect 636 1674 637 1675
rect 654 1675 660 1676
rect 654 1674 655 1675
rect 636 1672 655 1674
rect 636 1671 637 1672
rect 631 1670 637 1671
rect 654 1671 655 1672
rect 659 1671 660 1675
rect 654 1670 660 1671
rect 662 1675 668 1676
rect 662 1671 663 1675
rect 667 1674 668 1675
rect 695 1675 701 1676
rect 695 1674 696 1675
rect 667 1672 696 1674
rect 667 1671 668 1672
rect 662 1670 668 1671
rect 695 1671 696 1672
rect 700 1671 701 1675
rect 695 1670 701 1671
rect 719 1675 725 1676
rect 719 1671 720 1675
rect 724 1674 725 1675
rect 759 1675 765 1676
rect 759 1674 760 1675
rect 724 1672 760 1674
rect 724 1671 725 1672
rect 719 1670 725 1671
rect 759 1671 760 1672
rect 764 1671 765 1675
rect 790 1675 791 1679
rect 795 1678 796 1679
rect 824 1678 826 1680
rect 795 1676 826 1678
rect 795 1675 796 1676
rect 790 1674 796 1675
rect 831 1675 840 1676
rect 759 1670 765 1671
rect 831 1671 832 1675
rect 839 1671 840 1675
rect 844 1674 846 1680
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 903 1675 909 1676
rect 1094 1675 1100 1676
rect 1163 1675 1169 1676
rect 903 1674 904 1675
rect 844 1672 904 1674
rect 831 1670 840 1671
rect 903 1671 904 1672
rect 908 1671 909 1675
rect 903 1670 909 1671
rect 1163 1671 1164 1675
rect 1168 1674 1169 1675
rect 1186 1675 1192 1676
rect 1186 1674 1187 1675
rect 1168 1672 1187 1674
rect 1168 1671 1169 1672
rect 1163 1670 1169 1671
rect 1186 1671 1187 1672
rect 1191 1671 1192 1675
rect 1186 1670 1192 1671
rect 1194 1675 1200 1676
rect 1194 1671 1195 1675
rect 1199 1674 1200 1675
rect 1243 1675 1249 1676
rect 1243 1674 1244 1675
rect 1199 1672 1244 1674
rect 1199 1671 1200 1672
rect 1194 1670 1200 1671
rect 1243 1671 1244 1672
rect 1248 1671 1249 1675
rect 1243 1670 1249 1671
rect 1274 1675 1280 1676
rect 1274 1671 1275 1675
rect 1279 1674 1280 1675
rect 1331 1675 1337 1676
rect 1331 1674 1332 1675
rect 1279 1672 1332 1674
rect 1279 1671 1280 1672
rect 1274 1670 1280 1671
rect 1331 1671 1332 1672
rect 1336 1671 1337 1675
rect 1331 1670 1337 1671
rect 1362 1675 1368 1676
rect 1362 1671 1363 1675
rect 1367 1674 1368 1675
rect 1419 1675 1425 1676
rect 1419 1674 1420 1675
rect 1367 1672 1420 1674
rect 1367 1671 1368 1672
rect 1362 1670 1368 1671
rect 1419 1671 1420 1672
rect 1424 1671 1425 1675
rect 1419 1670 1425 1671
rect 1455 1675 1461 1676
rect 1455 1671 1456 1675
rect 1460 1674 1461 1675
rect 1507 1675 1513 1676
rect 1507 1674 1508 1675
rect 1460 1672 1508 1674
rect 1460 1671 1461 1672
rect 1455 1670 1461 1671
rect 1507 1671 1508 1672
rect 1512 1671 1513 1675
rect 1507 1670 1513 1671
rect 1595 1675 1601 1676
rect 1595 1671 1596 1675
rect 1600 1674 1601 1675
rect 1626 1675 1632 1676
rect 1600 1672 1622 1674
rect 1600 1671 1601 1672
rect 1595 1670 1601 1671
rect 1618 1671 1624 1672
rect 1618 1667 1619 1671
rect 1623 1667 1624 1671
rect 1626 1671 1627 1675
rect 1631 1674 1632 1675
rect 1675 1675 1681 1676
rect 1675 1674 1676 1675
rect 1631 1672 1676 1674
rect 1631 1671 1632 1672
rect 1626 1670 1632 1671
rect 1675 1671 1676 1672
rect 1680 1671 1681 1675
rect 1675 1670 1681 1671
rect 1747 1675 1753 1676
rect 1747 1671 1748 1675
rect 1752 1674 1753 1675
rect 1798 1675 1804 1676
rect 1798 1674 1799 1675
rect 1752 1672 1799 1674
rect 1752 1671 1753 1672
rect 1747 1670 1753 1671
rect 1798 1671 1799 1672
rect 1803 1671 1804 1675
rect 1798 1670 1804 1671
rect 1806 1675 1817 1676
rect 1806 1671 1807 1675
rect 1811 1671 1812 1675
rect 1816 1671 1817 1675
rect 1806 1670 1817 1671
rect 1867 1675 1873 1676
rect 1867 1671 1868 1675
rect 1872 1674 1873 1675
rect 1906 1675 1912 1676
rect 1872 1672 1902 1674
rect 1872 1671 1873 1672
rect 1867 1670 1873 1671
rect 1618 1666 1624 1667
rect 1166 1664 1172 1665
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 1094 1663 1100 1664
rect 110 1658 116 1659
rect 150 1660 156 1661
rect 150 1656 151 1660
rect 155 1656 156 1660
rect 150 1655 156 1656
rect 222 1660 228 1661
rect 222 1656 223 1660
rect 227 1656 228 1660
rect 222 1655 228 1656
rect 302 1660 308 1661
rect 302 1656 303 1660
rect 307 1656 308 1660
rect 302 1655 308 1656
rect 382 1660 388 1661
rect 382 1656 383 1660
rect 387 1656 388 1660
rect 382 1655 388 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 534 1660 540 1661
rect 534 1656 535 1660
rect 539 1656 540 1660
rect 534 1655 540 1656
rect 606 1660 612 1661
rect 606 1656 607 1660
rect 611 1656 612 1660
rect 606 1655 612 1656
rect 670 1660 676 1661
rect 670 1656 671 1660
rect 675 1656 676 1660
rect 670 1655 676 1656
rect 734 1660 740 1661
rect 734 1656 735 1660
rect 739 1656 740 1660
rect 734 1655 740 1656
rect 806 1660 812 1661
rect 806 1656 807 1660
rect 811 1656 812 1660
rect 806 1655 812 1656
rect 878 1660 884 1661
rect 878 1656 879 1660
rect 883 1656 884 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1166 1660 1167 1664
rect 1171 1660 1172 1664
rect 1166 1659 1172 1660
rect 1246 1664 1252 1665
rect 1246 1660 1247 1664
rect 1251 1660 1252 1664
rect 1246 1659 1252 1660
rect 1334 1664 1340 1665
rect 1334 1660 1335 1664
rect 1339 1660 1340 1664
rect 1334 1659 1340 1660
rect 1422 1664 1428 1665
rect 1422 1660 1423 1664
rect 1427 1660 1428 1664
rect 1422 1659 1428 1660
rect 1510 1664 1516 1665
rect 1510 1660 1511 1664
rect 1515 1660 1516 1664
rect 1510 1659 1516 1660
rect 1598 1664 1604 1665
rect 1598 1660 1599 1664
rect 1603 1660 1604 1664
rect 1598 1659 1604 1660
rect 1678 1664 1684 1665
rect 1678 1660 1679 1664
rect 1683 1660 1684 1664
rect 1678 1659 1684 1660
rect 1750 1664 1756 1665
rect 1750 1660 1751 1664
rect 1755 1660 1756 1664
rect 1750 1659 1756 1660
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 1094 1658 1100 1659
rect 1900 1658 1902 1672
rect 1906 1671 1907 1675
rect 1911 1674 1912 1675
rect 1923 1675 1929 1676
rect 1923 1674 1924 1675
rect 1911 1672 1924 1674
rect 1911 1671 1912 1672
rect 1906 1670 1912 1671
rect 1923 1671 1924 1672
rect 1928 1671 1929 1675
rect 1923 1670 1929 1671
rect 1959 1675 1965 1676
rect 1959 1671 1960 1675
rect 1964 1674 1965 1675
rect 1979 1675 1985 1676
rect 1979 1674 1980 1675
rect 1964 1672 1980 1674
rect 1964 1671 1965 1672
rect 1959 1670 1965 1671
rect 1979 1671 1980 1672
rect 1984 1671 1985 1675
rect 1979 1670 1985 1671
rect 2027 1675 2033 1676
rect 2027 1671 2028 1675
rect 2032 1674 2033 1675
rect 2067 1675 2073 1676
rect 2032 1672 2062 1674
rect 2032 1671 2033 1672
rect 2027 1670 2033 1671
rect 1926 1664 1932 1665
rect 1926 1660 1927 1664
rect 1931 1660 1932 1664
rect 1926 1659 1932 1660
rect 1982 1664 1988 1665
rect 1982 1660 1983 1664
rect 1987 1660 1988 1664
rect 1982 1659 1988 1660
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2060 1658 2062 1672
rect 2067 1671 2068 1675
rect 2072 1674 2073 1675
rect 2082 1675 2088 1676
rect 2082 1674 2083 1675
rect 2072 1672 2083 1674
rect 2072 1671 2073 1672
rect 2067 1670 2073 1671
rect 2082 1671 2083 1672
rect 2087 1671 2088 1675
rect 2082 1670 2088 1671
rect 2070 1664 2076 1665
rect 2070 1660 2071 1664
rect 2075 1660 2076 1664
rect 2070 1659 2076 1660
rect 878 1655 884 1656
rect 1134 1656 1140 1657
rect 1352 1656 1418 1658
rect 1134 1652 1135 1656
rect 1139 1652 1140 1656
rect 1302 1655 1308 1656
rect 470 1651 476 1652
rect 1134 1651 1140 1652
rect 1191 1651 1200 1652
rect 470 1647 471 1651
rect 475 1650 476 1651
rect 475 1648 634 1650
rect 475 1647 476 1648
rect 470 1646 476 1647
rect 174 1644 180 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 174 1640 175 1644
rect 179 1640 180 1644
rect 174 1639 180 1640
rect 214 1644 220 1645
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 254 1644 260 1645
rect 254 1640 255 1644
rect 259 1640 260 1644
rect 254 1639 260 1640
rect 302 1644 308 1645
rect 302 1640 303 1644
rect 307 1640 308 1644
rect 302 1639 308 1640
rect 358 1644 364 1645
rect 358 1640 359 1644
rect 363 1640 364 1644
rect 358 1639 364 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 454 1644 460 1645
rect 454 1640 455 1644
rect 459 1640 460 1644
rect 454 1639 460 1640
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 550 1644 556 1645
rect 550 1640 551 1644
rect 555 1640 556 1644
rect 550 1639 556 1640
rect 606 1644 612 1645
rect 606 1640 607 1644
rect 611 1640 612 1644
rect 606 1639 612 1640
rect 110 1636 116 1637
rect 330 1635 336 1636
rect 330 1631 331 1635
rect 335 1634 336 1635
rect 534 1635 540 1636
rect 335 1632 410 1634
rect 335 1631 336 1632
rect 330 1630 336 1631
rect 199 1627 208 1628
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 199 1623 200 1627
rect 207 1623 208 1627
rect 199 1622 208 1623
rect 239 1627 248 1628
rect 239 1623 240 1627
rect 247 1623 248 1627
rect 239 1622 248 1623
rect 278 1627 285 1628
rect 278 1623 279 1627
rect 284 1623 285 1627
rect 278 1622 285 1623
rect 322 1627 333 1628
rect 322 1623 323 1627
rect 327 1623 328 1627
rect 332 1623 333 1627
rect 322 1622 333 1623
rect 383 1627 389 1628
rect 383 1623 384 1627
rect 388 1626 389 1627
rect 398 1627 404 1628
rect 398 1626 399 1627
rect 388 1624 399 1626
rect 388 1623 389 1624
rect 383 1622 389 1623
rect 398 1623 399 1624
rect 403 1623 404 1627
rect 408 1626 410 1632
rect 534 1631 535 1635
rect 539 1634 540 1635
rect 632 1634 634 1648
rect 1191 1647 1192 1651
rect 1199 1647 1200 1651
rect 1191 1646 1200 1647
rect 1271 1651 1280 1652
rect 1271 1647 1272 1651
rect 1279 1647 1280 1651
rect 1302 1651 1303 1655
rect 1307 1654 1308 1655
rect 1352 1654 1354 1656
rect 1307 1652 1354 1654
rect 1416 1654 1418 1656
rect 1440 1656 1466 1658
rect 1900 1656 1922 1658
rect 1440 1654 1442 1656
rect 1416 1652 1442 1654
rect 1307 1651 1308 1652
rect 1302 1650 1308 1651
rect 1359 1651 1368 1652
rect 1271 1646 1280 1647
rect 1359 1647 1360 1651
rect 1367 1647 1368 1651
rect 1359 1646 1368 1647
rect 1447 1651 1453 1652
rect 1447 1647 1448 1651
rect 1452 1650 1453 1651
rect 1455 1651 1461 1652
rect 1455 1650 1456 1651
rect 1452 1648 1456 1650
rect 1452 1647 1453 1648
rect 1447 1646 1453 1647
rect 1455 1647 1456 1648
rect 1460 1647 1461 1651
rect 1464 1650 1466 1656
rect 1920 1654 1922 1656
rect 1944 1656 1970 1658
rect 1944 1654 1946 1656
rect 1920 1652 1946 1654
rect 1968 1654 1970 1656
rect 1999 1656 2026 1658
rect 2060 1656 2066 1658
rect 1999 1654 2001 1656
rect 1968 1652 2001 1654
rect 1535 1651 1541 1652
rect 1535 1650 1536 1651
rect 1464 1648 1536 1650
rect 1455 1646 1461 1647
rect 1535 1647 1536 1648
rect 1540 1647 1541 1651
rect 1535 1646 1541 1647
rect 1623 1651 1632 1652
rect 1623 1647 1624 1651
rect 1631 1647 1632 1651
rect 1623 1646 1632 1647
rect 1703 1651 1709 1652
rect 1703 1647 1704 1651
rect 1708 1650 1709 1651
rect 1742 1651 1748 1652
rect 1742 1650 1743 1651
rect 1708 1648 1743 1650
rect 1708 1647 1709 1648
rect 1703 1646 1709 1647
rect 1742 1647 1743 1648
rect 1747 1647 1748 1651
rect 1742 1646 1748 1647
rect 1774 1651 1781 1652
rect 1774 1647 1775 1651
rect 1780 1647 1781 1651
rect 1774 1646 1781 1647
rect 1798 1651 1804 1652
rect 1798 1647 1799 1651
rect 1803 1650 1804 1651
rect 1839 1651 1845 1652
rect 1839 1650 1840 1651
rect 1803 1648 1840 1650
rect 1803 1647 1804 1648
rect 1798 1646 1804 1647
rect 1839 1647 1840 1648
rect 1844 1647 1845 1651
rect 1839 1646 1845 1647
rect 1895 1651 1901 1652
rect 1895 1647 1896 1651
rect 1900 1650 1901 1651
rect 1906 1651 1912 1652
rect 1906 1650 1907 1651
rect 1900 1648 1907 1650
rect 1900 1647 1901 1648
rect 1895 1646 1901 1647
rect 1906 1647 1907 1648
rect 1911 1647 1912 1651
rect 1906 1646 1912 1647
rect 1951 1651 1957 1652
rect 1951 1647 1952 1651
rect 1956 1650 1957 1651
rect 1959 1651 1965 1652
rect 1959 1650 1960 1651
rect 1956 1648 1960 1650
rect 1956 1647 1957 1648
rect 1951 1646 1957 1647
rect 1959 1647 1960 1648
rect 1964 1647 1965 1651
rect 1959 1646 1965 1647
rect 2007 1651 2016 1652
rect 2007 1647 2008 1651
rect 2015 1647 2016 1651
rect 2024 1650 2026 1656
rect 2055 1651 2061 1652
rect 2055 1650 2056 1651
rect 2024 1648 2056 1650
rect 2007 1646 2016 1647
rect 2055 1647 2056 1648
rect 2060 1647 2061 1651
rect 2064 1650 2066 1656
rect 2118 1656 2124 1657
rect 2118 1652 2119 1656
rect 2123 1652 2124 1656
rect 2095 1651 2101 1652
rect 2118 1651 2124 1652
rect 2095 1650 2096 1651
rect 2064 1648 2096 1650
rect 2055 1646 2061 1647
rect 2095 1647 2096 1648
rect 2100 1647 2101 1651
rect 2095 1646 2101 1647
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 718 1644 724 1645
rect 718 1640 719 1644
rect 723 1640 724 1644
rect 718 1639 724 1640
rect 1094 1641 1100 1642
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1639 1140 1640
rect 1134 1635 1135 1639
rect 1139 1635 1140 1639
rect 2118 1639 2124 1640
rect 1134 1634 1140 1635
rect 1166 1636 1172 1637
rect 539 1632 610 1634
rect 632 1632 722 1634
rect 539 1631 540 1632
rect 534 1630 540 1631
rect 431 1627 437 1628
rect 431 1626 432 1627
rect 408 1624 432 1626
rect 398 1622 404 1623
rect 431 1623 432 1624
rect 436 1623 437 1627
rect 431 1622 437 1623
rect 479 1627 485 1628
rect 479 1623 480 1627
rect 484 1626 485 1627
rect 494 1627 500 1628
rect 494 1626 495 1627
rect 484 1624 495 1626
rect 484 1623 485 1624
rect 479 1622 485 1623
rect 494 1623 495 1624
rect 499 1623 500 1627
rect 494 1622 500 1623
rect 527 1627 533 1628
rect 527 1623 528 1627
rect 532 1626 533 1627
rect 542 1627 548 1628
rect 542 1626 543 1627
rect 532 1624 543 1626
rect 532 1623 533 1624
rect 527 1622 533 1623
rect 542 1623 543 1624
rect 547 1623 548 1627
rect 542 1622 548 1623
rect 575 1627 581 1628
rect 575 1623 576 1627
rect 580 1626 581 1627
rect 598 1627 604 1628
rect 598 1626 599 1627
rect 580 1624 599 1626
rect 580 1623 581 1624
rect 575 1622 581 1623
rect 598 1623 599 1624
rect 603 1623 604 1627
rect 608 1626 610 1632
rect 631 1627 637 1628
rect 631 1626 632 1627
rect 608 1624 632 1626
rect 598 1622 604 1623
rect 631 1623 632 1624
rect 636 1623 637 1627
rect 631 1622 637 1623
rect 687 1627 693 1628
rect 687 1623 688 1627
rect 692 1626 693 1627
rect 710 1627 716 1628
rect 710 1626 711 1627
rect 692 1624 711 1626
rect 692 1623 693 1624
rect 687 1622 693 1623
rect 710 1623 711 1624
rect 715 1623 716 1627
rect 720 1626 722 1632
rect 1166 1632 1167 1636
rect 1171 1632 1172 1636
rect 1166 1631 1172 1632
rect 1246 1636 1252 1637
rect 1246 1632 1247 1636
rect 1251 1632 1252 1636
rect 1246 1631 1252 1632
rect 1334 1636 1340 1637
rect 1334 1632 1335 1636
rect 1339 1632 1340 1636
rect 1334 1631 1340 1632
rect 1422 1636 1428 1637
rect 1422 1632 1423 1636
rect 1427 1632 1428 1636
rect 1422 1631 1428 1632
rect 1510 1636 1516 1637
rect 1510 1632 1511 1636
rect 1515 1632 1516 1636
rect 1510 1631 1516 1632
rect 1598 1636 1604 1637
rect 1598 1632 1599 1636
rect 1603 1632 1604 1636
rect 1598 1631 1604 1632
rect 1678 1636 1684 1637
rect 1678 1632 1679 1636
rect 1683 1632 1684 1636
rect 1678 1631 1684 1632
rect 1750 1636 1756 1637
rect 1750 1632 1751 1636
rect 1755 1632 1756 1636
rect 1750 1631 1756 1632
rect 1814 1636 1820 1637
rect 1814 1632 1815 1636
rect 1819 1632 1820 1636
rect 1814 1631 1820 1632
rect 1870 1636 1876 1637
rect 1870 1632 1871 1636
rect 1875 1632 1876 1636
rect 1870 1631 1876 1632
rect 1926 1636 1932 1637
rect 1926 1632 1927 1636
rect 1931 1632 1932 1636
rect 1926 1631 1932 1632
rect 1982 1636 1988 1637
rect 1982 1632 1983 1636
rect 1987 1632 1988 1636
rect 1982 1631 1988 1632
rect 2030 1636 2036 1637
rect 2030 1632 2031 1636
rect 2035 1632 2036 1636
rect 2030 1631 2036 1632
rect 2070 1636 2076 1637
rect 2070 1632 2071 1636
rect 2075 1632 2076 1636
rect 2118 1635 2119 1639
rect 2123 1635 2124 1639
rect 2118 1634 2124 1635
rect 2070 1631 2076 1632
rect 743 1627 749 1628
rect 743 1626 744 1627
rect 720 1624 744 1626
rect 710 1622 716 1623
rect 743 1623 744 1624
rect 748 1623 749 1627
rect 1178 1627 1184 1628
rect 743 1622 749 1623
rect 1094 1624 1100 1625
rect 110 1619 116 1620
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1178 1623 1179 1627
rect 1183 1626 1184 1627
rect 1470 1627 1476 1628
rect 1470 1626 1471 1627
rect 1183 1624 1471 1626
rect 1183 1623 1184 1624
rect 1178 1622 1184 1623
rect 1470 1623 1471 1624
rect 1475 1623 1476 1627
rect 1470 1622 1476 1623
rect 1618 1627 1624 1628
rect 1618 1623 1619 1627
rect 1623 1626 1624 1627
rect 1774 1627 1780 1628
rect 1774 1626 1775 1627
rect 1623 1624 1775 1626
rect 1623 1623 1624 1624
rect 1618 1622 1624 1623
rect 1774 1623 1775 1624
rect 1779 1623 1780 1627
rect 1774 1622 1780 1623
rect 1094 1619 1100 1620
rect 1158 1620 1164 1621
rect 1134 1617 1140 1618
rect 174 1616 180 1617
rect 174 1612 175 1616
rect 179 1612 180 1616
rect 174 1611 180 1612
rect 214 1616 220 1617
rect 214 1612 215 1616
rect 219 1612 220 1616
rect 214 1611 220 1612
rect 254 1616 260 1617
rect 254 1612 255 1616
rect 259 1612 260 1616
rect 254 1611 260 1612
rect 302 1616 308 1617
rect 302 1612 303 1616
rect 307 1612 308 1616
rect 302 1611 308 1612
rect 358 1616 364 1617
rect 358 1612 359 1616
rect 363 1612 364 1616
rect 358 1611 364 1612
rect 406 1616 412 1617
rect 406 1612 407 1616
rect 411 1612 412 1616
rect 406 1611 412 1612
rect 454 1616 460 1617
rect 454 1612 455 1616
rect 459 1612 460 1616
rect 454 1611 460 1612
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 550 1616 556 1617
rect 550 1612 551 1616
rect 555 1612 556 1616
rect 550 1611 556 1612
rect 606 1616 612 1617
rect 606 1612 607 1616
rect 611 1612 612 1616
rect 606 1611 612 1612
rect 662 1616 668 1617
rect 662 1612 663 1616
rect 667 1612 668 1616
rect 662 1611 668 1612
rect 718 1616 724 1617
rect 718 1612 719 1616
rect 723 1612 724 1616
rect 1134 1613 1135 1617
rect 1139 1613 1140 1617
rect 1158 1616 1159 1620
rect 1163 1616 1164 1620
rect 1158 1615 1164 1616
rect 1198 1620 1204 1621
rect 1198 1616 1199 1620
rect 1203 1616 1204 1620
rect 1198 1615 1204 1616
rect 1246 1620 1252 1621
rect 1246 1616 1247 1620
rect 1251 1616 1252 1620
rect 1246 1615 1252 1616
rect 1318 1620 1324 1621
rect 1318 1616 1319 1620
rect 1323 1616 1324 1620
rect 1318 1615 1324 1616
rect 1390 1620 1396 1621
rect 1390 1616 1391 1620
rect 1395 1616 1396 1620
rect 1390 1615 1396 1616
rect 1462 1620 1468 1621
rect 1462 1616 1463 1620
rect 1467 1616 1468 1620
rect 1462 1615 1468 1616
rect 1534 1620 1540 1621
rect 1534 1616 1535 1620
rect 1539 1616 1540 1620
rect 1534 1615 1540 1616
rect 1606 1620 1612 1621
rect 1606 1616 1607 1620
rect 1611 1616 1612 1620
rect 1606 1615 1612 1616
rect 1678 1620 1684 1621
rect 1678 1616 1679 1620
rect 1683 1616 1684 1620
rect 1678 1615 1684 1616
rect 1750 1620 1756 1621
rect 1750 1616 1751 1620
rect 1755 1616 1756 1620
rect 1750 1615 1756 1616
rect 1830 1620 1836 1621
rect 1830 1616 1831 1620
rect 1835 1616 1836 1620
rect 1830 1615 1836 1616
rect 2118 1617 2124 1618
rect 1134 1612 1140 1613
rect 2118 1613 2119 1617
rect 2123 1613 2124 1617
rect 2118 1612 2124 1613
rect 718 1611 724 1612
rect 1186 1611 1192 1612
rect 1186 1607 1187 1611
rect 1191 1610 1192 1611
rect 1558 1611 1564 1612
rect 1191 1608 1322 1610
rect 1191 1607 1192 1608
rect 1186 1606 1192 1607
rect 166 1603 177 1604
rect 166 1599 167 1603
rect 171 1599 172 1603
rect 176 1599 177 1603
rect 166 1598 177 1599
rect 202 1603 208 1604
rect 202 1599 203 1603
rect 207 1602 208 1603
rect 211 1603 217 1604
rect 211 1602 212 1603
rect 207 1600 212 1602
rect 207 1599 208 1600
rect 202 1598 208 1599
rect 211 1599 212 1600
rect 216 1599 217 1603
rect 211 1598 217 1599
rect 242 1603 248 1604
rect 242 1599 243 1603
rect 247 1602 248 1603
rect 251 1603 257 1604
rect 251 1602 252 1603
rect 247 1600 252 1602
rect 247 1599 248 1600
rect 242 1598 248 1599
rect 251 1599 252 1600
rect 256 1599 257 1603
rect 251 1598 257 1599
rect 299 1603 305 1604
rect 299 1599 300 1603
rect 304 1602 305 1603
rect 330 1603 336 1604
rect 330 1602 331 1603
rect 304 1600 331 1602
rect 304 1599 305 1600
rect 299 1598 305 1599
rect 330 1599 331 1600
rect 335 1599 336 1603
rect 330 1598 336 1599
rect 355 1603 361 1604
rect 355 1599 356 1603
rect 360 1602 361 1603
rect 374 1603 380 1604
rect 374 1602 375 1603
rect 360 1600 375 1602
rect 360 1599 361 1600
rect 355 1598 361 1599
rect 374 1599 375 1600
rect 379 1599 380 1603
rect 374 1598 380 1599
rect 398 1603 409 1604
rect 398 1599 399 1603
rect 403 1599 404 1603
rect 408 1599 409 1603
rect 398 1598 409 1599
rect 451 1603 457 1604
rect 451 1599 452 1603
rect 456 1602 457 1603
rect 470 1603 476 1604
rect 470 1602 471 1603
rect 456 1600 471 1602
rect 456 1599 457 1600
rect 451 1598 457 1599
rect 470 1599 471 1600
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 494 1603 505 1604
rect 494 1599 495 1603
rect 499 1599 500 1603
rect 504 1599 505 1603
rect 494 1598 505 1599
rect 542 1603 553 1604
rect 542 1599 543 1603
rect 547 1599 548 1603
rect 552 1599 553 1603
rect 542 1598 553 1599
rect 598 1603 609 1604
rect 598 1599 599 1603
rect 603 1599 604 1603
rect 608 1599 609 1603
rect 598 1598 609 1599
rect 654 1603 665 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 664 1599 665 1603
rect 654 1598 665 1599
rect 710 1603 721 1604
rect 710 1599 711 1603
rect 715 1599 716 1603
rect 720 1599 721 1603
rect 1183 1603 1192 1604
rect 710 1598 721 1599
rect 1134 1600 1140 1601
rect 1134 1596 1135 1600
rect 1139 1596 1140 1600
rect 1183 1599 1184 1603
rect 1191 1599 1192 1603
rect 1183 1598 1192 1599
rect 1223 1603 1229 1604
rect 1223 1599 1224 1603
rect 1228 1602 1229 1603
rect 1231 1603 1237 1604
rect 1231 1602 1232 1603
rect 1228 1600 1232 1602
rect 1228 1599 1229 1600
rect 1223 1598 1229 1599
rect 1231 1599 1232 1600
rect 1236 1599 1237 1603
rect 1231 1598 1237 1599
rect 1271 1603 1277 1604
rect 1271 1599 1272 1603
rect 1276 1602 1277 1603
rect 1310 1603 1316 1604
rect 1310 1602 1311 1603
rect 1276 1600 1311 1602
rect 1276 1599 1277 1600
rect 1271 1598 1277 1599
rect 1310 1599 1311 1600
rect 1315 1599 1316 1603
rect 1320 1602 1322 1608
rect 1558 1607 1559 1611
rect 1563 1610 1564 1611
rect 1702 1611 1708 1612
rect 1563 1608 1642 1610
rect 1563 1607 1564 1608
rect 1558 1606 1564 1607
rect 1343 1603 1349 1604
rect 1343 1602 1344 1603
rect 1320 1600 1344 1602
rect 1310 1598 1316 1599
rect 1343 1599 1344 1600
rect 1348 1599 1349 1603
rect 1343 1598 1349 1599
rect 1415 1603 1421 1604
rect 1415 1599 1416 1603
rect 1420 1602 1421 1603
rect 1454 1603 1460 1604
rect 1454 1602 1455 1603
rect 1420 1600 1455 1602
rect 1420 1599 1421 1600
rect 1415 1598 1421 1599
rect 1454 1599 1455 1600
rect 1459 1599 1460 1603
rect 1454 1598 1460 1599
rect 1470 1603 1476 1604
rect 1470 1599 1471 1603
rect 1475 1602 1476 1603
rect 1487 1603 1493 1604
rect 1487 1602 1488 1603
rect 1475 1600 1488 1602
rect 1475 1599 1476 1600
rect 1470 1598 1476 1599
rect 1487 1599 1488 1600
rect 1492 1599 1493 1603
rect 1487 1598 1493 1599
rect 1559 1603 1565 1604
rect 1559 1599 1560 1603
rect 1564 1602 1565 1603
rect 1598 1603 1604 1604
rect 1598 1602 1599 1603
rect 1564 1600 1599 1602
rect 1564 1599 1565 1600
rect 1559 1598 1565 1599
rect 1598 1599 1599 1600
rect 1603 1599 1604 1603
rect 1598 1598 1604 1599
rect 1630 1603 1637 1604
rect 1630 1599 1631 1603
rect 1636 1599 1637 1603
rect 1640 1602 1642 1608
rect 1702 1607 1703 1611
rect 1707 1610 1708 1611
rect 1707 1608 1834 1610
rect 1707 1607 1708 1608
rect 1702 1606 1708 1607
rect 1703 1603 1709 1604
rect 1703 1602 1704 1603
rect 1640 1600 1704 1602
rect 1630 1598 1637 1599
rect 1703 1599 1704 1600
rect 1708 1599 1709 1603
rect 1703 1598 1709 1599
rect 1775 1603 1781 1604
rect 1775 1599 1776 1603
rect 1780 1602 1781 1603
rect 1822 1603 1828 1604
rect 1822 1602 1823 1603
rect 1780 1600 1823 1602
rect 1780 1599 1781 1600
rect 1775 1598 1781 1599
rect 1822 1599 1823 1600
rect 1827 1599 1828 1603
rect 1832 1602 1834 1608
rect 1855 1603 1861 1604
rect 1855 1602 1856 1603
rect 1832 1600 1856 1602
rect 1822 1598 1828 1599
rect 1855 1599 1856 1600
rect 1860 1599 1861 1603
rect 1855 1598 1861 1599
rect 2118 1600 2124 1601
rect 1134 1595 1140 1596
rect 2118 1596 2119 1600
rect 2123 1596 2124 1600
rect 2118 1595 2124 1596
rect 1158 1592 1164 1593
rect 558 1591 564 1592
rect 558 1590 559 1591
rect 476 1588 559 1590
rect 476 1586 478 1588
rect 558 1587 559 1588
rect 563 1587 564 1591
rect 1158 1588 1159 1592
rect 1163 1588 1164 1592
rect 1158 1587 1164 1588
rect 1198 1592 1204 1593
rect 1198 1588 1199 1592
rect 1203 1588 1204 1592
rect 1198 1587 1204 1588
rect 1246 1592 1252 1593
rect 1246 1588 1247 1592
rect 1251 1588 1252 1592
rect 1246 1587 1252 1588
rect 1318 1592 1324 1593
rect 1318 1588 1319 1592
rect 1323 1588 1324 1592
rect 1318 1587 1324 1588
rect 1390 1592 1396 1593
rect 1390 1588 1391 1592
rect 1395 1588 1396 1592
rect 1390 1587 1396 1588
rect 1462 1592 1468 1593
rect 1462 1588 1463 1592
rect 1467 1588 1468 1592
rect 1462 1587 1468 1588
rect 1534 1592 1540 1593
rect 1534 1588 1535 1592
rect 1539 1588 1540 1592
rect 1534 1587 1540 1588
rect 1606 1592 1612 1593
rect 1606 1588 1607 1592
rect 1611 1588 1612 1592
rect 1606 1587 1612 1588
rect 1678 1592 1684 1593
rect 1678 1588 1679 1592
rect 1683 1588 1684 1592
rect 1678 1587 1684 1588
rect 1750 1592 1756 1593
rect 1750 1588 1751 1592
rect 1755 1588 1756 1592
rect 1750 1587 1756 1588
rect 1830 1592 1836 1593
rect 1830 1588 1831 1592
rect 1835 1588 1836 1592
rect 1830 1587 1836 1588
rect 558 1586 564 1587
rect 475 1585 481 1586
rect 139 1583 145 1584
rect 139 1579 140 1583
rect 144 1582 145 1583
rect 179 1583 185 1584
rect 144 1580 174 1582
rect 144 1579 145 1580
rect 139 1578 145 1579
rect 142 1572 148 1573
rect 142 1568 143 1572
rect 147 1568 148 1572
rect 142 1567 148 1568
rect 172 1566 174 1580
rect 179 1579 180 1583
rect 184 1582 185 1583
rect 215 1583 221 1584
rect 215 1582 216 1583
rect 184 1580 216 1582
rect 184 1579 185 1580
rect 179 1578 185 1579
rect 215 1579 216 1580
rect 220 1579 221 1583
rect 215 1578 221 1579
rect 227 1583 233 1584
rect 227 1579 228 1583
rect 232 1582 233 1583
rect 270 1583 276 1584
rect 270 1582 271 1583
rect 232 1580 271 1582
rect 232 1579 233 1580
rect 227 1578 233 1579
rect 270 1579 271 1580
rect 275 1579 276 1583
rect 270 1578 276 1579
rect 278 1583 289 1584
rect 278 1579 279 1583
rect 283 1579 284 1583
rect 288 1579 289 1583
rect 278 1578 289 1579
rect 347 1583 353 1584
rect 347 1579 348 1583
rect 352 1582 353 1583
rect 399 1583 405 1584
rect 399 1582 400 1583
rect 352 1580 400 1582
rect 352 1579 353 1580
rect 347 1578 353 1579
rect 399 1579 400 1580
rect 404 1579 405 1583
rect 399 1578 405 1579
rect 411 1583 417 1584
rect 411 1579 412 1583
rect 416 1582 417 1583
rect 466 1583 472 1584
rect 466 1582 467 1583
rect 416 1580 467 1582
rect 416 1579 417 1580
rect 411 1578 417 1579
rect 466 1579 467 1580
rect 471 1579 472 1583
rect 475 1581 476 1585
rect 480 1581 481 1585
rect 475 1580 481 1581
rect 534 1583 545 1584
rect 466 1578 472 1579
rect 534 1579 535 1583
rect 539 1579 540 1583
rect 544 1579 545 1583
rect 534 1578 545 1579
rect 570 1583 576 1584
rect 570 1579 571 1583
rect 575 1582 576 1583
rect 603 1583 609 1584
rect 603 1582 604 1583
rect 575 1580 604 1582
rect 575 1579 576 1580
rect 570 1578 576 1579
rect 603 1579 604 1580
rect 608 1579 609 1583
rect 603 1578 609 1579
rect 634 1583 640 1584
rect 634 1579 635 1583
rect 639 1582 640 1583
rect 659 1583 665 1584
rect 659 1582 660 1583
rect 639 1580 660 1582
rect 639 1579 640 1580
rect 634 1578 640 1579
rect 659 1579 660 1580
rect 664 1579 665 1583
rect 659 1578 665 1579
rect 690 1583 696 1584
rect 690 1579 691 1583
rect 695 1582 696 1583
rect 723 1583 729 1584
rect 723 1582 724 1583
rect 695 1580 724 1582
rect 695 1579 696 1580
rect 690 1578 696 1579
rect 723 1579 724 1580
rect 728 1579 729 1583
rect 723 1578 729 1579
rect 754 1583 760 1584
rect 754 1579 755 1583
rect 759 1582 760 1583
rect 787 1583 793 1584
rect 787 1582 788 1583
rect 759 1580 788 1582
rect 759 1579 760 1580
rect 754 1578 760 1579
rect 787 1579 788 1580
rect 792 1579 793 1583
rect 787 1578 793 1579
rect 818 1583 824 1584
rect 818 1579 819 1583
rect 823 1582 824 1583
rect 851 1583 857 1584
rect 851 1582 852 1583
rect 823 1580 852 1582
rect 823 1579 824 1580
rect 818 1578 824 1579
rect 851 1579 852 1580
rect 856 1579 857 1583
rect 851 1578 857 1579
rect 1155 1579 1161 1580
rect 1155 1575 1156 1579
rect 1160 1578 1161 1579
rect 1178 1579 1184 1580
rect 1178 1578 1179 1579
rect 1160 1576 1179 1578
rect 1160 1575 1161 1576
rect 1155 1574 1161 1575
rect 1178 1575 1179 1576
rect 1183 1575 1184 1579
rect 1178 1574 1184 1575
rect 1186 1579 1192 1580
rect 1186 1575 1187 1579
rect 1191 1578 1192 1579
rect 1195 1579 1201 1580
rect 1195 1578 1196 1579
rect 1191 1576 1196 1578
rect 1191 1575 1192 1576
rect 1186 1574 1192 1575
rect 1195 1575 1196 1576
rect 1200 1575 1201 1579
rect 1195 1574 1201 1575
rect 1231 1579 1237 1580
rect 1231 1575 1232 1579
rect 1236 1578 1237 1579
rect 1243 1579 1249 1580
rect 1243 1578 1244 1579
rect 1236 1576 1244 1578
rect 1236 1575 1237 1576
rect 1231 1574 1237 1575
rect 1243 1575 1244 1576
rect 1248 1575 1249 1579
rect 1243 1574 1249 1575
rect 1310 1579 1321 1580
rect 1310 1575 1311 1579
rect 1315 1575 1316 1579
rect 1320 1575 1321 1579
rect 1310 1574 1321 1575
rect 1354 1579 1360 1580
rect 1354 1575 1355 1579
rect 1359 1578 1360 1579
rect 1387 1579 1393 1580
rect 1387 1578 1388 1579
rect 1359 1576 1388 1578
rect 1359 1575 1360 1576
rect 1354 1574 1360 1575
rect 1387 1575 1388 1576
rect 1392 1575 1393 1579
rect 1387 1574 1393 1575
rect 1454 1579 1465 1580
rect 1454 1575 1455 1579
rect 1459 1575 1460 1579
rect 1464 1575 1465 1579
rect 1454 1574 1465 1575
rect 1531 1579 1537 1580
rect 1531 1575 1532 1579
rect 1536 1578 1537 1579
rect 1558 1579 1564 1580
rect 1558 1578 1559 1579
rect 1536 1576 1559 1578
rect 1536 1575 1537 1576
rect 1531 1574 1537 1575
rect 1558 1575 1559 1576
rect 1563 1575 1564 1579
rect 1558 1574 1564 1575
rect 1598 1579 1609 1580
rect 1598 1575 1599 1579
rect 1603 1575 1604 1579
rect 1608 1575 1609 1579
rect 1598 1574 1609 1575
rect 1675 1579 1681 1580
rect 1675 1575 1676 1579
rect 1680 1578 1681 1579
rect 1702 1579 1708 1580
rect 1702 1578 1703 1579
rect 1680 1576 1703 1578
rect 1680 1575 1681 1576
rect 1675 1574 1681 1575
rect 1702 1575 1703 1576
rect 1707 1575 1708 1579
rect 1702 1574 1708 1575
rect 1742 1579 1753 1580
rect 1742 1575 1743 1579
rect 1747 1575 1748 1579
rect 1752 1575 1753 1579
rect 1742 1574 1753 1575
rect 1822 1579 1833 1580
rect 1822 1575 1823 1579
rect 1827 1575 1828 1579
rect 1832 1575 1833 1579
rect 1822 1574 1833 1575
rect 182 1572 188 1573
rect 182 1568 183 1572
rect 187 1568 188 1572
rect 182 1567 188 1568
rect 230 1572 236 1573
rect 230 1568 231 1572
rect 235 1568 236 1572
rect 230 1567 236 1568
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 350 1572 356 1573
rect 350 1568 351 1572
rect 355 1568 356 1572
rect 350 1567 356 1568
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 478 1572 484 1573
rect 478 1568 479 1572
rect 483 1568 484 1572
rect 478 1567 484 1568
rect 542 1572 548 1573
rect 542 1568 543 1572
rect 547 1568 548 1572
rect 542 1567 548 1568
rect 606 1572 612 1573
rect 606 1568 607 1572
rect 611 1568 612 1572
rect 606 1567 612 1568
rect 662 1572 668 1573
rect 662 1568 663 1572
rect 667 1568 668 1572
rect 662 1567 668 1568
rect 726 1572 732 1573
rect 726 1568 727 1572
rect 731 1568 732 1572
rect 726 1567 732 1568
rect 790 1572 796 1573
rect 790 1568 791 1572
rect 795 1568 796 1572
rect 790 1567 796 1568
rect 854 1572 860 1573
rect 854 1568 855 1572
rect 859 1568 860 1572
rect 1469 1572 1527 1574
rect 1469 1570 1471 1572
rect 1525 1570 1527 1572
rect 1554 1571 1560 1572
rect 1554 1570 1555 1571
rect 1467 1569 1473 1570
rect 854 1567 860 1568
rect 1235 1567 1241 1568
rect 110 1564 116 1565
rect 172 1564 178 1566
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 110 1559 116 1560
rect 150 1559 156 1560
rect 150 1555 151 1559
rect 155 1558 156 1559
rect 167 1559 173 1560
rect 167 1558 168 1559
rect 155 1556 168 1558
rect 155 1555 156 1556
rect 150 1554 156 1555
rect 167 1555 168 1556
rect 172 1555 173 1559
rect 176 1558 178 1564
rect 1094 1564 1100 1565
rect 1094 1560 1095 1564
rect 1099 1560 1100 1564
rect 1235 1563 1236 1567
rect 1240 1566 1241 1567
rect 1258 1567 1264 1568
rect 1258 1566 1259 1567
rect 1240 1564 1259 1566
rect 1240 1563 1241 1564
rect 1235 1562 1241 1563
rect 1258 1563 1259 1564
rect 1263 1563 1264 1567
rect 1258 1562 1264 1563
rect 1266 1567 1272 1568
rect 1266 1563 1267 1567
rect 1271 1566 1272 1567
rect 1275 1567 1281 1568
rect 1275 1566 1276 1567
rect 1271 1564 1276 1566
rect 1271 1563 1272 1564
rect 1266 1562 1272 1563
rect 1275 1563 1276 1564
rect 1280 1563 1281 1567
rect 1275 1562 1281 1563
rect 1306 1567 1312 1568
rect 1306 1563 1307 1567
rect 1311 1566 1312 1567
rect 1323 1567 1329 1568
rect 1323 1566 1324 1567
rect 1311 1564 1324 1566
rect 1311 1563 1312 1564
rect 1306 1562 1312 1563
rect 1323 1563 1324 1564
rect 1328 1563 1329 1567
rect 1323 1562 1329 1563
rect 1371 1567 1377 1568
rect 1371 1563 1372 1567
rect 1376 1566 1377 1567
rect 1410 1567 1416 1568
rect 1410 1566 1411 1567
rect 1376 1564 1411 1566
rect 1376 1563 1377 1564
rect 1371 1562 1377 1563
rect 1410 1563 1411 1564
rect 1415 1563 1416 1567
rect 1410 1562 1416 1563
rect 1419 1567 1425 1568
rect 1419 1563 1420 1567
rect 1424 1566 1425 1567
rect 1430 1567 1436 1568
rect 1430 1566 1431 1567
rect 1424 1564 1431 1566
rect 1424 1563 1425 1564
rect 1419 1562 1425 1563
rect 1430 1563 1431 1564
rect 1435 1563 1436 1567
rect 1467 1565 1468 1569
rect 1472 1565 1473 1569
rect 1525 1568 1555 1570
rect 1467 1564 1473 1565
rect 1498 1567 1504 1568
rect 1430 1562 1436 1563
rect 1498 1563 1499 1567
rect 1503 1566 1504 1567
rect 1515 1567 1521 1568
rect 1515 1566 1516 1567
rect 1503 1564 1516 1566
rect 1503 1563 1504 1564
rect 1498 1562 1504 1563
rect 1515 1563 1516 1564
rect 1520 1563 1521 1567
rect 1554 1567 1555 1568
rect 1559 1567 1560 1571
rect 1554 1566 1560 1567
rect 1563 1567 1569 1568
rect 1515 1562 1521 1563
rect 1563 1563 1564 1567
rect 1568 1566 1569 1567
rect 1607 1567 1613 1568
rect 1607 1566 1608 1567
rect 1568 1564 1608 1566
rect 1568 1563 1569 1564
rect 1563 1562 1569 1563
rect 1607 1563 1608 1564
rect 1612 1563 1613 1567
rect 1607 1562 1613 1563
rect 1619 1567 1625 1568
rect 1619 1563 1620 1567
rect 1624 1566 1625 1567
rect 1630 1567 1636 1568
rect 1630 1566 1631 1567
rect 1624 1564 1631 1566
rect 1624 1563 1625 1564
rect 1619 1562 1625 1563
rect 1630 1563 1631 1564
rect 1635 1563 1636 1567
rect 1630 1562 1636 1563
rect 1650 1567 1656 1568
rect 1650 1563 1651 1567
rect 1655 1566 1656 1567
rect 1675 1567 1681 1568
rect 1675 1566 1676 1567
rect 1655 1564 1676 1566
rect 1655 1563 1656 1564
rect 1650 1562 1656 1563
rect 1675 1563 1676 1564
rect 1680 1563 1681 1567
rect 1675 1562 1681 1563
rect 1706 1567 1712 1568
rect 1706 1563 1707 1567
rect 1711 1566 1712 1567
rect 1731 1567 1737 1568
rect 1731 1566 1732 1567
rect 1711 1564 1732 1566
rect 1711 1563 1712 1564
rect 1706 1562 1712 1563
rect 1731 1563 1732 1564
rect 1736 1563 1737 1567
rect 1731 1562 1737 1563
rect 207 1559 213 1560
rect 207 1558 208 1559
rect 176 1556 208 1558
rect 167 1554 173 1555
rect 207 1555 208 1556
rect 212 1555 213 1559
rect 207 1554 213 1555
rect 215 1559 221 1560
rect 215 1555 216 1559
rect 220 1558 221 1559
rect 255 1559 261 1560
rect 255 1558 256 1559
rect 220 1556 256 1558
rect 220 1555 221 1556
rect 215 1554 221 1555
rect 255 1555 256 1556
rect 260 1555 261 1559
rect 255 1554 261 1555
rect 270 1559 276 1560
rect 270 1555 271 1559
rect 275 1558 276 1559
rect 311 1559 317 1560
rect 311 1558 312 1559
rect 275 1556 312 1558
rect 275 1555 276 1556
rect 270 1554 276 1555
rect 311 1555 312 1556
rect 316 1555 317 1559
rect 311 1554 317 1555
rect 374 1559 381 1560
rect 374 1555 375 1559
rect 380 1555 381 1559
rect 374 1554 381 1555
rect 399 1559 405 1560
rect 399 1555 400 1559
rect 404 1558 405 1559
rect 439 1559 445 1560
rect 439 1558 440 1559
rect 404 1556 440 1558
rect 404 1555 405 1556
rect 399 1554 405 1555
rect 439 1555 440 1556
rect 444 1555 445 1559
rect 439 1554 445 1555
rect 466 1559 472 1560
rect 466 1555 467 1559
rect 471 1558 472 1559
rect 503 1559 509 1560
rect 503 1558 504 1559
rect 471 1556 504 1558
rect 471 1555 472 1556
rect 466 1554 472 1555
rect 503 1555 504 1556
rect 508 1555 509 1559
rect 503 1554 509 1555
rect 567 1559 576 1560
rect 567 1555 568 1559
rect 575 1555 576 1559
rect 567 1554 576 1555
rect 631 1559 640 1560
rect 631 1555 632 1559
rect 639 1555 640 1559
rect 631 1554 640 1555
rect 687 1559 696 1560
rect 687 1555 688 1559
rect 695 1555 696 1559
rect 687 1554 696 1555
rect 751 1559 760 1560
rect 751 1555 752 1559
rect 759 1555 760 1559
rect 751 1554 760 1555
rect 815 1559 824 1560
rect 815 1555 816 1559
rect 823 1555 824 1559
rect 815 1554 824 1555
rect 838 1559 844 1560
rect 838 1555 839 1559
rect 843 1558 844 1559
rect 879 1559 885 1560
rect 1094 1559 1100 1560
rect 879 1558 880 1559
rect 843 1556 880 1558
rect 843 1555 844 1556
rect 838 1554 844 1555
rect 879 1555 880 1556
rect 884 1555 885 1559
rect 879 1554 885 1555
rect 1238 1556 1244 1557
rect 1238 1552 1239 1556
rect 1243 1552 1244 1556
rect 1238 1551 1244 1552
rect 1278 1556 1284 1557
rect 1278 1552 1279 1556
rect 1283 1552 1284 1556
rect 1278 1551 1284 1552
rect 1326 1556 1332 1557
rect 1326 1552 1327 1556
rect 1331 1552 1332 1556
rect 1326 1551 1332 1552
rect 1374 1556 1380 1557
rect 1374 1552 1375 1556
rect 1379 1552 1380 1556
rect 1374 1551 1380 1552
rect 1422 1556 1428 1557
rect 1422 1552 1423 1556
rect 1427 1552 1428 1556
rect 1422 1551 1428 1552
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1518 1556 1524 1557
rect 1518 1552 1519 1556
rect 1523 1552 1524 1556
rect 1518 1551 1524 1552
rect 1566 1556 1572 1557
rect 1566 1552 1567 1556
rect 1571 1552 1572 1556
rect 1566 1551 1572 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1678 1556 1684 1557
rect 1678 1552 1679 1556
rect 1683 1552 1684 1556
rect 1678 1551 1684 1552
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 1134 1548 1140 1549
rect 1640 1548 1674 1550
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 1094 1547 1100 1548
rect 110 1542 116 1543
rect 142 1544 148 1545
rect 142 1540 143 1544
rect 147 1540 148 1544
rect 142 1539 148 1540
rect 182 1544 188 1545
rect 182 1540 183 1544
rect 187 1540 188 1544
rect 182 1539 188 1540
rect 230 1544 236 1545
rect 230 1540 231 1544
rect 235 1540 236 1544
rect 230 1539 236 1540
rect 286 1544 292 1545
rect 286 1540 287 1544
rect 291 1540 292 1544
rect 286 1539 292 1540
rect 350 1544 356 1545
rect 350 1540 351 1544
rect 355 1540 356 1544
rect 350 1539 356 1540
rect 414 1544 420 1545
rect 414 1540 415 1544
rect 419 1540 420 1544
rect 414 1539 420 1540
rect 478 1544 484 1545
rect 478 1540 479 1544
rect 483 1540 484 1544
rect 478 1539 484 1540
rect 542 1544 548 1545
rect 542 1540 543 1544
rect 547 1540 548 1544
rect 542 1539 548 1540
rect 606 1544 612 1545
rect 606 1540 607 1544
rect 611 1540 612 1544
rect 606 1539 612 1540
rect 662 1544 668 1545
rect 662 1540 663 1544
rect 667 1540 668 1544
rect 662 1539 668 1540
rect 726 1544 732 1545
rect 726 1540 727 1544
rect 731 1540 732 1544
rect 726 1539 732 1540
rect 790 1544 796 1545
rect 790 1540 791 1544
rect 795 1540 796 1544
rect 790 1539 796 1540
rect 854 1544 860 1545
rect 854 1540 855 1544
rect 859 1540 860 1544
rect 1094 1543 1095 1547
rect 1099 1543 1100 1547
rect 1134 1544 1135 1548
rect 1139 1544 1140 1548
rect 1607 1547 1613 1548
rect 1134 1543 1140 1544
rect 1263 1543 1272 1544
rect 1094 1542 1100 1543
rect 854 1539 860 1540
rect 1263 1539 1264 1543
rect 1271 1539 1272 1543
rect 1263 1538 1272 1539
rect 1303 1543 1312 1544
rect 1303 1539 1304 1543
rect 1311 1539 1312 1543
rect 1303 1538 1312 1539
rect 1351 1543 1360 1544
rect 1351 1539 1352 1543
rect 1359 1539 1360 1543
rect 1351 1538 1360 1539
rect 1398 1543 1405 1544
rect 1398 1539 1399 1543
rect 1404 1539 1405 1543
rect 1398 1538 1405 1539
rect 1410 1543 1416 1544
rect 1410 1539 1411 1543
rect 1415 1542 1416 1543
rect 1447 1543 1453 1544
rect 1447 1542 1448 1543
rect 1415 1540 1448 1542
rect 1415 1539 1416 1540
rect 1410 1538 1416 1539
rect 1447 1539 1448 1540
rect 1452 1539 1453 1543
rect 1447 1538 1453 1539
rect 1495 1543 1504 1544
rect 1495 1539 1496 1543
rect 1503 1539 1504 1543
rect 1495 1538 1504 1539
rect 1543 1543 1552 1544
rect 1543 1539 1544 1543
rect 1551 1539 1552 1543
rect 1543 1538 1552 1539
rect 1554 1543 1560 1544
rect 1554 1539 1555 1543
rect 1559 1542 1560 1543
rect 1591 1543 1597 1544
rect 1591 1542 1592 1543
rect 1559 1540 1592 1542
rect 1559 1539 1560 1540
rect 1554 1538 1560 1539
rect 1591 1539 1592 1540
rect 1596 1539 1597 1543
rect 1607 1543 1608 1547
rect 1612 1546 1613 1547
rect 1640 1546 1642 1548
rect 1612 1544 1642 1546
rect 1672 1546 1674 1548
rect 1696 1548 1718 1550
rect 1696 1546 1698 1548
rect 1672 1544 1698 1546
rect 1612 1543 1613 1544
rect 1607 1542 1613 1543
rect 1647 1543 1656 1544
rect 1591 1538 1597 1539
rect 1647 1539 1648 1543
rect 1655 1539 1656 1543
rect 1647 1538 1656 1539
rect 1703 1543 1712 1544
rect 1703 1539 1704 1543
rect 1711 1539 1712 1543
rect 1716 1542 1718 1548
rect 2118 1548 2124 1549
rect 2118 1544 2119 1548
rect 2123 1544 2124 1548
rect 1759 1543 1765 1544
rect 2118 1543 2124 1544
rect 1759 1542 1760 1543
rect 1716 1540 1760 1542
rect 1703 1538 1712 1539
rect 1759 1539 1760 1540
rect 1764 1539 1765 1543
rect 1759 1538 1765 1539
rect 1134 1531 1140 1532
rect 1134 1527 1135 1531
rect 1139 1527 1140 1531
rect 2118 1531 2124 1532
rect 1134 1526 1140 1527
rect 1238 1528 1244 1529
rect 134 1524 140 1525
rect 110 1521 116 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 134 1520 135 1524
rect 139 1520 140 1524
rect 134 1519 140 1520
rect 174 1524 180 1525
rect 174 1520 175 1524
rect 179 1520 180 1524
rect 174 1519 180 1520
rect 214 1524 220 1525
rect 214 1520 215 1524
rect 219 1520 220 1524
rect 214 1519 220 1520
rect 254 1524 260 1525
rect 254 1520 255 1524
rect 259 1520 260 1524
rect 254 1519 260 1520
rect 294 1524 300 1525
rect 294 1520 295 1524
rect 299 1520 300 1524
rect 294 1519 300 1520
rect 334 1524 340 1525
rect 334 1520 335 1524
rect 339 1520 340 1524
rect 334 1519 340 1520
rect 374 1524 380 1525
rect 374 1520 375 1524
rect 379 1520 380 1524
rect 374 1519 380 1520
rect 414 1524 420 1525
rect 414 1520 415 1524
rect 419 1520 420 1524
rect 414 1519 420 1520
rect 454 1524 460 1525
rect 454 1520 455 1524
rect 459 1520 460 1524
rect 454 1519 460 1520
rect 494 1524 500 1525
rect 494 1520 495 1524
rect 499 1520 500 1524
rect 494 1519 500 1520
rect 534 1524 540 1525
rect 534 1520 535 1524
rect 539 1520 540 1524
rect 534 1519 540 1520
rect 574 1524 580 1525
rect 574 1520 575 1524
rect 579 1520 580 1524
rect 574 1519 580 1520
rect 614 1524 620 1525
rect 614 1520 615 1524
rect 619 1520 620 1524
rect 614 1519 620 1520
rect 654 1524 660 1525
rect 654 1520 655 1524
rect 659 1520 660 1524
rect 654 1519 660 1520
rect 694 1524 700 1525
rect 694 1520 695 1524
rect 699 1520 700 1524
rect 694 1519 700 1520
rect 734 1524 740 1525
rect 734 1520 735 1524
rect 739 1520 740 1524
rect 734 1519 740 1520
rect 774 1524 780 1525
rect 774 1520 775 1524
rect 779 1520 780 1524
rect 774 1519 780 1520
rect 830 1524 836 1525
rect 830 1520 831 1524
rect 835 1520 836 1524
rect 830 1519 836 1520
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1238 1523 1244 1524
rect 1278 1528 1284 1529
rect 1278 1524 1279 1528
rect 1283 1524 1284 1528
rect 1278 1523 1284 1524
rect 1326 1528 1332 1529
rect 1326 1524 1327 1528
rect 1331 1524 1332 1528
rect 1326 1523 1332 1524
rect 1374 1528 1380 1529
rect 1374 1524 1375 1528
rect 1379 1524 1380 1528
rect 1374 1523 1380 1524
rect 1422 1528 1428 1529
rect 1422 1524 1423 1528
rect 1427 1524 1428 1528
rect 1422 1523 1428 1524
rect 1470 1528 1476 1529
rect 1470 1524 1471 1528
rect 1475 1524 1476 1528
rect 1470 1523 1476 1524
rect 1518 1528 1524 1529
rect 1518 1524 1519 1528
rect 1523 1524 1524 1528
rect 1518 1523 1524 1524
rect 1566 1528 1572 1529
rect 1566 1524 1567 1528
rect 1571 1524 1572 1528
rect 1566 1523 1572 1524
rect 1622 1528 1628 1529
rect 1622 1524 1623 1528
rect 1627 1524 1628 1528
rect 1622 1523 1628 1524
rect 1678 1528 1684 1529
rect 1678 1524 1679 1528
rect 1683 1524 1684 1528
rect 1678 1523 1684 1524
rect 1734 1528 1740 1529
rect 1734 1524 1735 1528
rect 1739 1524 1740 1528
rect 2118 1527 2119 1531
rect 2123 1527 2124 1531
rect 2118 1526 2124 1527
rect 1734 1523 1740 1524
rect 886 1519 892 1520
rect 1094 1521 1100 1522
rect 110 1516 116 1517
rect 1094 1517 1095 1521
rect 1099 1517 1100 1521
rect 1094 1516 1100 1517
rect 1318 1512 1324 1513
rect 1134 1509 1140 1510
rect 159 1507 168 1508
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 159 1503 160 1507
rect 167 1503 168 1507
rect 159 1502 168 1503
rect 199 1507 208 1508
rect 199 1503 200 1507
rect 207 1503 208 1507
rect 199 1502 208 1503
rect 239 1507 248 1508
rect 239 1503 240 1507
rect 247 1503 248 1507
rect 239 1502 248 1503
rect 279 1507 288 1508
rect 279 1503 280 1507
rect 287 1503 288 1507
rect 279 1502 288 1503
rect 319 1507 328 1508
rect 319 1503 320 1507
rect 327 1503 328 1507
rect 319 1502 328 1503
rect 359 1507 368 1508
rect 359 1503 360 1507
rect 367 1503 368 1507
rect 359 1502 368 1503
rect 399 1507 408 1508
rect 399 1503 400 1507
rect 407 1503 408 1507
rect 399 1502 408 1503
rect 439 1507 448 1508
rect 439 1503 440 1507
rect 447 1503 448 1507
rect 439 1502 448 1503
rect 479 1507 488 1508
rect 479 1503 480 1507
rect 487 1503 488 1507
rect 479 1502 488 1503
rect 519 1507 528 1508
rect 519 1503 520 1507
rect 527 1503 528 1507
rect 519 1502 528 1503
rect 558 1507 565 1508
rect 558 1503 559 1507
rect 564 1503 565 1507
rect 558 1502 565 1503
rect 599 1507 608 1508
rect 599 1503 600 1507
rect 607 1503 608 1507
rect 599 1502 608 1503
rect 639 1507 648 1508
rect 639 1503 640 1507
rect 647 1503 648 1507
rect 639 1502 648 1503
rect 679 1507 688 1508
rect 679 1503 680 1507
rect 687 1503 688 1507
rect 679 1502 688 1503
rect 719 1507 728 1508
rect 719 1503 720 1507
rect 727 1503 728 1507
rect 719 1502 728 1503
rect 759 1507 768 1508
rect 759 1503 760 1507
rect 767 1503 768 1507
rect 759 1502 768 1503
rect 782 1507 788 1508
rect 782 1503 783 1507
rect 787 1506 788 1507
rect 799 1507 805 1508
rect 799 1506 800 1507
rect 787 1504 800 1506
rect 787 1503 788 1504
rect 782 1502 788 1503
rect 799 1503 800 1504
rect 804 1503 805 1507
rect 799 1502 805 1503
rect 855 1507 861 1508
rect 855 1503 856 1507
rect 860 1506 861 1507
rect 878 1507 884 1508
rect 878 1506 879 1507
rect 860 1504 879 1506
rect 860 1503 861 1504
rect 855 1502 861 1503
rect 878 1503 879 1504
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 911 1507 917 1508
rect 911 1503 912 1507
rect 916 1506 917 1507
rect 926 1507 932 1508
rect 926 1506 927 1507
rect 916 1504 927 1506
rect 916 1503 917 1504
rect 911 1502 917 1503
rect 926 1503 927 1504
rect 931 1503 932 1507
rect 1134 1505 1135 1509
rect 1139 1505 1140 1509
rect 1318 1508 1319 1512
rect 1323 1508 1324 1512
rect 1318 1507 1324 1508
rect 1358 1512 1364 1513
rect 1358 1508 1359 1512
rect 1363 1508 1364 1512
rect 1358 1507 1364 1508
rect 1398 1512 1404 1513
rect 1398 1508 1399 1512
rect 1403 1508 1404 1512
rect 1398 1507 1404 1508
rect 1438 1512 1444 1513
rect 1438 1508 1439 1512
rect 1443 1508 1444 1512
rect 1438 1507 1444 1508
rect 1478 1512 1484 1513
rect 1478 1508 1479 1512
rect 1483 1508 1484 1512
rect 1478 1507 1484 1508
rect 1518 1512 1524 1513
rect 1518 1508 1519 1512
rect 1523 1508 1524 1512
rect 1518 1507 1524 1508
rect 1558 1512 1564 1513
rect 1558 1508 1559 1512
rect 1563 1508 1564 1512
rect 1558 1507 1564 1508
rect 1606 1512 1612 1513
rect 1606 1508 1607 1512
rect 1611 1508 1612 1512
rect 1606 1507 1612 1508
rect 1662 1512 1668 1513
rect 1662 1508 1663 1512
rect 1667 1508 1668 1512
rect 1662 1507 1668 1508
rect 1734 1512 1740 1513
rect 1734 1508 1735 1512
rect 1739 1508 1740 1512
rect 1734 1507 1740 1508
rect 1814 1512 1820 1513
rect 1814 1508 1815 1512
rect 1819 1508 1820 1512
rect 1814 1507 1820 1508
rect 1902 1512 1908 1513
rect 1902 1508 1903 1512
rect 1907 1508 1908 1512
rect 1902 1507 1908 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2070 1512 2076 1513
rect 2070 1508 2071 1512
rect 2075 1508 2076 1512
rect 2070 1507 2076 1508
rect 2118 1509 2124 1510
rect 926 1502 932 1503
rect 1094 1504 1100 1505
rect 1134 1504 1140 1505
rect 2118 1505 2119 1509
rect 2123 1505 2124 1509
rect 2118 1504 2124 1505
rect 110 1499 116 1500
rect 1094 1500 1095 1504
rect 1099 1500 1100 1504
rect 1094 1499 1100 1500
rect 1430 1503 1436 1504
rect 1430 1499 1431 1503
rect 1435 1502 1436 1503
rect 1435 1500 1518 1502
rect 1435 1499 1436 1500
rect 1430 1498 1436 1499
rect 134 1496 140 1497
rect 134 1492 135 1496
rect 139 1492 140 1496
rect 134 1491 140 1492
rect 174 1496 180 1497
rect 174 1492 175 1496
rect 179 1492 180 1496
rect 174 1491 180 1492
rect 214 1496 220 1497
rect 214 1492 215 1496
rect 219 1492 220 1496
rect 214 1491 220 1492
rect 254 1496 260 1497
rect 254 1492 255 1496
rect 259 1492 260 1496
rect 254 1491 260 1492
rect 294 1496 300 1497
rect 294 1492 295 1496
rect 299 1492 300 1496
rect 294 1491 300 1492
rect 334 1496 340 1497
rect 334 1492 335 1496
rect 339 1492 340 1496
rect 334 1491 340 1492
rect 374 1496 380 1497
rect 374 1492 375 1496
rect 379 1492 380 1496
rect 374 1491 380 1492
rect 414 1496 420 1497
rect 414 1492 415 1496
rect 419 1492 420 1496
rect 414 1491 420 1492
rect 454 1496 460 1497
rect 454 1492 455 1496
rect 459 1492 460 1496
rect 454 1491 460 1492
rect 494 1496 500 1497
rect 494 1492 495 1496
rect 499 1492 500 1496
rect 494 1491 500 1492
rect 534 1496 540 1497
rect 534 1492 535 1496
rect 539 1492 540 1496
rect 534 1491 540 1492
rect 574 1496 580 1497
rect 574 1492 575 1496
rect 579 1492 580 1496
rect 574 1491 580 1492
rect 614 1496 620 1497
rect 614 1492 615 1496
rect 619 1492 620 1496
rect 614 1491 620 1492
rect 654 1496 660 1497
rect 654 1492 655 1496
rect 659 1492 660 1496
rect 654 1491 660 1492
rect 694 1496 700 1497
rect 694 1492 695 1496
rect 699 1492 700 1496
rect 694 1491 700 1492
rect 734 1496 740 1497
rect 734 1492 735 1496
rect 739 1492 740 1496
rect 734 1491 740 1492
rect 774 1496 780 1497
rect 774 1492 775 1496
rect 779 1492 780 1496
rect 774 1491 780 1492
rect 830 1496 836 1497
rect 830 1492 831 1496
rect 835 1492 836 1496
rect 830 1491 836 1492
rect 886 1496 892 1497
rect 886 1492 887 1496
rect 891 1492 892 1496
rect 1343 1495 1352 1496
rect 886 1491 892 1492
rect 1134 1492 1140 1493
rect 1134 1488 1135 1492
rect 1139 1488 1140 1492
rect 1343 1491 1344 1495
rect 1351 1491 1352 1495
rect 1343 1490 1352 1491
rect 1382 1495 1389 1496
rect 1382 1491 1383 1495
rect 1388 1491 1389 1495
rect 1382 1490 1389 1491
rect 1423 1495 1432 1496
rect 1423 1491 1424 1495
rect 1431 1491 1432 1495
rect 1423 1490 1432 1491
rect 1463 1495 1472 1496
rect 1463 1491 1464 1495
rect 1471 1491 1472 1495
rect 1463 1490 1472 1491
rect 1503 1495 1512 1496
rect 1503 1491 1504 1495
rect 1511 1491 1512 1495
rect 1516 1494 1518 1500
rect 1543 1495 1549 1496
rect 1543 1494 1544 1495
rect 1516 1492 1544 1494
rect 1503 1490 1512 1491
rect 1543 1491 1544 1492
rect 1548 1491 1549 1495
rect 1543 1490 1549 1491
rect 1583 1495 1589 1496
rect 1583 1491 1584 1495
rect 1588 1494 1589 1495
rect 1598 1495 1604 1496
rect 1598 1494 1599 1495
rect 1588 1492 1599 1494
rect 1588 1491 1589 1492
rect 1583 1490 1589 1491
rect 1598 1491 1599 1492
rect 1603 1491 1604 1495
rect 1598 1490 1604 1491
rect 1631 1495 1637 1496
rect 1631 1491 1632 1495
rect 1636 1494 1637 1495
rect 1654 1495 1660 1496
rect 1654 1494 1655 1495
rect 1636 1492 1655 1494
rect 1636 1491 1637 1492
rect 1631 1490 1637 1491
rect 1654 1491 1655 1492
rect 1659 1491 1660 1495
rect 1654 1490 1660 1491
rect 1687 1495 1693 1496
rect 1687 1491 1688 1495
rect 1692 1494 1693 1495
rect 1726 1495 1732 1496
rect 1726 1494 1727 1495
rect 1692 1492 1727 1494
rect 1692 1491 1693 1492
rect 1687 1490 1693 1491
rect 1726 1491 1727 1492
rect 1731 1491 1732 1495
rect 1726 1490 1732 1491
rect 1759 1495 1765 1496
rect 1759 1491 1760 1495
rect 1764 1494 1765 1495
rect 1799 1495 1805 1496
rect 1799 1494 1800 1495
rect 1764 1492 1800 1494
rect 1764 1491 1765 1492
rect 1759 1490 1765 1491
rect 1799 1491 1800 1492
rect 1804 1491 1805 1495
rect 1799 1490 1805 1491
rect 1839 1495 1845 1496
rect 1839 1491 1840 1495
rect 1844 1494 1845 1495
rect 1887 1495 1893 1496
rect 1887 1494 1888 1495
rect 1844 1492 1888 1494
rect 1844 1491 1845 1492
rect 1839 1490 1845 1491
rect 1887 1491 1888 1492
rect 1892 1491 1893 1495
rect 1887 1490 1893 1491
rect 1910 1495 1916 1496
rect 1910 1491 1911 1495
rect 1915 1494 1916 1495
rect 1927 1495 1933 1496
rect 1927 1494 1928 1495
rect 1915 1492 1928 1494
rect 1915 1491 1916 1492
rect 1910 1490 1916 1491
rect 1927 1491 1928 1492
rect 1932 1491 1933 1495
rect 1927 1490 1933 1491
rect 2015 1495 2021 1496
rect 2015 1491 2016 1495
rect 2020 1494 2021 1495
rect 2062 1495 2068 1496
rect 2062 1494 2063 1495
rect 2020 1492 2063 1494
rect 2020 1491 2021 1492
rect 2015 1490 2021 1491
rect 2062 1491 2063 1492
rect 2067 1491 2068 1495
rect 2062 1490 2068 1491
rect 2078 1495 2084 1496
rect 2078 1491 2079 1495
rect 2083 1494 2084 1495
rect 2095 1495 2101 1496
rect 2095 1494 2096 1495
rect 2083 1492 2096 1494
rect 2083 1491 2084 1492
rect 2078 1490 2084 1491
rect 2095 1491 2096 1492
rect 2100 1491 2101 1495
rect 2095 1490 2101 1491
rect 2118 1492 2124 1493
rect 1134 1487 1140 1488
rect 2118 1488 2119 1492
rect 2123 1488 2124 1492
rect 2118 1487 2124 1488
rect 1318 1484 1324 1485
rect 131 1483 137 1484
rect 131 1479 132 1483
rect 136 1482 137 1483
rect 150 1483 156 1484
rect 150 1482 151 1483
rect 136 1480 151 1482
rect 136 1479 137 1480
rect 131 1478 137 1479
rect 150 1479 151 1480
rect 155 1479 156 1483
rect 150 1478 156 1479
rect 162 1483 168 1484
rect 162 1479 163 1483
rect 167 1482 168 1483
rect 171 1483 177 1484
rect 171 1482 172 1483
rect 167 1480 172 1482
rect 167 1479 168 1480
rect 162 1478 168 1479
rect 171 1479 172 1480
rect 176 1479 177 1483
rect 171 1478 177 1479
rect 202 1483 208 1484
rect 202 1479 203 1483
rect 207 1482 208 1483
rect 211 1483 217 1484
rect 211 1482 212 1483
rect 207 1480 212 1482
rect 207 1479 208 1480
rect 202 1478 208 1479
rect 211 1479 212 1480
rect 216 1479 217 1483
rect 211 1478 217 1479
rect 242 1483 248 1484
rect 242 1479 243 1483
rect 247 1482 248 1483
rect 251 1483 257 1484
rect 251 1482 252 1483
rect 247 1480 252 1482
rect 247 1479 248 1480
rect 242 1478 248 1479
rect 251 1479 252 1480
rect 256 1479 257 1483
rect 251 1478 257 1479
rect 282 1483 288 1484
rect 282 1479 283 1483
rect 287 1482 288 1483
rect 291 1483 297 1484
rect 291 1482 292 1483
rect 287 1480 292 1482
rect 287 1479 288 1480
rect 282 1478 288 1479
rect 291 1479 292 1480
rect 296 1479 297 1483
rect 291 1478 297 1479
rect 322 1483 328 1484
rect 322 1479 323 1483
rect 327 1482 328 1483
rect 331 1483 337 1484
rect 331 1482 332 1483
rect 327 1480 332 1482
rect 327 1479 328 1480
rect 322 1478 328 1479
rect 331 1479 332 1480
rect 336 1479 337 1483
rect 331 1478 337 1479
rect 362 1483 368 1484
rect 362 1479 363 1483
rect 367 1482 368 1483
rect 371 1483 377 1484
rect 371 1482 372 1483
rect 367 1480 372 1482
rect 367 1479 368 1480
rect 362 1478 368 1479
rect 371 1479 372 1480
rect 376 1479 377 1483
rect 371 1478 377 1479
rect 402 1483 408 1484
rect 402 1479 403 1483
rect 407 1482 408 1483
rect 411 1483 417 1484
rect 411 1482 412 1483
rect 407 1480 412 1482
rect 407 1479 408 1480
rect 402 1478 408 1479
rect 411 1479 412 1480
rect 416 1479 417 1483
rect 411 1478 417 1479
rect 442 1483 448 1484
rect 442 1479 443 1483
rect 447 1482 448 1483
rect 451 1483 457 1484
rect 451 1482 452 1483
rect 447 1480 452 1482
rect 447 1479 448 1480
rect 442 1478 448 1479
rect 451 1479 452 1480
rect 456 1479 457 1483
rect 451 1478 457 1479
rect 482 1483 488 1484
rect 482 1479 483 1483
rect 487 1482 488 1483
rect 491 1483 497 1484
rect 491 1482 492 1483
rect 487 1480 492 1482
rect 487 1479 488 1480
rect 482 1478 488 1479
rect 491 1479 492 1480
rect 496 1479 497 1483
rect 491 1478 497 1479
rect 522 1483 528 1484
rect 522 1479 523 1483
rect 527 1482 528 1483
rect 531 1483 537 1484
rect 531 1482 532 1483
rect 527 1480 532 1482
rect 527 1479 528 1480
rect 522 1478 528 1479
rect 531 1479 532 1480
rect 536 1479 537 1483
rect 531 1478 537 1479
rect 546 1483 552 1484
rect 546 1479 547 1483
rect 551 1482 552 1483
rect 571 1483 577 1484
rect 571 1482 572 1483
rect 551 1480 572 1482
rect 551 1479 552 1480
rect 546 1478 552 1479
rect 571 1479 572 1480
rect 576 1479 577 1483
rect 571 1478 577 1479
rect 602 1483 608 1484
rect 602 1479 603 1483
rect 607 1482 608 1483
rect 611 1483 617 1484
rect 611 1482 612 1483
rect 607 1480 612 1482
rect 607 1479 608 1480
rect 602 1478 608 1479
rect 611 1479 612 1480
rect 616 1479 617 1483
rect 611 1478 617 1479
rect 642 1483 648 1484
rect 642 1479 643 1483
rect 647 1482 648 1483
rect 651 1483 657 1484
rect 651 1482 652 1483
rect 647 1480 652 1482
rect 647 1479 648 1480
rect 642 1478 648 1479
rect 651 1479 652 1480
rect 656 1479 657 1483
rect 651 1478 657 1479
rect 682 1483 688 1484
rect 682 1479 683 1483
rect 687 1482 688 1483
rect 691 1483 697 1484
rect 691 1482 692 1483
rect 687 1480 692 1482
rect 687 1479 688 1480
rect 682 1478 688 1479
rect 691 1479 692 1480
rect 696 1479 697 1483
rect 691 1478 697 1479
rect 722 1483 728 1484
rect 722 1479 723 1483
rect 727 1482 728 1483
rect 731 1483 737 1484
rect 731 1482 732 1483
rect 727 1480 732 1482
rect 727 1479 728 1480
rect 722 1478 728 1479
rect 731 1479 732 1480
rect 736 1479 737 1483
rect 731 1478 737 1479
rect 762 1483 768 1484
rect 762 1479 763 1483
rect 767 1482 768 1483
rect 771 1483 777 1484
rect 771 1482 772 1483
rect 767 1480 772 1482
rect 767 1479 768 1480
rect 762 1478 768 1479
rect 771 1479 772 1480
rect 776 1479 777 1483
rect 771 1478 777 1479
rect 827 1483 833 1484
rect 827 1479 828 1483
rect 832 1482 833 1483
rect 838 1483 844 1484
rect 838 1482 839 1483
rect 832 1480 839 1482
rect 832 1479 833 1480
rect 827 1478 833 1479
rect 838 1479 839 1480
rect 843 1479 844 1483
rect 838 1478 844 1479
rect 878 1483 889 1484
rect 878 1479 879 1483
rect 883 1479 884 1483
rect 888 1479 889 1483
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1358 1484 1364 1485
rect 1358 1480 1359 1484
rect 1363 1480 1364 1484
rect 1358 1479 1364 1480
rect 1398 1484 1404 1485
rect 1398 1480 1399 1484
rect 1403 1480 1404 1484
rect 1398 1479 1404 1480
rect 1438 1484 1444 1485
rect 1438 1480 1439 1484
rect 1443 1480 1444 1484
rect 1438 1479 1444 1480
rect 1478 1484 1484 1485
rect 1478 1480 1479 1484
rect 1483 1480 1484 1484
rect 1478 1479 1484 1480
rect 1518 1484 1524 1485
rect 1518 1480 1519 1484
rect 1523 1480 1524 1484
rect 1518 1479 1524 1480
rect 1558 1484 1564 1485
rect 1558 1480 1559 1484
rect 1563 1480 1564 1484
rect 1558 1479 1564 1480
rect 1606 1484 1612 1485
rect 1606 1480 1607 1484
rect 1611 1480 1612 1484
rect 1606 1479 1612 1480
rect 1662 1484 1668 1485
rect 1662 1480 1663 1484
rect 1667 1480 1668 1484
rect 1662 1479 1668 1480
rect 1734 1484 1740 1485
rect 1734 1480 1735 1484
rect 1739 1480 1740 1484
rect 1734 1479 1740 1480
rect 1814 1484 1820 1485
rect 1814 1480 1815 1484
rect 1819 1480 1820 1484
rect 1814 1479 1820 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 1990 1484 1996 1485
rect 1990 1480 1991 1484
rect 1995 1480 1996 1484
rect 1990 1479 1996 1480
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 878 1478 889 1479
rect 582 1471 588 1472
rect 582 1470 583 1471
rect 516 1468 583 1470
rect 516 1466 518 1468
rect 582 1467 583 1468
rect 587 1467 588 1471
rect 782 1471 788 1472
rect 782 1470 783 1471
rect 582 1466 588 1467
rect 644 1468 783 1470
rect 644 1466 646 1468
rect 782 1467 783 1468
rect 787 1467 788 1471
rect 782 1466 788 1467
rect 1315 1471 1321 1472
rect 1315 1467 1316 1471
rect 1320 1470 1321 1471
rect 1326 1471 1332 1472
rect 1326 1470 1327 1471
rect 1320 1468 1327 1470
rect 1320 1467 1321 1468
rect 1315 1466 1321 1467
rect 1326 1467 1327 1468
rect 1331 1467 1332 1471
rect 1326 1466 1332 1467
rect 1346 1471 1352 1472
rect 1346 1467 1347 1471
rect 1351 1470 1352 1471
rect 1355 1471 1361 1472
rect 1355 1470 1356 1471
rect 1351 1468 1356 1470
rect 1351 1467 1352 1468
rect 1346 1466 1352 1467
rect 1355 1467 1356 1468
rect 1360 1467 1361 1471
rect 1355 1466 1361 1467
rect 1382 1471 1388 1472
rect 1382 1467 1383 1471
rect 1387 1470 1388 1471
rect 1395 1471 1401 1472
rect 1395 1470 1396 1471
rect 1387 1468 1396 1470
rect 1387 1467 1388 1468
rect 1382 1466 1388 1467
rect 1395 1467 1396 1468
rect 1400 1467 1401 1471
rect 1395 1466 1401 1467
rect 1426 1471 1432 1472
rect 1426 1467 1427 1471
rect 1431 1470 1432 1471
rect 1435 1471 1441 1472
rect 1435 1470 1436 1471
rect 1431 1468 1436 1470
rect 1431 1467 1432 1468
rect 1426 1466 1432 1467
rect 1435 1467 1436 1468
rect 1440 1467 1441 1471
rect 1435 1466 1441 1467
rect 1466 1471 1472 1472
rect 1466 1467 1467 1471
rect 1471 1470 1472 1471
rect 1475 1471 1481 1472
rect 1475 1470 1476 1471
rect 1471 1468 1476 1470
rect 1471 1467 1472 1468
rect 1466 1466 1472 1467
rect 1475 1467 1476 1468
rect 1480 1467 1481 1471
rect 1475 1466 1481 1467
rect 1506 1471 1512 1472
rect 1506 1467 1507 1471
rect 1511 1470 1512 1471
rect 1515 1471 1521 1472
rect 1515 1470 1516 1471
rect 1511 1468 1516 1470
rect 1511 1467 1512 1468
rect 1506 1466 1512 1467
rect 1515 1467 1516 1468
rect 1520 1467 1521 1471
rect 1515 1466 1521 1467
rect 1546 1471 1552 1472
rect 1546 1467 1547 1471
rect 1551 1470 1552 1471
rect 1555 1471 1561 1472
rect 1555 1470 1556 1471
rect 1551 1468 1556 1470
rect 1551 1467 1552 1468
rect 1546 1466 1552 1467
rect 1555 1467 1556 1468
rect 1560 1467 1561 1471
rect 1555 1466 1561 1467
rect 1598 1471 1609 1472
rect 1598 1467 1599 1471
rect 1603 1467 1604 1471
rect 1608 1467 1609 1471
rect 1598 1466 1609 1467
rect 1654 1471 1665 1472
rect 1654 1467 1655 1471
rect 1659 1467 1660 1471
rect 1664 1467 1665 1471
rect 1654 1466 1665 1467
rect 1726 1471 1737 1472
rect 1726 1467 1727 1471
rect 1731 1467 1732 1471
rect 1736 1467 1737 1471
rect 1726 1466 1737 1467
rect 1799 1471 1805 1472
rect 1799 1467 1800 1471
rect 1804 1470 1805 1471
rect 1811 1471 1817 1472
rect 1811 1470 1812 1471
rect 1804 1468 1812 1470
rect 1804 1467 1805 1468
rect 1799 1466 1805 1467
rect 1811 1467 1812 1468
rect 1816 1467 1817 1471
rect 1811 1466 1817 1467
rect 1887 1471 1893 1472
rect 1887 1467 1888 1471
rect 1892 1470 1893 1471
rect 1899 1471 1905 1472
rect 1899 1470 1900 1471
rect 1892 1468 1900 1470
rect 1892 1467 1893 1468
rect 1887 1466 1893 1467
rect 1899 1467 1900 1468
rect 1904 1467 1905 1471
rect 1899 1466 1905 1467
rect 1987 1471 1993 1472
rect 1987 1467 1988 1471
rect 1992 1470 1993 1471
rect 2038 1471 2044 1472
rect 2038 1470 2039 1471
rect 1992 1468 2039 1470
rect 1992 1467 1993 1468
rect 1987 1466 1993 1467
rect 2038 1467 2039 1468
rect 2043 1467 2044 1471
rect 2038 1466 2044 1467
rect 2062 1471 2073 1472
rect 2062 1467 2063 1471
rect 2067 1467 2068 1471
rect 2072 1467 2073 1471
rect 2062 1466 2073 1467
rect 515 1465 521 1466
rect 515 1461 516 1465
rect 520 1461 521 1465
rect 643 1465 649 1466
rect 515 1460 521 1461
rect 555 1463 561 1464
rect 555 1459 556 1463
rect 560 1462 561 1463
rect 595 1463 601 1464
rect 560 1460 590 1462
rect 560 1459 561 1460
rect 555 1458 561 1459
rect 518 1452 524 1453
rect 518 1448 519 1452
rect 523 1448 524 1452
rect 518 1447 524 1448
rect 558 1452 564 1453
rect 558 1448 559 1452
rect 563 1448 564 1452
rect 558 1447 564 1448
rect 588 1446 590 1460
rect 595 1459 596 1463
rect 600 1462 601 1463
rect 600 1460 638 1462
rect 643 1461 644 1465
rect 648 1461 649 1465
rect 643 1460 649 1461
rect 674 1463 680 1464
rect 600 1459 601 1460
rect 595 1458 601 1459
rect 636 1458 638 1460
rect 654 1459 660 1460
rect 654 1458 655 1459
rect 636 1456 655 1458
rect 654 1455 655 1456
rect 659 1455 660 1459
rect 674 1459 675 1463
rect 679 1462 680 1463
rect 691 1463 697 1464
rect 691 1462 692 1463
rect 679 1460 692 1462
rect 679 1459 680 1460
rect 674 1458 680 1459
rect 691 1459 692 1460
rect 696 1459 697 1463
rect 691 1458 697 1459
rect 735 1463 741 1464
rect 735 1459 736 1463
rect 740 1462 741 1463
rect 747 1463 753 1464
rect 747 1462 748 1463
rect 740 1460 748 1462
rect 740 1459 741 1460
rect 735 1458 741 1459
rect 747 1459 748 1460
rect 752 1459 753 1463
rect 747 1458 753 1459
rect 786 1463 792 1464
rect 786 1459 787 1463
rect 791 1462 792 1463
rect 803 1463 809 1464
rect 803 1462 804 1463
rect 791 1460 804 1462
rect 791 1459 792 1460
rect 786 1458 792 1459
rect 803 1459 804 1460
rect 808 1459 809 1463
rect 803 1458 809 1459
rect 867 1463 873 1464
rect 867 1459 868 1463
rect 872 1462 873 1463
rect 918 1463 924 1464
rect 918 1462 919 1463
rect 872 1460 919 1462
rect 872 1459 873 1460
rect 867 1458 873 1459
rect 918 1459 919 1460
rect 923 1459 924 1463
rect 918 1458 924 1459
rect 926 1463 937 1464
rect 926 1459 927 1463
rect 931 1459 932 1463
rect 936 1459 937 1463
rect 926 1458 937 1459
rect 1227 1459 1233 1460
rect 654 1454 660 1455
rect 1227 1455 1228 1459
rect 1232 1458 1233 1459
rect 1250 1459 1256 1460
rect 1250 1458 1251 1459
rect 1232 1456 1251 1458
rect 1232 1455 1233 1456
rect 1227 1454 1233 1455
rect 1250 1455 1251 1456
rect 1255 1455 1256 1459
rect 1250 1454 1256 1455
rect 1258 1459 1264 1460
rect 1258 1455 1259 1459
rect 1263 1458 1264 1459
rect 1275 1459 1281 1460
rect 1275 1458 1276 1459
rect 1263 1456 1276 1458
rect 1263 1455 1264 1456
rect 1258 1454 1264 1455
rect 1275 1455 1276 1456
rect 1280 1455 1281 1459
rect 1275 1454 1281 1455
rect 1306 1459 1312 1460
rect 1306 1455 1307 1459
rect 1311 1458 1312 1459
rect 1331 1459 1337 1460
rect 1331 1458 1332 1459
rect 1311 1456 1332 1458
rect 1311 1455 1312 1456
rect 1306 1454 1312 1455
rect 1331 1455 1332 1456
rect 1336 1455 1337 1459
rect 1387 1459 1393 1460
rect 1331 1454 1337 1455
rect 1362 1455 1368 1456
rect 598 1452 604 1453
rect 598 1448 599 1452
rect 603 1448 604 1452
rect 598 1447 604 1448
rect 646 1452 652 1453
rect 646 1448 647 1452
rect 651 1448 652 1452
rect 646 1447 652 1448
rect 694 1452 700 1453
rect 694 1448 695 1452
rect 699 1448 700 1452
rect 694 1447 700 1448
rect 750 1452 756 1453
rect 750 1448 751 1452
rect 755 1448 756 1452
rect 750 1447 756 1448
rect 806 1452 812 1453
rect 806 1448 807 1452
rect 811 1448 812 1452
rect 806 1447 812 1448
rect 870 1452 876 1453
rect 870 1448 871 1452
rect 875 1448 876 1452
rect 870 1447 876 1448
rect 934 1452 940 1453
rect 934 1448 935 1452
rect 939 1448 940 1452
rect 1362 1451 1363 1455
rect 1367 1454 1368 1455
rect 1387 1455 1388 1459
rect 1392 1455 1393 1459
rect 1387 1454 1393 1455
rect 1418 1459 1424 1460
rect 1418 1455 1419 1459
rect 1423 1458 1424 1459
rect 1451 1459 1457 1460
rect 1451 1458 1452 1459
rect 1423 1456 1452 1458
rect 1423 1455 1424 1456
rect 1418 1454 1424 1455
rect 1451 1455 1452 1456
rect 1456 1455 1457 1459
rect 1451 1454 1457 1455
rect 1486 1459 1492 1460
rect 1486 1455 1487 1459
rect 1491 1458 1492 1459
rect 1515 1459 1521 1460
rect 1515 1458 1516 1459
rect 1491 1456 1516 1458
rect 1491 1455 1492 1456
rect 1486 1454 1492 1455
rect 1515 1455 1516 1456
rect 1520 1455 1521 1459
rect 1515 1454 1521 1455
rect 1579 1459 1585 1460
rect 1579 1455 1580 1459
rect 1584 1458 1585 1459
rect 1590 1459 1596 1460
rect 1590 1458 1591 1459
rect 1584 1456 1591 1458
rect 1584 1455 1585 1456
rect 1579 1454 1585 1455
rect 1590 1455 1591 1456
rect 1595 1455 1596 1459
rect 1590 1454 1596 1455
rect 1614 1459 1620 1460
rect 1614 1455 1615 1459
rect 1619 1458 1620 1459
rect 1643 1459 1649 1460
rect 1643 1458 1644 1459
rect 1619 1456 1644 1458
rect 1619 1455 1620 1456
rect 1614 1454 1620 1455
rect 1643 1455 1644 1456
rect 1648 1455 1649 1459
rect 1643 1454 1649 1455
rect 1674 1459 1680 1460
rect 1674 1455 1675 1459
rect 1679 1458 1680 1459
rect 1715 1459 1721 1460
rect 1715 1458 1716 1459
rect 1679 1456 1716 1458
rect 1679 1455 1680 1456
rect 1674 1454 1680 1455
rect 1715 1455 1716 1456
rect 1720 1455 1721 1459
rect 1715 1454 1721 1455
rect 1746 1459 1752 1460
rect 1746 1455 1747 1459
rect 1751 1458 1752 1459
rect 1803 1459 1809 1460
rect 1803 1458 1804 1459
rect 1751 1456 1804 1458
rect 1751 1455 1752 1456
rect 1746 1454 1752 1455
rect 1803 1455 1804 1456
rect 1808 1455 1809 1459
rect 1803 1454 1809 1455
rect 1834 1459 1840 1460
rect 1834 1455 1835 1459
rect 1839 1458 1840 1459
rect 1891 1459 1897 1460
rect 1891 1458 1892 1459
rect 1839 1456 1892 1458
rect 1839 1455 1840 1456
rect 1834 1454 1840 1455
rect 1891 1455 1892 1456
rect 1896 1455 1897 1459
rect 1891 1454 1897 1455
rect 1922 1459 1928 1460
rect 1922 1455 1923 1459
rect 1927 1458 1928 1459
rect 1987 1459 1993 1460
rect 1987 1458 1988 1459
rect 1927 1456 1988 1458
rect 1927 1455 1928 1456
rect 1922 1454 1928 1455
rect 1987 1455 1988 1456
rect 1992 1455 1993 1459
rect 1987 1454 1993 1455
rect 2067 1459 2073 1460
rect 2067 1455 2068 1459
rect 2072 1458 2073 1459
rect 2078 1459 2084 1460
rect 2078 1458 2079 1459
rect 2072 1456 2079 1458
rect 2072 1455 2073 1456
rect 2067 1454 2073 1455
rect 2078 1455 2079 1456
rect 2083 1455 2084 1459
rect 2078 1454 2084 1455
rect 1367 1452 1391 1454
rect 1367 1451 1368 1452
rect 1362 1450 1368 1451
rect 934 1447 940 1448
rect 1230 1448 1236 1449
rect 110 1444 116 1445
rect 588 1444 594 1446
rect 1094 1444 1100 1445
rect 110 1440 111 1444
rect 115 1440 116 1444
rect 110 1439 116 1440
rect 543 1439 552 1440
rect 543 1435 544 1439
rect 551 1435 552 1439
rect 543 1434 552 1435
rect 582 1439 589 1440
rect 582 1435 583 1439
rect 588 1435 589 1439
rect 592 1438 594 1444
rect 786 1443 792 1444
rect 786 1442 787 1443
rect 775 1441 787 1442
rect 623 1439 629 1440
rect 623 1438 624 1439
rect 592 1436 624 1438
rect 582 1434 589 1435
rect 623 1435 624 1436
rect 628 1435 629 1439
rect 623 1434 629 1435
rect 671 1439 680 1440
rect 671 1435 672 1439
rect 679 1435 680 1439
rect 671 1434 680 1435
rect 719 1439 725 1440
rect 719 1435 720 1439
rect 724 1438 725 1439
rect 735 1439 741 1440
rect 735 1438 736 1439
rect 724 1436 736 1438
rect 724 1435 725 1436
rect 719 1434 725 1435
rect 735 1435 736 1436
rect 740 1435 741 1439
rect 775 1437 776 1441
rect 780 1440 787 1441
rect 780 1437 781 1440
rect 786 1439 787 1440
rect 791 1439 792 1443
rect 1094 1440 1095 1444
rect 1099 1440 1100 1444
rect 1230 1444 1231 1448
rect 1235 1444 1236 1448
rect 1230 1443 1236 1444
rect 1278 1448 1284 1449
rect 1278 1444 1279 1448
rect 1283 1444 1284 1448
rect 1278 1443 1284 1444
rect 1334 1448 1340 1449
rect 1334 1444 1335 1448
rect 1339 1444 1340 1448
rect 1334 1443 1340 1444
rect 1390 1448 1396 1449
rect 1390 1444 1391 1448
rect 1395 1444 1396 1448
rect 1390 1443 1396 1444
rect 1454 1448 1460 1449
rect 1454 1444 1455 1448
rect 1459 1444 1460 1448
rect 1454 1443 1460 1444
rect 1518 1448 1524 1449
rect 1518 1444 1519 1448
rect 1523 1444 1524 1448
rect 1518 1443 1524 1444
rect 1582 1448 1588 1449
rect 1582 1444 1583 1448
rect 1587 1444 1588 1448
rect 1582 1443 1588 1444
rect 1646 1448 1652 1449
rect 1646 1444 1647 1448
rect 1651 1444 1652 1448
rect 1646 1443 1652 1444
rect 1718 1448 1724 1449
rect 1718 1444 1719 1448
rect 1723 1444 1724 1448
rect 1718 1443 1724 1444
rect 1806 1448 1812 1449
rect 1806 1444 1807 1448
rect 1811 1444 1812 1448
rect 1806 1443 1812 1444
rect 1894 1448 1900 1449
rect 1894 1444 1895 1448
rect 1899 1444 1900 1448
rect 1894 1443 1900 1444
rect 1990 1448 1996 1449
rect 1990 1444 1991 1448
rect 1995 1444 1996 1448
rect 1990 1443 1996 1444
rect 2070 1448 2076 1449
rect 2070 1444 2071 1448
rect 2075 1444 2076 1448
rect 2070 1443 2076 1444
rect 786 1438 792 1439
rect 830 1439 837 1440
rect 775 1436 781 1437
rect 735 1434 741 1435
rect 830 1435 831 1439
rect 836 1435 837 1439
rect 830 1434 837 1435
rect 886 1439 892 1440
rect 886 1435 887 1439
rect 891 1438 892 1439
rect 895 1439 901 1440
rect 895 1438 896 1439
rect 891 1436 896 1438
rect 891 1435 892 1436
rect 886 1434 892 1435
rect 895 1435 896 1436
rect 900 1435 901 1439
rect 895 1434 901 1435
rect 918 1439 924 1440
rect 918 1435 919 1439
rect 923 1438 924 1439
rect 959 1439 965 1440
rect 1094 1439 1100 1440
rect 1134 1440 1140 1441
rect 959 1438 960 1439
rect 923 1436 960 1438
rect 923 1435 924 1436
rect 918 1434 924 1435
rect 959 1435 960 1436
rect 964 1435 965 1439
rect 1134 1436 1135 1440
rect 1139 1436 1140 1440
rect 2118 1440 2124 1441
rect 2118 1436 2119 1440
rect 2123 1436 2124 1440
rect 1134 1435 1140 1436
rect 1255 1435 1264 1436
rect 959 1434 965 1435
rect 1255 1431 1256 1435
rect 1263 1431 1264 1435
rect 1255 1430 1264 1431
rect 1303 1435 1312 1436
rect 1303 1431 1304 1435
rect 1311 1431 1312 1435
rect 1303 1430 1312 1431
rect 1359 1435 1368 1436
rect 1359 1431 1360 1435
rect 1367 1431 1368 1435
rect 1359 1430 1368 1431
rect 1415 1435 1424 1436
rect 1415 1431 1416 1435
rect 1423 1431 1424 1435
rect 1415 1430 1424 1431
rect 1479 1435 1488 1436
rect 1479 1431 1480 1435
rect 1487 1431 1488 1435
rect 1479 1430 1488 1431
rect 1542 1435 1549 1436
rect 1542 1431 1543 1435
rect 1548 1431 1549 1435
rect 1542 1430 1549 1431
rect 1607 1435 1616 1436
rect 1607 1431 1608 1435
rect 1615 1431 1616 1435
rect 1607 1430 1616 1431
rect 1671 1435 1680 1436
rect 1671 1431 1672 1435
rect 1679 1431 1680 1435
rect 1671 1430 1680 1431
rect 1743 1435 1752 1436
rect 1743 1431 1744 1435
rect 1751 1431 1752 1435
rect 1743 1430 1752 1431
rect 1831 1435 1840 1436
rect 1831 1431 1832 1435
rect 1839 1431 1840 1435
rect 1831 1430 1840 1431
rect 1919 1435 1928 1436
rect 1919 1431 1920 1435
rect 1927 1431 1928 1435
rect 1919 1430 1928 1431
rect 1930 1435 1936 1436
rect 1930 1431 1931 1435
rect 1935 1434 1936 1435
rect 2015 1435 2021 1436
rect 2015 1434 2016 1435
rect 1935 1432 2016 1434
rect 1935 1431 1936 1432
rect 1930 1430 1936 1431
rect 2015 1431 2016 1432
rect 2020 1431 2021 1435
rect 2015 1430 2021 1431
rect 2090 1435 2101 1436
rect 2118 1435 2124 1436
rect 2090 1431 2091 1435
rect 2095 1431 2096 1435
rect 2100 1431 2101 1435
rect 2090 1430 2101 1431
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 1094 1427 1100 1428
rect 110 1422 116 1423
rect 518 1424 524 1425
rect 518 1420 519 1424
rect 523 1420 524 1424
rect 518 1419 524 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 646 1424 652 1425
rect 646 1420 647 1424
rect 651 1420 652 1424
rect 646 1419 652 1420
rect 694 1424 700 1425
rect 694 1420 695 1424
rect 699 1420 700 1424
rect 694 1419 700 1420
rect 750 1424 756 1425
rect 750 1420 751 1424
rect 755 1420 756 1424
rect 750 1419 756 1420
rect 806 1424 812 1425
rect 806 1420 807 1424
rect 811 1420 812 1424
rect 806 1419 812 1420
rect 870 1424 876 1425
rect 870 1420 871 1424
rect 875 1420 876 1424
rect 870 1419 876 1420
rect 934 1424 940 1425
rect 934 1420 935 1424
rect 939 1420 940 1424
rect 1094 1423 1095 1427
rect 1099 1423 1100 1427
rect 1094 1422 1100 1423
rect 1134 1423 1140 1424
rect 934 1419 940 1420
rect 1134 1419 1135 1423
rect 1139 1419 1140 1423
rect 2118 1423 2124 1424
rect 1134 1418 1140 1419
rect 1230 1420 1236 1421
rect 1230 1416 1231 1420
rect 1235 1416 1236 1420
rect 1230 1415 1236 1416
rect 1278 1420 1284 1421
rect 1278 1416 1279 1420
rect 1283 1416 1284 1420
rect 1278 1415 1284 1416
rect 1334 1420 1340 1421
rect 1334 1416 1335 1420
rect 1339 1416 1340 1420
rect 1334 1415 1340 1416
rect 1390 1420 1396 1421
rect 1390 1416 1391 1420
rect 1395 1416 1396 1420
rect 1390 1415 1396 1416
rect 1454 1420 1460 1421
rect 1454 1416 1455 1420
rect 1459 1416 1460 1420
rect 1454 1415 1460 1416
rect 1518 1420 1524 1421
rect 1518 1416 1519 1420
rect 1523 1416 1524 1420
rect 1518 1415 1524 1416
rect 1582 1420 1588 1421
rect 1582 1416 1583 1420
rect 1587 1416 1588 1420
rect 1582 1415 1588 1416
rect 1646 1420 1652 1421
rect 1646 1416 1647 1420
rect 1651 1416 1652 1420
rect 1646 1415 1652 1416
rect 1718 1420 1724 1421
rect 1718 1416 1719 1420
rect 1723 1416 1724 1420
rect 1718 1415 1724 1416
rect 1806 1420 1812 1421
rect 1806 1416 1807 1420
rect 1811 1416 1812 1420
rect 1806 1415 1812 1416
rect 1894 1420 1900 1421
rect 1894 1416 1895 1420
rect 1899 1416 1900 1420
rect 1894 1415 1900 1416
rect 1990 1420 1996 1421
rect 1990 1416 1991 1420
rect 1995 1416 1996 1420
rect 1990 1415 1996 1416
rect 2070 1420 2076 1421
rect 2070 1416 2071 1420
rect 2075 1416 2076 1420
rect 2118 1419 2119 1423
rect 2123 1419 2124 1423
rect 2118 1418 2124 1419
rect 2070 1415 2076 1416
rect 430 1408 436 1409
rect 110 1405 116 1406
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 430 1404 431 1408
rect 435 1404 436 1408
rect 430 1403 436 1404
rect 470 1408 476 1409
rect 470 1404 471 1408
rect 475 1404 476 1408
rect 470 1403 476 1404
rect 518 1408 524 1409
rect 518 1404 519 1408
rect 523 1404 524 1408
rect 518 1403 524 1404
rect 574 1408 580 1409
rect 574 1404 575 1408
rect 579 1404 580 1408
rect 574 1403 580 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 694 1408 700 1409
rect 694 1404 695 1408
rect 699 1404 700 1408
rect 694 1403 700 1404
rect 758 1408 764 1409
rect 758 1404 759 1408
rect 763 1404 764 1408
rect 758 1403 764 1404
rect 822 1408 828 1409
rect 822 1404 823 1408
rect 827 1404 828 1408
rect 822 1403 828 1404
rect 894 1408 900 1409
rect 894 1404 895 1408
rect 899 1404 900 1408
rect 894 1403 900 1404
rect 966 1408 972 1409
rect 966 1404 967 1408
rect 971 1404 972 1408
rect 966 1403 972 1404
rect 1094 1405 1100 1406
rect 110 1400 116 1401
rect 1094 1401 1095 1405
rect 1099 1401 1100 1405
rect 1158 1404 1164 1405
rect 1094 1400 1100 1401
rect 1134 1401 1140 1402
rect 1134 1397 1135 1401
rect 1139 1397 1140 1401
rect 1158 1400 1159 1404
rect 1163 1400 1164 1404
rect 1158 1399 1164 1400
rect 1198 1404 1204 1405
rect 1198 1400 1199 1404
rect 1203 1400 1204 1404
rect 1198 1399 1204 1400
rect 1262 1404 1268 1405
rect 1262 1400 1263 1404
rect 1267 1400 1268 1404
rect 1262 1399 1268 1400
rect 1350 1404 1356 1405
rect 1350 1400 1351 1404
rect 1355 1400 1356 1404
rect 1350 1399 1356 1400
rect 1446 1404 1452 1405
rect 1446 1400 1447 1404
rect 1451 1400 1452 1404
rect 1446 1399 1452 1400
rect 1542 1404 1548 1405
rect 1542 1400 1543 1404
rect 1547 1400 1548 1404
rect 1542 1399 1548 1400
rect 1630 1404 1636 1405
rect 1630 1400 1631 1404
rect 1635 1400 1636 1404
rect 1630 1399 1636 1400
rect 1718 1404 1724 1405
rect 1718 1400 1719 1404
rect 1723 1400 1724 1404
rect 1718 1399 1724 1400
rect 1798 1404 1804 1405
rect 1798 1400 1799 1404
rect 1803 1400 1804 1404
rect 1798 1399 1804 1400
rect 1870 1404 1876 1405
rect 1870 1400 1871 1404
rect 1875 1400 1876 1404
rect 1870 1399 1876 1400
rect 1942 1404 1948 1405
rect 1942 1400 1943 1404
rect 1947 1400 1948 1404
rect 1942 1399 1948 1400
rect 2014 1404 2020 1405
rect 2014 1400 2015 1404
rect 2019 1400 2020 1404
rect 2014 1399 2020 1400
rect 2070 1404 2076 1405
rect 2070 1400 2071 1404
rect 2075 1400 2076 1404
rect 2070 1399 2076 1400
rect 2118 1401 2124 1402
rect 1134 1396 1140 1397
rect 2118 1397 2119 1401
rect 2123 1397 2124 1401
rect 2118 1396 2124 1397
rect 1250 1395 1256 1396
rect 455 1391 464 1392
rect 110 1388 116 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 455 1387 456 1391
rect 463 1387 464 1391
rect 455 1386 464 1387
rect 495 1391 501 1392
rect 495 1387 496 1391
rect 500 1390 501 1391
rect 510 1391 516 1392
rect 510 1390 511 1391
rect 500 1388 511 1390
rect 500 1387 501 1388
rect 495 1386 501 1387
rect 510 1387 511 1388
rect 515 1387 516 1391
rect 510 1386 516 1387
rect 543 1391 549 1392
rect 543 1387 544 1391
rect 548 1390 549 1391
rect 566 1391 572 1392
rect 566 1390 567 1391
rect 548 1388 567 1390
rect 548 1387 549 1388
rect 543 1386 549 1387
rect 566 1387 567 1388
rect 571 1387 572 1391
rect 566 1386 572 1387
rect 599 1391 605 1392
rect 599 1387 600 1391
rect 604 1390 605 1391
rect 622 1391 628 1392
rect 622 1390 623 1391
rect 604 1388 623 1390
rect 604 1387 605 1388
rect 599 1386 605 1387
rect 622 1387 623 1388
rect 627 1387 628 1391
rect 622 1386 628 1387
rect 654 1391 661 1392
rect 654 1387 655 1391
rect 660 1387 661 1391
rect 654 1386 661 1387
rect 702 1391 708 1392
rect 702 1387 703 1391
rect 707 1390 708 1391
rect 719 1391 725 1392
rect 719 1390 720 1391
rect 707 1388 720 1390
rect 707 1387 708 1388
rect 702 1386 708 1387
rect 719 1387 720 1388
rect 724 1387 725 1391
rect 719 1386 725 1387
rect 727 1391 733 1392
rect 727 1387 728 1391
rect 732 1390 733 1391
rect 783 1391 789 1392
rect 783 1390 784 1391
rect 732 1388 784 1390
rect 732 1387 733 1388
rect 727 1386 733 1387
rect 783 1387 784 1388
rect 788 1387 789 1391
rect 783 1386 789 1387
rect 791 1391 797 1392
rect 791 1387 792 1391
rect 796 1390 797 1391
rect 847 1391 853 1392
rect 847 1390 848 1391
rect 796 1388 848 1390
rect 796 1387 797 1388
rect 791 1386 797 1387
rect 847 1387 848 1388
rect 852 1387 853 1391
rect 847 1386 853 1387
rect 919 1391 925 1392
rect 919 1387 920 1391
rect 924 1390 925 1391
rect 958 1391 964 1392
rect 958 1390 959 1391
rect 924 1388 959 1390
rect 924 1387 925 1388
rect 919 1386 925 1387
rect 958 1387 959 1388
rect 963 1387 964 1391
rect 958 1386 964 1387
rect 990 1391 997 1392
rect 990 1387 991 1391
rect 996 1387 997 1391
rect 1250 1391 1251 1395
rect 1255 1394 1256 1395
rect 1255 1392 1546 1394
rect 1255 1391 1256 1392
rect 1250 1390 1256 1391
rect 990 1386 997 1387
rect 1094 1388 1100 1389
rect 110 1383 116 1384
rect 1094 1384 1095 1388
rect 1099 1384 1100 1388
rect 1183 1387 1192 1388
rect 1094 1383 1100 1384
rect 1134 1384 1140 1385
rect 430 1380 436 1381
rect 430 1376 431 1380
rect 435 1376 436 1380
rect 430 1375 436 1376
rect 470 1380 476 1381
rect 470 1376 471 1380
rect 475 1376 476 1380
rect 470 1375 476 1376
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 574 1380 580 1381
rect 574 1376 575 1380
rect 579 1376 580 1380
rect 574 1375 580 1376
rect 630 1380 636 1381
rect 630 1376 631 1380
rect 635 1376 636 1380
rect 630 1375 636 1376
rect 694 1380 700 1381
rect 694 1376 695 1380
rect 699 1376 700 1380
rect 694 1375 700 1376
rect 758 1380 764 1381
rect 758 1376 759 1380
rect 763 1376 764 1380
rect 758 1375 764 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 894 1380 900 1381
rect 894 1376 895 1380
rect 899 1376 900 1380
rect 894 1375 900 1376
rect 966 1380 972 1381
rect 966 1376 967 1380
rect 971 1376 972 1380
rect 1134 1380 1135 1384
rect 1139 1380 1140 1384
rect 1183 1383 1184 1387
rect 1191 1383 1192 1387
rect 1183 1382 1192 1383
rect 1223 1387 1229 1388
rect 1223 1383 1224 1387
rect 1228 1386 1229 1387
rect 1254 1387 1260 1388
rect 1254 1386 1255 1387
rect 1228 1384 1255 1386
rect 1228 1383 1229 1384
rect 1223 1382 1229 1383
rect 1254 1383 1255 1384
rect 1259 1383 1260 1387
rect 1254 1382 1260 1383
rect 1287 1387 1293 1388
rect 1287 1383 1288 1387
rect 1292 1386 1293 1387
rect 1342 1387 1348 1388
rect 1342 1386 1343 1387
rect 1292 1384 1343 1386
rect 1292 1383 1293 1384
rect 1287 1382 1293 1383
rect 1342 1383 1343 1384
rect 1347 1383 1348 1387
rect 1342 1382 1348 1383
rect 1375 1387 1381 1388
rect 1375 1383 1376 1387
rect 1380 1386 1381 1387
rect 1438 1387 1444 1388
rect 1438 1386 1439 1387
rect 1380 1384 1439 1386
rect 1380 1383 1381 1384
rect 1375 1382 1381 1383
rect 1438 1383 1439 1384
rect 1443 1383 1444 1387
rect 1438 1382 1444 1383
rect 1471 1387 1477 1388
rect 1471 1383 1472 1387
rect 1476 1386 1477 1387
rect 1534 1387 1540 1388
rect 1534 1386 1535 1387
rect 1476 1384 1535 1386
rect 1476 1383 1477 1384
rect 1471 1382 1477 1383
rect 1534 1383 1535 1384
rect 1539 1383 1540 1387
rect 1544 1386 1546 1392
rect 1567 1387 1573 1388
rect 1567 1386 1568 1387
rect 1544 1384 1568 1386
rect 1534 1382 1540 1383
rect 1567 1383 1568 1384
rect 1572 1383 1573 1387
rect 1567 1382 1573 1383
rect 1655 1387 1661 1388
rect 1655 1383 1656 1387
rect 1660 1386 1661 1387
rect 1710 1387 1716 1388
rect 1710 1386 1711 1387
rect 1660 1384 1711 1386
rect 1660 1383 1661 1384
rect 1655 1382 1661 1383
rect 1710 1383 1711 1384
rect 1715 1383 1716 1387
rect 1710 1382 1716 1383
rect 1743 1387 1749 1388
rect 1743 1383 1744 1387
rect 1748 1386 1749 1387
rect 1790 1387 1796 1388
rect 1790 1386 1791 1387
rect 1748 1384 1791 1386
rect 1748 1383 1749 1384
rect 1743 1382 1749 1383
rect 1790 1383 1791 1384
rect 1795 1383 1796 1387
rect 1790 1382 1796 1383
rect 1823 1387 1829 1388
rect 1823 1383 1824 1387
rect 1828 1386 1829 1387
rect 1862 1387 1868 1388
rect 1862 1386 1863 1387
rect 1828 1384 1863 1386
rect 1828 1383 1829 1384
rect 1823 1382 1829 1383
rect 1862 1383 1863 1384
rect 1867 1383 1868 1387
rect 1862 1382 1868 1383
rect 1886 1387 1892 1388
rect 1886 1383 1887 1387
rect 1891 1386 1892 1387
rect 1895 1387 1901 1388
rect 1895 1386 1896 1387
rect 1891 1384 1896 1386
rect 1891 1383 1892 1384
rect 1886 1382 1892 1383
rect 1895 1383 1896 1384
rect 1900 1383 1901 1387
rect 1895 1382 1901 1383
rect 1967 1387 1973 1388
rect 1967 1383 1968 1387
rect 1972 1386 1973 1387
rect 2006 1387 2012 1388
rect 2006 1386 2007 1387
rect 1972 1384 2007 1386
rect 1972 1383 1973 1384
rect 1967 1382 1973 1383
rect 2006 1383 2007 1384
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2038 1387 2045 1388
rect 2038 1383 2039 1387
rect 2044 1383 2045 1387
rect 2038 1382 2045 1383
rect 2082 1387 2088 1388
rect 2082 1383 2083 1387
rect 2087 1386 2088 1387
rect 2095 1387 2101 1388
rect 2095 1386 2096 1387
rect 2087 1384 2096 1386
rect 2087 1383 2088 1384
rect 2082 1382 2088 1383
rect 2095 1383 2096 1384
rect 2100 1383 2101 1387
rect 2095 1382 2101 1383
rect 2118 1384 2124 1385
rect 1134 1379 1140 1380
rect 2118 1380 2119 1384
rect 2123 1380 2124 1384
rect 2118 1379 2124 1380
rect 966 1375 972 1376
rect 1158 1376 1164 1377
rect 1158 1372 1159 1376
rect 1163 1372 1164 1376
rect 1158 1371 1164 1372
rect 1198 1376 1204 1377
rect 1198 1372 1199 1376
rect 1203 1372 1204 1376
rect 1198 1371 1204 1372
rect 1262 1376 1268 1377
rect 1262 1372 1263 1376
rect 1267 1372 1268 1376
rect 1262 1371 1268 1372
rect 1350 1376 1356 1377
rect 1350 1372 1351 1376
rect 1355 1372 1356 1376
rect 1350 1371 1356 1372
rect 1446 1376 1452 1377
rect 1446 1372 1447 1376
rect 1451 1372 1452 1376
rect 1446 1371 1452 1372
rect 1542 1376 1548 1377
rect 1542 1372 1543 1376
rect 1547 1372 1548 1376
rect 1542 1371 1548 1372
rect 1630 1376 1636 1377
rect 1630 1372 1631 1376
rect 1635 1372 1636 1376
rect 1630 1371 1636 1372
rect 1718 1376 1724 1377
rect 1718 1372 1719 1376
rect 1723 1372 1724 1376
rect 1718 1371 1724 1372
rect 1798 1376 1804 1377
rect 1798 1372 1799 1376
rect 1803 1372 1804 1376
rect 1798 1371 1804 1372
rect 1870 1376 1876 1377
rect 1870 1372 1871 1376
rect 1875 1372 1876 1376
rect 1870 1371 1876 1372
rect 1942 1376 1948 1377
rect 1942 1372 1943 1376
rect 1947 1372 1948 1376
rect 1942 1371 1948 1372
rect 2014 1376 2020 1377
rect 2014 1372 2015 1376
rect 2019 1372 2020 1376
rect 2014 1371 2020 1372
rect 2070 1376 2076 1377
rect 2070 1372 2071 1376
rect 2075 1372 2076 1376
rect 2070 1371 2076 1372
rect 427 1367 433 1368
rect 427 1363 428 1367
rect 432 1366 433 1367
rect 442 1367 448 1368
rect 442 1366 443 1367
rect 432 1364 443 1366
rect 432 1363 433 1364
rect 427 1362 433 1363
rect 442 1363 443 1364
rect 447 1363 448 1367
rect 442 1362 448 1363
rect 458 1367 464 1368
rect 458 1363 459 1367
rect 463 1366 464 1367
rect 467 1367 473 1368
rect 467 1366 468 1367
rect 463 1364 468 1366
rect 463 1363 464 1364
rect 458 1362 464 1363
rect 467 1363 468 1364
rect 472 1363 473 1367
rect 467 1362 473 1363
rect 510 1367 521 1368
rect 510 1363 511 1367
rect 515 1363 516 1367
rect 520 1363 521 1367
rect 510 1362 521 1363
rect 566 1367 577 1368
rect 566 1363 567 1367
rect 571 1363 572 1367
rect 576 1363 577 1367
rect 566 1362 577 1363
rect 622 1367 633 1368
rect 622 1363 623 1367
rect 627 1363 628 1367
rect 632 1363 633 1367
rect 622 1362 633 1363
rect 691 1367 697 1368
rect 691 1363 692 1367
rect 696 1366 697 1367
rect 727 1367 733 1368
rect 727 1366 728 1367
rect 696 1364 728 1366
rect 696 1363 697 1364
rect 691 1362 697 1363
rect 727 1363 728 1364
rect 732 1363 733 1367
rect 727 1362 733 1363
rect 755 1367 761 1368
rect 755 1363 756 1367
rect 760 1366 761 1367
rect 791 1367 797 1368
rect 791 1366 792 1367
rect 760 1364 792 1366
rect 760 1363 761 1364
rect 755 1362 761 1363
rect 791 1363 792 1364
rect 796 1363 797 1367
rect 791 1362 797 1363
rect 819 1367 825 1368
rect 819 1363 820 1367
rect 824 1366 825 1367
rect 830 1367 836 1368
rect 830 1366 831 1367
rect 824 1364 831 1366
rect 824 1363 825 1364
rect 819 1362 825 1363
rect 830 1363 831 1364
rect 835 1363 836 1367
rect 830 1362 836 1363
rect 886 1367 897 1368
rect 886 1363 887 1367
rect 891 1363 892 1367
rect 896 1363 897 1367
rect 886 1362 897 1363
rect 958 1367 969 1368
rect 958 1363 959 1367
rect 963 1363 964 1367
rect 968 1363 969 1367
rect 958 1362 969 1363
rect 1155 1363 1161 1364
rect 1155 1359 1156 1363
rect 1160 1359 1161 1363
rect 1155 1358 1161 1359
rect 1186 1363 1192 1364
rect 1186 1359 1187 1363
rect 1191 1362 1192 1363
rect 1195 1363 1201 1364
rect 1195 1362 1196 1363
rect 1191 1360 1196 1362
rect 1191 1359 1192 1360
rect 1186 1358 1192 1359
rect 1195 1359 1196 1360
rect 1200 1359 1201 1363
rect 1195 1358 1201 1359
rect 1254 1363 1265 1364
rect 1254 1359 1255 1363
rect 1259 1359 1260 1363
rect 1264 1359 1265 1363
rect 1254 1358 1265 1359
rect 1342 1363 1353 1364
rect 1342 1359 1343 1363
rect 1347 1359 1348 1363
rect 1352 1359 1353 1363
rect 1342 1358 1353 1359
rect 1438 1363 1449 1364
rect 1438 1359 1439 1363
rect 1443 1359 1444 1363
rect 1448 1359 1449 1363
rect 1438 1358 1449 1359
rect 1534 1363 1545 1364
rect 1534 1359 1535 1363
rect 1539 1359 1540 1363
rect 1544 1359 1545 1363
rect 1534 1358 1545 1359
rect 1627 1363 1633 1364
rect 1627 1359 1628 1363
rect 1632 1362 1633 1363
rect 1670 1363 1676 1364
rect 1670 1362 1671 1363
rect 1632 1360 1671 1362
rect 1632 1359 1633 1360
rect 1627 1358 1633 1359
rect 1670 1359 1671 1360
rect 1675 1359 1676 1363
rect 1670 1358 1676 1359
rect 1710 1363 1721 1364
rect 1710 1359 1711 1363
rect 1715 1359 1716 1363
rect 1720 1359 1721 1363
rect 1710 1358 1721 1359
rect 1790 1363 1801 1364
rect 1790 1359 1791 1363
rect 1795 1359 1796 1363
rect 1800 1359 1801 1363
rect 1790 1358 1801 1359
rect 1862 1363 1873 1364
rect 1862 1359 1863 1363
rect 1867 1359 1868 1363
rect 1872 1359 1873 1363
rect 1862 1358 1873 1359
rect 1878 1363 1884 1364
rect 1878 1359 1879 1363
rect 1883 1362 1884 1363
rect 1939 1363 1945 1364
rect 1939 1362 1940 1363
rect 1883 1360 1940 1362
rect 1883 1359 1884 1360
rect 1878 1358 1884 1359
rect 1939 1359 1940 1360
rect 1944 1359 1945 1363
rect 1939 1358 1945 1359
rect 2006 1363 2017 1364
rect 2006 1359 2007 1363
rect 2011 1359 2012 1363
rect 2016 1359 2017 1363
rect 2006 1358 2017 1359
rect 2067 1363 2073 1364
rect 2067 1359 2068 1363
rect 2072 1362 2073 1363
rect 2090 1363 2096 1364
rect 2090 1362 2091 1363
rect 2072 1360 2091 1362
rect 2072 1359 2073 1360
rect 2067 1358 2073 1359
rect 2090 1359 2091 1360
rect 2095 1359 2096 1363
rect 2090 1358 2096 1359
rect 371 1355 377 1356
rect 371 1351 372 1355
rect 376 1354 377 1355
rect 382 1355 388 1356
rect 382 1354 383 1355
rect 376 1352 383 1354
rect 376 1351 377 1352
rect 371 1350 377 1351
rect 382 1351 383 1352
rect 387 1351 388 1355
rect 382 1350 388 1351
rect 402 1355 408 1356
rect 402 1351 403 1355
rect 407 1354 408 1355
rect 419 1355 425 1356
rect 419 1354 420 1355
rect 407 1352 420 1354
rect 407 1351 408 1352
rect 402 1350 408 1351
rect 419 1351 420 1352
rect 424 1351 425 1355
rect 419 1350 425 1351
rect 450 1355 456 1356
rect 450 1351 451 1355
rect 455 1354 456 1355
rect 475 1355 481 1356
rect 475 1354 476 1355
rect 455 1352 476 1354
rect 455 1351 456 1352
rect 450 1350 456 1351
rect 475 1351 476 1352
rect 480 1351 481 1355
rect 475 1350 481 1351
rect 506 1355 512 1356
rect 506 1351 507 1355
rect 511 1354 512 1355
rect 539 1355 545 1356
rect 539 1354 540 1355
rect 511 1352 540 1354
rect 511 1351 512 1352
rect 506 1350 512 1351
rect 539 1351 540 1352
rect 544 1351 545 1355
rect 539 1350 545 1351
rect 586 1355 592 1356
rect 586 1351 587 1355
rect 591 1354 592 1355
rect 603 1355 609 1356
rect 603 1354 604 1355
rect 591 1352 604 1354
rect 591 1351 592 1352
rect 586 1350 592 1351
rect 603 1351 604 1352
rect 608 1351 609 1355
rect 603 1350 609 1351
rect 667 1355 673 1356
rect 667 1351 668 1355
rect 672 1354 673 1355
rect 702 1355 708 1356
rect 702 1354 703 1355
rect 672 1352 703 1354
rect 672 1351 673 1352
rect 667 1350 673 1351
rect 702 1351 703 1352
rect 707 1351 708 1355
rect 702 1350 708 1351
rect 711 1355 717 1356
rect 711 1351 712 1355
rect 716 1354 717 1355
rect 731 1355 737 1356
rect 731 1354 732 1355
rect 716 1352 732 1354
rect 716 1351 717 1352
rect 711 1350 717 1351
rect 731 1351 732 1352
rect 736 1351 737 1355
rect 795 1355 801 1356
rect 795 1354 796 1355
rect 760 1352 796 1354
rect 731 1350 737 1351
rect 758 1351 764 1352
rect 758 1347 759 1351
rect 763 1347 764 1351
rect 795 1351 796 1352
rect 800 1351 801 1355
rect 795 1350 801 1351
rect 834 1355 840 1356
rect 834 1351 835 1355
rect 839 1354 840 1355
rect 859 1355 865 1356
rect 859 1354 860 1355
rect 839 1352 860 1354
rect 839 1351 840 1352
rect 834 1350 840 1351
rect 859 1351 860 1352
rect 864 1351 865 1355
rect 859 1350 865 1351
rect 923 1355 929 1356
rect 923 1351 924 1355
rect 928 1354 929 1355
rect 982 1355 988 1356
rect 982 1354 983 1355
rect 928 1352 983 1354
rect 928 1351 929 1352
rect 923 1350 929 1351
rect 982 1351 983 1352
rect 987 1351 988 1355
rect 982 1350 988 1351
rect 990 1355 1001 1356
rect 990 1351 991 1355
rect 995 1351 996 1355
rect 1000 1351 1001 1355
rect 990 1350 1001 1351
rect 1043 1355 1049 1356
rect 1043 1351 1044 1355
rect 1048 1354 1049 1355
rect 1070 1355 1076 1356
rect 1070 1354 1071 1355
rect 1048 1352 1071 1354
rect 1048 1351 1049 1352
rect 1043 1350 1049 1351
rect 1070 1351 1071 1352
rect 1075 1351 1076 1355
rect 1159 1354 1161 1358
rect 1510 1355 1516 1356
rect 1510 1354 1511 1355
rect 1159 1352 1511 1354
rect 1070 1350 1076 1351
rect 1510 1351 1511 1352
rect 1515 1351 1516 1355
rect 1886 1355 1892 1356
rect 1886 1354 1887 1355
rect 1510 1350 1516 1351
rect 1588 1352 1887 1354
rect 1588 1350 1590 1352
rect 1886 1351 1887 1352
rect 1891 1351 1892 1355
rect 1990 1355 1996 1356
rect 1990 1354 1991 1355
rect 1886 1350 1892 1351
rect 1900 1352 1991 1354
rect 1900 1350 1902 1352
rect 1990 1351 1991 1352
rect 1995 1351 1996 1355
rect 1990 1350 1996 1351
rect 1587 1349 1593 1350
rect 758 1346 764 1347
rect 1155 1347 1161 1348
rect 1155 1346 1156 1347
rect 374 1344 380 1345
rect 374 1340 375 1344
rect 379 1340 380 1344
rect 374 1339 380 1340
rect 422 1344 428 1345
rect 422 1340 423 1344
rect 427 1340 428 1344
rect 478 1344 484 1345
rect 478 1340 479 1344
rect 483 1340 484 1344
rect 422 1339 428 1340
rect 442 1339 448 1340
rect 478 1339 484 1340
rect 542 1344 548 1345
rect 542 1340 543 1344
rect 547 1340 548 1344
rect 542 1339 548 1340
rect 606 1344 612 1345
rect 606 1340 607 1344
rect 611 1340 612 1344
rect 606 1339 612 1340
rect 670 1344 676 1345
rect 670 1340 671 1344
rect 675 1340 676 1344
rect 670 1339 676 1340
rect 734 1344 740 1345
rect 734 1340 735 1344
rect 739 1340 740 1344
rect 734 1339 740 1340
rect 798 1344 804 1345
rect 798 1340 799 1344
rect 803 1340 804 1344
rect 798 1339 804 1340
rect 862 1344 868 1345
rect 862 1340 863 1344
rect 867 1340 868 1344
rect 862 1339 868 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1046 1339 1052 1340
rect 1088 1344 1156 1346
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 442 1335 443 1339
rect 447 1338 448 1339
rect 447 1336 474 1338
rect 447 1335 448 1336
rect 442 1334 448 1335
rect 472 1334 474 1336
rect 496 1336 538 1338
rect 496 1334 498 1336
rect 472 1332 498 1334
rect 536 1334 538 1336
rect 560 1336 598 1338
rect 560 1334 562 1336
rect 536 1332 562 1334
rect 110 1331 116 1332
rect 399 1331 408 1332
rect 399 1327 400 1331
rect 407 1327 408 1331
rect 399 1326 408 1327
rect 447 1331 456 1332
rect 447 1327 448 1331
rect 455 1327 456 1331
rect 447 1326 456 1327
rect 503 1331 512 1332
rect 503 1327 504 1331
rect 511 1327 512 1331
rect 503 1326 512 1327
rect 567 1331 573 1332
rect 567 1327 568 1331
rect 572 1330 573 1331
rect 586 1331 592 1332
rect 586 1330 587 1331
rect 572 1328 587 1330
rect 572 1327 573 1328
rect 567 1326 573 1327
rect 586 1327 587 1328
rect 591 1327 592 1331
rect 596 1330 598 1336
rect 631 1331 637 1332
rect 631 1330 632 1331
rect 596 1328 632 1330
rect 586 1326 592 1327
rect 631 1327 632 1328
rect 636 1327 637 1331
rect 631 1326 637 1327
rect 695 1331 701 1332
rect 695 1327 696 1331
rect 700 1330 701 1331
rect 711 1331 717 1332
rect 711 1330 712 1331
rect 700 1328 712 1330
rect 700 1327 701 1328
rect 695 1326 701 1327
rect 711 1327 712 1328
rect 716 1327 717 1331
rect 711 1326 717 1327
rect 758 1331 765 1332
rect 758 1327 759 1331
rect 764 1327 765 1331
rect 758 1326 765 1327
rect 823 1331 829 1332
rect 823 1327 824 1331
rect 828 1330 829 1331
rect 834 1331 840 1332
rect 834 1330 835 1331
rect 828 1328 835 1330
rect 828 1327 829 1328
rect 823 1326 829 1327
rect 834 1327 835 1328
rect 839 1327 840 1331
rect 834 1326 840 1327
rect 842 1331 848 1332
rect 842 1327 843 1331
rect 847 1330 848 1331
rect 887 1331 893 1332
rect 887 1330 888 1331
rect 847 1328 888 1330
rect 847 1327 848 1328
rect 842 1326 848 1327
rect 887 1327 888 1328
rect 892 1327 893 1331
rect 887 1326 893 1327
rect 951 1331 957 1332
rect 951 1327 952 1331
rect 956 1330 957 1331
rect 974 1331 980 1332
rect 974 1330 975 1331
rect 956 1328 975 1330
rect 956 1327 957 1328
rect 951 1326 957 1327
rect 974 1327 975 1328
rect 979 1327 980 1331
rect 974 1326 980 1327
rect 982 1331 988 1332
rect 982 1327 983 1331
rect 987 1330 988 1331
rect 1023 1331 1029 1332
rect 1023 1330 1024 1331
rect 987 1328 1024 1330
rect 987 1327 988 1328
rect 982 1326 988 1327
rect 1023 1327 1024 1328
rect 1028 1327 1029 1331
rect 1023 1326 1029 1327
rect 1071 1331 1077 1332
rect 1071 1327 1072 1331
rect 1076 1330 1077 1331
rect 1088 1330 1090 1344
rect 1155 1343 1156 1344
rect 1160 1343 1161 1347
rect 1155 1342 1161 1343
rect 1186 1347 1192 1348
rect 1186 1343 1187 1347
rect 1191 1346 1192 1347
rect 1251 1347 1257 1348
rect 1251 1346 1252 1347
rect 1191 1344 1252 1346
rect 1191 1343 1192 1344
rect 1186 1342 1192 1343
rect 1251 1343 1252 1344
rect 1256 1343 1257 1347
rect 1251 1342 1257 1343
rect 1282 1347 1288 1348
rect 1282 1343 1283 1347
rect 1287 1346 1288 1347
rect 1371 1347 1377 1348
rect 1371 1346 1372 1347
rect 1287 1344 1372 1346
rect 1287 1343 1288 1344
rect 1282 1342 1288 1343
rect 1371 1343 1372 1344
rect 1376 1343 1377 1347
rect 1371 1342 1377 1343
rect 1402 1347 1408 1348
rect 1402 1343 1403 1347
rect 1407 1346 1408 1347
rect 1483 1347 1489 1348
rect 1483 1346 1484 1347
rect 1407 1344 1484 1346
rect 1407 1343 1408 1344
rect 1402 1342 1408 1343
rect 1483 1343 1484 1344
rect 1488 1343 1489 1347
rect 1587 1345 1588 1349
rect 1592 1345 1593 1349
rect 1899 1349 1905 1350
rect 1587 1344 1593 1345
rect 1618 1347 1624 1348
rect 1483 1342 1489 1343
rect 1618 1343 1619 1347
rect 1623 1346 1624 1347
rect 1675 1347 1681 1348
rect 1675 1346 1676 1347
rect 1623 1344 1676 1346
rect 1623 1343 1624 1344
rect 1618 1342 1624 1343
rect 1675 1343 1676 1344
rect 1680 1343 1681 1347
rect 1675 1342 1681 1343
rect 1706 1347 1712 1348
rect 1706 1343 1707 1347
rect 1711 1346 1712 1347
rect 1755 1347 1761 1348
rect 1755 1346 1756 1347
rect 1711 1344 1756 1346
rect 1711 1343 1712 1344
rect 1706 1342 1712 1343
rect 1755 1343 1756 1344
rect 1760 1343 1761 1347
rect 1755 1342 1761 1343
rect 1786 1347 1792 1348
rect 1786 1343 1787 1347
rect 1791 1346 1792 1347
rect 1827 1347 1833 1348
rect 1827 1346 1828 1347
rect 1791 1344 1828 1346
rect 1791 1343 1792 1344
rect 1786 1342 1792 1343
rect 1827 1343 1828 1344
rect 1832 1343 1833 1347
rect 1899 1345 1900 1349
rect 1904 1345 1905 1349
rect 1899 1344 1905 1345
rect 1963 1347 1969 1348
rect 1827 1342 1833 1343
rect 1963 1343 1964 1347
rect 1968 1346 1969 1347
rect 2015 1347 2021 1348
rect 2015 1346 2016 1347
rect 1968 1344 2016 1346
rect 1968 1343 1969 1344
rect 1963 1342 1969 1343
rect 2015 1343 2016 1344
rect 2020 1343 2021 1347
rect 2015 1342 2021 1343
rect 2027 1347 2033 1348
rect 2027 1343 2028 1347
rect 2032 1346 2033 1347
rect 2046 1347 2052 1348
rect 2046 1346 2047 1347
rect 2032 1344 2047 1346
rect 2032 1343 2033 1344
rect 2027 1342 2033 1343
rect 2046 1343 2047 1344
rect 2051 1343 2052 1347
rect 2046 1342 2052 1343
rect 2067 1347 2073 1348
rect 2067 1343 2068 1347
rect 2072 1346 2073 1347
rect 2082 1347 2088 1348
rect 2082 1346 2083 1347
rect 2072 1344 2083 1346
rect 2072 1343 2073 1344
rect 2067 1342 2073 1343
rect 2082 1343 2083 1344
rect 2087 1343 2088 1347
rect 2082 1342 2088 1343
rect 1094 1336 1100 1337
rect 1094 1332 1095 1336
rect 1099 1332 1100 1336
rect 1094 1331 1100 1332
rect 1158 1336 1164 1337
rect 1158 1332 1159 1336
rect 1163 1332 1164 1336
rect 1158 1331 1164 1332
rect 1254 1336 1260 1337
rect 1254 1332 1255 1336
rect 1259 1332 1260 1336
rect 1254 1331 1260 1332
rect 1374 1336 1380 1337
rect 1374 1332 1375 1336
rect 1379 1332 1380 1336
rect 1374 1331 1380 1332
rect 1486 1336 1492 1337
rect 1486 1332 1487 1336
rect 1491 1332 1492 1336
rect 1486 1331 1492 1332
rect 1590 1336 1596 1337
rect 1590 1332 1591 1336
rect 1595 1332 1596 1336
rect 1590 1331 1596 1332
rect 1678 1336 1684 1337
rect 1678 1332 1679 1336
rect 1683 1332 1684 1336
rect 1678 1331 1684 1332
rect 1758 1336 1764 1337
rect 1758 1332 1759 1336
rect 1763 1332 1764 1336
rect 1758 1331 1764 1332
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 1902 1336 1908 1337
rect 1902 1332 1903 1336
rect 1907 1332 1908 1336
rect 1902 1331 1908 1332
rect 1966 1336 1972 1337
rect 1966 1332 1967 1336
rect 1971 1332 1972 1336
rect 1966 1331 1972 1332
rect 2030 1336 2036 1337
rect 2030 1332 2031 1336
rect 2035 1332 2036 1336
rect 2030 1331 2036 1332
rect 2070 1336 2076 1337
rect 2070 1332 2071 1336
rect 2075 1332 2076 1336
rect 2070 1331 2076 1332
rect 1076 1328 1090 1330
rect 1134 1328 1140 1329
rect 1076 1327 1077 1328
rect 1071 1326 1077 1327
rect 1134 1324 1135 1328
rect 1139 1324 1140 1328
rect 2118 1328 2124 1329
rect 2118 1324 2119 1328
rect 2123 1324 2124 1328
rect 1134 1323 1140 1324
rect 1183 1323 1192 1324
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 1094 1319 1100 1320
rect 110 1314 116 1315
rect 374 1316 380 1317
rect 374 1312 375 1316
rect 379 1312 380 1316
rect 374 1311 380 1312
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 478 1316 484 1317
rect 478 1312 479 1316
rect 483 1312 484 1316
rect 478 1311 484 1312
rect 542 1316 548 1317
rect 542 1312 543 1316
rect 547 1312 548 1316
rect 542 1311 548 1312
rect 606 1316 612 1317
rect 606 1312 607 1316
rect 611 1312 612 1316
rect 606 1311 612 1312
rect 670 1316 676 1317
rect 670 1312 671 1316
rect 675 1312 676 1316
rect 670 1311 676 1312
rect 734 1316 740 1317
rect 734 1312 735 1316
rect 739 1312 740 1316
rect 734 1311 740 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 998 1316 1004 1317
rect 998 1312 999 1316
rect 1003 1312 1004 1316
rect 998 1311 1004 1312
rect 1046 1316 1052 1317
rect 1046 1312 1047 1316
rect 1051 1312 1052 1316
rect 1094 1315 1095 1319
rect 1099 1315 1100 1319
rect 1183 1319 1184 1323
rect 1191 1319 1192 1323
rect 1183 1318 1192 1319
rect 1279 1323 1288 1324
rect 1279 1319 1280 1323
rect 1287 1319 1288 1323
rect 1279 1318 1288 1319
rect 1399 1323 1408 1324
rect 1399 1319 1400 1323
rect 1407 1319 1408 1323
rect 1399 1318 1408 1319
rect 1510 1323 1517 1324
rect 1510 1319 1511 1323
rect 1516 1319 1517 1323
rect 1510 1318 1517 1319
rect 1615 1323 1624 1324
rect 1615 1319 1616 1323
rect 1623 1319 1624 1323
rect 1615 1318 1624 1319
rect 1703 1323 1712 1324
rect 1703 1319 1704 1323
rect 1711 1319 1712 1323
rect 1703 1318 1712 1319
rect 1783 1323 1792 1324
rect 1783 1319 1784 1323
rect 1791 1319 1792 1323
rect 1783 1318 1792 1319
rect 1855 1323 1861 1324
rect 1855 1319 1856 1323
rect 1860 1322 1861 1323
rect 1878 1323 1884 1324
rect 1878 1322 1879 1323
rect 1860 1320 1879 1322
rect 1860 1319 1861 1320
rect 1855 1318 1861 1319
rect 1878 1319 1879 1320
rect 1883 1319 1884 1323
rect 1878 1318 1884 1319
rect 1927 1323 1933 1324
rect 1927 1319 1928 1323
rect 1932 1322 1933 1323
rect 1958 1323 1964 1324
rect 1958 1322 1959 1323
rect 1932 1320 1959 1322
rect 1932 1319 1933 1320
rect 1927 1318 1933 1319
rect 1958 1319 1959 1320
rect 1963 1319 1964 1323
rect 1958 1318 1964 1319
rect 1990 1323 1997 1324
rect 1990 1319 1991 1323
rect 1996 1319 1997 1323
rect 1990 1318 1997 1319
rect 2015 1323 2021 1324
rect 2015 1319 2016 1323
rect 2020 1322 2021 1323
rect 2055 1323 2061 1324
rect 2055 1322 2056 1323
rect 2020 1320 2056 1322
rect 2020 1319 2021 1320
rect 2015 1318 2021 1319
rect 2055 1319 2056 1320
rect 2060 1319 2061 1323
rect 2055 1318 2061 1319
rect 2082 1323 2088 1324
rect 2082 1319 2083 1323
rect 2087 1322 2088 1323
rect 2095 1323 2101 1324
rect 2118 1323 2124 1324
rect 2095 1322 2096 1323
rect 2087 1320 2096 1322
rect 2087 1319 2088 1320
rect 2082 1318 2088 1319
rect 2095 1319 2096 1320
rect 2100 1319 2101 1323
rect 2095 1318 2101 1319
rect 1094 1314 1100 1315
rect 1046 1311 1052 1312
rect 1134 1311 1140 1312
rect 1134 1307 1135 1311
rect 1139 1307 1140 1311
rect 2118 1311 2124 1312
rect 1134 1306 1140 1307
rect 1158 1308 1164 1309
rect 334 1304 340 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 334 1300 335 1304
rect 339 1300 340 1304
rect 334 1299 340 1300
rect 390 1304 396 1305
rect 390 1300 391 1304
rect 395 1300 396 1304
rect 390 1299 396 1300
rect 454 1304 460 1305
rect 454 1300 455 1304
rect 459 1300 460 1304
rect 454 1299 460 1300
rect 526 1304 532 1305
rect 526 1300 527 1304
rect 531 1300 532 1304
rect 526 1299 532 1300
rect 598 1304 604 1305
rect 598 1300 599 1304
rect 603 1300 604 1304
rect 598 1299 604 1300
rect 670 1304 676 1305
rect 670 1300 671 1304
rect 675 1300 676 1304
rect 670 1299 676 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 822 1304 828 1305
rect 822 1300 823 1304
rect 827 1300 828 1304
rect 822 1299 828 1300
rect 902 1304 908 1305
rect 902 1300 903 1304
rect 907 1300 908 1304
rect 902 1299 908 1300
rect 982 1304 988 1305
rect 982 1300 983 1304
rect 987 1300 988 1304
rect 982 1299 988 1300
rect 1046 1304 1052 1305
rect 1046 1300 1047 1304
rect 1051 1300 1052 1304
rect 1158 1304 1159 1308
rect 1163 1304 1164 1308
rect 1158 1303 1164 1304
rect 1254 1308 1260 1309
rect 1254 1304 1255 1308
rect 1259 1304 1260 1308
rect 1254 1303 1260 1304
rect 1374 1308 1380 1309
rect 1374 1304 1375 1308
rect 1379 1304 1380 1308
rect 1374 1303 1380 1304
rect 1486 1308 1492 1309
rect 1486 1304 1487 1308
rect 1491 1304 1492 1308
rect 1486 1303 1492 1304
rect 1590 1308 1596 1309
rect 1590 1304 1591 1308
rect 1595 1304 1596 1308
rect 1590 1303 1596 1304
rect 1678 1308 1684 1309
rect 1678 1304 1679 1308
rect 1683 1304 1684 1308
rect 1678 1303 1684 1304
rect 1758 1308 1764 1309
rect 1758 1304 1759 1308
rect 1763 1304 1764 1308
rect 1758 1303 1764 1304
rect 1830 1308 1836 1309
rect 1830 1304 1831 1308
rect 1835 1304 1836 1308
rect 1830 1303 1836 1304
rect 1902 1308 1908 1309
rect 1902 1304 1903 1308
rect 1907 1304 1908 1308
rect 1902 1303 1908 1304
rect 1966 1308 1972 1309
rect 1966 1304 1967 1308
rect 1971 1304 1972 1308
rect 1966 1303 1972 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2030 1303 2036 1304
rect 2070 1308 2076 1309
rect 2070 1304 2071 1308
rect 2075 1304 2076 1308
rect 2118 1307 2119 1311
rect 2123 1307 2124 1311
rect 2118 1306 2124 1307
rect 2070 1303 2076 1304
rect 1046 1299 1052 1300
rect 1094 1301 1100 1302
rect 110 1296 116 1297
rect 1094 1297 1095 1301
rect 1099 1297 1100 1301
rect 1094 1296 1100 1297
rect 382 1295 388 1296
rect 382 1291 383 1295
rect 387 1294 388 1295
rect 387 1292 602 1294
rect 387 1291 388 1292
rect 382 1290 388 1291
rect 359 1287 365 1288
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 359 1283 360 1287
rect 364 1286 365 1287
rect 382 1287 388 1288
rect 382 1286 383 1287
rect 364 1284 383 1286
rect 364 1283 365 1284
rect 359 1282 365 1283
rect 382 1283 383 1284
rect 387 1283 388 1287
rect 382 1282 388 1283
rect 415 1287 421 1288
rect 415 1283 416 1287
rect 420 1286 421 1287
rect 446 1287 452 1288
rect 446 1286 447 1287
rect 420 1284 447 1286
rect 420 1283 421 1284
rect 415 1282 421 1283
rect 446 1283 447 1284
rect 451 1283 452 1287
rect 446 1282 452 1283
rect 479 1287 485 1288
rect 479 1283 480 1287
rect 484 1286 485 1287
rect 518 1287 524 1288
rect 518 1286 519 1287
rect 484 1284 519 1286
rect 484 1283 485 1284
rect 479 1282 485 1283
rect 518 1283 519 1284
rect 523 1283 524 1287
rect 518 1282 524 1283
rect 551 1287 557 1288
rect 551 1283 552 1287
rect 556 1286 557 1287
rect 590 1287 596 1288
rect 590 1286 591 1287
rect 556 1284 591 1286
rect 556 1283 557 1284
rect 551 1282 557 1283
rect 590 1283 591 1284
rect 595 1283 596 1287
rect 600 1286 602 1292
rect 1158 1292 1164 1293
rect 1134 1289 1140 1290
rect 623 1287 629 1288
rect 623 1286 624 1287
rect 600 1284 624 1286
rect 590 1282 596 1283
rect 623 1283 624 1284
rect 628 1283 629 1287
rect 623 1282 629 1283
rect 695 1287 701 1288
rect 695 1283 696 1287
rect 700 1286 701 1287
rect 734 1287 740 1288
rect 734 1286 735 1287
rect 700 1284 735 1286
rect 700 1283 701 1284
rect 695 1282 701 1283
rect 734 1283 735 1284
rect 739 1283 740 1287
rect 734 1282 740 1283
rect 767 1287 773 1288
rect 767 1283 768 1287
rect 772 1286 773 1287
rect 790 1287 796 1288
rect 790 1286 791 1287
rect 772 1284 791 1286
rect 772 1283 773 1284
rect 767 1282 773 1283
rect 790 1283 791 1284
rect 795 1283 796 1287
rect 790 1282 796 1283
rect 799 1287 805 1288
rect 799 1283 800 1287
rect 804 1286 805 1287
rect 847 1287 853 1288
rect 847 1286 848 1287
rect 804 1284 848 1286
rect 804 1283 805 1284
rect 799 1282 805 1283
rect 847 1283 848 1284
rect 852 1283 853 1287
rect 847 1282 853 1283
rect 918 1287 924 1288
rect 918 1283 919 1287
rect 923 1286 924 1287
rect 927 1287 933 1288
rect 927 1286 928 1287
rect 923 1284 928 1286
rect 923 1283 924 1284
rect 918 1282 924 1283
rect 927 1283 928 1284
rect 932 1283 933 1287
rect 927 1282 933 1283
rect 935 1287 941 1288
rect 935 1283 936 1287
rect 940 1286 941 1287
rect 1007 1287 1013 1288
rect 1007 1286 1008 1287
rect 940 1284 1008 1286
rect 940 1283 941 1284
rect 935 1282 941 1283
rect 1007 1283 1008 1284
rect 1012 1283 1013 1287
rect 1007 1282 1013 1283
rect 1070 1287 1077 1288
rect 1070 1283 1071 1287
rect 1076 1283 1077 1287
rect 1134 1285 1135 1289
rect 1139 1285 1140 1289
rect 1158 1288 1159 1292
rect 1163 1288 1164 1292
rect 1158 1287 1164 1288
rect 1198 1292 1204 1293
rect 1198 1288 1199 1292
rect 1203 1288 1204 1292
rect 1198 1287 1204 1288
rect 1246 1292 1252 1293
rect 1246 1288 1247 1292
rect 1251 1288 1252 1292
rect 1246 1287 1252 1288
rect 1318 1292 1324 1293
rect 1318 1288 1319 1292
rect 1323 1288 1324 1292
rect 1318 1287 1324 1288
rect 1398 1292 1404 1293
rect 1398 1288 1399 1292
rect 1403 1288 1404 1292
rect 1398 1287 1404 1288
rect 1478 1292 1484 1293
rect 1478 1288 1479 1292
rect 1483 1288 1484 1292
rect 1478 1287 1484 1288
rect 1558 1292 1564 1293
rect 1558 1288 1559 1292
rect 1563 1288 1564 1292
rect 1558 1287 1564 1288
rect 1638 1292 1644 1293
rect 1638 1288 1639 1292
rect 1643 1288 1644 1292
rect 1638 1287 1644 1288
rect 1718 1292 1724 1293
rect 1718 1288 1719 1292
rect 1723 1288 1724 1292
rect 1718 1287 1724 1288
rect 1798 1292 1804 1293
rect 1798 1288 1799 1292
rect 1803 1288 1804 1292
rect 1798 1287 1804 1288
rect 1878 1292 1884 1293
rect 1878 1288 1879 1292
rect 1883 1288 1884 1292
rect 1878 1287 1884 1288
rect 1966 1292 1972 1293
rect 1966 1288 1967 1292
rect 1971 1288 1972 1292
rect 1966 1287 1972 1288
rect 2054 1292 2060 1293
rect 2054 1288 2055 1292
rect 2059 1288 2060 1292
rect 2054 1287 2060 1288
rect 2118 1289 2124 1290
rect 1070 1282 1077 1283
rect 1094 1284 1100 1285
rect 1134 1284 1140 1285
rect 2118 1285 2119 1289
rect 2123 1285 2124 1289
rect 2118 1284 2124 1285
rect 110 1279 116 1280
rect 1094 1280 1095 1284
rect 1099 1280 1100 1284
rect 1094 1279 1100 1280
rect 1270 1283 1276 1284
rect 1270 1279 1271 1283
rect 1275 1282 1276 1283
rect 1275 1280 1482 1282
rect 1275 1279 1276 1280
rect 1270 1278 1276 1279
rect 334 1276 340 1277
rect 334 1272 335 1276
rect 339 1272 340 1276
rect 334 1271 340 1272
rect 390 1276 396 1277
rect 390 1272 391 1276
rect 395 1272 396 1276
rect 390 1271 396 1272
rect 454 1276 460 1277
rect 454 1272 455 1276
rect 459 1272 460 1276
rect 454 1271 460 1272
rect 526 1276 532 1277
rect 526 1272 527 1276
rect 531 1272 532 1276
rect 526 1271 532 1272
rect 598 1276 604 1277
rect 598 1272 599 1276
rect 603 1272 604 1276
rect 598 1271 604 1272
rect 670 1276 676 1277
rect 670 1272 671 1276
rect 675 1272 676 1276
rect 670 1271 676 1272
rect 742 1276 748 1277
rect 742 1272 743 1276
rect 747 1272 748 1276
rect 742 1271 748 1272
rect 822 1276 828 1277
rect 822 1272 823 1276
rect 827 1272 828 1276
rect 822 1271 828 1272
rect 902 1276 908 1277
rect 902 1272 903 1276
rect 907 1272 908 1276
rect 902 1271 908 1272
rect 982 1276 988 1277
rect 982 1272 983 1276
rect 987 1272 988 1276
rect 982 1271 988 1272
rect 1046 1276 1052 1277
rect 1046 1272 1047 1276
rect 1051 1272 1052 1276
rect 1183 1275 1189 1276
rect 1183 1274 1184 1275
rect 1046 1271 1052 1272
rect 1134 1272 1140 1273
rect 1134 1268 1135 1272
rect 1139 1268 1140 1272
rect 1134 1267 1140 1268
rect 1144 1272 1184 1274
rect 331 1263 337 1264
rect 331 1259 332 1263
rect 336 1262 337 1263
rect 382 1263 393 1264
rect 336 1260 378 1262
rect 336 1259 337 1260
rect 331 1258 337 1259
rect 376 1254 378 1260
rect 382 1259 383 1263
rect 387 1259 388 1263
rect 392 1259 393 1263
rect 382 1258 393 1259
rect 446 1263 457 1264
rect 446 1259 447 1263
rect 451 1259 452 1263
rect 456 1259 457 1263
rect 446 1258 457 1259
rect 518 1263 529 1264
rect 518 1259 519 1263
rect 523 1259 524 1263
rect 528 1259 529 1263
rect 518 1258 529 1259
rect 590 1263 601 1264
rect 590 1259 591 1263
rect 595 1259 596 1263
rect 600 1259 601 1263
rect 590 1258 601 1259
rect 667 1263 673 1264
rect 667 1259 668 1263
rect 672 1262 673 1263
rect 734 1263 745 1264
rect 672 1260 681 1262
rect 672 1259 673 1260
rect 667 1258 673 1259
rect 566 1255 572 1256
rect 566 1254 567 1255
rect 376 1252 567 1254
rect 566 1251 567 1252
rect 571 1251 572 1255
rect 679 1254 681 1260
rect 734 1259 735 1263
rect 739 1259 740 1263
rect 744 1259 745 1263
rect 734 1258 745 1259
rect 819 1263 825 1264
rect 819 1259 820 1263
rect 824 1262 825 1263
rect 842 1263 848 1264
rect 842 1262 843 1263
rect 824 1260 843 1262
rect 824 1259 825 1260
rect 819 1258 825 1259
rect 842 1259 843 1260
rect 847 1259 848 1263
rect 842 1258 848 1259
rect 899 1263 905 1264
rect 899 1259 900 1263
rect 904 1262 905 1263
rect 935 1263 941 1264
rect 935 1262 936 1263
rect 904 1260 936 1262
rect 904 1259 905 1260
rect 899 1258 905 1259
rect 935 1259 936 1260
rect 940 1259 941 1263
rect 935 1258 941 1259
rect 974 1263 985 1264
rect 974 1259 975 1263
rect 979 1259 980 1263
rect 984 1259 985 1263
rect 974 1258 985 1259
rect 1043 1263 1049 1264
rect 1043 1259 1044 1263
rect 1048 1262 1049 1263
rect 1144 1262 1146 1272
rect 1183 1271 1184 1272
rect 1188 1271 1189 1275
rect 1223 1275 1229 1276
rect 1223 1274 1224 1275
rect 1183 1270 1189 1271
rect 1192 1272 1224 1274
rect 1048 1260 1146 1262
rect 1158 1264 1164 1265
rect 1158 1260 1159 1264
rect 1163 1260 1164 1264
rect 1048 1259 1049 1260
rect 1158 1259 1164 1260
rect 1043 1258 1049 1259
rect 1192 1258 1194 1272
rect 1223 1271 1224 1272
rect 1228 1271 1229 1275
rect 1223 1270 1229 1271
rect 1231 1275 1237 1276
rect 1231 1271 1232 1275
rect 1236 1274 1237 1275
rect 1271 1275 1277 1276
rect 1271 1274 1272 1275
rect 1236 1272 1272 1274
rect 1236 1271 1237 1272
rect 1231 1270 1237 1271
rect 1271 1271 1272 1272
rect 1276 1271 1277 1275
rect 1271 1270 1277 1271
rect 1343 1275 1349 1276
rect 1343 1271 1344 1275
rect 1348 1274 1349 1275
rect 1390 1275 1396 1276
rect 1390 1274 1391 1275
rect 1348 1272 1391 1274
rect 1348 1271 1349 1272
rect 1343 1270 1349 1271
rect 1390 1271 1391 1272
rect 1395 1271 1396 1275
rect 1390 1270 1396 1271
rect 1423 1275 1429 1276
rect 1423 1271 1424 1275
rect 1428 1274 1429 1275
rect 1470 1275 1476 1276
rect 1470 1274 1471 1275
rect 1428 1272 1471 1274
rect 1428 1271 1429 1272
rect 1423 1270 1429 1271
rect 1470 1271 1471 1272
rect 1475 1271 1476 1275
rect 1480 1274 1482 1280
rect 1503 1275 1509 1276
rect 1503 1274 1504 1275
rect 1480 1272 1504 1274
rect 1470 1270 1476 1271
rect 1503 1271 1504 1272
rect 1508 1271 1509 1275
rect 1503 1270 1509 1271
rect 1583 1275 1589 1276
rect 1583 1271 1584 1275
rect 1588 1274 1589 1275
rect 1630 1275 1636 1276
rect 1630 1274 1631 1275
rect 1588 1272 1631 1274
rect 1588 1271 1589 1272
rect 1583 1270 1589 1271
rect 1630 1271 1631 1272
rect 1635 1271 1636 1275
rect 1630 1270 1636 1271
rect 1663 1275 1669 1276
rect 1663 1271 1664 1275
rect 1668 1274 1669 1275
rect 1710 1275 1716 1276
rect 1710 1274 1711 1275
rect 1668 1272 1711 1274
rect 1668 1271 1669 1272
rect 1663 1270 1669 1271
rect 1710 1271 1711 1272
rect 1715 1271 1716 1275
rect 1710 1270 1716 1271
rect 1743 1275 1749 1276
rect 1743 1271 1744 1275
rect 1748 1274 1749 1275
rect 1814 1275 1820 1276
rect 1814 1274 1815 1275
rect 1748 1272 1815 1274
rect 1748 1271 1749 1272
rect 1743 1270 1749 1271
rect 1814 1271 1815 1272
rect 1819 1271 1820 1275
rect 1814 1270 1820 1271
rect 1822 1275 1829 1276
rect 1822 1271 1823 1275
rect 1828 1271 1829 1275
rect 1822 1270 1829 1271
rect 1834 1275 1840 1276
rect 1834 1271 1835 1275
rect 1839 1274 1840 1275
rect 1903 1275 1909 1276
rect 1903 1274 1904 1275
rect 1839 1272 1904 1274
rect 1839 1271 1840 1272
rect 1834 1270 1840 1271
rect 1903 1271 1904 1272
rect 1908 1271 1909 1275
rect 1903 1270 1909 1271
rect 1911 1275 1917 1276
rect 1911 1271 1912 1275
rect 1916 1274 1917 1275
rect 1991 1275 1997 1276
rect 1991 1274 1992 1275
rect 1916 1272 1992 1274
rect 1916 1271 1917 1272
rect 1911 1270 1917 1271
rect 1991 1271 1992 1272
rect 1996 1271 1997 1275
rect 1991 1270 1997 1271
rect 2046 1275 2052 1276
rect 2046 1271 2047 1275
rect 2051 1274 2052 1275
rect 2079 1275 2085 1276
rect 2079 1274 2080 1275
rect 2051 1272 2080 1274
rect 2051 1271 2052 1272
rect 2046 1270 2052 1271
rect 2079 1271 2080 1272
rect 2084 1271 2085 1275
rect 2079 1270 2085 1271
rect 2118 1272 2124 1273
rect 2118 1268 2119 1272
rect 2123 1268 2124 1272
rect 2118 1267 2124 1268
rect 1198 1264 1204 1265
rect 1198 1260 1199 1264
rect 1203 1260 1204 1264
rect 1198 1259 1204 1260
rect 1246 1264 1252 1265
rect 1246 1260 1247 1264
rect 1251 1260 1252 1264
rect 1318 1264 1324 1265
rect 1318 1260 1319 1264
rect 1323 1260 1324 1264
rect 1246 1259 1252 1260
rect 1270 1259 1276 1260
rect 1318 1259 1324 1260
rect 1398 1264 1404 1265
rect 1398 1260 1399 1264
rect 1403 1260 1404 1264
rect 1398 1259 1404 1260
rect 1478 1264 1484 1265
rect 1478 1260 1479 1264
rect 1483 1260 1484 1264
rect 1478 1259 1484 1260
rect 1558 1264 1564 1265
rect 1558 1260 1559 1264
rect 1563 1260 1564 1264
rect 1558 1259 1564 1260
rect 1638 1264 1644 1265
rect 1638 1260 1639 1264
rect 1643 1260 1644 1264
rect 1638 1259 1644 1260
rect 1718 1264 1724 1265
rect 1718 1260 1719 1264
rect 1723 1260 1724 1264
rect 1718 1259 1724 1260
rect 1798 1264 1804 1265
rect 1798 1260 1799 1264
rect 1803 1260 1804 1264
rect 1798 1259 1804 1260
rect 1878 1264 1884 1265
rect 1878 1260 1879 1264
rect 1883 1260 1884 1264
rect 1878 1259 1884 1260
rect 1966 1264 1972 1265
rect 1966 1260 1967 1264
rect 1971 1260 1972 1264
rect 1966 1259 1972 1260
rect 2054 1264 2060 1265
rect 2054 1260 2055 1264
rect 2059 1260 2060 1264
rect 2054 1259 2060 1260
rect 1270 1258 1271 1259
rect 1188 1256 1194 1258
rect 1256 1256 1271 1258
rect 799 1255 805 1256
rect 799 1254 800 1255
rect 679 1252 800 1254
rect 566 1250 572 1251
rect 799 1251 800 1252
rect 804 1251 805 1255
rect 1188 1254 1190 1256
rect 1256 1254 1258 1256
rect 1270 1255 1271 1256
rect 1275 1255 1276 1259
rect 1270 1254 1276 1255
rect 799 1250 805 1251
rect 1155 1253 1190 1254
rect 1155 1249 1156 1253
rect 1160 1252 1190 1253
rect 1243 1253 1258 1254
rect 1160 1249 1161 1252
rect 1155 1248 1161 1249
rect 1195 1251 1201 1252
rect 259 1247 265 1248
rect 259 1243 260 1247
rect 264 1246 265 1247
rect 270 1247 276 1248
rect 270 1246 271 1247
rect 264 1244 271 1246
rect 264 1243 265 1244
rect 259 1242 265 1243
rect 270 1243 271 1244
rect 275 1243 276 1247
rect 270 1242 276 1243
rect 290 1247 296 1248
rect 290 1243 291 1247
rect 295 1246 296 1247
rect 307 1247 313 1248
rect 307 1246 308 1247
rect 295 1244 308 1246
rect 295 1243 296 1244
rect 290 1242 296 1243
rect 307 1243 308 1244
rect 312 1243 313 1247
rect 307 1242 313 1243
rect 355 1247 361 1248
rect 355 1243 356 1247
rect 360 1243 361 1247
rect 355 1242 361 1243
rect 391 1247 397 1248
rect 391 1243 392 1247
rect 396 1246 397 1247
rect 411 1247 417 1248
rect 411 1246 412 1247
rect 396 1244 412 1246
rect 396 1243 397 1244
rect 391 1242 397 1243
rect 411 1243 412 1244
rect 416 1243 417 1247
rect 411 1242 417 1243
rect 442 1247 448 1248
rect 442 1243 443 1247
rect 447 1246 448 1247
rect 475 1247 481 1248
rect 475 1246 476 1247
rect 447 1244 476 1246
rect 447 1243 448 1244
rect 442 1242 448 1243
rect 475 1243 476 1244
rect 480 1243 481 1247
rect 475 1242 481 1243
rect 518 1247 524 1248
rect 518 1243 519 1247
rect 523 1246 524 1247
rect 539 1247 545 1248
rect 539 1246 540 1247
rect 523 1244 540 1246
rect 523 1243 524 1244
rect 518 1242 524 1243
rect 539 1243 540 1244
rect 544 1243 545 1247
rect 539 1242 545 1243
rect 603 1247 609 1248
rect 603 1243 604 1247
rect 608 1246 609 1247
rect 639 1247 645 1248
rect 639 1246 640 1247
rect 608 1244 640 1246
rect 608 1243 609 1244
rect 603 1242 609 1243
rect 639 1243 640 1244
rect 644 1243 645 1247
rect 639 1242 645 1243
rect 667 1247 673 1248
rect 667 1243 668 1247
rect 672 1246 673 1247
rect 722 1247 728 1248
rect 722 1246 723 1247
rect 672 1244 723 1246
rect 672 1243 673 1244
rect 667 1242 673 1243
rect 722 1243 723 1244
rect 727 1243 728 1247
rect 722 1242 728 1243
rect 731 1247 737 1248
rect 731 1243 732 1247
rect 736 1246 737 1247
rect 782 1247 788 1248
rect 782 1246 783 1247
rect 736 1244 783 1246
rect 736 1243 737 1244
rect 731 1242 737 1243
rect 782 1243 783 1244
rect 787 1243 788 1247
rect 782 1242 788 1243
rect 790 1247 801 1248
rect 790 1243 791 1247
rect 795 1243 796 1247
rect 800 1243 801 1247
rect 790 1242 801 1243
rect 859 1247 865 1248
rect 859 1243 860 1247
rect 864 1246 865 1247
rect 910 1247 916 1248
rect 910 1246 911 1247
rect 864 1244 911 1246
rect 864 1243 865 1244
rect 859 1242 865 1243
rect 910 1243 911 1244
rect 915 1243 916 1247
rect 910 1242 916 1243
rect 918 1247 929 1248
rect 918 1243 919 1247
rect 923 1243 924 1247
rect 928 1243 929 1247
rect 1195 1247 1196 1251
rect 1200 1250 1201 1251
rect 1231 1251 1237 1252
rect 1231 1250 1232 1251
rect 1200 1248 1232 1250
rect 1200 1247 1201 1248
rect 1195 1246 1201 1247
rect 1231 1247 1232 1248
rect 1236 1247 1237 1251
rect 1243 1249 1244 1253
rect 1248 1252 1258 1253
rect 1248 1249 1249 1252
rect 1243 1248 1249 1249
rect 1266 1251 1272 1252
rect 1231 1246 1237 1247
rect 1266 1247 1267 1251
rect 1271 1250 1272 1251
rect 1315 1251 1321 1252
rect 1315 1250 1316 1251
rect 1271 1248 1316 1250
rect 1271 1247 1272 1248
rect 1266 1246 1272 1247
rect 1315 1247 1316 1248
rect 1320 1247 1321 1251
rect 1315 1246 1321 1247
rect 1390 1251 1401 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1400 1247 1401 1251
rect 1390 1246 1401 1247
rect 1470 1251 1481 1252
rect 1470 1247 1471 1251
rect 1475 1247 1476 1251
rect 1480 1247 1481 1251
rect 1470 1246 1481 1247
rect 1555 1251 1561 1252
rect 1555 1247 1556 1251
rect 1560 1247 1561 1251
rect 1555 1246 1561 1247
rect 1630 1251 1641 1252
rect 1630 1247 1631 1251
rect 1635 1247 1636 1251
rect 1640 1247 1641 1251
rect 1630 1246 1641 1247
rect 1710 1251 1721 1252
rect 1710 1247 1711 1251
rect 1715 1247 1716 1251
rect 1720 1247 1721 1251
rect 1710 1246 1721 1247
rect 1795 1251 1801 1252
rect 1795 1247 1796 1251
rect 1800 1250 1801 1251
rect 1834 1251 1840 1252
rect 1834 1250 1835 1251
rect 1800 1248 1835 1250
rect 1800 1247 1801 1248
rect 1795 1246 1801 1247
rect 1834 1247 1835 1248
rect 1839 1247 1840 1251
rect 1834 1246 1840 1247
rect 1875 1251 1881 1252
rect 1875 1247 1876 1251
rect 1880 1250 1881 1251
rect 1911 1251 1917 1252
rect 1911 1250 1912 1251
rect 1880 1248 1912 1250
rect 1880 1247 1881 1248
rect 1875 1246 1881 1247
rect 1911 1247 1912 1248
rect 1916 1247 1917 1251
rect 1911 1246 1917 1247
rect 1958 1251 1969 1252
rect 1958 1247 1959 1251
rect 1963 1247 1964 1251
rect 1968 1247 1969 1251
rect 1958 1246 1969 1247
rect 2034 1251 2040 1252
rect 2034 1247 2035 1251
rect 2039 1250 2040 1251
rect 2051 1251 2057 1252
rect 2051 1250 2052 1251
rect 2039 1248 2052 1250
rect 2039 1247 2040 1248
rect 2034 1246 2040 1247
rect 2051 1247 2052 1248
rect 2056 1247 2057 1251
rect 2051 1246 2057 1247
rect 918 1242 929 1243
rect 1302 1243 1308 1244
rect 1302 1242 1303 1243
rect 337 1240 359 1242
rect 1156 1240 1303 1242
rect 262 1236 268 1237
rect 262 1232 263 1236
rect 267 1232 268 1236
rect 262 1231 268 1232
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 110 1228 116 1229
rect 110 1224 111 1228
rect 115 1224 116 1228
rect 337 1226 339 1240
rect 1156 1238 1158 1240
rect 1302 1239 1303 1240
rect 1307 1239 1308 1243
rect 1446 1243 1452 1244
rect 1446 1242 1447 1243
rect 1302 1238 1308 1239
rect 1325 1240 1447 1242
rect 1325 1238 1327 1240
rect 1446 1239 1447 1240
rect 1451 1239 1452 1243
rect 1546 1243 1552 1244
rect 1546 1242 1547 1243
rect 1446 1238 1452 1239
rect 1469 1240 1547 1242
rect 1469 1238 1471 1240
rect 1546 1239 1547 1240
rect 1551 1239 1552 1243
rect 1557 1242 1559 1246
rect 1822 1243 1828 1244
rect 1822 1242 1823 1243
rect 1557 1240 1823 1242
rect 1546 1238 1552 1239
rect 1822 1239 1823 1240
rect 1827 1239 1828 1243
rect 1822 1238 1828 1239
rect 1155 1237 1161 1238
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 414 1236 420 1237
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 542 1236 548 1237
rect 542 1232 543 1236
rect 547 1232 548 1236
rect 542 1231 548 1232
rect 606 1236 612 1237
rect 606 1232 607 1236
rect 611 1232 612 1236
rect 606 1231 612 1232
rect 670 1236 676 1237
rect 670 1232 671 1236
rect 675 1232 676 1236
rect 670 1231 676 1232
rect 734 1236 740 1237
rect 734 1232 735 1236
rect 739 1232 740 1236
rect 734 1231 740 1232
rect 798 1236 804 1237
rect 798 1232 799 1236
rect 803 1232 804 1236
rect 798 1231 804 1232
rect 862 1236 868 1237
rect 862 1232 863 1236
rect 867 1232 868 1236
rect 862 1231 868 1232
rect 926 1236 932 1237
rect 926 1232 927 1236
rect 931 1232 932 1236
rect 1155 1233 1156 1237
rect 1160 1233 1161 1237
rect 1323 1237 1329 1238
rect 1155 1232 1161 1233
rect 1186 1235 1192 1236
rect 926 1231 932 1232
rect 1186 1231 1187 1235
rect 1191 1234 1192 1235
rect 1195 1235 1201 1236
rect 1195 1234 1196 1235
rect 1191 1232 1196 1234
rect 1191 1231 1192 1232
rect 1186 1230 1192 1231
rect 1195 1231 1196 1232
rect 1200 1231 1201 1235
rect 1195 1230 1201 1231
rect 1226 1235 1232 1236
rect 1226 1231 1227 1235
rect 1231 1234 1232 1235
rect 1235 1235 1241 1236
rect 1235 1234 1236 1235
rect 1231 1232 1236 1234
rect 1231 1231 1232 1232
rect 1226 1230 1232 1231
rect 1235 1231 1236 1232
rect 1240 1231 1241 1235
rect 1235 1230 1241 1231
rect 1275 1235 1281 1236
rect 1275 1231 1276 1235
rect 1280 1234 1281 1235
rect 1311 1235 1317 1236
rect 1311 1234 1312 1235
rect 1280 1232 1312 1234
rect 1280 1231 1281 1232
rect 1275 1230 1281 1231
rect 1311 1231 1312 1232
rect 1316 1231 1317 1235
rect 1323 1233 1324 1237
rect 1328 1233 1329 1237
rect 1467 1237 1473 1238
rect 1323 1232 1329 1233
rect 1371 1235 1377 1236
rect 1311 1230 1317 1231
rect 1371 1231 1372 1235
rect 1376 1234 1377 1235
rect 1390 1235 1396 1236
rect 1390 1234 1391 1235
rect 1376 1232 1391 1234
rect 1376 1231 1377 1232
rect 1371 1230 1377 1231
rect 1390 1231 1391 1232
rect 1395 1231 1396 1235
rect 1390 1230 1396 1231
rect 1407 1235 1413 1236
rect 1407 1231 1408 1235
rect 1412 1234 1413 1235
rect 1419 1235 1425 1236
rect 1419 1234 1420 1235
rect 1412 1232 1420 1234
rect 1412 1231 1413 1232
rect 1407 1230 1413 1231
rect 1419 1231 1420 1232
rect 1424 1231 1425 1235
rect 1467 1233 1468 1237
rect 1472 1233 1473 1237
rect 1467 1232 1473 1233
rect 1498 1235 1504 1236
rect 1419 1230 1425 1231
rect 1498 1231 1499 1235
rect 1503 1234 1504 1235
rect 1531 1235 1537 1236
rect 1531 1234 1532 1235
rect 1503 1232 1532 1234
rect 1503 1231 1504 1232
rect 1498 1230 1504 1231
rect 1531 1231 1532 1232
rect 1536 1231 1537 1235
rect 1531 1230 1537 1231
rect 1570 1235 1576 1236
rect 1570 1231 1571 1235
rect 1575 1234 1576 1235
rect 1611 1235 1617 1236
rect 1611 1234 1612 1235
rect 1575 1232 1612 1234
rect 1575 1231 1576 1232
rect 1570 1230 1576 1231
rect 1611 1231 1612 1232
rect 1616 1231 1617 1235
rect 1611 1230 1617 1231
rect 1647 1235 1653 1236
rect 1647 1231 1648 1235
rect 1652 1234 1653 1235
rect 1715 1235 1721 1236
rect 1715 1234 1716 1235
rect 1652 1232 1716 1234
rect 1652 1231 1653 1232
rect 1647 1230 1653 1231
rect 1715 1231 1716 1232
rect 1720 1231 1721 1235
rect 1715 1230 1721 1231
rect 1814 1235 1820 1236
rect 1814 1231 1815 1235
rect 1819 1234 1820 1235
rect 1835 1235 1841 1236
rect 1835 1234 1836 1235
rect 1819 1232 1836 1234
rect 1819 1231 1820 1232
rect 1814 1230 1820 1231
rect 1835 1231 1836 1232
rect 1840 1231 1841 1235
rect 1835 1230 1841 1231
rect 1866 1235 1872 1236
rect 1866 1231 1867 1235
rect 1871 1234 1872 1235
rect 1963 1235 1969 1236
rect 1963 1234 1964 1235
rect 1871 1232 1964 1234
rect 1871 1231 1872 1232
rect 1866 1230 1872 1231
rect 1963 1231 1964 1232
rect 1968 1231 1969 1235
rect 1963 1230 1969 1231
rect 2067 1235 2073 1236
rect 2067 1231 2068 1235
rect 2072 1234 2073 1235
rect 2082 1235 2088 1236
rect 2082 1234 2083 1235
rect 2072 1232 2083 1234
rect 2072 1231 2073 1232
rect 2067 1230 2073 1231
rect 2082 1231 2083 1232
rect 2087 1231 2088 1235
rect 2082 1230 2088 1231
rect 1094 1228 1100 1229
rect 335 1225 341 1226
rect 110 1223 116 1224
rect 287 1223 296 1224
rect 287 1219 288 1223
rect 295 1219 296 1223
rect 335 1221 336 1225
rect 340 1221 341 1225
rect 1094 1224 1095 1228
rect 1099 1224 1100 1228
rect 335 1220 341 1221
rect 383 1223 389 1224
rect 287 1218 296 1219
rect 383 1219 384 1223
rect 388 1222 389 1223
rect 391 1223 397 1224
rect 391 1222 392 1223
rect 388 1220 392 1222
rect 388 1219 389 1220
rect 383 1218 389 1219
rect 391 1219 392 1220
rect 396 1219 397 1223
rect 391 1218 397 1219
rect 439 1223 448 1224
rect 439 1219 440 1223
rect 447 1219 448 1223
rect 439 1218 448 1219
rect 503 1223 509 1224
rect 503 1219 504 1223
rect 508 1222 509 1223
rect 518 1223 524 1224
rect 518 1222 519 1223
rect 508 1220 519 1222
rect 508 1219 509 1220
rect 503 1218 509 1219
rect 518 1219 519 1220
rect 523 1219 524 1223
rect 518 1218 524 1219
rect 566 1223 573 1224
rect 566 1219 567 1223
rect 572 1219 573 1223
rect 566 1218 573 1219
rect 578 1223 584 1224
rect 578 1219 579 1223
rect 583 1222 584 1223
rect 631 1223 637 1224
rect 631 1222 632 1223
rect 583 1220 632 1222
rect 583 1219 584 1220
rect 578 1218 584 1219
rect 631 1219 632 1220
rect 636 1219 637 1223
rect 631 1218 637 1219
rect 639 1223 645 1224
rect 639 1219 640 1223
rect 644 1222 645 1223
rect 695 1223 701 1224
rect 695 1222 696 1223
rect 644 1220 696 1222
rect 644 1219 645 1220
rect 639 1218 645 1219
rect 695 1219 696 1220
rect 700 1219 701 1223
rect 695 1218 701 1219
rect 722 1223 728 1224
rect 722 1219 723 1223
rect 727 1222 728 1223
rect 759 1223 765 1224
rect 759 1222 760 1223
rect 727 1220 760 1222
rect 727 1219 728 1220
rect 722 1218 728 1219
rect 759 1219 760 1220
rect 764 1219 765 1223
rect 759 1218 765 1219
rect 782 1223 788 1224
rect 782 1219 783 1223
rect 787 1222 788 1223
rect 823 1223 829 1224
rect 823 1222 824 1223
rect 787 1220 824 1222
rect 787 1219 788 1220
rect 782 1218 788 1219
rect 823 1219 824 1220
rect 828 1219 829 1223
rect 823 1218 829 1219
rect 886 1223 893 1224
rect 886 1219 887 1223
rect 892 1219 893 1223
rect 886 1218 893 1219
rect 910 1223 916 1224
rect 910 1219 911 1223
rect 915 1222 916 1223
rect 951 1223 957 1224
rect 1094 1223 1100 1224
rect 1158 1224 1164 1225
rect 951 1222 952 1223
rect 915 1220 952 1222
rect 915 1219 916 1220
rect 910 1218 916 1219
rect 951 1219 952 1220
rect 956 1219 957 1223
rect 1158 1220 1159 1224
rect 1163 1220 1164 1224
rect 1158 1219 1164 1220
rect 1198 1224 1204 1225
rect 1198 1220 1199 1224
rect 1203 1220 1204 1224
rect 1198 1219 1204 1220
rect 1238 1224 1244 1225
rect 1238 1220 1239 1224
rect 1243 1220 1244 1224
rect 1238 1219 1244 1220
rect 1278 1224 1284 1225
rect 1278 1220 1279 1224
rect 1283 1220 1284 1224
rect 1278 1219 1284 1220
rect 1326 1224 1332 1225
rect 1326 1220 1327 1224
rect 1331 1220 1332 1224
rect 1326 1219 1332 1220
rect 1374 1224 1380 1225
rect 1374 1220 1375 1224
rect 1379 1220 1380 1224
rect 1374 1219 1380 1220
rect 1422 1224 1428 1225
rect 1422 1220 1423 1224
rect 1427 1220 1428 1224
rect 1422 1219 1428 1220
rect 1470 1224 1476 1225
rect 1470 1220 1471 1224
rect 1475 1220 1476 1224
rect 1470 1219 1476 1220
rect 1534 1224 1540 1225
rect 1534 1220 1535 1224
rect 1539 1220 1540 1224
rect 1534 1219 1540 1220
rect 1614 1224 1620 1225
rect 1614 1220 1615 1224
rect 1619 1220 1620 1224
rect 1614 1219 1620 1220
rect 1718 1224 1724 1225
rect 1718 1220 1719 1224
rect 1723 1220 1724 1224
rect 1718 1219 1724 1220
rect 1838 1224 1844 1225
rect 1838 1220 1839 1224
rect 1843 1220 1844 1224
rect 1838 1219 1844 1220
rect 1966 1224 1972 1225
rect 1966 1220 1967 1224
rect 1971 1220 1972 1224
rect 1966 1219 1972 1220
rect 2070 1224 2076 1225
rect 2070 1220 2071 1224
rect 2075 1220 2076 1224
rect 2070 1219 2076 1220
rect 951 1218 957 1219
rect 1134 1216 1140 1217
rect 2118 1216 2124 1217
rect 1134 1212 1135 1216
rect 1139 1212 1140 1216
rect 1407 1215 1413 1216
rect 110 1211 116 1212
rect 110 1207 111 1211
rect 115 1207 116 1211
rect 1094 1211 1100 1212
rect 1134 1211 1140 1212
rect 1183 1211 1192 1212
rect 110 1206 116 1207
rect 262 1208 268 1209
rect 262 1204 263 1208
rect 267 1204 268 1208
rect 262 1203 268 1204
rect 310 1208 316 1209
rect 310 1204 311 1208
rect 315 1204 316 1208
rect 310 1203 316 1204
rect 358 1208 364 1209
rect 358 1204 359 1208
rect 363 1204 364 1208
rect 358 1203 364 1204
rect 414 1208 420 1209
rect 414 1204 415 1208
rect 419 1204 420 1208
rect 414 1203 420 1204
rect 478 1208 484 1209
rect 478 1204 479 1208
rect 483 1204 484 1208
rect 478 1203 484 1204
rect 542 1208 548 1209
rect 542 1204 543 1208
rect 547 1204 548 1208
rect 542 1203 548 1204
rect 606 1208 612 1209
rect 606 1204 607 1208
rect 611 1204 612 1208
rect 606 1203 612 1204
rect 670 1208 676 1209
rect 670 1204 671 1208
rect 675 1204 676 1208
rect 670 1203 676 1204
rect 734 1208 740 1209
rect 734 1204 735 1208
rect 739 1204 740 1208
rect 734 1203 740 1204
rect 798 1208 804 1209
rect 798 1204 799 1208
rect 803 1204 804 1208
rect 798 1203 804 1204
rect 862 1208 868 1209
rect 862 1204 863 1208
rect 867 1204 868 1208
rect 862 1203 868 1204
rect 926 1208 932 1209
rect 926 1204 927 1208
rect 931 1204 932 1208
rect 1094 1207 1095 1211
rect 1099 1207 1100 1211
rect 1094 1206 1100 1207
rect 1183 1207 1184 1211
rect 1191 1207 1192 1211
rect 1183 1206 1192 1207
rect 1223 1211 1232 1212
rect 1223 1207 1224 1211
rect 1231 1207 1232 1211
rect 1223 1206 1232 1207
rect 1263 1211 1272 1212
rect 1263 1207 1264 1211
rect 1271 1207 1272 1211
rect 1263 1206 1272 1207
rect 1302 1211 1309 1212
rect 1302 1207 1303 1211
rect 1308 1207 1309 1211
rect 1302 1206 1309 1207
rect 1311 1211 1317 1212
rect 1311 1207 1312 1211
rect 1316 1210 1317 1211
rect 1351 1211 1357 1212
rect 1351 1210 1352 1211
rect 1316 1208 1352 1210
rect 1316 1207 1317 1208
rect 1311 1206 1317 1207
rect 1351 1207 1352 1208
rect 1356 1207 1357 1211
rect 1351 1206 1357 1207
rect 1399 1211 1405 1212
rect 1399 1207 1400 1211
rect 1404 1210 1405 1211
rect 1407 1211 1408 1215
rect 1412 1211 1413 1215
rect 1647 1215 1653 1216
rect 1407 1210 1413 1211
rect 1446 1211 1453 1212
rect 1404 1208 1411 1210
rect 1404 1207 1405 1208
rect 1399 1206 1405 1207
rect 1446 1207 1447 1211
rect 1452 1207 1453 1211
rect 1446 1206 1453 1207
rect 1495 1211 1504 1212
rect 1495 1207 1496 1211
rect 1503 1207 1504 1211
rect 1495 1206 1504 1207
rect 1559 1211 1565 1212
rect 1559 1207 1560 1211
rect 1564 1210 1565 1211
rect 1570 1211 1576 1212
rect 1570 1210 1571 1211
rect 1564 1208 1571 1210
rect 1564 1207 1565 1208
rect 1559 1206 1565 1207
rect 1570 1207 1571 1208
rect 1575 1207 1576 1211
rect 1570 1206 1576 1207
rect 1639 1211 1645 1212
rect 1639 1207 1640 1211
rect 1644 1210 1645 1211
rect 1647 1211 1648 1215
rect 1652 1211 1653 1215
rect 2118 1212 2119 1216
rect 2123 1212 2124 1216
rect 1647 1210 1653 1211
rect 1663 1211 1669 1212
rect 1644 1208 1651 1210
rect 1644 1207 1645 1208
rect 1639 1206 1645 1207
rect 1663 1207 1664 1211
rect 1668 1210 1669 1211
rect 1743 1211 1749 1212
rect 1743 1210 1744 1211
rect 1668 1208 1744 1210
rect 1668 1207 1669 1208
rect 1663 1206 1669 1207
rect 1743 1207 1744 1208
rect 1748 1207 1749 1211
rect 1743 1206 1749 1207
rect 1863 1211 1872 1212
rect 1863 1207 1864 1211
rect 1871 1207 1872 1211
rect 1863 1206 1872 1207
rect 1990 1211 1997 1212
rect 1990 1207 1991 1211
rect 1996 1207 1997 1211
rect 1990 1206 1997 1207
rect 2086 1211 2092 1212
rect 2086 1207 2087 1211
rect 2091 1210 2092 1211
rect 2095 1211 2101 1212
rect 2118 1211 2124 1212
rect 2095 1210 2096 1211
rect 2091 1208 2096 1210
rect 2091 1207 2092 1208
rect 2086 1206 2092 1207
rect 2095 1207 2096 1208
rect 2100 1207 2101 1211
rect 2095 1206 2101 1207
rect 926 1203 932 1204
rect 1134 1199 1140 1200
rect 222 1196 228 1197
rect 110 1193 116 1194
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 222 1192 223 1196
rect 227 1192 228 1196
rect 222 1191 228 1192
rect 278 1196 284 1197
rect 278 1192 279 1196
rect 283 1192 284 1196
rect 278 1191 284 1192
rect 342 1196 348 1197
rect 342 1192 343 1196
rect 347 1192 348 1196
rect 342 1191 348 1192
rect 406 1196 412 1197
rect 406 1192 407 1196
rect 411 1192 412 1196
rect 406 1191 412 1192
rect 478 1196 484 1197
rect 478 1192 479 1196
rect 483 1192 484 1196
rect 478 1191 484 1192
rect 550 1196 556 1197
rect 550 1192 551 1196
rect 555 1192 556 1196
rect 550 1191 556 1192
rect 630 1196 636 1197
rect 630 1192 631 1196
rect 635 1192 636 1196
rect 630 1191 636 1192
rect 710 1196 716 1197
rect 710 1192 711 1196
rect 715 1192 716 1196
rect 710 1191 716 1192
rect 790 1196 796 1197
rect 790 1192 791 1196
rect 795 1192 796 1196
rect 790 1191 796 1192
rect 870 1196 876 1197
rect 870 1192 871 1196
rect 875 1192 876 1196
rect 870 1191 876 1192
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 1134 1195 1135 1199
rect 1139 1195 1140 1199
rect 2118 1199 2124 1200
rect 1134 1194 1140 1195
rect 1158 1196 1164 1197
rect 958 1191 964 1192
rect 1094 1193 1100 1194
rect 110 1188 116 1189
rect 1094 1189 1095 1193
rect 1099 1189 1100 1193
rect 1158 1192 1159 1196
rect 1163 1192 1164 1196
rect 1158 1191 1164 1192
rect 1198 1196 1204 1197
rect 1198 1192 1199 1196
rect 1203 1192 1204 1196
rect 1198 1191 1204 1192
rect 1238 1196 1244 1197
rect 1238 1192 1239 1196
rect 1243 1192 1244 1196
rect 1238 1191 1244 1192
rect 1278 1196 1284 1197
rect 1278 1192 1279 1196
rect 1283 1192 1284 1196
rect 1278 1191 1284 1192
rect 1326 1196 1332 1197
rect 1326 1192 1327 1196
rect 1331 1192 1332 1196
rect 1326 1191 1332 1192
rect 1374 1196 1380 1197
rect 1374 1192 1375 1196
rect 1379 1192 1380 1196
rect 1374 1191 1380 1192
rect 1422 1196 1428 1197
rect 1422 1192 1423 1196
rect 1427 1192 1428 1196
rect 1422 1191 1428 1192
rect 1470 1196 1476 1197
rect 1470 1192 1471 1196
rect 1475 1192 1476 1196
rect 1470 1191 1476 1192
rect 1534 1196 1540 1197
rect 1534 1192 1535 1196
rect 1539 1192 1540 1196
rect 1534 1191 1540 1192
rect 1614 1196 1620 1197
rect 1614 1192 1615 1196
rect 1619 1192 1620 1196
rect 1718 1196 1724 1197
rect 1718 1192 1719 1196
rect 1723 1192 1724 1196
rect 1614 1191 1620 1192
rect 1622 1191 1628 1192
rect 1094 1188 1100 1189
rect 270 1187 276 1188
rect 270 1183 271 1187
rect 275 1186 276 1187
rect 1622 1187 1623 1191
rect 1627 1190 1628 1191
rect 1663 1191 1669 1192
rect 1718 1191 1724 1192
rect 1838 1196 1844 1197
rect 1838 1192 1839 1196
rect 1843 1192 1844 1196
rect 1838 1191 1844 1192
rect 1966 1196 1972 1197
rect 1966 1192 1967 1196
rect 1971 1192 1972 1196
rect 1966 1191 1972 1192
rect 2070 1196 2076 1197
rect 2070 1192 2071 1196
rect 2075 1192 2076 1196
rect 2118 1195 2119 1199
rect 2123 1195 2124 1199
rect 2118 1194 2124 1195
rect 2070 1191 2076 1192
rect 1663 1190 1664 1191
rect 1627 1188 1664 1190
rect 1627 1187 1628 1188
rect 1622 1186 1628 1187
rect 1663 1187 1664 1188
rect 1668 1187 1669 1191
rect 1663 1186 1669 1187
rect 275 1184 482 1186
rect 275 1183 276 1184
rect 270 1182 276 1183
rect 247 1179 253 1180
rect 110 1176 116 1177
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 247 1175 248 1179
rect 252 1178 253 1179
rect 270 1179 276 1180
rect 270 1178 271 1179
rect 252 1176 271 1178
rect 252 1175 253 1176
rect 247 1174 253 1175
rect 270 1175 271 1176
rect 275 1175 276 1179
rect 270 1174 276 1175
rect 303 1179 309 1180
rect 303 1175 304 1179
rect 308 1178 309 1179
rect 334 1179 340 1180
rect 334 1178 335 1179
rect 308 1176 335 1178
rect 308 1175 309 1176
rect 303 1174 309 1175
rect 334 1175 335 1176
rect 339 1175 340 1179
rect 334 1174 340 1175
rect 367 1179 373 1180
rect 367 1175 368 1179
rect 372 1178 373 1179
rect 398 1179 404 1180
rect 398 1178 399 1179
rect 372 1176 399 1178
rect 372 1175 373 1176
rect 367 1174 373 1175
rect 398 1175 399 1176
rect 403 1175 404 1179
rect 398 1174 404 1175
rect 431 1179 437 1180
rect 431 1175 432 1179
rect 436 1178 437 1179
rect 470 1179 476 1180
rect 470 1178 471 1179
rect 436 1176 471 1178
rect 436 1175 437 1176
rect 431 1174 437 1175
rect 470 1175 471 1176
rect 475 1175 476 1179
rect 480 1178 482 1184
rect 1286 1184 1292 1185
rect 1134 1181 1140 1182
rect 503 1179 509 1180
rect 503 1178 504 1179
rect 480 1176 504 1178
rect 470 1174 476 1175
rect 503 1175 504 1176
rect 508 1175 509 1179
rect 503 1174 509 1175
rect 575 1179 581 1180
rect 575 1175 576 1179
rect 580 1178 581 1179
rect 622 1179 628 1180
rect 622 1178 623 1179
rect 580 1176 623 1178
rect 580 1175 581 1176
rect 575 1174 581 1175
rect 622 1175 623 1176
rect 627 1175 628 1179
rect 622 1174 628 1175
rect 655 1179 661 1180
rect 655 1175 656 1179
rect 660 1178 661 1179
rect 702 1179 708 1180
rect 702 1178 703 1179
rect 660 1176 703 1178
rect 660 1175 661 1176
rect 655 1174 661 1175
rect 702 1175 703 1176
rect 707 1175 708 1179
rect 702 1174 708 1175
rect 735 1179 741 1180
rect 735 1175 736 1179
rect 740 1178 741 1179
rect 782 1179 788 1180
rect 782 1178 783 1179
rect 740 1176 783 1178
rect 740 1175 741 1176
rect 735 1174 741 1175
rect 782 1175 783 1176
rect 787 1175 788 1179
rect 782 1174 788 1175
rect 798 1179 804 1180
rect 798 1175 799 1179
rect 803 1178 804 1179
rect 815 1179 821 1180
rect 815 1178 816 1179
rect 803 1176 816 1178
rect 803 1175 804 1176
rect 798 1174 804 1175
rect 815 1175 816 1176
rect 820 1175 821 1179
rect 815 1174 821 1175
rect 895 1179 901 1180
rect 895 1175 896 1179
rect 900 1178 901 1179
rect 950 1179 956 1180
rect 950 1178 951 1179
rect 900 1176 951 1178
rect 900 1175 901 1176
rect 895 1174 901 1175
rect 950 1175 951 1176
rect 955 1175 956 1179
rect 950 1174 956 1175
rect 982 1179 989 1180
rect 982 1175 983 1179
rect 988 1175 989 1179
rect 1134 1177 1135 1181
rect 1139 1177 1140 1181
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 1326 1184 1332 1185
rect 1326 1180 1327 1184
rect 1331 1180 1332 1184
rect 1326 1179 1332 1180
rect 1366 1184 1372 1185
rect 1366 1180 1367 1184
rect 1371 1180 1372 1184
rect 1366 1179 1372 1180
rect 1414 1184 1420 1185
rect 1414 1180 1415 1184
rect 1419 1180 1420 1184
rect 1414 1179 1420 1180
rect 1470 1184 1476 1185
rect 1470 1180 1471 1184
rect 1475 1180 1476 1184
rect 1470 1179 1476 1180
rect 1526 1184 1532 1185
rect 1526 1180 1527 1184
rect 1531 1180 1532 1184
rect 1526 1179 1532 1180
rect 1582 1184 1588 1185
rect 1582 1180 1583 1184
rect 1587 1180 1588 1184
rect 1582 1179 1588 1180
rect 1638 1184 1644 1185
rect 1638 1180 1639 1184
rect 1643 1180 1644 1184
rect 1638 1179 1644 1180
rect 1702 1184 1708 1185
rect 1702 1180 1703 1184
rect 1707 1180 1708 1184
rect 1702 1179 1708 1180
rect 1766 1184 1772 1185
rect 1766 1180 1767 1184
rect 1771 1180 1772 1184
rect 1766 1179 1772 1180
rect 1838 1184 1844 1185
rect 1838 1180 1839 1184
rect 1843 1180 1844 1184
rect 1838 1179 1844 1180
rect 1918 1184 1924 1185
rect 1918 1180 1919 1184
rect 1923 1180 1924 1184
rect 1918 1179 1924 1180
rect 2006 1184 2012 1185
rect 2006 1180 2007 1184
rect 2011 1180 2012 1184
rect 2006 1179 2012 1180
rect 2070 1184 2076 1185
rect 2070 1180 2071 1184
rect 2075 1180 2076 1184
rect 2070 1179 2076 1180
rect 2118 1181 2124 1182
rect 982 1174 989 1175
rect 1094 1176 1100 1177
rect 1134 1176 1140 1177
rect 2118 1177 2119 1181
rect 2123 1177 2124 1181
rect 2118 1176 2124 1177
rect 110 1171 116 1172
rect 1094 1172 1095 1176
rect 1099 1172 1100 1176
rect 1094 1171 1100 1172
rect 1438 1175 1444 1176
rect 1438 1171 1439 1175
rect 1443 1174 1444 1175
rect 1554 1175 1560 1176
rect 1443 1172 1530 1174
rect 1443 1171 1444 1172
rect 1438 1170 1444 1171
rect 222 1168 228 1169
rect 222 1164 223 1168
rect 227 1164 228 1168
rect 222 1163 228 1164
rect 278 1168 284 1169
rect 278 1164 279 1168
rect 283 1164 284 1168
rect 278 1163 284 1164
rect 342 1168 348 1169
rect 342 1164 343 1168
rect 347 1164 348 1168
rect 342 1163 348 1164
rect 406 1168 412 1169
rect 406 1164 407 1168
rect 411 1164 412 1168
rect 406 1163 412 1164
rect 478 1168 484 1169
rect 478 1164 479 1168
rect 483 1164 484 1168
rect 478 1163 484 1164
rect 550 1168 556 1169
rect 550 1164 551 1168
rect 555 1164 556 1168
rect 550 1163 556 1164
rect 630 1168 636 1169
rect 630 1164 631 1168
rect 635 1164 636 1168
rect 630 1163 636 1164
rect 710 1168 716 1169
rect 710 1164 711 1168
rect 715 1164 716 1168
rect 710 1163 716 1164
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 870 1168 876 1169
rect 870 1164 871 1168
rect 875 1164 876 1168
rect 870 1163 876 1164
rect 958 1168 964 1169
rect 958 1164 959 1168
rect 963 1164 964 1168
rect 1311 1167 1320 1168
rect 958 1163 964 1164
rect 1134 1164 1140 1165
rect 1134 1160 1135 1164
rect 1139 1160 1140 1164
rect 1311 1163 1312 1167
rect 1319 1163 1320 1167
rect 1311 1162 1320 1163
rect 1351 1167 1360 1168
rect 1351 1163 1352 1167
rect 1359 1163 1360 1167
rect 1351 1162 1360 1163
rect 1390 1167 1397 1168
rect 1390 1163 1391 1167
rect 1396 1163 1397 1167
rect 1390 1162 1397 1163
rect 1399 1167 1405 1168
rect 1399 1163 1400 1167
rect 1404 1166 1405 1167
rect 1439 1167 1445 1168
rect 1439 1166 1440 1167
rect 1404 1164 1440 1166
rect 1404 1163 1405 1164
rect 1399 1162 1405 1163
rect 1439 1163 1440 1164
rect 1444 1163 1445 1167
rect 1439 1162 1445 1163
rect 1495 1167 1501 1168
rect 1495 1163 1496 1167
rect 1500 1166 1501 1167
rect 1518 1167 1524 1168
rect 1518 1166 1519 1167
rect 1500 1164 1519 1166
rect 1500 1163 1501 1164
rect 1495 1162 1501 1163
rect 1518 1163 1519 1164
rect 1523 1163 1524 1167
rect 1528 1166 1530 1172
rect 1554 1171 1555 1175
rect 1559 1174 1560 1175
rect 1990 1175 1996 1176
rect 1990 1174 1991 1175
rect 1559 1172 1991 1174
rect 1559 1171 1560 1172
rect 1554 1170 1560 1171
rect 1990 1171 1991 1172
rect 1995 1171 1996 1175
rect 1990 1170 1996 1171
rect 1551 1167 1557 1168
rect 1551 1166 1552 1167
rect 1528 1164 1552 1166
rect 1518 1162 1524 1163
rect 1551 1163 1552 1164
rect 1556 1163 1557 1167
rect 1551 1162 1557 1163
rect 1607 1167 1613 1168
rect 1607 1163 1608 1167
rect 1612 1166 1613 1167
rect 1630 1167 1636 1168
rect 1630 1166 1631 1167
rect 1612 1164 1631 1166
rect 1612 1163 1613 1164
rect 1607 1162 1613 1163
rect 1630 1163 1631 1164
rect 1635 1163 1636 1167
rect 1630 1162 1636 1163
rect 1663 1167 1669 1168
rect 1663 1163 1664 1167
rect 1668 1166 1669 1167
rect 1694 1167 1700 1168
rect 1694 1166 1695 1167
rect 1668 1164 1695 1166
rect 1668 1163 1669 1164
rect 1663 1162 1669 1163
rect 1694 1163 1695 1164
rect 1699 1163 1700 1167
rect 1694 1162 1700 1163
rect 1727 1167 1733 1168
rect 1727 1163 1728 1167
rect 1732 1166 1733 1167
rect 1758 1167 1764 1168
rect 1758 1166 1759 1167
rect 1732 1164 1759 1166
rect 1732 1163 1733 1164
rect 1727 1162 1733 1163
rect 1758 1163 1759 1164
rect 1763 1163 1764 1167
rect 1758 1162 1764 1163
rect 1791 1167 1797 1168
rect 1791 1163 1792 1167
rect 1796 1166 1797 1167
rect 1830 1167 1836 1168
rect 1830 1166 1831 1167
rect 1796 1164 1831 1166
rect 1796 1163 1797 1164
rect 1791 1162 1797 1163
rect 1830 1163 1831 1164
rect 1835 1163 1836 1167
rect 1830 1162 1836 1163
rect 1863 1167 1869 1168
rect 1863 1163 1864 1167
rect 1868 1166 1869 1167
rect 1910 1167 1916 1168
rect 1910 1166 1911 1167
rect 1868 1164 1911 1166
rect 1868 1163 1869 1164
rect 1863 1162 1869 1163
rect 1910 1163 1911 1164
rect 1915 1163 1916 1167
rect 1910 1162 1916 1163
rect 1934 1167 1940 1168
rect 1934 1163 1935 1167
rect 1939 1166 1940 1167
rect 1943 1167 1949 1168
rect 1943 1166 1944 1167
rect 1939 1164 1944 1166
rect 1939 1163 1940 1164
rect 1934 1162 1940 1163
rect 1943 1163 1944 1164
rect 1948 1163 1949 1167
rect 1943 1162 1949 1163
rect 2031 1167 2040 1168
rect 2031 1163 2032 1167
rect 2039 1163 2040 1167
rect 2031 1162 2040 1163
rect 2078 1167 2084 1168
rect 2078 1163 2079 1167
rect 2083 1166 2084 1167
rect 2095 1167 2101 1168
rect 2095 1166 2096 1167
rect 2083 1164 2096 1166
rect 2083 1163 2084 1164
rect 2078 1162 2084 1163
rect 2095 1163 2096 1164
rect 2100 1163 2101 1167
rect 2095 1162 2101 1163
rect 2118 1164 2124 1165
rect 1134 1159 1140 1160
rect 2118 1160 2119 1164
rect 2123 1160 2124 1164
rect 2118 1159 2124 1160
rect 1286 1156 1292 1157
rect 219 1155 225 1156
rect 219 1151 220 1155
rect 224 1154 225 1155
rect 262 1155 268 1156
rect 262 1154 263 1155
rect 224 1152 263 1154
rect 224 1151 225 1152
rect 219 1150 225 1151
rect 262 1151 263 1152
rect 267 1151 268 1155
rect 262 1150 268 1151
rect 270 1155 281 1156
rect 270 1151 271 1155
rect 275 1151 276 1155
rect 280 1151 281 1155
rect 270 1150 281 1151
rect 334 1155 345 1156
rect 334 1151 335 1155
rect 339 1151 340 1155
rect 344 1151 345 1155
rect 334 1150 345 1151
rect 398 1155 409 1156
rect 398 1151 399 1155
rect 403 1151 404 1155
rect 408 1151 409 1155
rect 398 1150 409 1151
rect 470 1155 481 1156
rect 470 1151 471 1155
rect 475 1151 476 1155
rect 480 1151 481 1155
rect 470 1150 481 1151
rect 547 1155 553 1156
rect 547 1151 548 1155
rect 552 1154 553 1155
rect 578 1155 584 1156
rect 578 1154 579 1155
rect 552 1152 579 1154
rect 552 1151 553 1152
rect 547 1150 553 1151
rect 578 1151 579 1152
rect 583 1151 584 1155
rect 578 1150 584 1151
rect 622 1155 633 1156
rect 622 1151 623 1155
rect 627 1151 628 1155
rect 632 1151 633 1155
rect 622 1150 633 1151
rect 702 1155 713 1156
rect 702 1151 703 1155
rect 707 1151 708 1155
rect 712 1151 713 1155
rect 702 1150 713 1151
rect 782 1155 793 1156
rect 782 1151 783 1155
rect 787 1151 788 1155
rect 792 1151 793 1155
rect 782 1150 793 1151
rect 867 1155 873 1156
rect 867 1151 868 1155
rect 872 1154 873 1155
rect 886 1155 892 1156
rect 886 1154 887 1155
rect 872 1152 887 1154
rect 872 1151 873 1152
rect 867 1150 873 1151
rect 886 1151 887 1152
rect 891 1151 892 1155
rect 886 1150 892 1151
rect 950 1155 961 1156
rect 950 1151 951 1155
rect 955 1151 956 1155
rect 960 1151 961 1155
rect 1286 1152 1287 1156
rect 1291 1152 1292 1156
rect 1286 1151 1292 1152
rect 1326 1156 1332 1157
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1366 1156 1372 1157
rect 1366 1152 1367 1156
rect 1371 1152 1372 1156
rect 1366 1151 1372 1152
rect 1414 1156 1420 1157
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1414 1151 1420 1152
rect 1470 1156 1476 1157
rect 1470 1152 1471 1156
rect 1475 1152 1476 1156
rect 1470 1151 1476 1152
rect 1526 1156 1532 1157
rect 1526 1152 1527 1156
rect 1531 1152 1532 1156
rect 1526 1151 1532 1152
rect 1582 1156 1588 1157
rect 1582 1152 1583 1156
rect 1587 1152 1588 1156
rect 1582 1151 1588 1152
rect 1638 1156 1644 1157
rect 1638 1152 1639 1156
rect 1643 1152 1644 1156
rect 1638 1151 1644 1152
rect 1702 1156 1708 1157
rect 1702 1152 1703 1156
rect 1707 1152 1708 1156
rect 1702 1151 1708 1152
rect 1766 1156 1772 1157
rect 1766 1152 1767 1156
rect 1771 1152 1772 1156
rect 1766 1151 1772 1152
rect 1838 1156 1844 1157
rect 1838 1152 1839 1156
rect 1843 1152 1844 1156
rect 1838 1151 1844 1152
rect 1918 1156 1924 1157
rect 1918 1152 1919 1156
rect 1923 1152 1924 1156
rect 1918 1151 1924 1152
rect 2006 1156 2012 1157
rect 2006 1152 2007 1156
rect 2011 1152 2012 1156
rect 2006 1151 2012 1152
rect 2070 1156 2076 1157
rect 2070 1152 2071 1156
rect 2075 1152 2076 1156
rect 2070 1151 2076 1152
rect 950 1150 961 1151
rect 155 1143 161 1144
rect 155 1139 156 1143
rect 160 1142 161 1143
rect 174 1143 180 1144
rect 174 1142 175 1143
rect 160 1140 175 1142
rect 160 1139 161 1140
rect 155 1138 161 1139
rect 174 1139 175 1140
rect 179 1139 180 1143
rect 174 1138 180 1139
rect 182 1143 188 1144
rect 182 1139 183 1143
rect 187 1142 188 1143
rect 195 1143 201 1144
rect 195 1142 196 1143
rect 187 1140 196 1142
rect 187 1139 188 1140
rect 182 1138 188 1139
rect 195 1139 196 1140
rect 200 1139 201 1143
rect 195 1138 201 1139
rect 230 1143 236 1144
rect 230 1139 231 1143
rect 235 1142 236 1143
rect 243 1143 249 1144
rect 243 1142 244 1143
rect 235 1140 244 1142
rect 235 1139 236 1140
rect 230 1138 236 1139
rect 243 1139 244 1140
rect 248 1139 249 1143
rect 243 1138 249 1139
rect 286 1143 292 1144
rect 286 1139 287 1143
rect 291 1142 292 1143
rect 299 1143 305 1144
rect 299 1142 300 1143
rect 291 1140 300 1142
rect 291 1139 292 1140
rect 286 1138 292 1139
rect 299 1139 300 1140
rect 304 1139 305 1143
rect 299 1138 305 1139
rect 343 1143 349 1144
rect 343 1139 344 1143
rect 348 1142 349 1143
rect 363 1143 369 1144
rect 363 1142 364 1143
rect 348 1140 364 1142
rect 348 1139 349 1140
rect 343 1138 349 1139
rect 363 1139 364 1140
rect 368 1139 369 1143
rect 363 1138 369 1139
rect 394 1143 400 1144
rect 394 1139 395 1143
rect 399 1142 400 1143
rect 435 1143 441 1144
rect 435 1142 436 1143
rect 399 1140 436 1142
rect 399 1139 400 1140
rect 394 1138 400 1139
rect 435 1139 436 1140
rect 440 1139 441 1143
rect 435 1138 441 1139
rect 507 1143 513 1144
rect 507 1139 508 1143
rect 512 1142 513 1143
rect 578 1143 584 1144
rect 578 1142 579 1143
rect 512 1140 579 1142
rect 512 1139 513 1140
rect 507 1138 513 1139
rect 578 1139 579 1140
rect 583 1139 584 1143
rect 578 1138 584 1139
rect 587 1143 593 1144
rect 587 1139 588 1143
rect 592 1142 593 1143
rect 666 1143 672 1144
rect 666 1142 667 1143
rect 592 1140 667 1142
rect 592 1139 593 1140
rect 587 1138 593 1139
rect 666 1139 667 1140
rect 671 1139 672 1143
rect 666 1138 672 1139
rect 675 1143 681 1144
rect 675 1139 676 1143
rect 680 1142 681 1143
rect 762 1143 768 1144
rect 762 1142 763 1143
rect 680 1140 763 1142
rect 680 1139 681 1140
rect 675 1138 681 1139
rect 762 1139 763 1140
rect 767 1139 768 1143
rect 762 1138 768 1139
rect 771 1143 777 1144
rect 771 1139 772 1143
rect 776 1142 777 1143
rect 798 1143 804 1144
rect 798 1142 799 1143
rect 776 1140 799 1142
rect 776 1139 777 1140
rect 771 1138 777 1139
rect 798 1139 799 1140
rect 803 1139 804 1143
rect 798 1138 804 1139
rect 875 1143 881 1144
rect 875 1139 876 1143
rect 880 1142 881 1143
rect 974 1143 980 1144
rect 974 1142 975 1143
rect 880 1140 975 1142
rect 880 1139 881 1140
rect 875 1138 881 1139
rect 974 1139 975 1140
rect 979 1139 980 1143
rect 974 1138 980 1139
rect 982 1143 993 1144
rect 982 1139 983 1143
rect 987 1139 988 1143
rect 992 1139 993 1143
rect 982 1138 993 1139
rect 1283 1143 1289 1144
rect 1283 1139 1284 1143
rect 1288 1142 1289 1143
rect 1314 1143 1320 1144
rect 1288 1140 1310 1142
rect 1288 1139 1289 1140
rect 1283 1138 1289 1139
rect 1308 1134 1310 1140
rect 1314 1139 1315 1143
rect 1319 1142 1320 1143
rect 1323 1143 1329 1144
rect 1323 1142 1324 1143
rect 1319 1140 1324 1142
rect 1319 1139 1320 1140
rect 1314 1138 1320 1139
rect 1323 1139 1324 1140
rect 1328 1139 1329 1143
rect 1323 1138 1329 1139
rect 1354 1143 1360 1144
rect 1354 1139 1355 1143
rect 1359 1142 1360 1143
rect 1363 1143 1369 1144
rect 1363 1142 1364 1143
rect 1359 1140 1364 1142
rect 1359 1139 1360 1140
rect 1354 1138 1360 1139
rect 1363 1139 1364 1140
rect 1368 1139 1369 1143
rect 1363 1138 1369 1139
rect 1411 1143 1417 1144
rect 1411 1139 1412 1143
rect 1416 1142 1417 1143
rect 1438 1143 1444 1144
rect 1438 1142 1439 1143
rect 1416 1140 1439 1142
rect 1416 1139 1417 1140
rect 1411 1138 1417 1139
rect 1438 1139 1439 1140
rect 1443 1139 1444 1143
rect 1438 1138 1444 1139
rect 1467 1143 1473 1144
rect 1467 1139 1468 1143
rect 1472 1142 1473 1143
rect 1494 1143 1500 1144
rect 1494 1142 1495 1143
rect 1472 1140 1495 1142
rect 1472 1139 1473 1140
rect 1467 1138 1473 1139
rect 1494 1139 1495 1140
rect 1499 1139 1500 1143
rect 1494 1138 1500 1139
rect 1518 1143 1529 1144
rect 1518 1139 1519 1143
rect 1523 1139 1524 1143
rect 1528 1139 1529 1143
rect 1518 1138 1529 1139
rect 1579 1143 1585 1144
rect 1579 1139 1580 1143
rect 1584 1142 1585 1143
rect 1622 1143 1628 1144
rect 1622 1142 1623 1143
rect 1584 1140 1623 1142
rect 1584 1139 1585 1140
rect 1579 1138 1585 1139
rect 1622 1139 1623 1140
rect 1627 1139 1628 1143
rect 1622 1138 1628 1139
rect 1630 1143 1641 1144
rect 1630 1139 1631 1143
rect 1635 1139 1636 1143
rect 1640 1139 1641 1143
rect 1630 1138 1641 1139
rect 1694 1143 1705 1144
rect 1694 1139 1695 1143
rect 1699 1139 1700 1143
rect 1704 1139 1705 1143
rect 1694 1138 1705 1139
rect 1758 1143 1769 1144
rect 1758 1139 1759 1143
rect 1763 1139 1764 1143
rect 1768 1139 1769 1143
rect 1758 1138 1769 1139
rect 1830 1143 1841 1144
rect 1830 1139 1831 1143
rect 1835 1139 1836 1143
rect 1840 1139 1841 1143
rect 1830 1138 1841 1139
rect 1910 1143 1921 1144
rect 1910 1139 1911 1143
rect 1915 1139 1916 1143
rect 1920 1139 1921 1143
rect 1910 1138 1921 1139
rect 2003 1143 2009 1144
rect 2003 1139 2004 1143
rect 2008 1142 2009 1143
rect 2054 1143 2060 1144
rect 2054 1142 2055 1143
rect 2008 1140 2055 1142
rect 2008 1139 2009 1140
rect 2003 1138 2009 1139
rect 2054 1139 2055 1140
rect 2059 1139 2060 1143
rect 2054 1138 2060 1139
rect 2067 1143 2073 1144
rect 2067 1139 2068 1143
rect 2072 1142 2073 1143
rect 2086 1143 2092 1144
rect 2086 1142 2087 1143
rect 2072 1140 2087 1142
rect 2072 1139 2073 1140
rect 2067 1138 2073 1139
rect 2086 1139 2087 1140
rect 2091 1139 2092 1143
rect 2086 1138 2092 1139
rect 1399 1135 1405 1136
rect 1399 1134 1400 1135
rect 158 1132 164 1133
rect 158 1128 159 1132
rect 163 1128 164 1132
rect 158 1127 164 1128
rect 198 1132 204 1133
rect 198 1128 199 1132
rect 203 1128 204 1132
rect 198 1127 204 1128
rect 246 1132 252 1133
rect 246 1128 247 1132
rect 251 1128 252 1132
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 246 1127 252 1128
rect 262 1127 268 1128
rect 302 1127 308 1128
rect 366 1132 372 1133
rect 366 1128 367 1132
rect 371 1128 372 1132
rect 366 1127 372 1128
rect 438 1132 444 1133
rect 438 1128 439 1132
rect 443 1128 444 1132
rect 438 1127 444 1128
rect 510 1132 516 1133
rect 510 1128 511 1132
rect 515 1128 516 1132
rect 510 1127 516 1128
rect 590 1132 596 1133
rect 590 1128 591 1132
rect 595 1128 596 1132
rect 590 1127 596 1128
rect 678 1132 684 1133
rect 678 1128 679 1132
rect 683 1128 684 1132
rect 678 1127 684 1128
rect 774 1132 780 1133
rect 774 1128 775 1132
rect 779 1128 780 1132
rect 774 1127 780 1128
rect 878 1132 884 1133
rect 878 1128 879 1132
rect 883 1128 884 1132
rect 878 1127 884 1128
rect 990 1132 996 1133
rect 1308 1132 1400 1134
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 1399 1131 1400 1132
rect 1404 1131 1405 1135
rect 1399 1130 1405 1131
rect 1678 1131 1684 1132
rect 1678 1130 1679 1131
rect 990 1127 996 1128
rect 1524 1128 1679 1130
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 262 1123 263 1127
rect 267 1126 268 1127
rect 1524 1126 1526 1128
rect 1678 1127 1679 1128
rect 1683 1127 1684 1131
rect 1934 1131 1940 1132
rect 1934 1130 1935 1131
rect 1678 1126 1684 1127
rect 1708 1128 1935 1130
rect 1708 1126 1710 1128
rect 1934 1127 1935 1128
rect 1939 1127 1940 1131
rect 1934 1126 1940 1127
rect 267 1124 298 1126
rect 267 1123 268 1124
rect 262 1122 268 1123
rect 296 1122 298 1124
rect 319 1124 362 1126
rect 319 1122 321 1124
rect 296 1120 321 1122
rect 360 1122 362 1124
rect 384 1124 406 1126
rect 1523 1125 1529 1126
rect 384 1122 386 1124
rect 360 1120 386 1122
rect 110 1119 116 1120
rect 182 1119 189 1120
rect 182 1115 183 1119
rect 188 1115 189 1119
rect 182 1114 189 1115
rect 223 1119 232 1120
rect 223 1115 224 1119
rect 231 1115 232 1119
rect 223 1114 232 1115
rect 271 1119 277 1120
rect 271 1115 272 1119
rect 276 1118 277 1119
rect 286 1119 292 1120
rect 286 1118 287 1119
rect 276 1116 287 1118
rect 276 1115 277 1116
rect 271 1114 277 1115
rect 286 1115 287 1116
rect 291 1115 292 1119
rect 286 1114 292 1115
rect 327 1119 333 1120
rect 327 1115 328 1119
rect 332 1118 333 1119
rect 343 1119 349 1120
rect 343 1118 344 1119
rect 332 1116 344 1118
rect 332 1115 333 1116
rect 327 1114 333 1115
rect 343 1115 344 1116
rect 348 1115 349 1119
rect 343 1114 349 1115
rect 391 1119 400 1120
rect 391 1115 392 1119
rect 399 1115 400 1119
rect 404 1118 406 1124
rect 1094 1124 1100 1125
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 463 1119 469 1120
rect 463 1118 464 1119
rect 404 1116 464 1118
rect 391 1114 400 1115
rect 463 1115 464 1116
rect 468 1115 469 1119
rect 463 1114 469 1115
rect 518 1119 524 1120
rect 518 1115 519 1119
rect 523 1118 524 1119
rect 535 1119 541 1120
rect 535 1118 536 1119
rect 523 1116 536 1118
rect 523 1115 524 1116
rect 518 1114 524 1115
rect 535 1115 536 1116
rect 540 1115 541 1119
rect 535 1114 541 1115
rect 578 1119 584 1120
rect 578 1115 579 1119
rect 583 1118 584 1119
rect 615 1119 621 1120
rect 615 1118 616 1119
rect 583 1116 616 1118
rect 583 1115 584 1116
rect 578 1114 584 1115
rect 615 1115 616 1116
rect 620 1115 621 1119
rect 615 1114 621 1115
rect 666 1119 672 1120
rect 666 1115 667 1119
rect 671 1118 672 1119
rect 703 1119 709 1120
rect 703 1118 704 1119
rect 671 1116 704 1118
rect 671 1115 672 1116
rect 666 1114 672 1115
rect 703 1115 704 1116
rect 708 1115 709 1119
rect 703 1114 709 1115
rect 762 1119 768 1120
rect 762 1115 763 1119
rect 767 1118 768 1119
rect 799 1119 805 1120
rect 799 1118 800 1119
rect 767 1116 800 1118
rect 767 1115 768 1116
rect 762 1114 768 1115
rect 799 1115 800 1116
rect 804 1115 805 1119
rect 799 1114 805 1115
rect 810 1119 816 1120
rect 810 1115 811 1119
rect 815 1118 816 1119
rect 903 1119 909 1120
rect 903 1118 904 1119
rect 815 1116 904 1118
rect 815 1115 816 1116
rect 810 1114 816 1115
rect 903 1115 904 1116
rect 908 1115 909 1119
rect 903 1114 909 1115
rect 974 1119 980 1120
rect 974 1115 975 1119
rect 979 1118 980 1119
rect 1015 1119 1021 1120
rect 1094 1119 1100 1120
rect 1379 1123 1385 1124
rect 1379 1119 1380 1123
rect 1384 1122 1385 1123
rect 1398 1123 1404 1124
rect 1398 1122 1399 1123
rect 1384 1120 1399 1122
rect 1384 1119 1385 1120
rect 1015 1118 1016 1119
rect 979 1116 1016 1118
rect 979 1115 980 1116
rect 974 1114 980 1115
rect 1015 1115 1016 1116
rect 1020 1115 1021 1119
rect 1379 1118 1385 1119
rect 1398 1119 1399 1120
rect 1403 1119 1404 1123
rect 1398 1118 1404 1119
rect 1406 1123 1412 1124
rect 1406 1119 1407 1123
rect 1411 1122 1412 1123
rect 1419 1123 1425 1124
rect 1419 1122 1420 1123
rect 1411 1120 1420 1122
rect 1411 1119 1412 1120
rect 1406 1118 1412 1119
rect 1419 1119 1420 1120
rect 1424 1119 1425 1123
rect 1419 1118 1425 1119
rect 1450 1123 1456 1124
rect 1450 1119 1451 1123
rect 1455 1122 1456 1123
rect 1467 1123 1473 1124
rect 1467 1122 1468 1123
rect 1455 1120 1468 1122
rect 1455 1119 1456 1120
rect 1450 1118 1456 1119
rect 1467 1119 1468 1120
rect 1472 1119 1473 1123
rect 1523 1121 1524 1125
rect 1528 1121 1529 1125
rect 1707 1125 1713 1126
rect 1523 1120 1529 1121
rect 1587 1123 1593 1124
rect 1467 1118 1473 1119
rect 1587 1119 1588 1123
rect 1592 1122 1593 1123
rect 1598 1123 1604 1124
rect 1598 1122 1599 1123
rect 1592 1120 1599 1122
rect 1592 1119 1593 1120
rect 1587 1118 1593 1119
rect 1598 1119 1599 1120
rect 1603 1119 1604 1123
rect 1598 1118 1604 1119
rect 1618 1123 1624 1124
rect 1618 1119 1619 1123
rect 1623 1122 1624 1123
rect 1651 1123 1657 1124
rect 1651 1122 1652 1123
rect 1623 1120 1652 1122
rect 1623 1119 1624 1120
rect 1618 1118 1624 1119
rect 1651 1119 1652 1120
rect 1656 1119 1657 1123
rect 1707 1121 1708 1125
rect 1712 1121 1713 1125
rect 1707 1120 1713 1121
rect 1738 1123 1744 1124
rect 1651 1118 1657 1119
rect 1738 1119 1739 1123
rect 1743 1122 1744 1123
rect 1763 1123 1769 1124
rect 1763 1122 1764 1123
rect 1743 1120 1764 1122
rect 1743 1119 1744 1120
rect 1738 1118 1744 1119
rect 1763 1119 1764 1120
rect 1768 1119 1769 1123
rect 1763 1118 1769 1119
rect 1794 1123 1800 1124
rect 1794 1119 1795 1123
rect 1799 1122 1800 1123
rect 1819 1123 1825 1124
rect 1819 1122 1820 1123
rect 1799 1120 1820 1122
rect 1799 1119 1800 1120
rect 1794 1118 1800 1119
rect 1819 1119 1820 1120
rect 1824 1119 1825 1123
rect 1819 1118 1825 1119
rect 1850 1123 1856 1124
rect 1850 1119 1851 1123
rect 1855 1122 1856 1123
rect 1867 1123 1873 1124
rect 1867 1122 1868 1123
rect 1855 1120 1868 1122
rect 1855 1119 1856 1120
rect 1850 1118 1856 1119
rect 1867 1119 1868 1120
rect 1872 1119 1873 1123
rect 1867 1118 1873 1119
rect 1898 1123 1904 1124
rect 1898 1119 1899 1123
rect 1903 1122 1904 1123
rect 1923 1123 1929 1124
rect 1923 1122 1924 1123
rect 1903 1120 1924 1122
rect 1903 1119 1904 1120
rect 1898 1118 1904 1119
rect 1923 1119 1924 1120
rect 1928 1119 1929 1123
rect 1923 1118 1929 1119
rect 1954 1123 1960 1124
rect 1954 1119 1955 1123
rect 1959 1122 1960 1123
rect 1979 1123 1985 1124
rect 1979 1122 1980 1123
rect 1959 1120 1980 1122
rect 1959 1119 1960 1120
rect 1954 1118 1960 1119
rect 1979 1119 1980 1120
rect 1984 1119 1985 1123
rect 1979 1118 1985 1119
rect 2027 1123 2033 1124
rect 2027 1119 2028 1123
rect 2032 1122 2033 1123
rect 2046 1123 2052 1124
rect 2046 1122 2047 1123
rect 2032 1120 2047 1122
rect 2032 1119 2033 1120
rect 2027 1118 2033 1119
rect 2046 1119 2047 1120
rect 2051 1119 2052 1123
rect 2046 1118 2052 1119
rect 2067 1123 2073 1124
rect 2067 1119 2068 1123
rect 2072 1122 2073 1123
rect 2078 1123 2084 1124
rect 2078 1122 2079 1123
rect 2072 1120 2079 1122
rect 2072 1119 2073 1120
rect 2067 1118 2073 1119
rect 2078 1119 2079 1120
rect 2083 1119 2084 1123
rect 2078 1118 2084 1119
rect 1015 1114 1021 1115
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 110 1107 116 1108
rect 110 1103 111 1107
rect 115 1103 116 1107
rect 1094 1107 1100 1108
rect 1382 1107 1388 1108
rect 1422 1112 1428 1113
rect 1422 1108 1423 1112
rect 1427 1108 1428 1112
rect 1422 1107 1428 1108
rect 1470 1112 1476 1113
rect 1470 1108 1471 1112
rect 1475 1108 1476 1112
rect 1470 1107 1476 1108
rect 1526 1112 1532 1113
rect 1526 1108 1527 1112
rect 1531 1108 1532 1112
rect 1526 1107 1532 1108
rect 1590 1112 1596 1113
rect 1590 1108 1591 1112
rect 1595 1108 1596 1112
rect 1590 1107 1596 1108
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1710 1112 1716 1113
rect 1710 1108 1711 1112
rect 1715 1108 1716 1112
rect 1710 1107 1716 1108
rect 1766 1112 1772 1113
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1822 1112 1828 1113
rect 1822 1108 1823 1112
rect 1827 1108 1828 1112
rect 1822 1107 1828 1108
rect 1870 1112 1876 1113
rect 1870 1108 1871 1112
rect 1875 1108 1876 1112
rect 1870 1107 1876 1108
rect 1926 1112 1932 1113
rect 1926 1108 1927 1112
rect 1931 1108 1932 1112
rect 1926 1107 1932 1108
rect 1982 1112 1988 1113
rect 1982 1108 1983 1112
rect 1987 1108 1988 1112
rect 1982 1107 1988 1108
rect 2030 1112 2036 1113
rect 2030 1108 2031 1112
rect 2035 1108 2036 1112
rect 2030 1107 2036 1108
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 110 1102 116 1103
rect 158 1104 164 1105
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 246 1104 252 1105
rect 246 1100 247 1104
rect 251 1100 252 1104
rect 246 1099 252 1100
rect 302 1104 308 1105
rect 302 1100 303 1104
rect 307 1100 308 1104
rect 302 1099 308 1100
rect 366 1104 372 1105
rect 366 1100 367 1104
rect 371 1100 372 1104
rect 366 1099 372 1100
rect 438 1104 444 1105
rect 438 1100 439 1104
rect 443 1100 444 1104
rect 438 1099 444 1100
rect 510 1104 516 1105
rect 510 1100 511 1104
rect 515 1100 516 1104
rect 510 1099 516 1100
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 678 1104 684 1105
rect 678 1100 679 1104
rect 683 1100 684 1104
rect 678 1099 684 1100
rect 774 1104 780 1105
rect 774 1100 775 1104
rect 779 1100 780 1104
rect 774 1099 780 1100
rect 878 1104 884 1105
rect 878 1100 879 1104
rect 883 1100 884 1104
rect 878 1099 884 1100
rect 990 1104 996 1105
rect 990 1100 991 1104
rect 995 1100 996 1104
rect 1094 1103 1095 1107
rect 1099 1103 1100 1107
rect 1094 1102 1100 1103
rect 1134 1104 1140 1105
rect 990 1099 996 1100
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 1134 1099 1140 1100
rect 1406 1099 1413 1100
rect 1406 1095 1407 1099
rect 1412 1095 1413 1099
rect 1406 1094 1413 1095
rect 1447 1099 1456 1100
rect 1447 1095 1448 1099
rect 1455 1095 1456 1099
rect 1447 1094 1456 1095
rect 1494 1099 1501 1100
rect 1494 1095 1495 1099
rect 1500 1095 1501 1099
rect 1494 1094 1501 1095
rect 1550 1099 1557 1100
rect 1550 1095 1551 1099
rect 1556 1095 1557 1099
rect 1550 1094 1557 1095
rect 1615 1099 1624 1100
rect 1615 1095 1616 1099
rect 1623 1095 1624 1099
rect 1615 1094 1624 1095
rect 1678 1099 1685 1100
rect 1678 1095 1679 1099
rect 1684 1095 1685 1099
rect 1678 1094 1685 1095
rect 1735 1099 1744 1100
rect 1735 1095 1736 1099
rect 1743 1095 1744 1099
rect 1735 1094 1744 1095
rect 1791 1099 1800 1100
rect 1791 1095 1792 1099
rect 1799 1095 1800 1099
rect 1791 1094 1800 1095
rect 1847 1099 1856 1100
rect 1847 1095 1848 1099
rect 1855 1095 1856 1099
rect 1847 1094 1856 1095
rect 1895 1099 1904 1100
rect 1895 1095 1896 1099
rect 1903 1095 1904 1099
rect 1895 1094 1904 1095
rect 1951 1099 1960 1100
rect 1951 1095 1952 1099
rect 1959 1095 1960 1099
rect 1951 1094 1960 1095
rect 1998 1099 2004 1100
rect 1998 1095 1999 1099
rect 2003 1098 2004 1099
rect 2007 1099 2013 1100
rect 2007 1098 2008 1099
rect 2003 1096 2008 1098
rect 2003 1095 2004 1096
rect 1998 1094 2004 1095
rect 2007 1095 2008 1096
rect 2012 1095 2013 1099
rect 2007 1094 2013 1095
rect 2054 1099 2061 1100
rect 2054 1095 2055 1099
rect 2060 1095 2061 1099
rect 2054 1094 2061 1095
rect 2078 1099 2084 1100
rect 2078 1095 2079 1099
rect 2083 1098 2084 1099
rect 2095 1099 2101 1100
rect 2118 1099 2124 1100
rect 2095 1098 2096 1099
rect 2083 1096 2096 1098
rect 2083 1095 2084 1096
rect 2078 1094 2084 1095
rect 2095 1095 2096 1096
rect 2100 1095 2101 1099
rect 2095 1094 2101 1095
rect 1134 1087 1140 1088
rect 198 1084 204 1085
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 198 1080 199 1084
rect 203 1080 204 1084
rect 198 1079 204 1080
rect 246 1084 252 1085
rect 246 1080 247 1084
rect 251 1080 252 1084
rect 246 1079 252 1080
rect 302 1084 308 1085
rect 302 1080 303 1084
rect 307 1080 308 1084
rect 302 1079 308 1080
rect 366 1084 372 1085
rect 366 1080 367 1084
rect 371 1080 372 1084
rect 366 1079 372 1080
rect 430 1084 436 1085
rect 430 1080 431 1084
rect 435 1080 436 1084
rect 430 1079 436 1080
rect 502 1084 508 1085
rect 502 1080 503 1084
rect 507 1080 508 1084
rect 502 1079 508 1080
rect 574 1084 580 1085
rect 574 1080 575 1084
rect 579 1080 580 1084
rect 574 1079 580 1080
rect 646 1084 652 1085
rect 646 1080 647 1084
rect 651 1080 652 1084
rect 646 1079 652 1080
rect 718 1084 724 1085
rect 718 1080 719 1084
rect 723 1080 724 1084
rect 718 1079 724 1080
rect 782 1084 788 1085
rect 782 1080 783 1084
rect 787 1080 788 1084
rect 782 1079 788 1080
rect 838 1084 844 1085
rect 838 1080 839 1084
rect 843 1080 844 1084
rect 838 1079 844 1080
rect 894 1084 900 1085
rect 894 1080 895 1084
rect 899 1080 900 1084
rect 894 1079 900 1080
rect 950 1084 956 1085
rect 950 1080 951 1084
rect 955 1080 956 1084
rect 950 1079 956 1080
rect 1006 1084 1012 1085
rect 1006 1080 1007 1084
rect 1011 1080 1012 1084
rect 1006 1079 1012 1080
rect 1046 1084 1052 1085
rect 1046 1080 1047 1084
rect 1051 1080 1052 1084
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 2118 1087 2124 1088
rect 1134 1082 1140 1083
rect 1382 1084 1388 1085
rect 1046 1079 1052 1080
rect 1094 1081 1100 1082
rect 110 1076 116 1077
rect 1094 1077 1095 1081
rect 1099 1077 1100 1081
rect 1382 1080 1383 1084
rect 1387 1080 1388 1084
rect 1382 1079 1388 1080
rect 1422 1084 1428 1085
rect 1422 1080 1423 1084
rect 1427 1080 1428 1084
rect 1422 1079 1428 1080
rect 1470 1084 1476 1085
rect 1470 1080 1471 1084
rect 1475 1080 1476 1084
rect 1470 1079 1476 1080
rect 1526 1084 1532 1085
rect 1526 1080 1527 1084
rect 1531 1080 1532 1084
rect 1526 1079 1532 1080
rect 1590 1084 1596 1085
rect 1590 1080 1591 1084
rect 1595 1080 1596 1084
rect 1590 1079 1596 1080
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1710 1084 1716 1085
rect 1710 1080 1711 1084
rect 1715 1080 1716 1084
rect 1710 1079 1716 1080
rect 1766 1084 1772 1085
rect 1766 1080 1767 1084
rect 1771 1080 1772 1084
rect 1766 1079 1772 1080
rect 1822 1084 1828 1085
rect 1822 1080 1823 1084
rect 1827 1080 1828 1084
rect 1822 1079 1828 1080
rect 1870 1084 1876 1085
rect 1870 1080 1871 1084
rect 1875 1080 1876 1084
rect 1870 1079 1876 1080
rect 1926 1084 1932 1085
rect 1926 1080 1927 1084
rect 1931 1080 1932 1084
rect 1926 1079 1932 1080
rect 1982 1084 1988 1085
rect 1982 1080 1983 1084
rect 1987 1080 1988 1084
rect 1982 1079 1988 1080
rect 2030 1084 2036 1085
rect 2030 1080 2031 1084
rect 2035 1080 2036 1084
rect 2030 1079 2036 1080
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2070 1079 2076 1080
rect 1094 1076 1100 1077
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 174 1067 180 1068
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 174 1063 175 1067
rect 179 1066 180 1067
rect 223 1067 229 1068
rect 223 1066 224 1067
rect 179 1064 224 1066
rect 179 1063 180 1064
rect 174 1062 180 1063
rect 223 1063 224 1064
rect 228 1063 229 1067
rect 223 1062 229 1063
rect 231 1067 237 1068
rect 231 1063 232 1067
rect 236 1066 237 1067
rect 271 1067 277 1068
rect 271 1066 272 1067
rect 236 1064 272 1066
rect 236 1063 237 1064
rect 231 1062 237 1063
rect 271 1063 272 1064
rect 276 1063 277 1067
rect 271 1062 277 1063
rect 279 1067 285 1068
rect 279 1063 280 1067
rect 284 1066 285 1067
rect 327 1067 333 1068
rect 327 1066 328 1067
rect 284 1064 328 1066
rect 284 1063 285 1064
rect 279 1062 285 1063
rect 327 1063 328 1064
rect 332 1063 333 1067
rect 327 1062 333 1063
rect 346 1067 352 1068
rect 346 1063 347 1067
rect 351 1066 352 1067
rect 391 1067 397 1068
rect 391 1066 392 1067
rect 351 1064 392 1066
rect 351 1063 352 1064
rect 346 1062 352 1063
rect 391 1063 392 1064
rect 396 1063 397 1067
rect 391 1062 397 1063
rect 399 1067 405 1068
rect 399 1063 400 1067
rect 404 1066 405 1067
rect 455 1067 461 1068
rect 455 1066 456 1067
rect 404 1064 456 1066
rect 404 1063 405 1064
rect 399 1062 405 1063
rect 455 1063 456 1064
rect 460 1063 461 1067
rect 455 1062 461 1063
rect 527 1067 533 1068
rect 527 1063 528 1067
rect 532 1066 533 1067
rect 566 1067 572 1068
rect 566 1066 567 1067
rect 532 1064 567 1066
rect 532 1063 533 1064
rect 527 1062 533 1063
rect 566 1063 567 1064
rect 571 1063 572 1067
rect 566 1062 572 1063
rect 599 1067 605 1068
rect 599 1063 600 1067
rect 604 1066 605 1067
rect 638 1067 644 1068
rect 638 1066 639 1067
rect 604 1064 639 1066
rect 604 1063 605 1064
rect 599 1062 605 1063
rect 638 1063 639 1064
rect 643 1063 644 1067
rect 638 1062 644 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1066 660 1067
rect 671 1067 677 1068
rect 671 1066 672 1067
rect 659 1064 672 1066
rect 659 1063 660 1064
rect 654 1062 660 1063
rect 671 1063 672 1064
rect 676 1063 677 1067
rect 671 1062 677 1063
rect 743 1067 749 1068
rect 743 1063 744 1067
rect 748 1066 749 1067
rect 774 1067 780 1068
rect 774 1066 775 1067
rect 748 1064 775 1066
rect 748 1063 749 1064
rect 743 1062 749 1063
rect 774 1063 775 1064
rect 779 1063 780 1067
rect 774 1062 780 1063
rect 807 1067 813 1068
rect 807 1063 808 1067
rect 812 1066 813 1067
rect 830 1067 836 1068
rect 830 1066 831 1067
rect 812 1064 831 1066
rect 812 1063 813 1064
rect 807 1062 813 1063
rect 830 1063 831 1064
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 863 1067 869 1068
rect 863 1063 864 1067
rect 868 1066 869 1067
rect 910 1067 916 1068
rect 910 1066 911 1067
rect 868 1064 911 1066
rect 868 1063 869 1064
rect 863 1062 869 1063
rect 910 1063 911 1064
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 919 1067 925 1068
rect 919 1063 920 1067
rect 924 1066 925 1067
rect 942 1067 948 1068
rect 942 1066 943 1067
rect 924 1064 943 1066
rect 924 1063 925 1064
rect 919 1062 925 1063
rect 942 1063 943 1064
rect 947 1063 948 1067
rect 942 1062 948 1063
rect 975 1067 981 1068
rect 975 1063 976 1067
rect 980 1066 981 1067
rect 998 1067 1004 1068
rect 998 1066 999 1067
rect 980 1064 999 1066
rect 980 1063 981 1064
rect 975 1062 981 1063
rect 998 1063 999 1064
rect 1003 1063 1004 1067
rect 998 1062 1004 1063
rect 1031 1067 1040 1068
rect 1031 1063 1032 1067
rect 1039 1063 1040 1067
rect 1031 1062 1040 1063
rect 1071 1067 1077 1068
rect 1071 1063 1072 1067
rect 1076 1066 1077 1067
rect 1086 1067 1092 1068
rect 1086 1066 1087 1067
rect 1076 1064 1087 1066
rect 1076 1063 1077 1064
rect 1071 1062 1077 1063
rect 1086 1063 1087 1064
rect 1091 1063 1092 1067
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1358 1072 1364 1073
rect 1358 1068 1359 1072
rect 1363 1068 1364 1072
rect 1358 1067 1364 1068
rect 1470 1072 1476 1073
rect 1470 1068 1471 1072
rect 1475 1068 1476 1072
rect 1470 1067 1476 1068
rect 1574 1072 1580 1073
rect 1574 1068 1575 1072
rect 1579 1068 1580 1072
rect 1574 1067 1580 1068
rect 1670 1072 1676 1073
rect 1670 1068 1671 1072
rect 1675 1068 1676 1072
rect 1670 1067 1676 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1846 1072 1852 1073
rect 1846 1068 1847 1072
rect 1851 1068 1852 1072
rect 1846 1067 1852 1068
rect 1926 1072 1932 1073
rect 1926 1068 1927 1072
rect 1931 1068 1932 1072
rect 1926 1067 1932 1068
rect 2006 1072 2012 1073
rect 2006 1068 2007 1072
rect 2011 1068 2012 1072
rect 2006 1067 2012 1068
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 2118 1069 2124 1070
rect 1086 1062 1092 1063
rect 1094 1064 1100 1065
rect 1134 1064 1140 1065
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 110 1059 116 1060
rect 1094 1060 1095 1064
rect 1099 1060 1100 1064
rect 1702 1063 1708 1064
rect 1176 1060 1362 1062
rect 1094 1059 1100 1060
rect 1174 1059 1180 1060
rect 198 1056 204 1057
rect 198 1052 199 1056
rect 203 1052 204 1056
rect 198 1051 204 1052
rect 246 1056 252 1057
rect 246 1052 247 1056
rect 251 1052 252 1056
rect 246 1051 252 1052
rect 302 1056 308 1057
rect 302 1052 303 1056
rect 307 1052 308 1056
rect 302 1051 308 1052
rect 366 1056 372 1057
rect 366 1052 367 1056
rect 371 1052 372 1056
rect 366 1051 372 1052
rect 430 1056 436 1057
rect 430 1052 431 1056
rect 435 1052 436 1056
rect 430 1051 436 1052
rect 502 1056 508 1057
rect 502 1052 503 1056
rect 507 1052 508 1056
rect 502 1051 508 1052
rect 574 1056 580 1057
rect 574 1052 575 1056
rect 579 1052 580 1056
rect 574 1051 580 1052
rect 646 1056 652 1057
rect 646 1052 647 1056
rect 651 1052 652 1056
rect 646 1051 652 1052
rect 718 1056 724 1057
rect 718 1052 719 1056
rect 723 1052 724 1056
rect 718 1051 724 1052
rect 782 1056 788 1057
rect 782 1052 783 1056
rect 787 1052 788 1056
rect 782 1051 788 1052
rect 838 1056 844 1057
rect 838 1052 839 1056
rect 843 1052 844 1056
rect 838 1051 844 1052
rect 894 1056 900 1057
rect 894 1052 895 1056
rect 899 1052 900 1056
rect 894 1051 900 1052
rect 950 1056 956 1057
rect 950 1052 951 1056
rect 955 1052 956 1056
rect 950 1051 956 1052
rect 1006 1056 1012 1057
rect 1006 1052 1007 1056
rect 1011 1052 1012 1056
rect 1006 1051 1012 1052
rect 1046 1056 1052 1057
rect 1046 1052 1047 1056
rect 1051 1052 1052 1056
rect 1174 1055 1175 1059
rect 1179 1055 1180 1059
rect 1174 1054 1180 1055
rect 1183 1055 1189 1056
rect 1046 1051 1052 1052
rect 1134 1052 1140 1053
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1183 1051 1184 1055
rect 1188 1054 1189 1055
rect 1238 1055 1244 1056
rect 1238 1054 1239 1055
rect 1188 1052 1239 1054
rect 1188 1051 1189 1052
rect 1183 1050 1189 1051
rect 1238 1051 1239 1052
rect 1243 1051 1244 1055
rect 1238 1050 1244 1051
rect 1271 1055 1277 1056
rect 1271 1051 1272 1055
rect 1276 1054 1277 1055
rect 1350 1055 1356 1056
rect 1350 1054 1351 1055
rect 1276 1052 1351 1054
rect 1276 1051 1277 1052
rect 1271 1050 1277 1051
rect 1350 1051 1351 1052
rect 1355 1051 1356 1055
rect 1360 1054 1362 1060
rect 1702 1059 1703 1063
rect 1707 1062 1708 1063
rect 1707 1060 1826 1062
rect 1707 1059 1708 1060
rect 1702 1058 1708 1059
rect 1383 1055 1389 1056
rect 1383 1054 1384 1055
rect 1360 1052 1384 1054
rect 1350 1050 1356 1051
rect 1383 1051 1384 1052
rect 1388 1051 1389 1055
rect 1383 1050 1389 1051
rect 1495 1055 1501 1056
rect 1495 1051 1496 1055
rect 1500 1054 1501 1055
rect 1566 1055 1572 1056
rect 1566 1054 1567 1055
rect 1500 1052 1567 1054
rect 1500 1051 1501 1052
rect 1495 1050 1501 1051
rect 1566 1051 1567 1052
rect 1571 1051 1572 1055
rect 1566 1050 1572 1051
rect 1598 1055 1605 1056
rect 1598 1051 1599 1055
rect 1604 1051 1605 1055
rect 1598 1050 1605 1051
rect 1695 1055 1701 1056
rect 1695 1051 1696 1055
rect 1700 1054 1701 1055
rect 1750 1055 1756 1056
rect 1750 1054 1751 1055
rect 1700 1052 1751 1054
rect 1700 1051 1701 1052
rect 1695 1050 1701 1051
rect 1750 1051 1751 1052
rect 1755 1051 1756 1055
rect 1750 1050 1756 1051
rect 1783 1055 1789 1056
rect 1783 1051 1784 1055
rect 1788 1054 1789 1055
rect 1814 1055 1820 1056
rect 1814 1054 1815 1055
rect 1788 1052 1815 1054
rect 1788 1051 1789 1052
rect 1783 1050 1789 1051
rect 1814 1051 1815 1052
rect 1819 1051 1820 1055
rect 1824 1054 1826 1060
rect 1871 1055 1877 1056
rect 1871 1054 1872 1055
rect 1824 1052 1872 1054
rect 1814 1050 1820 1051
rect 1871 1051 1872 1052
rect 1876 1051 1877 1055
rect 1871 1050 1877 1051
rect 1879 1055 1885 1056
rect 1879 1051 1880 1055
rect 1884 1054 1885 1055
rect 1951 1055 1957 1056
rect 1951 1054 1952 1055
rect 1884 1052 1952 1054
rect 1884 1051 1885 1052
rect 1879 1050 1885 1051
rect 1951 1051 1952 1052
rect 1956 1051 1957 1055
rect 1951 1050 1957 1051
rect 1959 1055 1965 1056
rect 1959 1051 1960 1055
rect 1964 1054 1965 1055
rect 2031 1055 2037 1056
rect 2031 1054 2032 1055
rect 1964 1052 2032 1054
rect 1964 1051 1965 1052
rect 1959 1050 1965 1051
rect 2031 1051 2032 1052
rect 2036 1051 2037 1055
rect 2031 1050 2037 1051
rect 2046 1055 2052 1056
rect 2046 1051 2047 1055
rect 2051 1054 2052 1055
rect 2095 1055 2101 1056
rect 2095 1054 2096 1055
rect 2051 1052 2096 1054
rect 2051 1051 2052 1052
rect 2046 1050 2052 1051
rect 2095 1051 2096 1052
rect 2100 1051 2101 1055
rect 2095 1050 2101 1051
rect 2118 1052 2124 1053
rect 1134 1047 1140 1048
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 1158 1044 1164 1045
rect 195 1043 201 1044
rect 195 1039 196 1043
rect 200 1042 201 1043
rect 231 1043 237 1044
rect 231 1042 232 1043
rect 200 1040 232 1042
rect 200 1039 201 1040
rect 195 1038 201 1039
rect 231 1039 232 1040
rect 236 1039 237 1043
rect 231 1038 237 1039
rect 243 1043 249 1044
rect 243 1039 244 1043
rect 248 1042 249 1043
rect 279 1043 285 1044
rect 279 1042 280 1043
rect 248 1040 280 1042
rect 248 1039 249 1040
rect 243 1038 249 1039
rect 279 1039 280 1040
rect 284 1039 285 1043
rect 279 1038 285 1039
rect 299 1043 305 1044
rect 299 1039 300 1043
rect 304 1042 305 1043
rect 346 1043 352 1044
rect 346 1042 347 1043
rect 304 1040 347 1042
rect 304 1039 305 1040
rect 299 1038 305 1039
rect 346 1039 347 1040
rect 351 1039 352 1043
rect 346 1038 352 1039
rect 363 1043 369 1044
rect 363 1039 364 1043
rect 368 1042 369 1043
rect 399 1043 405 1044
rect 399 1042 400 1043
rect 368 1040 400 1042
rect 368 1039 369 1040
rect 363 1038 369 1039
rect 399 1039 400 1040
rect 404 1039 405 1043
rect 399 1038 405 1039
rect 422 1043 433 1044
rect 422 1039 423 1043
rect 427 1039 428 1043
rect 432 1039 433 1043
rect 422 1038 433 1039
rect 499 1043 505 1044
rect 499 1039 500 1043
rect 504 1042 505 1043
rect 518 1043 524 1044
rect 518 1042 519 1043
rect 504 1040 519 1042
rect 504 1039 505 1040
rect 499 1038 505 1039
rect 518 1039 519 1040
rect 523 1039 524 1043
rect 518 1038 524 1039
rect 566 1043 577 1044
rect 566 1039 567 1043
rect 571 1039 572 1043
rect 576 1039 577 1043
rect 566 1038 577 1039
rect 638 1043 649 1044
rect 638 1039 639 1043
rect 643 1039 644 1043
rect 648 1039 649 1043
rect 638 1038 649 1039
rect 715 1043 721 1044
rect 715 1039 716 1043
rect 720 1042 721 1043
rect 774 1043 785 1044
rect 720 1040 770 1042
rect 720 1039 721 1040
rect 715 1038 721 1039
rect 768 1034 770 1040
rect 774 1039 775 1043
rect 779 1039 780 1043
rect 784 1039 785 1043
rect 774 1038 785 1039
rect 830 1043 841 1044
rect 830 1039 831 1043
rect 835 1039 836 1043
rect 840 1039 841 1043
rect 830 1038 841 1039
rect 891 1043 897 1044
rect 891 1039 892 1043
rect 896 1042 897 1043
rect 926 1043 932 1044
rect 926 1042 927 1043
rect 896 1040 927 1042
rect 896 1039 897 1040
rect 891 1038 897 1039
rect 926 1039 927 1040
rect 931 1039 932 1043
rect 926 1038 932 1039
rect 942 1043 953 1044
rect 942 1039 943 1043
rect 947 1039 948 1043
rect 952 1039 953 1043
rect 942 1038 953 1039
rect 998 1043 1009 1044
rect 998 1039 999 1043
rect 1003 1039 1004 1043
rect 1008 1039 1009 1043
rect 998 1038 1009 1039
rect 1034 1043 1040 1044
rect 1034 1039 1035 1043
rect 1039 1042 1040 1043
rect 1043 1043 1049 1044
rect 1043 1042 1044 1043
rect 1039 1040 1044 1042
rect 1039 1039 1040 1040
rect 1034 1038 1040 1039
rect 1043 1039 1044 1040
rect 1048 1039 1049 1043
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1358 1044 1364 1045
rect 1358 1040 1359 1044
rect 1363 1040 1364 1044
rect 1358 1039 1364 1040
rect 1470 1044 1476 1045
rect 1470 1040 1471 1044
rect 1475 1040 1476 1044
rect 1470 1039 1476 1040
rect 1574 1044 1580 1045
rect 1574 1040 1575 1044
rect 1579 1040 1580 1044
rect 1574 1039 1580 1040
rect 1670 1044 1676 1045
rect 1670 1040 1671 1044
rect 1675 1040 1676 1044
rect 1670 1039 1676 1040
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1846 1044 1852 1045
rect 1846 1040 1847 1044
rect 1851 1040 1852 1044
rect 1846 1039 1852 1040
rect 1926 1044 1932 1045
rect 1926 1040 1927 1044
rect 1931 1040 1932 1044
rect 1926 1039 1932 1040
rect 2006 1044 2012 1045
rect 2006 1040 2007 1044
rect 2011 1040 2012 1044
rect 2006 1039 2012 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 1043 1038 1049 1039
rect 810 1035 816 1036
rect 810 1034 811 1035
rect 768 1032 811 1034
rect 810 1031 811 1032
rect 815 1031 816 1035
rect 810 1030 816 1031
rect 1086 1031 1092 1032
rect 219 1027 225 1028
rect 219 1023 220 1027
rect 224 1026 225 1027
rect 238 1027 244 1028
rect 238 1026 239 1027
rect 224 1024 239 1026
rect 224 1023 225 1024
rect 219 1022 225 1023
rect 238 1023 239 1024
rect 243 1023 244 1027
rect 238 1022 244 1023
rect 254 1027 260 1028
rect 254 1023 255 1027
rect 259 1026 260 1027
rect 267 1027 273 1028
rect 267 1026 268 1027
rect 259 1024 268 1026
rect 259 1023 260 1024
rect 254 1022 260 1023
rect 267 1023 268 1024
rect 272 1023 273 1027
rect 267 1022 273 1023
rect 303 1027 309 1028
rect 303 1023 304 1027
rect 308 1026 309 1027
rect 331 1027 337 1028
rect 331 1026 332 1027
rect 308 1024 332 1026
rect 308 1023 309 1024
rect 303 1022 309 1023
rect 331 1023 332 1024
rect 336 1023 337 1027
rect 331 1022 337 1023
rect 378 1027 384 1028
rect 378 1023 379 1027
rect 383 1026 384 1027
rect 403 1027 409 1028
rect 403 1026 404 1027
rect 383 1024 404 1026
rect 383 1023 384 1024
rect 378 1022 384 1023
rect 403 1023 404 1024
rect 408 1023 409 1027
rect 403 1022 409 1023
rect 475 1027 481 1028
rect 475 1023 476 1027
rect 480 1026 481 1027
rect 546 1027 552 1028
rect 546 1026 547 1027
rect 480 1024 547 1026
rect 480 1023 481 1024
rect 475 1022 481 1023
rect 546 1023 547 1024
rect 551 1023 552 1027
rect 546 1022 552 1023
rect 555 1027 561 1028
rect 555 1023 556 1027
rect 560 1026 561 1027
rect 618 1027 624 1028
rect 618 1026 619 1027
rect 560 1024 619 1026
rect 560 1023 561 1024
rect 555 1022 561 1023
rect 618 1023 619 1024
rect 623 1023 624 1027
rect 618 1022 624 1023
rect 627 1027 633 1028
rect 627 1023 628 1027
rect 632 1026 633 1027
rect 654 1027 660 1028
rect 654 1026 655 1027
rect 632 1024 655 1026
rect 632 1023 633 1024
rect 627 1022 633 1023
rect 654 1023 655 1024
rect 659 1023 660 1027
rect 654 1022 660 1023
rect 699 1027 705 1028
rect 699 1023 700 1027
rect 704 1026 705 1027
rect 710 1027 716 1028
rect 710 1026 711 1027
rect 704 1024 711 1026
rect 704 1023 705 1024
rect 699 1022 705 1023
rect 710 1023 711 1024
rect 715 1023 716 1027
rect 710 1022 716 1023
rect 730 1027 736 1028
rect 730 1023 731 1027
rect 735 1026 736 1027
rect 771 1027 777 1028
rect 771 1026 772 1027
rect 735 1024 772 1026
rect 735 1023 736 1024
rect 730 1022 736 1023
rect 771 1023 772 1024
rect 776 1023 777 1027
rect 771 1022 777 1023
rect 802 1027 808 1028
rect 802 1023 803 1027
rect 807 1026 808 1027
rect 835 1027 841 1028
rect 835 1026 836 1027
rect 807 1024 836 1026
rect 807 1023 808 1024
rect 802 1022 808 1023
rect 835 1023 836 1024
rect 840 1023 841 1027
rect 835 1022 841 1023
rect 866 1027 872 1028
rect 866 1023 867 1027
rect 871 1026 872 1027
rect 899 1027 905 1028
rect 899 1026 900 1027
rect 871 1024 900 1026
rect 871 1023 872 1024
rect 866 1022 872 1023
rect 899 1023 900 1024
rect 904 1023 905 1027
rect 899 1022 905 1023
rect 910 1027 916 1028
rect 910 1023 911 1027
rect 915 1026 916 1027
rect 963 1027 969 1028
rect 963 1026 964 1027
rect 915 1024 964 1026
rect 915 1023 916 1024
rect 910 1022 916 1023
rect 963 1023 964 1024
rect 968 1023 969 1027
rect 963 1022 969 1023
rect 994 1027 1000 1028
rect 994 1023 995 1027
rect 999 1026 1000 1027
rect 1035 1027 1041 1028
rect 1035 1026 1036 1027
rect 999 1024 1036 1026
rect 999 1023 1000 1024
rect 994 1022 1000 1023
rect 1035 1023 1036 1024
rect 1040 1023 1041 1027
rect 1086 1027 1087 1031
rect 1091 1030 1092 1031
rect 1155 1031 1161 1032
rect 1155 1030 1156 1031
rect 1091 1028 1156 1030
rect 1091 1027 1092 1028
rect 1086 1026 1092 1027
rect 1155 1027 1156 1028
rect 1160 1027 1161 1031
rect 1155 1026 1161 1027
rect 1238 1031 1249 1032
rect 1238 1027 1239 1031
rect 1243 1027 1244 1031
rect 1248 1027 1249 1031
rect 1238 1026 1249 1027
rect 1350 1031 1361 1032
rect 1350 1027 1351 1031
rect 1355 1027 1356 1031
rect 1360 1027 1361 1031
rect 1350 1026 1361 1027
rect 1467 1031 1473 1032
rect 1467 1027 1468 1031
rect 1472 1030 1473 1031
rect 1486 1031 1492 1032
rect 1486 1030 1487 1031
rect 1472 1028 1487 1030
rect 1472 1027 1473 1028
rect 1467 1026 1473 1027
rect 1486 1027 1487 1028
rect 1491 1027 1492 1031
rect 1486 1026 1492 1027
rect 1566 1031 1577 1032
rect 1566 1027 1567 1031
rect 1571 1027 1572 1031
rect 1576 1027 1577 1031
rect 1566 1026 1577 1027
rect 1667 1031 1673 1032
rect 1667 1027 1668 1031
rect 1672 1030 1673 1031
rect 1702 1031 1708 1032
rect 1702 1030 1703 1031
rect 1672 1028 1703 1030
rect 1672 1027 1673 1028
rect 1667 1026 1673 1027
rect 1702 1027 1703 1028
rect 1707 1027 1708 1031
rect 1702 1026 1708 1027
rect 1750 1031 1761 1032
rect 1750 1027 1751 1031
rect 1755 1027 1756 1031
rect 1760 1027 1761 1031
rect 1750 1026 1761 1027
rect 1843 1031 1849 1032
rect 1843 1027 1844 1031
rect 1848 1030 1849 1031
rect 1879 1031 1885 1032
rect 1879 1030 1880 1031
rect 1848 1028 1880 1030
rect 1848 1027 1849 1028
rect 1843 1026 1849 1027
rect 1879 1027 1880 1028
rect 1884 1027 1885 1031
rect 1879 1026 1885 1027
rect 1923 1031 1929 1032
rect 1923 1027 1924 1031
rect 1928 1030 1929 1031
rect 1959 1031 1965 1032
rect 1959 1030 1960 1031
rect 1928 1028 1960 1030
rect 1928 1027 1929 1028
rect 1923 1026 1929 1027
rect 1959 1027 1960 1028
rect 1964 1027 1965 1031
rect 1959 1026 1965 1027
rect 1998 1031 2009 1032
rect 1998 1027 1999 1031
rect 2003 1027 2004 1031
rect 2008 1027 2009 1031
rect 1998 1026 2009 1027
rect 2067 1031 2073 1032
rect 2067 1027 2068 1031
rect 2072 1030 2073 1031
rect 2078 1031 2084 1032
rect 2078 1030 2079 1031
rect 2072 1028 2079 1030
rect 2072 1027 2073 1028
rect 2067 1026 2073 1027
rect 2078 1027 2079 1028
rect 2083 1027 2084 1031
rect 2078 1026 2084 1027
rect 1035 1022 1041 1023
rect 1155 1019 1161 1020
rect 222 1016 228 1017
rect 222 1012 223 1016
rect 227 1012 228 1016
rect 222 1011 228 1012
rect 270 1016 276 1017
rect 270 1012 271 1016
rect 275 1012 276 1016
rect 270 1011 276 1012
rect 334 1016 340 1017
rect 334 1012 335 1016
rect 339 1012 340 1016
rect 334 1011 340 1012
rect 406 1016 412 1017
rect 406 1012 407 1016
rect 411 1012 412 1016
rect 406 1011 412 1012
rect 478 1016 484 1017
rect 478 1012 479 1016
rect 483 1012 484 1016
rect 478 1011 484 1012
rect 558 1016 564 1017
rect 558 1012 559 1016
rect 563 1012 564 1016
rect 558 1011 564 1012
rect 630 1016 636 1017
rect 630 1012 631 1016
rect 635 1012 636 1016
rect 630 1011 636 1012
rect 702 1016 708 1017
rect 702 1012 703 1016
rect 707 1012 708 1016
rect 702 1011 708 1012
rect 774 1016 780 1017
rect 774 1012 775 1016
rect 779 1012 780 1016
rect 774 1011 780 1012
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 902 1016 908 1017
rect 902 1012 903 1016
rect 907 1012 908 1016
rect 902 1011 908 1012
rect 966 1016 972 1017
rect 966 1012 967 1016
rect 971 1012 972 1016
rect 966 1011 972 1012
rect 1038 1016 1044 1017
rect 1038 1012 1039 1016
rect 1043 1012 1044 1016
rect 1155 1015 1156 1019
rect 1160 1018 1161 1019
rect 1174 1019 1180 1020
rect 1174 1018 1175 1019
rect 1160 1016 1175 1018
rect 1160 1015 1161 1016
rect 1155 1014 1161 1015
rect 1174 1015 1175 1016
rect 1179 1015 1180 1019
rect 1174 1014 1180 1015
rect 1186 1019 1192 1020
rect 1186 1015 1187 1019
rect 1191 1018 1192 1019
rect 1227 1019 1233 1020
rect 1227 1018 1228 1019
rect 1191 1016 1228 1018
rect 1191 1015 1192 1016
rect 1186 1014 1192 1015
rect 1227 1015 1228 1016
rect 1232 1015 1233 1019
rect 1227 1014 1233 1015
rect 1258 1019 1264 1020
rect 1258 1015 1259 1019
rect 1263 1018 1264 1019
rect 1299 1019 1305 1020
rect 1299 1018 1300 1019
rect 1263 1016 1300 1018
rect 1263 1015 1264 1016
rect 1258 1014 1264 1015
rect 1299 1015 1300 1016
rect 1304 1015 1305 1019
rect 1299 1014 1305 1015
rect 1330 1019 1336 1020
rect 1330 1015 1331 1019
rect 1335 1018 1336 1019
rect 1379 1019 1385 1020
rect 1379 1018 1380 1019
rect 1335 1016 1380 1018
rect 1335 1015 1336 1016
rect 1330 1014 1336 1015
rect 1379 1015 1380 1016
rect 1384 1015 1385 1019
rect 1379 1014 1385 1015
rect 1459 1019 1465 1020
rect 1459 1015 1460 1019
rect 1464 1018 1465 1019
rect 1526 1019 1532 1020
rect 1526 1018 1527 1019
rect 1464 1016 1527 1018
rect 1464 1015 1465 1016
rect 1459 1014 1465 1015
rect 1526 1015 1527 1016
rect 1531 1015 1532 1019
rect 1526 1014 1532 1015
rect 1534 1019 1545 1020
rect 1534 1015 1535 1019
rect 1539 1015 1540 1019
rect 1544 1015 1545 1019
rect 1534 1014 1545 1015
rect 1619 1019 1625 1020
rect 1619 1015 1620 1019
rect 1624 1018 1625 1019
rect 1650 1019 1656 1020
rect 1624 1016 1646 1018
rect 1624 1015 1625 1016
rect 1619 1014 1625 1015
rect 1038 1011 1044 1012
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 1094 1008 1100 1009
rect 1094 1004 1095 1008
rect 1099 1004 1100 1008
rect 110 1003 116 1004
rect 247 1003 256 1004
rect 247 999 248 1003
rect 255 999 256 1003
rect 247 998 256 999
rect 295 1003 301 1004
rect 295 999 296 1003
rect 300 1002 301 1003
rect 303 1003 309 1004
rect 303 1002 304 1003
rect 300 1000 304 1002
rect 300 999 301 1000
rect 295 998 301 999
rect 303 999 304 1000
rect 308 999 309 1003
rect 303 998 309 999
rect 359 1003 365 1004
rect 359 999 360 1003
rect 364 1002 365 1003
rect 378 1003 384 1004
rect 378 1002 379 1003
rect 364 1000 379 1002
rect 364 999 365 1000
rect 359 998 365 999
rect 378 999 379 1000
rect 383 999 384 1003
rect 378 998 384 999
rect 422 1003 428 1004
rect 422 999 423 1003
rect 427 1002 428 1003
rect 431 1003 437 1004
rect 431 1002 432 1003
rect 427 1000 432 1002
rect 427 999 428 1000
rect 422 998 428 999
rect 431 999 432 1000
rect 436 999 437 1003
rect 431 998 437 999
rect 503 1003 509 1004
rect 503 999 504 1003
rect 508 1002 509 1003
rect 518 1003 524 1004
rect 518 1002 519 1003
rect 508 1000 519 1002
rect 508 999 509 1000
rect 503 998 509 999
rect 518 999 519 1000
rect 523 999 524 1003
rect 518 998 524 999
rect 546 1003 552 1004
rect 546 999 547 1003
rect 551 1002 552 1003
rect 583 1003 589 1004
rect 583 1002 584 1003
rect 551 1000 584 1002
rect 551 999 552 1000
rect 546 998 552 999
rect 583 999 584 1000
rect 588 999 589 1003
rect 583 998 589 999
rect 618 1003 624 1004
rect 618 999 619 1003
rect 623 1002 624 1003
rect 655 1003 661 1004
rect 655 1002 656 1003
rect 623 1000 656 1002
rect 623 999 624 1000
rect 618 998 624 999
rect 655 999 656 1000
rect 660 999 661 1003
rect 655 998 661 999
rect 727 1003 736 1004
rect 727 999 728 1003
rect 735 999 736 1003
rect 727 998 736 999
rect 799 1003 808 1004
rect 799 999 800 1003
rect 807 999 808 1003
rect 799 998 808 999
rect 863 1003 872 1004
rect 863 999 864 1003
rect 871 999 872 1003
rect 863 998 872 999
rect 926 1003 933 1004
rect 926 999 927 1003
rect 932 999 933 1003
rect 926 998 933 999
rect 991 1003 1000 1004
rect 991 999 992 1003
rect 999 999 1000 1003
rect 991 998 1000 999
rect 1054 1003 1060 1004
rect 1054 999 1055 1003
rect 1059 1002 1060 1003
rect 1063 1003 1069 1004
rect 1094 1003 1100 1004
rect 1158 1008 1164 1009
rect 1158 1004 1159 1008
rect 1163 1004 1164 1008
rect 1158 1003 1164 1004
rect 1230 1008 1236 1009
rect 1230 1004 1231 1008
rect 1235 1004 1236 1008
rect 1230 1003 1236 1004
rect 1302 1008 1308 1009
rect 1302 1004 1303 1008
rect 1307 1004 1308 1008
rect 1302 1003 1308 1004
rect 1382 1008 1388 1009
rect 1382 1004 1383 1008
rect 1387 1004 1388 1008
rect 1382 1003 1388 1004
rect 1462 1008 1468 1009
rect 1462 1004 1463 1008
rect 1467 1004 1468 1008
rect 1462 1003 1468 1004
rect 1542 1008 1548 1009
rect 1542 1004 1543 1008
rect 1547 1004 1548 1008
rect 1542 1003 1548 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1063 1002 1064 1003
rect 1059 1000 1064 1002
rect 1059 999 1060 1000
rect 1054 998 1060 999
rect 1063 999 1064 1000
rect 1068 999 1069 1003
rect 1644 1002 1646 1016
rect 1650 1015 1651 1019
rect 1655 1018 1656 1019
rect 1691 1019 1697 1020
rect 1691 1018 1692 1019
rect 1655 1016 1692 1018
rect 1655 1015 1656 1016
rect 1650 1014 1656 1015
rect 1691 1015 1692 1016
rect 1696 1015 1697 1019
rect 1691 1014 1697 1015
rect 1722 1019 1728 1020
rect 1722 1015 1723 1019
rect 1727 1018 1728 1019
rect 1755 1019 1761 1020
rect 1755 1018 1756 1019
rect 1727 1016 1756 1018
rect 1727 1015 1728 1016
rect 1722 1014 1728 1015
rect 1755 1015 1756 1016
rect 1760 1015 1761 1019
rect 1755 1014 1761 1015
rect 1814 1019 1825 1020
rect 1814 1015 1815 1019
rect 1819 1015 1820 1019
rect 1824 1015 1825 1019
rect 1814 1014 1825 1015
rect 1866 1019 1872 1020
rect 1866 1015 1867 1019
rect 1871 1018 1872 1019
rect 1883 1019 1889 1020
rect 1883 1018 1884 1019
rect 1871 1016 1884 1018
rect 1871 1015 1872 1016
rect 1866 1014 1872 1015
rect 1883 1015 1884 1016
rect 1888 1015 1889 1019
rect 1883 1014 1889 1015
rect 1914 1019 1920 1020
rect 1914 1015 1915 1019
rect 1919 1018 1920 1019
rect 1947 1019 1953 1020
rect 1947 1018 1948 1019
rect 1919 1016 1948 1018
rect 1919 1015 1920 1016
rect 1914 1014 1920 1015
rect 1947 1015 1948 1016
rect 1952 1015 1953 1019
rect 1947 1014 1953 1015
rect 1694 1008 1700 1009
rect 1694 1004 1695 1008
rect 1699 1004 1700 1008
rect 1694 1003 1700 1004
rect 1758 1008 1764 1009
rect 1758 1004 1759 1008
rect 1763 1004 1764 1008
rect 1758 1003 1764 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1886 1008 1892 1009
rect 1822 1003 1828 1004
rect 1840 1004 1883 1006
rect 1063 998 1069 999
rect 1134 1000 1140 1001
rect 1644 1000 1690 1002
rect 1134 996 1135 1000
rect 1139 996 1140 1000
rect 1688 998 1690 1000
rect 1712 1000 1754 1002
rect 1712 998 1714 1000
rect 1688 996 1714 998
rect 1752 998 1754 1000
rect 1772 1000 1810 1002
rect 1772 998 1774 1000
rect 1752 996 1774 998
rect 1808 998 1810 1000
rect 1840 998 1842 1004
rect 1808 996 1842 998
rect 1866 999 1872 1000
rect 1134 995 1140 996
rect 1183 995 1192 996
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 1094 991 1100 992
rect 110 986 116 987
rect 222 988 228 989
rect 222 984 223 988
rect 227 984 228 988
rect 222 983 228 984
rect 270 988 276 989
rect 270 984 271 988
rect 275 984 276 988
rect 270 983 276 984
rect 334 988 340 989
rect 334 984 335 988
rect 339 984 340 988
rect 334 983 340 984
rect 406 988 412 989
rect 406 984 407 988
rect 411 984 412 988
rect 406 983 412 984
rect 478 988 484 989
rect 478 984 479 988
rect 483 984 484 988
rect 478 983 484 984
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 630 988 636 989
rect 630 984 631 988
rect 635 984 636 988
rect 630 983 636 984
rect 702 988 708 989
rect 702 984 703 988
rect 707 984 708 988
rect 702 983 708 984
rect 774 988 780 989
rect 774 984 775 988
rect 779 984 780 988
rect 774 983 780 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 902 988 908 989
rect 902 984 903 988
rect 907 984 908 988
rect 902 983 908 984
rect 966 988 972 989
rect 966 984 967 988
rect 971 984 972 988
rect 966 983 972 984
rect 1038 988 1044 989
rect 1038 984 1039 988
rect 1043 984 1044 988
rect 1094 987 1095 991
rect 1099 987 1100 991
rect 1183 991 1184 995
rect 1191 991 1192 995
rect 1183 990 1192 991
rect 1255 995 1264 996
rect 1255 991 1256 995
rect 1263 991 1264 995
rect 1255 990 1264 991
rect 1327 995 1336 996
rect 1327 991 1328 995
rect 1335 991 1336 995
rect 1327 990 1336 991
rect 1338 995 1344 996
rect 1338 991 1339 995
rect 1343 994 1344 995
rect 1407 995 1413 996
rect 1407 994 1408 995
rect 1343 992 1408 994
rect 1343 991 1344 992
rect 1338 990 1344 991
rect 1407 991 1408 992
rect 1412 991 1413 995
rect 1407 990 1413 991
rect 1486 995 1493 996
rect 1486 991 1487 995
rect 1492 991 1493 995
rect 1486 990 1493 991
rect 1526 995 1532 996
rect 1526 991 1527 995
rect 1531 994 1532 995
rect 1567 995 1573 996
rect 1567 994 1568 995
rect 1531 992 1568 994
rect 1531 991 1532 992
rect 1526 990 1532 991
rect 1567 991 1568 992
rect 1572 991 1573 995
rect 1567 990 1573 991
rect 1647 995 1656 996
rect 1647 991 1648 995
rect 1655 991 1656 995
rect 1647 990 1656 991
rect 1719 995 1728 996
rect 1719 991 1720 995
rect 1727 991 1728 995
rect 1719 990 1728 991
rect 1783 995 1792 996
rect 1783 991 1784 995
rect 1791 991 1792 995
rect 1783 990 1792 991
rect 1847 995 1853 996
rect 1847 991 1848 995
rect 1852 994 1853 995
rect 1866 995 1867 999
rect 1871 995 1872 999
rect 1881 998 1883 1004
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 1904 1000 1926 1002
rect 1904 998 1906 1000
rect 1881 996 1906 998
rect 1866 994 1872 995
rect 1911 995 1920 996
rect 1852 992 1870 994
rect 1852 991 1853 992
rect 1847 990 1853 991
rect 1911 991 1912 995
rect 1919 991 1920 995
rect 1924 994 1926 1000
rect 2118 1000 2124 1001
rect 2118 996 2119 1000
rect 2123 996 2124 1000
rect 1975 995 1981 996
rect 2118 995 2124 996
rect 1975 994 1976 995
rect 1924 992 1976 994
rect 1911 990 1920 991
rect 1975 991 1976 992
rect 1980 991 1981 995
rect 1975 990 1981 991
rect 1094 986 1100 987
rect 1038 983 1044 984
rect 1134 983 1140 984
rect 1134 979 1135 983
rect 1139 979 1140 983
rect 2118 983 2124 984
rect 1134 978 1140 979
rect 1158 980 1164 981
rect 1158 976 1159 980
rect 1163 976 1164 980
rect 1158 975 1164 976
rect 1230 980 1236 981
rect 1230 976 1231 980
rect 1235 976 1236 980
rect 1230 975 1236 976
rect 1302 980 1308 981
rect 1302 976 1303 980
rect 1307 976 1308 980
rect 1302 975 1308 976
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1462 980 1468 981
rect 1462 976 1463 980
rect 1467 976 1468 980
rect 1462 975 1468 976
rect 1542 980 1548 981
rect 1542 976 1543 980
rect 1547 976 1548 980
rect 1542 975 1548 976
rect 1622 980 1628 981
rect 1622 976 1623 980
rect 1627 976 1628 980
rect 1622 975 1628 976
rect 1694 980 1700 981
rect 1694 976 1695 980
rect 1699 976 1700 980
rect 1694 975 1700 976
rect 1758 980 1764 981
rect 1758 976 1759 980
rect 1763 976 1764 980
rect 1758 975 1764 976
rect 1822 980 1828 981
rect 1822 976 1823 980
rect 1827 976 1828 980
rect 1822 975 1828 976
rect 1886 980 1892 981
rect 1886 976 1887 980
rect 1891 976 1892 980
rect 1886 975 1892 976
rect 1950 980 1956 981
rect 1950 976 1951 980
rect 1955 976 1956 980
rect 2118 979 2119 983
rect 2123 979 2124 983
rect 2118 978 2124 979
rect 1950 975 1956 976
rect 150 972 156 973
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 150 968 151 972
rect 155 968 156 972
rect 150 967 156 968
rect 214 972 220 973
rect 214 968 215 972
rect 219 968 220 972
rect 214 967 220 968
rect 286 972 292 973
rect 286 968 287 972
rect 291 968 292 972
rect 286 967 292 968
rect 366 972 372 973
rect 366 968 367 972
rect 371 968 372 972
rect 366 967 372 968
rect 446 972 452 973
rect 446 968 447 972
rect 451 968 452 972
rect 446 967 452 968
rect 526 972 532 973
rect 526 968 527 972
rect 531 968 532 972
rect 526 967 532 968
rect 598 972 604 973
rect 598 968 599 972
rect 603 968 604 972
rect 598 967 604 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 798 972 804 973
rect 798 968 799 972
rect 803 968 804 972
rect 798 967 804 968
rect 862 972 868 973
rect 862 968 863 972
rect 867 968 868 972
rect 862 967 868 968
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 990 972 996 973
rect 990 968 991 972
rect 995 968 996 972
rect 990 967 996 968
rect 1046 972 1052 973
rect 1046 968 1047 972
rect 1051 968 1052 972
rect 1046 967 1052 968
rect 1094 969 1100 970
rect 110 964 116 965
rect 1094 965 1095 969
rect 1099 965 1100 969
rect 1238 968 1244 969
rect 1094 964 1100 965
rect 1134 965 1140 966
rect 238 963 244 964
rect 238 959 239 963
rect 243 962 244 963
rect 710 963 716 964
rect 243 960 370 962
rect 243 959 244 960
rect 238 958 244 959
rect 175 955 181 956
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 175 951 176 955
rect 180 954 181 955
rect 206 955 212 956
rect 206 954 207 955
rect 180 952 207 954
rect 180 951 181 952
rect 175 950 181 951
rect 206 951 207 952
rect 211 951 212 955
rect 206 950 212 951
rect 239 955 245 956
rect 239 951 240 955
rect 244 954 245 955
rect 278 955 284 956
rect 278 954 279 955
rect 244 952 279 954
rect 244 951 245 952
rect 239 950 245 951
rect 278 951 279 952
rect 283 951 284 955
rect 278 950 284 951
rect 311 955 317 956
rect 311 951 312 955
rect 316 954 317 955
rect 358 955 364 956
rect 358 954 359 955
rect 316 952 359 954
rect 316 951 317 952
rect 311 950 317 951
rect 358 951 359 952
rect 363 951 364 955
rect 368 954 370 960
rect 710 959 711 963
rect 715 962 716 963
rect 715 960 930 962
rect 1134 961 1135 965
rect 1139 961 1140 965
rect 1238 964 1239 968
rect 1243 964 1244 968
rect 1238 963 1244 964
rect 1302 968 1308 969
rect 1302 964 1303 968
rect 1307 964 1308 968
rect 1302 963 1308 964
rect 1374 968 1380 969
rect 1374 964 1375 968
rect 1379 964 1380 968
rect 1374 963 1380 964
rect 1438 968 1444 969
rect 1438 964 1439 968
rect 1443 964 1444 968
rect 1438 963 1444 964
rect 1510 968 1516 969
rect 1510 964 1511 968
rect 1515 964 1516 968
rect 1510 963 1516 964
rect 1582 968 1588 969
rect 1582 964 1583 968
rect 1587 964 1588 968
rect 1582 963 1588 964
rect 1654 968 1660 969
rect 1654 964 1655 968
rect 1659 964 1660 968
rect 1654 963 1660 964
rect 1726 968 1732 969
rect 1726 964 1727 968
rect 1731 964 1732 968
rect 1726 963 1732 964
rect 1798 968 1804 969
rect 1798 964 1799 968
rect 1803 964 1804 968
rect 1798 963 1804 964
rect 1870 968 1876 969
rect 1870 964 1871 968
rect 1875 964 1876 968
rect 1870 963 1876 964
rect 1942 968 1948 969
rect 1942 964 1943 968
rect 1947 964 1948 968
rect 1942 963 1948 964
rect 2014 968 2020 969
rect 2014 964 2015 968
rect 2019 964 2020 968
rect 2014 963 2020 964
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2070 963 2076 964
rect 2118 965 2124 966
rect 1134 960 1140 961
rect 2118 961 2119 965
rect 2123 961 2124 965
rect 2118 960 2124 961
rect 715 959 716 960
rect 710 958 716 959
rect 391 955 397 956
rect 391 954 392 955
rect 368 952 392 954
rect 358 950 364 951
rect 391 951 392 952
rect 396 951 397 955
rect 391 950 397 951
rect 470 955 477 956
rect 470 951 471 955
rect 476 951 477 955
rect 470 950 477 951
rect 482 955 488 956
rect 482 951 483 955
rect 487 954 488 955
rect 551 955 557 956
rect 551 954 552 955
rect 487 952 552 954
rect 487 951 488 952
rect 482 950 488 951
rect 551 951 552 952
rect 556 951 557 955
rect 551 950 557 951
rect 623 955 629 956
rect 623 951 624 955
rect 628 954 629 955
rect 662 955 668 956
rect 662 954 663 955
rect 628 952 663 954
rect 628 951 629 952
rect 623 950 629 951
rect 662 951 663 952
rect 667 951 668 955
rect 662 950 668 951
rect 695 955 701 956
rect 695 951 696 955
rect 700 954 701 955
rect 726 955 732 956
rect 726 954 727 955
rect 700 952 727 954
rect 700 951 701 952
rect 695 950 701 951
rect 726 951 727 952
rect 731 951 732 955
rect 726 950 732 951
rect 759 955 765 956
rect 759 951 760 955
rect 764 954 765 955
rect 790 955 796 956
rect 790 954 791 955
rect 764 952 791 954
rect 764 951 765 952
rect 759 950 765 951
rect 790 951 791 952
rect 795 951 796 955
rect 790 950 796 951
rect 823 955 829 956
rect 823 951 824 955
rect 828 954 829 955
rect 854 955 860 956
rect 854 954 855 955
rect 828 952 855 954
rect 828 951 829 952
rect 823 950 829 951
rect 854 951 855 952
rect 859 951 860 955
rect 854 950 860 951
rect 887 955 893 956
rect 887 951 888 955
rect 892 954 893 955
rect 918 955 924 956
rect 918 954 919 955
rect 892 952 919 954
rect 892 951 893 952
rect 887 950 893 951
rect 918 951 919 952
rect 923 951 924 955
rect 928 954 930 960
rect 1610 959 1616 960
rect 951 955 957 956
rect 951 954 952 955
rect 928 952 952 954
rect 918 950 924 951
rect 951 951 952 952
rect 956 951 957 955
rect 951 950 957 951
rect 998 955 1004 956
rect 998 951 999 955
rect 1003 954 1004 955
rect 1015 955 1021 956
rect 1015 954 1016 955
rect 1003 952 1016 954
rect 1003 951 1004 952
rect 998 950 1004 951
rect 1015 951 1016 952
rect 1020 951 1021 955
rect 1015 950 1021 951
rect 1026 955 1032 956
rect 1026 951 1027 955
rect 1031 954 1032 955
rect 1071 955 1077 956
rect 1071 954 1072 955
rect 1031 952 1072 954
rect 1031 951 1032 952
rect 1026 950 1032 951
rect 1071 951 1072 952
rect 1076 951 1077 955
rect 1610 955 1611 959
rect 1615 958 1616 959
rect 1615 956 1874 958
rect 1615 955 1616 956
rect 1610 954 1616 955
rect 1071 950 1077 951
rect 1094 952 1100 953
rect 110 947 116 948
rect 1094 948 1095 952
rect 1099 948 1100 952
rect 1263 951 1269 952
rect 1094 947 1100 948
rect 1134 948 1140 949
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 214 944 220 945
rect 214 940 215 944
rect 219 940 220 944
rect 214 939 220 940
rect 286 944 292 945
rect 286 940 287 944
rect 291 940 292 944
rect 286 939 292 940
rect 366 944 372 945
rect 366 940 367 944
rect 371 940 372 944
rect 366 939 372 940
rect 446 944 452 945
rect 446 940 447 944
rect 451 940 452 944
rect 446 939 452 940
rect 526 944 532 945
rect 526 940 527 944
rect 531 940 532 944
rect 526 939 532 940
rect 598 944 604 945
rect 598 940 599 944
rect 603 940 604 944
rect 598 939 604 940
rect 670 944 676 945
rect 670 940 671 944
rect 675 940 676 944
rect 670 939 676 940
rect 734 944 740 945
rect 734 940 735 944
rect 739 940 740 944
rect 734 939 740 940
rect 798 944 804 945
rect 798 940 799 944
rect 803 940 804 944
rect 798 939 804 940
rect 862 944 868 945
rect 862 940 863 944
rect 867 940 868 944
rect 862 939 868 940
rect 926 944 932 945
rect 926 940 927 944
rect 931 940 932 944
rect 926 939 932 940
rect 990 944 996 945
rect 990 940 991 944
rect 995 940 996 944
rect 990 939 996 940
rect 1046 944 1052 945
rect 1046 940 1047 944
rect 1051 940 1052 944
rect 1134 944 1135 948
rect 1139 944 1140 948
rect 1263 947 1264 951
rect 1268 950 1269 951
rect 1294 951 1300 952
rect 1294 950 1295 951
rect 1268 948 1295 950
rect 1268 947 1269 948
rect 1263 946 1269 947
rect 1294 947 1295 948
rect 1299 947 1300 951
rect 1294 946 1300 947
rect 1327 951 1333 952
rect 1327 947 1328 951
rect 1332 950 1333 951
rect 1366 951 1372 952
rect 1366 950 1367 951
rect 1332 948 1367 950
rect 1332 947 1333 948
rect 1327 946 1333 947
rect 1366 947 1367 948
rect 1371 947 1372 951
rect 1366 946 1372 947
rect 1382 951 1388 952
rect 1382 947 1383 951
rect 1387 950 1388 951
rect 1399 951 1405 952
rect 1399 950 1400 951
rect 1387 948 1400 950
rect 1387 947 1388 948
rect 1382 946 1388 947
rect 1399 947 1400 948
rect 1404 947 1405 951
rect 1399 946 1405 947
rect 1463 951 1469 952
rect 1463 947 1464 951
rect 1468 950 1469 951
rect 1502 951 1508 952
rect 1502 950 1503 951
rect 1468 948 1503 950
rect 1468 947 1469 948
rect 1463 946 1469 947
rect 1502 947 1503 948
rect 1507 947 1508 951
rect 1502 946 1508 947
rect 1534 951 1541 952
rect 1534 947 1535 951
rect 1540 947 1541 951
rect 1534 946 1541 947
rect 1607 951 1613 952
rect 1607 947 1608 951
rect 1612 950 1613 951
rect 1646 951 1652 952
rect 1646 950 1647 951
rect 1612 948 1647 950
rect 1612 947 1613 948
rect 1607 946 1613 947
rect 1646 947 1647 948
rect 1651 947 1652 951
rect 1646 946 1652 947
rect 1679 951 1685 952
rect 1679 947 1680 951
rect 1684 950 1685 951
rect 1718 951 1724 952
rect 1718 950 1719 951
rect 1684 948 1719 950
rect 1684 947 1685 948
rect 1679 946 1685 947
rect 1718 947 1719 948
rect 1723 947 1724 951
rect 1718 946 1724 947
rect 1751 951 1757 952
rect 1751 947 1752 951
rect 1756 950 1757 951
rect 1778 951 1784 952
rect 1778 950 1779 951
rect 1756 948 1779 950
rect 1756 947 1757 948
rect 1751 946 1757 947
rect 1778 947 1779 948
rect 1783 947 1784 951
rect 1778 946 1784 947
rect 1823 951 1829 952
rect 1823 947 1824 951
rect 1828 950 1829 951
rect 1862 951 1868 952
rect 1862 950 1863 951
rect 1828 948 1863 950
rect 1828 947 1829 948
rect 1823 946 1829 947
rect 1862 947 1863 948
rect 1867 947 1868 951
rect 1872 950 1874 956
rect 1895 951 1901 952
rect 1895 950 1896 951
rect 1872 948 1896 950
rect 1862 946 1868 947
rect 1895 947 1896 948
rect 1900 947 1901 951
rect 1895 946 1901 947
rect 1967 951 1973 952
rect 1967 947 1968 951
rect 1972 950 1973 951
rect 1990 951 1996 952
rect 1972 948 1986 950
rect 1972 947 1973 948
rect 1967 946 1973 947
rect 1134 943 1140 944
rect 1984 942 1986 948
rect 1990 947 1991 951
rect 1995 950 1996 951
rect 2039 951 2045 952
rect 2039 950 2040 951
rect 1995 948 2040 950
rect 1995 947 1996 948
rect 1990 946 1996 947
rect 2039 947 2040 948
rect 2044 947 2045 951
rect 2039 946 2045 947
rect 2047 951 2053 952
rect 2047 947 2048 951
rect 2052 950 2053 951
rect 2095 951 2101 952
rect 2095 950 2096 951
rect 2052 948 2096 950
rect 2052 947 2053 948
rect 2047 946 2053 947
rect 2095 947 2096 948
rect 2100 947 2101 951
rect 2095 946 2101 947
rect 2118 948 2124 949
rect 2118 944 2119 948
rect 2123 944 2124 948
rect 2006 943 2012 944
rect 2118 943 2124 944
rect 2006 942 2007 943
rect 1046 939 1052 940
rect 1238 940 1244 941
rect 1238 936 1239 940
rect 1243 936 1244 940
rect 1238 935 1244 936
rect 1302 940 1308 941
rect 1302 936 1303 940
rect 1307 936 1308 940
rect 1302 935 1308 936
rect 1374 940 1380 941
rect 1374 936 1375 940
rect 1379 936 1380 940
rect 1374 935 1380 936
rect 1438 940 1444 941
rect 1438 936 1439 940
rect 1443 936 1444 940
rect 1438 935 1444 936
rect 1510 940 1516 941
rect 1510 936 1511 940
rect 1515 936 1516 940
rect 1510 935 1516 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1654 940 1660 941
rect 1654 936 1655 940
rect 1659 936 1660 940
rect 1654 935 1660 936
rect 1726 940 1732 941
rect 1726 936 1727 940
rect 1731 936 1732 940
rect 1726 935 1732 936
rect 1798 940 1804 941
rect 1798 936 1799 940
rect 1803 936 1804 940
rect 1798 935 1804 936
rect 1870 940 1876 941
rect 1870 936 1871 940
rect 1875 936 1876 940
rect 1870 935 1876 936
rect 1942 940 1948 941
rect 1984 940 2007 942
rect 1942 936 1943 940
rect 1947 936 1948 940
rect 2006 939 2007 940
rect 2011 939 2012 943
rect 2006 938 2012 939
rect 2014 940 2020 941
rect 1942 935 1948 936
rect 2014 936 2015 940
rect 2019 936 2020 940
rect 2014 935 2020 936
rect 2070 940 2076 941
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 147 931 153 932
rect 147 927 148 931
rect 152 930 153 931
rect 158 931 164 932
rect 158 930 159 931
rect 152 928 159 930
rect 152 927 153 928
rect 147 926 153 927
rect 158 927 159 928
rect 163 927 164 931
rect 158 926 164 927
rect 206 931 217 932
rect 206 927 207 931
rect 211 927 212 931
rect 216 927 217 931
rect 206 926 217 927
rect 278 931 289 932
rect 278 927 279 931
rect 283 927 284 931
rect 288 927 289 931
rect 278 926 289 927
rect 358 931 369 932
rect 358 927 359 931
rect 363 927 364 931
rect 368 927 369 931
rect 358 926 369 927
rect 443 931 449 932
rect 443 927 444 931
rect 448 930 449 931
rect 482 931 488 932
rect 482 930 483 931
rect 448 928 483 930
rect 448 927 449 928
rect 443 926 449 927
rect 482 927 483 928
rect 487 927 488 931
rect 482 926 488 927
rect 518 931 529 932
rect 518 927 519 931
rect 523 927 524 931
rect 528 927 529 931
rect 518 926 529 927
rect 595 931 601 932
rect 595 927 596 931
rect 600 930 601 931
rect 654 931 660 932
rect 654 930 655 931
rect 600 928 655 930
rect 600 927 601 928
rect 595 926 601 927
rect 654 927 655 928
rect 659 927 660 931
rect 654 926 660 927
rect 662 931 673 932
rect 662 927 663 931
rect 667 927 668 931
rect 672 927 673 931
rect 662 926 673 927
rect 726 931 737 932
rect 726 927 727 931
rect 731 927 732 931
rect 736 927 737 931
rect 726 926 737 927
rect 790 931 801 932
rect 790 927 791 931
rect 795 927 796 931
rect 800 927 801 931
rect 790 926 801 927
rect 854 931 865 932
rect 854 927 855 931
rect 859 927 860 931
rect 864 927 865 931
rect 854 926 865 927
rect 918 931 929 932
rect 918 927 919 931
rect 923 927 924 931
rect 928 927 929 931
rect 918 926 929 927
rect 987 931 993 932
rect 987 927 988 931
rect 992 930 993 931
rect 1026 931 1032 932
rect 1026 930 1027 931
rect 992 928 1027 930
rect 992 927 993 928
rect 987 926 993 927
rect 1026 927 1027 928
rect 1031 927 1032 931
rect 1026 926 1032 927
rect 1043 931 1049 932
rect 1043 927 1044 931
rect 1048 930 1049 931
rect 1054 931 1060 932
rect 1054 930 1055 931
rect 1048 928 1055 930
rect 1048 927 1049 928
rect 1043 926 1049 927
rect 1054 927 1055 928
rect 1059 927 1060 931
rect 1054 926 1060 927
rect 1235 927 1241 928
rect 1235 923 1236 927
rect 1240 926 1241 927
rect 1294 927 1305 928
rect 1240 924 1290 926
rect 1240 923 1241 924
rect 1235 922 1241 923
rect 131 919 137 920
rect 131 915 132 919
rect 136 918 137 919
rect 170 919 176 920
rect 170 918 171 919
rect 136 916 171 918
rect 136 915 137 916
rect 131 914 137 915
rect 170 915 171 916
rect 175 915 176 919
rect 170 914 176 915
rect 179 919 185 920
rect 179 915 180 919
rect 184 918 185 919
rect 242 919 248 920
rect 242 918 243 919
rect 184 916 243 918
rect 184 915 185 916
rect 179 914 185 915
rect 242 915 243 916
rect 247 915 248 919
rect 242 914 248 915
rect 251 919 257 920
rect 251 915 252 919
rect 256 918 257 919
rect 302 919 308 920
rect 302 918 303 919
rect 256 916 303 918
rect 256 915 257 916
rect 251 914 257 915
rect 302 915 303 916
rect 307 915 308 919
rect 302 914 308 915
rect 323 919 329 920
rect 323 915 324 919
rect 328 918 329 919
rect 386 919 392 920
rect 386 918 387 919
rect 328 916 387 918
rect 328 915 329 916
rect 323 914 329 915
rect 386 915 387 916
rect 391 915 392 919
rect 386 914 392 915
rect 395 919 401 920
rect 395 915 396 919
rect 400 918 401 919
rect 447 919 453 920
rect 447 918 448 919
rect 400 916 448 918
rect 400 915 401 916
rect 395 914 401 915
rect 447 915 448 916
rect 452 915 453 919
rect 447 914 453 915
rect 459 919 465 920
rect 459 915 460 919
rect 464 918 465 919
rect 470 919 476 920
rect 470 918 471 919
rect 464 916 471 918
rect 464 915 465 916
rect 459 914 465 915
rect 470 915 471 916
rect 475 915 476 919
rect 470 914 476 915
rect 523 919 529 920
rect 523 915 524 919
rect 528 918 529 919
rect 546 919 552 920
rect 546 918 547 919
rect 528 916 547 918
rect 528 915 529 916
rect 523 914 529 915
rect 546 915 547 916
rect 551 915 552 919
rect 546 914 552 915
rect 554 919 560 920
rect 554 915 555 919
rect 559 918 560 919
rect 595 919 601 920
rect 595 918 596 919
rect 559 916 596 918
rect 559 915 560 916
rect 554 914 560 915
rect 595 915 596 916
rect 600 915 601 919
rect 595 914 601 915
rect 626 919 632 920
rect 626 915 627 919
rect 631 918 632 919
rect 667 919 673 920
rect 667 918 668 919
rect 631 916 668 918
rect 631 915 632 916
rect 626 914 632 915
rect 667 915 668 916
rect 672 915 673 919
rect 667 914 673 915
rect 698 919 704 920
rect 698 915 699 919
rect 703 918 704 919
rect 739 919 745 920
rect 739 918 740 919
rect 703 916 740 918
rect 703 915 704 916
rect 698 914 704 915
rect 739 915 740 916
rect 744 915 745 919
rect 739 914 745 915
rect 770 919 776 920
rect 770 915 771 919
rect 775 918 776 919
rect 811 919 817 920
rect 811 918 812 919
rect 775 916 812 918
rect 775 915 776 916
rect 770 914 776 915
rect 811 915 812 916
rect 816 915 817 919
rect 811 914 817 915
rect 842 919 848 920
rect 842 915 843 919
rect 847 918 848 919
rect 891 919 897 920
rect 891 918 892 919
rect 847 916 892 918
rect 847 915 848 916
rect 842 914 848 915
rect 891 915 892 916
rect 896 915 897 919
rect 891 914 897 915
rect 979 919 985 920
rect 979 915 980 919
rect 984 918 985 919
rect 998 919 1004 920
rect 998 918 999 919
rect 984 916 999 918
rect 984 915 985 916
rect 979 914 985 915
rect 998 915 999 916
rect 1003 915 1004 919
rect 998 914 1004 915
rect 1026 919 1032 920
rect 1026 915 1027 919
rect 1031 918 1032 919
rect 1043 919 1049 920
rect 1043 918 1044 919
rect 1031 916 1044 918
rect 1031 915 1032 916
rect 1026 914 1032 915
rect 1043 915 1044 916
rect 1048 915 1049 919
rect 1288 918 1290 924
rect 1294 923 1295 927
rect 1299 923 1300 927
rect 1304 923 1305 927
rect 1294 922 1305 923
rect 1366 927 1377 928
rect 1366 923 1367 927
rect 1371 923 1372 927
rect 1376 923 1377 927
rect 1366 922 1377 923
rect 1435 927 1441 928
rect 1435 923 1436 927
rect 1440 926 1441 927
rect 1446 927 1452 928
rect 1446 926 1447 927
rect 1440 924 1447 926
rect 1440 923 1441 924
rect 1435 922 1441 923
rect 1446 923 1447 924
rect 1451 923 1452 927
rect 1446 922 1452 923
rect 1502 927 1513 928
rect 1502 923 1503 927
rect 1507 923 1508 927
rect 1512 923 1513 927
rect 1502 922 1513 923
rect 1579 927 1585 928
rect 1579 923 1580 927
rect 1584 926 1585 927
rect 1610 927 1616 928
rect 1610 926 1611 927
rect 1584 924 1611 926
rect 1584 923 1585 924
rect 1579 922 1585 923
rect 1610 923 1611 924
rect 1615 923 1616 927
rect 1610 922 1616 923
rect 1646 927 1657 928
rect 1646 923 1647 927
rect 1651 923 1652 927
rect 1656 923 1657 927
rect 1646 922 1657 923
rect 1718 927 1729 928
rect 1718 923 1719 927
rect 1723 923 1724 927
rect 1728 923 1729 927
rect 1718 922 1729 923
rect 1786 927 1792 928
rect 1786 923 1787 927
rect 1791 926 1792 927
rect 1795 927 1801 928
rect 1795 926 1796 927
rect 1791 924 1796 926
rect 1791 923 1792 924
rect 1786 922 1792 923
rect 1795 923 1796 924
rect 1800 923 1801 927
rect 1795 922 1801 923
rect 1862 927 1873 928
rect 1862 923 1863 927
rect 1867 923 1868 927
rect 1872 923 1873 927
rect 1862 922 1873 923
rect 1939 927 1945 928
rect 1939 923 1940 927
rect 1944 926 1945 927
rect 1990 927 1996 928
rect 1990 926 1991 927
rect 1944 924 1991 926
rect 1944 923 1945 924
rect 1939 922 1945 923
rect 1990 923 1991 924
rect 1995 923 1996 927
rect 1990 922 1996 923
rect 2011 927 2017 928
rect 2011 923 2012 927
rect 2016 926 2017 927
rect 2047 927 2053 928
rect 2047 926 2048 927
rect 2016 924 2048 926
rect 2016 923 2017 924
rect 2011 922 2017 923
rect 2047 923 2048 924
rect 2052 923 2053 927
rect 2047 922 2053 923
rect 2067 927 2073 928
rect 2067 923 2068 927
rect 2072 926 2073 927
rect 2086 927 2092 928
rect 2086 926 2087 927
rect 2072 924 2087 926
rect 2072 923 2073 924
rect 2067 922 2073 923
rect 2086 923 2087 924
rect 2091 923 2092 927
rect 2086 922 2092 923
rect 1338 919 1344 920
rect 1338 918 1339 919
rect 1288 916 1339 918
rect 1043 914 1049 915
rect 1338 915 1339 916
rect 1343 915 1344 919
rect 1338 914 1344 915
rect 1283 911 1289 912
rect 134 908 140 909
rect 134 904 135 908
rect 139 904 140 908
rect 134 903 140 904
rect 182 908 188 909
rect 182 904 183 908
rect 187 904 188 908
rect 182 903 188 904
rect 254 908 260 909
rect 254 904 255 908
rect 259 904 260 908
rect 254 903 260 904
rect 326 908 332 909
rect 326 904 327 908
rect 331 904 332 908
rect 326 903 332 904
rect 398 908 404 909
rect 398 904 399 908
rect 403 904 404 908
rect 398 903 404 904
rect 462 908 468 909
rect 462 904 463 908
rect 467 904 468 908
rect 462 903 468 904
rect 526 908 532 909
rect 526 904 527 908
rect 531 904 532 908
rect 526 903 532 904
rect 598 908 604 909
rect 598 904 599 908
rect 603 904 604 908
rect 598 903 604 904
rect 670 908 676 909
rect 670 904 671 908
rect 675 904 676 908
rect 670 903 676 904
rect 742 908 748 909
rect 742 904 743 908
rect 747 904 748 908
rect 742 903 748 904
rect 814 908 820 909
rect 814 904 815 908
rect 819 904 820 908
rect 814 903 820 904
rect 894 908 900 909
rect 894 904 895 908
rect 899 904 900 908
rect 894 903 900 904
rect 982 908 988 909
rect 982 904 983 908
rect 987 904 988 908
rect 982 903 988 904
rect 1046 908 1052 909
rect 1046 904 1047 908
rect 1051 904 1052 908
rect 1283 907 1284 911
rect 1288 910 1289 911
rect 1323 911 1329 912
rect 1288 908 1318 910
rect 1288 907 1289 908
rect 1283 906 1289 907
rect 1046 903 1052 904
rect 110 900 116 901
rect 110 896 111 900
rect 115 896 116 900
rect 1094 900 1100 901
rect 1094 896 1095 900
rect 1099 896 1100 900
rect 110 895 116 896
rect 158 895 165 896
rect 158 891 159 895
rect 164 891 165 895
rect 158 890 165 891
rect 170 895 176 896
rect 170 891 171 895
rect 175 894 176 895
rect 207 895 213 896
rect 207 894 208 895
rect 175 892 208 894
rect 175 891 176 892
rect 170 890 176 891
rect 207 891 208 892
rect 212 891 213 895
rect 207 890 213 891
rect 242 895 248 896
rect 242 891 243 895
rect 247 894 248 895
rect 279 895 285 896
rect 279 894 280 895
rect 247 892 280 894
rect 247 891 248 892
rect 242 890 248 891
rect 279 891 280 892
rect 284 891 285 895
rect 279 890 285 891
rect 350 895 357 896
rect 350 891 351 895
rect 356 891 357 895
rect 350 890 357 891
rect 386 895 392 896
rect 386 891 387 895
rect 391 894 392 895
rect 423 895 429 896
rect 423 894 424 895
rect 391 892 424 894
rect 391 891 392 892
rect 386 890 392 891
rect 423 891 424 892
rect 428 891 429 895
rect 423 890 429 891
rect 447 895 453 896
rect 447 891 448 895
rect 452 894 453 895
rect 487 895 493 896
rect 487 894 488 895
rect 452 892 488 894
rect 452 891 453 892
rect 447 890 453 891
rect 487 891 488 892
rect 492 891 493 895
rect 487 890 493 891
rect 551 895 560 896
rect 551 891 552 895
rect 559 891 560 895
rect 551 890 560 891
rect 623 895 632 896
rect 623 891 624 895
rect 631 891 632 895
rect 623 890 632 891
rect 695 895 704 896
rect 695 891 696 895
rect 703 891 704 895
rect 695 890 704 891
rect 767 895 776 896
rect 767 891 768 895
rect 775 891 776 895
rect 767 890 776 891
rect 839 895 848 896
rect 839 891 840 895
rect 847 891 848 895
rect 839 890 848 891
rect 918 895 925 896
rect 918 891 919 895
rect 924 891 925 895
rect 918 890 925 891
rect 1007 895 1013 896
rect 1007 891 1008 895
rect 1012 894 1013 895
rect 1026 895 1032 896
rect 1026 894 1027 895
rect 1012 892 1027 894
rect 1012 891 1013 892
rect 1007 890 1013 891
rect 1026 891 1027 892
rect 1031 891 1032 895
rect 1026 890 1032 891
rect 1071 895 1077 896
rect 1071 891 1072 895
rect 1076 894 1077 895
rect 1086 895 1092 896
rect 1094 895 1100 896
rect 1286 900 1292 901
rect 1286 896 1287 900
rect 1291 896 1292 900
rect 1286 895 1292 896
rect 1086 894 1087 895
rect 1076 892 1087 894
rect 1076 891 1077 892
rect 1071 890 1077 891
rect 1086 891 1087 892
rect 1091 891 1092 895
rect 1316 894 1318 908
rect 1323 907 1324 911
rect 1328 910 1329 911
rect 1362 911 1368 912
rect 1362 910 1363 911
rect 1328 908 1363 910
rect 1328 907 1329 908
rect 1323 906 1329 907
rect 1362 907 1363 908
rect 1367 907 1368 911
rect 1362 906 1368 907
rect 1371 911 1377 912
rect 1371 907 1372 911
rect 1376 910 1377 911
rect 1382 911 1388 912
rect 1382 910 1383 911
rect 1376 908 1383 910
rect 1376 907 1377 908
rect 1371 906 1377 907
rect 1382 907 1383 908
rect 1387 907 1388 911
rect 1382 906 1388 907
rect 1419 911 1425 912
rect 1419 907 1420 911
rect 1424 910 1425 911
rect 1466 911 1472 912
rect 1466 910 1467 911
rect 1424 908 1467 910
rect 1424 907 1425 908
rect 1419 906 1425 907
rect 1466 907 1467 908
rect 1471 907 1472 911
rect 1466 906 1472 907
rect 1475 911 1481 912
rect 1475 907 1476 911
rect 1480 910 1481 911
rect 1494 911 1500 912
rect 1494 910 1495 911
rect 1480 908 1495 910
rect 1480 907 1481 908
rect 1475 906 1481 907
rect 1494 907 1495 908
rect 1499 907 1500 911
rect 1494 906 1500 907
rect 1547 911 1553 912
rect 1547 907 1548 911
rect 1552 910 1553 911
rect 1610 911 1616 912
rect 1610 910 1611 911
rect 1552 908 1611 910
rect 1552 907 1553 908
rect 1547 906 1553 907
rect 1610 907 1611 908
rect 1615 907 1616 911
rect 1610 906 1616 907
rect 1619 911 1625 912
rect 1619 907 1620 911
rect 1624 910 1625 911
rect 1690 911 1696 912
rect 1690 910 1691 911
rect 1624 908 1691 910
rect 1624 907 1625 908
rect 1619 906 1625 907
rect 1690 907 1691 908
rect 1695 907 1696 911
rect 1690 906 1696 907
rect 1699 911 1705 912
rect 1699 907 1700 911
rect 1704 910 1705 911
rect 1770 911 1776 912
rect 1770 910 1771 911
rect 1704 908 1771 910
rect 1704 907 1705 908
rect 1699 906 1705 907
rect 1770 907 1771 908
rect 1775 907 1776 911
rect 1770 906 1776 907
rect 1778 911 1784 912
rect 1778 907 1779 911
rect 1783 910 1784 911
rect 1787 911 1793 912
rect 1787 910 1788 911
rect 1783 908 1788 910
rect 1783 907 1784 908
rect 1778 906 1784 907
rect 1787 907 1788 908
rect 1792 907 1793 911
rect 1875 911 1881 912
rect 1875 908 1876 911
rect 1787 906 1793 907
rect 1870 907 1876 908
rect 1880 907 1881 911
rect 1870 903 1871 907
rect 1875 906 1881 907
rect 1906 911 1912 912
rect 1906 907 1907 911
rect 1911 910 1912 911
rect 1963 911 1969 912
rect 1963 910 1964 911
rect 1911 908 1964 910
rect 1911 907 1912 908
rect 1906 906 1912 907
rect 1963 907 1964 908
rect 1968 907 1969 911
rect 1963 906 1969 907
rect 1994 911 2000 912
rect 1994 907 1995 911
rect 1999 910 2000 911
rect 2059 911 2065 912
rect 2059 910 2060 911
rect 1999 908 2060 910
rect 1999 907 2000 908
rect 1994 906 2000 907
rect 2059 907 2060 908
rect 2064 907 2065 911
rect 2059 906 2065 907
rect 1875 904 1879 906
rect 1875 903 1876 904
rect 1870 902 1876 903
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1374 900 1380 901
rect 1374 896 1375 900
rect 1379 896 1380 900
rect 1374 895 1380 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1478 900 1484 901
rect 1478 896 1479 900
rect 1483 896 1484 900
rect 1478 895 1484 896
rect 1550 900 1556 901
rect 1550 896 1551 900
rect 1555 896 1556 900
rect 1550 895 1556 896
rect 1622 900 1628 901
rect 1622 896 1623 900
rect 1627 896 1628 900
rect 1622 895 1628 896
rect 1702 900 1708 901
rect 1702 896 1703 900
rect 1707 896 1708 900
rect 1702 895 1708 896
rect 1790 900 1796 901
rect 1790 896 1791 900
rect 1795 896 1796 900
rect 1790 895 1796 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1966 900 1972 901
rect 1966 896 1967 900
rect 1971 896 1972 900
rect 1966 895 1972 896
rect 2062 900 2068 901
rect 2062 896 2063 900
rect 2067 896 2068 900
rect 2062 895 2068 896
rect 1086 890 1092 891
rect 1134 892 1140 893
rect 1316 892 1322 894
rect 1134 888 1135 892
rect 1139 888 1140 892
rect 1134 887 1140 888
rect 1206 887 1212 888
rect 110 883 116 884
rect 110 879 111 883
rect 115 879 116 883
rect 1094 883 1100 884
rect 110 878 116 879
rect 134 880 140 881
rect 134 876 135 880
rect 139 876 140 880
rect 134 875 140 876
rect 182 880 188 881
rect 182 876 183 880
rect 187 876 188 880
rect 182 875 188 876
rect 254 880 260 881
rect 254 876 255 880
rect 259 876 260 880
rect 254 875 260 876
rect 326 880 332 881
rect 326 876 327 880
rect 331 876 332 880
rect 326 875 332 876
rect 398 880 404 881
rect 398 876 399 880
rect 403 876 404 880
rect 398 875 404 876
rect 462 880 468 881
rect 462 876 463 880
rect 467 876 468 880
rect 462 875 468 876
rect 526 880 532 881
rect 526 876 527 880
rect 531 876 532 880
rect 526 875 532 876
rect 598 880 604 881
rect 598 876 599 880
rect 603 876 604 880
rect 598 875 604 876
rect 670 880 676 881
rect 670 876 671 880
rect 675 876 676 880
rect 670 875 676 876
rect 742 880 748 881
rect 742 876 743 880
rect 747 876 748 880
rect 742 875 748 876
rect 814 880 820 881
rect 814 876 815 880
rect 819 876 820 880
rect 814 875 820 876
rect 894 880 900 881
rect 894 876 895 880
rect 899 876 900 880
rect 894 875 900 876
rect 982 880 988 881
rect 982 876 983 880
rect 987 876 988 880
rect 982 875 988 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1094 879 1095 883
rect 1099 879 1100 883
rect 1206 883 1207 887
rect 1211 886 1212 887
rect 1311 887 1317 888
rect 1311 886 1312 887
rect 1211 884 1312 886
rect 1211 883 1212 884
rect 1206 882 1212 883
rect 1311 883 1312 884
rect 1316 883 1317 887
rect 1320 886 1322 892
rect 2118 892 2124 893
rect 2118 888 2119 892
rect 2123 888 2124 892
rect 1351 887 1357 888
rect 1351 886 1352 887
rect 1320 884 1352 886
rect 1311 882 1317 883
rect 1351 883 1352 884
rect 1356 883 1357 887
rect 1351 882 1357 883
rect 1362 887 1368 888
rect 1362 883 1363 887
rect 1367 886 1368 887
rect 1399 887 1405 888
rect 1399 886 1400 887
rect 1367 884 1400 886
rect 1367 883 1368 884
rect 1362 882 1368 883
rect 1399 883 1400 884
rect 1404 883 1405 887
rect 1399 882 1405 883
rect 1446 887 1453 888
rect 1446 883 1447 887
rect 1452 883 1453 887
rect 1446 882 1453 883
rect 1466 887 1472 888
rect 1466 883 1467 887
rect 1471 886 1472 887
rect 1503 887 1509 888
rect 1503 886 1504 887
rect 1471 884 1504 886
rect 1471 883 1472 884
rect 1466 882 1472 883
rect 1503 883 1504 884
rect 1508 883 1509 887
rect 1503 882 1509 883
rect 1558 887 1564 888
rect 1558 883 1559 887
rect 1563 886 1564 887
rect 1575 887 1581 888
rect 1575 886 1576 887
rect 1563 884 1576 886
rect 1563 883 1564 884
rect 1558 882 1564 883
rect 1575 883 1576 884
rect 1580 883 1581 887
rect 1575 882 1581 883
rect 1610 887 1616 888
rect 1610 883 1611 887
rect 1615 886 1616 887
rect 1647 887 1653 888
rect 1647 886 1648 887
rect 1615 884 1648 886
rect 1615 883 1616 884
rect 1610 882 1616 883
rect 1647 883 1648 884
rect 1652 883 1653 887
rect 1647 882 1653 883
rect 1690 887 1696 888
rect 1690 883 1691 887
rect 1695 886 1696 887
rect 1727 887 1733 888
rect 1727 886 1728 887
rect 1695 884 1728 886
rect 1695 883 1696 884
rect 1690 882 1696 883
rect 1727 883 1728 884
rect 1732 883 1733 887
rect 1727 882 1733 883
rect 1770 887 1776 888
rect 1770 883 1771 887
rect 1775 886 1776 887
rect 1815 887 1821 888
rect 1815 886 1816 887
rect 1775 884 1816 886
rect 1775 883 1776 884
rect 1770 882 1776 883
rect 1815 883 1816 884
rect 1820 883 1821 887
rect 1815 882 1821 883
rect 1903 887 1912 888
rect 1903 883 1904 887
rect 1911 883 1912 887
rect 1903 882 1912 883
rect 1991 887 2000 888
rect 1991 883 1992 887
rect 1999 883 2000 887
rect 1991 882 2000 883
rect 2086 887 2093 888
rect 2118 887 2124 888
rect 2086 883 2087 887
rect 2092 883 2093 887
rect 2086 882 2093 883
rect 1094 878 1100 879
rect 1046 875 1052 876
rect 1134 875 1140 876
rect 654 871 660 872
rect 654 867 655 871
rect 659 870 660 871
rect 918 871 924 872
rect 918 870 919 871
rect 659 868 919 870
rect 659 867 660 868
rect 654 866 660 867
rect 918 867 919 868
rect 923 867 924 871
rect 1134 871 1135 875
rect 1139 871 1140 875
rect 2118 875 2124 876
rect 1134 870 1140 871
rect 1286 872 1292 873
rect 1286 868 1287 872
rect 1291 868 1292 872
rect 1286 867 1292 868
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 1326 867 1332 868
rect 1374 872 1380 873
rect 1374 868 1375 872
rect 1379 868 1380 872
rect 1374 867 1380 868
rect 1422 872 1428 873
rect 1422 868 1423 872
rect 1427 868 1428 872
rect 1422 867 1428 868
rect 1478 872 1484 873
rect 1478 868 1479 872
rect 1483 868 1484 872
rect 1478 867 1484 868
rect 1550 872 1556 873
rect 1550 868 1551 872
rect 1555 868 1556 872
rect 1550 867 1556 868
rect 1622 872 1628 873
rect 1622 868 1623 872
rect 1627 868 1628 872
rect 1622 867 1628 868
rect 1702 872 1708 873
rect 1702 868 1703 872
rect 1707 868 1708 872
rect 1702 867 1708 868
rect 1790 872 1796 873
rect 1790 868 1791 872
rect 1795 868 1796 872
rect 1790 867 1796 868
rect 1878 872 1884 873
rect 1878 868 1879 872
rect 1883 868 1884 872
rect 1878 867 1884 868
rect 1966 872 1972 873
rect 1966 868 1967 872
rect 1971 868 1972 872
rect 1966 867 1972 868
rect 2062 872 2068 873
rect 2062 868 2063 872
rect 2067 868 2068 872
rect 2118 871 2119 875
rect 2123 871 2124 875
rect 2118 870 2124 871
rect 2062 867 2068 868
rect 918 866 924 867
rect 134 864 140 865
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 134 860 135 864
rect 139 860 140 864
rect 134 859 140 860
rect 174 864 180 865
rect 174 860 175 864
rect 179 860 180 864
rect 174 859 180 860
rect 214 864 220 865
rect 214 860 215 864
rect 219 860 220 864
rect 214 859 220 860
rect 278 864 284 865
rect 278 860 279 864
rect 283 860 284 864
rect 278 859 284 860
rect 342 864 348 865
rect 342 860 343 864
rect 347 860 348 864
rect 342 859 348 860
rect 398 864 404 865
rect 398 860 399 864
rect 403 860 404 864
rect 398 859 404 860
rect 462 864 468 865
rect 462 860 463 864
rect 467 860 468 864
rect 462 859 468 860
rect 534 864 540 865
rect 534 860 535 864
rect 539 860 540 864
rect 534 859 540 860
rect 614 864 620 865
rect 614 860 615 864
rect 619 860 620 864
rect 614 859 620 860
rect 710 864 716 865
rect 710 860 711 864
rect 715 860 716 864
rect 710 859 716 860
rect 822 864 828 865
rect 822 860 823 864
rect 827 860 828 864
rect 822 859 828 860
rect 942 864 948 865
rect 942 860 943 864
rect 947 860 948 864
rect 942 859 948 860
rect 1046 864 1052 865
rect 1046 860 1047 864
rect 1051 860 1052 864
rect 1046 859 1052 860
rect 1094 861 1100 862
rect 110 856 116 857
rect 1094 857 1095 861
rect 1099 857 1100 861
rect 1158 860 1164 861
rect 1094 856 1100 857
rect 1134 857 1140 858
rect 902 855 908 856
rect 902 851 903 855
rect 907 854 908 855
rect 907 852 987 854
rect 1134 853 1135 857
rect 1139 853 1140 857
rect 1158 856 1159 860
rect 1163 856 1164 860
rect 1158 855 1164 856
rect 1198 860 1204 861
rect 1198 856 1199 860
rect 1203 856 1204 860
rect 1198 855 1204 856
rect 1262 860 1268 861
rect 1262 856 1263 860
rect 1267 856 1268 860
rect 1262 855 1268 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1398 860 1404 861
rect 1398 856 1399 860
rect 1403 856 1404 860
rect 1398 855 1404 856
rect 1470 860 1476 861
rect 1470 856 1471 860
rect 1475 856 1476 860
rect 1470 855 1476 856
rect 1542 860 1548 861
rect 1542 856 1543 860
rect 1547 856 1548 860
rect 1542 855 1548 856
rect 1622 860 1628 861
rect 1622 856 1623 860
rect 1627 856 1628 860
rect 1622 855 1628 856
rect 1702 860 1708 861
rect 1702 856 1703 860
rect 1707 856 1708 860
rect 1702 855 1708 856
rect 1774 860 1780 861
rect 1774 856 1775 860
rect 1779 856 1780 860
rect 1774 855 1780 856
rect 1854 860 1860 861
rect 1854 856 1855 860
rect 1859 856 1860 860
rect 1854 855 1860 856
rect 1934 860 1940 861
rect 1934 856 1935 860
rect 1939 856 1940 860
rect 1934 855 1940 856
rect 2014 860 2020 861
rect 2014 856 2015 860
rect 2019 856 2020 860
rect 2014 855 2020 856
rect 2070 860 2076 861
rect 2070 856 2071 860
rect 2075 856 2076 860
rect 2070 855 2076 856
rect 2118 857 2124 858
rect 1134 852 1140 853
rect 2118 853 2119 857
rect 2123 853 2124 857
rect 2118 852 2124 853
rect 907 851 908 852
rect 902 850 908 851
rect 159 847 168 848
rect 110 844 116 845
rect 110 840 111 844
rect 115 840 116 844
rect 159 843 160 847
rect 167 843 168 847
rect 159 842 168 843
rect 199 847 208 848
rect 199 843 200 847
rect 207 843 208 847
rect 199 842 208 843
rect 239 847 245 848
rect 239 843 240 847
rect 244 846 245 847
rect 270 847 276 848
rect 270 846 271 847
rect 244 844 271 846
rect 244 843 245 844
rect 239 842 245 843
rect 270 843 271 844
rect 275 843 276 847
rect 270 842 276 843
rect 302 847 309 848
rect 302 843 303 847
rect 308 843 309 847
rect 302 842 309 843
rect 367 847 373 848
rect 367 843 368 847
rect 372 846 373 847
rect 383 847 389 848
rect 383 846 384 847
rect 372 844 384 846
rect 372 843 373 844
rect 367 842 373 843
rect 383 843 384 844
rect 388 843 389 847
rect 383 842 389 843
rect 406 847 412 848
rect 406 843 407 847
rect 411 846 412 847
rect 423 847 429 848
rect 423 846 424 847
rect 411 844 424 846
rect 411 843 412 844
rect 406 842 412 843
rect 423 843 424 844
rect 428 843 429 847
rect 423 842 429 843
rect 470 847 476 848
rect 470 843 471 847
rect 475 846 476 847
rect 487 847 493 848
rect 487 846 488 847
rect 475 844 488 846
rect 475 843 476 844
rect 470 842 476 843
rect 487 843 488 844
rect 492 843 493 847
rect 487 842 493 843
rect 559 847 565 848
rect 559 843 560 847
rect 564 846 565 847
rect 606 847 612 848
rect 606 846 607 847
rect 564 844 607 846
rect 564 843 565 844
rect 559 842 565 843
rect 606 843 607 844
rect 611 843 612 847
rect 606 842 612 843
rect 639 847 645 848
rect 639 843 640 847
rect 644 846 645 847
rect 702 847 708 848
rect 702 846 703 847
rect 644 844 703 846
rect 644 843 645 844
rect 639 842 645 843
rect 702 843 703 844
rect 707 843 708 847
rect 702 842 708 843
rect 735 847 741 848
rect 735 843 736 847
rect 740 846 741 847
rect 807 847 813 848
rect 807 846 808 847
rect 740 844 808 846
rect 740 843 741 844
rect 735 842 741 843
rect 807 843 808 844
rect 812 843 813 847
rect 807 842 813 843
rect 846 847 853 848
rect 846 843 847 847
rect 852 843 853 847
rect 846 842 853 843
rect 858 847 864 848
rect 858 843 859 847
rect 863 846 864 847
rect 967 847 973 848
rect 967 846 968 847
rect 863 844 968 846
rect 863 843 864 844
rect 858 842 864 843
rect 967 843 968 844
rect 972 843 973 847
rect 985 846 987 852
rect 1071 847 1077 848
rect 1071 846 1072 847
rect 985 844 1072 846
rect 967 842 973 843
rect 1071 843 1072 844
rect 1076 843 1077 847
rect 1071 842 1077 843
rect 1094 844 1100 845
rect 110 839 116 840
rect 1094 840 1095 844
rect 1099 840 1100 844
rect 1142 843 1148 844
rect 1094 839 1100 840
rect 1134 840 1140 841
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 174 836 180 837
rect 174 832 175 836
rect 179 832 180 836
rect 174 831 180 832
rect 214 836 220 837
rect 214 832 215 836
rect 219 832 220 836
rect 214 831 220 832
rect 278 836 284 837
rect 278 832 279 836
rect 283 832 284 836
rect 278 831 284 832
rect 342 836 348 837
rect 342 832 343 836
rect 347 832 348 836
rect 342 831 348 832
rect 398 836 404 837
rect 398 832 399 836
rect 403 832 404 836
rect 398 831 404 832
rect 462 836 468 837
rect 462 832 463 836
rect 467 832 468 836
rect 462 831 468 832
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 614 836 620 837
rect 614 832 615 836
rect 619 832 620 836
rect 614 831 620 832
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 822 836 828 837
rect 822 832 823 836
rect 827 832 828 836
rect 822 831 828 832
rect 942 836 948 837
rect 942 832 943 836
rect 947 832 948 836
rect 942 831 948 832
rect 1046 836 1052 837
rect 1046 832 1047 836
rect 1051 832 1052 836
rect 1134 836 1135 840
rect 1139 836 1140 840
rect 1142 839 1143 843
rect 1147 842 1148 843
rect 1183 843 1189 844
rect 1183 842 1184 843
rect 1147 840 1184 842
rect 1147 839 1148 840
rect 1142 838 1148 839
rect 1183 839 1184 840
rect 1188 839 1189 843
rect 1183 838 1189 839
rect 1223 843 1229 844
rect 1223 839 1224 843
rect 1228 842 1229 843
rect 1254 843 1260 844
rect 1254 842 1255 843
rect 1228 840 1255 842
rect 1228 839 1229 840
rect 1223 838 1229 839
rect 1254 839 1255 840
rect 1259 839 1260 843
rect 1254 838 1260 839
rect 1287 843 1293 844
rect 1287 839 1288 843
rect 1292 842 1293 843
rect 1318 843 1324 844
rect 1318 842 1319 843
rect 1292 840 1319 842
rect 1292 839 1293 840
rect 1287 838 1293 839
rect 1318 839 1319 840
rect 1323 839 1324 843
rect 1318 838 1324 839
rect 1351 843 1357 844
rect 1351 839 1352 843
rect 1356 842 1357 843
rect 1390 843 1396 844
rect 1390 842 1391 843
rect 1356 840 1391 842
rect 1356 839 1357 840
rect 1351 838 1357 839
rect 1390 839 1391 840
rect 1395 839 1396 843
rect 1390 838 1396 839
rect 1423 843 1429 844
rect 1423 839 1424 843
rect 1428 842 1429 843
rect 1462 843 1468 844
rect 1462 842 1463 843
rect 1428 840 1463 842
rect 1428 839 1429 840
rect 1423 838 1429 839
rect 1462 839 1463 840
rect 1467 839 1468 843
rect 1462 838 1468 839
rect 1494 843 1501 844
rect 1494 839 1495 843
rect 1500 839 1501 843
rect 1494 838 1501 839
rect 1567 843 1573 844
rect 1567 839 1568 843
rect 1572 842 1573 843
rect 1614 843 1620 844
rect 1614 842 1615 843
rect 1572 840 1615 842
rect 1572 839 1573 840
rect 1567 838 1573 839
rect 1614 839 1615 840
rect 1619 839 1620 843
rect 1614 838 1620 839
rect 1647 843 1653 844
rect 1647 839 1648 843
rect 1652 842 1653 843
rect 1694 843 1700 844
rect 1694 842 1695 843
rect 1652 840 1695 842
rect 1652 839 1653 840
rect 1647 838 1653 839
rect 1694 839 1695 840
rect 1699 839 1700 843
rect 1694 838 1700 839
rect 1727 843 1733 844
rect 1727 839 1728 843
rect 1732 842 1733 843
rect 1766 843 1772 844
rect 1766 842 1767 843
rect 1732 840 1767 842
rect 1732 839 1733 840
rect 1727 838 1733 839
rect 1766 839 1767 840
rect 1771 839 1772 843
rect 1766 838 1772 839
rect 1782 843 1788 844
rect 1782 839 1783 843
rect 1787 842 1788 843
rect 1799 843 1805 844
rect 1799 842 1800 843
rect 1787 840 1800 842
rect 1787 839 1788 840
rect 1782 838 1788 839
rect 1799 839 1800 840
rect 1804 839 1805 843
rect 1799 838 1805 839
rect 1870 843 1876 844
rect 1870 839 1871 843
rect 1875 842 1876 843
rect 1879 843 1885 844
rect 1879 842 1880 843
rect 1875 840 1880 842
rect 1875 839 1876 840
rect 1870 838 1876 839
rect 1879 839 1880 840
rect 1884 839 1885 843
rect 1879 838 1885 839
rect 1898 843 1904 844
rect 1898 839 1899 843
rect 1903 842 1904 843
rect 1959 843 1965 844
rect 1959 842 1960 843
rect 1903 840 1960 842
rect 1903 839 1904 840
rect 1898 838 1904 839
rect 1959 839 1960 840
rect 1964 839 1965 843
rect 1959 838 1965 839
rect 2039 843 2045 844
rect 2039 839 2040 843
rect 2044 842 2045 843
rect 2062 843 2068 844
rect 2062 842 2063 843
rect 2044 840 2063 842
rect 2044 839 2045 840
rect 2039 838 2045 839
rect 2062 839 2063 840
rect 2067 839 2068 843
rect 2062 838 2068 839
rect 2078 843 2084 844
rect 2078 839 2079 843
rect 2083 842 2084 843
rect 2095 843 2101 844
rect 2095 842 2096 843
rect 2083 840 2096 842
rect 2083 839 2084 840
rect 2078 838 2084 839
rect 2095 839 2096 840
rect 2100 839 2101 843
rect 2095 838 2101 839
rect 2118 840 2124 841
rect 1134 835 1140 836
rect 2118 836 2119 840
rect 2123 836 2124 840
rect 2118 835 2124 836
rect 1158 832 1164 833
rect 1046 831 1052 832
rect 1086 831 1092 832
rect 1086 827 1087 831
rect 1091 830 1092 831
rect 1091 828 1154 830
rect 1091 827 1092 828
rect 1086 826 1092 827
rect 131 823 137 824
rect 131 819 132 823
rect 136 822 137 823
rect 154 823 160 824
rect 154 822 155 823
rect 136 820 155 822
rect 136 819 137 820
rect 131 818 137 819
rect 154 819 155 820
rect 159 819 160 823
rect 154 818 160 819
rect 162 823 168 824
rect 162 819 163 823
rect 167 822 168 823
rect 171 823 177 824
rect 171 822 172 823
rect 167 820 172 822
rect 167 819 168 820
rect 162 818 168 819
rect 171 819 172 820
rect 176 819 177 823
rect 171 818 177 819
rect 202 823 208 824
rect 202 819 203 823
rect 207 822 208 823
rect 211 823 217 824
rect 211 822 212 823
rect 207 820 212 822
rect 207 819 208 820
rect 202 818 208 819
rect 211 819 212 820
rect 216 819 217 823
rect 211 818 217 819
rect 270 823 281 824
rect 270 819 271 823
rect 275 819 276 823
rect 280 819 281 823
rect 270 818 281 819
rect 339 823 345 824
rect 339 819 340 823
rect 344 822 345 823
rect 350 823 356 824
rect 350 822 351 823
rect 344 820 351 822
rect 344 819 345 820
rect 339 818 345 819
rect 350 819 351 820
rect 355 819 356 823
rect 350 818 356 819
rect 383 823 389 824
rect 383 819 384 823
rect 388 822 389 823
rect 395 823 401 824
rect 395 822 396 823
rect 388 820 396 822
rect 388 819 389 820
rect 383 818 389 819
rect 395 819 396 820
rect 400 819 401 823
rect 395 818 401 819
rect 459 823 465 824
rect 459 819 460 823
rect 464 822 465 823
rect 478 823 484 824
rect 478 822 479 823
rect 464 820 479 822
rect 464 819 465 820
rect 459 818 465 819
rect 478 819 479 820
rect 483 819 484 823
rect 478 818 484 819
rect 531 823 537 824
rect 531 819 532 823
rect 536 822 537 823
rect 598 823 604 824
rect 598 822 599 823
rect 536 820 599 822
rect 536 819 537 820
rect 531 818 537 819
rect 598 819 599 820
rect 603 819 604 823
rect 598 818 604 819
rect 606 823 617 824
rect 606 819 607 823
rect 611 819 612 823
rect 616 819 617 823
rect 606 818 617 819
rect 702 823 713 824
rect 702 819 703 823
rect 707 819 708 823
rect 712 819 713 823
rect 702 818 713 819
rect 807 823 813 824
rect 807 819 808 823
rect 812 822 813 823
rect 819 823 825 824
rect 819 822 820 823
rect 812 820 820 822
rect 812 819 813 820
rect 807 818 813 819
rect 819 819 820 820
rect 824 819 825 823
rect 819 818 825 819
rect 842 823 848 824
rect 842 819 843 823
rect 847 822 848 823
rect 939 823 945 824
rect 939 822 940 823
rect 847 820 940 822
rect 847 819 848 820
rect 842 818 848 819
rect 939 819 940 820
rect 944 819 945 823
rect 939 818 945 819
rect 1043 823 1049 824
rect 1043 819 1044 823
rect 1048 822 1049 823
rect 1142 823 1148 824
rect 1142 822 1143 823
rect 1048 820 1143 822
rect 1048 819 1049 820
rect 1043 818 1049 819
rect 1142 819 1143 820
rect 1147 819 1148 823
rect 1152 822 1154 828
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1158 827 1164 828
rect 1198 832 1204 833
rect 1198 828 1199 832
rect 1203 828 1204 832
rect 1198 827 1204 828
rect 1262 832 1268 833
rect 1262 828 1263 832
rect 1267 828 1268 832
rect 1262 827 1268 828
rect 1326 832 1332 833
rect 1326 828 1327 832
rect 1331 828 1332 832
rect 1326 827 1332 828
rect 1398 832 1404 833
rect 1398 828 1399 832
rect 1403 828 1404 832
rect 1398 827 1404 828
rect 1470 832 1476 833
rect 1470 828 1471 832
rect 1475 828 1476 832
rect 1470 827 1476 828
rect 1542 832 1548 833
rect 1542 828 1543 832
rect 1547 828 1548 832
rect 1542 827 1548 828
rect 1622 832 1628 833
rect 1622 828 1623 832
rect 1627 828 1628 832
rect 1622 827 1628 828
rect 1702 832 1708 833
rect 1702 828 1703 832
rect 1707 828 1708 832
rect 1702 827 1708 828
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1854 832 1860 833
rect 1854 828 1855 832
rect 1859 828 1860 832
rect 1854 827 1860 828
rect 1934 832 1940 833
rect 1934 828 1935 832
rect 1939 828 1940 832
rect 1934 827 1940 828
rect 2014 832 2020 833
rect 2014 828 2015 832
rect 2019 828 2020 832
rect 2014 827 2020 828
rect 2070 832 2076 833
rect 2070 828 2071 832
rect 2075 828 2076 832
rect 2070 827 2076 828
rect 1152 821 1161 822
rect 1152 820 1156 821
rect 1142 818 1148 819
rect 1155 817 1156 820
rect 1160 817 1161 821
rect 1155 816 1161 817
rect 1195 819 1201 820
rect 1195 815 1196 819
rect 1200 818 1201 819
rect 1206 819 1212 820
rect 1206 818 1207 819
rect 1200 816 1207 818
rect 1200 815 1201 816
rect 1195 814 1201 815
rect 1206 815 1207 816
rect 1211 815 1212 819
rect 1206 814 1212 815
rect 1254 819 1265 820
rect 1254 815 1255 819
rect 1259 815 1260 819
rect 1264 815 1265 819
rect 1254 814 1265 815
rect 1318 819 1329 820
rect 1318 815 1319 819
rect 1323 815 1324 819
rect 1328 815 1329 819
rect 1318 814 1329 815
rect 1390 819 1401 820
rect 1390 815 1391 819
rect 1395 815 1396 819
rect 1400 815 1401 819
rect 1390 814 1401 815
rect 1462 819 1473 820
rect 1462 815 1463 819
rect 1467 815 1468 819
rect 1472 815 1473 819
rect 1462 814 1473 815
rect 1539 819 1545 820
rect 1539 815 1540 819
rect 1544 818 1545 819
rect 1558 819 1564 820
rect 1558 818 1559 819
rect 1544 816 1559 818
rect 1544 815 1545 816
rect 1539 814 1545 815
rect 1558 815 1559 816
rect 1563 815 1564 819
rect 1558 814 1564 815
rect 1614 819 1625 820
rect 1614 815 1615 819
rect 1619 815 1620 819
rect 1624 815 1625 819
rect 1614 814 1625 815
rect 1694 819 1705 820
rect 1694 815 1695 819
rect 1699 815 1700 819
rect 1704 815 1705 819
rect 1694 814 1705 815
rect 1766 819 1777 820
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1776 815 1777 819
rect 1766 814 1777 815
rect 1851 819 1857 820
rect 1851 815 1852 819
rect 1856 818 1857 819
rect 1898 819 1904 820
rect 1898 818 1899 819
rect 1856 816 1899 818
rect 1856 815 1857 816
rect 1851 814 1857 815
rect 1898 815 1899 816
rect 1903 815 1904 819
rect 1898 814 1904 815
rect 1931 819 1937 820
rect 1931 815 1932 819
rect 1936 818 1937 819
rect 1998 819 2004 820
rect 1998 818 1999 819
rect 1936 816 1999 818
rect 1936 815 1937 816
rect 1931 814 1937 815
rect 1998 815 1999 816
rect 2003 815 2004 819
rect 1998 814 2004 815
rect 2006 819 2017 820
rect 2006 815 2007 819
rect 2011 815 2012 819
rect 2016 815 2017 819
rect 2006 814 2017 815
rect 2062 819 2073 820
rect 2062 815 2063 819
rect 2067 815 2068 819
rect 2072 815 2073 819
rect 2062 814 2073 815
rect 131 811 137 812
rect 131 807 132 811
rect 136 810 137 811
rect 162 811 168 812
rect 136 808 158 810
rect 136 807 137 808
rect 131 806 137 807
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 156 794 158 808
rect 162 807 163 811
rect 167 810 168 811
rect 171 811 177 812
rect 171 810 172 811
rect 167 808 172 810
rect 167 807 168 808
rect 162 806 168 807
rect 171 807 172 808
rect 176 807 177 811
rect 171 806 177 807
rect 202 811 208 812
rect 202 807 203 811
rect 207 810 208 811
rect 211 811 217 812
rect 211 810 212 811
rect 207 808 212 810
rect 207 807 208 808
rect 202 806 208 807
rect 211 807 212 808
rect 216 807 217 811
rect 211 806 217 807
rect 275 811 281 812
rect 275 807 276 811
rect 280 810 281 811
rect 322 811 328 812
rect 322 810 323 811
rect 280 808 323 810
rect 280 807 281 808
rect 275 806 281 807
rect 322 807 323 808
rect 327 807 328 811
rect 322 806 328 807
rect 331 811 337 812
rect 331 807 332 811
rect 336 810 337 811
rect 378 811 384 812
rect 378 810 379 811
rect 336 808 379 810
rect 336 807 337 808
rect 331 806 337 807
rect 378 807 379 808
rect 383 807 384 811
rect 378 806 384 807
rect 387 811 393 812
rect 387 807 388 811
rect 392 810 393 811
rect 406 811 412 812
rect 406 810 407 811
rect 392 808 407 810
rect 392 807 393 808
rect 387 806 393 807
rect 406 807 407 808
rect 411 807 412 811
rect 406 806 412 807
rect 451 811 457 812
rect 451 807 452 811
rect 456 810 457 811
rect 470 811 476 812
rect 470 810 471 811
rect 456 808 471 810
rect 456 807 457 808
rect 451 806 457 807
rect 470 807 471 808
rect 475 807 476 811
rect 470 806 476 807
rect 482 811 488 812
rect 482 807 483 811
rect 487 810 488 811
rect 515 811 521 812
rect 515 810 516 811
rect 487 808 516 810
rect 487 807 488 808
rect 482 806 488 807
rect 515 807 516 808
rect 520 807 521 811
rect 515 806 521 807
rect 546 811 552 812
rect 546 807 547 811
rect 551 810 552 811
rect 579 811 585 812
rect 579 810 580 811
rect 551 808 580 810
rect 551 807 552 808
rect 546 806 552 807
rect 579 807 580 808
rect 584 807 585 811
rect 579 806 585 807
rect 615 811 621 812
rect 615 807 616 811
rect 620 810 621 811
rect 651 811 657 812
rect 651 810 652 811
rect 620 808 652 810
rect 620 807 621 808
rect 615 806 621 807
rect 651 807 652 808
rect 656 807 657 811
rect 651 806 657 807
rect 718 811 724 812
rect 718 807 719 811
rect 723 810 724 811
rect 731 811 737 812
rect 731 810 732 811
rect 723 808 732 810
rect 723 807 724 808
rect 718 806 724 807
rect 731 807 732 808
rect 736 807 737 811
rect 731 806 737 807
rect 762 811 768 812
rect 762 807 763 811
rect 767 810 768 811
rect 811 811 817 812
rect 811 810 812 811
rect 767 808 812 810
rect 767 807 768 808
rect 762 806 768 807
rect 811 807 812 808
rect 816 807 817 811
rect 811 806 817 807
rect 891 811 897 812
rect 891 807 892 811
rect 896 810 897 811
rect 902 811 908 812
rect 902 810 903 811
rect 896 808 903 810
rect 896 807 897 808
rect 891 806 897 807
rect 902 807 903 808
rect 907 807 908 811
rect 902 806 908 807
rect 922 811 928 812
rect 922 807 923 811
rect 927 810 928 811
rect 979 811 985 812
rect 979 810 980 811
rect 927 808 980 810
rect 927 807 928 808
rect 922 806 928 807
rect 979 807 980 808
rect 984 807 985 811
rect 979 806 985 807
rect 1010 811 1016 812
rect 1010 807 1011 811
rect 1015 810 1016 811
rect 1043 811 1049 812
rect 1043 810 1044 811
rect 1015 808 1044 810
rect 1015 807 1016 808
rect 1010 806 1016 807
rect 1043 807 1044 808
rect 1048 807 1049 811
rect 1043 806 1049 807
rect 174 800 180 801
rect 174 796 175 800
rect 179 796 180 800
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 174 795 180 796
rect 199 795 205 796
rect 214 795 220 796
rect 278 800 284 801
rect 278 796 279 800
rect 283 796 284 800
rect 278 795 284 796
rect 334 800 340 801
rect 334 796 335 800
rect 339 796 340 800
rect 334 795 340 796
rect 390 800 396 801
rect 390 796 391 800
rect 395 796 396 800
rect 390 795 396 796
rect 454 800 460 801
rect 454 796 455 800
rect 459 796 460 800
rect 454 795 460 796
rect 518 800 524 801
rect 518 796 519 800
rect 523 796 524 800
rect 518 795 524 796
rect 582 800 588 801
rect 582 796 583 800
rect 587 796 588 800
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 582 795 588 796
rect 598 795 604 796
rect 654 795 660 796
rect 734 800 740 801
rect 734 796 735 800
rect 739 796 740 800
rect 734 795 740 796
rect 814 800 820 801
rect 814 796 815 800
rect 819 796 820 800
rect 814 795 820 796
rect 894 800 900 801
rect 894 796 895 800
rect 899 796 900 800
rect 894 795 900 796
rect 982 800 988 801
rect 982 796 983 800
rect 987 796 988 800
rect 982 795 988 796
rect 1046 800 1052 801
rect 1046 796 1047 800
rect 1051 796 1052 800
rect 1155 799 1161 800
rect 1155 798 1156 799
rect 1046 795 1052 796
rect 1088 796 1156 798
rect 199 794 200 795
rect 110 792 116 793
rect 156 792 170 794
rect 110 788 111 792
rect 115 788 116 792
rect 168 790 170 792
rect 193 792 200 794
rect 193 790 195 792
rect 199 791 200 792
rect 204 791 205 795
rect 199 790 205 791
rect 598 791 599 795
rect 603 794 604 795
rect 603 792 618 794
rect 603 791 604 792
rect 598 790 604 791
rect 168 788 195 790
rect 110 787 116 788
rect 154 787 165 788
rect 154 783 155 787
rect 159 783 160 787
rect 164 783 165 787
rect 154 782 165 783
rect 199 787 208 788
rect 199 783 200 787
rect 207 783 208 787
rect 199 782 208 783
rect 215 787 221 788
rect 215 783 216 787
rect 220 786 221 787
rect 239 787 245 788
rect 239 786 240 787
rect 220 784 240 786
rect 220 783 221 784
rect 215 782 221 783
rect 239 783 240 784
rect 244 783 245 787
rect 239 782 245 783
rect 247 787 253 788
rect 247 783 248 787
rect 252 786 253 787
rect 303 787 309 788
rect 303 786 304 787
rect 252 784 304 786
rect 252 783 253 784
rect 247 782 253 783
rect 303 783 304 784
rect 308 783 309 787
rect 303 782 309 783
rect 322 787 328 788
rect 322 783 323 787
rect 327 786 328 787
rect 359 787 365 788
rect 359 786 360 787
rect 327 784 360 786
rect 327 783 328 784
rect 322 782 328 783
rect 359 783 360 784
rect 364 783 365 787
rect 359 782 365 783
rect 378 787 384 788
rect 378 783 379 787
rect 383 786 384 787
rect 415 787 421 788
rect 415 786 416 787
rect 383 784 416 786
rect 383 783 384 784
rect 378 782 384 783
rect 415 783 416 784
rect 420 783 421 787
rect 415 782 421 783
rect 479 787 488 788
rect 479 783 480 787
rect 487 783 488 787
rect 479 782 488 783
rect 543 787 552 788
rect 543 783 544 787
rect 551 783 552 787
rect 543 782 552 783
rect 554 787 560 788
rect 554 783 555 787
rect 559 786 560 787
rect 607 787 613 788
rect 607 786 608 787
rect 559 784 608 786
rect 559 783 560 784
rect 554 782 560 783
rect 607 783 608 784
rect 612 783 613 787
rect 616 786 618 792
rect 679 787 685 788
rect 679 786 680 787
rect 616 784 680 786
rect 607 782 613 783
rect 679 783 680 784
rect 684 783 685 787
rect 679 782 685 783
rect 759 787 768 788
rect 759 783 760 787
rect 767 783 768 787
rect 759 782 768 783
rect 839 787 848 788
rect 839 783 840 787
rect 847 783 848 787
rect 839 782 848 783
rect 919 787 928 788
rect 919 783 920 787
rect 927 783 928 787
rect 919 782 928 783
rect 1007 787 1016 788
rect 1007 783 1008 787
rect 1015 783 1016 787
rect 1007 782 1016 783
rect 1071 787 1077 788
rect 1071 783 1072 787
rect 1076 786 1077 787
rect 1088 786 1090 796
rect 1155 795 1156 796
rect 1160 795 1161 799
rect 1155 794 1161 795
rect 1186 799 1192 800
rect 1186 795 1187 799
rect 1191 798 1192 799
rect 1235 799 1241 800
rect 1235 798 1236 799
rect 1191 796 1236 798
rect 1191 795 1192 796
rect 1186 794 1192 795
rect 1235 795 1236 796
rect 1240 795 1241 799
rect 1235 794 1241 795
rect 1302 799 1308 800
rect 1302 795 1303 799
rect 1307 798 1308 799
rect 1339 799 1345 800
rect 1339 798 1340 799
rect 1307 796 1340 798
rect 1307 795 1308 796
rect 1302 794 1308 795
rect 1339 795 1340 796
rect 1344 795 1345 799
rect 1339 794 1345 795
rect 1443 799 1449 800
rect 1443 795 1444 799
rect 1448 798 1449 799
rect 1535 799 1541 800
rect 1535 798 1536 799
rect 1448 796 1536 798
rect 1448 795 1449 796
rect 1443 794 1449 795
rect 1535 795 1536 796
rect 1540 795 1541 799
rect 1535 794 1541 795
rect 1547 799 1553 800
rect 1547 795 1548 799
rect 1552 798 1553 799
rect 1642 799 1648 800
rect 1642 798 1643 799
rect 1552 796 1643 798
rect 1552 795 1553 796
rect 1547 794 1553 795
rect 1642 795 1643 796
rect 1647 795 1648 799
rect 1642 794 1648 795
rect 1651 799 1657 800
rect 1651 795 1652 799
rect 1656 798 1657 799
rect 1738 799 1744 800
rect 1738 798 1739 799
rect 1656 796 1739 798
rect 1656 795 1657 796
rect 1651 794 1657 795
rect 1738 795 1739 796
rect 1743 795 1744 799
rect 1738 794 1744 795
rect 1747 799 1753 800
rect 1747 795 1748 799
rect 1752 798 1753 799
rect 1782 799 1788 800
rect 1782 798 1783 799
rect 1752 796 1783 798
rect 1752 795 1753 796
rect 1747 794 1753 795
rect 1782 795 1783 796
rect 1787 795 1788 799
rect 1782 794 1788 795
rect 1830 799 1841 800
rect 1830 795 1831 799
rect 1835 795 1836 799
rect 1840 795 1841 799
rect 1830 794 1841 795
rect 1866 799 1872 800
rect 1866 795 1867 799
rect 1871 798 1872 799
rect 1915 799 1921 800
rect 1915 798 1916 799
rect 1871 796 1916 798
rect 1871 795 1872 796
rect 1866 794 1872 795
rect 1915 795 1916 796
rect 1920 795 1921 799
rect 1915 794 1921 795
rect 1946 799 1952 800
rect 1946 795 1947 799
rect 1951 798 1952 799
rect 2003 799 2009 800
rect 2003 798 2004 799
rect 1951 796 2004 798
rect 1951 795 1952 796
rect 1946 794 1952 795
rect 2003 795 2004 796
rect 2008 795 2009 799
rect 2003 794 2009 795
rect 2067 799 2073 800
rect 2067 795 2068 799
rect 2072 798 2073 799
rect 2078 799 2084 800
rect 2078 798 2079 799
rect 2072 796 2079 798
rect 2072 795 2073 796
rect 2067 794 2073 795
rect 2078 795 2079 796
rect 2083 795 2084 799
rect 2078 794 2084 795
rect 1094 792 1100 793
rect 1094 788 1095 792
rect 1099 788 1100 792
rect 1094 787 1100 788
rect 1158 788 1164 789
rect 1076 784 1090 786
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1076 783 1077 784
rect 1158 783 1164 784
rect 1238 788 1244 789
rect 1238 784 1239 788
rect 1243 784 1244 788
rect 1238 783 1244 784
rect 1342 788 1348 789
rect 1342 784 1343 788
rect 1347 784 1348 788
rect 1342 783 1348 784
rect 1446 788 1452 789
rect 1446 784 1447 788
rect 1451 784 1452 788
rect 1446 783 1452 784
rect 1550 788 1556 789
rect 1550 784 1551 788
rect 1555 784 1556 788
rect 1550 783 1556 784
rect 1654 788 1660 789
rect 1654 784 1655 788
rect 1659 784 1660 788
rect 1654 783 1660 784
rect 1750 788 1756 789
rect 1750 784 1751 788
rect 1755 784 1756 788
rect 1750 783 1756 784
rect 1838 788 1844 789
rect 1838 784 1839 788
rect 1843 784 1844 788
rect 1838 783 1844 784
rect 1918 788 1924 789
rect 1918 784 1919 788
rect 1923 784 1924 788
rect 1918 783 1924 784
rect 2006 788 2012 789
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 1071 782 1077 783
rect 1134 780 1140 781
rect 2118 780 2124 781
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 1302 779 1308 780
rect 110 775 116 776
rect 110 771 111 775
rect 115 771 116 775
rect 1094 775 1100 776
rect 1134 775 1140 776
rect 1183 775 1192 776
rect 110 770 116 771
rect 134 772 140 773
rect 134 768 135 772
rect 139 768 140 772
rect 134 767 140 768
rect 174 772 180 773
rect 174 768 175 772
rect 179 768 180 772
rect 174 767 180 768
rect 214 772 220 773
rect 214 768 215 772
rect 219 768 220 772
rect 214 767 220 768
rect 278 772 284 773
rect 278 768 279 772
rect 283 768 284 772
rect 278 767 284 768
rect 334 772 340 773
rect 334 768 335 772
rect 339 768 340 772
rect 334 767 340 768
rect 390 772 396 773
rect 390 768 391 772
rect 395 768 396 772
rect 390 767 396 768
rect 454 772 460 773
rect 454 768 455 772
rect 459 768 460 772
rect 454 767 460 768
rect 518 772 524 773
rect 518 768 519 772
rect 523 768 524 772
rect 518 767 524 768
rect 582 772 588 773
rect 582 768 583 772
rect 587 768 588 772
rect 582 767 588 768
rect 654 772 660 773
rect 654 768 655 772
rect 659 768 660 772
rect 654 767 660 768
rect 734 772 740 773
rect 734 768 735 772
rect 739 768 740 772
rect 734 767 740 768
rect 814 772 820 773
rect 814 768 815 772
rect 819 768 820 772
rect 814 767 820 768
rect 894 772 900 773
rect 894 768 895 772
rect 899 768 900 772
rect 894 767 900 768
rect 982 772 988 773
rect 982 768 983 772
rect 987 768 988 772
rect 982 767 988 768
rect 1046 772 1052 773
rect 1046 768 1047 772
rect 1051 768 1052 772
rect 1094 771 1095 775
rect 1099 771 1100 775
rect 1094 770 1100 771
rect 1183 771 1184 775
rect 1191 771 1192 775
rect 1183 770 1192 771
rect 1263 775 1269 776
rect 1263 771 1264 775
rect 1268 774 1269 775
rect 1302 775 1303 779
rect 1307 775 1308 779
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 1302 774 1308 775
rect 1310 775 1316 776
rect 1268 772 1306 774
rect 1268 771 1269 772
rect 1263 770 1269 771
rect 1310 771 1311 775
rect 1315 774 1316 775
rect 1367 775 1373 776
rect 1367 774 1368 775
rect 1315 772 1368 774
rect 1315 771 1316 772
rect 1310 770 1316 771
rect 1367 771 1368 772
rect 1372 771 1373 775
rect 1367 770 1373 771
rect 1471 775 1477 776
rect 1471 771 1472 775
rect 1476 774 1477 775
rect 1518 775 1524 776
rect 1518 774 1519 775
rect 1476 772 1519 774
rect 1476 771 1477 772
rect 1471 770 1477 771
rect 1518 771 1519 772
rect 1523 771 1524 775
rect 1518 770 1524 771
rect 1535 775 1541 776
rect 1535 771 1536 775
rect 1540 774 1541 775
rect 1575 775 1581 776
rect 1575 774 1576 775
rect 1540 772 1576 774
rect 1540 771 1541 772
rect 1535 770 1541 771
rect 1575 771 1576 772
rect 1580 771 1581 775
rect 1575 770 1581 771
rect 1642 775 1648 776
rect 1642 771 1643 775
rect 1647 774 1648 775
rect 1679 775 1685 776
rect 1679 774 1680 775
rect 1647 772 1680 774
rect 1647 771 1648 772
rect 1642 770 1648 771
rect 1679 771 1680 772
rect 1684 771 1685 775
rect 1679 770 1685 771
rect 1738 775 1744 776
rect 1738 771 1739 775
rect 1743 774 1744 775
rect 1775 775 1781 776
rect 1775 774 1776 775
rect 1743 772 1776 774
rect 1743 771 1744 772
rect 1738 770 1744 771
rect 1775 771 1776 772
rect 1780 771 1781 775
rect 1775 770 1781 771
rect 1863 775 1872 776
rect 1863 771 1864 775
rect 1871 771 1872 775
rect 1863 770 1872 771
rect 1943 775 1952 776
rect 1943 771 1944 775
rect 1951 771 1952 775
rect 1943 770 1952 771
rect 1998 775 2004 776
rect 1998 771 1999 775
rect 2003 774 2004 775
rect 2031 775 2037 776
rect 2031 774 2032 775
rect 2003 772 2032 774
rect 2003 771 2004 772
rect 1998 770 2004 771
rect 2031 771 2032 772
rect 2036 771 2037 775
rect 2031 770 2037 771
rect 2086 775 2092 776
rect 2086 771 2087 775
rect 2091 774 2092 775
rect 2095 775 2101 776
rect 2118 775 2124 776
rect 2095 774 2096 775
rect 2091 772 2096 774
rect 2091 771 2092 772
rect 2086 770 2092 771
rect 2095 771 2096 772
rect 2100 771 2101 775
rect 2095 770 2101 771
rect 1046 767 1052 768
rect 1134 763 1140 764
rect 134 760 140 761
rect 110 757 116 758
rect 110 753 111 757
rect 115 753 116 757
rect 134 756 135 760
rect 139 756 140 760
rect 134 755 140 756
rect 206 760 212 761
rect 206 756 207 760
rect 211 756 212 760
rect 206 755 212 756
rect 294 760 300 761
rect 294 756 295 760
rect 299 756 300 760
rect 294 755 300 756
rect 374 760 380 761
rect 374 756 375 760
rect 379 756 380 760
rect 374 755 380 756
rect 446 760 452 761
rect 446 756 447 760
rect 451 756 452 760
rect 446 755 452 756
rect 518 760 524 761
rect 518 756 519 760
rect 523 756 524 760
rect 518 755 524 756
rect 582 760 588 761
rect 582 756 583 760
rect 587 756 588 760
rect 582 755 588 756
rect 638 760 644 761
rect 638 756 639 760
rect 643 756 644 760
rect 638 755 644 756
rect 686 760 692 761
rect 686 756 687 760
rect 691 756 692 760
rect 686 755 692 756
rect 742 760 748 761
rect 742 756 743 760
rect 747 756 748 760
rect 742 755 748 756
rect 798 760 804 761
rect 798 756 799 760
rect 803 756 804 760
rect 798 755 804 756
rect 854 760 860 761
rect 854 756 855 760
rect 859 756 860 760
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 2118 763 2124 764
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 854 755 860 756
rect 1094 757 1100 758
rect 110 752 116 753
rect 1094 753 1095 757
rect 1099 753 1100 757
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1238 760 1244 761
rect 1238 756 1239 760
rect 1243 756 1244 760
rect 1238 755 1244 756
rect 1342 760 1348 761
rect 1342 756 1343 760
rect 1347 756 1348 760
rect 1342 755 1348 756
rect 1446 760 1452 761
rect 1446 756 1447 760
rect 1451 756 1452 760
rect 1446 755 1452 756
rect 1550 760 1556 761
rect 1550 756 1551 760
rect 1555 756 1556 760
rect 1550 755 1556 756
rect 1654 760 1660 761
rect 1654 756 1655 760
rect 1659 756 1660 760
rect 1654 755 1660 756
rect 1750 760 1756 761
rect 1750 756 1751 760
rect 1755 756 1756 760
rect 1750 755 1756 756
rect 1838 760 1844 761
rect 1838 756 1839 760
rect 1843 756 1844 760
rect 1838 755 1844 756
rect 1918 760 1924 761
rect 1918 756 1919 760
rect 1923 756 1924 760
rect 1918 755 1924 756
rect 2006 760 2012 761
rect 2006 756 2007 760
rect 2011 756 2012 760
rect 2006 755 2012 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2070 755 2076 756
rect 1094 752 1100 753
rect 1158 748 1164 749
rect 1134 745 1140 746
rect 159 743 168 744
rect 110 740 116 741
rect 110 736 111 740
rect 115 736 116 740
rect 159 739 160 743
rect 167 739 168 743
rect 159 738 168 739
rect 231 743 237 744
rect 231 739 232 743
rect 236 742 237 743
rect 286 743 292 744
rect 286 742 287 743
rect 236 740 287 742
rect 236 739 237 740
rect 231 738 237 739
rect 286 739 287 740
rect 291 739 292 743
rect 286 738 292 739
rect 318 743 325 744
rect 318 739 319 743
rect 324 739 325 743
rect 318 738 325 739
rect 390 743 396 744
rect 390 739 391 743
rect 395 742 396 743
rect 399 743 405 744
rect 399 742 400 743
rect 395 740 400 742
rect 395 739 396 740
rect 390 738 396 739
rect 399 739 400 740
rect 404 739 405 743
rect 399 738 405 739
rect 418 743 424 744
rect 418 739 419 743
rect 423 742 424 743
rect 471 743 477 744
rect 471 742 472 743
rect 423 740 472 742
rect 423 739 424 740
rect 418 738 424 739
rect 471 739 472 740
rect 476 739 477 743
rect 471 738 477 739
rect 479 743 485 744
rect 479 739 480 743
rect 484 742 485 743
rect 543 743 549 744
rect 543 742 544 743
rect 484 740 544 742
rect 484 739 485 740
rect 479 738 485 739
rect 543 739 544 740
rect 548 739 549 743
rect 543 738 549 739
rect 607 743 613 744
rect 607 739 608 743
rect 612 742 613 743
rect 615 743 621 744
rect 615 742 616 743
rect 612 740 616 742
rect 612 739 613 740
rect 607 738 613 739
rect 615 739 616 740
rect 620 739 621 743
rect 615 738 621 739
rect 663 743 669 744
rect 663 739 664 743
rect 668 742 669 743
rect 678 743 684 744
rect 678 742 679 743
rect 668 740 679 742
rect 668 739 669 740
rect 663 738 669 739
rect 678 739 679 740
rect 683 739 684 743
rect 678 738 684 739
rect 711 743 720 744
rect 711 739 712 743
rect 719 739 720 743
rect 711 738 720 739
rect 726 743 732 744
rect 726 739 727 743
rect 731 742 732 743
rect 767 743 773 744
rect 767 742 768 743
rect 731 740 768 742
rect 731 739 732 740
rect 726 738 732 739
rect 767 739 768 740
rect 772 739 773 743
rect 767 738 773 739
rect 823 743 829 744
rect 823 739 824 743
rect 828 742 829 743
rect 846 743 852 744
rect 846 742 847 743
rect 828 740 847 742
rect 828 739 829 740
rect 823 738 829 739
rect 846 739 847 740
rect 851 739 852 743
rect 846 738 852 739
rect 862 743 868 744
rect 862 739 863 743
rect 867 742 868 743
rect 879 743 885 744
rect 879 742 880 743
rect 867 740 880 742
rect 867 739 868 740
rect 862 738 868 739
rect 879 739 880 740
rect 884 739 885 743
rect 1134 741 1135 745
rect 1139 741 1140 745
rect 1158 744 1159 748
rect 1163 744 1164 748
rect 1158 743 1164 744
rect 1198 748 1204 749
rect 1198 744 1199 748
rect 1203 744 1204 748
rect 1198 743 1204 744
rect 1238 748 1244 749
rect 1238 744 1239 748
rect 1243 744 1244 748
rect 1238 743 1244 744
rect 1286 748 1292 749
rect 1286 744 1287 748
rect 1291 744 1292 748
rect 1286 743 1292 744
rect 1358 748 1364 749
rect 1358 744 1359 748
rect 1363 744 1364 748
rect 1358 743 1364 744
rect 1438 748 1444 749
rect 1438 744 1439 748
rect 1443 744 1444 748
rect 1438 743 1444 744
rect 1526 748 1532 749
rect 1526 744 1527 748
rect 1531 744 1532 748
rect 1526 743 1532 744
rect 1614 748 1620 749
rect 1614 744 1615 748
rect 1619 744 1620 748
rect 1614 743 1620 744
rect 1710 748 1716 749
rect 1710 744 1711 748
rect 1715 744 1716 748
rect 1710 743 1716 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1806 743 1812 744
rect 1902 748 1908 749
rect 1902 744 1903 748
rect 1907 744 1908 748
rect 1902 743 1908 744
rect 1998 748 2004 749
rect 1998 744 1999 748
rect 2003 744 2004 748
rect 1998 743 2004 744
rect 2070 748 2076 749
rect 2070 744 2071 748
rect 2075 744 2076 748
rect 2070 743 2076 744
rect 2118 745 2124 746
rect 879 738 885 739
rect 1094 740 1100 741
rect 1134 740 1140 741
rect 2118 741 2119 745
rect 2123 741 2124 745
rect 2118 740 2124 741
rect 110 735 116 736
rect 1094 736 1095 740
rect 1099 736 1100 740
rect 1094 735 1100 736
rect 1342 739 1348 740
rect 1342 735 1343 739
rect 1347 738 1348 739
rect 1347 736 1467 738
rect 1347 735 1348 736
rect 1342 734 1348 735
rect 134 732 140 733
rect 134 728 135 732
rect 139 728 140 732
rect 134 727 140 728
rect 206 732 212 733
rect 206 728 207 732
rect 211 728 212 732
rect 206 727 212 728
rect 294 732 300 733
rect 294 728 295 732
rect 299 728 300 732
rect 294 727 300 728
rect 374 732 380 733
rect 374 728 375 732
rect 379 728 380 732
rect 374 727 380 728
rect 446 732 452 733
rect 446 728 447 732
rect 451 728 452 732
rect 446 727 452 728
rect 518 732 524 733
rect 518 728 519 732
rect 523 728 524 732
rect 518 727 524 728
rect 582 732 588 733
rect 582 728 583 732
rect 587 728 588 732
rect 582 727 588 728
rect 638 732 644 733
rect 638 728 639 732
rect 643 728 644 732
rect 638 727 644 728
rect 686 732 692 733
rect 686 728 687 732
rect 691 728 692 732
rect 686 727 692 728
rect 742 732 748 733
rect 742 728 743 732
rect 747 728 748 732
rect 742 727 748 728
rect 798 732 804 733
rect 798 728 799 732
rect 803 728 804 732
rect 798 727 804 728
rect 854 732 860 733
rect 1465 732 1467 736
rect 854 728 855 732
rect 859 728 860 732
rect 1183 731 1192 732
rect 854 727 860 728
rect 1134 728 1140 729
rect 1134 724 1135 728
rect 1139 724 1140 728
rect 1183 727 1184 731
rect 1191 727 1192 731
rect 1183 726 1192 727
rect 1223 731 1232 732
rect 1223 727 1224 731
rect 1231 727 1232 731
rect 1223 726 1232 727
rect 1263 731 1269 732
rect 1263 727 1264 731
rect 1268 730 1269 731
rect 1278 731 1284 732
rect 1278 730 1279 731
rect 1268 728 1279 730
rect 1268 727 1269 728
rect 1263 726 1269 727
rect 1278 727 1279 728
rect 1283 727 1284 731
rect 1278 726 1284 727
rect 1311 731 1317 732
rect 1311 727 1312 731
rect 1316 730 1317 731
rect 1350 731 1356 732
rect 1350 730 1351 731
rect 1316 728 1351 730
rect 1316 727 1317 728
rect 1311 726 1317 727
rect 1350 727 1351 728
rect 1355 727 1356 731
rect 1350 726 1356 727
rect 1383 731 1389 732
rect 1383 727 1384 731
rect 1388 730 1389 731
rect 1430 731 1436 732
rect 1430 730 1431 731
rect 1388 728 1431 730
rect 1388 727 1389 728
rect 1383 726 1389 727
rect 1430 727 1431 728
rect 1435 727 1436 731
rect 1430 726 1436 727
rect 1463 731 1469 732
rect 1463 727 1464 731
rect 1468 727 1469 731
rect 1463 726 1469 727
rect 1551 731 1557 732
rect 1551 727 1552 731
rect 1556 730 1557 731
rect 1606 731 1612 732
rect 1606 730 1607 731
rect 1556 728 1607 730
rect 1556 727 1557 728
rect 1551 726 1557 727
rect 1606 727 1607 728
rect 1611 727 1612 731
rect 1606 726 1612 727
rect 1639 731 1645 732
rect 1639 727 1640 731
rect 1644 730 1645 731
rect 1702 731 1708 732
rect 1702 730 1703 731
rect 1644 728 1703 730
rect 1644 727 1645 728
rect 1639 726 1645 727
rect 1702 727 1703 728
rect 1707 727 1708 731
rect 1702 726 1708 727
rect 1718 731 1724 732
rect 1718 727 1719 731
rect 1723 730 1724 731
rect 1735 731 1741 732
rect 1735 730 1736 731
rect 1723 728 1736 730
rect 1723 727 1724 728
rect 1718 726 1724 727
rect 1735 727 1736 728
rect 1740 727 1741 731
rect 1735 726 1741 727
rect 1830 731 1837 732
rect 1830 727 1831 731
rect 1836 727 1837 731
rect 1830 726 1837 727
rect 1839 731 1845 732
rect 1839 727 1840 731
rect 1844 730 1845 731
rect 1927 731 1933 732
rect 1927 730 1928 731
rect 1844 728 1928 730
rect 1844 727 1845 728
rect 1839 726 1845 727
rect 1927 727 1928 728
rect 1932 727 1933 731
rect 1927 726 1933 727
rect 1935 731 1941 732
rect 1935 727 1936 731
rect 1940 730 1941 731
rect 2023 731 2029 732
rect 2023 730 2024 731
rect 1940 728 2024 730
rect 1940 727 1941 728
rect 1935 726 1941 727
rect 2023 727 2024 728
rect 2028 727 2029 731
rect 2023 726 2029 727
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 730 2084 731
rect 2095 731 2101 732
rect 2095 730 2096 731
rect 2083 728 2096 730
rect 2083 727 2084 728
rect 2078 726 2084 727
rect 2095 727 2096 728
rect 2100 727 2101 731
rect 2095 726 2101 727
rect 2118 728 2124 729
rect 1134 723 1140 724
rect 2118 724 2119 728
rect 2123 724 2124 728
rect 2118 723 2124 724
rect 1158 720 1164 721
rect 131 719 137 720
rect 131 715 132 719
rect 136 718 137 719
rect 158 719 164 720
rect 158 718 159 719
rect 136 716 159 718
rect 136 715 137 716
rect 131 714 137 715
rect 158 715 159 716
rect 163 715 164 719
rect 158 714 164 715
rect 203 719 209 720
rect 203 715 204 719
rect 208 718 209 719
rect 247 719 253 720
rect 247 718 248 719
rect 208 716 248 718
rect 208 715 209 716
rect 203 714 209 715
rect 247 715 248 716
rect 252 715 253 719
rect 247 714 253 715
rect 286 719 297 720
rect 286 715 287 719
rect 291 715 292 719
rect 296 715 297 719
rect 286 714 297 715
rect 371 719 377 720
rect 371 715 372 719
rect 376 718 377 719
rect 418 719 424 720
rect 418 718 419 719
rect 376 716 419 718
rect 376 715 377 716
rect 371 714 377 715
rect 418 715 419 716
rect 423 715 424 719
rect 418 714 424 715
rect 443 719 449 720
rect 443 715 444 719
rect 448 718 449 719
rect 479 719 485 720
rect 479 718 480 719
rect 448 716 480 718
rect 448 715 449 716
rect 443 714 449 715
rect 479 715 480 716
rect 484 715 485 719
rect 479 714 485 715
rect 515 719 521 720
rect 515 715 516 719
rect 520 718 521 719
rect 554 719 560 720
rect 554 718 555 719
rect 520 716 555 718
rect 520 715 521 716
rect 515 714 521 715
rect 554 715 555 716
rect 559 715 560 719
rect 554 714 560 715
rect 579 719 585 720
rect 579 715 580 719
rect 584 718 585 719
rect 606 719 612 720
rect 606 718 607 719
rect 584 716 607 718
rect 584 715 585 716
rect 579 714 585 715
rect 606 715 607 716
rect 611 715 612 719
rect 606 714 612 715
rect 635 719 641 720
rect 635 715 636 719
rect 640 718 641 719
rect 678 719 689 720
rect 640 716 674 718
rect 640 715 641 716
rect 635 714 641 715
rect 672 710 674 716
rect 678 715 679 719
rect 683 715 684 719
rect 688 715 689 719
rect 678 714 689 715
rect 739 719 745 720
rect 739 715 740 719
rect 744 718 745 719
rect 790 719 801 720
rect 744 715 746 718
rect 739 714 746 715
rect 790 715 791 719
rect 795 715 796 719
rect 800 715 801 719
rect 790 714 801 715
rect 846 719 857 720
rect 846 715 847 719
rect 851 715 852 719
rect 856 715 857 719
rect 1158 716 1159 720
rect 1163 716 1164 720
rect 1158 715 1164 716
rect 1198 720 1204 721
rect 1198 716 1199 720
rect 1203 716 1204 720
rect 1198 715 1204 716
rect 1238 720 1244 721
rect 1238 716 1239 720
rect 1243 716 1244 720
rect 1238 715 1244 716
rect 1286 720 1292 721
rect 1286 716 1287 720
rect 1291 716 1292 720
rect 1286 715 1292 716
rect 1358 720 1364 721
rect 1358 716 1359 720
rect 1363 716 1364 720
rect 1358 715 1364 716
rect 1438 720 1444 721
rect 1438 716 1439 720
rect 1443 716 1444 720
rect 1438 715 1444 716
rect 1526 720 1532 721
rect 1526 716 1527 720
rect 1531 716 1532 720
rect 1526 715 1532 716
rect 1614 720 1620 721
rect 1614 716 1615 720
rect 1619 716 1620 720
rect 1614 715 1620 716
rect 1710 720 1716 721
rect 1710 716 1711 720
rect 1715 716 1716 720
rect 1710 715 1716 716
rect 1806 720 1812 721
rect 1806 716 1807 720
rect 1811 716 1812 720
rect 1806 715 1812 716
rect 1902 720 1908 721
rect 1902 716 1903 720
rect 1907 716 1908 720
rect 1902 715 1908 716
rect 1998 720 2004 721
rect 1998 716 1999 720
rect 2003 716 2004 720
rect 1998 715 2004 716
rect 2070 720 2076 721
rect 2070 716 2071 720
rect 2075 716 2076 720
rect 2070 715 2076 716
rect 846 714 857 715
rect 726 711 732 712
rect 726 710 727 711
rect 672 708 727 710
rect 726 707 727 708
rect 731 707 732 711
rect 744 710 746 714
rect 862 711 868 712
rect 862 710 863 711
rect 744 708 863 710
rect 726 706 732 707
rect 862 707 863 708
rect 867 707 868 711
rect 862 706 868 707
rect 1155 707 1161 708
rect 131 703 137 704
rect 131 699 132 703
rect 136 702 137 703
rect 170 703 176 704
rect 170 702 171 703
rect 136 700 171 702
rect 136 699 137 700
rect 131 698 137 699
rect 170 699 171 700
rect 175 699 176 703
rect 170 698 176 699
rect 179 703 185 704
rect 179 699 180 703
rect 184 702 185 703
rect 234 703 240 704
rect 234 702 235 703
rect 184 700 235 702
rect 184 699 185 700
rect 179 698 185 699
rect 234 699 235 700
rect 239 699 240 703
rect 234 698 240 699
rect 243 703 249 704
rect 243 699 244 703
rect 248 702 249 703
rect 282 703 288 704
rect 282 702 283 703
rect 248 700 283 702
rect 248 699 249 700
rect 243 698 249 699
rect 282 699 283 700
rect 287 699 288 703
rect 282 698 288 699
rect 307 703 313 704
rect 307 699 308 703
rect 312 702 313 703
rect 318 703 324 704
rect 318 702 319 703
rect 312 700 319 702
rect 312 699 313 700
rect 307 698 313 699
rect 318 699 319 700
rect 323 699 324 703
rect 318 698 324 699
rect 379 703 385 704
rect 379 699 380 703
rect 384 702 385 703
rect 390 703 396 704
rect 390 702 391 703
rect 384 700 391 702
rect 384 699 385 700
rect 379 698 385 699
rect 390 699 391 700
rect 395 699 396 703
rect 390 698 396 699
rect 410 703 416 704
rect 410 699 411 703
rect 415 702 416 703
rect 451 703 457 704
rect 451 702 452 703
rect 415 700 452 702
rect 415 699 416 700
rect 410 698 416 699
rect 451 699 452 700
rect 456 699 457 703
rect 451 698 457 699
rect 482 703 488 704
rect 482 699 483 703
rect 487 702 488 703
rect 515 703 521 704
rect 515 702 516 703
rect 487 700 516 702
rect 487 699 488 700
rect 482 698 488 699
rect 515 699 516 700
rect 520 699 521 703
rect 515 698 521 699
rect 579 703 585 704
rect 579 699 580 703
rect 584 702 585 703
rect 630 703 636 704
rect 630 702 631 703
rect 584 700 631 702
rect 584 699 585 700
rect 579 698 585 699
rect 630 699 631 700
rect 635 699 636 703
rect 630 698 636 699
rect 643 703 649 704
rect 643 699 644 703
rect 648 702 649 703
rect 654 703 660 704
rect 654 702 655 703
rect 648 700 655 702
rect 648 699 649 700
rect 643 698 649 699
rect 654 699 655 700
rect 659 699 660 703
rect 654 698 660 699
rect 707 703 713 704
rect 707 699 708 703
rect 712 702 713 703
rect 734 703 740 704
rect 734 702 735 703
rect 712 700 735 702
rect 712 699 713 700
rect 707 698 713 699
rect 734 699 735 700
rect 739 699 740 703
rect 734 698 740 699
rect 743 703 749 704
rect 743 699 744 703
rect 748 702 749 703
rect 763 703 769 704
rect 763 702 764 703
rect 748 700 764 702
rect 748 699 749 700
rect 743 698 749 699
rect 763 699 764 700
rect 768 699 769 703
rect 763 698 769 699
rect 814 703 825 704
rect 814 699 815 703
rect 819 699 820 703
rect 824 699 825 703
rect 814 698 825 699
rect 855 703 861 704
rect 855 699 856 703
rect 860 702 861 703
rect 875 703 881 704
rect 875 702 876 703
rect 860 700 876 702
rect 860 699 861 700
rect 855 698 861 699
rect 875 699 876 700
rect 880 699 881 703
rect 875 698 881 699
rect 906 703 912 704
rect 906 699 907 703
rect 911 702 912 703
rect 939 703 945 704
rect 939 702 940 703
rect 911 700 940 702
rect 911 699 912 700
rect 906 698 912 699
rect 939 699 940 700
rect 944 699 945 703
rect 1155 703 1156 707
rect 1160 703 1161 707
rect 1155 702 1161 703
rect 1186 707 1192 708
rect 1186 703 1187 707
rect 1191 706 1192 707
rect 1195 707 1201 708
rect 1195 706 1196 707
rect 1191 704 1196 706
rect 1191 703 1192 704
rect 1186 702 1192 703
rect 1195 703 1196 704
rect 1200 703 1201 707
rect 1195 702 1201 703
rect 1226 707 1232 708
rect 1226 703 1227 707
rect 1231 706 1232 707
rect 1235 707 1241 708
rect 1235 706 1236 707
rect 1231 704 1236 706
rect 1231 703 1232 704
rect 1226 702 1232 703
rect 1235 703 1236 704
rect 1240 703 1241 707
rect 1235 702 1241 703
rect 1278 707 1289 708
rect 1278 703 1279 707
rect 1283 703 1284 707
rect 1288 703 1289 707
rect 1278 702 1289 703
rect 1350 707 1361 708
rect 1350 703 1351 707
rect 1355 703 1356 707
rect 1360 703 1361 707
rect 1350 702 1361 703
rect 1430 707 1441 708
rect 1430 703 1431 707
rect 1435 703 1436 707
rect 1440 703 1441 707
rect 1430 702 1441 703
rect 1518 707 1529 708
rect 1518 703 1519 707
rect 1523 703 1524 707
rect 1528 703 1529 707
rect 1518 702 1529 703
rect 1606 707 1617 708
rect 1606 703 1607 707
rect 1611 703 1612 707
rect 1616 703 1617 707
rect 1606 702 1617 703
rect 1702 707 1713 708
rect 1702 703 1703 707
rect 1707 703 1708 707
rect 1712 703 1713 707
rect 1702 702 1713 703
rect 1803 707 1809 708
rect 1803 703 1804 707
rect 1808 706 1809 707
rect 1839 707 1845 708
rect 1839 706 1840 707
rect 1808 704 1840 706
rect 1808 703 1809 704
rect 1803 702 1809 703
rect 1839 703 1840 704
rect 1844 703 1845 707
rect 1839 702 1845 703
rect 1899 707 1905 708
rect 1899 703 1900 707
rect 1904 706 1905 707
rect 1935 707 1941 708
rect 1935 706 1936 707
rect 1904 704 1936 706
rect 1904 703 1905 704
rect 1899 702 1905 703
rect 1935 703 1936 704
rect 1940 703 1941 707
rect 1935 702 1941 703
rect 1986 707 1992 708
rect 1986 703 1987 707
rect 1991 706 1992 707
rect 1995 707 2001 708
rect 1995 706 1996 707
rect 1991 704 1996 706
rect 1991 703 1992 704
rect 1986 702 1992 703
rect 1995 703 1996 704
rect 2000 703 2001 707
rect 1995 702 2001 703
rect 2067 707 2073 708
rect 2067 703 2068 707
rect 2072 706 2073 707
rect 2086 707 2092 708
rect 2086 706 2087 707
rect 2072 704 2087 706
rect 2072 703 2073 704
rect 2067 702 2073 703
rect 2086 703 2087 704
rect 2091 703 2092 707
rect 2086 702 2092 703
rect 939 698 945 699
rect 1159 698 1161 702
rect 1310 699 1316 700
rect 1310 698 1311 699
rect 1159 696 1311 698
rect 1310 695 1311 696
rect 1315 695 1316 699
rect 1534 699 1540 700
rect 1534 698 1535 699
rect 1310 694 1316 695
rect 1388 696 1535 698
rect 1388 694 1390 696
rect 1534 695 1535 696
rect 1539 695 1540 699
rect 1718 699 1724 700
rect 1718 698 1719 699
rect 1534 694 1540 695
rect 1636 696 1719 698
rect 1636 694 1638 696
rect 1718 695 1719 696
rect 1723 695 1724 699
rect 1718 694 1724 695
rect 1387 693 1393 694
rect 134 692 140 693
rect 134 688 135 692
rect 139 688 140 692
rect 134 687 140 688
rect 182 692 188 693
rect 182 688 183 692
rect 187 688 188 692
rect 182 687 188 688
rect 246 692 252 693
rect 246 688 247 692
rect 251 688 252 692
rect 246 687 252 688
rect 310 692 316 693
rect 310 688 311 692
rect 315 688 316 692
rect 310 687 316 688
rect 382 692 388 693
rect 382 688 383 692
rect 387 688 388 692
rect 382 687 388 688
rect 454 692 460 693
rect 454 688 455 692
rect 459 688 460 692
rect 454 687 460 688
rect 518 692 524 693
rect 518 688 519 692
rect 523 688 524 692
rect 518 687 524 688
rect 582 692 588 693
rect 582 688 583 692
rect 587 688 588 692
rect 582 687 588 688
rect 646 692 652 693
rect 646 688 647 692
rect 651 688 652 692
rect 646 687 652 688
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 766 692 772 693
rect 766 688 767 692
rect 771 688 772 692
rect 766 687 772 688
rect 822 692 828 693
rect 822 688 823 692
rect 827 688 828 692
rect 822 687 828 688
rect 878 692 884 693
rect 878 688 879 692
rect 883 688 884 692
rect 878 687 884 688
rect 942 692 948 693
rect 942 688 943 692
rect 947 688 948 692
rect 942 687 948 688
rect 1235 691 1241 692
rect 1235 687 1236 691
rect 1240 690 1241 691
rect 1274 691 1280 692
rect 1274 690 1275 691
rect 1240 688 1275 690
rect 1240 687 1241 688
rect 1235 686 1241 687
rect 1274 687 1275 688
rect 1279 687 1280 691
rect 1274 686 1280 687
rect 1283 691 1289 692
rect 1283 687 1284 691
rect 1288 690 1289 691
rect 1322 691 1328 692
rect 1322 690 1323 691
rect 1288 688 1323 690
rect 1288 687 1289 688
rect 1283 686 1289 687
rect 1322 687 1323 688
rect 1327 687 1328 691
rect 1322 686 1328 687
rect 1331 691 1337 692
rect 1331 687 1332 691
rect 1336 690 1337 691
rect 1342 691 1348 692
rect 1342 690 1343 691
rect 1336 688 1343 690
rect 1336 687 1337 688
rect 1331 686 1337 687
rect 1342 687 1343 688
rect 1347 687 1348 691
rect 1387 689 1388 693
rect 1392 689 1393 693
rect 1635 693 1641 694
rect 1387 688 1393 689
rect 1423 691 1429 692
rect 1342 686 1348 687
rect 1423 687 1424 691
rect 1428 690 1429 691
rect 1443 691 1449 692
rect 1443 690 1444 691
rect 1428 688 1444 690
rect 1428 687 1429 688
rect 1423 686 1429 687
rect 1443 687 1444 688
rect 1448 687 1449 691
rect 1443 686 1449 687
rect 1507 691 1513 692
rect 1507 687 1508 691
rect 1512 690 1513 691
rect 1562 691 1568 692
rect 1562 690 1563 691
rect 1512 688 1563 690
rect 1512 687 1513 688
rect 1507 686 1513 687
rect 1562 687 1563 688
rect 1567 687 1568 691
rect 1562 686 1568 687
rect 1571 691 1577 692
rect 1571 687 1572 691
rect 1576 690 1577 691
rect 1626 691 1632 692
rect 1626 690 1627 691
rect 1576 688 1627 690
rect 1576 687 1577 688
rect 1571 686 1577 687
rect 1626 687 1627 688
rect 1631 687 1632 691
rect 1635 689 1636 693
rect 1640 689 1641 693
rect 1635 688 1641 689
rect 1699 691 1705 692
rect 1626 686 1632 687
rect 1699 687 1700 691
rect 1704 690 1705 691
rect 1730 691 1736 692
rect 1704 688 1714 690
rect 1704 687 1705 688
rect 1699 686 1705 687
rect 1710 687 1716 688
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 1094 684 1100 685
rect 1094 680 1095 684
rect 1099 680 1100 684
rect 1710 683 1711 687
rect 1715 683 1716 687
rect 1730 687 1731 691
rect 1735 690 1736 691
rect 1763 691 1769 692
rect 1763 690 1764 691
rect 1735 688 1764 690
rect 1735 687 1736 688
rect 1730 686 1736 687
rect 1763 687 1764 688
rect 1768 687 1769 691
rect 1763 686 1769 687
rect 1807 691 1813 692
rect 1807 687 1808 691
rect 1812 690 1813 691
rect 1827 691 1833 692
rect 1827 690 1828 691
rect 1812 688 1828 690
rect 1812 687 1813 688
rect 1807 686 1813 687
rect 1827 687 1828 688
rect 1832 687 1833 691
rect 1827 686 1833 687
rect 1858 691 1864 692
rect 1858 687 1859 691
rect 1863 690 1864 691
rect 1891 691 1897 692
rect 1891 690 1892 691
rect 1863 688 1892 690
rect 1863 687 1864 688
rect 1858 686 1864 687
rect 1891 687 1892 688
rect 1896 687 1897 691
rect 1891 686 1897 687
rect 1930 691 1936 692
rect 1930 687 1931 691
rect 1935 690 1936 691
rect 1955 691 1961 692
rect 1955 690 1956 691
rect 1935 688 1956 690
rect 1935 687 1936 688
rect 1930 686 1936 687
rect 1955 687 1956 688
rect 1960 687 1961 691
rect 1955 686 1961 687
rect 2019 691 2025 692
rect 2019 687 2020 691
rect 2024 690 2025 691
rect 2058 691 2064 692
rect 2058 690 2059 691
rect 2024 688 2059 690
rect 2024 687 2025 688
rect 2019 686 2025 687
rect 2058 687 2059 688
rect 2063 687 2064 691
rect 2058 686 2064 687
rect 2067 691 2073 692
rect 2067 687 2068 691
rect 2072 690 2073 691
rect 2078 691 2084 692
rect 2078 690 2079 691
rect 2072 688 2079 690
rect 2072 687 2073 688
rect 2067 686 2073 687
rect 2078 687 2079 688
rect 2083 687 2084 691
rect 2078 686 2084 687
rect 1710 682 1716 683
rect 110 679 116 680
rect 158 679 165 680
rect 158 675 159 679
rect 164 675 165 679
rect 158 674 165 675
rect 170 679 176 680
rect 170 675 171 679
rect 175 678 176 679
rect 207 679 213 680
rect 207 678 208 679
rect 175 676 208 678
rect 175 675 176 676
rect 170 674 176 675
rect 207 675 208 676
rect 212 675 213 679
rect 207 674 213 675
rect 271 679 280 680
rect 271 675 272 679
rect 279 675 280 679
rect 271 674 280 675
rect 282 679 288 680
rect 282 675 283 679
rect 287 678 288 679
rect 335 679 341 680
rect 335 678 336 679
rect 287 676 336 678
rect 287 675 288 676
rect 282 674 288 675
rect 335 675 336 676
rect 340 675 341 679
rect 335 674 341 675
rect 407 679 416 680
rect 407 675 408 679
rect 415 675 416 679
rect 407 674 416 675
rect 479 679 488 680
rect 479 675 480 679
rect 487 675 488 679
rect 479 674 488 675
rect 534 679 540 680
rect 534 675 535 679
rect 539 678 540 679
rect 543 679 549 680
rect 543 678 544 679
rect 539 676 544 678
rect 539 675 540 676
rect 534 674 540 675
rect 543 675 544 676
rect 548 675 549 679
rect 543 674 549 675
rect 606 679 613 680
rect 606 675 607 679
rect 612 675 613 679
rect 606 674 613 675
rect 630 679 636 680
rect 630 675 631 679
rect 635 678 636 679
rect 671 679 677 680
rect 671 678 672 679
rect 635 676 672 678
rect 635 675 636 676
rect 630 674 636 675
rect 671 675 672 676
rect 676 675 677 679
rect 671 674 677 675
rect 735 679 741 680
rect 735 675 736 679
rect 740 678 741 679
rect 743 679 749 680
rect 743 678 744 679
rect 740 676 744 678
rect 740 675 741 676
rect 735 674 741 675
rect 743 675 744 676
rect 748 675 749 679
rect 743 674 749 675
rect 790 679 797 680
rect 790 675 791 679
rect 796 675 797 679
rect 790 674 797 675
rect 847 679 853 680
rect 847 675 848 679
rect 852 678 853 679
rect 855 679 861 680
rect 855 678 856 679
rect 852 676 856 678
rect 852 675 853 676
rect 847 674 853 675
rect 855 675 856 676
rect 860 675 861 679
rect 855 674 861 675
rect 903 679 912 680
rect 903 675 904 679
rect 911 675 912 679
rect 903 674 912 675
rect 966 679 973 680
rect 1094 679 1100 680
rect 1238 680 1244 681
rect 966 675 967 679
rect 972 675 973 679
rect 1238 676 1239 680
rect 1243 676 1244 680
rect 1238 675 1244 676
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1574 680 1580 681
rect 1574 676 1575 680
rect 1579 676 1580 680
rect 1574 675 1580 676
rect 1638 680 1644 681
rect 1638 676 1639 680
rect 1643 676 1644 680
rect 1638 675 1644 676
rect 1702 680 1708 681
rect 1702 676 1703 680
rect 1707 676 1708 680
rect 1702 675 1708 676
rect 1766 680 1772 681
rect 1766 676 1767 680
rect 1771 676 1772 680
rect 1766 675 1772 676
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1894 680 1900 681
rect 1894 676 1895 680
rect 1899 676 1900 680
rect 1894 675 1900 676
rect 1958 680 1964 681
rect 1958 676 1959 680
rect 1963 676 1964 680
rect 1958 675 1964 676
rect 2022 680 2028 681
rect 2022 676 2023 680
rect 2027 676 2028 680
rect 2022 675 2028 676
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 966 674 973 675
rect 1134 672 1140 673
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 1094 667 1100 668
rect 1134 667 1140 668
rect 1263 667 1272 668
rect 110 662 116 663
rect 134 664 140 665
rect 134 660 135 664
rect 139 660 140 664
rect 134 659 140 660
rect 182 664 188 665
rect 182 660 183 664
rect 187 660 188 664
rect 182 659 188 660
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 310 664 316 665
rect 310 660 311 664
rect 315 660 316 664
rect 310 659 316 660
rect 382 664 388 665
rect 382 660 383 664
rect 387 660 388 664
rect 382 659 388 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 518 664 524 665
rect 518 660 519 664
rect 523 660 524 664
rect 518 659 524 660
rect 582 664 588 665
rect 582 660 583 664
rect 587 660 588 664
rect 582 659 588 660
rect 646 664 652 665
rect 646 660 647 664
rect 651 660 652 664
rect 646 659 652 660
rect 710 664 716 665
rect 710 660 711 664
rect 715 660 716 664
rect 710 659 716 660
rect 766 664 772 665
rect 766 660 767 664
rect 771 660 772 664
rect 766 659 772 660
rect 822 664 828 665
rect 822 660 823 664
rect 827 660 828 664
rect 822 659 828 660
rect 878 664 884 665
rect 878 660 879 664
rect 883 660 884 664
rect 878 659 884 660
rect 942 664 948 665
rect 942 660 943 664
rect 947 660 948 664
rect 1094 663 1095 667
rect 1099 663 1100 667
rect 1094 662 1100 663
rect 1263 663 1264 667
rect 1271 663 1272 667
rect 1263 662 1272 663
rect 1274 667 1280 668
rect 1274 663 1275 667
rect 1279 666 1280 667
rect 1311 667 1317 668
rect 1311 666 1312 667
rect 1279 664 1312 666
rect 1279 663 1280 664
rect 1274 662 1280 663
rect 1311 663 1312 664
rect 1316 663 1317 667
rect 1311 662 1317 663
rect 1322 667 1328 668
rect 1322 663 1323 667
rect 1327 666 1328 667
rect 1359 667 1365 668
rect 1359 666 1360 667
rect 1327 664 1360 666
rect 1327 663 1328 664
rect 1322 662 1328 663
rect 1359 663 1360 664
rect 1364 663 1365 667
rect 1359 662 1365 663
rect 1415 667 1421 668
rect 1415 663 1416 667
rect 1420 666 1421 667
rect 1423 667 1429 668
rect 1423 666 1424 667
rect 1420 664 1424 666
rect 1420 663 1421 664
rect 1415 662 1421 663
rect 1423 663 1424 664
rect 1428 663 1429 667
rect 1423 662 1429 663
rect 1470 667 1477 668
rect 1470 663 1471 667
rect 1476 663 1477 667
rect 1470 662 1477 663
rect 1534 667 1541 668
rect 1534 663 1535 667
rect 1540 663 1541 667
rect 1534 662 1541 663
rect 1562 667 1568 668
rect 1562 663 1563 667
rect 1567 666 1568 667
rect 1599 667 1605 668
rect 1599 666 1600 667
rect 1567 664 1600 666
rect 1567 663 1568 664
rect 1562 662 1568 663
rect 1599 663 1600 664
rect 1604 663 1605 667
rect 1599 662 1605 663
rect 1626 667 1632 668
rect 1626 663 1627 667
rect 1631 666 1632 667
rect 1663 667 1669 668
rect 1663 666 1664 667
rect 1631 664 1664 666
rect 1631 663 1632 664
rect 1626 662 1632 663
rect 1663 663 1664 664
rect 1668 663 1669 667
rect 1663 662 1669 663
rect 1727 667 1736 668
rect 1727 663 1728 667
rect 1735 663 1736 667
rect 1727 662 1736 663
rect 1791 667 1797 668
rect 1791 663 1792 667
rect 1796 666 1797 667
rect 1807 667 1813 668
rect 1807 666 1808 667
rect 1796 664 1808 666
rect 1796 663 1797 664
rect 1791 662 1797 663
rect 1807 663 1808 664
rect 1812 663 1813 667
rect 1807 662 1813 663
rect 1855 667 1864 668
rect 1855 663 1856 667
rect 1863 663 1864 667
rect 1855 662 1864 663
rect 1919 667 1925 668
rect 1919 663 1920 667
rect 1924 666 1925 667
rect 1930 667 1936 668
rect 1930 666 1931 667
rect 1924 664 1931 666
rect 1924 663 1925 664
rect 1919 662 1925 663
rect 1930 663 1931 664
rect 1935 663 1936 667
rect 1930 662 1936 663
rect 1983 667 1992 668
rect 1983 663 1984 667
rect 1991 663 1992 667
rect 1983 662 1992 663
rect 2047 667 2056 668
rect 2047 663 2048 667
rect 2055 663 2056 667
rect 2047 662 2056 663
rect 2058 667 2064 668
rect 2058 663 2059 667
rect 2063 666 2064 667
rect 2095 667 2101 668
rect 2118 667 2124 668
rect 2095 666 2096 667
rect 2063 664 2096 666
rect 2063 663 2064 664
rect 2058 662 2064 663
rect 2095 663 2096 664
rect 2100 663 2101 667
rect 2095 662 2101 663
rect 942 659 948 660
rect 1134 655 1140 656
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 2118 655 2124 656
rect 1134 650 1140 651
rect 1238 652 1244 653
rect 1238 648 1239 652
rect 1243 648 1244 652
rect 1238 647 1244 648
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1574 652 1580 653
rect 1574 648 1575 652
rect 1579 648 1580 652
rect 1574 647 1580 648
rect 1638 652 1644 653
rect 1638 648 1639 652
rect 1643 648 1644 652
rect 1638 647 1644 648
rect 1702 652 1708 653
rect 1702 648 1703 652
rect 1707 648 1708 652
rect 1702 647 1708 648
rect 1766 652 1772 653
rect 1766 648 1767 652
rect 1771 648 1772 652
rect 1766 647 1772 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1830 647 1836 648
rect 1894 652 1900 653
rect 1894 648 1895 652
rect 1899 648 1900 652
rect 1894 647 1900 648
rect 1958 652 1964 653
rect 1958 648 1959 652
rect 1963 648 1964 652
rect 1958 647 1964 648
rect 2022 652 2028 653
rect 2022 648 2023 652
rect 2027 648 2028 652
rect 2022 647 2028 648
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 158 644 164 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 158 640 159 644
rect 163 640 164 644
rect 158 639 164 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 454 644 460 645
rect 454 640 455 644
rect 459 640 460 644
rect 454 639 460 640
rect 542 644 548 645
rect 542 640 543 644
rect 547 640 548 644
rect 542 639 548 640
rect 630 644 636 645
rect 630 640 631 644
rect 635 640 636 644
rect 630 639 636 640
rect 718 644 724 645
rect 718 640 719 644
rect 723 640 724 644
rect 718 639 724 640
rect 798 644 804 645
rect 798 640 799 644
rect 803 640 804 644
rect 798 639 804 640
rect 870 644 876 645
rect 870 640 871 644
rect 875 640 876 644
rect 870 639 876 640
rect 950 644 956 645
rect 950 640 951 644
rect 955 640 956 644
rect 950 639 956 640
rect 1030 644 1036 645
rect 1030 640 1031 644
rect 1035 640 1036 644
rect 1030 639 1036 640
rect 1094 641 1100 642
rect 110 636 116 637
rect 1094 637 1095 641
rect 1099 637 1100 641
rect 1278 640 1284 641
rect 1094 636 1100 637
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1318 640 1324 641
rect 1318 636 1319 640
rect 1323 636 1324 640
rect 1318 635 1324 636
rect 1366 640 1372 641
rect 1366 636 1367 640
rect 1371 636 1372 640
rect 1366 635 1372 636
rect 1422 640 1428 641
rect 1422 636 1423 640
rect 1427 636 1428 640
rect 1422 635 1428 636
rect 1478 640 1484 641
rect 1478 636 1479 640
rect 1483 636 1484 640
rect 1478 635 1484 636
rect 1534 640 1540 641
rect 1534 636 1535 640
rect 1539 636 1540 640
rect 1534 635 1540 636
rect 1590 640 1596 641
rect 1590 636 1591 640
rect 1595 636 1596 640
rect 1590 635 1596 636
rect 1646 640 1652 641
rect 1646 636 1647 640
rect 1651 636 1652 640
rect 1646 635 1652 636
rect 1718 640 1724 641
rect 1718 636 1719 640
rect 1723 636 1724 640
rect 1718 635 1724 636
rect 1798 640 1804 641
rect 1798 636 1799 640
rect 1803 636 1804 640
rect 1798 635 1804 636
rect 1878 640 1884 641
rect 1878 636 1879 640
rect 1883 636 1884 640
rect 1878 635 1884 636
rect 1966 640 1972 641
rect 1966 636 1967 640
rect 1971 636 1972 640
rect 1966 635 1972 636
rect 2062 640 2068 641
rect 2062 636 2063 640
rect 2067 636 2068 640
rect 2062 635 2068 636
rect 2118 637 2124 638
rect 1134 632 1140 633
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 1342 631 1348 632
rect 183 627 189 628
rect 110 624 116 625
rect 110 620 111 624
rect 115 620 116 624
rect 183 623 184 627
rect 188 626 189 627
rect 206 627 212 628
rect 206 626 207 627
rect 188 624 207 626
rect 188 623 189 624
rect 183 622 189 623
rect 206 623 207 624
rect 211 623 212 627
rect 206 622 212 623
rect 234 627 245 628
rect 234 623 235 627
rect 239 623 240 627
rect 244 623 245 627
rect 234 622 245 623
rect 262 627 268 628
rect 262 623 263 627
rect 267 626 268 627
rect 311 627 317 628
rect 311 626 312 627
rect 267 624 312 626
rect 267 623 268 624
rect 262 622 268 623
rect 311 623 312 624
rect 316 623 317 627
rect 311 622 317 623
rect 390 627 397 628
rect 390 623 391 627
rect 396 623 397 627
rect 390 622 397 623
rect 402 627 408 628
rect 402 623 403 627
rect 407 626 408 627
rect 479 627 485 628
rect 479 626 480 627
rect 407 624 480 626
rect 407 623 408 624
rect 402 622 408 623
rect 479 623 480 624
rect 484 623 485 627
rect 479 622 485 623
rect 487 627 493 628
rect 487 623 488 627
rect 492 626 493 627
rect 567 627 573 628
rect 567 626 568 627
rect 492 624 568 626
rect 492 623 493 624
rect 487 622 493 623
rect 567 623 568 624
rect 572 623 573 627
rect 567 622 573 623
rect 654 627 661 628
rect 654 623 655 627
rect 660 623 661 627
rect 654 622 661 623
rect 743 627 749 628
rect 743 623 744 627
rect 748 626 749 627
rect 790 627 796 628
rect 790 626 791 627
rect 748 624 791 626
rect 748 623 749 624
rect 743 622 749 623
rect 790 623 791 624
rect 795 623 796 627
rect 790 622 796 623
rect 814 627 820 628
rect 814 623 815 627
rect 819 626 820 627
rect 823 627 829 628
rect 823 626 824 627
rect 819 624 824 626
rect 819 623 820 624
rect 814 622 820 623
rect 823 623 824 624
rect 828 623 829 627
rect 823 622 829 623
rect 895 627 901 628
rect 895 623 896 627
rect 900 626 901 627
rect 942 627 948 628
rect 942 626 943 627
rect 900 624 943 626
rect 900 623 901 624
rect 895 622 901 623
rect 942 623 943 624
rect 947 623 948 627
rect 942 622 948 623
rect 975 627 981 628
rect 975 623 976 627
rect 980 626 981 627
rect 1022 627 1028 628
rect 1022 626 1023 627
rect 980 624 1023 626
rect 980 623 981 624
rect 975 622 981 623
rect 1022 623 1023 624
rect 1027 623 1028 627
rect 1022 622 1028 623
rect 1038 627 1044 628
rect 1038 623 1039 627
rect 1043 626 1044 627
rect 1055 627 1061 628
rect 1055 626 1056 627
rect 1043 624 1056 626
rect 1043 623 1044 624
rect 1038 622 1044 623
rect 1055 623 1056 624
rect 1060 623 1061 627
rect 1342 627 1343 631
rect 1347 630 1348 631
rect 1710 631 1716 632
rect 1347 628 1418 630
rect 1347 627 1348 628
rect 1342 626 1348 627
rect 1055 622 1061 623
rect 1094 624 1100 625
rect 110 619 116 620
rect 1094 620 1095 624
rect 1099 620 1100 624
rect 1303 623 1312 624
rect 1094 619 1100 620
rect 1134 620 1140 621
rect 158 616 164 617
rect 158 612 159 616
rect 163 612 164 616
rect 158 611 164 612
rect 214 616 220 617
rect 214 612 215 616
rect 219 612 220 616
rect 214 611 220 612
rect 286 616 292 617
rect 286 612 287 616
rect 291 612 292 616
rect 286 611 292 612
rect 366 616 372 617
rect 366 612 367 616
rect 371 612 372 616
rect 366 611 372 612
rect 454 616 460 617
rect 454 612 455 616
rect 459 612 460 616
rect 454 611 460 612
rect 542 616 548 617
rect 542 612 543 616
rect 547 612 548 616
rect 542 611 548 612
rect 630 616 636 617
rect 630 612 631 616
rect 635 612 636 616
rect 630 611 636 612
rect 718 616 724 617
rect 718 612 719 616
rect 723 612 724 616
rect 718 611 724 612
rect 798 616 804 617
rect 798 612 799 616
rect 803 612 804 616
rect 798 611 804 612
rect 870 616 876 617
rect 870 612 871 616
rect 875 612 876 616
rect 870 611 876 612
rect 950 616 956 617
rect 950 612 951 616
rect 955 612 956 616
rect 950 611 956 612
rect 1030 616 1036 617
rect 1030 612 1031 616
rect 1035 612 1036 616
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1303 619 1304 623
rect 1311 619 1312 623
rect 1303 618 1312 619
rect 1343 623 1349 624
rect 1343 619 1344 623
rect 1348 622 1349 623
rect 1358 623 1364 624
rect 1358 622 1359 623
rect 1348 620 1359 622
rect 1348 619 1349 620
rect 1343 618 1349 619
rect 1358 619 1359 620
rect 1363 619 1364 623
rect 1358 618 1364 619
rect 1391 623 1397 624
rect 1391 619 1392 623
rect 1396 622 1397 623
rect 1406 623 1412 624
rect 1406 622 1407 623
rect 1396 620 1407 622
rect 1396 619 1397 620
rect 1391 618 1397 619
rect 1406 619 1407 620
rect 1411 619 1412 623
rect 1416 622 1418 628
rect 1710 627 1711 631
rect 1715 630 1716 631
rect 1715 628 1970 630
rect 1715 627 1716 628
rect 1710 626 1716 627
rect 1447 623 1453 624
rect 1447 622 1448 623
rect 1416 620 1448 622
rect 1406 618 1412 619
rect 1447 619 1448 620
rect 1452 619 1453 623
rect 1447 618 1453 619
rect 1503 623 1509 624
rect 1503 619 1504 623
rect 1508 622 1509 623
rect 1526 623 1532 624
rect 1526 622 1527 623
rect 1508 620 1527 622
rect 1508 619 1509 620
rect 1503 618 1509 619
rect 1526 619 1527 620
rect 1531 619 1532 623
rect 1526 618 1532 619
rect 1559 623 1565 624
rect 1559 619 1560 623
rect 1564 622 1565 623
rect 1574 623 1580 624
rect 1574 622 1575 623
rect 1564 620 1575 622
rect 1564 619 1565 620
rect 1559 618 1565 619
rect 1574 619 1575 620
rect 1579 619 1580 623
rect 1574 618 1580 619
rect 1615 623 1621 624
rect 1615 619 1616 623
rect 1620 622 1621 623
rect 1638 623 1644 624
rect 1638 622 1639 623
rect 1620 620 1639 622
rect 1620 619 1621 620
rect 1615 618 1621 619
rect 1638 619 1639 620
rect 1643 619 1644 623
rect 1638 618 1644 619
rect 1671 623 1677 624
rect 1671 619 1672 623
rect 1676 622 1677 623
rect 1710 623 1716 624
rect 1710 622 1711 623
rect 1676 620 1711 622
rect 1676 619 1677 620
rect 1671 618 1677 619
rect 1710 619 1711 620
rect 1715 619 1716 623
rect 1710 618 1716 619
rect 1743 623 1749 624
rect 1743 619 1744 623
rect 1748 622 1749 623
rect 1790 623 1796 624
rect 1790 622 1791 623
rect 1748 620 1791 622
rect 1748 619 1749 620
rect 1743 618 1749 619
rect 1790 619 1791 620
rect 1795 619 1796 623
rect 1790 618 1796 619
rect 1823 623 1829 624
rect 1823 619 1824 623
rect 1828 622 1829 623
rect 1870 623 1876 624
rect 1870 622 1871 623
rect 1828 620 1871 622
rect 1828 619 1829 620
rect 1823 618 1829 619
rect 1870 619 1871 620
rect 1875 619 1876 623
rect 1870 618 1876 619
rect 1903 623 1909 624
rect 1903 619 1904 623
rect 1908 622 1909 623
rect 1958 623 1964 624
rect 1958 622 1959 623
rect 1908 620 1959 622
rect 1908 619 1909 620
rect 1903 618 1909 619
rect 1958 619 1959 620
rect 1963 619 1964 623
rect 1968 622 1970 628
rect 1991 623 1997 624
rect 1991 622 1992 623
rect 1968 620 1992 622
rect 1958 618 1964 619
rect 1991 619 1992 620
rect 1996 619 1997 623
rect 1991 618 1997 619
rect 2070 623 2076 624
rect 2070 619 2071 623
rect 2075 622 2076 623
rect 2087 623 2093 624
rect 2087 622 2088 623
rect 2075 620 2088 622
rect 2075 619 2076 620
rect 2070 618 2076 619
rect 2087 619 2088 620
rect 2092 619 2093 623
rect 2087 618 2093 619
rect 2118 620 2124 621
rect 1134 615 1140 616
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 1030 611 1036 612
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1318 612 1324 613
rect 1318 608 1319 612
rect 1323 608 1324 612
rect 1318 607 1324 608
rect 1366 612 1372 613
rect 1366 608 1367 612
rect 1371 608 1372 612
rect 1366 607 1372 608
rect 1422 612 1428 613
rect 1422 608 1423 612
rect 1427 608 1428 612
rect 1422 607 1428 608
rect 1478 612 1484 613
rect 1478 608 1479 612
rect 1483 608 1484 612
rect 1478 607 1484 608
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1646 612 1652 613
rect 1646 608 1647 612
rect 1651 608 1652 612
rect 1646 607 1652 608
rect 1718 612 1724 613
rect 1718 608 1719 612
rect 1723 608 1724 612
rect 1718 607 1724 608
rect 1798 612 1804 613
rect 1798 608 1799 612
rect 1803 608 1804 612
rect 1798 607 1804 608
rect 1878 612 1884 613
rect 1878 608 1879 612
rect 1883 608 1884 612
rect 1878 607 1884 608
rect 1966 612 1972 613
rect 1966 608 1967 612
rect 1971 608 1972 612
rect 1966 607 1972 608
rect 2062 612 2068 613
rect 2062 608 2063 612
rect 2067 608 2068 612
rect 2062 607 2068 608
rect 155 603 161 604
rect 155 599 156 603
rect 160 602 161 603
rect 182 603 188 604
rect 182 602 183 603
rect 160 600 183 602
rect 160 599 161 600
rect 155 598 161 599
rect 182 599 183 600
rect 187 599 188 603
rect 182 598 188 599
rect 206 603 217 604
rect 206 599 207 603
rect 211 599 212 603
rect 216 599 217 603
rect 206 598 217 599
rect 274 603 280 604
rect 274 599 275 603
rect 279 602 280 603
rect 283 603 289 604
rect 283 602 284 603
rect 279 600 284 602
rect 279 599 280 600
rect 274 598 280 599
rect 283 599 284 600
rect 288 599 289 603
rect 283 598 289 599
rect 363 603 369 604
rect 363 599 364 603
rect 368 602 369 603
rect 402 603 408 604
rect 402 602 403 603
rect 368 600 403 602
rect 368 599 369 600
rect 363 598 369 599
rect 402 599 403 600
rect 407 599 408 603
rect 402 598 408 599
rect 451 603 457 604
rect 451 599 452 603
rect 456 602 457 603
rect 487 603 493 604
rect 487 602 488 603
rect 456 600 488 602
rect 456 599 457 600
rect 451 598 457 599
rect 487 599 488 600
rect 492 599 493 603
rect 487 598 493 599
rect 534 603 545 604
rect 534 599 535 603
rect 539 599 540 603
rect 544 599 545 603
rect 534 598 545 599
rect 627 603 633 604
rect 627 599 628 603
rect 632 602 633 603
rect 646 603 652 604
rect 646 602 647 603
rect 632 600 647 602
rect 632 599 633 600
rect 627 598 633 599
rect 646 599 647 600
rect 651 599 652 603
rect 646 598 652 599
rect 715 603 721 604
rect 715 599 716 603
rect 720 602 721 603
rect 726 603 732 604
rect 726 602 727 603
rect 720 600 727 602
rect 720 599 721 600
rect 715 598 721 599
rect 726 599 727 600
rect 731 599 732 603
rect 726 598 732 599
rect 790 603 801 604
rect 790 599 791 603
rect 795 599 796 603
rect 800 599 801 603
rect 790 598 801 599
rect 867 603 873 604
rect 867 599 868 603
rect 872 602 873 603
rect 878 603 884 604
rect 878 602 879 603
rect 872 600 879 602
rect 872 599 873 600
rect 867 598 873 599
rect 878 599 879 600
rect 883 599 884 603
rect 878 598 884 599
rect 942 603 953 604
rect 942 599 943 603
rect 947 599 948 603
rect 952 599 953 603
rect 942 598 953 599
rect 1022 603 1033 604
rect 1022 599 1023 603
rect 1027 599 1028 603
rect 1032 599 1033 603
rect 1022 598 1033 599
rect 1266 599 1272 600
rect 334 595 340 596
rect 334 594 335 595
rect 156 592 335 594
rect 156 590 158 592
rect 334 591 335 592
rect 339 591 340 595
rect 942 595 948 596
rect 942 594 943 595
rect 334 590 340 591
rect 780 592 943 594
rect 780 590 782 592
rect 942 591 943 592
rect 947 591 948 595
rect 1266 595 1267 599
rect 1271 598 1272 599
rect 1275 599 1281 600
rect 1275 598 1276 599
rect 1271 596 1276 598
rect 1271 595 1272 596
rect 1266 594 1272 595
rect 1275 595 1276 596
rect 1280 595 1281 599
rect 1275 594 1281 595
rect 1306 599 1312 600
rect 1306 595 1307 599
rect 1311 598 1312 599
rect 1315 599 1321 600
rect 1315 598 1316 599
rect 1311 596 1316 598
rect 1311 595 1312 596
rect 1306 594 1312 595
rect 1315 595 1316 596
rect 1320 595 1321 599
rect 1315 594 1321 595
rect 1358 599 1369 600
rect 1358 595 1359 599
rect 1363 595 1364 599
rect 1368 595 1369 599
rect 1358 594 1369 595
rect 1406 599 1412 600
rect 1406 595 1407 599
rect 1411 598 1412 599
rect 1419 599 1425 600
rect 1419 598 1420 599
rect 1411 596 1420 598
rect 1411 595 1412 596
rect 1406 594 1412 595
rect 1419 595 1420 596
rect 1424 595 1425 599
rect 1419 594 1425 595
rect 1470 599 1481 600
rect 1470 595 1471 599
rect 1475 595 1476 599
rect 1480 595 1481 599
rect 1470 594 1481 595
rect 1526 599 1537 600
rect 1526 595 1527 599
rect 1531 595 1532 599
rect 1536 595 1537 599
rect 1526 594 1537 595
rect 1587 599 1593 600
rect 1587 595 1588 599
rect 1592 598 1593 599
rect 1630 599 1636 600
rect 1630 598 1631 599
rect 1592 596 1631 598
rect 1592 595 1593 596
rect 1587 594 1593 595
rect 1630 595 1631 596
rect 1635 595 1636 599
rect 1630 594 1636 595
rect 1638 599 1649 600
rect 1638 595 1639 599
rect 1643 595 1644 599
rect 1648 595 1649 599
rect 1638 594 1649 595
rect 1710 599 1721 600
rect 1710 595 1711 599
rect 1715 595 1716 599
rect 1720 595 1721 599
rect 1710 594 1721 595
rect 1790 599 1801 600
rect 1790 595 1791 599
rect 1795 595 1796 599
rect 1800 595 1801 599
rect 1790 594 1801 595
rect 1870 599 1881 600
rect 1870 595 1871 599
rect 1875 595 1876 599
rect 1880 595 1881 599
rect 1870 594 1881 595
rect 1958 599 1969 600
rect 1958 595 1959 599
rect 1963 595 1964 599
rect 1968 595 1969 599
rect 1958 594 1969 595
rect 2050 599 2056 600
rect 2050 595 2051 599
rect 2055 598 2056 599
rect 2059 599 2065 600
rect 2059 598 2060 599
rect 2055 596 2060 598
rect 2055 595 2056 596
rect 2050 594 2056 595
rect 2059 595 2060 596
rect 2064 595 2065 599
rect 2059 594 2065 595
rect 942 590 948 591
rect 155 589 161 590
rect 155 585 156 589
rect 160 585 161 589
rect 779 589 785 590
rect 155 584 161 585
rect 203 587 209 588
rect 203 583 204 587
rect 208 586 209 587
rect 242 587 248 588
rect 242 586 243 587
rect 208 584 243 586
rect 208 583 209 584
rect 203 582 209 583
rect 242 583 243 584
rect 247 583 248 587
rect 242 582 248 583
rect 251 587 257 588
rect 251 583 252 587
rect 256 586 257 587
rect 262 587 268 588
rect 262 586 263 587
rect 256 584 263 586
rect 256 583 257 584
rect 251 582 257 583
rect 262 583 263 584
rect 267 583 268 587
rect 262 582 268 583
rect 307 587 313 588
rect 307 583 308 587
rect 312 586 313 587
rect 379 587 385 588
rect 312 584 321 586
rect 312 583 313 584
rect 307 582 313 583
rect 319 582 321 584
rect 370 583 376 584
rect 370 582 371 583
rect 319 580 371 582
rect 370 579 371 580
rect 375 579 376 583
rect 379 583 380 587
rect 384 586 385 587
rect 390 587 396 588
rect 390 586 391 587
rect 384 584 391 586
rect 384 583 385 584
rect 379 582 385 583
rect 390 583 391 584
rect 395 583 396 587
rect 390 582 396 583
rect 410 587 416 588
rect 410 583 411 587
rect 415 586 416 587
rect 459 587 465 588
rect 459 586 460 587
rect 415 584 460 586
rect 415 583 416 584
rect 410 582 416 583
rect 459 583 460 584
rect 464 583 465 587
rect 459 582 465 583
rect 490 587 496 588
rect 490 583 491 587
rect 495 586 496 587
rect 539 587 545 588
rect 539 586 540 587
rect 495 584 540 586
rect 495 583 496 584
rect 490 582 496 583
rect 539 583 540 584
rect 544 583 545 587
rect 539 582 545 583
rect 619 587 625 588
rect 619 583 620 587
rect 624 586 625 587
rect 682 587 688 588
rect 682 586 683 587
rect 624 584 683 586
rect 624 583 625 584
rect 619 582 625 583
rect 682 583 683 584
rect 687 583 688 587
rect 682 582 688 583
rect 690 587 696 588
rect 690 583 691 587
rect 695 586 696 587
rect 699 587 705 588
rect 699 586 700 587
rect 695 584 700 586
rect 695 583 696 584
rect 690 582 696 583
rect 699 583 700 584
rect 704 583 705 587
rect 779 585 780 589
rect 784 585 785 589
rect 779 584 785 585
rect 810 587 816 588
rect 699 582 705 583
rect 810 583 811 587
rect 815 586 816 587
rect 851 587 857 588
rect 851 586 852 587
rect 815 584 852 586
rect 815 583 816 584
rect 810 582 816 583
rect 851 583 852 584
rect 856 583 857 587
rect 851 582 857 583
rect 923 587 929 588
rect 923 583 924 587
rect 928 586 929 587
rect 986 587 992 588
rect 986 586 987 587
rect 928 584 987 586
rect 928 583 929 584
rect 923 582 929 583
rect 986 583 987 584
rect 991 583 992 587
rect 986 582 992 583
rect 995 587 1001 588
rect 995 583 996 587
rect 1000 586 1001 587
rect 1031 587 1037 588
rect 1031 586 1032 587
rect 1000 584 1032 586
rect 1000 583 1001 584
rect 995 582 1001 583
rect 1031 583 1032 584
rect 1036 583 1037 587
rect 1031 582 1037 583
rect 1043 587 1049 588
rect 1043 583 1044 587
rect 1048 586 1049 587
rect 1070 587 1076 588
rect 1070 586 1071 587
rect 1048 584 1071 586
rect 1048 583 1049 584
rect 1043 582 1049 583
rect 1070 583 1071 584
rect 1075 583 1076 587
rect 1070 582 1076 583
rect 1331 587 1337 588
rect 1331 583 1332 587
rect 1336 586 1337 587
rect 1342 587 1348 588
rect 1342 586 1343 587
rect 1336 584 1343 586
rect 1336 583 1337 584
rect 1331 582 1337 583
rect 1342 583 1343 584
rect 1347 583 1348 587
rect 1342 582 1348 583
rect 1358 587 1364 588
rect 1358 583 1359 587
rect 1363 586 1364 587
rect 1371 587 1377 588
rect 1371 586 1372 587
rect 1363 584 1372 586
rect 1363 583 1364 584
rect 1358 582 1364 583
rect 1371 583 1372 584
rect 1376 583 1377 587
rect 1371 582 1377 583
rect 1402 587 1408 588
rect 1402 583 1403 587
rect 1407 586 1408 587
rect 1411 587 1417 588
rect 1411 586 1412 587
rect 1407 584 1412 586
rect 1407 583 1408 584
rect 1402 582 1408 583
rect 1411 583 1412 584
rect 1416 583 1417 587
rect 1411 582 1417 583
rect 1442 587 1448 588
rect 1442 583 1443 587
rect 1447 586 1448 587
rect 1459 587 1465 588
rect 1459 586 1460 587
rect 1447 584 1460 586
rect 1447 583 1448 584
rect 1442 582 1448 583
rect 1459 583 1460 584
rect 1464 583 1465 587
rect 1459 582 1465 583
rect 1490 587 1496 588
rect 1490 583 1491 587
rect 1495 586 1496 587
rect 1515 587 1521 588
rect 1515 586 1516 587
rect 1495 584 1516 586
rect 1495 583 1496 584
rect 1490 582 1496 583
rect 1515 583 1516 584
rect 1520 583 1521 587
rect 1515 582 1521 583
rect 1574 587 1585 588
rect 1574 583 1575 587
rect 1579 583 1580 587
rect 1584 583 1585 587
rect 1574 582 1585 583
rect 1610 587 1616 588
rect 1610 583 1611 587
rect 1615 586 1616 587
rect 1651 587 1657 588
rect 1651 586 1652 587
rect 1615 584 1652 586
rect 1615 583 1616 584
rect 1610 582 1616 583
rect 1651 583 1652 584
rect 1656 583 1657 587
rect 1651 582 1657 583
rect 1723 587 1729 588
rect 1723 583 1724 587
rect 1728 586 1729 587
rect 1790 587 1796 588
rect 1790 586 1791 587
rect 1728 584 1791 586
rect 1728 583 1729 584
rect 1723 582 1729 583
rect 1790 583 1791 584
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1803 587 1809 588
rect 1803 583 1804 587
rect 1808 586 1809 587
rect 1870 587 1876 588
rect 1870 586 1871 587
rect 1808 584 1871 586
rect 1808 583 1809 584
rect 1803 582 1809 583
rect 1870 583 1871 584
rect 1875 583 1876 587
rect 1883 587 1889 588
rect 1883 584 1884 587
rect 1870 582 1876 583
rect 1878 583 1884 584
rect 1888 583 1889 587
rect 370 578 376 579
rect 1878 579 1879 583
rect 1883 582 1889 583
rect 1971 587 1977 588
rect 1971 583 1972 587
rect 1976 586 1977 587
rect 2050 587 2056 588
rect 2050 586 2051 587
rect 1976 584 2051 586
rect 1976 583 1977 584
rect 1971 582 1977 583
rect 2050 583 2051 584
rect 2055 583 2056 587
rect 2050 582 2056 583
rect 2059 587 2065 588
rect 2059 583 2060 587
rect 2064 586 2065 587
rect 2070 587 2076 588
rect 2070 586 2071 587
rect 2064 584 2071 586
rect 2064 583 2065 584
rect 2059 582 2065 583
rect 2070 583 2071 584
rect 2075 583 2076 587
rect 2070 582 2076 583
rect 1883 580 1887 582
rect 1883 579 1884 580
rect 1878 578 1884 579
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 206 576 212 577
rect 206 572 207 576
rect 211 572 212 576
rect 206 571 212 572
rect 254 576 260 577
rect 254 572 255 576
rect 259 572 260 576
rect 254 571 260 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 462 571 468 572
rect 542 576 548 577
rect 542 572 543 576
rect 547 572 548 576
rect 542 571 548 572
rect 622 576 628 577
rect 622 572 623 576
rect 627 572 628 576
rect 622 571 628 572
rect 702 576 708 577
rect 702 572 703 576
rect 707 572 708 576
rect 702 571 708 572
rect 782 576 788 577
rect 782 572 783 576
rect 787 572 788 576
rect 782 571 788 572
rect 854 576 860 577
rect 854 572 855 576
rect 859 572 860 576
rect 854 571 860 572
rect 926 576 932 577
rect 926 572 927 576
rect 931 572 932 576
rect 926 571 932 572
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1046 576 1052 577
rect 1046 572 1047 576
rect 1051 572 1052 576
rect 1046 571 1052 572
rect 1334 576 1340 577
rect 1334 572 1335 576
rect 1339 572 1340 576
rect 1334 571 1340 572
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1414 576 1420 577
rect 1414 572 1415 576
rect 1419 572 1420 576
rect 1414 571 1420 572
rect 1462 576 1468 577
rect 1462 572 1463 576
rect 1467 572 1468 576
rect 1462 571 1468 572
rect 1518 576 1524 577
rect 1518 572 1519 576
rect 1523 572 1524 576
rect 1518 571 1524 572
rect 1582 576 1588 577
rect 1582 572 1583 576
rect 1587 572 1588 576
rect 1582 571 1588 572
rect 1654 576 1660 577
rect 1654 572 1655 576
rect 1659 572 1660 576
rect 1654 571 1660 572
rect 1726 576 1732 577
rect 1726 572 1727 576
rect 1731 572 1732 576
rect 1726 571 1732 572
rect 1806 576 1812 577
rect 1806 572 1807 576
rect 1811 572 1812 576
rect 1806 571 1812 572
rect 1886 576 1892 577
rect 1886 572 1887 576
rect 1891 572 1892 576
rect 1886 571 1892 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2062 576 2068 577
rect 2062 572 2063 576
rect 2067 572 2068 576
rect 2062 571 2068 572
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 110 563 116 564
rect 182 563 189 564
rect 182 559 183 563
rect 188 559 189 563
rect 182 558 189 559
rect 230 563 237 564
rect 230 559 231 563
rect 236 559 237 563
rect 230 558 237 559
rect 242 563 248 564
rect 242 559 243 563
rect 247 562 248 563
rect 279 563 285 564
rect 279 562 280 563
rect 247 560 280 562
rect 247 559 248 560
rect 242 558 248 559
rect 279 559 280 560
rect 284 559 285 563
rect 279 558 285 559
rect 334 563 341 564
rect 334 559 335 563
rect 340 559 341 563
rect 334 558 341 559
rect 407 563 416 564
rect 407 559 408 563
rect 415 559 416 563
rect 407 558 416 559
rect 487 563 496 564
rect 487 559 488 563
rect 495 559 496 563
rect 487 558 496 559
rect 567 563 573 564
rect 567 559 568 563
rect 572 562 573 563
rect 582 563 588 564
rect 582 562 583 563
rect 572 560 583 562
rect 572 559 573 560
rect 567 558 573 559
rect 582 559 583 560
rect 587 559 588 563
rect 582 558 588 559
rect 646 563 653 564
rect 646 559 647 563
rect 652 559 653 563
rect 646 558 653 559
rect 682 563 688 564
rect 682 559 683 563
rect 687 562 688 563
rect 727 563 733 564
rect 727 562 728 563
rect 687 560 728 562
rect 687 559 688 560
rect 682 558 688 559
rect 727 559 728 560
rect 732 559 733 563
rect 727 558 733 559
rect 807 563 816 564
rect 807 559 808 563
rect 815 559 816 563
rect 807 558 816 559
rect 878 563 885 564
rect 878 559 879 563
rect 884 559 885 563
rect 878 558 885 559
rect 942 563 948 564
rect 942 559 943 563
rect 947 562 948 563
rect 951 563 957 564
rect 951 562 952 563
rect 947 560 952 562
rect 947 559 948 560
rect 942 558 948 559
rect 951 559 952 560
rect 956 559 957 563
rect 951 558 957 559
rect 986 563 992 564
rect 986 559 987 563
rect 991 562 992 563
rect 1023 563 1029 564
rect 1023 562 1024 563
rect 991 560 1024 562
rect 991 559 992 560
rect 986 558 992 559
rect 1023 559 1024 560
rect 1028 559 1029 563
rect 1023 558 1029 559
rect 1031 563 1037 564
rect 1031 559 1032 563
rect 1036 562 1037 563
rect 1071 563 1077 564
rect 1094 563 1100 564
rect 1134 568 1140 569
rect 1672 568 1690 570
rect 1134 564 1135 568
rect 1139 564 1140 568
rect 1630 567 1636 568
rect 1134 563 1140 564
rect 1358 563 1365 564
rect 1071 562 1072 563
rect 1036 560 1072 562
rect 1036 559 1037 560
rect 1031 558 1037 559
rect 1071 559 1072 560
rect 1076 559 1077 563
rect 1071 558 1077 559
rect 1358 559 1359 563
rect 1364 559 1365 563
rect 1358 558 1365 559
rect 1399 563 1408 564
rect 1399 559 1400 563
rect 1407 559 1408 563
rect 1399 558 1408 559
rect 1439 563 1448 564
rect 1439 559 1440 563
rect 1447 559 1448 563
rect 1439 558 1448 559
rect 1487 563 1496 564
rect 1487 559 1488 563
rect 1495 559 1496 563
rect 1487 558 1496 559
rect 1502 563 1508 564
rect 1502 559 1503 563
rect 1507 562 1508 563
rect 1543 563 1549 564
rect 1543 562 1544 563
rect 1507 560 1544 562
rect 1507 559 1508 560
rect 1502 558 1508 559
rect 1543 559 1544 560
rect 1548 559 1549 563
rect 1543 558 1549 559
rect 1607 563 1616 564
rect 1607 559 1608 563
rect 1615 559 1616 563
rect 1630 563 1631 567
rect 1635 566 1636 567
rect 1672 566 1674 568
rect 1635 564 1674 566
rect 1635 563 1636 564
rect 1630 562 1636 563
rect 1678 563 1685 564
rect 1607 558 1616 559
rect 1678 559 1679 563
rect 1684 559 1685 563
rect 1688 562 1690 568
rect 2118 568 2124 569
rect 2118 564 2119 568
rect 2123 564 2124 568
rect 1751 563 1757 564
rect 1751 562 1752 563
rect 1688 560 1752 562
rect 1678 558 1685 559
rect 1751 559 1752 560
rect 1756 559 1757 563
rect 1751 558 1757 559
rect 1790 563 1796 564
rect 1790 559 1791 563
rect 1795 562 1796 563
rect 1831 563 1837 564
rect 1831 562 1832 563
rect 1795 560 1832 562
rect 1795 559 1796 560
rect 1790 558 1796 559
rect 1831 559 1832 560
rect 1836 559 1837 563
rect 1831 558 1837 559
rect 1870 563 1876 564
rect 1870 559 1871 563
rect 1875 562 1876 563
rect 1911 563 1917 564
rect 1911 562 1912 563
rect 1875 560 1912 562
rect 1875 559 1876 560
rect 1870 558 1876 559
rect 1911 559 1912 560
rect 1916 559 1917 563
rect 1911 558 1917 559
rect 1998 563 2005 564
rect 1998 559 1999 563
rect 2004 559 2005 563
rect 1998 558 2005 559
rect 2050 563 2056 564
rect 2050 559 2051 563
rect 2055 562 2056 563
rect 2087 563 2093 564
rect 2118 563 2124 564
rect 2087 562 2088 563
rect 2055 560 2088 562
rect 2055 559 2056 560
rect 2050 558 2056 559
rect 2087 559 2088 560
rect 2092 559 2093 563
rect 2087 558 2093 559
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 1094 551 1100 552
rect 110 546 116 547
rect 158 548 164 549
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 206 548 212 549
rect 206 544 207 548
rect 211 544 212 548
rect 206 543 212 544
rect 254 548 260 549
rect 254 544 255 548
rect 259 544 260 548
rect 254 543 260 544
rect 310 548 316 549
rect 310 544 311 548
rect 315 544 316 548
rect 310 543 316 544
rect 382 548 388 549
rect 382 544 383 548
rect 387 544 388 548
rect 382 543 388 544
rect 462 548 468 549
rect 462 544 463 548
rect 467 544 468 548
rect 462 543 468 544
rect 542 548 548 549
rect 542 544 543 548
rect 547 544 548 548
rect 542 543 548 544
rect 622 548 628 549
rect 622 544 623 548
rect 627 544 628 548
rect 622 543 628 544
rect 702 548 708 549
rect 702 544 703 548
rect 707 544 708 548
rect 702 543 708 544
rect 782 548 788 549
rect 782 544 783 548
rect 787 544 788 548
rect 782 543 788 544
rect 854 548 860 549
rect 854 544 855 548
rect 859 544 860 548
rect 854 543 860 544
rect 926 548 932 549
rect 926 544 927 548
rect 931 544 932 548
rect 926 543 932 544
rect 998 548 1004 549
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1046 548 1052 549
rect 1046 544 1047 548
rect 1051 544 1052 548
rect 1094 547 1095 551
rect 1099 547 1100 551
rect 1094 546 1100 547
rect 1134 551 1140 552
rect 1134 547 1135 551
rect 1139 547 1140 551
rect 2118 551 2124 552
rect 1134 546 1140 547
rect 1334 548 1340 549
rect 1046 543 1052 544
rect 1334 544 1335 548
rect 1339 544 1340 548
rect 1334 543 1340 544
rect 1374 548 1380 549
rect 1374 544 1375 548
rect 1379 544 1380 548
rect 1374 543 1380 544
rect 1414 548 1420 549
rect 1414 544 1415 548
rect 1419 544 1420 548
rect 1414 543 1420 544
rect 1462 548 1468 549
rect 1462 544 1463 548
rect 1467 544 1468 548
rect 1462 543 1468 544
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1582 548 1588 549
rect 1582 544 1583 548
rect 1587 544 1588 548
rect 1582 543 1588 544
rect 1654 548 1660 549
rect 1654 544 1655 548
rect 1659 544 1660 548
rect 1654 543 1660 544
rect 1726 548 1732 549
rect 1726 544 1727 548
rect 1731 544 1732 548
rect 1726 543 1732 544
rect 1806 548 1812 549
rect 1806 544 1807 548
rect 1811 544 1812 548
rect 1806 543 1812 544
rect 1886 548 1892 549
rect 1886 544 1887 548
rect 1891 544 1892 548
rect 1886 543 1892 544
rect 1974 548 1980 549
rect 1974 544 1975 548
rect 1979 544 1980 548
rect 1974 543 1980 544
rect 2062 548 2068 549
rect 2062 544 2063 548
rect 2067 544 2068 548
rect 2118 547 2119 551
rect 2123 547 2124 551
rect 2118 546 2124 547
rect 2062 543 2068 544
rect 1550 539 1556 540
rect 1550 535 1551 539
rect 1555 538 1556 539
rect 1678 539 1684 540
rect 1678 538 1679 539
rect 1555 536 1679 538
rect 1555 535 1556 536
rect 1550 534 1556 535
rect 1678 535 1679 536
rect 1683 535 1684 539
rect 1678 534 1684 535
rect 1190 532 1196 533
rect 1134 529 1140 530
rect 166 528 172 529
rect 110 525 116 526
rect 110 521 111 525
rect 115 521 116 525
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 286 528 292 529
rect 286 524 287 528
rect 291 524 292 528
rect 286 523 292 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 430 528 436 529
rect 430 524 431 528
rect 435 524 436 528
rect 430 523 436 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 590 528 596 529
rect 590 524 591 528
rect 595 524 596 528
rect 590 523 596 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 734 528 740 529
rect 734 524 735 528
rect 739 524 740 528
rect 734 523 740 524
rect 806 528 812 529
rect 806 524 807 528
rect 811 524 812 528
rect 806 523 812 524
rect 870 528 876 529
rect 870 524 871 528
rect 875 524 876 528
rect 870 523 876 524
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 998 528 1004 529
rect 998 524 999 528
rect 1003 524 1004 528
rect 998 523 1004 524
rect 1046 528 1052 529
rect 1046 524 1047 528
rect 1051 524 1052 528
rect 1046 523 1052 524
rect 1094 525 1100 526
rect 110 520 116 521
rect 1094 521 1095 525
rect 1099 521 1100 525
rect 1134 525 1135 529
rect 1139 525 1140 529
rect 1190 528 1191 532
rect 1195 528 1196 532
rect 1190 527 1196 528
rect 1238 532 1244 533
rect 1238 528 1239 532
rect 1243 528 1244 532
rect 1238 527 1244 528
rect 1286 532 1292 533
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1286 527 1292 528
rect 1342 532 1348 533
rect 1342 528 1343 532
rect 1347 528 1348 532
rect 1342 527 1348 528
rect 1406 532 1412 533
rect 1406 528 1407 532
rect 1411 528 1412 532
rect 1406 527 1412 528
rect 1478 532 1484 533
rect 1478 528 1479 532
rect 1483 528 1484 532
rect 1478 527 1484 528
rect 1542 532 1548 533
rect 1542 528 1543 532
rect 1547 528 1548 532
rect 1542 527 1548 528
rect 1606 532 1612 533
rect 1606 528 1607 532
rect 1611 528 1612 532
rect 1606 527 1612 528
rect 1670 532 1676 533
rect 1670 528 1671 532
rect 1675 528 1676 532
rect 1670 527 1676 528
rect 1734 532 1740 533
rect 1734 528 1735 532
rect 1739 528 1740 532
rect 1734 527 1740 528
rect 1798 532 1804 533
rect 1798 528 1799 532
rect 1803 528 1804 532
rect 1798 527 1804 528
rect 1862 532 1868 533
rect 1862 528 1863 532
rect 1867 528 1868 532
rect 1862 527 1868 528
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 1934 527 1940 528
rect 2006 532 2012 533
rect 2006 528 2007 532
rect 2011 528 2012 532
rect 2006 527 2012 528
rect 2070 532 2076 533
rect 2070 528 2071 532
rect 2075 528 2076 532
rect 2070 527 2076 528
rect 2118 529 2124 530
rect 1134 524 1140 525
rect 1888 524 1906 526
rect 2118 525 2119 529
rect 2123 525 2124 529
rect 2118 524 2124 525
rect 1094 520 1100 521
rect 1214 523 1220 524
rect 966 519 972 520
rect 966 515 967 519
rect 971 518 972 519
rect 1206 519 1212 520
rect 1206 518 1207 519
rect 971 516 1207 518
rect 971 515 972 516
rect 966 514 972 515
rect 1206 515 1207 516
rect 1211 515 1212 519
rect 1214 519 1215 523
rect 1219 522 1220 523
rect 1758 523 1764 524
rect 1219 520 1371 522
rect 1219 519 1220 520
rect 1214 518 1220 519
rect 1369 516 1371 520
rect 1758 519 1759 523
rect 1763 522 1764 523
rect 1888 522 1890 524
rect 1763 520 1890 522
rect 1763 519 1764 520
rect 1758 518 1764 519
rect 1887 516 1893 517
rect 1206 514 1212 515
rect 1215 515 1221 516
rect 1134 512 1140 513
rect 174 511 180 512
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 174 507 175 511
rect 179 510 180 511
rect 191 511 197 512
rect 191 510 192 511
rect 179 508 192 510
rect 179 507 180 508
rect 174 506 180 507
rect 191 507 192 508
rect 196 507 197 511
rect 191 506 197 507
rect 199 511 205 512
rect 199 507 200 511
rect 204 510 205 511
rect 247 511 253 512
rect 247 510 248 511
rect 204 508 248 510
rect 204 507 205 508
rect 199 506 205 507
rect 247 507 248 508
rect 252 507 253 511
rect 247 506 253 507
rect 311 511 317 512
rect 311 507 312 511
rect 316 510 317 511
rect 350 511 356 512
rect 350 510 351 511
rect 316 508 351 510
rect 316 507 317 508
rect 311 506 317 507
rect 350 507 351 508
rect 355 507 356 511
rect 350 506 356 507
rect 370 511 376 512
rect 370 507 371 511
rect 375 510 376 511
rect 383 511 389 512
rect 383 510 384 511
rect 375 508 384 510
rect 375 507 376 508
rect 370 506 376 507
rect 383 507 384 508
rect 388 507 389 511
rect 383 506 389 507
rect 394 511 400 512
rect 394 507 395 511
rect 399 510 400 511
rect 455 511 461 512
rect 455 510 456 511
rect 399 508 456 510
rect 399 507 400 508
rect 394 506 400 507
rect 455 507 456 508
rect 460 507 461 511
rect 455 506 461 507
rect 463 511 469 512
rect 463 507 464 511
rect 468 510 469 511
rect 535 511 541 512
rect 535 510 536 511
rect 468 508 536 510
rect 468 507 469 508
rect 463 506 469 507
rect 535 507 536 508
rect 540 507 541 511
rect 535 506 541 507
rect 546 511 552 512
rect 546 507 547 511
rect 551 510 552 511
rect 615 511 621 512
rect 615 510 616 511
rect 551 508 616 510
rect 551 507 552 508
rect 546 506 552 507
rect 615 507 616 508
rect 620 507 621 511
rect 615 506 621 507
rect 687 511 696 512
rect 687 507 688 511
rect 695 507 696 511
rect 687 506 696 507
rect 759 511 765 512
rect 759 507 760 511
rect 764 510 765 511
rect 791 511 797 512
rect 791 510 792 511
rect 764 508 792 510
rect 764 507 765 508
rect 759 506 765 507
rect 791 507 792 508
rect 796 507 797 511
rect 791 506 797 507
rect 831 511 837 512
rect 831 507 832 511
rect 836 510 837 511
rect 862 511 868 512
rect 862 510 863 511
rect 836 508 863 510
rect 836 507 837 508
rect 831 506 837 507
rect 862 507 863 508
rect 867 507 868 511
rect 862 506 868 507
rect 895 511 901 512
rect 895 507 896 511
rect 900 510 901 511
rect 926 511 932 512
rect 926 510 927 511
rect 900 508 927 510
rect 900 507 901 508
rect 895 506 901 507
rect 926 507 927 508
rect 931 507 932 511
rect 926 506 932 507
rect 959 511 965 512
rect 959 507 960 511
rect 964 510 965 511
rect 990 511 996 512
rect 990 510 991 511
rect 964 508 991 510
rect 964 507 965 508
rect 959 506 965 507
rect 990 507 991 508
rect 995 507 996 511
rect 990 506 996 507
rect 1023 511 1029 512
rect 1023 507 1024 511
rect 1028 510 1029 511
rect 1038 511 1044 512
rect 1038 510 1039 511
rect 1028 508 1039 510
rect 1028 507 1029 508
rect 1023 506 1029 507
rect 1038 507 1039 508
rect 1043 507 1044 511
rect 1038 506 1044 507
rect 1070 511 1077 512
rect 1070 507 1071 511
rect 1076 507 1077 511
rect 1070 506 1077 507
rect 1094 508 1100 509
rect 110 503 116 504
rect 1094 504 1095 508
rect 1099 504 1100 508
rect 1134 508 1135 512
rect 1139 508 1140 512
rect 1215 511 1216 515
rect 1220 514 1221 515
rect 1230 515 1236 516
rect 1230 514 1231 515
rect 1220 512 1231 514
rect 1220 511 1221 512
rect 1215 510 1221 511
rect 1230 511 1231 512
rect 1235 511 1236 515
rect 1230 510 1236 511
rect 1263 515 1269 516
rect 1263 511 1264 515
rect 1268 514 1269 515
rect 1278 515 1284 516
rect 1278 514 1279 515
rect 1268 512 1279 514
rect 1268 511 1269 512
rect 1263 510 1269 511
rect 1278 511 1279 512
rect 1283 511 1284 515
rect 1278 510 1284 511
rect 1311 515 1317 516
rect 1311 511 1312 515
rect 1316 514 1317 515
rect 1358 515 1364 516
rect 1358 514 1359 515
rect 1316 512 1359 514
rect 1316 511 1317 512
rect 1311 510 1317 511
rect 1358 511 1359 512
rect 1363 511 1364 515
rect 1358 510 1364 511
rect 1367 515 1373 516
rect 1367 511 1368 515
rect 1372 511 1373 515
rect 1367 510 1373 511
rect 1375 515 1381 516
rect 1375 511 1376 515
rect 1380 514 1381 515
rect 1431 515 1437 516
rect 1431 514 1432 515
rect 1380 512 1432 514
rect 1380 511 1381 512
rect 1375 510 1381 511
rect 1431 511 1432 512
rect 1436 511 1437 515
rect 1431 510 1437 511
rect 1442 515 1448 516
rect 1442 511 1443 515
rect 1447 514 1448 515
rect 1503 515 1509 516
rect 1503 514 1504 515
rect 1447 512 1504 514
rect 1447 511 1448 512
rect 1442 510 1448 511
rect 1503 511 1504 512
rect 1508 511 1509 515
rect 1503 510 1509 511
rect 1567 515 1573 516
rect 1567 511 1568 515
rect 1572 514 1573 515
rect 1590 515 1596 516
rect 1590 514 1591 515
rect 1572 512 1591 514
rect 1572 511 1573 512
rect 1567 510 1573 511
rect 1590 511 1591 512
rect 1595 511 1596 515
rect 1590 510 1596 511
rect 1631 515 1637 516
rect 1631 511 1632 515
rect 1636 514 1637 515
rect 1662 515 1668 516
rect 1662 514 1663 515
rect 1636 512 1663 514
rect 1636 511 1637 512
rect 1631 510 1637 511
rect 1662 511 1663 512
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1694 515 1701 516
rect 1694 511 1695 515
rect 1700 511 1701 515
rect 1694 510 1701 511
rect 1759 515 1765 516
rect 1759 511 1760 515
rect 1764 514 1765 515
rect 1790 515 1796 516
rect 1790 514 1791 515
rect 1764 512 1791 514
rect 1764 511 1765 512
rect 1759 510 1765 511
rect 1790 511 1791 512
rect 1795 511 1796 515
rect 1790 510 1796 511
rect 1823 515 1829 516
rect 1823 511 1824 515
rect 1828 514 1829 515
rect 1854 515 1860 516
rect 1854 514 1855 515
rect 1828 512 1855 514
rect 1828 511 1829 512
rect 1823 510 1829 511
rect 1854 511 1855 512
rect 1859 511 1860 515
rect 1854 510 1860 511
rect 1878 515 1884 516
rect 1878 511 1879 515
rect 1883 514 1884 515
rect 1887 514 1888 516
rect 1883 512 1888 514
rect 1892 512 1893 516
rect 1904 514 1906 524
rect 1959 515 1965 516
rect 1959 514 1960 515
rect 1904 512 1960 514
rect 1883 511 1884 512
rect 1887 511 1893 512
rect 1959 511 1960 512
rect 1964 511 1965 515
rect 1878 510 1884 511
rect 1959 510 1965 511
rect 2031 515 2037 516
rect 2031 511 2032 515
rect 2036 514 2037 515
rect 2062 515 2068 516
rect 2062 514 2063 515
rect 2036 512 2063 514
rect 2036 511 2037 512
rect 2031 510 2037 511
rect 2062 511 2063 512
rect 2067 511 2068 515
rect 2062 510 2068 511
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 514 2084 515
rect 2095 515 2101 516
rect 2095 514 2096 515
rect 2083 512 2096 514
rect 2083 511 2084 512
rect 2078 510 2084 511
rect 2095 511 2096 512
rect 2100 511 2101 515
rect 2095 510 2101 511
rect 2118 512 2124 513
rect 1134 507 1140 508
rect 2118 508 2119 512
rect 2123 508 2124 512
rect 2118 507 2124 508
rect 1094 503 1100 504
rect 1190 504 1196 505
rect 166 500 172 501
rect 166 496 167 500
rect 171 496 172 500
rect 166 495 172 496
rect 222 500 228 501
rect 222 496 223 500
rect 227 496 228 500
rect 222 495 228 496
rect 286 500 292 501
rect 286 496 287 500
rect 291 496 292 500
rect 286 495 292 496
rect 358 500 364 501
rect 358 496 359 500
rect 363 496 364 500
rect 358 495 364 496
rect 430 500 436 501
rect 430 496 431 500
rect 435 496 436 500
rect 430 495 436 496
rect 510 500 516 501
rect 510 496 511 500
rect 515 496 516 500
rect 510 495 516 496
rect 590 500 596 501
rect 590 496 591 500
rect 595 496 596 500
rect 590 495 596 496
rect 662 500 668 501
rect 662 496 663 500
rect 667 496 668 500
rect 662 495 668 496
rect 734 500 740 501
rect 734 496 735 500
rect 739 496 740 500
rect 734 495 740 496
rect 806 500 812 501
rect 806 496 807 500
rect 811 496 812 500
rect 806 495 812 496
rect 870 500 876 501
rect 870 496 871 500
rect 875 496 876 500
rect 870 495 876 496
rect 934 500 940 501
rect 934 496 935 500
rect 939 496 940 500
rect 934 495 940 496
rect 998 500 1004 501
rect 998 496 999 500
rect 1003 496 1004 500
rect 998 495 1004 496
rect 1046 500 1052 501
rect 1046 496 1047 500
rect 1051 496 1052 500
rect 1190 500 1191 504
rect 1195 500 1196 504
rect 1190 499 1196 500
rect 1238 504 1244 505
rect 1238 500 1239 504
rect 1243 500 1244 504
rect 1238 499 1244 500
rect 1286 504 1292 505
rect 1286 500 1287 504
rect 1291 500 1292 504
rect 1286 499 1292 500
rect 1342 504 1348 505
rect 1342 500 1343 504
rect 1347 500 1348 504
rect 1342 499 1348 500
rect 1406 504 1412 505
rect 1406 500 1407 504
rect 1411 500 1412 504
rect 1406 499 1412 500
rect 1478 504 1484 505
rect 1478 500 1479 504
rect 1483 500 1484 504
rect 1478 499 1484 500
rect 1542 504 1548 505
rect 1542 500 1543 504
rect 1547 500 1548 504
rect 1542 499 1548 500
rect 1606 504 1612 505
rect 1606 500 1607 504
rect 1611 500 1612 504
rect 1606 499 1612 500
rect 1670 504 1676 505
rect 1670 500 1671 504
rect 1675 500 1676 504
rect 1670 499 1676 500
rect 1734 504 1740 505
rect 1734 500 1735 504
rect 1739 500 1740 504
rect 1734 499 1740 500
rect 1798 504 1804 505
rect 1798 500 1799 504
rect 1803 500 1804 504
rect 1798 499 1804 500
rect 1862 504 1868 505
rect 1862 500 1863 504
rect 1867 500 1868 504
rect 1862 499 1868 500
rect 1934 504 1940 505
rect 1934 500 1935 504
rect 1939 500 1940 504
rect 1934 499 1940 500
rect 2006 504 2012 505
rect 2006 500 2007 504
rect 2011 500 2012 504
rect 2006 499 2012 500
rect 2070 504 2076 505
rect 2070 500 2071 504
rect 2075 500 2076 504
rect 2070 499 2076 500
rect 1046 495 1052 496
rect 230 491 236 492
rect 230 490 231 491
rect 219 489 231 490
rect 163 487 169 488
rect 163 483 164 487
rect 168 486 169 487
rect 199 487 205 488
rect 199 486 200 487
rect 168 484 200 486
rect 168 483 169 484
rect 163 482 169 483
rect 199 483 200 484
rect 204 483 205 487
rect 219 485 220 489
rect 224 488 231 489
rect 224 485 225 488
rect 230 487 231 488
rect 235 487 236 491
rect 1187 491 1193 492
rect 230 486 236 487
rect 258 487 264 488
rect 219 484 225 485
rect 199 482 205 483
rect 258 483 259 487
rect 263 486 264 487
rect 283 487 289 488
rect 283 486 284 487
rect 263 484 284 486
rect 263 483 264 484
rect 258 482 264 483
rect 283 483 284 484
rect 288 483 289 487
rect 283 482 289 483
rect 350 487 361 488
rect 350 483 351 487
rect 355 483 356 487
rect 360 483 361 487
rect 350 482 361 483
rect 427 487 433 488
rect 427 483 428 487
rect 432 486 433 487
rect 463 487 469 488
rect 463 486 464 487
rect 432 484 464 486
rect 432 483 433 484
rect 427 482 433 483
rect 463 483 464 484
rect 468 483 469 487
rect 463 482 469 483
rect 507 487 513 488
rect 507 483 508 487
rect 512 486 513 487
rect 546 487 552 488
rect 546 486 547 487
rect 512 484 547 486
rect 512 483 513 484
rect 507 482 513 483
rect 546 483 547 484
rect 551 483 552 487
rect 546 482 552 483
rect 582 487 593 488
rect 582 483 583 487
rect 587 483 588 487
rect 592 483 593 487
rect 582 482 593 483
rect 634 487 640 488
rect 634 483 635 487
rect 639 486 640 487
rect 659 487 665 488
rect 659 486 660 487
rect 639 484 660 486
rect 639 483 640 484
rect 634 482 640 483
rect 659 483 660 484
rect 664 483 665 487
rect 659 482 665 483
rect 731 487 737 488
rect 731 483 732 487
rect 736 486 737 487
rect 783 487 789 488
rect 783 486 784 487
rect 736 484 784 486
rect 736 483 737 484
rect 731 482 737 483
rect 783 483 784 484
rect 788 483 789 487
rect 783 482 789 483
rect 791 487 797 488
rect 791 483 792 487
rect 796 486 797 487
rect 803 487 809 488
rect 803 486 804 487
rect 796 484 804 486
rect 796 483 797 484
rect 791 482 797 483
rect 803 483 804 484
rect 808 483 809 487
rect 803 482 809 483
rect 862 487 873 488
rect 862 483 863 487
rect 867 483 868 487
rect 872 483 873 487
rect 862 482 873 483
rect 926 487 937 488
rect 926 483 927 487
rect 931 483 932 487
rect 936 483 937 487
rect 926 482 937 483
rect 990 487 1001 488
rect 990 483 991 487
rect 995 483 996 487
rect 1000 483 1001 487
rect 990 482 1001 483
rect 1038 487 1049 488
rect 1038 483 1039 487
rect 1043 483 1044 487
rect 1048 483 1049 487
rect 1187 487 1188 491
rect 1192 490 1193 491
rect 1214 491 1220 492
rect 1214 490 1215 491
rect 1192 488 1215 490
rect 1192 487 1193 488
rect 1187 486 1193 487
rect 1214 487 1215 488
rect 1219 487 1220 491
rect 1214 486 1220 487
rect 1230 491 1241 492
rect 1230 487 1231 491
rect 1235 487 1236 491
rect 1240 487 1241 491
rect 1230 486 1241 487
rect 1278 491 1289 492
rect 1278 487 1279 491
rect 1283 487 1284 491
rect 1288 487 1289 491
rect 1278 486 1289 487
rect 1339 491 1345 492
rect 1339 487 1340 491
rect 1344 490 1345 491
rect 1375 491 1381 492
rect 1375 490 1376 491
rect 1344 488 1376 490
rect 1344 487 1345 488
rect 1339 486 1345 487
rect 1375 487 1376 488
rect 1380 487 1381 491
rect 1375 486 1381 487
rect 1403 491 1409 492
rect 1403 487 1404 491
rect 1408 490 1409 491
rect 1442 491 1448 492
rect 1442 490 1443 491
rect 1408 488 1443 490
rect 1408 487 1409 488
rect 1403 486 1409 487
rect 1442 487 1443 488
rect 1447 487 1448 491
rect 1442 486 1448 487
rect 1475 491 1481 492
rect 1475 487 1476 491
rect 1480 490 1481 491
rect 1502 491 1508 492
rect 1502 490 1503 491
rect 1480 488 1503 490
rect 1480 487 1481 488
rect 1475 486 1481 487
rect 1502 487 1503 488
rect 1507 487 1508 491
rect 1502 486 1508 487
rect 1539 491 1545 492
rect 1539 487 1540 491
rect 1544 490 1545 491
rect 1550 491 1556 492
rect 1550 490 1551 491
rect 1544 488 1551 490
rect 1544 487 1545 488
rect 1539 486 1545 487
rect 1550 487 1551 488
rect 1555 487 1556 491
rect 1550 486 1556 487
rect 1590 491 1596 492
rect 1590 487 1591 491
rect 1595 490 1596 491
rect 1603 491 1609 492
rect 1603 490 1604 491
rect 1595 488 1604 490
rect 1595 487 1596 488
rect 1590 486 1596 487
rect 1603 487 1604 488
rect 1608 487 1609 491
rect 1603 486 1609 487
rect 1662 491 1673 492
rect 1662 487 1663 491
rect 1667 487 1668 491
rect 1672 487 1673 491
rect 1662 486 1673 487
rect 1731 491 1737 492
rect 1731 487 1732 491
rect 1736 490 1737 491
rect 1758 491 1764 492
rect 1758 490 1759 491
rect 1736 488 1759 490
rect 1736 487 1737 488
rect 1731 486 1737 487
rect 1758 487 1759 488
rect 1763 487 1764 491
rect 1758 486 1764 487
rect 1790 491 1801 492
rect 1790 487 1791 491
rect 1795 487 1796 491
rect 1800 487 1801 491
rect 1790 486 1801 487
rect 1854 491 1865 492
rect 1854 487 1855 491
rect 1859 487 1860 491
rect 1864 487 1865 491
rect 1854 486 1865 487
rect 1931 491 1937 492
rect 1931 487 1932 491
rect 1936 490 1937 491
rect 1966 491 1972 492
rect 1966 490 1967 491
rect 1936 488 1967 490
rect 1936 487 1937 488
rect 1931 486 1937 487
rect 1966 487 1967 488
rect 1971 487 1972 491
rect 1966 486 1972 487
rect 1998 491 2009 492
rect 1998 487 1999 491
rect 2003 487 2004 491
rect 2008 487 2009 491
rect 1998 486 2009 487
rect 2062 491 2073 492
rect 2062 487 2063 491
rect 2067 487 2068 491
rect 2072 487 2073 491
rect 2062 486 2073 487
rect 1038 482 1049 483
rect 1074 479 1080 480
rect 163 475 169 476
rect 163 471 164 475
rect 168 474 169 475
rect 174 475 180 476
rect 174 474 175 475
rect 168 472 175 474
rect 168 471 169 472
rect 163 470 169 471
rect 174 471 175 472
rect 179 471 180 475
rect 174 470 180 471
rect 227 475 233 476
rect 227 471 228 475
rect 232 474 233 475
rect 271 475 277 476
rect 271 474 272 475
rect 232 472 272 474
rect 232 471 233 472
rect 227 470 233 471
rect 271 471 272 472
rect 276 471 277 475
rect 271 470 277 471
rect 294 475 305 476
rect 294 471 295 475
rect 299 471 300 475
rect 304 471 305 475
rect 294 470 305 471
rect 371 475 377 476
rect 371 471 372 475
rect 376 474 377 475
rect 394 475 400 476
rect 394 474 395 475
rect 376 472 395 474
rect 376 471 377 472
rect 371 470 377 471
rect 394 471 395 472
rect 399 471 400 475
rect 394 470 400 471
rect 402 475 408 476
rect 402 471 403 475
rect 407 474 408 475
rect 451 475 457 476
rect 451 474 452 475
rect 407 472 452 474
rect 407 471 408 472
rect 402 470 408 471
rect 451 471 452 472
rect 456 471 457 475
rect 451 470 457 471
rect 482 475 488 476
rect 482 471 483 475
rect 487 474 488 475
rect 531 475 537 476
rect 531 474 532 475
rect 487 472 532 474
rect 487 471 488 472
rect 482 470 488 471
rect 531 471 532 472
rect 536 471 537 475
rect 531 470 537 471
rect 578 475 584 476
rect 578 471 579 475
rect 583 474 584 475
rect 603 475 609 476
rect 603 474 604 475
rect 583 472 604 474
rect 583 471 584 472
rect 578 470 584 471
rect 603 471 604 472
rect 608 471 609 475
rect 603 470 609 471
rect 675 475 681 476
rect 675 471 676 475
rect 680 474 681 475
rect 698 475 704 476
rect 698 474 699 475
rect 680 472 699 474
rect 680 471 681 472
rect 675 470 681 471
rect 698 471 699 472
rect 703 471 704 475
rect 698 470 704 471
rect 706 475 712 476
rect 706 471 707 475
rect 711 474 712 475
rect 739 475 745 476
rect 739 474 740 475
rect 711 472 740 474
rect 711 471 712 472
rect 706 470 712 471
rect 739 471 740 472
rect 744 471 745 475
rect 739 470 745 471
rect 770 475 776 476
rect 770 471 771 475
rect 775 474 776 475
rect 795 475 801 476
rect 795 474 796 475
rect 775 472 796 474
rect 775 471 776 472
rect 770 470 776 471
rect 795 471 796 472
rect 800 471 801 475
rect 795 470 801 471
rect 826 475 832 476
rect 826 471 827 475
rect 831 474 832 475
rect 851 475 857 476
rect 851 474 852 475
rect 831 472 852 474
rect 831 471 832 472
rect 826 470 832 471
rect 851 471 852 472
rect 856 471 857 475
rect 851 470 857 471
rect 882 475 888 476
rect 882 471 883 475
rect 887 474 888 475
rect 899 475 905 476
rect 899 474 900 475
rect 887 472 900 474
rect 887 471 888 472
rect 882 470 888 471
rect 899 471 900 472
rect 904 471 905 475
rect 899 470 905 471
rect 955 475 961 476
rect 955 471 956 475
rect 960 474 961 475
rect 966 475 972 476
rect 966 474 967 475
rect 960 472 967 474
rect 960 471 961 472
rect 955 470 961 471
rect 966 471 967 472
rect 971 471 972 475
rect 966 470 972 471
rect 986 475 992 476
rect 986 471 987 475
rect 991 474 992 475
rect 1003 475 1009 476
rect 1003 474 1004 475
rect 991 472 1004 474
rect 991 471 992 472
rect 986 470 992 471
rect 1003 471 1004 472
rect 1008 471 1009 475
rect 1003 470 1009 471
rect 1034 475 1040 476
rect 1034 471 1035 475
rect 1039 474 1040 475
rect 1043 475 1049 476
rect 1043 474 1044 475
rect 1039 472 1044 474
rect 1039 471 1040 472
rect 1034 470 1040 471
rect 1043 471 1044 472
rect 1048 471 1049 475
rect 1074 475 1075 479
rect 1079 478 1080 479
rect 1155 479 1161 480
rect 1155 478 1156 479
rect 1079 476 1156 478
rect 1079 475 1080 476
rect 1074 474 1080 475
rect 1155 475 1156 476
rect 1160 475 1161 479
rect 1155 474 1161 475
rect 1259 479 1265 480
rect 1259 475 1260 479
rect 1264 478 1265 479
rect 1350 479 1356 480
rect 1350 478 1351 479
rect 1264 476 1351 478
rect 1264 475 1265 476
rect 1259 474 1265 475
rect 1350 475 1351 476
rect 1355 475 1356 479
rect 1350 474 1356 475
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 478 1364 479
rect 1379 479 1385 480
rect 1379 478 1380 479
rect 1363 476 1380 478
rect 1363 475 1364 476
rect 1358 474 1364 475
rect 1379 475 1380 476
rect 1384 475 1385 479
rect 1379 474 1385 475
rect 1491 479 1497 480
rect 1491 475 1492 479
rect 1496 478 1497 479
rect 1586 479 1592 480
rect 1586 478 1587 479
rect 1496 476 1587 478
rect 1496 475 1497 476
rect 1491 474 1497 475
rect 1586 475 1587 476
rect 1591 475 1592 479
rect 1586 474 1592 475
rect 1595 479 1601 480
rect 1595 475 1596 479
rect 1600 478 1601 479
rect 1686 479 1692 480
rect 1686 478 1687 479
rect 1600 476 1687 478
rect 1600 475 1601 476
rect 1595 474 1601 475
rect 1686 475 1687 476
rect 1691 475 1692 479
rect 1686 474 1692 475
rect 1694 479 1705 480
rect 1694 475 1695 479
rect 1699 475 1700 479
rect 1704 475 1705 479
rect 1694 474 1705 475
rect 1795 479 1801 480
rect 1795 475 1796 479
rect 1800 478 1801 479
rect 1826 479 1832 480
rect 1800 476 1822 478
rect 1800 475 1801 476
rect 1795 474 1801 475
rect 1043 470 1049 471
rect 1820 470 1822 476
rect 1826 475 1827 479
rect 1831 478 1832 479
rect 1883 479 1889 480
rect 1883 478 1884 479
rect 1831 476 1884 478
rect 1831 475 1832 476
rect 1826 474 1832 475
rect 1883 475 1884 476
rect 1888 475 1889 479
rect 1883 474 1889 475
rect 1914 479 1920 480
rect 1914 475 1915 479
rect 1919 478 1920 479
rect 1979 479 1985 480
rect 1979 478 1980 479
rect 1919 476 1980 478
rect 1919 475 1920 476
rect 1914 474 1920 475
rect 1979 475 1980 476
rect 1984 475 1985 479
rect 1979 474 1985 475
rect 2067 479 2073 480
rect 2067 475 2068 479
rect 2072 478 2073 479
rect 2078 479 2084 480
rect 2078 478 2079 479
rect 2072 476 2079 478
rect 2072 475 2073 476
rect 2067 474 2073 475
rect 2078 475 2079 476
rect 2083 475 2084 479
rect 2078 474 2084 475
rect 1846 471 1852 472
rect 1846 470 1847 471
rect 1158 468 1164 469
rect 166 464 172 465
rect 166 460 167 464
rect 171 460 172 464
rect 166 459 172 460
rect 230 464 236 465
rect 230 460 231 464
rect 235 460 236 464
rect 230 459 236 460
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 374 464 380 465
rect 374 460 375 464
rect 379 460 380 464
rect 374 459 380 460
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 534 464 540 465
rect 534 460 535 464
rect 539 460 540 464
rect 534 459 540 460
rect 606 464 612 465
rect 606 460 607 464
rect 611 460 612 464
rect 606 459 612 460
rect 678 464 684 465
rect 678 460 679 464
rect 683 460 684 464
rect 678 459 684 460
rect 742 464 748 465
rect 742 460 743 464
rect 747 460 748 464
rect 742 459 748 460
rect 798 464 804 465
rect 798 460 799 464
rect 803 460 804 464
rect 798 459 804 460
rect 854 464 860 465
rect 854 460 855 464
rect 859 460 860 464
rect 854 459 860 460
rect 902 464 908 465
rect 902 460 903 464
rect 907 460 908 464
rect 902 459 908 460
rect 958 464 964 465
rect 958 460 959 464
rect 963 460 964 464
rect 958 459 964 460
rect 1006 464 1012 465
rect 1006 460 1007 464
rect 1011 460 1012 464
rect 1006 459 1012 460
rect 1046 464 1052 465
rect 1046 460 1047 464
rect 1051 460 1052 464
rect 1158 464 1159 468
rect 1163 464 1164 468
rect 1158 463 1164 464
rect 1262 468 1268 469
rect 1262 464 1263 468
rect 1267 464 1268 468
rect 1262 463 1268 464
rect 1382 468 1388 469
rect 1382 464 1383 468
rect 1387 464 1388 468
rect 1382 463 1388 464
rect 1494 468 1500 469
rect 1494 464 1495 468
rect 1499 464 1500 468
rect 1494 463 1500 464
rect 1598 468 1604 469
rect 1598 464 1599 468
rect 1603 464 1604 468
rect 1598 463 1604 464
rect 1702 468 1708 469
rect 1702 464 1703 468
rect 1707 464 1708 468
rect 1702 463 1708 464
rect 1798 468 1804 469
rect 1820 468 1847 470
rect 1798 464 1799 468
rect 1803 464 1804 468
rect 1846 467 1847 468
rect 1851 467 1852 471
rect 1846 466 1852 467
rect 1886 468 1892 469
rect 1798 463 1804 464
rect 1886 464 1887 468
rect 1891 464 1892 468
rect 1886 463 1892 464
rect 1982 468 1988 469
rect 1982 464 1983 468
rect 1987 464 1988 468
rect 1982 463 1988 464
rect 2070 468 2076 469
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 1046 459 1052 460
rect 1134 460 1140 461
rect 110 456 116 457
rect 817 456 850 458
rect 110 452 111 456
rect 115 452 116 456
rect 783 455 789 456
rect 110 451 116 452
rect 158 451 164 452
rect 158 447 159 451
rect 163 450 164 451
rect 191 451 197 452
rect 191 450 192 451
rect 163 448 192 450
rect 163 447 164 448
rect 158 446 164 447
rect 191 447 192 448
rect 196 447 197 451
rect 191 446 197 447
rect 255 451 264 452
rect 255 447 256 451
rect 263 447 264 451
rect 255 446 264 447
rect 271 451 277 452
rect 271 447 272 451
rect 276 450 277 451
rect 327 451 333 452
rect 327 450 328 451
rect 276 448 328 450
rect 276 447 277 448
rect 271 446 277 447
rect 327 447 328 448
rect 332 447 333 451
rect 327 446 333 447
rect 399 451 408 452
rect 399 447 400 451
rect 407 447 408 451
rect 399 446 408 447
rect 479 451 488 452
rect 479 447 480 451
rect 487 447 488 451
rect 479 446 488 447
rect 494 451 500 452
rect 494 447 495 451
rect 499 450 500 451
rect 559 451 565 452
rect 559 450 560 451
rect 499 448 560 450
rect 499 447 500 448
rect 494 446 500 447
rect 559 447 560 448
rect 564 447 565 451
rect 559 446 565 447
rect 631 451 640 452
rect 631 447 632 451
rect 639 447 640 451
rect 631 446 640 447
rect 703 451 712 452
rect 703 447 704 451
rect 711 447 712 451
rect 703 446 712 447
rect 767 451 776 452
rect 767 447 768 451
rect 775 447 776 451
rect 783 451 784 455
rect 788 454 789 455
rect 817 454 819 456
rect 788 452 819 454
rect 848 454 850 456
rect 872 456 894 458
rect 872 454 874 456
rect 848 452 874 454
rect 788 451 789 452
rect 783 450 789 451
rect 823 451 832 452
rect 767 446 776 447
rect 823 447 824 451
rect 831 447 832 451
rect 823 446 832 447
rect 879 451 888 452
rect 879 447 880 451
rect 887 447 888 451
rect 892 450 894 456
rect 1094 456 1100 457
rect 1094 452 1095 456
rect 1099 452 1100 456
rect 1134 456 1135 460
rect 1139 456 1140 460
rect 2118 460 2124 461
rect 2118 456 2119 460
rect 2123 456 2124 460
rect 1134 455 1140 456
rect 1166 455 1172 456
rect 927 451 933 452
rect 927 450 928 451
rect 892 448 928 450
rect 879 446 888 447
rect 927 447 928 448
rect 932 447 933 451
rect 927 446 933 447
rect 983 451 992 452
rect 983 447 984 451
rect 991 447 992 451
rect 983 446 992 447
rect 1031 451 1040 452
rect 1031 447 1032 451
rect 1039 447 1040 451
rect 1031 446 1040 447
rect 1071 451 1080 452
rect 1094 451 1100 452
rect 1166 451 1167 455
rect 1171 454 1172 455
rect 1183 455 1189 456
rect 1183 454 1184 455
rect 1171 452 1184 454
rect 1171 451 1172 452
rect 1071 447 1072 451
rect 1079 447 1080 451
rect 1166 450 1172 451
rect 1183 451 1184 452
rect 1188 451 1189 455
rect 1183 450 1189 451
rect 1206 455 1212 456
rect 1206 451 1207 455
rect 1211 454 1212 455
rect 1287 455 1293 456
rect 1287 454 1288 455
rect 1211 452 1288 454
rect 1211 451 1212 452
rect 1206 450 1212 451
rect 1287 451 1288 452
rect 1292 451 1293 455
rect 1287 450 1293 451
rect 1350 455 1356 456
rect 1350 451 1351 455
rect 1355 454 1356 455
rect 1407 455 1413 456
rect 1407 454 1408 455
rect 1355 452 1408 454
rect 1355 451 1356 452
rect 1350 450 1356 451
rect 1407 451 1408 452
rect 1412 451 1413 455
rect 1407 450 1413 451
rect 1519 455 1525 456
rect 1519 451 1520 455
rect 1524 454 1525 455
rect 1582 455 1588 456
rect 1582 454 1583 455
rect 1524 452 1583 454
rect 1524 451 1525 452
rect 1519 450 1525 451
rect 1582 451 1583 452
rect 1587 451 1588 455
rect 1582 450 1588 451
rect 1590 455 1596 456
rect 1590 451 1591 455
rect 1595 454 1596 455
rect 1623 455 1629 456
rect 1623 454 1624 455
rect 1595 452 1624 454
rect 1595 451 1596 452
rect 1590 450 1596 451
rect 1623 451 1624 452
rect 1628 451 1629 455
rect 1623 450 1629 451
rect 1686 455 1692 456
rect 1686 451 1687 455
rect 1691 454 1692 455
rect 1727 455 1733 456
rect 1727 454 1728 455
rect 1691 452 1728 454
rect 1691 451 1692 452
rect 1686 450 1692 451
rect 1727 451 1728 452
rect 1732 451 1733 455
rect 1727 450 1733 451
rect 1823 455 1832 456
rect 1823 451 1824 455
rect 1831 451 1832 455
rect 1823 450 1832 451
rect 1911 455 1920 456
rect 1911 451 1912 455
rect 1919 451 1920 455
rect 1911 450 1920 451
rect 1966 455 1972 456
rect 1966 451 1967 455
rect 1971 454 1972 455
rect 2007 455 2013 456
rect 2007 454 2008 455
rect 1971 452 2008 454
rect 1971 451 1972 452
rect 1966 450 1972 451
rect 2007 451 2008 452
rect 2012 451 2013 455
rect 2007 450 2013 451
rect 2030 455 2036 456
rect 2030 451 2031 455
rect 2035 454 2036 455
rect 2095 455 2101 456
rect 2118 455 2124 456
rect 2095 454 2096 455
rect 2035 452 2096 454
rect 2035 451 2036 452
rect 2030 450 2036 451
rect 2095 451 2096 452
rect 2100 451 2101 455
rect 2095 450 2101 451
rect 1071 446 1080 447
rect 1134 443 1140 444
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 1094 439 1100 440
rect 110 434 116 435
rect 166 436 172 437
rect 166 432 167 436
rect 171 432 172 436
rect 166 431 172 432
rect 230 436 236 437
rect 230 432 231 436
rect 235 432 236 436
rect 230 431 236 432
rect 302 436 308 437
rect 302 432 303 436
rect 307 432 308 436
rect 302 431 308 432
rect 374 436 380 437
rect 374 432 375 436
rect 379 432 380 436
rect 374 431 380 432
rect 454 436 460 437
rect 454 432 455 436
rect 459 432 460 436
rect 454 431 460 432
rect 534 436 540 437
rect 534 432 535 436
rect 539 432 540 436
rect 534 431 540 432
rect 606 436 612 437
rect 606 432 607 436
rect 611 432 612 436
rect 606 431 612 432
rect 678 436 684 437
rect 678 432 679 436
rect 683 432 684 436
rect 678 431 684 432
rect 742 436 748 437
rect 742 432 743 436
rect 747 432 748 436
rect 742 431 748 432
rect 798 436 804 437
rect 798 432 799 436
rect 803 432 804 436
rect 798 431 804 432
rect 854 436 860 437
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 902 436 908 437
rect 902 432 903 436
rect 907 432 908 436
rect 902 431 908 432
rect 958 436 964 437
rect 958 432 959 436
rect 963 432 964 436
rect 958 431 964 432
rect 1006 436 1012 437
rect 1006 432 1007 436
rect 1011 432 1012 436
rect 1006 431 1012 432
rect 1046 436 1052 437
rect 1046 432 1047 436
rect 1051 432 1052 436
rect 1094 435 1095 439
rect 1099 435 1100 439
rect 1134 439 1135 443
rect 1139 439 1140 443
rect 2118 443 2124 444
rect 1134 438 1140 439
rect 1158 440 1164 441
rect 1158 436 1159 440
rect 1163 436 1164 440
rect 1158 435 1164 436
rect 1262 440 1268 441
rect 1262 436 1263 440
rect 1267 436 1268 440
rect 1262 435 1268 436
rect 1382 440 1388 441
rect 1382 436 1383 440
rect 1387 436 1388 440
rect 1382 435 1388 436
rect 1494 440 1500 441
rect 1494 436 1495 440
rect 1499 436 1500 440
rect 1494 435 1500 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1702 440 1708 441
rect 1702 436 1703 440
rect 1707 436 1708 440
rect 1702 435 1708 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1886 440 1892 441
rect 1886 436 1887 440
rect 1891 436 1892 440
rect 1886 435 1892 436
rect 1982 440 1988 441
rect 1982 436 1983 440
rect 1987 436 1988 440
rect 1982 435 1988 436
rect 2070 440 2076 441
rect 2070 436 2071 440
rect 2075 436 2076 440
rect 2118 439 2119 443
rect 2123 439 2124 443
rect 2118 438 2124 439
rect 2070 435 2076 436
rect 1094 434 1100 435
rect 1046 431 1052 432
rect 1158 428 1164 429
rect 1134 425 1140 426
rect 150 424 156 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 150 420 151 424
rect 155 420 156 424
rect 150 419 156 420
rect 214 424 220 425
rect 214 420 215 424
rect 219 420 220 424
rect 214 419 220 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 350 424 356 425
rect 350 420 351 424
rect 355 420 356 424
rect 350 419 356 420
rect 422 424 428 425
rect 422 420 423 424
rect 427 420 428 424
rect 422 419 428 420
rect 486 424 492 425
rect 486 420 487 424
rect 491 420 492 424
rect 486 419 492 420
rect 550 424 556 425
rect 550 420 551 424
rect 555 420 556 424
rect 550 419 556 420
rect 614 424 620 425
rect 614 420 615 424
rect 619 420 620 424
rect 614 419 620 420
rect 670 424 676 425
rect 670 420 671 424
rect 675 420 676 424
rect 670 419 676 420
rect 726 424 732 425
rect 726 420 727 424
rect 731 420 732 424
rect 726 419 732 420
rect 790 424 796 425
rect 790 420 791 424
rect 795 420 796 424
rect 790 419 796 420
rect 854 424 860 425
rect 854 420 855 424
rect 859 420 860 424
rect 854 419 860 420
rect 1094 421 1100 422
rect 110 416 116 417
rect 1094 417 1095 421
rect 1099 417 1100 421
rect 1134 421 1135 425
rect 1139 421 1140 425
rect 1158 424 1159 428
rect 1163 424 1164 428
rect 1158 423 1164 424
rect 1198 428 1204 429
rect 1198 424 1199 428
rect 1203 424 1204 428
rect 1198 423 1204 424
rect 1254 428 1260 429
rect 1254 424 1255 428
rect 1259 424 1260 428
rect 1254 423 1260 424
rect 1334 428 1340 429
rect 1334 424 1335 428
rect 1339 424 1340 428
rect 1334 423 1340 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1502 428 1508 429
rect 1502 424 1503 428
rect 1507 424 1508 428
rect 1502 423 1508 424
rect 1590 428 1596 429
rect 1590 424 1591 428
rect 1595 424 1596 428
rect 1590 423 1596 424
rect 1670 428 1676 429
rect 1670 424 1671 428
rect 1675 424 1676 428
rect 1670 423 1676 424
rect 1750 428 1756 429
rect 1750 424 1751 428
rect 1755 424 1756 428
rect 1750 423 1756 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1822 423 1828 424
rect 1886 428 1892 429
rect 1886 424 1887 428
rect 1891 424 1892 428
rect 1886 423 1892 424
rect 1950 428 1956 429
rect 1950 424 1951 428
rect 1955 424 1956 428
rect 1950 423 1956 424
rect 2022 428 2028 429
rect 2022 424 2023 428
rect 2027 424 2028 428
rect 2022 423 2028 424
rect 2070 428 2076 429
rect 2070 424 2071 428
rect 2075 424 2076 428
rect 2070 423 2076 424
rect 2118 425 2124 426
rect 1134 420 1140 421
rect 2118 421 2119 425
rect 2123 421 2124 425
rect 2118 420 2124 421
rect 1094 416 1100 417
rect 698 415 704 416
rect 698 411 699 415
rect 703 414 704 415
rect 703 412 858 414
rect 703 411 704 412
rect 698 410 704 411
rect 175 407 181 408
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 175 403 176 407
rect 180 406 181 407
rect 206 407 212 408
rect 206 406 207 407
rect 180 404 207 406
rect 180 403 181 404
rect 175 402 181 403
rect 206 403 207 404
rect 211 403 212 407
rect 206 402 212 403
rect 239 407 245 408
rect 239 403 240 407
rect 244 406 245 407
rect 263 407 269 408
rect 263 406 264 407
rect 244 404 264 406
rect 244 403 245 404
rect 239 402 245 403
rect 263 403 264 404
rect 268 403 269 407
rect 263 402 269 403
rect 294 407 300 408
rect 294 403 295 407
rect 299 406 300 407
rect 303 407 309 408
rect 303 406 304 407
rect 299 404 304 406
rect 299 403 300 404
rect 294 402 300 403
rect 303 403 304 404
rect 308 403 309 407
rect 303 402 309 403
rect 375 407 381 408
rect 375 403 376 407
rect 380 406 381 407
rect 390 407 396 408
rect 390 406 391 407
rect 380 404 391 406
rect 380 403 381 404
rect 375 402 381 403
rect 390 403 391 404
rect 395 403 396 407
rect 390 402 396 403
rect 399 407 405 408
rect 399 403 400 407
rect 404 406 405 407
rect 447 407 453 408
rect 447 406 448 407
rect 404 404 448 406
rect 404 403 405 404
rect 399 402 405 403
rect 447 403 448 404
rect 452 403 453 407
rect 447 402 453 403
rect 455 407 461 408
rect 455 403 456 407
rect 460 406 461 407
rect 511 407 517 408
rect 511 406 512 407
rect 460 404 512 406
rect 460 403 461 404
rect 455 402 461 403
rect 511 403 512 404
rect 516 403 517 407
rect 511 402 517 403
rect 575 407 584 408
rect 575 403 576 407
rect 583 403 584 407
rect 575 402 584 403
rect 639 407 645 408
rect 639 403 640 407
rect 644 406 645 407
rect 662 407 668 408
rect 662 406 663 407
rect 644 404 663 406
rect 644 403 645 404
rect 639 402 645 403
rect 662 403 663 404
rect 667 403 668 407
rect 662 402 668 403
rect 695 407 701 408
rect 695 403 696 407
rect 700 406 701 407
rect 718 407 724 408
rect 718 406 719 407
rect 700 404 719 406
rect 700 403 701 404
rect 695 402 701 403
rect 718 403 719 404
rect 723 403 724 407
rect 718 402 724 403
rect 751 407 757 408
rect 751 403 752 407
rect 756 406 757 407
rect 782 407 788 408
rect 782 406 783 407
rect 756 404 783 406
rect 756 403 757 404
rect 751 402 757 403
rect 782 403 783 404
rect 787 403 788 407
rect 782 402 788 403
rect 815 407 821 408
rect 815 403 816 407
rect 820 406 821 407
rect 846 407 852 408
rect 846 406 847 407
rect 820 404 847 406
rect 820 403 821 404
rect 815 402 821 403
rect 846 403 847 404
rect 851 403 852 407
rect 856 406 858 412
rect 1183 411 1192 412
rect 1134 408 1140 409
rect 879 407 885 408
rect 879 406 880 407
rect 856 404 880 406
rect 846 402 852 403
rect 879 403 880 404
rect 884 403 885 407
rect 879 402 885 403
rect 1094 404 1100 405
rect 110 399 116 400
rect 1094 400 1095 404
rect 1099 400 1100 404
rect 1134 404 1135 408
rect 1139 404 1140 408
rect 1183 407 1184 411
rect 1191 407 1192 411
rect 1183 406 1192 407
rect 1223 411 1229 412
rect 1223 407 1224 411
rect 1228 410 1229 411
rect 1246 411 1252 412
rect 1246 410 1247 411
rect 1228 408 1247 410
rect 1228 407 1229 408
rect 1223 406 1229 407
rect 1246 407 1247 408
rect 1251 407 1252 411
rect 1246 406 1252 407
rect 1279 411 1285 412
rect 1279 407 1280 411
rect 1284 410 1285 411
rect 1326 411 1332 412
rect 1326 410 1327 411
rect 1284 408 1327 410
rect 1284 407 1285 408
rect 1279 406 1285 407
rect 1326 407 1327 408
rect 1331 407 1332 411
rect 1326 406 1332 407
rect 1359 411 1365 412
rect 1359 407 1360 411
rect 1364 410 1365 411
rect 1406 411 1412 412
rect 1406 410 1407 411
rect 1364 408 1407 410
rect 1364 407 1365 408
rect 1359 406 1365 407
rect 1406 407 1407 408
rect 1411 407 1412 411
rect 1406 406 1412 407
rect 1439 411 1445 412
rect 1439 407 1440 411
rect 1444 410 1445 411
rect 1494 411 1500 412
rect 1494 410 1495 411
rect 1444 408 1495 410
rect 1444 407 1445 408
rect 1439 406 1445 407
rect 1494 407 1495 408
rect 1499 407 1500 411
rect 1494 406 1500 407
rect 1510 411 1516 412
rect 1510 407 1511 411
rect 1515 410 1516 411
rect 1527 411 1533 412
rect 1527 410 1528 411
rect 1515 408 1528 410
rect 1515 407 1516 408
rect 1510 406 1516 407
rect 1527 407 1528 408
rect 1532 407 1533 411
rect 1527 406 1533 407
rect 1615 411 1621 412
rect 1615 407 1616 411
rect 1620 410 1621 411
rect 1662 411 1668 412
rect 1662 410 1663 411
rect 1620 408 1663 410
rect 1620 407 1621 408
rect 1615 406 1621 407
rect 1662 407 1663 408
rect 1667 407 1668 411
rect 1662 406 1668 407
rect 1695 411 1701 412
rect 1695 407 1696 411
rect 1700 410 1701 411
rect 1742 411 1748 412
rect 1742 410 1743 411
rect 1700 408 1743 410
rect 1700 407 1701 408
rect 1695 406 1701 407
rect 1742 407 1743 408
rect 1747 407 1748 411
rect 1742 406 1748 407
rect 1775 411 1781 412
rect 1775 407 1776 411
rect 1780 410 1781 411
rect 1814 411 1820 412
rect 1814 410 1815 411
rect 1780 408 1815 410
rect 1780 407 1781 408
rect 1775 406 1781 407
rect 1814 407 1815 408
rect 1819 407 1820 411
rect 1814 406 1820 407
rect 1846 411 1853 412
rect 1846 407 1847 411
rect 1852 407 1853 411
rect 1846 406 1853 407
rect 1855 411 1861 412
rect 1855 407 1856 411
rect 1860 410 1861 411
rect 1911 411 1917 412
rect 1911 410 1912 411
rect 1860 408 1912 410
rect 1860 407 1861 408
rect 1855 406 1861 407
rect 1911 407 1912 408
rect 1916 407 1917 411
rect 1911 406 1917 407
rect 1922 411 1928 412
rect 1922 407 1923 411
rect 1927 410 1928 411
rect 1975 411 1981 412
rect 1975 410 1976 411
rect 1927 408 1976 410
rect 1927 407 1928 408
rect 1922 406 1928 407
rect 1975 407 1976 408
rect 1980 407 1981 411
rect 1975 406 1981 407
rect 2047 411 2053 412
rect 2047 407 2048 411
rect 2052 410 2053 411
rect 2062 411 2068 412
rect 2062 410 2063 411
rect 2052 408 2063 410
rect 2052 407 2053 408
rect 2047 406 2053 407
rect 2062 407 2063 408
rect 2067 407 2068 411
rect 2062 406 2068 407
rect 2082 411 2088 412
rect 2082 407 2083 411
rect 2087 410 2088 411
rect 2095 411 2101 412
rect 2095 410 2096 411
rect 2087 408 2096 410
rect 2087 407 2088 408
rect 2082 406 2088 407
rect 2095 407 2096 408
rect 2100 407 2101 411
rect 2095 406 2101 407
rect 2118 408 2124 409
rect 1134 403 1140 404
rect 2118 404 2119 408
rect 2123 404 2124 408
rect 2118 403 2124 404
rect 1094 399 1100 400
rect 1158 400 1164 401
rect 150 396 156 397
rect 150 392 151 396
rect 155 392 156 396
rect 150 391 156 392
rect 214 396 220 397
rect 214 392 215 396
rect 219 392 220 396
rect 214 391 220 392
rect 278 396 284 397
rect 278 392 279 396
rect 283 392 284 396
rect 278 391 284 392
rect 350 396 356 397
rect 350 392 351 396
rect 355 392 356 396
rect 350 391 356 392
rect 422 396 428 397
rect 422 392 423 396
rect 427 392 428 396
rect 422 391 428 392
rect 486 396 492 397
rect 486 392 487 396
rect 491 392 492 396
rect 486 391 492 392
rect 550 396 556 397
rect 550 392 551 396
rect 555 392 556 396
rect 550 391 556 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 726 396 732 397
rect 726 392 727 396
rect 731 392 732 396
rect 726 391 732 392
rect 790 396 796 397
rect 790 392 791 396
rect 795 392 796 396
rect 790 391 796 392
rect 854 396 860 397
rect 854 392 855 396
rect 859 392 860 396
rect 1158 396 1159 400
rect 1163 396 1164 400
rect 1158 395 1164 396
rect 1198 400 1204 401
rect 1198 396 1199 400
rect 1203 396 1204 400
rect 1198 395 1204 396
rect 1254 400 1260 401
rect 1254 396 1255 400
rect 1259 396 1260 400
rect 1254 395 1260 396
rect 1334 400 1340 401
rect 1334 396 1335 400
rect 1339 396 1340 400
rect 1334 395 1340 396
rect 1414 400 1420 401
rect 1414 396 1415 400
rect 1419 396 1420 400
rect 1414 395 1420 396
rect 1502 400 1508 401
rect 1502 396 1503 400
rect 1507 396 1508 400
rect 1502 395 1508 396
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1670 400 1676 401
rect 1670 396 1671 400
rect 1675 396 1676 400
rect 1670 395 1676 396
rect 1750 400 1756 401
rect 1750 396 1751 400
rect 1755 396 1756 400
rect 1750 395 1756 396
rect 1822 400 1828 401
rect 1822 396 1823 400
rect 1827 396 1828 400
rect 1822 395 1828 396
rect 1886 400 1892 401
rect 1886 396 1887 400
rect 1891 396 1892 400
rect 1886 395 1892 396
rect 1950 400 1956 401
rect 1950 396 1951 400
rect 1955 396 1956 400
rect 1950 395 1956 396
rect 2022 400 2028 401
rect 2022 396 2023 400
rect 2027 396 2028 400
rect 2022 395 2028 396
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 854 391 860 392
rect 1155 387 1161 388
rect 147 383 153 384
rect 147 379 148 383
rect 152 382 153 383
rect 158 383 164 384
rect 158 382 159 383
rect 152 380 159 382
rect 152 379 153 380
rect 147 378 153 379
rect 158 379 159 380
rect 163 379 164 383
rect 158 378 164 379
rect 211 383 217 384
rect 211 379 212 383
rect 216 382 217 383
rect 255 383 261 384
rect 255 382 256 383
rect 216 380 256 382
rect 216 379 217 380
rect 211 378 217 379
rect 255 379 256 380
rect 260 379 261 383
rect 255 378 261 379
rect 263 383 269 384
rect 263 379 264 383
rect 268 382 269 383
rect 275 383 281 384
rect 275 382 276 383
rect 268 380 276 382
rect 268 379 269 380
rect 263 378 269 379
rect 275 379 276 380
rect 280 379 281 383
rect 275 378 281 379
rect 347 383 353 384
rect 347 379 348 383
rect 352 382 353 383
rect 399 383 405 384
rect 399 382 400 383
rect 352 380 400 382
rect 352 379 353 380
rect 347 378 353 379
rect 399 379 400 380
rect 404 379 405 383
rect 399 378 405 379
rect 419 383 425 384
rect 419 379 420 383
rect 424 382 425 383
rect 455 383 461 384
rect 455 382 456 383
rect 424 380 456 382
rect 424 379 425 380
rect 419 378 425 379
rect 455 379 456 380
rect 460 379 461 383
rect 455 378 461 379
rect 483 383 489 384
rect 483 379 484 383
rect 488 382 489 383
rect 494 383 500 384
rect 494 382 495 383
rect 488 380 495 382
rect 488 379 489 380
rect 483 378 489 379
rect 494 379 495 380
rect 499 379 500 383
rect 494 378 500 379
rect 542 383 553 384
rect 542 379 543 383
rect 547 379 548 383
rect 552 379 553 383
rect 542 378 553 379
rect 602 383 608 384
rect 602 379 603 383
rect 607 382 608 383
rect 611 383 617 384
rect 611 382 612 383
rect 607 380 612 382
rect 607 379 608 380
rect 602 378 608 379
rect 611 379 612 380
rect 616 379 617 383
rect 611 378 617 379
rect 662 383 673 384
rect 662 379 663 383
rect 667 379 668 383
rect 672 379 673 383
rect 662 378 673 379
rect 718 383 729 384
rect 718 379 719 383
rect 723 379 724 383
rect 728 379 729 383
rect 718 378 729 379
rect 782 383 793 384
rect 782 379 783 383
rect 787 379 788 383
rect 792 379 793 383
rect 782 378 793 379
rect 846 383 857 384
rect 846 379 847 383
rect 851 379 852 383
rect 856 379 857 383
rect 1155 383 1156 387
rect 1160 386 1161 387
rect 1166 387 1172 388
rect 1166 386 1167 387
rect 1160 384 1167 386
rect 1160 383 1161 384
rect 1155 382 1161 383
rect 1166 383 1167 384
rect 1171 383 1172 387
rect 1166 382 1172 383
rect 1186 387 1192 388
rect 1186 383 1187 387
rect 1191 386 1192 387
rect 1195 387 1201 388
rect 1195 386 1196 387
rect 1191 384 1196 386
rect 1191 383 1192 384
rect 1186 382 1192 383
rect 1195 383 1196 384
rect 1200 383 1201 387
rect 1195 382 1201 383
rect 1246 387 1257 388
rect 1246 383 1247 387
rect 1251 383 1252 387
rect 1256 383 1257 387
rect 1246 382 1257 383
rect 1326 387 1337 388
rect 1326 383 1327 387
rect 1331 383 1332 387
rect 1336 383 1337 387
rect 1326 382 1337 383
rect 1406 387 1417 388
rect 1406 383 1407 387
rect 1411 383 1412 387
rect 1416 383 1417 387
rect 1406 382 1417 383
rect 1494 387 1505 388
rect 1494 383 1495 387
rect 1499 383 1500 387
rect 1504 383 1505 387
rect 1494 382 1505 383
rect 1582 387 1593 388
rect 1582 383 1583 387
rect 1587 383 1588 387
rect 1592 383 1593 387
rect 1582 382 1593 383
rect 1662 387 1673 388
rect 1662 383 1663 387
rect 1667 383 1668 387
rect 1672 383 1673 387
rect 1662 382 1673 383
rect 1742 387 1753 388
rect 1742 383 1743 387
rect 1747 383 1748 387
rect 1752 383 1753 387
rect 1742 382 1753 383
rect 1819 387 1825 388
rect 1819 383 1820 387
rect 1824 386 1825 387
rect 1855 387 1861 388
rect 1855 386 1856 387
rect 1824 384 1856 386
rect 1824 383 1825 384
rect 1819 382 1825 383
rect 1855 383 1856 384
rect 1860 383 1861 387
rect 1855 382 1861 383
rect 1883 387 1889 388
rect 1883 383 1884 387
rect 1888 386 1889 387
rect 1922 387 1928 388
rect 1922 386 1923 387
rect 1888 384 1923 386
rect 1888 383 1889 384
rect 1883 382 1889 383
rect 1922 383 1923 384
rect 1927 383 1928 387
rect 1922 382 1928 383
rect 1947 387 1953 388
rect 1947 383 1948 387
rect 1952 386 1953 387
rect 1998 387 2004 388
rect 1998 386 1999 387
rect 1952 384 1999 386
rect 1952 383 1953 384
rect 1947 382 1953 383
rect 1998 383 1999 384
rect 2003 383 2004 387
rect 1998 382 2004 383
rect 2019 387 2025 388
rect 2019 383 2020 387
rect 2024 386 2025 387
rect 2030 387 2036 388
rect 2030 386 2031 387
rect 2024 384 2031 386
rect 2024 383 2025 384
rect 2019 382 2025 383
rect 2030 383 2031 384
rect 2035 383 2036 387
rect 2030 382 2036 383
rect 2062 387 2073 388
rect 2062 383 2063 387
rect 2067 383 2068 387
rect 2072 383 2073 387
rect 2062 382 2073 383
rect 846 378 857 379
rect 1510 379 1516 380
rect 1510 378 1511 379
rect 1300 376 1511 378
rect 1300 374 1302 376
rect 1510 375 1511 376
rect 1515 375 1516 379
rect 1510 374 1516 375
rect 1299 373 1305 374
rect 131 371 137 372
rect 131 367 132 371
rect 136 370 137 371
rect 171 371 177 372
rect 136 368 166 370
rect 136 367 137 368
rect 131 366 137 367
rect 134 360 140 361
rect 134 356 135 360
rect 139 356 140 360
rect 134 355 140 356
rect 164 354 166 368
rect 171 367 172 371
rect 176 370 177 371
rect 206 371 217 372
rect 176 368 202 370
rect 176 367 177 368
rect 171 366 177 367
rect 174 360 180 361
rect 174 356 175 360
rect 179 356 180 360
rect 174 355 180 356
rect 200 354 202 368
rect 206 367 207 371
rect 211 367 212 371
rect 216 367 217 371
rect 206 366 217 367
rect 242 371 248 372
rect 242 367 243 371
rect 247 370 248 371
rect 267 371 273 372
rect 267 370 268 371
rect 247 368 268 370
rect 247 367 248 368
rect 242 366 248 367
rect 267 367 268 368
rect 272 367 273 371
rect 267 366 273 367
rect 298 371 304 372
rect 298 367 299 371
rect 303 370 304 371
rect 331 371 337 372
rect 331 370 332 371
rect 303 368 332 370
rect 303 367 304 368
rect 298 366 304 367
rect 331 367 332 368
rect 336 367 337 371
rect 331 366 337 367
rect 390 371 401 372
rect 390 367 391 371
rect 395 367 396 371
rect 400 367 401 371
rect 390 366 401 367
rect 410 371 416 372
rect 410 367 411 371
rect 415 370 416 371
rect 459 371 465 372
rect 459 370 460 371
rect 415 368 460 370
rect 415 367 416 368
rect 410 366 416 367
rect 459 367 460 368
rect 464 367 465 371
rect 459 366 465 367
rect 498 371 504 372
rect 498 367 499 371
rect 503 370 504 371
rect 515 371 521 372
rect 515 370 516 371
rect 503 368 516 370
rect 503 367 504 368
rect 498 366 504 367
rect 515 367 516 368
rect 520 367 521 371
rect 515 366 521 367
rect 571 371 577 372
rect 571 367 572 371
rect 576 370 577 371
rect 615 371 621 372
rect 615 370 616 371
rect 576 368 616 370
rect 576 367 577 368
rect 571 366 577 367
rect 615 367 616 368
rect 620 367 621 371
rect 615 366 621 367
rect 627 371 633 372
rect 627 367 628 371
rect 632 370 633 371
rect 646 371 652 372
rect 646 370 647 371
rect 632 368 647 370
rect 632 367 633 368
rect 627 366 633 367
rect 646 367 647 368
rect 651 367 652 371
rect 646 366 652 367
rect 658 371 664 372
rect 658 367 659 371
rect 663 370 664 371
rect 683 371 689 372
rect 683 370 684 371
rect 663 368 684 370
rect 663 367 664 368
rect 658 366 664 367
rect 683 367 684 368
rect 688 367 689 371
rect 683 366 689 367
rect 714 371 720 372
rect 714 367 715 371
rect 719 370 720 371
rect 747 371 753 372
rect 747 370 748 371
rect 719 368 748 370
rect 719 367 720 368
rect 714 366 720 367
rect 747 367 748 368
rect 752 367 753 371
rect 1299 369 1300 373
rect 1304 369 1305 373
rect 1299 368 1305 369
rect 1326 371 1332 372
rect 747 366 753 367
rect 1326 367 1327 371
rect 1331 370 1332 371
rect 1339 371 1345 372
rect 1339 370 1340 371
rect 1331 368 1340 370
rect 1331 367 1332 368
rect 1326 366 1332 367
rect 1339 367 1340 368
rect 1344 367 1345 371
rect 1339 366 1345 367
rect 1370 371 1376 372
rect 1370 367 1371 371
rect 1375 370 1376 371
rect 1379 371 1385 372
rect 1379 370 1380 371
rect 1375 368 1380 370
rect 1375 367 1376 368
rect 1370 366 1376 367
rect 1379 367 1380 368
rect 1384 367 1385 371
rect 1379 366 1385 367
rect 1406 371 1412 372
rect 1406 367 1407 371
rect 1411 370 1412 371
rect 1419 371 1425 372
rect 1419 370 1420 371
rect 1411 368 1420 370
rect 1411 367 1412 368
rect 1406 366 1412 367
rect 1419 367 1420 368
rect 1424 367 1425 371
rect 1419 366 1425 367
rect 1450 371 1456 372
rect 1450 367 1451 371
rect 1455 370 1456 371
rect 1459 371 1465 372
rect 1459 370 1460 371
rect 1455 368 1460 370
rect 1455 367 1456 368
rect 1450 366 1456 367
rect 1459 367 1460 368
rect 1464 367 1465 371
rect 1459 366 1465 367
rect 1490 371 1496 372
rect 1490 367 1491 371
rect 1495 370 1496 371
rect 1499 371 1505 372
rect 1499 370 1500 371
rect 1495 368 1500 370
rect 1495 367 1496 368
rect 1490 366 1496 367
rect 1499 367 1500 368
rect 1504 367 1505 371
rect 1499 366 1505 367
rect 1547 371 1553 372
rect 1547 367 1548 371
rect 1552 370 1553 371
rect 1570 371 1576 372
rect 1570 370 1571 371
rect 1552 368 1571 370
rect 1552 367 1553 368
rect 1547 366 1553 367
rect 1570 367 1571 368
rect 1575 367 1576 371
rect 1570 366 1576 367
rect 1578 371 1584 372
rect 1578 367 1579 371
rect 1583 370 1584 371
rect 1611 371 1617 372
rect 1611 370 1612 371
rect 1583 368 1612 370
rect 1583 367 1584 368
rect 1578 366 1584 367
rect 1611 367 1612 368
rect 1616 367 1617 371
rect 1611 366 1617 367
rect 1642 371 1648 372
rect 1642 367 1643 371
rect 1647 370 1648 371
rect 1675 371 1681 372
rect 1675 370 1676 371
rect 1647 368 1676 370
rect 1647 367 1648 368
rect 1642 366 1648 367
rect 1675 367 1676 368
rect 1680 367 1681 371
rect 1675 366 1681 367
rect 1706 371 1712 372
rect 1706 367 1707 371
rect 1711 370 1712 371
rect 1747 371 1753 372
rect 1747 370 1748 371
rect 1711 368 1748 370
rect 1711 367 1712 368
rect 1706 366 1712 367
rect 1747 367 1748 368
rect 1752 367 1753 371
rect 1747 366 1753 367
rect 1814 371 1820 372
rect 1814 367 1815 371
rect 1819 370 1820 371
rect 1827 371 1833 372
rect 1827 370 1828 371
rect 1819 368 1828 370
rect 1819 367 1820 368
rect 1814 366 1820 367
rect 1827 367 1828 368
rect 1832 367 1833 371
rect 1827 366 1833 367
rect 1915 371 1921 372
rect 1915 367 1916 371
rect 1920 370 1921 371
rect 1942 371 1948 372
rect 1942 370 1943 371
rect 1920 368 1943 370
rect 1920 367 1921 368
rect 1915 366 1921 367
rect 1942 367 1943 368
rect 1947 367 1948 371
rect 1942 366 1948 367
rect 1951 371 1957 372
rect 1951 367 1952 371
rect 1956 370 1957 371
rect 2003 371 2009 372
rect 2003 370 2004 371
rect 1956 368 2004 370
rect 1956 367 1957 368
rect 1951 366 1957 367
rect 2003 367 2004 368
rect 2008 367 2009 371
rect 2003 366 2009 367
rect 2067 371 2073 372
rect 2067 367 2068 371
rect 2072 370 2073 371
rect 2082 371 2088 372
rect 2082 370 2083 371
rect 2072 368 2083 370
rect 2072 367 2073 368
rect 2067 366 2073 367
rect 2082 367 2083 368
rect 2087 367 2088 371
rect 2082 366 2088 367
rect 214 360 220 361
rect 214 356 215 360
rect 219 356 220 360
rect 214 355 220 356
rect 270 360 276 361
rect 270 356 271 360
rect 275 356 276 360
rect 270 355 276 356
rect 334 360 340 361
rect 334 356 335 360
rect 339 356 340 360
rect 334 355 340 356
rect 398 360 404 361
rect 398 356 399 360
rect 403 356 404 360
rect 398 355 404 356
rect 462 360 468 361
rect 462 356 463 360
rect 467 356 468 360
rect 462 355 468 356
rect 518 360 524 361
rect 518 356 519 360
rect 523 356 524 360
rect 518 355 524 356
rect 574 360 580 361
rect 574 356 575 360
rect 579 356 580 360
rect 574 355 580 356
rect 630 360 636 361
rect 630 356 631 360
rect 635 356 636 360
rect 630 355 636 356
rect 686 360 692 361
rect 686 356 687 360
rect 691 356 692 360
rect 686 355 692 356
rect 750 360 756 361
rect 750 356 751 360
rect 755 356 756 360
rect 750 355 756 356
rect 1302 360 1308 361
rect 1302 356 1303 360
rect 1307 356 1308 360
rect 1302 355 1308 356
rect 1342 360 1348 361
rect 1342 356 1343 360
rect 1347 356 1348 360
rect 1342 355 1348 356
rect 1382 360 1388 361
rect 1382 356 1383 360
rect 1387 356 1388 360
rect 1382 355 1388 356
rect 1422 360 1428 361
rect 1422 356 1423 360
rect 1427 356 1428 360
rect 1422 355 1428 356
rect 1462 360 1468 361
rect 1462 356 1463 360
rect 1467 356 1468 360
rect 1462 355 1468 356
rect 1502 360 1508 361
rect 1502 356 1503 360
rect 1507 356 1508 360
rect 1502 355 1508 356
rect 1550 360 1556 361
rect 1550 356 1551 360
rect 1555 356 1556 360
rect 1550 355 1556 356
rect 1614 360 1620 361
rect 1614 356 1615 360
rect 1619 356 1620 360
rect 1614 355 1620 356
rect 1678 360 1684 361
rect 1678 356 1679 360
rect 1683 356 1684 360
rect 1678 355 1684 356
rect 1750 360 1756 361
rect 1750 356 1751 360
rect 1755 356 1756 360
rect 1750 355 1756 356
rect 1830 360 1836 361
rect 1830 356 1831 360
rect 1835 356 1836 360
rect 1830 355 1836 356
rect 1918 360 1924 361
rect 1918 356 1919 360
rect 1923 356 1924 360
rect 1918 355 1924 356
rect 2006 360 2012 361
rect 2006 356 2007 360
rect 2011 356 2012 360
rect 2006 355 2012 356
rect 2070 360 2076 361
rect 2070 356 2071 360
rect 2075 356 2076 360
rect 2070 355 2076 356
rect 110 352 116 353
rect 164 352 170 354
rect 200 352 210 354
rect 110 348 111 352
rect 115 348 116 352
rect 110 347 116 348
rect 142 347 148 348
rect 142 343 143 347
rect 147 346 148 347
rect 159 347 165 348
rect 159 346 160 347
rect 147 344 160 346
rect 147 343 148 344
rect 142 342 148 343
rect 159 343 160 344
rect 164 343 165 347
rect 168 346 170 352
rect 208 350 210 352
rect 233 352 266 354
rect 233 350 235 352
rect 208 348 235 350
rect 264 350 266 352
rect 288 352 321 354
rect 649 352 682 354
rect 288 350 290 352
rect 264 348 290 350
rect 199 347 205 348
rect 199 346 200 347
rect 168 344 200 346
rect 159 342 165 343
rect 199 343 200 344
rect 204 343 205 347
rect 199 342 205 343
rect 239 347 248 348
rect 239 343 240 347
rect 247 343 248 347
rect 239 342 248 343
rect 295 347 304 348
rect 295 343 296 347
rect 303 343 304 347
rect 319 346 321 352
rect 615 351 621 352
rect 359 347 365 348
rect 359 346 360 347
rect 319 344 360 346
rect 295 342 304 343
rect 359 343 360 344
rect 364 343 365 347
rect 359 342 365 343
rect 370 347 376 348
rect 370 343 371 347
rect 375 346 376 347
rect 423 347 429 348
rect 423 346 424 347
rect 375 344 424 346
rect 375 343 376 344
rect 370 342 376 343
rect 423 343 424 344
rect 428 343 429 347
rect 423 342 429 343
rect 487 347 493 348
rect 487 343 488 347
rect 492 346 493 347
rect 498 347 504 348
rect 498 346 499 347
rect 492 344 499 346
rect 492 343 493 344
rect 487 342 493 343
rect 498 343 499 344
rect 503 343 504 347
rect 498 342 504 343
rect 542 347 549 348
rect 542 343 543 347
rect 548 343 549 347
rect 542 342 549 343
rect 599 347 608 348
rect 599 343 600 347
rect 607 343 608 347
rect 615 347 616 351
rect 620 350 621 351
rect 649 350 651 352
rect 620 348 651 350
rect 680 350 682 352
rect 704 352 726 354
rect 704 350 706 352
rect 680 348 706 350
rect 620 347 621 348
rect 615 346 621 347
rect 655 347 664 348
rect 599 342 608 343
rect 655 343 656 347
rect 663 343 664 347
rect 655 342 664 343
rect 711 347 720 348
rect 711 343 712 347
rect 719 343 720 347
rect 724 346 726 352
rect 1094 352 1100 353
rect 1094 348 1095 352
rect 1099 348 1100 352
rect 775 347 781 348
rect 1094 347 1100 348
rect 1134 352 1140 353
rect 1134 348 1135 352
rect 1139 348 1140 352
rect 2118 352 2124 353
rect 2118 348 2119 352
rect 2123 348 2124 352
rect 1134 347 1140 348
rect 1326 347 1333 348
rect 775 346 776 347
rect 724 344 776 346
rect 711 342 720 343
rect 775 343 776 344
rect 780 343 781 347
rect 775 342 781 343
rect 1326 343 1327 347
rect 1332 343 1333 347
rect 1326 342 1333 343
rect 1367 347 1376 348
rect 1367 343 1368 347
rect 1375 343 1376 347
rect 1367 342 1376 343
rect 1406 347 1413 348
rect 1406 343 1407 347
rect 1412 343 1413 347
rect 1406 342 1413 343
rect 1447 347 1456 348
rect 1447 343 1448 347
rect 1455 343 1456 347
rect 1447 342 1456 343
rect 1487 347 1496 348
rect 1487 343 1488 347
rect 1495 343 1496 347
rect 1487 342 1496 343
rect 1527 347 1533 348
rect 1527 343 1528 347
rect 1532 346 1533 347
rect 1542 347 1548 348
rect 1542 346 1543 347
rect 1532 344 1543 346
rect 1532 343 1533 344
rect 1527 342 1533 343
rect 1542 343 1543 344
rect 1547 343 1548 347
rect 1542 342 1548 343
rect 1575 347 1584 348
rect 1575 343 1576 347
rect 1583 343 1584 347
rect 1575 342 1584 343
rect 1639 347 1648 348
rect 1639 343 1640 347
rect 1647 343 1648 347
rect 1639 342 1648 343
rect 1703 347 1712 348
rect 1703 343 1704 347
rect 1711 343 1712 347
rect 1703 342 1712 343
rect 1714 347 1720 348
rect 1714 343 1715 347
rect 1719 346 1720 347
rect 1775 347 1781 348
rect 1775 346 1776 347
rect 1719 344 1776 346
rect 1719 343 1720 344
rect 1714 342 1720 343
rect 1775 343 1776 344
rect 1780 343 1781 347
rect 1775 342 1781 343
rect 1786 347 1792 348
rect 1786 343 1787 347
rect 1791 346 1792 347
rect 1855 347 1861 348
rect 1855 346 1856 347
rect 1791 344 1856 346
rect 1791 343 1792 344
rect 1786 342 1792 343
rect 1855 343 1856 344
rect 1860 343 1861 347
rect 1855 342 1861 343
rect 1943 347 1949 348
rect 1943 343 1944 347
rect 1948 346 1949 347
rect 1951 347 1957 348
rect 1951 346 1952 347
rect 1948 344 1952 346
rect 1948 343 1949 344
rect 1943 342 1949 343
rect 1951 343 1952 344
rect 1956 343 1957 347
rect 1951 342 1957 343
rect 1998 347 2004 348
rect 1998 343 1999 347
rect 2003 346 2004 347
rect 2031 347 2037 348
rect 2031 346 2032 347
rect 2003 344 2032 346
rect 2003 343 2004 344
rect 1998 342 2004 343
rect 2031 343 2032 344
rect 2036 343 2037 347
rect 2031 342 2037 343
rect 2078 347 2084 348
rect 2078 343 2079 347
rect 2083 346 2084 347
rect 2095 347 2101 348
rect 2118 347 2124 348
rect 2095 346 2096 347
rect 2083 344 2096 346
rect 2083 343 2084 344
rect 2078 342 2084 343
rect 2095 343 2096 344
rect 2100 343 2101 347
rect 2095 342 2101 343
rect 110 335 116 336
rect 110 331 111 335
rect 115 331 116 335
rect 1094 335 1100 336
rect 110 330 116 331
rect 134 332 140 333
rect 134 328 135 332
rect 139 328 140 332
rect 134 327 140 328
rect 174 332 180 333
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 214 332 220 333
rect 214 328 215 332
rect 219 328 220 332
rect 214 327 220 328
rect 270 332 276 333
rect 270 328 271 332
rect 275 328 276 332
rect 270 327 276 328
rect 334 332 340 333
rect 334 328 335 332
rect 339 328 340 332
rect 334 327 340 328
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 462 332 468 333
rect 462 328 463 332
rect 467 328 468 332
rect 462 327 468 328
rect 518 332 524 333
rect 518 328 519 332
rect 523 328 524 332
rect 518 327 524 328
rect 574 332 580 333
rect 574 328 575 332
rect 579 328 580 332
rect 574 327 580 328
rect 630 332 636 333
rect 630 328 631 332
rect 635 328 636 332
rect 630 327 636 328
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 750 332 756 333
rect 750 328 751 332
rect 755 328 756 332
rect 1094 331 1095 335
rect 1099 331 1100 335
rect 1094 330 1100 331
rect 1134 335 1140 336
rect 1134 331 1135 335
rect 1139 331 1140 335
rect 2118 335 2124 336
rect 1134 330 1140 331
rect 1302 332 1308 333
rect 750 327 756 328
rect 1302 328 1303 332
rect 1307 328 1308 332
rect 1302 327 1308 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1342 327 1348 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1422 332 1428 333
rect 1422 328 1423 332
rect 1427 328 1428 332
rect 1422 327 1428 328
rect 1462 332 1468 333
rect 1462 328 1463 332
rect 1467 328 1468 332
rect 1462 327 1468 328
rect 1502 332 1508 333
rect 1502 328 1503 332
rect 1507 328 1508 332
rect 1502 327 1508 328
rect 1550 332 1556 333
rect 1550 328 1551 332
rect 1555 328 1556 332
rect 1550 327 1556 328
rect 1614 332 1620 333
rect 1614 328 1615 332
rect 1619 328 1620 332
rect 1614 327 1620 328
rect 1678 332 1684 333
rect 1678 328 1679 332
rect 1683 328 1684 332
rect 1678 327 1684 328
rect 1750 332 1756 333
rect 1750 328 1751 332
rect 1755 328 1756 332
rect 1750 327 1756 328
rect 1830 332 1836 333
rect 1830 328 1831 332
rect 1835 328 1836 332
rect 1830 327 1836 328
rect 1918 332 1924 333
rect 1918 328 1919 332
rect 1923 328 1924 332
rect 1918 327 1924 328
rect 2006 332 2012 333
rect 2006 328 2007 332
rect 2011 328 2012 332
rect 2006 327 2012 328
rect 2070 332 2076 333
rect 2070 328 2071 332
rect 2075 328 2076 332
rect 2118 331 2119 335
rect 2123 331 2124 335
rect 2118 330 2124 331
rect 2070 327 2076 328
rect 255 323 261 324
rect 255 319 256 323
rect 260 322 261 323
rect 370 323 376 324
rect 370 322 371 323
rect 260 320 371 322
rect 260 319 261 320
rect 255 318 261 319
rect 370 319 371 320
rect 375 319 376 323
rect 370 318 376 319
rect 134 316 140 317
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 134 312 135 316
rect 139 312 140 316
rect 134 311 140 312
rect 206 316 212 317
rect 206 312 207 316
rect 211 312 212 316
rect 206 311 212 312
rect 294 316 300 317
rect 294 312 295 316
rect 299 312 300 316
rect 294 311 300 312
rect 382 316 388 317
rect 382 312 383 316
rect 387 312 388 316
rect 382 311 388 312
rect 470 316 476 317
rect 470 312 471 316
rect 475 312 476 316
rect 470 311 476 312
rect 550 316 556 317
rect 550 312 551 316
rect 555 312 556 316
rect 550 311 556 312
rect 622 316 628 317
rect 622 312 623 316
rect 627 312 628 316
rect 622 311 628 312
rect 686 316 692 317
rect 686 312 687 316
rect 691 312 692 316
rect 686 311 692 312
rect 750 316 756 317
rect 750 312 751 316
rect 755 312 756 316
rect 750 311 756 312
rect 806 316 812 317
rect 806 312 807 316
rect 811 312 812 316
rect 806 311 812 312
rect 870 316 876 317
rect 870 312 871 316
rect 875 312 876 316
rect 870 311 876 312
rect 934 316 940 317
rect 934 312 935 316
rect 939 312 940 316
rect 1166 316 1172 317
rect 934 311 940 312
rect 1094 313 1100 314
rect 110 308 116 309
rect 1094 309 1095 313
rect 1099 309 1100 313
rect 1094 308 1100 309
rect 1134 313 1140 314
rect 1134 309 1135 313
rect 1139 309 1140 313
rect 1166 312 1167 316
rect 1171 312 1172 316
rect 1166 311 1172 312
rect 1206 316 1212 317
rect 1206 312 1207 316
rect 1211 312 1212 316
rect 1206 311 1212 312
rect 1246 316 1252 317
rect 1246 312 1247 316
rect 1251 312 1252 316
rect 1246 311 1252 312
rect 1294 316 1300 317
rect 1294 312 1295 316
rect 1299 312 1300 316
rect 1294 311 1300 312
rect 1342 316 1348 317
rect 1342 312 1343 316
rect 1347 312 1348 316
rect 1342 311 1348 312
rect 1390 316 1396 317
rect 1390 312 1391 316
rect 1395 312 1396 316
rect 1390 311 1396 312
rect 1438 316 1444 317
rect 1438 312 1439 316
rect 1443 312 1444 316
rect 1438 311 1444 312
rect 1494 316 1500 317
rect 1494 312 1495 316
rect 1499 312 1500 316
rect 1494 311 1500 312
rect 1558 316 1564 317
rect 1558 312 1559 316
rect 1563 312 1564 316
rect 1558 311 1564 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1694 316 1700 317
rect 1694 312 1695 316
rect 1699 312 1700 316
rect 1694 311 1700 312
rect 1774 316 1780 317
rect 1774 312 1775 316
rect 1779 312 1780 316
rect 1774 311 1780 312
rect 1854 316 1860 317
rect 1854 312 1855 316
rect 1859 312 1860 316
rect 1854 311 1860 312
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 1934 311 1940 312
rect 2014 316 2020 317
rect 2014 312 2015 316
rect 2019 312 2020 316
rect 2014 311 2020 312
rect 2070 316 2076 317
rect 2070 312 2071 316
rect 2075 312 2076 316
rect 2070 311 2076 312
rect 2118 313 2124 314
rect 1134 308 1140 309
rect 2118 309 2119 313
rect 2123 309 2124 313
rect 2118 308 2124 309
rect 1318 307 1324 308
rect 1318 303 1319 307
rect 1323 306 1324 307
rect 1462 307 1468 308
rect 1323 304 1394 306
rect 1323 303 1324 304
rect 1318 302 1324 303
rect 159 299 165 300
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 159 295 160 299
rect 164 298 165 299
rect 191 299 197 300
rect 191 298 192 299
rect 164 296 192 298
rect 164 295 165 296
rect 159 294 165 295
rect 191 295 192 296
rect 196 295 197 299
rect 191 294 197 295
rect 231 299 237 300
rect 231 295 232 299
rect 236 298 237 299
rect 286 299 292 300
rect 286 298 287 299
rect 236 296 287 298
rect 236 295 237 296
rect 231 294 237 295
rect 286 295 287 296
rect 291 295 292 299
rect 286 294 292 295
rect 302 299 308 300
rect 302 295 303 299
rect 307 298 308 299
rect 319 299 325 300
rect 319 298 320 299
rect 307 296 320 298
rect 307 295 308 296
rect 302 294 308 295
rect 319 295 320 296
rect 324 295 325 299
rect 319 294 325 295
rect 407 299 416 300
rect 407 295 408 299
rect 415 295 416 299
rect 407 294 416 295
rect 418 299 424 300
rect 418 295 419 299
rect 423 298 424 299
rect 495 299 501 300
rect 495 298 496 299
rect 423 296 496 298
rect 423 295 424 296
rect 418 294 424 295
rect 495 295 496 296
rect 500 295 501 299
rect 495 294 501 295
rect 503 299 509 300
rect 503 295 504 299
rect 508 298 509 299
rect 575 299 581 300
rect 575 298 576 299
rect 508 296 576 298
rect 508 295 509 296
rect 503 294 509 295
rect 575 295 576 296
rect 580 295 581 299
rect 575 294 581 295
rect 646 299 653 300
rect 646 295 647 299
rect 652 295 653 299
rect 646 294 653 295
rect 655 299 661 300
rect 655 295 656 299
rect 660 298 661 299
rect 711 299 717 300
rect 711 298 712 299
rect 660 296 712 298
rect 660 295 661 296
rect 655 294 661 295
rect 711 295 712 296
rect 716 295 717 299
rect 711 294 717 295
rect 722 299 728 300
rect 722 295 723 299
rect 727 298 728 299
rect 775 299 781 300
rect 775 298 776 299
rect 727 296 776 298
rect 727 295 728 296
rect 722 294 728 295
rect 775 295 776 296
rect 780 295 781 299
rect 775 294 781 295
rect 783 299 789 300
rect 783 295 784 299
rect 788 298 789 299
rect 831 299 837 300
rect 831 298 832 299
rect 788 296 832 298
rect 788 295 789 296
rect 783 294 789 295
rect 831 295 832 296
rect 836 295 837 299
rect 831 294 837 295
rect 839 299 845 300
rect 839 295 840 299
rect 844 298 845 299
rect 895 299 901 300
rect 895 298 896 299
rect 844 296 896 298
rect 844 295 845 296
rect 839 294 845 295
rect 895 295 896 296
rect 900 295 901 299
rect 959 299 965 300
rect 959 298 960 299
rect 895 294 901 295
rect 916 296 960 298
rect 110 291 116 292
rect 916 290 918 296
rect 959 295 960 296
rect 964 295 965 299
rect 1174 299 1180 300
rect 959 294 965 295
rect 1094 296 1100 297
rect 1094 292 1095 296
rect 1099 292 1100 296
rect 1094 291 1100 292
rect 1134 296 1140 297
rect 1134 292 1135 296
rect 1139 292 1140 296
rect 1174 295 1175 299
rect 1179 298 1180 299
rect 1191 299 1197 300
rect 1191 298 1192 299
rect 1179 296 1192 298
rect 1179 295 1180 296
rect 1174 294 1180 295
rect 1191 295 1192 296
rect 1196 295 1197 299
rect 1231 299 1237 300
rect 1231 298 1232 299
rect 1191 294 1197 295
rect 1200 296 1232 298
rect 1134 291 1140 292
rect 134 288 140 289
rect 134 284 135 288
rect 139 284 140 288
rect 134 283 140 284
rect 206 288 212 289
rect 206 284 207 288
rect 211 284 212 288
rect 206 283 212 284
rect 294 288 300 289
rect 294 284 295 288
rect 299 284 300 288
rect 294 283 300 284
rect 382 288 388 289
rect 382 284 383 288
rect 387 284 388 288
rect 382 283 388 284
rect 470 288 476 289
rect 470 284 471 288
rect 475 284 476 288
rect 470 283 476 284
rect 550 288 556 289
rect 550 284 551 288
rect 555 284 556 288
rect 550 283 556 284
rect 622 288 628 289
rect 622 284 623 288
rect 627 284 628 288
rect 622 283 628 284
rect 686 288 692 289
rect 686 284 687 288
rect 691 284 692 288
rect 686 283 692 284
rect 750 288 756 289
rect 750 284 751 288
rect 755 284 756 288
rect 750 283 756 284
rect 806 288 812 289
rect 806 284 807 288
rect 811 284 812 288
rect 806 283 812 284
rect 870 288 876 289
rect 870 284 871 288
rect 875 284 876 288
rect 870 283 876 284
rect 880 288 918 290
rect 934 288 940 289
rect 880 278 882 288
rect 934 284 935 288
rect 939 284 940 288
rect 934 283 940 284
rect 1166 288 1172 289
rect 1166 284 1167 288
rect 1171 284 1172 288
rect 1200 286 1202 296
rect 1231 295 1232 296
rect 1236 295 1237 299
rect 1271 299 1277 300
rect 1271 298 1272 299
rect 1231 294 1237 295
rect 1240 296 1272 298
rect 1166 283 1172 284
rect 1176 284 1202 286
rect 1206 288 1212 289
rect 1206 284 1207 288
rect 1211 284 1212 288
rect 1176 278 1178 284
rect 1206 283 1212 284
rect 1240 282 1242 296
rect 1271 295 1272 296
rect 1276 295 1277 299
rect 1271 294 1277 295
rect 1279 299 1285 300
rect 1279 295 1280 299
rect 1284 298 1285 299
rect 1319 299 1325 300
rect 1319 298 1320 299
rect 1284 296 1320 298
rect 1284 295 1285 296
rect 1279 294 1285 295
rect 1319 295 1320 296
rect 1324 295 1325 299
rect 1319 294 1325 295
rect 1367 299 1373 300
rect 1367 295 1368 299
rect 1372 298 1373 299
rect 1382 299 1388 300
rect 1382 298 1383 299
rect 1372 296 1383 298
rect 1372 295 1373 296
rect 1367 294 1373 295
rect 1382 295 1383 296
rect 1387 295 1388 299
rect 1392 298 1394 304
rect 1462 303 1463 307
rect 1467 306 1468 307
rect 1467 304 1594 306
rect 1467 303 1468 304
rect 1462 302 1468 303
rect 1415 299 1421 300
rect 1415 298 1416 299
rect 1392 296 1416 298
rect 1382 294 1388 295
rect 1415 295 1416 296
rect 1420 295 1421 299
rect 1415 294 1421 295
rect 1463 299 1469 300
rect 1463 295 1464 299
rect 1468 298 1469 299
rect 1486 299 1492 300
rect 1486 298 1487 299
rect 1468 296 1487 298
rect 1468 295 1469 296
rect 1463 294 1469 295
rect 1486 295 1487 296
rect 1491 295 1492 299
rect 1486 294 1492 295
rect 1518 299 1525 300
rect 1518 295 1519 299
rect 1524 295 1525 299
rect 1518 294 1525 295
rect 1570 299 1576 300
rect 1570 295 1571 299
rect 1575 298 1576 299
rect 1583 299 1589 300
rect 1583 298 1584 299
rect 1575 296 1584 298
rect 1575 295 1576 296
rect 1570 294 1576 295
rect 1583 295 1584 296
rect 1588 295 1589 299
rect 1592 298 1594 304
rect 1647 299 1653 300
rect 1647 298 1648 299
rect 1592 296 1648 298
rect 1583 294 1589 295
rect 1647 295 1648 296
rect 1652 295 1653 299
rect 1647 294 1653 295
rect 1655 299 1661 300
rect 1655 295 1656 299
rect 1660 298 1661 299
rect 1719 299 1725 300
rect 1719 298 1720 299
rect 1660 296 1720 298
rect 1660 295 1661 296
rect 1655 294 1661 295
rect 1719 295 1720 296
rect 1724 295 1725 299
rect 1719 294 1725 295
rect 1730 299 1736 300
rect 1730 295 1731 299
rect 1735 298 1736 299
rect 1799 299 1805 300
rect 1799 298 1800 299
rect 1735 296 1800 298
rect 1735 295 1736 296
rect 1730 294 1736 295
rect 1799 295 1800 296
rect 1804 295 1805 299
rect 1799 294 1805 295
rect 1879 299 1885 300
rect 1879 295 1880 299
rect 1884 298 1885 299
rect 1926 299 1932 300
rect 1926 298 1927 299
rect 1884 296 1927 298
rect 1884 295 1885 296
rect 1879 294 1885 295
rect 1926 295 1927 296
rect 1931 295 1932 299
rect 1926 294 1932 295
rect 1942 299 1948 300
rect 1942 295 1943 299
rect 1947 298 1948 299
rect 1959 299 1965 300
rect 1959 298 1960 299
rect 1947 296 1960 298
rect 1947 295 1948 296
rect 1942 294 1948 295
rect 1959 295 1960 296
rect 1964 295 1965 299
rect 1959 294 1965 295
rect 2006 299 2012 300
rect 2006 295 2007 299
rect 2011 298 2012 299
rect 2039 299 2045 300
rect 2039 298 2040 299
rect 2011 296 2040 298
rect 2011 295 2012 296
rect 2006 294 2012 295
rect 2039 295 2040 296
rect 2044 295 2045 299
rect 2039 294 2045 295
rect 2047 299 2053 300
rect 2047 295 2048 299
rect 2052 298 2053 299
rect 2095 299 2101 300
rect 2095 298 2096 299
rect 2052 296 2096 298
rect 2052 295 2053 296
rect 2047 294 2053 295
rect 2095 295 2096 296
rect 2100 295 2101 299
rect 2095 294 2101 295
rect 2118 296 2124 297
rect 2118 292 2119 296
rect 2123 292 2124 296
rect 2118 291 2124 292
rect 1246 288 1252 289
rect 1246 284 1247 288
rect 1251 284 1252 288
rect 1246 283 1252 284
rect 1294 288 1300 289
rect 1294 284 1295 288
rect 1299 284 1300 288
rect 1294 283 1300 284
rect 1342 288 1348 289
rect 1342 284 1343 288
rect 1347 284 1348 288
rect 1342 283 1348 284
rect 1390 288 1396 289
rect 1390 284 1391 288
rect 1395 284 1396 288
rect 1390 283 1396 284
rect 1438 288 1444 289
rect 1438 284 1439 288
rect 1443 284 1444 288
rect 1438 283 1444 284
rect 1494 288 1500 289
rect 1494 284 1495 288
rect 1499 284 1500 288
rect 1494 283 1500 284
rect 1558 288 1564 289
rect 1558 284 1559 288
rect 1563 284 1564 288
rect 1558 283 1564 284
rect 1622 288 1628 289
rect 1622 284 1623 288
rect 1627 284 1628 288
rect 1622 283 1628 284
rect 1694 288 1700 289
rect 1694 284 1695 288
rect 1699 284 1700 288
rect 1694 283 1700 284
rect 1774 288 1780 289
rect 1774 284 1775 288
rect 1779 284 1780 288
rect 1774 283 1780 284
rect 1854 288 1860 289
rect 1854 284 1855 288
rect 1859 284 1860 288
rect 1854 283 1860 284
rect 1934 288 1940 289
rect 1934 284 1935 288
rect 1939 284 1940 288
rect 1934 283 1940 284
rect 2014 288 2020 289
rect 2014 284 2015 288
rect 2019 284 2020 288
rect 2014 283 2020 284
rect 2070 288 2076 289
rect 2070 284 2071 288
rect 2075 284 2076 288
rect 2070 283 2076 284
rect 1228 280 1242 282
rect 1228 278 1230 280
rect 867 277 882 278
rect 131 275 137 276
rect 131 271 132 275
rect 136 274 137 275
rect 142 275 148 276
rect 142 274 143 275
rect 136 272 143 274
rect 136 271 137 272
rect 131 270 137 271
rect 142 271 143 272
rect 147 271 148 275
rect 142 270 148 271
rect 191 275 197 276
rect 191 271 192 275
rect 196 274 197 275
rect 203 275 209 276
rect 203 274 204 275
rect 196 272 204 274
rect 196 271 197 272
rect 191 270 197 271
rect 203 271 204 272
rect 208 271 209 275
rect 203 270 209 271
rect 286 275 297 276
rect 286 271 287 275
rect 291 271 292 275
rect 296 271 297 275
rect 286 270 297 271
rect 379 275 385 276
rect 379 271 380 275
rect 384 274 385 275
rect 418 275 424 276
rect 418 274 419 275
rect 384 272 419 274
rect 384 271 385 272
rect 379 270 385 271
rect 418 271 419 272
rect 423 271 424 275
rect 418 270 424 271
rect 467 275 473 276
rect 467 271 468 275
rect 472 274 473 275
rect 503 275 509 276
rect 503 274 504 275
rect 472 272 504 274
rect 472 271 473 272
rect 467 270 473 271
rect 503 271 504 272
rect 508 271 509 275
rect 503 270 509 271
rect 538 275 544 276
rect 538 271 539 275
rect 543 274 544 275
rect 547 275 553 276
rect 547 274 548 275
rect 543 272 548 274
rect 543 271 544 272
rect 538 270 544 271
rect 547 271 548 272
rect 552 271 553 275
rect 547 270 553 271
rect 619 275 625 276
rect 619 271 620 275
rect 624 274 625 275
rect 655 275 661 276
rect 655 274 656 275
rect 624 272 656 274
rect 624 271 625 272
rect 619 270 625 271
rect 655 271 656 272
rect 660 271 661 275
rect 655 270 661 271
rect 683 275 689 276
rect 683 271 684 275
rect 688 274 689 275
rect 722 275 728 276
rect 722 274 723 275
rect 688 272 723 274
rect 688 271 689 272
rect 683 270 689 271
rect 722 271 723 272
rect 727 271 728 275
rect 722 270 728 271
rect 747 275 753 276
rect 747 271 748 275
rect 752 274 753 275
rect 783 275 789 276
rect 783 274 784 275
rect 752 272 784 274
rect 752 271 753 272
rect 747 270 753 271
rect 783 271 784 272
rect 788 271 789 275
rect 783 270 789 271
rect 803 275 809 276
rect 803 271 804 275
rect 808 274 809 275
rect 839 275 845 276
rect 839 274 840 275
rect 808 272 840 274
rect 808 271 809 272
rect 803 270 809 271
rect 839 271 840 272
rect 844 271 845 275
rect 867 273 868 277
rect 872 276 882 277
rect 1163 277 1178 278
rect 872 273 873 276
rect 867 272 873 273
rect 906 275 912 276
rect 839 270 845 271
rect 906 271 907 275
rect 911 274 912 275
rect 931 275 937 276
rect 931 274 932 275
rect 911 272 932 274
rect 911 271 912 272
rect 906 270 912 271
rect 931 271 932 272
rect 936 271 937 275
rect 1163 273 1164 277
rect 1168 276 1178 277
rect 1203 277 1230 278
rect 1168 273 1169 276
rect 1163 272 1169 273
rect 1203 273 1204 277
rect 1208 276 1230 277
rect 1208 273 1209 276
rect 1203 272 1209 273
rect 1243 275 1249 276
rect 931 270 937 271
rect 1243 271 1244 275
rect 1248 274 1249 275
rect 1279 275 1285 276
rect 1279 274 1280 275
rect 1248 272 1280 274
rect 1248 271 1249 272
rect 1243 270 1249 271
rect 1279 271 1280 272
rect 1284 271 1285 275
rect 1279 270 1285 271
rect 1291 275 1297 276
rect 1291 271 1292 275
rect 1296 274 1297 275
rect 1318 275 1324 276
rect 1318 274 1319 275
rect 1296 272 1319 274
rect 1296 271 1297 272
rect 1291 270 1297 271
rect 1318 271 1319 272
rect 1323 271 1324 275
rect 1318 270 1324 271
rect 1339 275 1345 276
rect 1339 271 1340 275
rect 1344 274 1345 275
rect 1350 275 1356 276
rect 1350 274 1351 275
rect 1344 272 1351 274
rect 1344 271 1345 272
rect 1339 270 1345 271
rect 1350 271 1351 272
rect 1355 271 1356 275
rect 1350 270 1356 271
rect 1382 275 1393 276
rect 1382 271 1383 275
rect 1387 271 1388 275
rect 1392 271 1393 275
rect 1382 270 1393 271
rect 1435 275 1441 276
rect 1435 271 1436 275
rect 1440 274 1441 275
rect 1462 275 1468 276
rect 1462 274 1463 275
rect 1440 272 1463 274
rect 1440 271 1441 272
rect 1435 270 1441 271
rect 1462 271 1463 272
rect 1467 271 1468 275
rect 1462 270 1468 271
rect 1486 275 1497 276
rect 1486 271 1487 275
rect 1491 271 1492 275
rect 1496 271 1497 275
rect 1486 270 1497 271
rect 1542 275 1548 276
rect 1542 271 1543 275
rect 1547 274 1548 275
rect 1555 275 1561 276
rect 1555 274 1556 275
rect 1547 272 1556 274
rect 1547 271 1548 272
rect 1542 270 1548 271
rect 1555 271 1556 272
rect 1560 271 1561 275
rect 1555 270 1561 271
rect 1619 275 1625 276
rect 1619 271 1620 275
rect 1624 274 1625 275
rect 1691 275 1697 276
rect 1624 272 1670 274
rect 1624 271 1625 272
rect 1619 270 1625 271
rect 1668 266 1670 272
rect 1691 271 1692 275
rect 1696 274 1697 275
rect 1730 275 1736 276
rect 1730 274 1731 275
rect 1696 272 1731 274
rect 1696 271 1697 272
rect 1691 270 1697 271
rect 1730 271 1731 272
rect 1735 271 1736 275
rect 1730 270 1736 271
rect 1771 275 1777 276
rect 1771 271 1772 275
rect 1776 274 1777 275
rect 1786 275 1792 276
rect 1786 274 1787 275
rect 1776 272 1787 274
rect 1776 271 1777 272
rect 1771 270 1777 271
rect 1786 271 1787 272
rect 1791 271 1792 275
rect 1786 270 1792 271
rect 1851 275 1857 276
rect 1851 271 1852 275
rect 1856 274 1857 275
rect 1862 275 1868 276
rect 1862 274 1863 275
rect 1856 272 1863 274
rect 1856 271 1857 272
rect 1851 270 1857 271
rect 1862 271 1863 272
rect 1867 271 1868 275
rect 1862 270 1868 271
rect 1926 275 1937 276
rect 1926 271 1927 275
rect 1931 271 1932 275
rect 1936 271 1937 275
rect 1926 270 1937 271
rect 2011 275 2017 276
rect 2011 271 2012 275
rect 2016 274 2017 275
rect 2047 275 2053 276
rect 2047 274 2048 275
rect 2016 272 2048 274
rect 2016 271 2017 272
rect 2011 270 2017 271
rect 2047 271 2048 272
rect 2052 271 2053 275
rect 2047 270 2053 271
rect 2067 275 2073 276
rect 2067 271 2068 275
rect 2072 274 2073 275
rect 2078 275 2084 276
rect 2078 274 2079 275
rect 2072 272 2079 274
rect 2072 271 2073 272
rect 2067 270 2073 271
rect 2078 271 2079 272
rect 2083 271 2084 275
rect 2078 270 2084 271
rect 1714 267 1720 268
rect 1714 266 1715 267
rect 1668 264 1715 266
rect 131 263 137 264
rect 131 259 132 263
rect 136 262 137 263
rect 186 263 192 264
rect 186 262 187 263
rect 136 260 187 262
rect 136 259 137 260
rect 131 258 137 259
rect 186 259 187 260
rect 191 259 192 263
rect 186 258 192 259
rect 195 263 201 264
rect 195 259 196 263
rect 200 262 201 263
rect 266 263 272 264
rect 266 262 267 263
rect 200 260 267 262
rect 200 259 201 260
rect 195 258 201 259
rect 266 259 267 260
rect 271 259 272 263
rect 266 258 272 259
rect 275 263 281 264
rect 275 259 276 263
rect 280 262 281 263
rect 302 263 308 264
rect 302 262 303 263
rect 280 260 303 262
rect 280 259 281 260
rect 275 258 281 259
rect 302 259 303 260
rect 307 259 308 263
rect 302 258 308 259
rect 350 263 361 264
rect 350 259 351 263
rect 355 259 356 263
rect 360 259 361 263
rect 350 258 361 259
rect 390 263 396 264
rect 390 259 391 263
rect 395 262 396 263
rect 435 263 441 264
rect 435 262 436 263
rect 395 260 436 262
rect 395 259 396 260
rect 390 258 396 259
rect 435 259 436 260
rect 440 259 441 263
rect 435 258 441 259
rect 471 263 477 264
rect 471 259 472 263
rect 476 262 477 263
rect 507 263 513 264
rect 507 262 508 263
rect 476 260 508 262
rect 476 259 477 260
rect 471 258 477 259
rect 507 259 508 260
rect 512 259 513 263
rect 507 258 513 259
rect 579 263 585 264
rect 579 259 580 263
rect 584 262 585 263
rect 590 263 596 264
rect 590 262 591 263
rect 584 260 591 262
rect 584 259 585 260
rect 579 258 585 259
rect 590 259 591 260
rect 595 259 596 263
rect 590 258 596 259
rect 610 263 616 264
rect 610 259 611 263
rect 615 262 616 263
rect 643 263 649 264
rect 643 262 644 263
rect 615 260 644 262
rect 615 259 616 260
rect 610 258 616 259
rect 643 259 644 260
rect 648 259 649 263
rect 643 258 649 259
rect 679 263 685 264
rect 679 259 680 263
rect 684 262 685 263
rect 699 263 705 264
rect 699 262 700 263
rect 684 260 700 262
rect 684 259 685 260
rect 679 258 685 259
rect 699 259 700 260
rect 704 259 705 263
rect 699 258 705 259
rect 730 263 736 264
rect 730 259 731 263
rect 735 262 736 263
rect 755 263 761 264
rect 755 262 756 263
rect 735 260 756 262
rect 735 259 736 260
rect 730 258 736 259
rect 755 259 756 260
rect 760 259 761 263
rect 755 258 761 259
rect 786 263 792 264
rect 786 259 787 263
rect 791 262 792 263
rect 811 263 817 264
rect 811 262 812 263
rect 791 260 812 262
rect 791 259 792 260
rect 786 258 792 259
rect 811 259 812 260
rect 816 259 817 263
rect 811 258 817 259
rect 842 263 848 264
rect 842 259 843 263
rect 847 262 848 263
rect 875 263 881 264
rect 875 262 876 263
rect 847 260 876 262
rect 847 259 848 260
rect 842 258 848 259
rect 875 259 876 260
rect 880 259 881 263
rect 1655 263 1661 264
rect 1655 262 1656 263
rect 875 258 881 259
rect 1604 260 1656 262
rect 1604 258 1606 260
rect 1655 259 1656 260
rect 1660 259 1661 263
rect 1714 263 1715 264
rect 1719 263 1720 267
rect 1714 262 1720 263
rect 1655 258 1661 259
rect 1603 257 1609 258
rect 1155 255 1161 256
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 198 252 204 253
rect 198 248 199 252
rect 203 248 204 252
rect 198 247 204 248
rect 278 252 284 253
rect 278 248 279 252
rect 283 248 284 252
rect 278 247 284 248
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 438 252 444 253
rect 438 248 439 252
rect 443 248 444 252
rect 438 247 444 248
rect 510 252 516 253
rect 510 248 511 252
rect 515 248 516 252
rect 510 247 516 248
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 646 252 652 253
rect 646 248 647 252
rect 651 248 652 252
rect 646 247 652 248
rect 702 252 708 253
rect 702 248 703 252
rect 707 248 708 252
rect 702 247 708 248
rect 758 252 764 253
rect 758 248 759 252
rect 763 248 764 252
rect 758 247 764 248
rect 814 252 820 253
rect 814 248 815 252
rect 819 248 820 252
rect 814 247 820 248
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 1155 251 1156 255
rect 1160 254 1161 255
rect 1174 255 1180 256
rect 1174 254 1175 255
rect 1160 252 1175 254
rect 1160 251 1161 252
rect 1155 250 1161 251
rect 1174 251 1175 252
rect 1179 251 1180 255
rect 1174 250 1180 251
rect 1186 255 1192 256
rect 1186 251 1187 255
rect 1191 254 1192 255
rect 1203 255 1209 256
rect 1203 254 1204 255
rect 1191 252 1204 254
rect 1191 251 1192 252
rect 1186 250 1192 251
rect 1203 251 1204 252
rect 1208 251 1209 255
rect 1203 250 1209 251
rect 1234 255 1240 256
rect 1234 251 1235 255
rect 1239 254 1240 255
rect 1267 255 1273 256
rect 1267 254 1268 255
rect 1239 252 1268 254
rect 1239 251 1240 252
rect 1234 250 1240 251
rect 1267 251 1268 252
rect 1272 251 1273 255
rect 1267 250 1273 251
rect 1323 255 1329 256
rect 1323 251 1324 255
rect 1328 254 1329 255
rect 1378 255 1384 256
rect 1378 254 1379 255
rect 1328 252 1379 254
rect 1328 251 1329 252
rect 1323 250 1329 251
rect 1378 251 1379 252
rect 1383 251 1384 255
rect 1378 250 1384 251
rect 1387 255 1393 256
rect 1387 251 1388 255
rect 1392 254 1393 255
rect 1422 255 1428 256
rect 1422 254 1423 255
rect 1392 252 1423 254
rect 1392 251 1393 252
rect 1387 250 1393 251
rect 1422 251 1423 252
rect 1427 251 1428 255
rect 1422 250 1428 251
rect 1451 255 1457 256
rect 1451 251 1452 255
rect 1456 254 1457 255
rect 1510 255 1516 256
rect 1510 254 1511 255
rect 1456 252 1511 254
rect 1456 251 1457 252
rect 1451 250 1457 251
rect 1510 251 1511 252
rect 1515 251 1516 255
rect 1510 250 1516 251
rect 1518 255 1529 256
rect 1518 251 1519 255
rect 1523 251 1524 255
rect 1528 251 1529 255
rect 1603 253 1604 257
rect 1608 253 1609 257
rect 1603 252 1609 253
rect 1634 255 1640 256
rect 1518 250 1529 251
rect 1634 251 1635 255
rect 1639 254 1640 255
rect 1683 255 1689 256
rect 1683 254 1684 255
rect 1639 252 1684 254
rect 1639 251 1640 252
rect 1634 250 1640 251
rect 1683 251 1684 252
rect 1688 251 1689 255
rect 1683 250 1689 251
rect 1714 255 1720 256
rect 1714 251 1715 255
rect 1719 254 1720 255
rect 1763 255 1769 256
rect 1763 254 1764 255
rect 1719 252 1764 254
rect 1719 251 1720 252
rect 1714 250 1720 251
rect 1763 251 1764 252
rect 1768 251 1769 255
rect 1763 250 1769 251
rect 1835 255 1841 256
rect 1835 251 1836 255
rect 1840 254 1841 255
rect 1906 255 1912 256
rect 1906 254 1907 255
rect 1840 252 1907 254
rect 1840 251 1841 252
rect 1835 250 1841 251
rect 1906 251 1907 252
rect 1911 251 1912 255
rect 1906 250 1912 251
rect 1915 255 1921 256
rect 1915 251 1916 255
rect 1920 254 1921 255
rect 1974 255 1980 256
rect 1974 254 1975 255
rect 1920 252 1975 254
rect 1920 251 1921 252
rect 1915 250 1921 251
rect 1974 251 1975 252
rect 1979 251 1980 255
rect 1974 250 1980 251
rect 1995 255 2001 256
rect 1995 251 1996 255
rect 2000 254 2001 255
rect 2006 255 2012 256
rect 2006 254 2007 255
rect 2000 252 2007 254
rect 2000 251 2001 252
rect 1995 250 2001 251
rect 2006 251 2007 252
rect 2011 251 2012 255
rect 2006 250 2012 251
rect 2026 255 2032 256
rect 2026 251 2027 255
rect 2031 254 2032 255
rect 2067 255 2073 256
rect 2067 254 2068 255
rect 2031 252 2068 254
rect 2031 251 2032 252
rect 2026 250 2032 251
rect 2067 251 2068 252
rect 2072 251 2073 255
rect 2067 250 2073 251
rect 878 247 884 248
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 110 239 116 240
rect 142 239 148 240
rect 142 235 143 239
rect 147 238 148 239
rect 159 239 165 240
rect 159 238 160 239
rect 147 236 160 238
rect 147 235 148 236
rect 142 234 148 235
rect 159 235 160 236
rect 164 235 165 239
rect 159 234 165 235
rect 186 239 192 240
rect 186 235 187 239
rect 191 238 192 239
rect 223 239 229 240
rect 223 238 224 239
rect 191 236 224 238
rect 191 235 192 236
rect 186 234 192 235
rect 223 235 224 236
rect 228 235 229 239
rect 223 234 229 235
rect 266 239 272 240
rect 266 235 267 239
rect 271 238 272 239
rect 303 239 309 240
rect 303 238 304 239
rect 271 236 304 238
rect 271 235 272 236
rect 266 234 272 235
rect 303 235 304 236
rect 308 235 309 239
rect 303 234 309 235
rect 383 239 392 240
rect 383 235 384 239
rect 391 235 392 239
rect 383 234 392 235
rect 463 239 469 240
rect 463 235 464 239
rect 468 238 469 239
rect 471 239 477 240
rect 471 238 472 239
rect 468 236 472 238
rect 468 235 469 236
rect 463 234 469 235
rect 471 235 472 236
rect 476 235 477 239
rect 471 234 477 235
rect 535 239 544 240
rect 535 235 536 239
rect 543 235 544 239
rect 535 234 544 235
rect 607 239 616 240
rect 607 235 608 239
rect 615 235 616 239
rect 607 234 616 235
rect 671 239 677 240
rect 671 235 672 239
rect 676 238 677 239
rect 679 239 685 240
rect 679 238 680 239
rect 676 236 680 238
rect 676 235 677 236
rect 671 234 677 235
rect 679 235 680 236
rect 684 235 685 239
rect 679 234 685 235
rect 727 239 736 240
rect 727 235 728 239
rect 735 235 736 239
rect 727 234 736 235
rect 783 239 792 240
rect 783 235 784 239
rect 791 235 792 239
rect 783 234 792 235
rect 839 239 848 240
rect 839 235 840 239
rect 847 235 848 239
rect 839 234 848 235
rect 903 239 912 240
rect 1094 239 1100 240
rect 1158 244 1164 245
rect 1158 240 1159 244
rect 1163 240 1164 244
rect 1158 239 1164 240
rect 1206 244 1212 245
rect 1206 240 1207 244
rect 1211 240 1212 244
rect 1206 239 1212 240
rect 1270 244 1276 245
rect 1270 240 1271 244
rect 1275 240 1276 244
rect 1270 239 1276 240
rect 1326 244 1332 245
rect 1326 240 1327 244
rect 1331 240 1332 244
rect 1326 239 1332 240
rect 1390 244 1396 245
rect 1390 240 1391 244
rect 1395 240 1396 244
rect 1390 239 1396 240
rect 1454 244 1460 245
rect 1454 240 1455 244
rect 1459 240 1460 244
rect 1454 239 1460 240
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1606 244 1612 245
rect 1606 240 1607 244
rect 1611 240 1612 244
rect 1606 239 1612 240
rect 1686 244 1692 245
rect 1686 240 1687 244
rect 1691 240 1692 244
rect 1686 239 1692 240
rect 1766 244 1772 245
rect 1766 240 1767 244
rect 1771 240 1772 244
rect 1766 239 1772 240
rect 1838 244 1844 245
rect 1838 240 1839 244
rect 1843 240 1844 244
rect 1838 239 1844 240
rect 1918 244 1924 245
rect 1918 240 1919 244
rect 1923 240 1924 244
rect 1918 239 1924 240
rect 1998 244 2004 245
rect 1998 240 1999 244
rect 2003 240 2004 244
rect 1998 239 2004 240
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 903 235 904 239
rect 911 235 912 239
rect 903 234 912 235
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 1134 231 1140 232
rect 1183 231 1192 232
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1094 227 1100 228
rect 110 222 116 223
rect 134 224 140 225
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 198 224 204 225
rect 198 220 199 224
rect 203 220 204 224
rect 198 219 204 220
rect 278 224 284 225
rect 278 220 279 224
rect 283 220 284 224
rect 278 219 284 220
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 438 224 444 225
rect 438 220 439 224
rect 443 220 444 224
rect 438 219 444 220
rect 510 224 516 225
rect 510 220 511 224
rect 515 220 516 224
rect 510 219 516 220
rect 582 224 588 225
rect 582 220 583 224
rect 587 220 588 224
rect 582 219 588 220
rect 646 224 652 225
rect 646 220 647 224
rect 651 220 652 224
rect 646 219 652 220
rect 702 224 708 225
rect 702 220 703 224
rect 707 220 708 224
rect 702 219 708 220
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 878 224 884 225
rect 878 220 879 224
rect 883 220 884 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1183 227 1184 231
rect 1191 227 1192 231
rect 1183 226 1192 227
rect 1231 231 1240 232
rect 1231 227 1232 231
rect 1239 227 1240 231
rect 1231 226 1240 227
rect 1278 231 1284 232
rect 1278 227 1279 231
rect 1283 230 1284 231
rect 1295 231 1301 232
rect 1295 230 1296 231
rect 1283 228 1296 230
rect 1283 227 1284 228
rect 1278 226 1284 227
rect 1295 227 1296 228
rect 1300 227 1301 231
rect 1295 226 1301 227
rect 1350 231 1357 232
rect 1350 227 1351 231
rect 1356 227 1357 231
rect 1350 226 1357 227
rect 1378 231 1384 232
rect 1378 227 1379 231
rect 1383 230 1384 231
rect 1415 231 1421 232
rect 1415 230 1416 231
rect 1383 228 1416 230
rect 1383 227 1384 228
rect 1378 226 1384 227
rect 1415 227 1416 228
rect 1420 227 1421 231
rect 1415 226 1421 227
rect 1478 231 1485 232
rect 1478 227 1479 231
rect 1484 227 1485 231
rect 1478 226 1485 227
rect 1510 231 1516 232
rect 1510 227 1511 231
rect 1515 230 1516 231
rect 1551 231 1557 232
rect 1551 230 1552 231
rect 1515 228 1552 230
rect 1515 227 1516 228
rect 1510 226 1516 227
rect 1551 227 1552 228
rect 1556 227 1557 231
rect 1551 226 1557 227
rect 1631 231 1640 232
rect 1631 227 1632 231
rect 1639 227 1640 231
rect 1631 226 1640 227
rect 1711 231 1720 232
rect 1711 227 1712 231
rect 1719 227 1720 231
rect 1711 226 1720 227
rect 1742 231 1748 232
rect 1742 227 1743 231
rect 1747 230 1748 231
rect 1791 231 1797 232
rect 1791 230 1792 231
rect 1747 228 1792 230
rect 1747 227 1748 228
rect 1742 226 1748 227
rect 1791 227 1792 228
rect 1796 227 1797 231
rect 1791 226 1797 227
rect 1862 231 1869 232
rect 1862 227 1863 231
rect 1868 227 1869 231
rect 1862 226 1869 227
rect 1906 231 1912 232
rect 1906 227 1907 231
rect 1911 230 1912 231
rect 1943 231 1949 232
rect 1943 230 1944 231
rect 1911 228 1944 230
rect 1911 227 1912 228
rect 1906 226 1912 227
rect 1943 227 1944 228
rect 1948 227 1949 231
rect 1943 226 1949 227
rect 2023 231 2032 232
rect 2023 227 2024 231
rect 2031 227 2032 231
rect 2023 226 2032 227
rect 2086 231 2092 232
rect 2086 227 2087 231
rect 2091 230 2092 231
rect 2095 231 2101 232
rect 2118 231 2124 232
rect 2095 230 2096 231
rect 2091 228 2096 230
rect 2091 227 2092 228
rect 2086 226 2092 227
rect 2095 227 2096 228
rect 2100 227 2101 231
rect 2095 226 2101 227
rect 1094 222 1100 223
rect 878 219 884 220
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 2118 219 2124 220
rect 1134 214 1140 215
rect 1158 216 1164 217
rect 1158 212 1159 216
rect 1163 212 1164 216
rect 1158 211 1164 212
rect 1206 216 1212 217
rect 1206 212 1207 216
rect 1211 212 1212 216
rect 1206 211 1212 212
rect 1270 216 1276 217
rect 1270 212 1271 216
rect 1275 212 1276 216
rect 1270 211 1276 212
rect 1326 216 1332 217
rect 1326 212 1327 216
rect 1331 212 1332 216
rect 1326 211 1332 212
rect 1390 216 1396 217
rect 1390 212 1391 216
rect 1395 212 1396 216
rect 1390 211 1396 212
rect 1454 216 1460 217
rect 1454 212 1455 216
rect 1459 212 1460 216
rect 1454 211 1460 212
rect 1526 216 1532 217
rect 1526 212 1527 216
rect 1531 212 1532 216
rect 1526 211 1532 212
rect 1606 216 1612 217
rect 1606 212 1607 216
rect 1611 212 1612 216
rect 1606 211 1612 212
rect 1686 216 1692 217
rect 1686 212 1687 216
rect 1691 212 1692 216
rect 1686 211 1692 212
rect 1766 216 1772 217
rect 1766 212 1767 216
rect 1771 212 1772 216
rect 1766 211 1772 212
rect 1838 216 1844 217
rect 1838 212 1839 216
rect 1843 212 1844 216
rect 1838 211 1844 212
rect 1918 216 1924 217
rect 1918 212 1919 216
rect 1923 212 1924 216
rect 1918 211 1924 212
rect 1998 216 2004 217
rect 1998 212 1999 216
rect 2003 212 2004 216
rect 1998 211 2004 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2070 211 2076 212
rect 134 208 140 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 134 204 135 208
rect 139 204 140 208
rect 134 203 140 204
rect 182 208 188 209
rect 182 204 183 208
rect 187 204 188 208
rect 182 203 188 204
rect 230 208 236 209
rect 230 204 231 208
rect 235 204 236 208
rect 230 203 236 204
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 326 208 332 209
rect 326 204 327 208
rect 331 204 332 208
rect 326 203 332 204
rect 374 208 380 209
rect 374 204 375 208
rect 379 204 380 208
rect 374 203 380 204
rect 414 208 420 209
rect 414 204 415 208
rect 419 204 420 208
rect 414 203 420 204
rect 454 208 460 209
rect 454 204 455 208
rect 459 204 460 208
rect 454 203 460 204
rect 502 208 508 209
rect 502 204 503 208
rect 507 204 508 208
rect 502 203 508 204
rect 550 208 556 209
rect 550 204 551 208
rect 555 204 556 208
rect 550 203 556 204
rect 598 208 604 209
rect 598 204 599 208
rect 603 204 604 208
rect 598 203 604 204
rect 646 208 652 209
rect 646 204 647 208
rect 651 204 652 208
rect 646 203 652 204
rect 694 208 700 209
rect 694 204 695 208
rect 699 204 700 208
rect 694 203 700 204
rect 742 208 748 209
rect 742 204 743 208
rect 747 204 748 208
rect 742 203 748 204
rect 1094 205 1100 206
rect 110 200 116 201
rect 1094 201 1095 205
rect 1099 201 1100 205
rect 1158 204 1164 205
rect 1094 200 1100 201
rect 1134 201 1140 202
rect 590 199 596 200
rect 590 195 591 199
rect 595 198 596 199
rect 595 196 746 198
rect 1134 197 1135 201
rect 1139 197 1140 201
rect 1158 200 1159 204
rect 1163 200 1164 204
rect 1158 199 1164 200
rect 1198 204 1204 205
rect 1198 200 1199 204
rect 1203 200 1204 204
rect 1198 199 1204 200
rect 1262 204 1268 205
rect 1262 200 1263 204
rect 1267 200 1268 204
rect 1262 199 1268 200
rect 1326 204 1332 205
rect 1326 200 1327 204
rect 1331 200 1332 204
rect 1326 199 1332 200
rect 1398 204 1404 205
rect 1398 200 1399 204
rect 1403 200 1404 204
rect 1398 199 1404 200
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1542 204 1548 205
rect 1542 200 1543 204
rect 1547 200 1548 204
rect 1542 199 1548 200
rect 1606 204 1612 205
rect 1606 200 1607 204
rect 1611 200 1612 204
rect 1606 199 1612 200
rect 1670 204 1676 205
rect 1670 200 1671 204
rect 1675 200 1676 204
rect 1670 199 1676 200
rect 1734 204 1740 205
rect 1734 200 1735 204
rect 1739 200 1740 204
rect 1734 199 1740 200
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1878 204 1884 205
rect 1878 200 1879 204
rect 1883 200 1884 204
rect 1878 199 1884 200
rect 1950 204 1956 205
rect 1950 200 1951 204
rect 1955 200 1956 204
rect 1950 199 1956 200
rect 2022 204 2028 205
rect 2022 200 2023 204
rect 2027 200 2028 204
rect 2022 199 2028 200
rect 2070 204 2076 205
rect 2070 200 2071 204
rect 2075 200 2076 204
rect 2070 199 2076 200
rect 2118 201 2124 202
rect 1134 196 1140 197
rect 2118 197 2119 201
rect 2123 197 2124 201
rect 2118 196 2124 197
rect 595 195 596 196
rect 590 194 596 195
rect 159 191 165 192
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 159 187 160 191
rect 164 190 165 191
rect 174 191 180 192
rect 174 190 175 191
rect 164 188 175 190
rect 164 187 165 188
rect 159 186 165 187
rect 174 187 175 188
rect 179 187 180 191
rect 174 186 180 187
rect 207 191 213 192
rect 207 187 208 191
rect 212 190 213 191
rect 222 191 228 192
rect 222 190 223 191
rect 212 188 223 190
rect 212 187 213 188
rect 207 186 213 187
rect 222 187 223 188
rect 227 187 228 191
rect 222 186 228 187
rect 255 191 261 192
rect 255 187 256 191
rect 260 190 261 191
rect 270 191 276 192
rect 270 190 271 191
rect 260 188 271 190
rect 260 187 261 188
rect 255 186 261 187
rect 270 187 271 188
rect 275 187 276 191
rect 270 186 276 187
rect 286 191 292 192
rect 286 187 287 191
rect 291 190 292 191
rect 303 191 309 192
rect 303 190 304 191
rect 291 188 304 190
rect 291 187 292 188
rect 286 186 292 187
rect 303 187 304 188
rect 308 187 309 191
rect 303 186 309 187
rect 350 191 357 192
rect 350 187 351 191
rect 356 187 357 191
rect 350 186 357 187
rect 359 191 365 192
rect 359 187 360 191
rect 364 190 365 191
rect 399 191 405 192
rect 399 190 400 191
rect 364 188 400 190
rect 364 187 365 188
rect 359 186 365 187
rect 399 187 400 188
rect 404 187 405 191
rect 439 191 445 192
rect 439 190 440 191
rect 399 186 405 187
rect 408 188 440 190
rect 110 183 116 184
rect 134 180 140 181
rect 134 176 135 180
rect 139 176 140 180
rect 134 175 140 176
rect 182 180 188 181
rect 182 176 183 180
rect 187 176 188 180
rect 182 175 188 176
rect 230 180 236 181
rect 230 176 231 180
rect 235 176 236 180
rect 230 175 236 176
rect 278 180 284 181
rect 278 176 279 180
rect 283 176 284 180
rect 278 175 284 176
rect 326 180 332 181
rect 326 176 327 180
rect 331 176 332 180
rect 326 175 332 176
rect 374 180 380 181
rect 374 176 375 180
rect 379 176 380 180
rect 374 175 380 176
rect 408 174 410 188
rect 439 187 440 188
rect 444 187 445 191
rect 439 186 445 187
rect 479 191 485 192
rect 479 187 480 191
rect 484 190 485 191
rect 494 191 500 192
rect 494 190 495 191
rect 484 188 495 190
rect 484 187 485 188
rect 479 186 485 187
rect 494 187 495 188
rect 499 187 500 191
rect 494 186 500 187
rect 527 191 533 192
rect 527 187 528 191
rect 532 190 533 191
rect 542 191 548 192
rect 542 190 543 191
rect 532 188 543 190
rect 532 187 533 188
rect 527 186 533 187
rect 542 187 543 188
rect 547 187 548 191
rect 542 186 548 187
rect 575 191 581 192
rect 575 187 576 191
rect 580 190 581 191
rect 590 191 596 192
rect 590 190 591 191
rect 580 188 591 190
rect 580 187 581 188
rect 575 186 581 187
rect 590 187 591 188
rect 595 187 596 191
rect 590 186 596 187
rect 623 191 629 192
rect 623 187 624 191
rect 628 190 629 191
rect 638 191 644 192
rect 638 190 639 191
rect 628 188 639 190
rect 628 187 629 188
rect 623 186 629 187
rect 638 187 639 188
rect 643 187 644 191
rect 638 186 644 187
rect 671 191 677 192
rect 671 187 672 191
rect 676 190 677 191
rect 686 191 692 192
rect 686 190 687 191
rect 676 188 687 190
rect 676 187 677 188
rect 671 186 677 187
rect 686 187 687 188
rect 691 187 692 191
rect 686 186 692 187
rect 719 191 725 192
rect 719 187 720 191
rect 724 190 725 191
rect 734 191 740 192
rect 734 190 735 191
rect 724 188 735 190
rect 724 187 725 188
rect 719 186 725 187
rect 734 187 735 188
rect 739 187 740 191
rect 744 190 746 196
rect 1974 195 1980 196
rect 767 191 773 192
rect 767 190 768 191
rect 744 188 768 190
rect 734 186 740 187
rect 767 187 768 188
rect 772 187 773 191
rect 1974 191 1975 195
rect 1979 194 1980 195
rect 1979 192 2026 194
rect 1979 191 1980 192
rect 1974 190 1980 191
rect 767 186 773 187
rect 1094 188 1100 189
rect 1094 184 1095 188
rect 1099 184 1100 188
rect 1170 187 1176 188
rect 1094 183 1100 184
rect 1134 184 1140 185
rect 414 180 420 181
rect 414 176 415 180
rect 419 176 420 180
rect 414 175 420 176
rect 454 180 460 181
rect 454 176 455 180
rect 459 176 460 180
rect 454 175 460 176
rect 502 180 508 181
rect 502 176 503 180
rect 507 176 508 180
rect 502 175 508 176
rect 550 180 556 181
rect 550 176 551 180
rect 555 176 556 180
rect 550 175 556 176
rect 598 180 604 181
rect 598 176 599 180
rect 603 176 604 180
rect 598 175 604 176
rect 646 180 652 181
rect 646 176 647 180
rect 651 176 652 180
rect 646 175 652 176
rect 694 180 700 181
rect 694 176 695 180
rect 699 176 700 180
rect 694 175 700 176
rect 742 180 748 181
rect 742 176 743 180
rect 747 176 748 180
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1170 183 1171 187
rect 1175 186 1176 187
rect 1183 187 1189 188
rect 1183 186 1184 187
rect 1175 184 1184 186
rect 1175 183 1176 184
rect 1170 182 1176 183
rect 1183 183 1184 184
rect 1188 183 1189 187
rect 1223 187 1229 188
rect 1223 186 1224 187
rect 1183 182 1189 183
rect 1192 184 1224 186
rect 1134 179 1140 180
rect 742 175 748 176
rect 1158 176 1164 177
rect 400 172 410 174
rect 1158 172 1159 176
rect 1163 172 1164 176
rect 400 170 402 172
rect 1158 171 1164 172
rect 1192 170 1194 184
rect 1223 183 1224 184
rect 1228 183 1229 187
rect 1223 182 1229 183
rect 1231 187 1237 188
rect 1231 183 1232 187
rect 1236 186 1237 187
rect 1287 187 1293 188
rect 1287 186 1288 187
rect 1236 184 1288 186
rect 1236 183 1237 184
rect 1231 182 1237 183
rect 1287 183 1288 184
rect 1292 183 1293 187
rect 1287 182 1293 183
rect 1351 187 1357 188
rect 1351 183 1352 187
rect 1356 186 1357 187
rect 1390 187 1396 188
rect 1390 186 1391 187
rect 1356 184 1391 186
rect 1356 183 1357 184
rect 1351 182 1357 183
rect 1390 183 1391 184
rect 1395 183 1396 187
rect 1390 182 1396 183
rect 1422 187 1429 188
rect 1422 183 1423 187
rect 1428 183 1429 187
rect 1422 182 1429 183
rect 1495 187 1501 188
rect 1495 183 1496 187
rect 1500 186 1501 187
rect 1534 187 1540 188
rect 1534 186 1535 187
rect 1500 184 1535 186
rect 1500 183 1501 184
rect 1495 182 1501 183
rect 1534 183 1535 184
rect 1539 183 1540 187
rect 1534 182 1540 183
rect 1550 187 1556 188
rect 1550 183 1551 187
rect 1555 186 1556 187
rect 1567 187 1573 188
rect 1567 186 1568 187
rect 1555 184 1568 186
rect 1555 183 1556 184
rect 1550 182 1556 183
rect 1567 183 1568 184
rect 1572 183 1573 187
rect 1567 182 1573 183
rect 1578 187 1584 188
rect 1578 183 1579 187
rect 1583 186 1584 187
rect 1631 187 1637 188
rect 1631 186 1632 187
rect 1583 184 1632 186
rect 1583 183 1584 184
rect 1578 182 1584 183
rect 1631 183 1632 184
rect 1636 183 1637 187
rect 1631 182 1637 183
rect 1639 187 1645 188
rect 1639 183 1640 187
rect 1644 186 1645 187
rect 1695 187 1701 188
rect 1695 186 1696 187
rect 1644 184 1696 186
rect 1644 183 1645 184
rect 1639 182 1645 183
rect 1695 183 1696 184
rect 1700 183 1701 187
rect 1695 182 1701 183
rect 1703 187 1709 188
rect 1703 183 1704 187
rect 1708 186 1709 187
rect 1759 187 1765 188
rect 1759 186 1760 187
rect 1708 184 1760 186
rect 1708 183 1709 184
rect 1703 182 1709 183
rect 1759 183 1760 184
rect 1764 183 1765 187
rect 1759 182 1765 183
rect 1831 187 1837 188
rect 1831 183 1832 187
rect 1836 186 1837 187
rect 1870 187 1876 188
rect 1870 186 1871 187
rect 1836 184 1871 186
rect 1836 183 1837 184
rect 1831 182 1837 183
rect 1870 183 1871 184
rect 1875 183 1876 187
rect 1870 182 1876 183
rect 1903 187 1909 188
rect 1903 183 1904 187
rect 1908 186 1909 187
rect 1942 187 1948 188
rect 1942 186 1943 187
rect 1908 184 1943 186
rect 1908 183 1909 184
rect 1903 182 1909 183
rect 1942 183 1943 184
rect 1947 183 1948 187
rect 1942 182 1948 183
rect 1975 187 1981 188
rect 1975 183 1976 187
rect 1980 186 1981 187
rect 2014 187 2020 188
rect 2014 186 2015 187
rect 1980 184 2015 186
rect 1980 183 1981 184
rect 1975 182 1981 183
rect 2014 183 2015 184
rect 2019 183 2020 187
rect 2024 186 2026 192
rect 2047 187 2053 188
rect 2047 186 2048 187
rect 2024 184 2048 186
rect 2014 182 2020 183
rect 2047 183 2048 184
rect 2052 183 2053 187
rect 2047 182 2053 183
rect 2078 187 2084 188
rect 2078 183 2079 187
rect 2083 186 2084 187
rect 2095 187 2101 188
rect 2095 186 2096 187
rect 2083 184 2096 186
rect 2083 183 2084 184
rect 2078 182 2084 183
rect 2095 183 2096 184
rect 2100 183 2101 187
rect 2095 182 2101 183
rect 2118 184 2124 185
rect 2118 180 2119 184
rect 2123 180 2124 184
rect 2118 179 2124 180
rect 1198 176 1204 177
rect 1198 172 1199 176
rect 1203 172 1204 176
rect 1198 171 1204 172
rect 1262 176 1268 177
rect 1262 172 1263 176
rect 1267 172 1268 176
rect 1262 171 1268 172
rect 1326 176 1332 177
rect 1326 172 1327 176
rect 1331 172 1332 176
rect 1326 171 1332 172
rect 1398 176 1404 177
rect 1398 172 1399 176
rect 1403 172 1404 176
rect 1398 171 1404 172
rect 1470 176 1476 177
rect 1470 172 1471 176
rect 1475 172 1476 176
rect 1470 171 1476 172
rect 1542 176 1548 177
rect 1542 172 1543 176
rect 1547 172 1548 176
rect 1542 171 1548 172
rect 1606 176 1612 177
rect 1606 172 1607 176
rect 1611 172 1612 176
rect 1606 171 1612 172
rect 1670 176 1676 177
rect 1670 172 1671 176
rect 1675 172 1676 176
rect 1670 171 1676 172
rect 1734 176 1740 177
rect 1734 172 1735 176
rect 1739 172 1740 176
rect 1734 171 1740 172
rect 1806 176 1812 177
rect 1806 172 1807 176
rect 1811 172 1812 176
rect 1806 171 1812 172
rect 1878 176 1884 177
rect 1878 172 1879 176
rect 1883 172 1884 176
rect 1878 171 1884 172
rect 1950 176 1956 177
rect 1950 172 1951 176
rect 1955 172 1956 176
rect 1950 171 1956 172
rect 2022 176 2028 177
rect 2022 172 2023 176
rect 2027 172 2028 176
rect 2022 171 2028 172
rect 2070 176 2076 177
rect 2070 172 2071 176
rect 2075 172 2076 176
rect 2070 171 2076 172
rect 371 169 402 170
rect 131 167 137 168
rect 131 163 132 167
rect 136 166 137 167
rect 142 167 148 168
rect 142 166 143 167
rect 136 164 143 166
rect 136 163 137 164
rect 131 162 137 163
rect 142 163 143 164
rect 147 163 148 167
rect 142 162 148 163
rect 174 167 185 168
rect 174 163 175 167
rect 179 163 180 167
rect 184 163 185 167
rect 174 162 185 163
rect 222 167 233 168
rect 222 163 223 167
rect 227 163 228 167
rect 232 163 233 167
rect 222 162 233 163
rect 270 167 281 168
rect 270 163 271 167
rect 275 163 276 167
rect 280 163 281 167
rect 270 162 281 163
rect 323 167 329 168
rect 323 163 324 167
rect 328 166 329 167
rect 359 167 365 168
rect 359 166 360 167
rect 328 164 360 166
rect 328 163 329 164
rect 323 162 329 163
rect 359 163 360 164
rect 364 163 365 167
rect 371 165 372 169
rect 376 168 402 169
rect 1188 168 1194 170
rect 376 165 377 168
rect 371 164 377 165
rect 411 167 417 168
rect 359 162 365 163
rect 411 163 412 167
rect 416 166 417 167
rect 451 167 457 168
rect 416 164 446 166
rect 416 163 417 164
rect 411 162 417 163
rect 444 150 446 164
rect 451 163 452 167
rect 456 166 457 167
rect 494 167 505 168
rect 456 164 490 166
rect 456 163 457 164
rect 451 162 457 163
rect 488 158 490 164
rect 494 163 495 167
rect 499 163 500 167
rect 504 163 505 167
rect 494 162 505 163
rect 542 167 553 168
rect 542 163 543 167
rect 547 163 548 167
rect 552 163 553 167
rect 542 162 553 163
rect 590 167 601 168
rect 590 163 591 167
rect 595 163 596 167
rect 600 163 601 167
rect 590 162 601 163
rect 638 167 649 168
rect 638 163 639 167
rect 643 163 644 167
rect 648 163 649 167
rect 638 162 649 163
rect 686 167 697 168
rect 686 163 687 167
rect 691 163 692 167
rect 696 163 697 167
rect 686 162 697 163
rect 734 167 745 168
rect 734 163 735 167
rect 739 163 740 167
rect 744 163 745 167
rect 1188 166 1190 168
rect 734 162 745 163
rect 1155 165 1190 166
rect 1155 161 1156 165
rect 1160 164 1190 165
rect 1160 161 1161 164
rect 1155 160 1161 161
rect 1195 163 1201 164
rect 566 159 572 160
rect 566 158 567 159
rect 488 156 567 158
rect 566 155 567 156
rect 571 155 572 159
rect 1195 159 1196 163
rect 1200 162 1201 163
rect 1231 163 1237 164
rect 1231 162 1232 163
rect 1200 160 1232 162
rect 1200 159 1201 160
rect 1195 158 1201 159
rect 1231 159 1232 160
rect 1236 159 1237 163
rect 1231 158 1237 159
rect 1259 163 1265 164
rect 1259 159 1260 163
rect 1264 162 1265 163
rect 1278 163 1284 164
rect 1278 162 1279 163
rect 1264 160 1279 162
rect 1264 159 1265 160
rect 1259 158 1265 159
rect 1278 159 1279 160
rect 1283 159 1284 163
rect 1278 158 1284 159
rect 1298 163 1304 164
rect 1298 159 1299 163
rect 1303 162 1304 163
rect 1323 163 1329 164
rect 1323 162 1324 163
rect 1303 160 1324 162
rect 1303 159 1304 160
rect 1298 158 1304 159
rect 1323 159 1324 160
rect 1328 159 1329 163
rect 1323 158 1329 159
rect 1390 163 1401 164
rect 1390 159 1391 163
rect 1395 159 1396 163
rect 1400 159 1401 163
rect 1390 158 1401 159
rect 1467 163 1473 164
rect 1467 159 1468 163
rect 1472 162 1473 163
rect 1478 163 1484 164
rect 1478 162 1479 163
rect 1472 160 1479 162
rect 1472 159 1473 160
rect 1467 158 1473 159
rect 1478 159 1479 160
rect 1483 159 1484 163
rect 1478 158 1484 159
rect 1534 163 1545 164
rect 1534 159 1535 163
rect 1539 159 1540 163
rect 1544 159 1545 163
rect 1534 158 1545 159
rect 1603 163 1609 164
rect 1603 159 1604 163
rect 1608 162 1609 163
rect 1639 163 1645 164
rect 1639 162 1640 163
rect 1608 160 1640 162
rect 1608 159 1609 160
rect 1603 158 1609 159
rect 1639 159 1640 160
rect 1644 159 1645 163
rect 1639 158 1645 159
rect 1667 163 1673 164
rect 1667 159 1668 163
rect 1672 162 1673 163
rect 1703 163 1709 164
rect 1703 162 1704 163
rect 1672 160 1704 162
rect 1672 159 1673 160
rect 1667 158 1673 159
rect 1703 159 1704 160
rect 1708 159 1709 163
rect 1703 158 1709 159
rect 1731 163 1737 164
rect 1731 159 1732 163
rect 1736 162 1737 163
rect 1742 163 1748 164
rect 1742 162 1743 163
rect 1736 160 1743 162
rect 1736 159 1737 160
rect 1731 158 1737 159
rect 1742 159 1743 160
rect 1747 159 1748 163
rect 1742 158 1748 159
rect 1803 163 1809 164
rect 1803 159 1804 163
rect 1808 162 1809 163
rect 1870 163 1881 164
rect 1808 160 1866 162
rect 1808 159 1809 160
rect 1803 158 1809 159
rect 566 154 572 155
rect 1864 154 1866 160
rect 1870 159 1871 163
rect 1875 159 1876 163
rect 1880 159 1881 163
rect 1870 158 1881 159
rect 1942 163 1953 164
rect 1942 159 1943 163
rect 1947 159 1948 163
rect 1952 159 1953 163
rect 1942 158 1953 159
rect 2014 163 2025 164
rect 2014 159 2015 163
rect 2019 159 2020 163
rect 2024 159 2025 163
rect 2014 158 2025 159
rect 2067 163 2073 164
rect 2067 159 2068 163
rect 2072 162 2073 163
rect 2086 163 2092 164
rect 2086 162 2087 163
rect 2072 160 2087 162
rect 2072 159 2073 160
rect 2067 158 2073 159
rect 2086 159 2087 160
rect 2091 159 2092 163
rect 2086 158 2092 159
rect 1974 155 1980 156
rect 1974 154 1975 155
rect 1864 152 1975 154
rect 526 151 532 152
rect 526 150 527 151
rect 444 148 527 150
rect 526 147 527 148
rect 531 147 532 151
rect 1974 151 1975 152
rect 1979 151 1980 155
rect 1974 150 1980 151
rect 526 146 532 147
rect 286 139 292 140
rect 286 138 287 139
rect 140 136 287 138
rect 140 134 142 136
rect 286 135 287 136
rect 291 135 292 139
rect 1358 139 1364 140
rect 1358 138 1359 139
rect 286 134 292 135
rect 1204 136 1359 138
rect 1204 134 1206 136
rect 1358 135 1359 136
rect 1363 135 1364 139
rect 1550 139 1556 140
rect 1550 138 1551 139
rect 1358 134 1364 135
rect 1508 136 1551 138
rect 1508 134 1510 136
rect 1550 135 1551 136
rect 1555 135 1556 139
rect 1550 134 1556 135
rect 139 133 145 134
rect 139 129 140 133
rect 144 129 145 133
rect 1203 133 1209 134
rect 139 128 145 129
rect 170 131 176 132
rect 170 127 171 131
rect 175 130 176 131
rect 179 131 185 132
rect 179 130 180 131
rect 175 128 180 130
rect 175 127 176 128
rect 170 126 176 127
rect 179 127 180 128
rect 184 127 185 131
rect 179 126 185 127
rect 210 131 216 132
rect 210 127 211 131
rect 215 130 216 131
rect 219 131 225 132
rect 219 130 220 131
rect 215 128 220 130
rect 215 127 216 128
rect 210 126 216 127
rect 219 127 220 128
rect 224 127 225 131
rect 219 126 225 127
rect 246 131 252 132
rect 246 127 247 131
rect 251 130 252 131
rect 259 131 265 132
rect 259 130 260 131
rect 251 128 260 130
rect 251 127 252 128
rect 246 126 252 127
rect 259 127 260 128
rect 264 127 265 131
rect 259 126 265 127
rect 290 131 296 132
rect 290 127 291 131
rect 295 130 296 131
rect 299 131 305 132
rect 299 130 300 131
rect 295 128 300 130
rect 295 127 296 128
rect 290 126 296 127
rect 299 127 300 128
rect 304 127 305 131
rect 299 126 305 127
rect 334 131 345 132
rect 334 127 335 131
rect 339 127 340 131
rect 344 127 345 131
rect 334 126 345 127
rect 366 131 372 132
rect 366 127 367 131
rect 371 130 372 131
rect 379 131 385 132
rect 379 130 380 131
rect 371 128 380 130
rect 371 127 372 128
rect 366 126 372 127
rect 379 127 380 128
rect 384 127 385 131
rect 379 126 385 127
rect 406 131 412 132
rect 406 127 407 131
rect 411 130 412 131
rect 419 131 425 132
rect 419 130 420 131
rect 411 128 420 130
rect 411 127 412 128
rect 406 126 412 127
rect 419 127 420 128
rect 424 127 425 131
rect 419 126 425 127
rect 446 131 452 132
rect 446 127 447 131
rect 451 130 452 131
rect 459 131 465 132
rect 459 130 460 131
rect 451 128 460 130
rect 451 127 452 128
rect 446 126 452 127
rect 459 127 460 128
rect 464 127 465 131
rect 459 126 465 127
rect 490 131 496 132
rect 490 127 491 131
rect 495 130 496 131
rect 499 131 505 132
rect 499 130 500 131
rect 495 128 500 130
rect 495 127 496 128
rect 490 126 496 127
rect 499 127 500 128
rect 504 127 505 131
rect 499 126 505 127
rect 539 131 545 132
rect 539 127 540 131
rect 544 130 545 131
rect 579 131 585 132
rect 544 128 574 130
rect 544 127 545 128
rect 539 126 545 127
rect 142 120 148 121
rect 142 116 143 120
rect 147 116 148 120
rect 142 115 148 116
rect 182 120 188 121
rect 182 116 183 120
rect 187 116 188 120
rect 182 115 188 116
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 262 120 268 121
rect 262 116 263 120
rect 267 116 268 120
rect 262 115 268 116
rect 302 120 308 121
rect 302 116 303 120
rect 307 116 308 120
rect 302 115 308 116
rect 342 120 348 121
rect 342 116 343 120
rect 347 116 348 120
rect 342 115 348 116
rect 382 120 388 121
rect 382 116 383 120
rect 387 116 388 120
rect 382 115 388 116
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 462 120 468 121
rect 462 116 463 120
rect 467 116 468 120
rect 462 115 468 116
rect 502 120 508 121
rect 502 116 503 120
rect 507 116 508 120
rect 502 115 508 116
rect 542 120 548 121
rect 542 116 543 120
rect 547 116 548 120
rect 542 115 548 116
rect 572 114 574 128
rect 579 127 580 131
rect 584 130 585 131
rect 619 131 625 132
rect 584 128 614 130
rect 584 127 585 128
rect 579 126 585 127
rect 582 120 588 121
rect 582 116 583 120
rect 587 116 588 120
rect 582 115 588 116
rect 612 114 614 128
rect 619 127 620 131
rect 624 130 625 131
rect 659 131 665 132
rect 624 128 654 130
rect 624 127 625 128
rect 619 126 625 127
rect 622 120 628 121
rect 622 116 623 120
rect 627 116 628 120
rect 622 115 628 116
rect 652 114 654 128
rect 659 127 660 131
rect 664 130 665 131
rect 699 131 705 132
rect 664 128 694 130
rect 664 127 665 128
rect 659 126 665 127
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 692 114 694 128
rect 699 127 700 131
rect 704 130 705 131
rect 739 131 745 132
rect 704 128 734 130
rect 704 127 705 128
rect 699 126 705 127
rect 702 120 708 121
rect 702 116 703 120
rect 707 116 708 120
rect 702 115 708 116
rect 732 114 734 128
rect 739 127 740 131
rect 744 130 745 131
rect 779 131 785 132
rect 744 128 774 130
rect 744 127 745 128
rect 739 126 745 127
rect 742 120 748 121
rect 742 116 743 120
rect 747 116 748 120
rect 742 115 748 116
rect 772 114 774 128
rect 779 127 780 131
rect 784 130 785 131
rect 818 131 824 132
rect 818 130 819 131
rect 784 128 819 130
rect 784 127 785 128
rect 779 126 785 127
rect 818 127 819 128
rect 823 127 824 131
rect 818 126 824 127
rect 827 131 833 132
rect 827 127 828 131
rect 832 130 833 131
rect 866 131 872 132
rect 866 130 867 131
rect 832 128 867 130
rect 832 127 833 128
rect 827 126 833 127
rect 866 127 867 128
rect 871 127 872 131
rect 866 126 872 127
rect 875 131 881 132
rect 875 127 876 131
rect 880 130 881 131
rect 911 131 917 132
rect 911 130 912 131
rect 880 128 912 130
rect 880 127 881 128
rect 875 126 881 127
rect 911 127 912 128
rect 916 127 917 131
rect 911 126 917 127
rect 923 131 929 132
rect 923 127 924 131
rect 928 130 929 131
rect 963 131 969 132
rect 928 128 958 130
rect 928 127 929 128
rect 923 126 929 127
rect 782 120 788 121
rect 782 116 783 120
rect 787 116 788 120
rect 782 115 788 116
rect 830 120 836 121
rect 830 116 831 120
rect 835 116 836 120
rect 830 115 836 116
rect 878 120 884 121
rect 878 116 879 120
rect 883 116 884 120
rect 878 115 884 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 956 114 958 128
rect 963 127 964 131
rect 968 130 969 131
rect 1003 131 1009 132
rect 968 128 998 130
rect 968 127 969 128
rect 963 126 969 127
rect 966 120 972 121
rect 966 116 967 120
rect 971 116 972 120
rect 966 115 972 116
rect 996 114 998 128
rect 1003 127 1004 131
rect 1008 130 1009 131
rect 1043 131 1049 132
rect 1008 128 1038 130
rect 1008 127 1009 128
rect 1003 126 1009 127
rect 1006 120 1012 121
rect 1006 116 1007 120
rect 1011 116 1012 120
rect 1006 115 1012 116
rect 1036 114 1038 128
rect 1043 127 1044 131
rect 1048 130 1049 131
rect 1142 131 1148 132
rect 1142 130 1143 131
rect 1048 128 1143 130
rect 1048 127 1049 128
rect 1043 126 1049 127
rect 1142 127 1143 128
rect 1147 127 1148 131
rect 1142 126 1148 127
rect 1155 131 1161 132
rect 1155 127 1156 131
rect 1160 130 1161 131
rect 1170 131 1176 132
rect 1170 130 1171 131
rect 1160 128 1171 130
rect 1160 127 1161 128
rect 1155 126 1161 127
rect 1170 127 1171 128
rect 1175 127 1176 131
rect 1203 129 1204 133
rect 1208 129 1209 133
rect 1507 133 1513 134
rect 1203 128 1209 129
rect 1234 131 1240 132
rect 1170 126 1176 127
rect 1234 127 1235 131
rect 1239 130 1240 131
rect 1267 131 1273 132
rect 1267 130 1268 131
rect 1239 128 1268 130
rect 1239 127 1240 128
rect 1234 126 1240 127
rect 1267 127 1268 128
rect 1272 127 1273 131
rect 1267 126 1273 127
rect 1331 131 1337 132
rect 1331 127 1332 131
rect 1336 130 1337 131
rect 1386 131 1392 132
rect 1386 130 1387 131
rect 1336 128 1387 130
rect 1336 127 1337 128
rect 1331 126 1337 127
rect 1386 127 1387 128
rect 1391 127 1392 131
rect 1386 126 1392 127
rect 1395 131 1401 132
rect 1395 127 1396 131
rect 1400 130 1401 131
rect 1438 131 1444 132
rect 1438 130 1439 131
rect 1400 128 1439 130
rect 1400 127 1401 128
rect 1395 126 1401 127
rect 1438 127 1439 128
rect 1443 127 1444 131
rect 1438 126 1444 127
rect 1451 131 1457 132
rect 1451 127 1452 131
rect 1456 130 1457 131
rect 1498 131 1504 132
rect 1498 130 1499 131
rect 1456 128 1499 130
rect 1456 127 1457 128
rect 1451 126 1457 127
rect 1498 127 1499 128
rect 1503 127 1504 131
rect 1507 129 1508 133
rect 1512 129 1513 133
rect 1507 128 1513 129
rect 1555 131 1561 132
rect 1498 126 1504 127
rect 1555 127 1556 131
rect 1560 130 1561 131
rect 1578 131 1584 132
rect 1578 130 1579 131
rect 1560 128 1579 130
rect 1560 127 1561 128
rect 1555 126 1561 127
rect 1578 127 1579 128
rect 1583 127 1584 131
rect 1578 126 1584 127
rect 1586 131 1592 132
rect 1586 127 1587 131
rect 1591 130 1592 131
rect 1603 131 1609 132
rect 1603 130 1604 131
rect 1591 128 1604 130
rect 1591 127 1592 128
rect 1586 126 1592 127
rect 1603 127 1604 128
rect 1608 127 1609 131
rect 1603 126 1609 127
rect 1634 131 1640 132
rect 1634 127 1635 131
rect 1639 130 1640 131
rect 1643 131 1649 132
rect 1643 130 1644 131
rect 1639 128 1644 130
rect 1639 127 1640 128
rect 1634 126 1640 127
rect 1643 127 1644 128
rect 1648 127 1649 131
rect 1643 126 1649 127
rect 1678 131 1689 132
rect 1678 127 1679 131
rect 1683 127 1684 131
rect 1688 127 1689 131
rect 1678 126 1689 127
rect 1714 131 1720 132
rect 1714 127 1715 131
rect 1719 130 1720 131
rect 1723 131 1729 132
rect 1723 130 1724 131
rect 1719 128 1724 130
rect 1719 127 1720 128
rect 1714 126 1720 127
rect 1723 127 1724 128
rect 1728 127 1729 131
rect 1723 126 1729 127
rect 1754 131 1760 132
rect 1754 127 1755 131
rect 1759 130 1760 131
rect 1763 131 1769 132
rect 1763 130 1764 131
rect 1759 128 1764 130
rect 1759 127 1760 128
rect 1754 126 1760 127
rect 1763 127 1764 128
rect 1768 127 1769 131
rect 1763 126 1769 127
rect 1794 131 1800 132
rect 1794 127 1795 131
rect 1799 130 1800 131
rect 1803 131 1809 132
rect 1803 130 1804 131
rect 1799 128 1804 130
rect 1799 127 1800 128
rect 1794 126 1800 127
rect 1803 127 1804 128
rect 1808 127 1809 131
rect 1803 126 1809 127
rect 1834 131 1840 132
rect 1834 127 1835 131
rect 1839 130 1840 131
rect 1851 131 1857 132
rect 1851 130 1852 131
rect 1839 128 1852 130
rect 1839 127 1840 128
rect 1834 126 1840 127
rect 1851 127 1852 128
rect 1856 127 1857 131
rect 1851 126 1857 127
rect 1887 131 1893 132
rect 1887 127 1888 131
rect 1892 130 1893 131
rect 1899 131 1905 132
rect 1899 130 1900 131
rect 1892 128 1900 130
rect 1892 127 1893 128
rect 1887 126 1893 127
rect 1899 127 1900 128
rect 1904 127 1905 131
rect 1899 126 1905 127
rect 1930 131 1936 132
rect 1930 127 1931 131
rect 1935 130 1936 131
rect 1947 131 1953 132
rect 1947 130 1948 131
rect 1935 128 1948 130
rect 1935 127 1936 128
rect 1930 126 1936 127
rect 1947 127 1948 128
rect 1952 127 1953 131
rect 1947 126 1953 127
rect 1987 131 1993 132
rect 1987 127 1988 131
rect 1992 130 1993 131
rect 2014 131 2020 132
rect 2014 130 2015 131
rect 1992 128 2015 130
rect 1992 127 1993 128
rect 1987 126 1993 127
rect 2014 127 2015 128
rect 2019 127 2020 131
rect 2014 126 2020 127
rect 2027 131 2033 132
rect 2027 127 2028 131
rect 2032 130 2033 131
rect 2067 131 2073 132
rect 2032 128 2062 130
rect 2032 127 2033 128
rect 2027 126 2033 127
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1158 120 1164 121
rect 1158 116 1159 120
rect 1163 116 1164 120
rect 1158 115 1164 116
rect 1206 120 1212 121
rect 1206 116 1207 120
rect 1211 116 1212 120
rect 1206 115 1212 116
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1334 120 1340 121
rect 1334 116 1335 120
rect 1339 116 1340 120
rect 1334 115 1340 116
rect 1398 120 1404 121
rect 1398 116 1399 120
rect 1403 116 1404 120
rect 1398 115 1404 116
rect 1454 120 1460 121
rect 1454 116 1455 120
rect 1459 116 1460 120
rect 1454 115 1460 116
rect 1510 120 1516 121
rect 1510 116 1511 120
rect 1515 116 1516 120
rect 1510 115 1516 116
rect 1558 120 1564 121
rect 1558 116 1559 120
rect 1563 116 1564 120
rect 1558 115 1564 116
rect 1606 120 1612 121
rect 1606 116 1607 120
rect 1611 116 1612 120
rect 1606 115 1612 116
rect 1646 120 1652 121
rect 1646 116 1647 120
rect 1651 116 1652 120
rect 1646 115 1652 116
rect 1686 120 1692 121
rect 1686 116 1687 120
rect 1691 116 1692 120
rect 1686 115 1692 116
rect 1726 120 1732 121
rect 1726 116 1727 120
rect 1731 116 1732 120
rect 1726 115 1732 116
rect 1766 120 1772 121
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1854 120 1860 121
rect 1854 116 1855 120
rect 1859 116 1860 120
rect 1854 115 1860 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 1902 115 1908 116
rect 1950 120 1956 121
rect 1950 116 1951 120
rect 1955 116 1956 120
rect 1950 115 1956 116
rect 1990 120 1996 121
rect 1990 116 1991 120
rect 1995 116 1996 120
rect 1990 115 1996 116
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2030 115 2036 116
rect 2060 114 2062 128
rect 2067 127 2068 131
rect 2072 130 2073 131
rect 2078 131 2084 132
rect 2078 130 2079 131
rect 2072 128 2079 130
rect 2072 127 2073 128
rect 2067 126 2073 127
rect 2078 127 2079 128
rect 2083 127 2084 131
rect 2078 126 2084 127
rect 2070 120 2076 121
rect 2070 116 2071 120
rect 2075 116 2076 120
rect 2070 115 2076 116
rect 110 112 116 113
rect 572 112 578 114
rect 612 112 618 114
rect 652 112 658 114
rect 692 112 698 114
rect 732 112 738 114
rect 772 112 778 114
rect 956 112 962 114
rect 996 112 1002 114
rect 1036 112 1042 114
rect 110 108 111 112
rect 115 108 116 112
rect 110 107 116 108
rect 167 107 176 108
rect 167 103 168 107
rect 175 103 176 107
rect 167 102 176 103
rect 207 107 216 108
rect 207 103 208 107
rect 215 103 216 107
rect 207 102 216 103
rect 246 107 253 108
rect 246 103 247 107
rect 252 103 253 107
rect 246 102 253 103
rect 287 107 296 108
rect 287 103 288 107
rect 295 103 296 107
rect 287 102 296 103
rect 327 107 336 108
rect 327 103 328 107
rect 335 103 336 107
rect 327 102 336 103
rect 366 107 373 108
rect 366 103 367 107
rect 372 103 373 107
rect 366 102 373 103
rect 406 107 413 108
rect 406 103 407 107
rect 412 103 413 107
rect 406 102 413 103
rect 446 107 453 108
rect 446 103 447 107
rect 452 103 453 107
rect 446 102 453 103
rect 487 107 496 108
rect 487 103 488 107
rect 495 103 496 107
rect 487 102 496 103
rect 526 107 533 108
rect 526 103 527 107
rect 532 103 533 107
rect 526 102 533 103
rect 566 107 573 108
rect 566 103 567 107
rect 572 103 573 107
rect 576 106 578 112
rect 607 107 613 108
rect 607 106 608 107
rect 576 104 608 106
rect 566 102 573 103
rect 607 103 608 104
rect 612 103 613 107
rect 616 106 618 112
rect 647 107 653 108
rect 647 106 648 107
rect 616 104 648 106
rect 607 102 613 103
rect 647 103 648 104
rect 652 103 653 107
rect 656 106 658 112
rect 687 107 693 108
rect 687 106 688 107
rect 656 104 688 106
rect 647 102 653 103
rect 687 103 688 104
rect 692 103 693 107
rect 696 106 698 112
rect 727 107 733 108
rect 727 106 728 107
rect 696 104 728 106
rect 687 102 693 103
rect 727 103 728 104
rect 732 103 733 107
rect 736 106 738 112
rect 767 107 773 108
rect 767 106 768 107
rect 736 104 768 106
rect 727 102 733 103
rect 767 103 768 104
rect 772 103 773 107
rect 776 106 778 112
rect 807 107 813 108
rect 807 106 808 107
rect 776 104 808 106
rect 767 102 773 103
rect 807 103 808 104
rect 812 103 813 107
rect 807 102 813 103
rect 818 107 824 108
rect 818 103 819 107
rect 823 106 824 107
rect 855 107 861 108
rect 855 106 856 107
rect 823 104 856 106
rect 823 103 824 104
rect 818 102 824 103
rect 855 103 856 104
rect 860 103 861 107
rect 855 102 861 103
rect 866 107 872 108
rect 866 103 867 107
rect 871 106 872 107
rect 903 107 909 108
rect 903 106 904 107
rect 871 104 904 106
rect 871 103 872 104
rect 866 102 872 103
rect 903 103 904 104
rect 908 103 909 107
rect 903 102 909 103
rect 911 107 917 108
rect 911 103 912 107
rect 916 106 917 107
rect 951 107 957 108
rect 951 106 952 107
rect 916 104 952 106
rect 916 103 917 104
rect 911 102 917 103
rect 951 103 952 104
rect 956 103 957 107
rect 960 106 962 112
rect 991 107 997 108
rect 991 106 992 107
rect 960 104 992 106
rect 951 102 957 103
rect 991 103 992 104
rect 996 103 997 107
rect 1000 106 1002 112
rect 1031 107 1037 108
rect 1031 106 1032 107
rect 1000 104 1032 106
rect 991 102 997 103
rect 1031 103 1032 104
rect 1036 103 1037 107
rect 1040 106 1042 112
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 1071 107 1077 108
rect 1094 107 1100 108
rect 1134 112 1140 113
rect 2060 112 2066 114
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1134 107 1140 108
rect 1142 107 1148 108
rect 1071 106 1072 107
rect 1040 104 1072 106
rect 1031 102 1037 103
rect 1071 103 1072 104
rect 1076 103 1077 107
rect 1071 102 1077 103
rect 1142 103 1143 107
rect 1147 106 1148 107
rect 1183 107 1189 108
rect 1183 106 1184 107
rect 1147 104 1184 106
rect 1147 103 1148 104
rect 1142 102 1148 103
rect 1183 103 1184 104
rect 1188 103 1189 107
rect 1183 102 1189 103
rect 1231 107 1240 108
rect 1231 103 1232 107
rect 1239 103 1240 107
rect 1231 102 1240 103
rect 1295 107 1304 108
rect 1295 103 1296 107
rect 1303 103 1304 107
rect 1295 102 1304 103
rect 1358 107 1365 108
rect 1358 103 1359 107
rect 1364 103 1365 107
rect 1358 102 1365 103
rect 1386 107 1392 108
rect 1386 103 1387 107
rect 1391 106 1392 107
rect 1423 107 1429 108
rect 1423 106 1424 107
rect 1391 104 1424 106
rect 1391 103 1392 104
rect 1386 102 1392 103
rect 1423 103 1424 104
rect 1428 103 1429 107
rect 1423 102 1429 103
rect 1438 107 1444 108
rect 1438 103 1439 107
rect 1443 106 1444 107
rect 1479 107 1485 108
rect 1479 106 1480 107
rect 1443 104 1480 106
rect 1443 103 1444 104
rect 1438 102 1444 103
rect 1479 103 1480 104
rect 1484 103 1485 107
rect 1479 102 1485 103
rect 1498 107 1504 108
rect 1498 103 1499 107
rect 1503 106 1504 107
rect 1535 107 1541 108
rect 1535 106 1536 107
rect 1503 104 1536 106
rect 1503 103 1504 104
rect 1498 102 1504 103
rect 1535 103 1536 104
rect 1540 103 1541 107
rect 1535 102 1541 103
rect 1583 107 1592 108
rect 1583 103 1584 107
rect 1591 103 1592 107
rect 1583 102 1592 103
rect 1631 107 1640 108
rect 1631 103 1632 107
rect 1639 103 1640 107
rect 1631 102 1640 103
rect 1671 107 1680 108
rect 1671 103 1672 107
rect 1679 103 1680 107
rect 1671 102 1680 103
rect 1711 107 1720 108
rect 1711 103 1712 107
rect 1719 103 1720 107
rect 1711 102 1720 103
rect 1751 107 1760 108
rect 1751 103 1752 107
rect 1759 103 1760 107
rect 1751 102 1760 103
rect 1791 107 1800 108
rect 1791 103 1792 107
rect 1799 103 1800 107
rect 1791 102 1800 103
rect 1831 107 1840 108
rect 1831 103 1832 107
rect 1839 103 1840 107
rect 1831 102 1840 103
rect 1879 107 1885 108
rect 1879 103 1880 107
rect 1884 106 1885 107
rect 1887 107 1893 108
rect 1887 106 1888 107
rect 1884 104 1888 106
rect 1884 103 1885 104
rect 1879 102 1885 103
rect 1887 103 1888 104
rect 1892 103 1893 107
rect 1887 102 1893 103
rect 1927 107 1936 108
rect 1927 103 1928 107
rect 1935 103 1936 107
rect 1927 102 1936 103
rect 1974 107 1981 108
rect 1974 103 1975 107
rect 1980 103 1981 107
rect 1974 102 1981 103
rect 2014 107 2020 108
rect 2014 103 2015 107
rect 2019 106 2020 107
rect 2055 107 2061 108
rect 2055 106 2056 107
rect 2019 104 2056 106
rect 2019 103 2020 104
rect 2014 102 2020 103
rect 2055 103 2056 104
rect 2060 103 2061 107
rect 2064 106 2066 112
rect 2118 112 2124 113
rect 2118 108 2119 112
rect 2123 108 2124 112
rect 2095 107 2101 108
rect 2118 107 2124 108
rect 2095 106 2096 107
rect 2064 104 2096 106
rect 2055 102 2061 103
rect 2095 103 2096 104
rect 2100 103 2101 107
rect 2095 102 2101 103
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 142 92 148 93
rect 142 88 143 92
rect 147 88 148 92
rect 142 87 148 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 222 92 228 93
rect 222 88 223 92
rect 227 88 228 92
rect 222 87 228 88
rect 262 92 268 93
rect 262 88 263 92
rect 267 88 268 92
rect 262 87 268 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 342 92 348 93
rect 342 88 343 92
rect 347 88 348 92
rect 342 87 348 88
rect 382 92 388 93
rect 382 88 383 92
rect 387 88 388 92
rect 382 87 388 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 502 92 508 93
rect 502 88 503 92
rect 507 88 508 92
rect 502 87 508 88
rect 542 92 548 93
rect 542 88 543 92
rect 547 88 548 92
rect 542 87 548 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 622 92 628 93
rect 622 88 623 92
rect 627 88 628 92
rect 622 87 628 88
rect 662 92 668 93
rect 662 88 663 92
rect 667 88 668 92
rect 662 87 668 88
rect 702 92 708 93
rect 702 88 703 92
rect 707 88 708 92
rect 702 87 708 88
rect 742 92 748 93
rect 742 88 743 92
rect 747 88 748 92
rect 742 87 748 88
rect 782 92 788 93
rect 782 88 783 92
rect 787 88 788 92
rect 782 87 788 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 878 92 884 93
rect 878 88 879 92
rect 883 88 884 92
rect 878 87 884 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 966 92 972 93
rect 966 88 967 92
rect 971 88 972 92
rect 966 87 972 88
rect 1006 92 1012 93
rect 1006 88 1007 92
rect 1011 88 1012 92
rect 1006 87 1012 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1134 95 1140 96
rect 1134 91 1135 95
rect 1139 91 1140 95
rect 2118 95 2124 96
rect 1134 90 1140 91
rect 1158 92 1164 93
rect 1046 87 1052 88
rect 1158 88 1159 92
rect 1163 88 1164 92
rect 1158 87 1164 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1398 92 1404 93
rect 1398 88 1399 92
rect 1403 88 1404 92
rect 1398 87 1404 88
rect 1454 92 1460 93
rect 1454 88 1455 92
rect 1459 88 1460 92
rect 1454 87 1460 88
rect 1510 92 1516 93
rect 1510 88 1511 92
rect 1515 88 1516 92
rect 1510 87 1516 88
rect 1558 92 1564 93
rect 1558 88 1559 92
rect 1563 88 1564 92
rect 1558 87 1564 88
rect 1606 92 1612 93
rect 1606 88 1607 92
rect 1611 88 1612 92
rect 1606 87 1612 88
rect 1646 92 1652 93
rect 1646 88 1647 92
rect 1651 88 1652 92
rect 1646 87 1652 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1726 92 1732 93
rect 1726 88 1727 92
rect 1731 88 1732 92
rect 1726 87 1732 88
rect 1766 92 1772 93
rect 1766 88 1767 92
rect 1771 88 1772 92
rect 1766 87 1772 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1902 92 1908 93
rect 1902 88 1903 92
rect 1907 88 1908 92
rect 1902 87 1908 88
rect 1950 92 1956 93
rect 1950 88 1951 92
rect 1955 88 1956 92
rect 1950 87 1956 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2030 92 2036 93
rect 2030 88 2031 92
rect 2035 88 2036 92
rect 2030 87 2036 88
rect 2070 92 2076 93
rect 2070 88 2071 92
rect 2075 88 2076 92
rect 2118 91 2119 95
rect 2123 91 2124 95
rect 2118 90 2124 91
rect 2070 87 2076 88
<< m3c >>
rect 1679 2219 1683 2223
rect 1715 2219 1719 2223
rect 1751 2219 1755 2223
rect 1795 2219 1799 2223
rect 111 2201 115 2205
rect 135 2204 139 2208
rect 175 2204 179 2208
rect 215 2204 219 2208
rect 255 2204 259 2208
rect 319 2204 323 2208
rect 383 2204 387 2208
rect 447 2204 451 2208
rect 511 2204 515 2208
rect 575 2204 579 2208
rect 631 2204 635 2208
rect 687 2204 691 2208
rect 735 2204 739 2208
rect 791 2204 795 2208
rect 847 2204 851 2208
rect 903 2204 907 2208
rect 1687 2208 1691 2212
rect 1727 2208 1731 2212
rect 1767 2208 1771 2212
rect 1807 2208 1811 2212
rect 1095 2201 1099 2205
rect 1135 2200 1139 2204
rect 2119 2200 2123 2204
rect 1715 2195 1716 2199
rect 1716 2195 1719 2199
rect 1751 2195 1752 2199
rect 1752 2195 1755 2199
rect 1795 2195 1796 2199
rect 1796 2195 1799 2199
rect 1815 2195 1819 2199
rect 111 2184 115 2188
rect 163 2187 164 2191
rect 164 2187 167 2191
rect 203 2187 204 2191
rect 204 2187 207 2191
rect 243 2187 244 2191
rect 244 2187 247 2191
rect 311 2187 315 2191
rect 375 2187 379 2191
rect 439 2187 443 2191
rect 455 2187 459 2191
rect 567 2187 571 2191
rect 623 2187 627 2191
rect 679 2187 683 2191
rect 727 2187 731 2191
rect 783 2187 787 2191
rect 839 2187 843 2191
rect 895 2187 899 2191
rect 911 2187 915 2191
rect 1095 2184 1099 2188
rect 1135 2183 1139 2187
rect 135 2176 139 2180
rect 175 2176 179 2180
rect 215 2176 219 2180
rect 255 2176 259 2180
rect 319 2176 323 2180
rect 383 2176 387 2180
rect 447 2176 451 2180
rect 511 2176 515 2180
rect 575 2176 579 2180
rect 631 2176 635 2180
rect 687 2176 691 2180
rect 735 2176 739 2180
rect 791 2176 795 2180
rect 847 2176 851 2180
rect 903 2176 907 2180
rect 1687 2180 1691 2184
rect 1727 2180 1731 2184
rect 1767 2180 1771 2184
rect 1807 2180 1811 2184
rect 2119 2183 2123 2187
rect 163 2163 167 2167
rect 203 2163 207 2167
rect 243 2163 247 2167
rect 311 2163 315 2167
rect 375 2163 379 2167
rect 439 2163 443 2167
rect 567 2163 571 2167
rect 623 2163 627 2167
rect 679 2163 683 2167
rect 727 2163 731 2167
rect 783 2163 787 2167
rect 839 2163 843 2167
rect 895 2163 899 2167
rect 1135 2165 1139 2169
rect 1159 2168 1163 2172
rect 1199 2168 1203 2172
rect 1239 2168 1243 2172
rect 1279 2168 1283 2172
rect 1335 2168 1339 2172
rect 1391 2168 1395 2172
rect 1455 2168 1459 2172
rect 1527 2168 1531 2172
rect 1591 2168 1595 2172
rect 1663 2168 1667 2172
rect 1735 2168 1739 2172
rect 1807 2168 1811 2172
rect 1879 2168 1883 2172
rect 2119 2165 2123 2169
rect 455 2151 459 2155
rect 911 2151 915 2155
rect 1175 2155 1179 2159
rect 1319 2159 1323 2163
rect 1767 2159 1771 2163
rect 299 2143 303 2147
rect 339 2143 343 2147
rect 231 2132 235 2136
rect 111 2124 115 2128
rect 383 2139 387 2143
rect 727 2143 731 2147
rect 1135 2148 1139 2152
rect 1187 2151 1188 2155
rect 1188 2151 1191 2155
rect 1227 2151 1228 2155
rect 1228 2151 1231 2155
rect 1267 2151 1268 2155
rect 1268 2151 1271 2155
rect 1327 2151 1331 2155
rect 1383 2151 1387 2155
rect 1447 2151 1451 2155
rect 1499 2151 1503 2155
rect 1535 2151 1539 2155
rect 1655 2151 1659 2155
rect 1679 2151 1683 2155
rect 1759 2151 1760 2155
rect 1760 2151 1763 2155
rect 1871 2151 1875 2155
rect 827 2143 831 2147
rect 2119 2148 2123 2152
rect 271 2132 275 2136
rect 311 2132 315 2136
rect 359 2132 363 2136
rect 423 2132 427 2136
rect 487 2132 491 2136
rect 559 2132 563 2136
rect 639 2132 643 2136
rect 719 2132 723 2136
rect 799 2132 803 2136
rect 879 2132 883 2136
rect 1159 2140 1163 2144
rect 1199 2140 1203 2144
rect 1239 2140 1243 2144
rect 1279 2140 1283 2144
rect 1335 2140 1339 2144
rect 1391 2140 1395 2144
rect 1455 2140 1459 2144
rect 1527 2140 1531 2144
rect 1591 2140 1595 2144
rect 1663 2140 1667 2144
rect 1735 2140 1739 2144
rect 1807 2140 1811 2144
rect 1879 2140 1883 2144
rect 967 2132 971 2136
rect 299 2119 300 2123
rect 300 2119 303 2123
rect 339 2119 340 2123
rect 340 2119 343 2123
rect 383 2119 384 2123
rect 384 2119 387 2123
rect 479 2119 483 2123
rect 827 2119 828 2123
rect 828 2119 831 2123
rect 1095 2124 1099 2128
rect 1175 2127 1179 2131
rect 1187 2127 1191 2131
rect 1227 2127 1231 2131
rect 1267 2127 1271 2131
rect 1327 2127 1331 2131
rect 1383 2127 1387 2131
rect 1447 2127 1451 2131
rect 1499 2127 1503 2131
rect 1647 2127 1651 2131
rect 1655 2127 1659 2131
rect 1767 2127 1771 2131
rect 1815 2127 1819 2131
rect 1871 2127 1875 2131
rect 1031 2119 1035 2123
rect 1179 2115 1183 2119
rect 1187 2115 1191 2119
rect 1227 2115 1231 2119
rect 1267 2115 1271 2119
rect 111 2107 115 2111
rect 231 2104 235 2108
rect 271 2104 275 2108
rect 311 2104 315 2108
rect 359 2104 363 2108
rect 423 2104 427 2108
rect 487 2104 491 2108
rect 559 2104 563 2108
rect 639 2104 643 2108
rect 719 2104 723 2108
rect 799 2104 803 2108
rect 879 2104 883 2108
rect 967 2104 971 2108
rect 1095 2107 1099 2111
rect 1159 2104 1163 2108
rect 1199 2104 1203 2108
rect 1239 2104 1243 2108
rect 1295 2104 1299 2108
rect 1367 2104 1371 2108
rect 1403 2115 1407 2119
rect 1535 2115 1539 2119
rect 1615 2115 1619 2119
rect 1627 2115 1631 2119
rect 1759 2115 1763 2119
rect 1799 2115 1803 2119
rect 1867 2115 1871 2119
rect 1983 2115 1987 2119
rect 1995 2115 1999 2119
rect 2051 2115 2055 2119
rect 1135 2096 1139 2100
rect 1439 2104 1443 2108
rect 1519 2104 1523 2108
rect 1599 2104 1603 2108
rect 1679 2104 1683 2108
rect 1751 2104 1755 2108
rect 1823 2104 1827 2108
rect 1887 2104 1891 2108
rect 1951 2104 1955 2108
rect 2023 2104 2027 2108
rect 2071 2104 2075 2108
rect 111 2085 115 2089
rect 303 2088 307 2092
rect 351 2088 355 2092
rect 407 2088 411 2092
rect 471 2088 475 2092
rect 543 2088 547 2092
rect 623 2088 627 2092
rect 703 2088 707 2092
rect 783 2088 787 2092
rect 863 2088 867 2092
rect 951 2088 955 2092
rect 1039 2088 1043 2092
rect 1187 2091 1188 2095
rect 1188 2091 1191 2095
rect 1227 2091 1228 2095
rect 1228 2091 1231 2095
rect 1267 2091 1268 2095
rect 1268 2091 1271 2095
rect 1319 2091 1320 2095
rect 1320 2091 1323 2095
rect 1403 2091 1407 2095
rect 1487 2091 1491 2095
rect 2119 2096 2123 2100
rect 1627 2091 1628 2095
rect 1628 2091 1631 2095
rect 1647 2091 1651 2095
rect 1799 2091 1803 2095
rect 1867 2091 1871 2095
rect 1903 2091 1907 2095
rect 1995 2091 1999 2095
rect 2051 2091 2052 2095
rect 2052 2091 2055 2095
rect 2059 2091 2063 2095
rect 1095 2085 1099 2089
rect 1135 2079 1139 2083
rect 1159 2076 1163 2080
rect 111 2068 115 2072
rect 287 2071 291 2075
rect 399 2071 403 2075
rect 463 2071 467 2075
rect 535 2071 539 2075
rect 615 2071 619 2075
rect 631 2071 635 2075
rect 727 2071 728 2075
rect 728 2071 731 2075
rect 823 2071 827 2075
rect 1199 2076 1203 2080
rect 1239 2076 1243 2080
rect 1295 2076 1299 2080
rect 1367 2076 1371 2080
rect 1439 2076 1443 2080
rect 1519 2076 1523 2080
rect 1599 2076 1603 2080
rect 1679 2076 1683 2080
rect 1751 2076 1755 2080
rect 1823 2076 1827 2080
rect 1887 2076 1891 2080
rect 1951 2076 1955 2080
rect 2023 2076 2027 2080
rect 2071 2076 2075 2080
rect 2119 2079 2123 2083
rect 1095 2068 1099 2072
rect 303 2060 307 2064
rect 351 2060 355 2064
rect 407 2060 411 2064
rect 471 2060 475 2064
rect 543 2060 547 2064
rect 623 2060 627 2064
rect 703 2060 707 2064
rect 783 2060 787 2064
rect 863 2060 867 2064
rect 951 2060 955 2064
rect 1039 2060 1043 2064
rect 1135 2061 1139 2065
rect 1159 2064 1163 2068
rect 1215 2064 1219 2068
rect 1303 2064 1307 2068
rect 1399 2064 1403 2068
rect 1495 2064 1499 2068
rect 1591 2064 1595 2068
rect 1679 2064 1683 2068
rect 1759 2064 1763 2068
rect 1831 2064 1835 2068
rect 1895 2064 1899 2068
rect 1959 2064 1963 2068
rect 2023 2064 2027 2068
rect 2071 2064 2075 2068
rect 2119 2061 2123 2065
rect 391 2047 395 2051
rect 399 2047 403 2051
rect 463 2047 467 2051
rect 535 2047 539 2051
rect 615 2047 619 2051
rect 775 2047 779 2051
rect 1031 2047 1035 2051
rect 1135 2044 1139 2048
rect 1179 2047 1183 2051
rect 1359 2047 1363 2051
rect 1615 2047 1616 2051
rect 1616 2047 1619 2051
rect 1647 2047 1651 2051
rect 1751 2047 1755 2051
rect 1983 2047 1984 2051
rect 1984 2047 1987 2051
rect 2063 2047 2067 2051
rect 2079 2047 2083 2051
rect 479 2039 483 2043
rect 2119 2044 2123 2048
rect 631 2039 635 2043
rect 255 2031 259 2035
rect 287 2031 291 2035
rect 399 2031 403 2035
rect 531 2031 535 2035
rect 1159 2036 1163 2040
rect 643 2031 647 2035
rect 651 2031 655 2035
rect 723 2031 727 2035
rect 823 2031 827 2035
rect 843 2031 847 2035
rect 891 2031 895 2035
rect 939 2031 943 2035
rect 987 2031 991 2035
rect 1031 2031 1035 2035
rect 1215 2036 1219 2040
rect 1303 2036 1307 2040
rect 1399 2036 1403 2040
rect 1495 2036 1499 2040
rect 1591 2036 1595 2040
rect 1679 2036 1683 2040
rect 1759 2036 1763 2040
rect 1831 2036 1835 2040
rect 1895 2036 1899 2040
rect 1959 2036 1963 2040
rect 2023 2036 2027 2040
rect 2071 2036 2075 2040
rect 183 2020 187 2024
rect 279 2020 283 2024
rect 375 2020 379 2024
rect 463 2020 467 2024
rect 543 2020 547 2024
rect 623 2020 627 2024
rect 695 2020 699 2024
rect 759 2020 763 2024
rect 815 2020 819 2024
rect 863 2020 867 2024
rect 911 2020 915 2024
rect 959 2020 963 2024
rect 1007 2020 1011 2024
rect 1047 2020 1051 2024
rect 1267 2023 1271 2027
rect 1487 2023 1491 2027
rect 1647 2023 1651 2027
rect 1671 2023 1675 2027
rect 1903 2023 1907 2027
rect 2055 2023 2059 2027
rect 2063 2023 2067 2027
rect 111 2012 115 2016
rect 1095 2012 1099 2016
rect 167 2007 171 2011
rect 255 2007 259 2011
rect 391 2007 395 2011
rect 455 2007 459 2011
rect 531 2007 535 2011
rect 651 2007 652 2011
rect 652 2007 655 2011
rect 723 2007 724 2011
rect 724 2007 727 2011
rect 775 2007 779 2011
rect 843 2007 844 2011
rect 844 2007 847 2011
rect 891 2007 892 2011
rect 892 2007 895 2011
rect 939 2007 940 2011
rect 940 2007 943 2011
rect 987 2007 988 2011
rect 988 2007 991 2011
rect 1031 2007 1032 2011
rect 1032 2007 1035 2011
rect 1187 2011 1191 2015
rect 1359 2011 1363 2015
rect 1379 2011 1383 2015
rect 1647 2011 1651 2015
rect 1751 2011 1755 2015
rect 1771 2011 1775 2015
rect 1851 2011 1855 2015
rect 1939 2011 1943 2015
rect 1987 2011 1991 2015
rect 2079 2011 2083 2015
rect 1159 2000 1163 2004
rect 111 1995 115 1999
rect 1239 2000 1243 2004
rect 1351 2000 1355 2004
rect 1455 2000 1459 2004
rect 1559 2000 1563 2004
rect 1655 2000 1659 2004
rect 1743 2000 1747 2004
rect 1823 2000 1827 2004
rect 1895 2000 1899 2004
rect 1959 2000 1963 2004
rect 2023 2000 2027 2004
rect 2071 2000 2075 2004
rect 183 1992 187 1996
rect 279 1992 283 1996
rect 375 1992 379 1996
rect 463 1992 467 1996
rect 543 1992 547 1996
rect 623 1992 627 1996
rect 695 1992 699 1996
rect 759 1992 763 1996
rect 815 1992 819 1996
rect 863 1992 867 1996
rect 911 1992 915 1996
rect 959 1992 963 1996
rect 1007 1992 1011 1996
rect 1047 1992 1051 1996
rect 1095 1995 1099 1999
rect 1135 1992 1139 1996
rect 2119 1992 2123 1996
rect 1187 1987 1188 1991
rect 1188 1987 1191 1991
rect 1267 1987 1268 1991
rect 1268 1987 1271 1991
rect 1379 1987 1380 1991
rect 1380 1987 1383 1991
rect 1567 1987 1571 1991
rect 1671 1987 1675 1991
rect 1771 1987 1772 1991
rect 1772 1987 1775 1991
rect 1851 1987 1852 1991
rect 1852 1987 1855 1991
rect 1939 1987 1943 1991
rect 1987 1987 1988 1991
rect 1988 1987 1991 1991
rect 2059 1987 2063 1991
rect 111 1977 115 1981
rect 159 1980 163 1984
rect 231 1980 235 1984
rect 303 1980 307 1984
rect 375 1980 379 1984
rect 447 1980 451 1984
rect 527 1980 531 1984
rect 607 1980 611 1984
rect 687 1980 691 1984
rect 759 1980 763 1984
rect 831 1980 835 1984
rect 911 1980 915 1984
rect 991 1980 995 1984
rect 1095 1977 1099 1981
rect 643 1971 647 1975
rect 111 1960 115 1964
rect 183 1963 184 1967
rect 184 1963 187 1967
rect 295 1963 299 1967
rect 367 1963 371 1967
rect 399 1963 400 1967
rect 400 1963 403 1967
rect 519 1963 523 1967
rect 599 1963 603 1967
rect 679 1963 683 1967
rect 711 1963 712 1967
rect 712 1963 715 1967
rect 859 1971 863 1975
rect 1135 1975 1139 1979
rect 983 1963 987 1967
rect 1159 1972 1163 1976
rect 1239 1972 1243 1976
rect 1351 1972 1355 1976
rect 1455 1972 1459 1976
rect 1559 1972 1563 1976
rect 1655 1972 1659 1976
rect 1743 1972 1747 1976
rect 1823 1972 1827 1976
rect 1895 1972 1899 1976
rect 1959 1972 1963 1976
rect 2023 1972 2027 1976
rect 2071 1972 2075 1976
rect 2119 1975 2123 1979
rect 1095 1960 1099 1964
rect 159 1952 163 1956
rect 231 1952 235 1956
rect 303 1952 307 1956
rect 375 1952 379 1956
rect 447 1952 451 1956
rect 527 1952 531 1956
rect 607 1952 611 1956
rect 687 1952 691 1956
rect 759 1952 763 1956
rect 831 1952 835 1956
rect 911 1952 915 1956
rect 991 1952 995 1956
rect 1135 1945 1139 1949
rect 1359 1948 1363 1952
rect 1423 1948 1427 1952
rect 1487 1948 1491 1952
rect 1559 1948 1563 1952
rect 1631 1948 1635 1952
rect 1703 1948 1707 1952
rect 1775 1948 1779 1952
rect 1847 1948 1851 1952
rect 1927 1948 1931 1952
rect 2007 1948 2011 1952
rect 2071 1948 2075 1952
rect 2119 1945 2123 1949
rect 167 1939 171 1943
rect 199 1931 203 1935
rect 295 1939 299 1943
rect 367 1939 371 1943
rect 455 1939 459 1943
rect 519 1939 523 1943
rect 599 1939 603 1943
rect 679 1939 683 1943
rect 859 1939 863 1943
rect 903 1939 907 1943
rect 983 1939 987 1943
rect 1383 1939 1387 1943
rect 471 1931 475 1935
rect 727 1931 731 1935
rect 183 1923 187 1927
rect 259 1923 263 1927
rect 323 1923 327 1927
rect 395 1923 399 1927
rect 1135 1928 1139 1932
rect 1415 1931 1419 1935
rect 1447 1931 1448 1935
rect 1448 1931 1451 1935
rect 1647 1931 1651 1935
rect 2063 1931 2067 1935
rect 2079 1931 2083 1935
rect 555 1923 559 1927
rect 711 1923 715 1927
rect 811 1923 815 1927
rect 819 1923 823 1927
rect 2119 1928 2123 1932
rect 1359 1920 1363 1924
rect 1423 1920 1427 1924
rect 1487 1920 1491 1924
rect 1559 1920 1563 1924
rect 1631 1920 1635 1924
rect 1703 1920 1707 1924
rect 1775 1920 1779 1924
rect 1847 1920 1851 1924
rect 1927 1920 1931 1924
rect 2007 1920 2011 1924
rect 2071 1920 2075 1924
rect 135 1912 139 1916
rect 175 1912 179 1916
rect 231 1912 235 1916
rect 295 1912 299 1916
rect 367 1912 371 1916
rect 447 1912 451 1916
rect 527 1912 531 1916
rect 615 1912 619 1916
rect 703 1912 707 1916
rect 791 1912 795 1916
rect 879 1912 883 1916
rect 111 1904 115 1908
rect 1095 1904 1099 1908
rect 163 1899 164 1903
rect 164 1899 167 1903
rect 199 1899 200 1903
rect 200 1899 203 1903
rect 259 1899 260 1903
rect 260 1899 263 1903
rect 323 1899 324 1903
rect 324 1899 327 1903
rect 395 1899 396 1903
rect 396 1899 399 1903
rect 471 1899 472 1903
rect 472 1899 475 1903
rect 555 1899 556 1903
rect 556 1899 559 1903
rect 639 1899 640 1903
rect 640 1899 643 1903
rect 727 1899 728 1903
rect 728 1899 731 1903
rect 819 1899 820 1903
rect 820 1899 823 1903
rect 903 1899 904 1903
rect 904 1899 907 1903
rect 1343 1903 1347 1907
rect 1383 1907 1387 1911
rect 1415 1907 1419 1911
rect 1475 1903 1479 1907
rect 1567 1907 1571 1911
rect 1987 1907 1991 1911
rect 2055 1907 2059 1911
rect 2063 1907 2067 1911
rect 1259 1895 1263 1899
rect 1447 1895 1451 1899
rect 1467 1895 1471 1899
rect 1567 1895 1571 1899
rect 1603 1895 1607 1899
rect 1683 1895 1687 1899
rect 111 1887 115 1891
rect 135 1884 139 1888
rect 175 1884 179 1888
rect 231 1884 235 1888
rect 295 1884 299 1888
rect 367 1884 371 1888
rect 447 1884 451 1888
rect 527 1884 531 1888
rect 615 1884 619 1888
rect 703 1884 707 1888
rect 791 1884 795 1888
rect 879 1884 883 1888
rect 1095 1887 1099 1891
rect 1775 1891 1779 1895
rect 1891 1895 1895 1899
rect 2079 1895 2083 1899
rect 1231 1884 1235 1888
rect 1271 1884 1275 1888
rect 1319 1884 1323 1888
rect 1375 1884 1379 1888
rect 1439 1884 1443 1888
rect 1503 1884 1507 1888
rect 1575 1884 1579 1888
rect 1655 1884 1659 1888
rect 1751 1884 1755 1888
rect 1863 1884 1867 1888
rect 1975 1884 1979 1888
rect 2071 1884 2075 1888
rect 1135 1876 1139 1880
rect 2119 1876 2123 1880
rect 111 1865 115 1869
rect 135 1868 139 1872
rect 175 1868 179 1872
rect 223 1868 227 1872
rect 287 1868 291 1872
rect 359 1868 363 1872
rect 431 1868 435 1872
rect 503 1868 507 1872
rect 567 1868 571 1872
rect 631 1868 635 1872
rect 695 1868 699 1872
rect 759 1868 763 1872
rect 831 1868 835 1872
rect 1259 1871 1260 1875
rect 1260 1871 1263 1875
rect 1295 1871 1296 1875
rect 1296 1871 1299 1875
rect 1343 1871 1344 1875
rect 1344 1871 1347 1875
rect 1467 1871 1468 1875
rect 1468 1871 1471 1875
rect 1475 1871 1479 1875
rect 1603 1871 1604 1875
rect 1604 1871 1607 1875
rect 1683 1871 1684 1875
rect 1684 1871 1687 1875
rect 1775 1871 1776 1875
rect 1776 1871 1779 1875
rect 1891 1871 1892 1875
rect 1892 1871 1895 1875
rect 1987 1871 1991 1875
rect 1095 1865 1099 1869
rect 311 1859 315 1863
rect 111 1848 115 1852
rect 143 1851 147 1855
rect 215 1851 219 1855
rect 231 1851 235 1855
rect 423 1851 427 1855
rect 527 1859 531 1863
rect 559 1851 563 1855
rect 595 1851 596 1855
rect 596 1851 599 1855
rect 811 1859 815 1863
rect 1135 1859 1139 1863
rect 1231 1856 1235 1860
rect 751 1851 755 1855
rect 823 1851 827 1855
rect 1271 1856 1275 1860
rect 1319 1856 1323 1860
rect 1375 1856 1379 1860
rect 1439 1856 1443 1860
rect 1503 1856 1507 1860
rect 1575 1856 1579 1860
rect 1655 1856 1659 1860
rect 1751 1856 1755 1860
rect 1863 1856 1867 1860
rect 1975 1856 1979 1860
rect 2071 1856 2075 1860
rect 2119 1859 2123 1863
rect 1095 1848 1099 1852
rect 135 1840 139 1844
rect 175 1840 179 1844
rect 223 1840 227 1844
rect 287 1840 291 1844
rect 359 1840 363 1844
rect 431 1840 435 1844
rect 503 1840 507 1844
rect 567 1840 571 1844
rect 631 1840 635 1844
rect 695 1840 699 1844
rect 759 1840 763 1844
rect 831 1840 835 1844
rect 1135 1837 1139 1841
rect 1159 1840 1163 1844
rect 1199 1840 1203 1844
rect 1239 1840 1243 1844
rect 1303 1840 1307 1844
rect 1367 1840 1371 1844
rect 1431 1840 1435 1844
rect 1503 1840 1507 1844
rect 1583 1840 1587 1844
rect 1671 1840 1675 1844
rect 1767 1840 1771 1844
rect 1871 1840 1875 1844
rect 1983 1840 1987 1844
rect 2071 1840 2075 1844
rect 2119 1837 2123 1841
rect 163 1827 167 1831
rect 215 1827 219 1831
rect 311 1827 315 1831
rect 375 1827 379 1831
rect 423 1827 427 1831
rect 527 1827 531 1831
rect 559 1827 563 1831
rect 639 1827 643 1831
rect 743 1827 747 1831
rect 751 1827 755 1831
rect 823 1827 827 1831
rect 1567 1831 1571 1835
rect 231 1819 235 1823
rect 463 1819 467 1823
rect 1015 1819 1019 1823
rect 1135 1820 1139 1824
rect 143 1811 147 1815
rect 163 1811 167 1815
rect 299 1811 303 1815
rect 511 1811 515 1815
rect 519 1811 523 1815
rect 595 1811 599 1815
rect 715 1811 719 1815
rect 867 1811 871 1815
rect 1035 1811 1039 1815
rect 1159 1812 1163 1816
rect 1199 1812 1203 1816
rect 1359 1823 1363 1827
rect 1375 1823 1379 1827
rect 1495 1823 1499 1827
rect 1575 1823 1579 1827
rect 1663 1823 1667 1827
rect 1759 1823 1763 1827
rect 1863 1823 1867 1827
rect 2063 1823 2067 1827
rect 2079 1823 2083 1827
rect 2119 1820 2123 1824
rect 1239 1812 1243 1816
rect 1303 1812 1307 1816
rect 1367 1812 1371 1816
rect 1431 1812 1435 1816
rect 1503 1812 1507 1816
rect 1583 1812 1587 1816
rect 1671 1812 1675 1816
rect 1767 1812 1771 1816
rect 1871 1812 1875 1816
rect 1983 1812 1987 1816
rect 2071 1812 2075 1816
rect 135 1800 139 1804
rect 183 1800 187 1804
rect 263 1800 267 1804
rect 351 1800 355 1804
rect 439 1800 443 1804
rect 527 1800 531 1804
rect 607 1800 611 1804
rect 687 1800 691 1804
rect 767 1800 771 1804
rect 839 1800 843 1804
rect 911 1800 915 1804
rect 991 1800 995 1804
rect 1047 1800 1051 1804
rect 1295 1799 1299 1803
rect 1359 1799 1363 1803
rect 1439 1799 1443 1803
rect 1495 1799 1499 1803
rect 1575 1799 1579 1803
rect 1663 1799 1667 1803
rect 1759 1799 1763 1803
rect 1863 1799 1867 1803
rect 2063 1799 2067 1803
rect 111 1792 115 1796
rect 1095 1792 1099 1796
rect 163 1787 164 1791
rect 164 1787 167 1791
rect 171 1787 175 1791
rect 299 1787 303 1791
rect 375 1787 376 1791
rect 376 1787 379 1791
rect 463 1787 464 1791
rect 464 1787 467 1791
rect 511 1787 515 1791
rect 715 1787 716 1791
rect 716 1787 719 1791
rect 743 1787 747 1791
rect 867 1787 868 1791
rect 868 1787 871 1791
rect 951 1787 955 1791
rect 1015 1787 1016 1791
rect 1016 1787 1019 1791
rect 1035 1787 1039 1791
rect 1375 1791 1379 1795
rect 111 1775 115 1779
rect 135 1772 139 1776
rect 183 1772 187 1776
rect 263 1772 267 1776
rect 351 1772 355 1776
rect 439 1772 443 1776
rect 527 1772 531 1776
rect 607 1772 611 1776
rect 687 1772 691 1776
rect 767 1772 771 1776
rect 839 1772 843 1776
rect 911 1772 915 1776
rect 991 1772 995 1776
rect 1047 1772 1051 1776
rect 1095 1775 1099 1779
rect 1331 1779 1335 1783
rect 1339 1779 1343 1783
rect 1379 1779 1383 1783
rect 1419 1779 1423 1783
rect 1455 1779 1459 1783
rect 1495 1779 1499 1783
rect 1539 1779 1543 1783
rect 1635 1779 1639 1783
rect 1707 1779 1711 1783
rect 1795 1779 1799 1783
rect 1899 1779 1903 1783
rect 2079 1779 2083 1783
rect 1311 1768 1315 1772
rect 1351 1768 1355 1772
rect 1391 1768 1395 1772
rect 1431 1768 1435 1772
rect 1471 1768 1475 1772
rect 1511 1768 1515 1772
rect 1551 1768 1555 1772
rect 1607 1768 1611 1772
rect 1679 1768 1683 1772
rect 1767 1768 1771 1772
rect 1871 1768 1875 1772
rect 1983 1768 1987 1772
rect 2071 1768 2075 1772
rect 1135 1760 1139 1764
rect 2119 1760 2123 1764
rect 111 1749 115 1753
rect 135 1752 139 1756
rect 199 1752 203 1756
rect 295 1752 299 1756
rect 399 1752 403 1756
rect 495 1752 499 1756
rect 591 1752 595 1756
rect 671 1752 675 1756
rect 751 1752 755 1756
rect 823 1752 827 1756
rect 887 1752 891 1756
rect 959 1752 963 1756
rect 1031 1752 1035 1756
rect 1339 1755 1340 1759
rect 1340 1755 1343 1759
rect 1379 1755 1380 1759
rect 1380 1755 1383 1759
rect 1419 1755 1420 1759
rect 1420 1755 1423 1759
rect 1455 1755 1456 1759
rect 1456 1755 1459 1759
rect 1495 1755 1496 1759
rect 1496 1755 1499 1759
rect 1539 1755 1540 1759
rect 1540 1755 1543 1759
rect 1635 1755 1636 1759
rect 1636 1755 1639 1759
rect 1707 1755 1708 1759
rect 1708 1755 1711 1759
rect 1795 1755 1796 1759
rect 1796 1755 1799 1759
rect 1899 1755 1900 1759
rect 1900 1755 1903 1759
rect 2007 1755 2008 1759
rect 2008 1755 2011 1759
rect 2091 1755 2095 1759
rect 1095 1749 1099 1753
rect 431 1743 435 1747
rect 111 1732 115 1736
rect 183 1735 187 1739
rect 287 1735 291 1739
rect 311 1735 315 1739
rect 487 1735 491 1739
rect 519 1735 520 1739
rect 520 1735 523 1739
rect 911 1743 915 1747
rect 743 1735 747 1739
rect 799 1735 803 1739
rect 1023 1735 1027 1739
rect 1135 1743 1139 1747
rect 1311 1740 1315 1744
rect 1351 1740 1355 1744
rect 1391 1740 1395 1744
rect 1431 1740 1435 1744
rect 1471 1740 1475 1744
rect 1511 1740 1515 1744
rect 1551 1740 1555 1744
rect 1607 1740 1611 1744
rect 1679 1740 1683 1744
rect 1767 1740 1771 1744
rect 1871 1740 1875 1744
rect 1983 1740 1987 1744
rect 2071 1740 2075 1744
rect 2119 1743 2123 1747
rect 1095 1732 1099 1736
rect 135 1724 139 1728
rect 199 1724 203 1728
rect 295 1724 299 1728
rect 399 1724 403 1728
rect 495 1724 499 1728
rect 591 1724 595 1728
rect 671 1724 675 1728
rect 751 1724 755 1728
rect 823 1724 827 1728
rect 887 1724 891 1728
rect 959 1724 963 1728
rect 1031 1724 1035 1728
rect 1135 1721 1139 1725
rect 1263 1724 1267 1728
rect 1319 1724 1323 1728
rect 1383 1724 1387 1728
rect 1455 1724 1459 1728
rect 1535 1724 1539 1728
rect 1615 1724 1619 1728
rect 1687 1724 1691 1728
rect 1759 1724 1763 1728
rect 1831 1724 1835 1728
rect 1895 1724 1899 1728
rect 1959 1724 1963 1728
rect 2023 1724 2027 1728
rect 2071 1724 2075 1728
rect 2119 1721 2123 1725
rect 171 1711 175 1715
rect 183 1711 187 1715
rect 287 1711 291 1715
rect 431 1711 435 1715
rect 487 1711 491 1715
rect 563 1711 567 1715
rect 311 1703 315 1707
rect 743 1711 747 1715
rect 911 1711 915 1715
rect 951 1711 955 1715
rect 1023 1711 1027 1715
rect 1135 1704 1139 1708
rect 1311 1707 1315 1711
rect 1331 1711 1335 1715
rect 1375 1707 1379 1711
rect 1447 1707 1451 1711
rect 1527 1707 1531 1711
rect 1607 1707 1611 1711
rect 1711 1715 1715 1719
rect 1743 1707 1747 1711
rect 1807 1707 1811 1711
rect 2083 1707 2087 1711
rect 2119 1704 2123 1708
rect 211 1695 215 1699
rect 323 1695 327 1699
rect 331 1695 335 1699
rect 411 1695 415 1699
rect 659 1695 663 1699
rect 791 1695 795 1699
rect 799 1695 803 1699
rect 835 1695 839 1699
rect 1263 1696 1267 1700
rect 1319 1696 1323 1700
rect 1383 1696 1387 1700
rect 1455 1696 1459 1700
rect 1535 1696 1539 1700
rect 1615 1696 1619 1700
rect 1687 1696 1691 1700
rect 1759 1696 1763 1700
rect 1831 1696 1835 1700
rect 1895 1696 1899 1700
rect 1959 1696 1963 1700
rect 2023 1696 2027 1700
rect 2071 1696 2075 1700
rect 151 1684 155 1688
rect 223 1684 227 1688
rect 303 1684 307 1688
rect 383 1684 387 1688
rect 463 1684 467 1688
rect 535 1684 539 1688
rect 607 1684 611 1688
rect 671 1684 675 1688
rect 735 1684 739 1688
rect 807 1684 811 1688
rect 879 1684 883 1688
rect 1303 1683 1307 1687
rect 1311 1683 1315 1687
rect 1375 1683 1379 1687
rect 1447 1683 1451 1687
rect 1527 1683 1531 1687
rect 1607 1683 1611 1687
rect 1711 1683 1715 1687
rect 1743 1683 1747 1687
rect 2011 1683 2015 1687
rect 2091 1683 2095 1687
rect 111 1676 115 1680
rect 167 1671 171 1675
rect 211 1671 215 1675
rect 331 1671 332 1675
rect 332 1671 335 1675
rect 411 1671 412 1675
rect 412 1671 415 1675
rect 563 1671 564 1675
rect 564 1671 567 1675
rect 655 1671 659 1675
rect 663 1671 667 1675
rect 791 1675 795 1679
rect 835 1671 836 1675
rect 836 1671 839 1675
rect 1095 1676 1099 1680
rect 1187 1671 1191 1675
rect 1195 1671 1199 1675
rect 1275 1671 1279 1675
rect 1363 1671 1367 1675
rect 1619 1667 1623 1671
rect 1627 1671 1631 1675
rect 1799 1671 1803 1675
rect 1807 1671 1811 1675
rect 111 1659 115 1663
rect 151 1656 155 1660
rect 223 1656 227 1660
rect 303 1656 307 1660
rect 383 1656 387 1660
rect 463 1656 467 1660
rect 535 1656 539 1660
rect 607 1656 611 1660
rect 671 1656 675 1660
rect 735 1656 739 1660
rect 807 1656 811 1660
rect 879 1656 883 1660
rect 1095 1659 1099 1663
rect 1167 1660 1171 1664
rect 1247 1660 1251 1664
rect 1335 1660 1339 1664
rect 1423 1660 1427 1664
rect 1511 1660 1515 1664
rect 1599 1660 1603 1664
rect 1679 1660 1683 1664
rect 1751 1660 1755 1664
rect 1815 1660 1819 1664
rect 1871 1660 1875 1664
rect 1907 1671 1911 1675
rect 1927 1660 1931 1664
rect 1983 1660 1987 1664
rect 2031 1660 2035 1664
rect 2083 1671 2087 1675
rect 2071 1660 2075 1664
rect 1135 1652 1139 1656
rect 471 1647 475 1651
rect 111 1637 115 1641
rect 175 1640 179 1644
rect 215 1640 219 1644
rect 255 1640 259 1644
rect 303 1640 307 1644
rect 359 1640 363 1644
rect 407 1640 411 1644
rect 455 1640 459 1644
rect 503 1640 507 1644
rect 551 1640 555 1644
rect 607 1640 611 1644
rect 331 1631 335 1635
rect 111 1620 115 1624
rect 203 1623 204 1627
rect 204 1623 207 1627
rect 243 1623 244 1627
rect 244 1623 247 1627
rect 279 1623 280 1627
rect 280 1623 283 1627
rect 323 1623 327 1627
rect 399 1623 403 1627
rect 535 1631 539 1635
rect 1195 1647 1196 1651
rect 1196 1647 1199 1651
rect 1275 1647 1276 1651
rect 1276 1647 1279 1651
rect 1303 1651 1307 1655
rect 1363 1647 1364 1651
rect 1364 1647 1367 1651
rect 1627 1647 1628 1651
rect 1628 1647 1631 1651
rect 1743 1647 1747 1651
rect 1775 1647 1776 1651
rect 1776 1647 1779 1651
rect 1799 1647 1803 1651
rect 1907 1647 1911 1651
rect 2011 1647 2012 1651
rect 2012 1647 2015 1651
rect 2119 1652 2123 1656
rect 663 1640 667 1644
rect 719 1640 723 1644
rect 1095 1637 1099 1641
rect 1135 1635 1139 1639
rect 495 1623 499 1627
rect 543 1623 547 1627
rect 599 1623 603 1627
rect 711 1623 715 1627
rect 1167 1632 1171 1636
rect 1247 1632 1251 1636
rect 1335 1632 1339 1636
rect 1423 1632 1427 1636
rect 1511 1632 1515 1636
rect 1599 1632 1603 1636
rect 1679 1632 1683 1636
rect 1751 1632 1755 1636
rect 1815 1632 1819 1636
rect 1871 1632 1875 1636
rect 1927 1632 1931 1636
rect 1983 1632 1987 1636
rect 2031 1632 2035 1636
rect 2071 1632 2075 1636
rect 2119 1635 2123 1639
rect 1095 1620 1099 1624
rect 1179 1623 1183 1627
rect 1471 1623 1475 1627
rect 1619 1623 1623 1627
rect 1775 1623 1779 1627
rect 175 1612 179 1616
rect 215 1612 219 1616
rect 255 1612 259 1616
rect 303 1612 307 1616
rect 359 1612 363 1616
rect 407 1612 411 1616
rect 455 1612 459 1616
rect 503 1612 507 1616
rect 551 1612 555 1616
rect 607 1612 611 1616
rect 663 1612 667 1616
rect 719 1612 723 1616
rect 1135 1613 1139 1617
rect 1159 1616 1163 1620
rect 1199 1616 1203 1620
rect 1247 1616 1251 1620
rect 1319 1616 1323 1620
rect 1391 1616 1395 1620
rect 1463 1616 1467 1620
rect 1535 1616 1539 1620
rect 1607 1616 1611 1620
rect 1679 1616 1683 1620
rect 1751 1616 1755 1620
rect 1831 1616 1835 1620
rect 2119 1613 2123 1617
rect 1187 1607 1191 1611
rect 167 1599 171 1603
rect 203 1599 207 1603
rect 243 1599 247 1603
rect 331 1599 335 1603
rect 375 1599 379 1603
rect 399 1599 403 1603
rect 471 1599 475 1603
rect 495 1599 499 1603
rect 543 1599 547 1603
rect 599 1599 603 1603
rect 655 1599 659 1603
rect 711 1599 715 1603
rect 1135 1596 1139 1600
rect 1187 1599 1188 1603
rect 1188 1599 1191 1603
rect 1311 1599 1315 1603
rect 1559 1607 1563 1611
rect 1455 1599 1459 1603
rect 1471 1599 1475 1603
rect 1599 1599 1603 1603
rect 1631 1599 1632 1603
rect 1632 1599 1635 1603
rect 1703 1607 1707 1611
rect 1823 1599 1827 1603
rect 2119 1596 2123 1600
rect 559 1587 563 1591
rect 1159 1588 1163 1592
rect 1199 1588 1203 1592
rect 1247 1588 1251 1592
rect 1319 1588 1323 1592
rect 1391 1588 1395 1592
rect 1463 1588 1467 1592
rect 1535 1588 1539 1592
rect 1607 1588 1611 1592
rect 1679 1588 1683 1592
rect 1751 1588 1755 1592
rect 1831 1588 1835 1592
rect 143 1568 147 1572
rect 271 1579 275 1583
rect 279 1579 283 1583
rect 467 1579 471 1583
rect 535 1579 539 1583
rect 571 1579 575 1583
rect 635 1579 639 1583
rect 691 1579 695 1583
rect 755 1579 759 1583
rect 819 1579 823 1583
rect 1179 1575 1183 1579
rect 1187 1575 1191 1579
rect 1311 1575 1315 1579
rect 1355 1575 1359 1579
rect 1455 1575 1459 1579
rect 1559 1575 1563 1579
rect 1599 1575 1603 1579
rect 1703 1575 1707 1579
rect 1743 1575 1747 1579
rect 1823 1575 1827 1579
rect 183 1568 187 1572
rect 231 1568 235 1572
rect 287 1568 291 1572
rect 351 1568 355 1572
rect 415 1568 419 1572
rect 479 1568 483 1572
rect 543 1568 547 1572
rect 607 1568 611 1572
rect 663 1568 667 1572
rect 727 1568 731 1572
rect 791 1568 795 1572
rect 855 1568 859 1572
rect 111 1560 115 1564
rect 151 1555 155 1559
rect 1095 1560 1099 1564
rect 1259 1563 1263 1567
rect 1267 1563 1271 1567
rect 1307 1563 1311 1567
rect 1411 1563 1415 1567
rect 1431 1563 1435 1567
rect 1499 1563 1503 1567
rect 1555 1567 1559 1571
rect 1631 1563 1635 1567
rect 1651 1563 1655 1567
rect 1707 1563 1711 1567
rect 271 1555 275 1559
rect 375 1555 376 1559
rect 376 1555 379 1559
rect 467 1555 471 1559
rect 571 1555 572 1559
rect 572 1555 575 1559
rect 635 1555 636 1559
rect 636 1555 639 1559
rect 691 1555 692 1559
rect 692 1555 695 1559
rect 755 1555 756 1559
rect 756 1555 759 1559
rect 819 1555 820 1559
rect 820 1555 823 1559
rect 839 1555 843 1559
rect 1239 1552 1243 1556
rect 1279 1552 1283 1556
rect 1327 1552 1331 1556
rect 1375 1552 1379 1556
rect 1423 1552 1427 1556
rect 1471 1552 1475 1556
rect 1519 1552 1523 1556
rect 1567 1552 1571 1556
rect 1623 1552 1627 1556
rect 1679 1552 1683 1556
rect 1735 1552 1739 1556
rect 111 1543 115 1547
rect 143 1540 147 1544
rect 183 1540 187 1544
rect 231 1540 235 1544
rect 287 1540 291 1544
rect 351 1540 355 1544
rect 415 1540 419 1544
rect 479 1540 483 1544
rect 543 1540 547 1544
rect 607 1540 611 1544
rect 663 1540 667 1544
rect 727 1540 731 1544
rect 791 1540 795 1544
rect 855 1540 859 1544
rect 1095 1543 1099 1547
rect 1135 1544 1139 1548
rect 1267 1539 1268 1543
rect 1268 1539 1271 1543
rect 1307 1539 1308 1543
rect 1308 1539 1311 1543
rect 1355 1539 1356 1543
rect 1356 1539 1359 1543
rect 1399 1539 1400 1543
rect 1400 1539 1403 1543
rect 1411 1539 1415 1543
rect 1499 1539 1500 1543
rect 1500 1539 1503 1543
rect 1547 1539 1548 1543
rect 1548 1539 1551 1543
rect 1555 1539 1559 1543
rect 1651 1539 1652 1543
rect 1652 1539 1655 1543
rect 1707 1539 1708 1543
rect 1708 1539 1711 1543
rect 2119 1544 2123 1548
rect 1135 1527 1139 1531
rect 111 1517 115 1521
rect 135 1520 139 1524
rect 175 1520 179 1524
rect 215 1520 219 1524
rect 255 1520 259 1524
rect 295 1520 299 1524
rect 335 1520 339 1524
rect 375 1520 379 1524
rect 415 1520 419 1524
rect 455 1520 459 1524
rect 495 1520 499 1524
rect 535 1520 539 1524
rect 575 1520 579 1524
rect 615 1520 619 1524
rect 655 1520 659 1524
rect 695 1520 699 1524
rect 735 1520 739 1524
rect 775 1520 779 1524
rect 831 1520 835 1524
rect 887 1520 891 1524
rect 1239 1524 1243 1528
rect 1279 1524 1283 1528
rect 1327 1524 1331 1528
rect 1375 1524 1379 1528
rect 1423 1524 1427 1528
rect 1471 1524 1475 1528
rect 1519 1524 1523 1528
rect 1567 1524 1571 1528
rect 1623 1524 1627 1528
rect 1679 1524 1683 1528
rect 1735 1524 1739 1528
rect 2119 1527 2123 1531
rect 1095 1517 1099 1521
rect 111 1500 115 1504
rect 163 1503 164 1507
rect 164 1503 167 1507
rect 203 1503 204 1507
rect 204 1503 207 1507
rect 243 1503 244 1507
rect 244 1503 247 1507
rect 283 1503 284 1507
rect 284 1503 287 1507
rect 323 1503 324 1507
rect 324 1503 327 1507
rect 363 1503 364 1507
rect 364 1503 367 1507
rect 403 1503 404 1507
rect 404 1503 407 1507
rect 443 1503 444 1507
rect 444 1503 447 1507
rect 483 1503 484 1507
rect 484 1503 487 1507
rect 523 1503 524 1507
rect 524 1503 527 1507
rect 559 1503 560 1507
rect 560 1503 563 1507
rect 603 1503 604 1507
rect 604 1503 607 1507
rect 643 1503 644 1507
rect 644 1503 647 1507
rect 683 1503 684 1507
rect 684 1503 687 1507
rect 723 1503 724 1507
rect 724 1503 727 1507
rect 763 1503 764 1507
rect 764 1503 767 1507
rect 783 1503 787 1507
rect 879 1503 883 1507
rect 927 1503 931 1507
rect 1135 1505 1139 1509
rect 1319 1508 1323 1512
rect 1359 1508 1363 1512
rect 1399 1508 1403 1512
rect 1439 1508 1443 1512
rect 1479 1508 1483 1512
rect 1519 1508 1523 1512
rect 1559 1508 1563 1512
rect 1607 1508 1611 1512
rect 1663 1508 1667 1512
rect 1735 1508 1739 1512
rect 1815 1508 1819 1512
rect 1903 1508 1907 1512
rect 1991 1508 1995 1512
rect 2071 1508 2075 1512
rect 2119 1505 2123 1509
rect 1095 1500 1099 1504
rect 1431 1499 1435 1503
rect 135 1492 139 1496
rect 175 1492 179 1496
rect 215 1492 219 1496
rect 255 1492 259 1496
rect 295 1492 299 1496
rect 335 1492 339 1496
rect 375 1492 379 1496
rect 415 1492 419 1496
rect 455 1492 459 1496
rect 495 1492 499 1496
rect 535 1492 539 1496
rect 575 1492 579 1496
rect 615 1492 619 1496
rect 655 1492 659 1496
rect 695 1492 699 1496
rect 735 1492 739 1496
rect 775 1492 779 1496
rect 831 1492 835 1496
rect 887 1492 891 1496
rect 1135 1488 1139 1492
rect 1347 1491 1348 1495
rect 1348 1491 1351 1495
rect 1383 1491 1384 1495
rect 1384 1491 1387 1495
rect 1427 1491 1428 1495
rect 1428 1491 1431 1495
rect 1467 1491 1468 1495
rect 1468 1491 1471 1495
rect 1507 1491 1508 1495
rect 1508 1491 1511 1495
rect 1599 1491 1603 1495
rect 1655 1491 1659 1495
rect 1727 1491 1731 1495
rect 1911 1491 1915 1495
rect 2063 1491 2067 1495
rect 2079 1491 2083 1495
rect 2119 1488 2123 1492
rect 151 1479 155 1483
rect 163 1479 167 1483
rect 203 1479 207 1483
rect 243 1479 247 1483
rect 283 1479 287 1483
rect 323 1479 327 1483
rect 363 1479 367 1483
rect 403 1479 407 1483
rect 443 1479 447 1483
rect 483 1479 487 1483
rect 523 1479 527 1483
rect 547 1479 551 1483
rect 603 1479 607 1483
rect 643 1479 647 1483
rect 683 1479 687 1483
rect 723 1479 727 1483
rect 763 1479 767 1483
rect 839 1479 843 1483
rect 879 1479 883 1483
rect 1319 1480 1323 1484
rect 1359 1480 1363 1484
rect 1399 1480 1403 1484
rect 1439 1480 1443 1484
rect 1479 1480 1483 1484
rect 1519 1480 1523 1484
rect 1559 1480 1563 1484
rect 1607 1480 1611 1484
rect 1663 1480 1667 1484
rect 1735 1480 1739 1484
rect 1815 1480 1819 1484
rect 1903 1480 1907 1484
rect 1991 1480 1995 1484
rect 2071 1480 2075 1484
rect 583 1467 587 1471
rect 783 1467 787 1471
rect 1327 1467 1331 1471
rect 1347 1467 1351 1471
rect 1383 1467 1387 1471
rect 1427 1467 1431 1471
rect 1467 1467 1471 1471
rect 1507 1467 1511 1471
rect 1547 1467 1551 1471
rect 1599 1467 1603 1471
rect 1655 1467 1659 1471
rect 1727 1467 1731 1471
rect 2039 1467 2043 1471
rect 2063 1467 2067 1471
rect 519 1448 523 1452
rect 559 1448 563 1452
rect 655 1455 659 1459
rect 675 1459 679 1463
rect 787 1459 791 1463
rect 919 1459 923 1463
rect 927 1459 931 1463
rect 1251 1455 1255 1459
rect 1259 1455 1263 1459
rect 1307 1455 1311 1459
rect 599 1448 603 1452
rect 647 1448 651 1452
rect 695 1448 699 1452
rect 751 1448 755 1452
rect 807 1448 811 1452
rect 871 1448 875 1452
rect 935 1448 939 1452
rect 1363 1451 1367 1455
rect 1419 1455 1423 1459
rect 1487 1455 1491 1459
rect 1591 1455 1595 1459
rect 1615 1455 1619 1459
rect 1675 1455 1679 1459
rect 1747 1455 1751 1459
rect 1835 1455 1839 1459
rect 1923 1455 1927 1459
rect 2079 1455 2083 1459
rect 111 1440 115 1444
rect 547 1435 548 1439
rect 548 1435 551 1439
rect 583 1435 584 1439
rect 584 1435 587 1439
rect 675 1435 676 1439
rect 676 1435 679 1439
rect 787 1439 791 1443
rect 1095 1440 1099 1444
rect 1231 1444 1235 1448
rect 1279 1444 1283 1448
rect 1335 1444 1339 1448
rect 1391 1444 1395 1448
rect 1455 1444 1459 1448
rect 1519 1444 1523 1448
rect 1583 1444 1587 1448
rect 1647 1444 1651 1448
rect 1719 1444 1723 1448
rect 1807 1444 1811 1448
rect 1895 1444 1899 1448
rect 1991 1444 1995 1448
rect 2071 1444 2075 1448
rect 831 1435 832 1439
rect 832 1435 835 1439
rect 887 1435 891 1439
rect 919 1435 923 1439
rect 1135 1436 1139 1440
rect 2119 1436 2123 1440
rect 1259 1431 1260 1435
rect 1260 1431 1263 1435
rect 1307 1431 1308 1435
rect 1308 1431 1311 1435
rect 1363 1431 1364 1435
rect 1364 1431 1367 1435
rect 1419 1431 1420 1435
rect 1420 1431 1423 1435
rect 1483 1431 1484 1435
rect 1484 1431 1487 1435
rect 1543 1431 1544 1435
rect 1544 1431 1547 1435
rect 1611 1431 1612 1435
rect 1612 1431 1615 1435
rect 1675 1431 1676 1435
rect 1676 1431 1679 1435
rect 1747 1431 1748 1435
rect 1748 1431 1751 1435
rect 1835 1431 1836 1435
rect 1836 1431 1839 1435
rect 1923 1431 1924 1435
rect 1924 1431 1927 1435
rect 1931 1431 1935 1435
rect 2091 1431 2095 1435
rect 111 1423 115 1427
rect 519 1420 523 1424
rect 559 1420 563 1424
rect 599 1420 603 1424
rect 647 1420 651 1424
rect 695 1420 699 1424
rect 751 1420 755 1424
rect 807 1420 811 1424
rect 871 1420 875 1424
rect 935 1420 939 1424
rect 1095 1423 1099 1427
rect 1135 1419 1139 1423
rect 1231 1416 1235 1420
rect 1279 1416 1283 1420
rect 1335 1416 1339 1420
rect 1391 1416 1395 1420
rect 1455 1416 1459 1420
rect 1519 1416 1523 1420
rect 1583 1416 1587 1420
rect 1647 1416 1651 1420
rect 1719 1416 1723 1420
rect 1807 1416 1811 1420
rect 1895 1416 1899 1420
rect 1991 1416 1995 1420
rect 2071 1416 2075 1420
rect 2119 1419 2123 1423
rect 111 1401 115 1405
rect 431 1404 435 1408
rect 471 1404 475 1408
rect 519 1404 523 1408
rect 575 1404 579 1408
rect 631 1404 635 1408
rect 695 1404 699 1408
rect 759 1404 763 1408
rect 823 1404 827 1408
rect 895 1404 899 1408
rect 967 1404 971 1408
rect 1095 1401 1099 1405
rect 1135 1397 1139 1401
rect 1159 1400 1163 1404
rect 1199 1400 1203 1404
rect 1263 1400 1267 1404
rect 1351 1400 1355 1404
rect 1447 1400 1451 1404
rect 1543 1400 1547 1404
rect 1631 1400 1635 1404
rect 1719 1400 1723 1404
rect 1799 1400 1803 1404
rect 1871 1400 1875 1404
rect 1943 1400 1947 1404
rect 2015 1400 2019 1404
rect 2071 1400 2075 1404
rect 2119 1397 2123 1401
rect 111 1384 115 1388
rect 459 1387 460 1391
rect 460 1387 463 1391
rect 511 1387 515 1391
rect 567 1387 571 1391
rect 623 1387 627 1391
rect 655 1387 656 1391
rect 656 1387 659 1391
rect 703 1387 707 1391
rect 959 1387 963 1391
rect 991 1387 992 1391
rect 992 1387 995 1391
rect 1251 1391 1255 1395
rect 1095 1384 1099 1388
rect 431 1376 435 1380
rect 471 1376 475 1380
rect 519 1376 523 1380
rect 575 1376 579 1380
rect 631 1376 635 1380
rect 695 1376 699 1380
rect 759 1376 763 1380
rect 823 1376 827 1380
rect 895 1376 899 1380
rect 967 1376 971 1380
rect 1135 1380 1139 1384
rect 1187 1383 1188 1387
rect 1188 1383 1191 1387
rect 1255 1383 1259 1387
rect 1343 1383 1347 1387
rect 1439 1383 1443 1387
rect 1535 1383 1539 1387
rect 1711 1383 1715 1387
rect 1791 1383 1795 1387
rect 1863 1383 1867 1387
rect 1887 1383 1891 1387
rect 2007 1383 2011 1387
rect 2039 1383 2040 1387
rect 2040 1383 2043 1387
rect 2083 1383 2087 1387
rect 2119 1380 2123 1384
rect 1159 1372 1163 1376
rect 1199 1372 1203 1376
rect 1263 1372 1267 1376
rect 1351 1372 1355 1376
rect 1447 1372 1451 1376
rect 1543 1372 1547 1376
rect 1631 1372 1635 1376
rect 1719 1372 1723 1376
rect 1799 1372 1803 1376
rect 1871 1372 1875 1376
rect 1943 1372 1947 1376
rect 2015 1372 2019 1376
rect 2071 1372 2075 1376
rect 443 1363 447 1367
rect 459 1363 463 1367
rect 511 1363 515 1367
rect 567 1363 571 1367
rect 623 1363 627 1367
rect 831 1363 835 1367
rect 887 1363 891 1367
rect 959 1363 963 1367
rect 1187 1359 1191 1363
rect 1255 1359 1259 1363
rect 1343 1359 1347 1363
rect 1439 1359 1443 1363
rect 1535 1359 1539 1363
rect 1671 1359 1675 1363
rect 1711 1359 1715 1363
rect 1791 1359 1795 1363
rect 1863 1359 1867 1363
rect 1879 1359 1883 1363
rect 2007 1359 2011 1363
rect 2091 1359 2095 1363
rect 383 1351 387 1355
rect 403 1351 407 1355
rect 451 1351 455 1355
rect 507 1351 511 1355
rect 587 1351 591 1355
rect 703 1351 707 1355
rect 759 1347 763 1351
rect 835 1351 839 1355
rect 983 1351 987 1355
rect 991 1351 995 1355
rect 1071 1351 1075 1355
rect 1511 1351 1515 1355
rect 1887 1351 1891 1355
rect 1991 1351 1995 1355
rect 375 1340 379 1344
rect 423 1340 427 1344
rect 479 1340 483 1344
rect 543 1340 547 1344
rect 607 1340 611 1344
rect 671 1340 675 1344
rect 735 1340 739 1344
rect 799 1340 803 1344
rect 863 1340 867 1344
rect 927 1340 931 1344
rect 999 1340 1003 1344
rect 1047 1340 1051 1344
rect 111 1332 115 1336
rect 443 1335 447 1339
rect 403 1327 404 1331
rect 404 1327 407 1331
rect 451 1327 452 1331
rect 452 1327 455 1331
rect 507 1327 508 1331
rect 508 1327 511 1331
rect 587 1327 591 1331
rect 759 1327 760 1331
rect 760 1327 763 1331
rect 835 1327 839 1331
rect 843 1327 847 1331
rect 975 1327 979 1331
rect 983 1327 987 1331
rect 1187 1343 1191 1347
rect 1283 1343 1287 1347
rect 1403 1343 1407 1347
rect 1619 1343 1623 1347
rect 1707 1343 1711 1347
rect 1787 1343 1791 1347
rect 2047 1343 2051 1347
rect 2083 1343 2087 1347
rect 1095 1332 1099 1336
rect 1159 1332 1163 1336
rect 1255 1332 1259 1336
rect 1375 1332 1379 1336
rect 1487 1332 1491 1336
rect 1591 1332 1595 1336
rect 1679 1332 1683 1336
rect 1759 1332 1763 1336
rect 1831 1332 1835 1336
rect 1903 1332 1907 1336
rect 1967 1332 1971 1336
rect 2031 1332 2035 1336
rect 2071 1332 2075 1336
rect 1135 1324 1139 1328
rect 2119 1324 2123 1328
rect 111 1315 115 1319
rect 375 1312 379 1316
rect 423 1312 427 1316
rect 479 1312 483 1316
rect 543 1312 547 1316
rect 607 1312 611 1316
rect 671 1312 675 1316
rect 735 1312 739 1316
rect 799 1312 803 1316
rect 863 1312 867 1316
rect 927 1312 931 1316
rect 999 1312 1003 1316
rect 1047 1312 1051 1316
rect 1095 1315 1099 1319
rect 1187 1319 1188 1323
rect 1188 1319 1191 1323
rect 1283 1319 1284 1323
rect 1284 1319 1287 1323
rect 1403 1319 1404 1323
rect 1404 1319 1407 1323
rect 1511 1319 1512 1323
rect 1512 1319 1515 1323
rect 1619 1319 1620 1323
rect 1620 1319 1623 1323
rect 1707 1319 1708 1323
rect 1708 1319 1711 1323
rect 1787 1319 1788 1323
rect 1788 1319 1791 1323
rect 1879 1319 1883 1323
rect 1959 1319 1963 1323
rect 1991 1319 1992 1323
rect 1992 1319 1995 1323
rect 2083 1319 2087 1323
rect 1135 1307 1139 1311
rect 111 1297 115 1301
rect 335 1300 339 1304
rect 391 1300 395 1304
rect 455 1300 459 1304
rect 527 1300 531 1304
rect 599 1300 603 1304
rect 671 1300 675 1304
rect 743 1300 747 1304
rect 823 1300 827 1304
rect 903 1300 907 1304
rect 983 1300 987 1304
rect 1047 1300 1051 1304
rect 1159 1304 1163 1308
rect 1255 1304 1259 1308
rect 1375 1304 1379 1308
rect 1487 1304 1491 1308
rect 1591 1304 1595 1308
rect 1679 1304 1683 1308
rect 1759 1304 1763 1308
rect 1831 1304 1835 1308
rect 1903 1304 1907 1308
rect 1967 1304 1971 1308
rect 2031 1304 2035 1308
rect 2071 1304 2075 1308
rect 2119 1307 2123 1311
rect 1095 1297 1099 1301
rect 383 1291 387 1295
rect 111 1280 115 1284
rect 383 1283 387 1287
rect 447 1283 451 1287
rect 519 1283 523 1287
rect 591 1283 595 1287
rect 735 1283 739 1287
rect 791 1283 795 1287
rect 919 1283 923 1287
rect 1071 1283 1072 1287
rect 1072 1283 1075 1287
rect 1135 1285 1139 1289
rect 1159 1288 1163 1292
rect 1199 1288 1203 1292
rect 1247 1288 1251 1292
rect 1319 1288 1323 1292
rect 1399 1288 1403 1292
rect 1479 1288 1483 1292
rect 1559 1288 1563 1292
rect 1639 1288 1643 1292
rect 1719 1288 1723 1292
rect 1799 1288 1803 1292
rect 1879 1288 1883 1292
rect 1967 1288 1971 1292
rect 2055 1288 2059 1292
rect 2119 1285 2123 1289
rect 1095 1280 1099 1284
rect 1271 1279 1275 1283
rect 335 1272 339 1276
rect 391 1272 395 1276
rect 455 1272 459 1276
rect 527 1272 531 1276
rect 599 1272 603 1276
rect 671 1272 675 1276
rect 743 1272 747 1276
rect 823 1272 827 1276
rect 903 1272 907 1276
rect 983 1272 987 1276
rect 1047 1272 1051 1276
rect 1135 1268 1139 1272
rect 383 1259 387 1263
rect 447 1259 451 1263
rect 519 1259 523 1263
rect 591 1259 595 1263
rect 567 1251 571 1255
rect 735 1259 739 1263
rect 843 1259 847 1263
rect 975 1259 979 1263
rect 1159 1260 1163 1264
rect 1391 1271 1395 1275
rect 1471 1271 1475 1275
rect 1631 1271 1635 1275
rect 1711 1271 1715 1275
rect 1815 1271 1819 1275
rect 1823 1271 1824 1275
rect 1824 1271 1827 1275
rect 1835 1271 1839 1275
rect 2047 1271 2051 1275
rect 2119 1268 2123 1272
rect 1199 1260 1203 1264
rect 1247 1260 1251 1264
rect 1319 1260 1323 1264
rect 1399 1260 1403 1264
rect 1479 1260 1483 1264
rect 1559 1260 1563 1264
rect 1639 1260 1643 1264
rect 1719 1260 1723 1264
rect 1799 1260 1803 1264
rect 1879 1260 1883 1264
rect 1967 1260 1971 1264
rect 2055 1260 2059 1264
rect 1271 1255 1275 1259
rect 271 1243 275 1247
rect 291 1243 295 1247
rect 443 1243 447 1247
rect 519 1243 523 1247
rect 723 1243 727 1247
rect 783 1243 787 1247
rect 791 1243 795 1247
rect 911 1243 915 1247
rect 919 1243 923 1247
rect 1267 1247 1271 1251
rect 1391 1247 1395 1251
rect 1471 1247 1475 1251
rect 1631 1247 1635 1251
rect 1711 1247 1715 1251
rect 1835 1247 1839 1251
rect 1959 1247 1963 1251
rect 2035 1247 2039 1251
rect 263 1232 267 1236
rect 311 1232 315 1236
rect 111 1224 115 1228
rect 1303 1239 1307 1243
rect 1447 1239 1451 1243
rect 1547 1239 1551 1243
rect 1823 1239 1827 1243
rect 359 1232 363 1236
rect 415 1232 419 1236
rect 479 1232 483 1236
rect 543 1232 547 1236
rect 607 1232 611 1236
rect 671 1232 675 1236
rect 735 1232 739 1236
rect 799 1232 803 1236
rect 863 1232 867 1236
rect 927 1232 931 1236
rect 1187 1231 1191 1235
rect 1227 1231 1231 1235
rect 1391 1231 1395 1235
rect 1499 1231 1503 1235
rect 1571 1231 1575 1235
rect 1815 1231 1819 1235
rect 1867 1231 1871 1235
rect 2083 1231 2087 1235
rect 291 1219 292 1223
rect 292 1219 295 1223
rect 1095 1224 1099 1228
rect 443 1219 444 1223
rect 444 1219 447 1223
rect 519 1219 523 1223
rect 567 1219 568 1223
rect 568 1219 571 1223
rect 579 1219 583 1223
rect 723 1219 727 1223
rect 783 1219 787 1223
rect 887 1219 888 1223
rect 888 1219 891 1223
rect 911 1219 915 1223
rect 1159 1220 1163 1224
rect 1199 1220 1203 1224
rect 1239 1220 1243 1224
rect 1279 1220 1283 1224
rect 1327 1220 1331 1224
rect 1375 1220 1379 1224
rect 1423 1220 1427 1224
rect 1471 1220 1475 1224
rect 1535 1220 1539 1224
rect 1615 1220 1619 1224
rect 1719 1220 1723 1224
rect 1839 1220 1843 1224
rect 1967 1220 1971 1224
rect 2071 1220 2075 1224
rect 1135 1212 1139 1216
rect 111 1207 115 1211
rect 263 1204 267 1208
rect 311 1204 315 1208
rect 359 1204 363 1208
rect 415 1204 419 1208
rect 479 1204 483 1208
rect 543 1204 547 1208
rect 607 1204 611 1208
rect 671 1204 675 1208
rect 735 1204 739 1208
rect 799 1204 803 1208
rect 863 1204 867 1208
rect 927 1204 931 1208
rect 1095 1207 1099 1211
rect 1187 1207 1188 1211
rect 1188 1207 1191 1211
rect 1227 1207 1228 1211
rect 1228 1207 1231 1211
rect 1267 1207 1268 1211
rect 1268 1207 1271 1211
rect 1303 1207 1304 1211
rect 1304 1207 1307 1211
rect 1447 1207 1448 1211
rect 1448 1207 1451 1211
rect 1499 1207 1500 1211
rect 1500 1207 1503 1211
rect 1571 1207 1575 1211
rect 2119 1212 2123 1216
rect 1867 1207 1868 1211
rect 1868 1207 1871 1211
rect 1991 1207 1992 1211
rect 1992 1207 1995 1211
rect 2087 1207 2091 1211
rect 111 1189 115 1193
rect 223 1192 227 1196
rect 279 1192 283 1196
rect 343 1192 347 1196
rect 407 1192 411 1196
rect 479 1192 483 1196
rect 551 1192 555 1196
rect 631 1192 635 1196
rect 711 1192 715 1196
rect 791 1192 795 1196
rect 871 1192 875 1196
rect 959 1192 963 1196
rect 1135 1195 1139 1199
rect 1095 1189 1099 1193
rect 1159 1192 1163 1196
rect 1199 1192 1203 1196
rect 1239 1192 1243 1196
rect 1279 1192 1283 1196
rect 1327 1192 1331 1196
rect 1375 1192 1379 1196
rect 1423 1192 1427 1196
rect 1471 1192 1475 1196
rect 1535 1192 1539 1196
rect 1615 1192 1619 1196
rect 1719 1192 1723 1196
rect 271 1183 275 1187
rect 1623 1187 1627 1191
rect 1839 1192 1843 1196
rect 1967 1192 1971 1196
rect 2071 1192 2075 1196
rect 2119 1195 2123 1199
rect 111 1172 115 1176
rect 271 1175 275 1179
rect 335 1175 339 1179
rect 399 1175 403 1179
rect 471 1175 475 1179
rect 623 1175 627 1179
rect 703 1175 707 1179
rect 783 1175 787 1179
rect 799 1175 803 1179
rect 951 1175 955 1179
rect 983 1175 984 1179
rect 984 1175 987 1179
rect 1135 1177 1139 1181
rect 1287 1180 1291 1184
rect 1327 1180 1331 1184
rect 1367 1180 1371 1184
rect 1415 1180 1419 1184
rect 1471 1180 1475 1184
rect 1527 1180 1531 1184
rect 1583 1180 1587 1184
rect 1639 1180 1643 1184
rect 1703 1180 1707 1184
rect 1767 1180 1771 1184
rect 1839 1180 1843 1184
rect 1919 1180 1923 1184
rect 2007 1180 2011 1184
rect 2071 1180 2075 1184
rect 2119 1177 2123 1181
rect 1095 1172 1099 1176
rect 1439 1171 1443 1175
rect 223 1164 227 1168
rect 279 1164 283 1168
rect 343 1164 347 1168
rect 407 1164 411 1168
rect 479 1164 483 1168
rect 551 1164 555 1168
rect 631 1164 635 1168
rect 711 1164 715 1168
rect 791 1164 795 1168
rect 871 1164 875 1168
rect 959 1164 963 1168
rect 1135 1160 1139 1164
rect 1315 1163 1316 1167
rect 1316 1163 1319 1167
rect 1355 1163 1356 1167
rect 1356 1163 1359 1167
rect 1391 1163 1392 1167
rect 1392 1163 1395 1167
rect 1519 1163 1523 1167
rect 1555 1171 1559 1175
rect 1991 1171 1995 1175
rect 1631 1163 1635 1167
rect 1695 1163 1699 1167
rect 1759 1163 1763 1167
rect 1831 1163 1835 1167
rect 1911 1163 1915 1167
rect 1935 1163 1939 1167
rect 2035 1163 2036 1167
rect 2036 1163 2039 1167
rect 2079 1163 2083 1167
rect 2119 1160 2123 1164
rect 263 1151 267 1155
rect 271 1151 275 1155
rect 335 1151 339 1155
rect 399 1151 403 1155
rect 471 1151 475 1155
rect 579 1151 583 1155
rect 623 1151 627 1155
rect 703 1151 707 1155
rect 783 1151 787 1155
rect 887 1151 891 1155
rect 951 1151 955 1155
rect 1287 1152 1291 1156
rect 1327 1152 1331 1156
rect 1367 1152 1371 1156
rect 1415 1152 1419 1156
rect 1471 1152 1475 1156
rect 1527 1152 1531 1156
rect 1583 1152 1587 1156
rect 1639 1152 1643 1156
rect 1703 1152 1707 1156
rect 1767 1152 1771 1156
rect 1839 1152 1843 1156
rect 1919 1152 1923 1156
rect 2007 1152 2011 1156
rect 2071 1152 2075 1156
rect 175 1139 179 1143
rect 183 1139 187 1143
rect 231 1139 235 1143
rect 287 1139 291 1143
rect 395 1139 399 1143
rect 579 1139 583 1143
rect 667 1139 671 1143
rect 763 1139 767 1143
rect 799 1139 803 1143
rect 975 1139 979 1143
rect 983 1139 987 1143
rect 1315 1139 1319 1143
rect 1355 1139 1359 1143
rect 1439 1139 1443 1143
rect 1495 1139 1499 1143
rect 1519 1139 1523 1143
rect 1623 1139 1627 1143
rect 1631 1139 1635 1143
rect 1695 1139 1699 1143
rect 1759 1139 1763 1143
rect 1831 1139 1835 1143
rect 1911 1139 1915 1143
rect 2055 1139 2059 1143
rect 2087 1139 2091 1143
rect 159 1128 163 1132
rect 199 1128 203 1132
rect 247 1128 251 1132
rect 303 1128 307 1132
rect 367 1128 371 1132
rect 439 1128 443 1132
rect 511 1128 515 1132
rect 591 1128 595 1132
rect 679 1128 683 1132
rect 775 1128 779 1132
rect 879 1128 883 1132
rect 991 1128 995 1132
rect 111 1120 115 1124
rect 263 1123 267 1127
rect 1679 1127 1683 1131
rect 1935 1127 1939 1131
rect 183 1115 184 1119
rect 184 1115 187 1119
rect 227 1115 228 1119
rect 228 1115 231 1119
rect 287 1115 291 1119
rect 395 1115 396 1119
rect 396 1115 399 1119
rect 1095 1120 1099 1124
rect 519 1115 523 1119
rect 579 1115 583 1119
rect 667 1115 671 1119
rect 763 1115 767 1119
rect 811 1115 815 1119
rect 975 1115 979 1119
rect 1399 1119 1403 1123
rect 1407 1119 1411 1123
rect 1451 1119 1455 1123
rect 1599 1119 1603 1123
rect 1619 1119 1623 1123
rect 1739 1119 1743 1123
rect 1795 1119 1799 1123
rect 1851 1119 1855 1123
rect 1899 1119 1903 1123
rect 1955 1119 1959 1123
rect 2047 1119 2051 1123
rect 2079 1119 2083 1123
rect 1383 1108 1387 1112
rect 111 1103 115 1107
rect 1423 1108 1427 1112
rect 1471 1108 1475 1112
rect 1527 1108 1531 1112
rect 1591 1108 1595 1112
rect 1655 1108 1659 1112
rect 1711 1108 1715 1112
rect 1767 1108 1771 1112
rect 1823 1108 1827 1112
rect 1871 1108 1875 1112
rect 1927 1108 1931 1112
rect 1983 1108 1987 1112
rect 2031 1108 2035 1112
rect 2071 1108 2075 1112
rect 159 1100 163 1104
rect 199 1100 203 1104
rect 247 1100 251 1104
rect 303 1100 307 1104
rect 367 1100 371 1104
rect 439 1100 443 1104
rect 511 1100 515 1104
rect 591 1100 595 1104
rect 679 1100 683 1104
rect 775 1100 779 1104
rect 879 1100 883 1104
rect 991 1100 995 1104
rect 1095 1103 1099 1107
rect 1135 1100 1139 1104
rect 2119 1100 2123 1104
rect 1407 1095 1408 1099
rect 1408 1095 1411 1099
rect 1451 1095 1452 1099
rect 1452 1095 1455 1099
rect 1495 1095 1496 1099
rect 1496 1095 1499 1099
rect 1551 1095 1552 1099
rect 1552 1095 1555 1099
rect 1619 1095 1620 1099
rect 1620 1095 1623 1099
rect 1679 1095 1680 1099
rect 1680 1095 1683 1099
rect 1739 1095 1740 1099
rect 1740 1095 1743 1099
rect 1795 1095 1796 1099
rect 1796 1095 1799 1099
rect 1851 1095 1852 1099
rect 1852 1095 1855 1099
rect 1899 1095 1900 1099
rect 1900 1095 1903 1099
rect 1955 1095 1956 1099
rect 1956 1095 1959 1099
rect 1999 1095 2003 1099
rect 2055 1095 2056 1099
rect 2056 1095 2059 1099
rect 2079 1095 2083 1099
rect 111 1077 115 1081
rect 199 1080 203 1084
rect 247 1080 251 1084
rect 303 1080 307 1084
rect 367 1080 371 1084
rect 431 1080 435 1084
rect 503 1080 507 1084
rect 575 1080 579 1084
rect 647 1080 651 1084
rect 719 1080 723 1084
rect 783 1080 787 1084
rect 839 1080 843 1084
rect 895 1080 899 1084
rect 951 1080 955 1084
rect 1007 1080 1011 1084
rect 1047 1080 1051 1084
rect 1135 1083 1139 1087
rect 1095 1077 1099 1081
rect 1383 1080 1387 1084
rect 1423 1080 1427 1084
rect 1471 1080 1475 1084
rect 1527 1080 1531 1084
rect 1591 1080 1595 1084
rect 1655 1080 1659 1084
rect 1711 1080 1715 1084
rect 1767 1080 1771 1084
rect 1823 1080 1827 1084
rect 1871 1080 1875 1084
rect 1927 1080 1931 1084
rect 1983 1080 1987 1084
rect 2031 1080 2035 1084
rect 2071 1080 2075 1084
rect 2119 1083 2123 1087
rect 111 1060 115 1064
rect 175 1063 179 1067
rect 347 1063 351 1067
rect 567 1063 571 1067
rect 639 1063 643 1067
rect 655 1063 659 1067
rect 775 1063 779 1067
rect 831 1063 835 1067
rect 911 1063 915 1067
rect 943 1063 947 1067
rect 999 1063 1003 1067
rect 1035 1063 1036 1067
rect 1036 1063 1039 1067
rect 1087 1063 1091 1067
rect 1135 1065 1139 1069
rect 1159 1068 1163 1072
rect 1247 1068 1251 1072
rect 1359 1068 1363 1072
rect 1471 1068 1475 1072
rect 1575 1068 1579 1072
rect 1671 1068 1675 1072
rect 1759 1068 1763 1072
rect 1847 1068 1851 1072
rect 1927 1068 1931 1072
rect 2007 1068 2011 1072
rect 2071 1068 2075 1072
rect 2119 1065 2123 1069
rect 1095 1060 1099 1064
rect 199 1052 203 1056
rect 247 1052 251 1056
rect 303 1052 307 1056
rect 367 1052 371 1056
rect 431 1052 435 1056
rect 503 1052 507 1056
rect 575 1052 579 1056
rect 647 1052 651 1056
rect 719 1052 723 1056
rect 783 1052 787 1056
rect 839 1052 843 1056
rect 895 1052 899 1056
rect 951 1052 955 1056
rect 1007 1052 1011 1056
rect 1047 1052 1051 1056
rect 1175 1055 1179 1059
rect 1135 1048 1139 1052
rect 1239 1051 1243 1055
rect 1351 1051 1355 1055
rect 1703 1059 1707 1063
rect 1567 1051 1571 1055
rect 1599 1051 1600 1055
rect 1600 1051 1603 1055
rect 1751 1051 1755 1055
rect 1815 1051 1819 1055
rect 2047 1051 2051 1055
rect 2119 1048 2123 1052
rect 347 1039 351 1043
rect 423 1039 427 1043
rect 519 1039 523 1043
rect 567 1039 571 1043
rect 639 1039 643 1043
rect 775 1039 779 1043
rect 831 1039 835 1043
rect 927 1039 931 1043
rect 943 1039 947 1043
rect 999 1039 1003 1043
rect 1035 1039 1039 1043
rect 1159 1040 1163 1044
rect 1247 1040 1251 1044
rect 1359 1040 1363 1044
rect 1471 1040 1475 1044
rect 1575 1040 1579 1044
rect 1671 1040 1675 1044
rect 1759 1040 1763 1044
rect 1847 1040 1851 1044
rect 1927 1040 1931 1044
rect 2007 1040 2011 1044
rect 2071 1040 2075 1044
rect 811 1031 815 1035
rect 239 1023 243 1027
rect 255 1023 259 1027
rect 379 1023 383 1027
rect 547 1023 551 1027
rect 619 1023 623 1027
rect 655 1023 659 1027
rect 711 1023 715 1027
rect 731 1023 735 1027
rect 803 1023 807 1027
rect 867 1023 871 1027
rect 911 1023 915 1027
rect 995 1023 999 1027
rect 1087 1027 1091 1031
rect 1239 1027 1243 1031
rect 1351 1027 1355 1031
rect 1487 1027 1491 1031
rect 1567 1027 1571 1031
rect 1703 1027 1707 1031
rect 1751 1027 1755 1031
rect 1999 1027 2003 1031
rect 2079 1027 2083 1031
rect 223 1012 227 1016
rect 271 1012 275 1016
rect 335 1012 339 1016
rect 407 1012 411 1016
rect 479 1012 483 1016
rect 559 1012 563 1016
rect 631 1012 635 1016
rect 703 1012 707 1016
rect 775 1012 779 1016
rect 839 1012 843 1016
rect 903 1012 907 1016
rect 967 1012 971 1016
rect 1039 1012 1043 1016
rect 1175 1015 1179 1019
rect 1187 1015 1191 1019
rect 1259 1015 1263 1019
rect 1331 1015 1335 1019
rect 1527 1015 1531 1019
rect 1535 1015 1539 1019
rect 111 1004 115 1008
rect 1095 1004 1099 1008
rect 251 999 252 1003
rect 252 999 255 1003
rect 379 999 383 1003
rect 423 999 427 1003
rect 519 999 523 1003
rect 547 999 551 1003
rect 619 999 623 1003
rect 731 999 732 1003
rect 732 999 735 1003
rect 803 999 804 1003
rect 804 999 807 1003
rect 867 999 868 1003
rect 868 999 871 1003
rect 927 999 928 1003
rect 928 999 931 1003
rect 995 999 996 1003
rect 996 999 999 1003
rect 1055 999 1059 1003
rect 1159 1004 1163 1008
rect 1231 1004 1235 1008
rect 1303 1004 1307 1008
rect 1383 1004 1387 1008
rect 1463 1004 1467 1008
rect 1543 1004 1547 1008
rect 1623 1004 1627 1008
rect 1651 1015 1655 1019
rect 1723 1015 1727 1019
rect 1815 1015 1819 1019
rect 1867 1015 1871 1019
rect 1915 1015 1919 1019
rect 1695 1004 1699 1008
rect 1759 1004 1763 1008
rect 1823 1004 1827 1008
rect 1135 996 1139 1000
rect 111 987 115 991
rect 223 984 227 988
rect 271 984 275 988
rect 335 984 339 988
rect 407 984 411 988
rect 479 984 483 988
rect 559 984 563 988
rect 631 984 635 988
rect 703 984 707 988
rect 775 984 779 988
rect 839 984 843 988
rect 903 984 907 988
rect 967 984 971 988
rect 1039 984 1043 988
rect 1095 987 1099 991
rect 1187 991 1188 995
rect 1188 991 1191 995
rect 1259 991 1260 995
rect 1260 991 1263 995
rect 1331 991 1332 995
rect 1332 991 1335 995
rect 1339 991 1343 995
rect 1487 991 1488 995
rect 1488 991 1491 995
rect 1527 991 1531 995
rect 1651 991 1652 995
rect 1652 991 1655 995
rect 1723 991 1724 995
rect 1724 991 1727 995
rect 1787 991 1788 995
rect 1788 991 1791 995
rect 1867 995 1871 999
rect 1887 1004 1891 1008
rect 1951 1004 1955 1008
rect 1915 991 1916 995
rect 1916 991 1919 995
rect 2119 996 2123 1000
rect 1135 979 1139 983
rect 1159 976 1163 980
rect 1231 976 1235 980
rect 1303 976 1307 980
rect 1383 976 1387 980
rect 1463 976 1467 980
rect 1543 976 1547 980
rect 1623 976 1627 980
rect 1695 976 1699 980
rect 1759 976 1763 980
rect 1823 976 1827 980
rect 1887 976 1891 980
rect 1951 976 1955 980
rect 2119 979 2123 983
rect 111 965 115 969
rect 151 968 155 972
rect 215 968 219 972
rect 287 968 291 972
rect 367 968 371 972
rect 447 968 451 972
rect 527 968 531 972
rect 599 968 603 972
rect 671 968 675 972
rect 735 968 739 972
rect 799 968 803 972
rect 863 968 867 972
rect 927 968 931 972
rect 991 968 995 972
rect 1047 968 1051 972
rect 1095 965 1099 969
rect 239 959 243 963
rect 111 948 115 952
rect 207 951 211 955
rect 279 951 283 955
rect 359 951 363 955
rect 711 959 715 963
rect 1135 961 1139 965
rect 1239 964 1243 968
rect 1303 964 1307 968
rect 1375 964 1379 968
rect 1439 964 1443 968
rect 1511 964 1515 968
rect 1583 964 1587 968
rect 1655 964 1659 968
rect 1727 964 1731 968
rect 1799 964 1803 968
rect 1871 964 1875 968
rect 1943 964 1947 968
rect 2015 964 2019 968
rect 2071 964 2075 968
rect 2119 961 2123 965
rect 471 951 472 955
rect 472 951 475 955
rect 483 951 487 955
rect 663 951 667 955
rect 727 951 731 955
rect 791 951 795 955
rect 855 951 859 955
rect 919 951 923 955
rect 999 951 1003 955
rect 1027 951 1031 955
rect 1611 955 1615 959
rect 1095 948 1099 952
rect 151 940 155 944
rect 215 940 219 944
rect 287 940 291 944
rect 367 940 371 944
rect 447 940 451 944
rect 527 940 531 944
rect 599 940 603 944
rect 671 940 675 944
rect 735 940 739 944
rect 799 940 803 944
rect 863 940 867 944
rect 927 940 931 944
rect 991 940 995 944
rect 1047 940 1051 944
rect 1135 944 1139 948
rect 1295 947 1299 951
rect 1367 947 1371 951
rect 1383 947 1387 951
rect 1503 947 1507 951
rect 1535 947 1536 951
rect 1536 947 1539 951
rect 1647 947 1651 951
rect 1719 947 1723 951
rect 1779 947 1783 951
rect 1863 947 1867 951
rect 1991 947 1995 951
rect 2119 944 2123 948
rect 1239 936 1243 940
rect 1303 936 1307 940
rect 1375 936 1379 940
rect 1439 936 1443 940
rect 1511 936 1515 940
rect 1583 936 1587 940
rect 1655 936 1659 940
rect 1727 936 1731 940
rect 1799 936 1803 940
rect 1871 936 1875 940
rect 1943 936 1947 940
rect 2007 939 2011 943
rect 2015 936 2019 940
rect 2071 936 2075 940
rect 159 927 163 931
rect 207 927 211 931
rect 279 927 283 931
rect 359 927 363 931
rect 483 927 487 931
rect 519 927 523 931
rect 655 927 659 931
rect 663 927 667 931
rect 727 927 731 931
rect 791 927 795 931
rect 855 927 859 931
rect 919 927 923 931
rect 1027 927 1031 931
rect 1055 927 1059 931
rect 171 915 175 919
rect 243 915 247 919
rect 303 915 307 919
rect 387 915 391 919
rect 471 915 475 919
rect 547 915 551 919
rect 555 915 559 919
rect 627 915 631 919
rect 699 915 703 919
rect 771 915 775 919
rect 843 915 847 919
rect 999 915 1003 919
rect 1027 915 1031 919
rect 1295 923 1299 927
rect 1367 923 1371 927
rect 1447 923 1451 927
rect 1503 923 1507 927
rect 1611 923 1615 927
rect 1647 923 1651 927
rect 1719 923 1723 927
rect 1787 923 1791 927
rect 1863 923 1867 927
rect 1991 923 1995 927
rect 2087 923 2091 927
rect 1339 915 1343 919
rect 135 904 139 908
rect 183 904 187 908
rect 255 904 259 908
rect 327 904 331 908
rect 399 904 403 908
rect 463 904 467 908
rect 527 904 531 908
rect 599 904 603 908
rect 671 904 675 908
rect 743 904 747 908
rect 815 904 819 908
rect 895 904 899 908
rect 983 904 987 908
rect 1047 904 1051 908
rect 111 896 115 900
rect 1095 896 1099 900
rect 159 891 160 895
rect 160 891 163 895
rect 171 891 175 895
rect 243 891 247 895
rect 351 891 352 895
rect 352 891 355 895
rect 387 891 391 895
rect 555 891 556 895
rect 556 891 559 895
rect 627 891 628 895
rect 628 891 631 895
rect 699 891 700 895
rect 700 891 703 895
rect 771 891 772 895
rect 772 891 775 895
rect 843 891 844 895
rect 844 891 847 895
rect 919 891 920 895
rect 920 891 923 895
rect 1027 891 1031 895
rect 1287 896 1291 900
rect 1087 891 1091 895
rect 1363 907 1367 911
rect 1383 907 1387 911
rect 1467 907 1471 911
rect 1495 907 1499 911
rect 1611 907 1615 911
rect 1691 907 1695 911
rect 1771 907 1775 911
rect 1779 907 1783 911
rect 1871 903 1875 907
rect 1907 907 1911 911
rect 1995 907 1999 911
rect 1327 896 1331 900
rect 1375 896 1379 900
rect 1423 896 1427 900
rect 1479 896 1483 900
rect 1551 896 1555 900
rect 1623 896 1627 900
rect 1703 896 1707 900
rect 1791 896 1795 900
rect 1879 896 1883 900
rect 1967 896 1971 900
rect 2063 896 2067 900
rect 1135 888 1139 892
rect 111 879 115 883
rect 135 876 139 880
rect 183 876 187 880
rect 255 876 259 880
rect 327 876 331 880
rect 399 876 403 880
rect 463 876 467 880
rect 527 876 531 880
rect 599 876 603 880
rect 671 876 675 880
rect 743 876 747 880
rect 815 876 819 880
rect 895 876 899 880
rect 983 876 987 880
rect 1047 876 1051 880
rect 1095 879 1099 883
rect 1207 883 1211 887
rect 2119 888 2123 892
rect 1363 883 1367 887
rect 1447 883 1448 887
rect 1448 883 1451 887
rect 1467 883 1471 887
rect 1559 883 1563 887
rect 1611 883 1615 887
rect 1691 883 1695 887
rect 1771 883 1775 887
rect 1907 883 1908 887
rect 1908 883 1911 887
rect 1995 883 1996 887
rect 1996 883 1999 887
rect 2087 883 2088 887
rect 2088 883 2091 887
rect 655 867 659 871
rect 919 867 923 871
rect 1135 871 1139 875
rect 1287 868 1291 872
rect 1327 868 1331 872
rect 1375 868 1379 872
rect 1423 868 1427 872
rect 1479 868 1483 872
rect 1551 868 1555 872
rect 1623 868 1627 872
rect 1703 868 1707 872
rect 1791 868 1795 872
rect 1879 868 1883 872
rect 1967 868 1971 872
rect 2063 868 2067 872
rect 2119 871 2123 875
rect 111 857 115 861
rect 135 860 139 864
rect 175 860 179 864
rect 215 860 219 864
rect 279 860 283 864
rect 343 860 347 864
rect 399 860 403 864
rect 463 860 467 864
rect 535 860 539 864
rect 615 860 619 864
rect 711 860 715 864
rect 823 860 827 864
rect 943 860 947 864
rect 1047 860 1051 864
rect 1095 857 1099 861
rect 903 851 907 855
rect 1135 853 1139 857
rect 1159 856 1163 860
rect 1199 856 1203 860
rect 1263 856 1267 860
rect 1327 856 1331 860
rect 1399 856 1403 860
rect 1471 856 1475 860
rect 1543 856 1547 860
rect 1623 856 1627 860
rect 1703 856 1707 860
rect 1775 856 1779 860
rect 1855 856 1859 860
rect 1935 856 1939 860
rect 2015 856 2019 860
rect 2071 856 2075 860
rect 2119 853 2123 857
rect 111 840 115 844
rect 163 843 164 847
rect 164 843 167 847
rect 203 843 204 847
rect 204 843 207 847
rect 271 843 275 847
rect 303 843 304 847
rect 304 843 307 847
rect 407 843 411 847
rect 471 843 475 847
rect 607 843 611 847
rect 703 843 707 847
rect 847 843 848 847
rect 848 843 851 847
rect 859 843 863 847
rect 1095 840 1099 844
rect 135 832 139 836
rect 175 832 179 836
rect 215 832 219 836
rect 279 832 283 836
rect 343 832 347 836
rect 399 832 403 836
rect 463 832 467 836
rect 535 832 539 836
rect 615 832 619 836
rect 711 832 715 836
rect 823 832 827 836
rect 943 832 947 836
rect 1047 832 1051 836
rect 1135 836 1139 840
rect 1143 839 1147 843
rect 1255 839 1259 843
rect 1319 839 1323 843
rect 1391 839 1395 843
rect 1463 839 1467 843
rect 1495 839 1496 843
rect 1496 839 1499 843
rect 1615 839 1619 843
rect 1695 839 1699 843
rect 1767 839 1771 843
rect 1783 839 1787 843
rect 1871 839 1875 843
rect 1899 839 1903 843
rect 2063 839 2067 843
rect 2079 839 2083 843
rect 2119 836 2123 840
rect 1087 827 1091 831
rect 155 819 159 823
rect 163 819 167 823
rect 203 819 207 823
rect 271 819 275 823
rect 351 819 355 823
rect 479 819 483 823
rect 599 819 603 823
rect 607 819 611 823
rect 703 819 707 823
rect 843 819 847 823
rect 1143 819 1147 823
rect 1159 828 1163 832
rect 1199 828 1203 832
rect 1263 828 1267 832
rect 1327 828 1331 832
rect 1399 828 1403 832
rect 1471 828 1475 832
rect 1543 828 1547 832
rect 1623 828 1627 832
rect 1703 828 1707 832
rect 1775 828 1779 832
rect 1855 828 1859 832
rect 1935 828 1939 832
rect 2015 828 2019 832
rect 2071 828 2075 832
rect 1207 815 1211 819
rect 1255 815 1259 819
rect 1319 815 1323 819
rect 1391 815 1395 819
rect 1463 815 1467 819
rect 1559 815 1563 819
rect 1615 815 1619 819
rect 1695 815 1699 819
rect 1767 815 1771 819
rect 1899 815 1903 819
rect 1999 815 2003 819
rect 2007 815 2011 819
rect 2063 815 2067 819
rect 135 796 139 800
rect 163 807 167 811
rect 203 807 207 811
rect 323 807 327 811
rect 379 807 383 811
rect 407 807 411 811
rect 471 807 475 811
rect 483 807 487 811
rect 547 807 551 811
rect 719 807 723 811
rect 763 807 767 811
rect 903 807 907 811
rect 923 807 927 811
rect 1011 807 1015 811
rect 175 796 179 800
rect 215 796 219 800
rect 279 796 283 800
rect 335 796 339 800
rect 391 796 395 800
rect 455 796 459 800
rect 519 796 523 800
rect 583 796 587 800
rect 655 796 659 800
rect 735 796 739 800
rect 815 796 819 800
rect 895 796 899 800
rect 983 796 987 800
rect 1047 796 1051 800
rect 111 788 115 792
rect 599 791 603 795
rect 155 783 159 787
rect 203 783 204 787
rect 204 783 207 787
rect 323 783 327 787
rect 379 783 383 787
rect 483 783 484 787
rect 484 783 487 787
rect 547 783 548 787
rect 548 783 551 787
rect 555 783 559 787
rect 763 783 764 787
rect 764 783 767 787
rect 843 783 844 787
rect 844 783 847 787
rect 923 783 924 787
rect 924 783 927 787
rect 1011 783 1012 787
rect 1012 783 1015 787
rect 1187 795 1191 799
rect 1303 795 1307 799
rect 1643 795 1647 799
rect 1739 795 1743 799
rect 1783 795 1787 799
rect 1831 795 1835 799
rect 1867 795 1871 799
rect 1947 795 1951 799
rect 2079 795 2083 799
rect 1095 788 1099 792
rect 1159 784 1163 788
rect 1239 784 1243 788
rect 1343 784 1347 788
rect 1447 784 1451 788
rect 1551 784 1555 788
rect 1655 784 1659 788
rect 1751 784 1755 788
rect 1839 784 1843 788
rect 1919 784 1923 788
rect 2007 784 2011 788
rect 2071 784 2075 788
rect 1135 776 1139 780
rect 111 771 115 775
rect 135 768 139 772
rect 175 768 179 772
rect 215 768 219 772
rect 279 768 283 772
rect 335 768 339 772
rect 391 768 395 772
rect 455 768 459 772
rect 519 768 523 772
rect 583 768 587 772
rect 655 768 659 772
rect 735 768 739 772
rect 815 768 819 772
rect 895 768 899 772
rect 983 768 987 772
rect 1047 768 1051 772
rect 1095 771 1099 775
rect 1187 771 1188 775
rect 1188 771 1191 775
rect 1303 775 1307 779
rect 2119 776 2123 780
rect 1311 771 1315 775
rect 1519 771 1523 775
rect 1643 771 1647 775
rect 1739 771 1743 775
rect 1867 771 1868 775
rect 1868 771 1871 775
rect 1947 771 1948 775
rect 1948 771 1951 775
rect 1999 771 2003 775
rect 2087 771 2091 775
rect 111 753 115 757
rect 135 756 139 760
rect 207 756 211 760
rect 295 756 299 760
rect 375 756 379 760
rect 447 756 451 760
rect 519 756 523 760
rect 583 756 587 760
rect 639 756 643 760
rect 687 756 691 760
rect 743 756 747 760
rect 799 756 803 760
rect 855 756 859 760
rect 1135 759 1139 763
rect 1095 753 1099 757
rect 1159 756 1163 760
rect 1239 756 1243 760
rect 1343 756 1347 760
rect 1447 756 1451 760
rect 1551 756 1555 760
rect 1655 756 1659 760
rect 1751 756 1755 760
rect 1839 756 1843 760
rect 1919 756 1923 760
rect 2007 756 2011 760
rect 2071 756 2075 760
rect 2119 759 2123 763
rect 111 736 115 740
rect 163 739 164 743
rect 164 739 167 743
rect 287 739 291 743
rect 319 739 320 743
rect 320 739 323 743
rect 391 739 395 743
rect 419 739 423 743
rect 679 739 683 743
rect 715 739 716 743
rect 716 739 719 743
rect 727 739 731 743
rect 847 739 851 743
rect 863 739 867 743
rect 1135 741 1139 745
rect 1159 744 1163 748
rect 1199 744 1203 748
rect 1239 744 1243 748
rect 1287 744 1291 748
rect 1359 744 1363 748
rect 1439 744 1443 748
rect 1527 744 1531 748
rect 1615 744 1619 748
rect 1711 744 1715 748
rect 1807 744 1811 748
rect 1903 744 1907 748
rect 1999 744 2003 748
rect 2071 744 2075 748
rect 2119 741 2123 745
rect 1095 736 1099 740
rect 1343 735 1347 739
rect 135 728 139 732
rect 207 728 211 732
rect 295 728 299 732
rect 375 728 379 732
rect 447 728 451 732
rect 519 728 523 732
rect 583 728 587 732
rect 639 728 643 732
rect 687 728 691 732
rect 743 728 747 732
rect 799 728 803 732
rect 855 728 859 732
rect 1135 724 1139 728
rect 1187 727 1188 731
rect 1188 727 1191 731
rect 1227 727 1228 731
rect 1228 727 1231 731
rect 1279 727 1283 731
rect 1351 727 1355 731
rect 1431 727 1435 731
rect 1607 727 1611 731
rect 1703 727 1707 731
rect 1719 727 1723 731
rect 1831 727 1832 731
rect 1832 727 1835 731
rect 2079 727 2083 731
rect 2119 724 2123 728
rect 159 715 163 719
rect 287 715 291 719
rect 419 715 423 719
rect 555 715 559 719
rect 607 715 611 719
rect 679 715 683 719
rect 791 715 795 719
rect 847 715 851 719
rect 1159 716 1163 720
rect 1199 716 1203 720
rect 1239 716 1243 720
rect 1287 716 1291 720
rect 1359 716 1363 720
rect 1439 716 1443 720
rect 1527 716 1531 720
rect 1615 716 1619 720
rect 1711 716 1715 720
rect 1807 716 1811 720
rect 1903 716 1907 720
rect 1999 716 2003 720
rect 2071 716 2075 720
rect 727 707 731 711
rect 863 707 867 711
rect 171 699 175 703
rect 235 699 239 703
rect 283 699 287 703
rect 319 699 323 703
rect 391 699 395 703
rect 411 699 415 703
rect 483 699 487 703
rect 631 699 635 703
rect 655 699 659 703
rect 735 699 739 703
rect 815 699 819 703
rect 907 699 911 703
rect 1187 703 1191 707
rect 1227 703 1231 707
rect 1279 703 1283 707
rect 1351 703 1355 707
rect 1431 703 1435 707
rect 1519 703 1523 707
rect 1607 703 1611 707
rect 1703 703 1707 707
rect 1987 703 1991 707
rect 2087 703 2091 707
rect 1311 695 1315 699
rect 1535 695 1539 699
rect 1719 695 1723 699
rect 135 688 139 692
rect 183 688 187 692
rect 247 688 251 692
rect 311 688 315 692
rect 383 688 387 692
rect 455 688 459 692
rect 519 688 523 692
rect 583 688 587 692
rect 647 688 651 692
rect 711 688 715 692
rect 767 688 771 692
rect 823 688 827 692
rect 879 688 883 692
rect 943 688 947 692
rect 1275 687 1279 691
rect 1323 687 1327 691
rect 1343 687 1347 691
rect 1563 687 1567 691
rect 1627 687 1631 691
rect 111 680 115 684
rect 1095 680 1099 684
rect 1711 683 1715 687
rect 1731 687 1735 691
rect 1859 687 1863 691
rect 1931 687 1935 691
rect 2059 687 2063 691
rect 2079 687 2083 691
rect 159 675 160 679
rect 160 675 163 679
rect 171 675 175 679
rect 275 675 276 679
rect 276 675 279 679
rect 283 675 287 679
rect 411 675 412 679
rect 412 675 415 679
rect 483 675 484 679
rect 484 675 487 679
rect 535 675 539 679
rect 607 675 608 679
rect 608 675 611 679
rect 631 675 635 679
rect 791 675 792 679
rect 792 675 795 679
rect 907 675 908 679
rect 908 675 911 679
rect 967 675 968 679
rect 968 675 971 679
rect 1239 676 1243 680
rect 1287 676 1291 680
rect 1335 676 1339 680
rect 1391 676 1395 680
rect 1447 676 1451 680
rect 1511 676 1515 680
rect 1575 676 1579 680
rect 1639 676 1643 680
rect 1703 676 1707 680
rect 1767 676 1771 680
rect 1831 676 1835 680
rect 1895 676 1899 680
rect 1959 676 1963 680
rect 2023 676 2027 680
rect 2071 676 2075 680
rect 1135 668 1139 672
rect 2119 668 2123 672
rect 111 663 115 667
rect 135 660 139 664
rect 183 660 187 664
rect 247 660 251 664
rect 311 660 315 664
rect 383 660 387 664
rect 455 660 459 664
rect 519 660 523 664
rect 583 660 587 664
rect 647 660 651 664
rect 711 660 715 664
rect 767 660 771 664
rect 823 660 827 664
rect 879 660 883 664
rect 943 660 947 664
rect 1095 663 1099 667
rect 1267 663 1268 667
rect 1268 663 1271 667
rect 1275 663 1279 667
rect 1323 663 1327 667
rect 1471 663 1472 667
rect 1472 663 1475 667
rect 1535 663 1536 667
rect 1536 663 1539 667
rect 1563 663 1567 667
rect 1627 663 1631 667
rect 1731 663 1732 667
rect 1732 663 1735 667
rect 1859 663 1860 667
rect 1860 663 1863 667
rect 1931 663 1935 667
rect 1987 663 1988 667
rect 1988 663 1991 667
rect 2051 663 2052 667
rect 2052 663 2055 667
rect 2059 663 2063 667
rect 1135 651 1139 655
rect 1239 648 1243 652
rect 1287 648 1291 652
rect 1335 648 1339 652
rect 1391 648 1395 652
rect 1447 648 1451 652
rect 1511 648 1515 652
rect 1575 648 1579 652
rect 1639 648 1643 652
rect 1703 648 1707 652
rect 1767 648 1771 652
rect 1831 648 1835 652
rect 1895 648 1899 652
rect 1959 648 1963 652
rect 2023 648 2027 652
rect 2071 648 2075 652
rect 2119 651 2123 655
rect 111 637 115 641
rect 159 640 163 644
rect 215 640 219 644
rect 287 640 291 644
rect 367 640 371 644
rect 455 640 459 644
rect 543 640 547 644
rect 631 640 635 644
rect 719 640 723 644
rect 799 640 803 644
rect 871 640 875 644
rect 951 640 955 644
rect 1031 640 1035 644
rect 1095 637 1099 641
rect 1135 633 1139 637
rect 1279 636 1283 640
rect 1319 636 1323 640
rect 1367 636 1371 640
rect 1423 636 1427 640
rect 1479 636 1483 640
rect 1535 636 1539 640
rect 1591 636 1595 640
rect 1647 636 1651 640
rect 1719 636 1723 640
rect 1799 636 1803 640
rect 1879 636 1883 640
rect 1967 636 1971 640
rect 2063 636 2067 640
rect 2119 633 2123 637
rect 111 620 115 624
rect 207 623 211 627
rect 235 623 239 627
rect 263 623 267 627
rect 391 623 392 627
rect 392 623 395 627
rect 403 623 407 627
rect 655 623 656 627
rect 656 623 659 627
rect 791 623 795 627
rect 815 623 819 627
rect 943 623 947 627
rect 1023 623 1027 627
rect 1039 623 1043 627
rect 1343 627 1347 631
rect 1095 620 1099 624
rect 159 612 163 616
rect 215 612 219 616
rect 287 612 291 616
rect 367 612 371 616
rect 455 612 459 616
rect 543 612 547 616
rect 631 612 635 616
rect 719 612 723 616
rect 799 612 803 616
rect 871 612 875 616
rect 951 612 955 616
rect 1031 612 1035 616
rect 1135 616 1139 620
rect 1307 619 1308 623
rect 1308 619 1311 623
rect 1359 619 1363 623
rect 1407 619 1411 623
rect 1711 627 1715 631
rect 1527 619 1531 623
rect 1575 619 1579 623
rect 1639 619 1643 623
rect 1711 619 1715 623
rect 1791 619 1795 623
rect 1871 619 1875 623
rect 1959 619 1963 623
rect 2071 619 2075 623
rect 2119 616 2123 620
rect 1279 608 1283 612
rect 1319 608 1323 612
rect 1367 608 1371 612
rect 1423 608 1427 612
rect 1479 608 1483 612
rect 1535 608 1539 612
rect 1591 608 1595 612
rect 1647 608 1651 612
rect 1719 608 1723 612
rect 1799 608 1803 612
rect 1879 608 1883 612
rect 1967 608 1971 612
rect 2063 608 2067 612
rect 183 599 187 603
rect 207 599 211 603
rect 275 599 279 603
rect 403 599 407 603
rect 535 599 539 603
rect 647 599 651 603
rect 727 599 731 603
rect 791 599 795 603
rect 879 599 883 603
rect 943 599 947 603
rect 1023 599 1027 603
rect 335 591 339 595
rect 943 591 947 595
rect 1267 595 1271 599
rect 1307 595 1311 599
rect 1359 595 1363 599
rect 1407 595 1411 599
rect 1471 595 1475 599
rect 1527 595 1531 599
rect 1631 595 1635 599
rect 1639 595 1643 599
rect 1711 595 1715 599
rect 1791 595 1795 599
rect 1871 595 1875 599
rect 1959 595 1963 599
rect 2051 595 2055 599
rect 243 583 247 587
rect 263 583 267 587
rect 371 579 375 583
rect 391 583 395 587
rect 411 583 415 587
rect 491 583 495 587
rect 683 583 687 587
rect 691 583 695 587
rect 811 583 815 587
rect 987 583 991 587
rect 1071 583 1075 587
rect 1343 583 1347 587
rect 1359 583 1363 587
rect 1403 583 1407 587
rect 1443 583 1447 587
rect 1491 583 1495 587
rect 1575 583 1579 587
rect 1611 583 1615 587
rect 1791 583 1795 587
rect 1871 583 1875 587
rect 1879 579 1883 583
rect 2051 583 2055 587
rect 2071 583 2075 587
rect 159 572 163 576
rect 207 572 211 576
rect 255 572 259 576
rect 311 572 315 576
rect 383 572 387 576
rect 463 572 467 576
rect 543 572 547 576
rect 623 572 627 576
rect 703 572 707 576
rect 783 572 787 576
rect 855 572 859 576
rect 927 572 931 576
rect 999 572 1003 576
rect 1047 572 1051 576
rect 1335 572 1339 576
rect 1375 572 1379 576
rect 1415 572 1419 576
rect 1463 572 1467 576
rect 1519 572 1523 576
rect 1583 572 1587 576
rect 1655 572 1659 576
rect 1727 572 1731 576
rect 1807 572 1811 576
rect 1887 572 1891 576
rect 1975 572 1979 576
rect 2063 572 2067 576
rect 111 564 115 568
rect 1095 564 1099 568
rect 183 559 184 563
rect 184 559 187 563
rect 231 559 232 563
rect 232 559 235 563
rect 243 559 247 563
rect 335 559 336 563
rect 336 559 339 563
rect 411 559 412 563
rect 412 559 415 563
rect 491 559 492 563
rect 492 559 495 563
rect 583 559 587 563
rect 647 559 648 563
rect 648 559 651 563
rect 683 559 687 563
rect 811 559 812 563
rect 812 559 815 563
rect 879 559 880 563
rect 880 559 883 563
rect 943 559 947 563
rect 987 559 991 563
rect 1135 564 1139 568
rect 1359 559 1360 563
rect 1360 559 1363 563
rect 1403 559 1404 563
rect 1404 559 1407 563
rect 1443 559 1444 563
rect 1444 559 1447 563
rect 1491 559 1492 563
rect 1492 559 1495 563
rect 1503 559 1507 563
rect 1611 559 1612 563
rect 1612 559 1615 563
rect 1631 563 1635 567
rect 1679 559 1680 563
rect 1680 559 1683 563
rect 2119 564 2123 568
rect 1791 559 1795 563
rect 1871 559 1875 563
rect 1999 559 2000 563
rect 2000 559 2003 563
rect 2051 559 2055 563
rect 111 547 115 551
rect 159 544 163 548
rect 207 544 211 548
rect 255 544 259 548
rect 311 544 315 548
rect 383 544 387 548
rect 463 544 467 548
rect 543 544 547 548
rect 623 544 627 548
rect 703 544 707 548
rect 783 544 787 548
rect 855 544 859 548
rect 927 544 931 548
rect 999 544 1003 548
rect 1047 544 1051 548
rect 1095 547 1099 551
rect 1135 547 1139 551
rect 1335 544 1339 548
rect 1375 544 1379 548
rect 1415 544 1419 548
rect 1463 544 1467 548
rect 1519 544 1523 548
rect 1583 544 1587 548
rect 1655 544 1659 548
rect 1727 544 1731 548
rect 1807 544 1811 548
rect 1887 544 1891 548
rect 1975 544 1979 548
rect 2063 544 2067 548
rect 2119 547 2123 551
rect 1551 535 1555 539
rect 1679 535 1683 539
rect 111 521 115 525
rect 167 524 171 528
rect 223 524 227 528
rect 287 524 291 528
rect 359 524 363 528
rect 431 524 435 528
rect 511 524 515 528
rect 591 524 595 528
rect 663 524 667 528
rect 735 524 739 528
rect 807 524 811 528
rect 871 524 875 528
rect 935 524 939 528
rect 999 524 1003 528
rect 1047 524 1051 528
rect 1095 521 1099 525
rect 1135 525 1139 529
rect 1191 528 1195 532
rect 1239 528 1243 532
rect 1287 528 1291 532
rect 1343 528 1347 532
rect 1407 528 1411 532
rect 1479 528 1483 532
rect 1543 528 1547 532
rect 1607 528 1611 532
rect 1671 528 1675 532
rect 1735 528 1739 532
rect 1799 528 1803 532
rect 1863 528 1867 532
rect 1935 528 1939 532
rect 2007 528 2011 532
rect 2071 528 2075 532
rect 2119 525 2123 529
rect 967 515 971 519
rect 1207 515 1211 519
rect 1215 519 1219 523
rect 1759 519 1763 523
rect 111 504 115 508
rect 175 507 179 511
rect 351 507 355 511
rect 371 507 375 511
rect 395 507 399 511
rect 547 507 551 511
rect 691 507 692 511
rect 692 507 695 511
rect 863 507 867 511
rect 927 507 931 511
rect 991 507 995 511
rect 1039 507 1043 511
rect 1071 507 1072 511
rect 1072 507 1075 511
rect 1095 504 1099 508
rect 1135 508 1139 512
rect 1231 511 1235 515
rect 1279 511 1283 515
rect 1359 511 1363 515
rect 1443 511 1447 515
rect 1591 511 1595 515
rect 1663 511 1667 515
rect 1695 511 1696 515
rect 1696 511 1699 515
rect 1791 511 1795 515
rect 1855 511 1859 515
rect 1879 511 1883 515
rect 2063 511 2067 515
rect 2079 511 2083 515
rect 2119 508 2123 512
rect 167 496 171 500
rect 223 496 227 500
rect 287 496 291 500
rect 359 496 363 500
rect 431 496 435 500
rect 511 496 515 500
rect 591 496 595 500
rect 663 496 667 500
rect 735 496 739 500
rect 807 496 811 500
rect 871 496 875 500
rect 935 496 939 500
rect 999 496 1003 500
rect 1047 496 1051 500
rect 1191 500 1195 504
rect 1239 500 1243 504
rect 1287 500 1291 504
rect 1343 500 1347 504
rect 1407 500 1411 504
rect 1479 500 1483 504
rect 1543 500 1547 504
rect 1607 500 1611 504
rect 1671 500 1675 504
rect 1735 500 1739 504
rect 1799 500 1803 504
rect 1863 500 1867 504
rect 1935 500 1939 504
rect 2007 500 2011 504
rect 2071 500 2075 504
rect 231 487 235 491
rect 259 483 263 487
rect 351 483 355 487
rect 547 483 551 487
rect 583 483 587 487
rect 635 483 639 487
rect 863 483 867 487
rect 927 483 931 487
rect 991 483 995 487
rect 1039 483 1043 487
rect 1215 487 1219 491
rect 1231 487 1235 491
rect 1279 487 1283 491
rect 1443 487 1447 491
rect 1503 487 1507 491
rect 1551 487 1555 491
rect 1591 487 1595 491
rect 1663 487 1667 491
rect 1759 487 1763 491
rect 1791 487 1795 491
rect 1855 487 1859 491
rect 1967 487 1971 491
rect 1999 487 2003 491
rect 2063 487 2067 491
rect 175 471 179 475
rect 295 471 299 475
rect 395 471 399 475
rect 403 471 407 475
rect 483 471 487 475
rect 579 471 583 475
rect 699 471 703 475
rect 707 471 711 475
rect 771 471 775 475
rect 827 471 831 475
rect 883 471 887 475
rect 967 471 971 475
rect 987 471 991 475
rect 1035 471 1039 475
rect 1075 475 1079 479
rect 1351 475 1355 479
rect 1359 475 1363 479
rect 1587 475 1591 479
rect 1687 475 1691 479
rect 1695 475 1699 479
rect 1827 475 1831 479
rect 1915 475 1919 479
rect 2079 475 2083 479
rect 167 460 171 464
rect 231 460 235 464
rect 303 460 307 464
rect 375 460 379 464
rect 455 460 459 464
rect 535 460 539 464
rect 607 460 611 464
rect 679 460 683 464
rect 743 460 747 464
rect 799 460 803 464
rect 855 460 859 464
rect 903 460 907 464
rect 959 460 963 464
rect 1007 460 1011 464
rect 1047 460 1051 464
rect 1159 464 1163 468
rect 1263 464 1267 468
rect 1383 464 1387 468
rect 1495 464 1499 468
rect 1599 464 1603 468
rect 1703 464 1707 468
rect 1799 464 1803 468
rect 1847 467 1851 471
rect 1887 464 1891 468
rect 1983 464 1987 468
rect 2071 464 2075 468
rect 111 452 115 456
rect 159 447 163 451
rect 259 447 260 451
rect 260 447 263 451
rect 403 447 404 451
rect 404 447 407 451
rect 483 447 484 451
rect 484 447 487 451
rect 495 447 499 451
rect 635 447 636 451
rect 636 447 639 451
rect 707 447 708 451
rect 708 447 711 451
rect 771 447 772 451
rect 772 447 775 451
rect 827 447 828 451
rect 828 447 831 451
rect 883 447 884 451
rect 884 447 887 451
rect 1095 452 1099 456
rect 1135 456 1139 460
rect 2119 456 2123 460
rect 987 447 988 451
rect 988 447 991 451
rect 1035 447 1036 451
rect 1036 447 1039 451
rect 1167 451 1171 455
rect 1075 447 1076 451
rect 1076 447 1079 451
rect 1207 451 1211 455
rect 1351 451 1355 455
rect 1583 451 1587 455
rect 1591 451 1595 455
rect 1687 451 1691 455
rect 1827 451 1828 455
rect 1828 451 1831 455
rect 1915 451 1916 455
rect 1916 451 1919 455
rect 1967 451 1971 455
rect 2031 451 2035 455
rect 111 435 115 439
rect 167 432 171 436
rect 231 432 235 436
rect 303 432 307 436
rect 375 432 379 436
rect 455 432 459 436
rect 535 432 539 436
rect 607 432 611 436
rect 679 432 683 436
rect 743 432 747 436
rect 799 432 803 436
rect 855 432 859 436
rect 903 432 907 436
rect 959 432 963 436
rect 1007 432 1011 436
rect 1047 432 1051 436
rect 1095 435 1099 439
rect 1135 439 1139 443
rect 1159 436 1163 440
rect 1263 436 1267 440
rect 1383 436 1387 440
rect 1495 436 1499 440
rect 1599 436 1603 440
rect 1703 436 1707 440
rect 1799 436 1803 440
rect 1887 436 1891 440
rect 1983 436 1987 440
rect 2071 436 2075 440
rect 2119 439 2123 443
rect 111 417 115 421
rect 151 420 155 424
rect 215 420 219 424
rect 279 420 283 424
rect 351 420 355 424
rect 423 420 427 424
rect 487 420 491 424
rect 551 420 555 424
rect 615 420 619 424
rect 671 420 675 424
rect 727 420 731 424
rect 791 420 795 424
rect 855 420 859 424
rect 1095 417 1099 421
rect 1135 421 1139 425
rect 1159 424 1163 428
rect 1199 424 1203 428
rect 1255 424 1259 428
rect 1335 424 1339 428
rect 1415 424 1419 428
rect 1503 424 1507 428
rect 1591 424 1595 428
rect 1671 424 1675 428
rect 1751 424 1755 428
rect 1823 424 1827 428
rect 1887 424 1891 428
rect 1951 424 1955 428
rect 2023 424 2027 428
rect 2071 424 2075 428
rect 2119 421 2123 425
rect 699 411 703 415
rect 111 400 115 404
rect 207 403 211 407
rect 295 403 299 407
rect 391 403 395 407
rect 579 403 580 407
rect 580 403 583 407
rect 663 403 667 407
rect 719 403 723 407
rect 783 403 787 407
rect 847 403 851 407
rect 1095 400 1099 404
rect 1135 404 1139 408
rect 1187 407 1188 411
rect 1188 407 1191 411
rect 1247 407 1251 411
rect 1327 407 1331 411
rect 1407 407 1411 411
rect 1495 407 1499 411
rect 1511 407 1515 411
rect 1663 407 1667 411
rect 1743 407 1747 411
rect 1815 407 1819 411
rect 1847 407 1848 411
rect 1848 407 1851 411
rect 1923 407 1927 411
rect 2063 407 2067 411
rect 2083 407 2087 411
rect 2119 404 2123 408
rect 151 392 155 396
rect 215 392 219 396
rect 279 392 283 396
rect 351 392 355 396
rect 423 392 427 396
rect 487 392 491 396
rect 551 392 555 396
rect 615 392 619 396
rect 671 392 675 396
rect 727 392 731 396
rect 791 392 795 396
rect 855 392 859 396
rect 1159 396 1163 400
rect 1199 396 1203 400
rect 1255 396 1259 400
rect 1335 396 1339 400
rect 1415 396 1419 400
rect 1503 396 1507 400
rect 1591 396 1595 400
rect 1671 396 1675 400
rect 1751 396 1755 400
rect 1823 396 1827 400
rect 1887 396 1891 400
rect 1951 396 1955 400
rect 2023 396 2027 400
rect 2071 396 2075 400
rect 159 379 163 383
rect 495 379 499 383
rect 543 379 547 383
rect 603 379 607 383
rect 663 379 667 383
rect 719 379 723 383
rect 783 379 787 383
rect 847 379 851 383
rect 1167 383 1171 387
rect 1187 383 1191 387
rect 1247 383 1251 387
rect 1327 383 1331 387
rect 1407 383 1411 387
rect 1495 383 1499 387
rect 1583 383 1587 387
rect 1663 383 1667 387
rect 1743 383 1747 387
rect 1923 383 1927 387
rect 1999 383 2003 387
rect 2031 383 2035 387
rect 2063 383 2067 387
rect 1511 375 1515 379
rect 135 356 139 360
rect 175 356 179 360
rect 207 367 211 371
rect 243 367 247 371
rect 299 367 303 371
rect 391 367 395 371
rect 411 367 415 371
rect 499 367 503 371
rect 647 367 651 371
rect 659 367 663 371
rect 715 367 719 371
rect 1327 367 1331 371
rect 1371 367 1375 371
rect 1407 367 1411 371
rect 1451 367 1455 371
rect 1491 367 1495 371
rect 1571 367 1575 371
rect 1579 367 1583 371
rect 1643 367 1647 371
rect 1707 367 1711 371
rect 1815 367 1819 371
rect 1943 367 1947 371
rect 2083 367 2087 371
rect 215 356 219 360
rect 271 356 275 360
rect 335 356 339 360
rect 399 356 403 360
rect 463 356 467 360
rect 519 356 523 360
rect 575 356 579 360
rect 631 356 635 360
rect 687 356 691 360
rect 751 356 755 360
rect 1303 356 1307 360
rect 1343 356 1347 360
rect 1383 356 1387 360
rect 1423 356 1427 360
rect 1463 356 1467 360
rect 1503 356 1507 360
rect 1551 356 1555 360
rect 1615 356 1619 360
rect 1679 356 1683 360
rect 1751 356 1755 360
rect 1831 356 1835 360
rect 1919 356 1923 360
rect 2007 356 2011 360
rect 2071 356 2075 360
rect 111 348 115 352
rect 143 343 147 347
rect 243 343 244 347
rect 244 343 247 347
rect 299 343 300 347
rect 300 343 303 347
rect 371 343 375 347
rect 499 343 503 347
rect 543 343 544 347
rect 544 343 547 347
rect 603 343 604 347
rect 604 343 607 347
rect 659 343 660 347
rect 660 343 663 347
rect 715 343 716 347
rect 716 343 719 347
rect 1095 348 1099 352
rect 1135 348 1139 352
rect 2119 348 2123 352
rect 1327 343 1328 347
rect 1328 343 1331 347
rect 1371 343 1372 347
rect 1372 343 1375 347
rect 1407 343 1408 347
rect 1408 343 1411 347
rect 1451 343 1452 347
rect 1452 343 1455 347
rect 1491 343 1492 347
rect 1492 343 1495 347
rect 1543 343 1547 347
rect 1579 343 1580 347
rect 1580 343 1583 347
rect 1643 343 1644 347
rect 1644 343 1647 347
rect 1707 343 1708 347
rect 1708 343 1711 347
rect 1715 343 1719 347
rect 1787 343 1791 347
rect 1999 343 2003 347
rect 2079 343 2083 347
rect 111 331 115 335
rect 135 328 139 332
rect 175 328 179 332
rect 215 328 219 332
rect 271 328 275 332
rect 335 328 339 332
rect 399 328 403 332
rect 463 328 467 332
rect 519 328 523 332
rect 575 328 579 332
rect 631 328 635 332
rect 687 328 691 332
rect 751 328 755 332
rect 1095 331 1099 335
rect 1135 331 1139 335
rect 1303 328 1307 332
rect 1343 328 1347 332
rect 1383 328 1387 332
rect 1423 328 1427 332
rect 1463 328 1467 332
rect 1503 328 1507 332
rect 1551 328 1555 332
rect 1615 328 1619 332
rect 1679 328 1683 332
rect 1751 328 1755 332
rect 1831 328 1835 332
rect 1919 328 1923 332
rect 2007 328 2011 332
rect 2071 328 2075 332
rect 2119 331 2123 335
rect 371 319 375 323
rect 111 309 115 313
rect 135 312 139 316
rect 207 312 211 316
rect 295 312 299 316
rect 383 312 387 316
rect 471 312 475 316
rect 551 312 555 316
rect 623 312 627 316
rect 687 312 691 316
rect 751 312 755 316
rect 807 312 811 316
rect 871 312 875 316
rect 935 312 939 316
rect 1095 309 1099 313
rect 1135 309 1139 313
rect 1167 312 1171 316
rect 1207 312 1211 316
rect 1247 312 1251 316
rect 1295 312 1299 316
rect 1343 312 1347 316
rect 1391 312 1395 316
rect 1439 312 1443 316
rect 1495 312 1499 316
rect 1559 312 1563 316
rect 1623 312 1627 316
rect 1695 312 1699 316
rect 1775 312 1779 316
rect 1855 312 1859 316
rect 1935 312 1939 316
rect 2015 312 2019 316
rect 2071 312 2075 316
rect 2119 309 2123 313
rect 1319 303 1323 307
rect 111 292 115 296
rect 287 295 291 299
rect 303 295 307 299
rect 411 295 412 299
rect 412 295 415 299
rect 419 295 423 299
rect 647 295 648 299
rect 648 295 651 299
rect 723 295 727 299
rect 1095 292 1099 296
rect 1135 292 1139 296
rect 1175 295 1179 299
rect 135 284 139 288
rect 207 284 211 288
rect 295 284 299 288
rect 383 284 387 288
rect 471 284 475 288
rect 551 284 555 288
rect 623 284 627 288
rect 687 284 691 288
rect 751 284 755 288
rect 807 284 811 288
rect 871 284 875 288
rect 935 284 939 288
rect 1167 284 1171 288
rect 1207 284 1211 288
rect 1383 295 1387 299
rect 1463 303 1467 307
rect 1487 295 1491 299
rect 1519 295 1520 299
rect 1520 295 1523 299
rect 1571 295 1575 299
rect 1731 295 1735 299
rect 1927 295 1931 299
rect 1943 295 1947 299
rect 2007 295 2011 299
rect 2119 292 2123 296
rect 1247 284 1251 288
rect 1295 284 1299 288
rect 1343 284 1347 288
rect 1391 284 1395 288
rect 1439 284 1443 288
rect 1495 284 1499 288
rect 1559 284 1563 288
rect 1623 284 1627 288
rect 1695 284 1699 288
rect 1775 284 1779 288
rect 1855 284 1859 288
rect 1935 284 1939 288
rect 2015 284 2019 288
rect 2071 284 2075 288
rect 143 271 147 275
rect 287 271 291 275
rect 419 271 423 275
rect 539 271 543 275
rect 723 271 727 275
rect 907 271 911 275
rect 1319 271 1323 275
rect 1351 271 1355 275
rect 1383 271 1387 275
rect 1463 271 1467 275
rect 1487 271 1491 275
rect 1543 271 1547 275
rect 1731 271 1735 275
rect 1787 271 1791 275
rect 1863 271 1867 275
rect 1927 271 1931 275
rect 2079 271 2083 275
rect 187 259 191 263
rect 267 259 271 263
rect 303 259 307 263
rect 351 259 355 263
rect 391 259 395 263
rect 591 259 595 263
rect 611 259 615 263
rect 731 259 735 263
rect 787 259 791 263
rect 843 259 847 263
rect 1715 263 1719 267
rect 135 248 139 252
rect 199 248 203 252
rect 279 248 283 252
rect 359 248 363 252
rect 439 248 443 252
rect 511 248 515 252
rect 583 248 587 252
rect 647 248 651 252
rect 703 248 707 252
rect 759 248 763 252
rect 815 248 819 252
rect 879 248 883 252
rect 1175 251 1179 255
rect 1187 251 1191 255
rect 1235 251 1239 255
rect 1379 251 1383 255
rect 1423 251 1427 255
rect 1511 251 1515 255
rect 1519 251 1523 255
rect 1635 251 1639 255
rect 1715 251 1719 255
rect 1907 251 1911 255
rect 1975 251 1979 255
rect 2007 251 2011 255
rect 2027 251 2031 255
rect 111 240 115 244
rect 1095 240 1099 244
rect 143 235 147 239
rect 187 235 191 239
rect 267 235 271 239
rect 387 235 388 239
rect 388 235 391 239
rect 539 235 540 239
rect 540 235 543 239
rect 611 235 612 239
rect 612 235 615 239
rect 731 235 732 239
rect 732 235 735 239
rect 787 235 788 239
rect 788 235 791 239
rect 843 235 844 239
rect 844 235 847 239
rect 1159 240 1163 244
rect 1207 240 1211 244
rect 1271 240 1275 244
rect 1327 240 1331 244
rect 1391 240 1395 244
rect 1455 240 1459 244
rect 1527 240 1531 244
rect 1607 240 1611 244
rect 1687 240 1691 244
rect 1767 240 1771 244
rect 1839 240 1843 244
rect 1919 240 1923 244
rect 1999 240 2003 244
rect 2071 240 2075 244
rect 907 235 908 239
rect 908 235 911 239
rect 1135 232 1139 236
rect 2119 232 2123 236
rect 111 223 115 227
rect 135 220 139 224
rect 199 220 203 224
rect 279 220 283 224
rect 359 220 363 224
rect 439 220 443 224
rect 511 220 515 224
rect 583 220 587 224
rect 647 220 651 224
rect 703 220 707 224
rect 759 220 763 224
rect 815 220 819 224
rect 879 220 883 224
rect 1095 223 1099 227
rect 1187 227 1188 231
rect 1188 227 1191 231
rect 1235 227 1236 231
rect 1236 227 1239 231
rect 1279 227 1283 231
rect 1351 227 1352 231
rect 1352 227 1355 231
rect 1379 227 1383 231
rect 1479 227 1480 231
rect 1480 227 1483 231
rect 1511 227 1515 231
rect 1635 227 1636 231
rect 1636 227 1639 231
rect 1715 227 1716 231
rect 1716 227 1719 231
rect 1743 227 1747 231
rect 1863 227 1864 231
rect 1864 227 1867 231
rect 1907 227 1911 231
rect 2027 227 2028 231
rect 2028 227 2031 231
rect 2087 227 2091 231
rect 1135 215 1139 219
rect 1159 212 1163 216
rect 1207 212 1211 216
rect 1271 212 1275 216
rect 1327 212 1331 216
rect 1391 212 1395 216
rect 1455 212 1459 216
rect 1527 212 1531 216
rect 1607 212 1611 216
rect 1687 212 1691 216
rect 1767 212 1771 216
rect 1839 212 1843 216
rect 1919 212 1923 216
rect 1999 212 2003 216
rect 2071 212 2075 216
rect 2119 215 2123 219
rect 111 201 115 205
rect 135 204 139 208
rect 183 204 187 208
rect 231 204 235 208
rect 279 204 283 208
rect 327 204 331 208
rect 375 204 379 208
rect 415 204 419 208
rect 455 204 459 208
rect 503 204 507 208
rect 551 204 555 208
rect 599 204 603 208
rect 647 204 651 208
rect 695 204 699 208
rect 743 204 747 208
rect 1095 201 1099 205
rect 591 195 595 199
rect 1135 197 1139 201
rect 1159 200 1163 204
rect 1199 200 1203 204
rect 1263 200 1267 204
rect 1327 200 1331 204
rect 1399 200 1403 204
rect 1471 200 1475 204
rect 1543 200 1547 204
rect 1607 200 1611 204
rect 1671 200 1675 204
rect 1735 200 1739 204
rect 1807 200 1811 204
rect 1879 200 1883 204
rect 1951 200 1955 204
rect 2023 200 2027 204
rect 2071 200 2075 204
rect 2119 197 2123 201
rect 111 184 115 188
rect 175 187 179 191
rect 223 187 227 191
rect 271 187 275 191
rect 287 187 291 191
rect 351 187 352 191
rect 352 187 355 191
rect 135 176 139 180
rect 183 176 187 180
rect 231 176 235 180
rect 279 176 283 180
rect 327 176 331 180
rect 375 176 379 180
rect 495 187 499 191
rect 543 187 547 191
rect 591 187 595 191
rect 639 187 643 191
rect 687 187 691 191
rect 735 187 739 191
rect 1975 191 1979 195
rect 1095 184 1099 188
rect 415 176 419 180
rect 455 176 459 180
rect 503 176 507 180
rect 551 176 555 180
rect 599 176 603 180
rect 647 176 651 180
rect 695 176 699 180
rect 743 176 747 180
rect 1135 180 1139 184
rect 1171 183 1175 187
rect 1159 172 1163 176
rect 1391 183 1395 187
rect 1423 183 1424 187
rect 1424 183 1427 187
rect 1535 183 1539 187
rect 1551 183 1555 187
rect 1579 183 1583 187
rect 1871 183 1875 187
rect 1943 183 1947 187
rect 2015 183 2019 187
rect 2079 183 2083 187
rect 2119 180 2123 184
rect 1199 172 1203 176
rect 1263 172 1267 176
rect 1327 172 1331 176
rect 1399 172 1403 176
rect 1471 172 1475 176
rect 1543 172 1547 176
rect 1607 172 1611 176
rect 1671 172 1675 176
rect 1735 172 1739 176
rect 1807 172 1811 176
rect 1879 172 1883 176
rect 1951 172 1955 176
rect 2023 172 2027 176
rect 2071 172 2075 176
rect 143 163 147 167
rect 175 163 179 167
rect 223 163 227 167
rect 271 163 275 167
rect 495 163 499 167
rect 543 163 547 167
rect 591 163 595 167
rect 639 163 643 167
rect 687 163 691 167
rect 735 163 739 167
rect 567 155 571 159
rect 1279 159 1283 163
rect 1299 159 1303 163
rect 1391 159 1395 163
rect 1479 159 1483 163
rect 1535 159 1539 163
rect 1743 159 1747 163
rect 1871 159 1875 163
rect 1943 159 1947 163
rect 2015 159 2019 163
rect 2087 159 2091 163
rect 527 147 531 151
rect 1975 151 1979 155
rect 287 135 291 139
rect 1359 135 1363 139
rect 1551 135 1555 139
rect 171 127 175 131
rect 211 127 215 131
rect 247 127 251 131
rect 291 127 295 131
rect 335 127 339 131
rect 367 127 371 131
rect 407 127 411 131
rect 447 127 451 131
rect 491 127 495 131
rect 143 116 147 120
rect 183 116 187 120
rect 223 116 227 120
rect 263 116 267 120
rect 303 116 307 120
rect 343 116 347 120
rect 383 116 387 120
rect 423 116 427 120
rect 463 116 467 120
rect 503 116 507 120
rect 543 116 547 120
rect 583 116 587 120
rect 623 116 627 120
rect 663 116 667 120
rect 703 116 707 120
rect 743 116 747 120
rect 819 127 823 131
rect 867 127 871 131
rect 783 116 787 120
rect 831 116 835 120
rect 879 116 883 120
rect 927 116 931 120
rect 967 116 971 120
rect 1007 116 1011 120
rect 1143 127 1147 131
rect 1171 127 1175 131
rect 1235 127 1239 131
rect 1387 127 1391 131
rect 1439 127 1443 131
rect 1499 127 1503 131
rect 1579 127 1583 131
rect 1587 127 1591 131
rect 1635 127 1639 131
rect 1679 127 1683 131
rect 1715 127 1719 131
rect 1755 127 1759 131
rect 1795 127 1799 131
rect 1835 127 1839 131
rect 1931 127 1935 131
rect 2015 127 2019 131
rect 1047 116 1051 120
rect 1159 116 1163 120
rect 1207 116 1211 120
rect 1271 116 1275 120
rect 1335 116 1339 120
rect 1399 116 1403 120
rect 1455 116 1459 120
rect 1511 116 1515 120
rect 1559 116 1563 120
rect 1607 116 1611 120
rect 1647 116 1651 120
rect 1687 116 1691 120
rect 1727 116 1731 120
rect 1767 116 1771 120
rect 1807 116 1811 120
rect 1855 116 1859 120
rect 1903 116 1907 120
rect 1951 116 1955 120
rect 1991 116 1995 120
rect 2031 116 2035 120
rect 2079 127 2083 131
rect 2071 116 2075 120
rect 111 108 115 112
rect 171 103 172 107
rect 172 103 175 107
rect 211 103 212 107
rect 212 103 215 107
rect 247 103 248 107
rect 248 103 251 107
rect 291 103 292 107
rect 292 103 295 107
rect 331 103 332 107
rect 332 103 335 107
rect 367 103 368 107
rect 368 103 371 107
rect 407 103 408 107
rect 408 103 411 107
rect 447 103 448 107
rect 448 103 451 107
rect 491 103 492 107
rect 492 103 495 107
rect 527 103 528 107
rect 528 103 531 107
rect 567 103 568 107
rect 568 103 571 107
rect 819 103 823 107
rect 867 103 871 107
rect 1095 108 1099 112
rect 1135 108 1139 112
rect 1143 103 1147 107
rect 1235 103 1236 107
rect 1236 103 1239 107
rect 1299 103 1300 107
rect 1300 103 1303 107
rect 1359 103 1360 107
rect 1360 103 1363 107
rect 1387 103 1391 107
rect 1439 103 1443 107
rect 1499 103 1503 107
rect 1587 103 1588 107
rect 1588 103 1591 107
rect 1635 103 1636 107
rect 1636 103 1639 107
rect 1675 103 1676 107
rect 1676 103 1679 107
rect 1715 103 1716 107
rect 1716 103 1719 107
rect 1755 103 1756 107
rect 1756 103 1759 107
rect 1795 103 1796 107
rect 1796 103 1799 107
rect 1835 103 1836 107
rect 1836 103 1839 107
rect 1931 103 1932 107
rect 1932 103 1935 107
rect 1975 103 1976 107
rect 1976 103 1979 107
rect 2015 103 2019 107
rect 2119 108 2123 112
rect 111 91 115 95
rect 143 88 147 92
rect 183 88 187 92
rect 223 88 227 92
rect 263 88 267 92
rect 303 88 307 92
rect 343 88 347 92
rect 383 88 387 92
rect 423 88 427 92
rect 463 88 467 92
rect 503 88 507 92
rect 543 88 547 92
rect 583 88 587 92
rect 623 88 627 92
rect 663 88 667 92
rect 703 88 707 92
rect 743 88 747 92
rect 783 88 787 92
rect 831 88 835 92
rect 879 88 883 92
rect 927 88 931 92
rect 967 88 971 92
rect 1007 88 1011 92
rect 1047 88 1051 92
rect 1095 91 1099 95
rect 1135 91 1139 95
rect 1159 88 1163 92
rect 1207 88 1211 92
rect 1271 88 1275 92
rect 1335 88 1339 92
rect 1399 88 1403 92
rect 1455 88 1459 92
rect 1511 88 1515 92
rect 1559 88 1563 92
rect 1607 88 1611 92
rect 1647 88 1651 92
rect 1687 88 1691 92
rect 1727 88 1731 92
rect 1767 88 1771 92
rect 1807 88 1811 92
rect 1855 88 1859 92
rect 1903 88 1907 92
rect 1951 88 1955 92
rect 1991 88 1995 92
rect 2031 88 2035 92
rect 2071 88 2075 92
rect 2119 91 2123 95
<< m3 >>
rect 1135 2230 1139 2231
rect 1135 2225 1139 2226
rect 1687 2230 1691 2231
rect 1687 2225 1691 2226
rect 1727 2230 1731 2231
rect 1727 2225 1731 2226
rect 1767 2230 1771 2231
rect 1767 2225 1771 2226
rect 1807 2230 1811 2231
rect 1807 2225 1811 2226
rect 2119 2230 2123 2231
rect 2119 2225 2123 2226
rect 111 2214 115 2215
rect 111 2209 115 2210
rect 135 2214 139 2215
rect 135 2209 139 2210
rect 175 2214 179 2215
rect 175 2209 179 2210
rect 215 2214 219 2215
rect 215 2209 219 2210
rect 255 2214 259 2215
rect 255 2209 259 2210
rect 319 2214 323 2215
rect 319 2209 323 2210
rect 383 2214 387 2215
rect 383 2209 387 2210
rect 447 2214 451 2215
rect 447 2209 451 2210
rect 511 2214 515 2215
rect 511 2209 515 2210
rect 575 2214 579 2215
rect 575 2209 579 2210
rect 631 2214 635 2215
rect 631 2209 635 2210
rect 687 2214 691 2215
rect 687 2209 691 2210
rect 735 2214 739 2215
rect 735 2209 739 2210
rect 791 2214 795 2215
rect 791 2209 795 2210
rect 847 2214 851 2215
rect 847 2209 851 2210
rect 903 2214 907 2215
rect 903 2209 907 2210
rect 1095 2214 1099 2215
rect 1095 2209 1099 2210
rect 112 2206 114 2209
rect 134 2208 140 2209
rect 110 2205 116 2206
rect 110 2201 111 2205
rect 115 2201 116 2205
rect 134 2204 135 2208
rect 139 2204 140 2208
rect 134 2203 140 2204
rect 174 2208 180 2209
rect 174 2204 175 2208
rect 179 2204 180 2208
rect 174 2203 180 2204
rect 214 2208 220 2209
rect 214 2204 215 2208
rect 219 2204 220 2208
rect 214 2203 220 2204
rect 254 2208 260 2209
rect 254 2204 255 2208
rect 259 2204 260 2208
rect 254 2203 260 2204
rect 318 2208 324 2209
rect 318 2204 319 2208
rect 323 2204 324 2208
rect 318 2203 324 2204
rect 382 2208 388 2209
rect 382 2204 383 2208
rect 387 2204 388 2208
rect 382 2203 388 2204
rect 446 2208 452 2209
rect 446 2204 447 2208
rect 451 2204 452 2208
rect 446 2203 452 2204
rect 510 2208 516 2209
rect 510 2204 511 2208
rect 515 2204 516 2208
rect 510 2203 516 2204
rect 574 2208 580 2209
rect 574 2204 575 2208
rect 579 2204 580 2208
rect 574 2203 580 2204
rect 630 2208 636 2209
rect 630 2204 631 2208
rect 635 2204 636 2208
rect 630 2203 636 2204
rect 686 2208 692 2209
rect 686 2204 687 2208
rect 691 2204 692 2208
rect 686 2203 692 2204
rect 734 2208 740 2209
rect 734 2204 735 2208
rect 739 2204 740 2208
rect 734 2203 740 2204
rect 790 2208 796 2209
rect 790 2204 791 2208
rect 795 2204 796 2208
rect 790 2203 796 2204
rect 846 2208 852 2209
rect 846 2204 847 2208
rect 851 2204 852 2208
rect 846 2203 852 2204
rect 902 2208 908 2209
rect 902 2204 903 2208
rect 907 2204 908 2208
rect 1096 2206 1098 2209
rect 902 2203 908 2204
rect 1094 2205 1100 2206
rect 1136 2205 1138 2225
rect 1678 2223 1684 2224
rect 1678 2219 1679 2223
rect 1683 2219 1684 2223
rect 1678 2218 1684 2219
rect 110 2200 116 2201
rect 1094 2201 1095 2205
rect 1099 2201 1100 2205
rect 1094 2200 1100 2201
rect 1134 2204 1140 2205
rect 1134 2200 1135 2204
rect 1139 2200 1140 2204
rect 1134 2199 1140 2200
rect 162 2191 168 2192
rect 110 2188 116 2189
rect 110 2184 111 2188
rect 115 2184 116 2188
rect 162 2187 163 2191
rect 167 2187 168 2191
rect 162 2186 168 2187
rect 202 2191 208 2192
rect 202 2187 203 2191
rect 207 2187 208 2191
rect 202 2186 208 2187
rect 242 2191 248 2192
rect 242 2187 243 2191
rect 247 2187 248 2191
rect 242 2186 248 2187
rect 310 2191 316 2192
rect 310 2187 311 2191
rect 315 2187 316 2191
rect 310 2186 316 2187
rect 374 2191 380 2192
rect 374 2187 375 2191
rect 379 2187 380 2191
rect 374 2186 380 2187
rect 438 2191 444 2192
rect 438 2187 439 2191
rect 443 2187 444 2191
rect 438 2186 444 2187
rect 454 2191 460 2192
rect 454 2187 455 2191
rect 459 2187 460 2191
rect 454 2186 460 2187
rect 566 2191 572 2192
rect 566 2187 567 2191
rect 571 2187 572 2191
rect 566 2186 572 2187
rect 622 2191 628 2192
rect 622 2187 623 2191
rect 627 2187 628 2191
rect 622 2186 628 2187
rect 678 2191 684 2192
rect 678 2187 679 2191
rect 683 2187 684 2191
rect 678 2186 684 2187
rect 726 2191 732 2192
rect 726 2187 727 2191
rect 731 2187 732 2191
rect 726 2186 732 2187
rect 782 2191 788 2192
rect 782 2187 783 2191
rect 787 2187 788 2191
rect 782 2186 788 2187
rect 838 2191 844 2192
rect 838 2187 839 2191
rect 843 2187 844 2191
rect 838 2186 844 2187
rect 894 2191 900 2192
rect 894 2187 895 2191
rect 899 2187 900 2191
rect 894 2186 900 2187
rect 910 2191 916 2192
rect 910 2187 911 2191
rect 915 2187 916 2191
rect 910 2186 916 2187
rect 1094 2188 1100 2189
rect 110 2183 116 2184
rect 112 2155 114 2183
rect 134 2180 140 2181
rect 134 2176 135 2180
rect 139 2176 140 2180
rect 134 2175 140 2176
rect 136 2155 138 2175
rect 164 2168 166 2186
rect 174 2180 180 2181
rect 174 2176 175 2180
rect 179 2176 180 2180
rect 174 2175 180 2176
rect 162 2167 168 2168
rect 162 2163 163 2167
rect 167 2163 168 2167
rect 162 2162 168 2163
rect 176 2155 178 2175
rect 204 2168 206 2186
rect 214 2180 220 2181
rect 214 2176 215 2180
rect 219 2176 220 2180
rect 214 2175 220 2176
rect 202 2167 208 2168
rect 202 2163 203 2167
rect 207 2163 208 2167
rect 202 2162 208 2163
rect 216 2155 218 2175
rect 244 2168 246 2186
rect 254 2180 260 2181
rect 254 2176 255 2180
rect 259 2176 260 2180
rect 254 2175 260 2176
rect 242 2167 248 2168
rect 242 2163 243 2167
rect 247 2163 248 2167
rect 242 2162 248 2163
rect 256 2155 258 2175
rect 312 2168 314 2186
rect 318 2180 324 2181
rect 318 2176 319 2180
rect 323 2176 324 2180
rect 318 2175 324 2176
rect 310 2167 316 2168
rect 310 2163 311 2167
rect 315 2163 316 2167
rect 310 2162 316 2163
rect 320 2155 322 2175
rect 376 2168 378 2186
rect 382 2180 388 2181
rect 382 2176 383 2180
rect 387 2176 388 2180
rect 382 2175 388 2176
rect 374 2167 380 2168
rect 374 2163 375 2167
rect 379 2163 380 2167
rect 374 2162 380 2163
rect 384 2155 386 2175
rect 440 2168 442 2186
rect 446 2180 452 2181
rect 446 2176 447 2180
rect 451 2176 452 2180
rect 446 2175 452 2176
rect 438 2167 444 2168
rect 438 2163 439 2167
rect 443 2163 444 2167
rect 438 2162 444 2163
rect 448 2155 450 2175
rect 456 2156 458 2186
rect 510 2180 516 2181
rect 510 2176 511 2180
rect 515 2176 516 2180
rect 510 2175 516 2176
rect 454 2155 460 2156
rect 512 2155 514 2175
rect 568 2168 570 2186
rect 574 2180 580 2181
rect 574 2176 575 2180
rect 579 2176 580 2180
rect 574 2175 580 2176
rect 566 2167 572 2168
rect 566 2163 567 2167
rect 571 2163 572 2167
rect 566 2162 572 2163
rect 576 2155 578 2175
rect 624 2168 626 2186
rect 630 2180 636 2181
rect 630 2176 631 2180
rect 635 2176 636 2180
rect 630 2175 636 2176
rect 622 2167 628 2168
rect 622 2163 623 2167
rect 627 2163 628 2167
rect 622 2162 628 2163
rect 632 2155 634 2175
rect 680 2168 682 2186
rect 686 2180 692 2181
rect 686 2176 687 2180
rect 691 2176 692 2180
rect 686 2175 692 2176
rect 678 2167 684 2168
rect 678 2163 679 2167
rect 683 2163 684 2167
rect 678 2162 684 2163
rect 688 2155 690 2175
rect 728 2168 730 2186
rect 734 2180 740 2181
rect 734 2176 735 2180
rect 739 2176 740 2180
rect 734 2175 740 2176
rect 726 2167 732 2168
rect 726 2163 727 2167
rect 731 2163 732 2167
rect 726 2162 732 2163
rect 736 2155 738 2175
rect 784 2168 786 2186
rect 790 2180 796 2181
rect 790 2176 791 2180
rect 795 2176 796 2180
rect 790 2175 796 2176
rect 782 2167 788 2168
rect 782 2163 783 2167
rect 787 2163 788 2167
rect 782 2162 788 2163
rect 792 2155 794 2175
rect 840 2168 842 2186
rect 846 2180 852 2181
rect 846 2176 847 2180
rect 851 2176 852 2180
rect 846 2175 852 2176
rect 838 2167 844 2168
rect 838 2163 839 2167
rect 843 2163 844 2167
rect 838 2162 844 2163
rect 848 2155 850 2175
rect 896 2168 898 2186
rect 902 2180 908 2181
rect 902 2176 903 2180
rect 907 2176 908 2180
rect 902 2175 908 2176
rect 894 2167 900 2168
rect 894 2163 895 2167
rect 899 2163 900 2167
rect 894 2162 900 2163
rect 904 2155 906 2175
rect 912 2156 914 2186
rect 1094 2184 1095 2188
rect 1099 2184 1100 2188
rect 1094 2183 1100 2184
rect 1134 2187 1140 2188
rect 1134 2183 1135 2187
rect 1139 2183 1140 2187
rect 910 2155 916 2156
rect 1096 2155 1098 2183
rect 1134 2182 1140 2183
rect 1136 2179 1138 2182
rect 1135 2178 1139 2179
rect 1135 2173 1139 2174
rect 1159 2178 1163 2179
rect 1159 2173 1163 2174
rect 1199 2178 1203 2179
rect 1199 2173 1203 2174
rect 1239 2178 1243 2179
rect 1239 2173 1243 2174
rect 1279 2178 1283 2179
rect 1279 2173 1283 2174
rect 1335 2178 1339 2179
rect 1335 2173 1339 2174
rect 1391 2178 1395 2179
rect 1391 2173 1395 2174
rect 1455 2178 1459 2179
rect 1455 2173 1459 2174
rect 1527 2178 1531 2179
rect 1527 2173 1531 2174
rect 1591 2178 1595 2179
rect 1591 2173 1595 2174
rect 1663 2178 1667 2179
rect 1663 2173 1667 2174
rect 1136 2170 1138 2173
rect 1158 2172 1164 2173
rect 1134 2169 1140 2170
rect 1134 2165 1135 2169
rect 1139 2165 1140 2169
rect 1158 2168 1159 2172
rect 1163 2168 1164 2172
rect 1158 2167 1164 2168
rect 1198 2172 1204 2173
rect 1198 2168 1199 2172
rect 1203 2168 1204 2172
rect 1198 2167 1204 2168
rect 1238 2172 1244 2173
rect 1238 2168 1239 2172
rect 1243 2168 1244 2172
rect 1238 2167 1244 2168
rect 1278 2172 1284 2173
rect 1278 2168 1279 2172
rect 1283 2168 1284 2172
rect 1278 2167 1284 2168
rect 1334 2172 1340 2173
rect 1334 2168 1335 2172
rect 1339 2168 1340 2172
rect 1334 2167 1340 2168
rect 1390 2172 1396 2173
rect 1390 2168 1391 2172
rect 1395 2168 1396 2172
rect 1390 2167 1396 2168
rect 1454 2172 1460 2173
rect 1454 2168 1455 2172
rect 1459 2168 1460 2172
rect 1454 2167 1460 2168
rect 1526 2172 1532 2173
rect 1526 2168 1527 2172
rect 1531 2168 1532 2172
rect 1526 2167 1532 2168
rect 1590 2172 1596 2173
rect 1590 2168 1591 2172
rect 1595 2168 1596 2172
rect 1590 2167 1596 2168
rect 1662 2172 1668 2173
rect 1662 2168 1663 2172
rect 1667 2168 1668 2172
rect 1662 2167 1668 2168
rect 1134 2164 1140 2165
rect 1318 2163 1324 2164
rect 1174 2159 1180 2160
rect 1174 2155 1175 2159
rect 1179 2155 1180 2159
rect 1318 2159 1319 2163
rect 1323 2159 1324 2163
rect 1318 2158 1324 2159
rect 111 2154 115 2155
rect 111 2149 115 2150
rect 135 2154 139 2155
rect 135 2149 139 2150
rect 175 2154 179 2155
rect 175 2149 179 2150
rect 215 2154 219 2155
rect 215 2149 219 2150
rect 231 2154 235 2155
rect 231 2149 235 2150
rect 255 2154 259 2155
rect 255 2149 259 2150
rect 271 2154 275 2155
rect 271 2149 275 2150
rect 311 2154 315 2155
rect 311 2149 315 2150
rect 319 2154 323 2155
rect 319 2149 323 2150
rect 359 2154 363 2155
rect 359 2149 363 2150
rect 383 2154 387 2155
rect 383 2149 387 2150
rect 423 2154 427 2155
rect 423 2149 427 2150
rect 447 2154 451 2155
rect 454 2151 455 2155
rect 459 2151 460 2155
rect 454 2150 460 2151
rect 487 2154 491 2155
rect 447 2149 451 2150
rect 487 2149 491 2150
rect 511 2154 515 2155
rect 511 2149 515 2150
rect 559 2154 563 2155
rect 559 2149 563 2150
rect 575 2154 579 2155
rect 575 2149 579 2150
rect 631 2154 635 2155
rect 631 2149 635 2150
rect 639 2154 643 2155
rect 639 2149 643 2150
rect 687 2154 691 2155
rect 687 2149 691 2150
rect 719 2154 723 2155
rect 719 2149 723 2150
rect 735 2154 739 2155
rect 735 2149 739 2150
rect 791 2154 795 2155
rect 791 2149 795 2150
rect 799 2154 803 2155
rect 799 2149 803 2150
rect 847 2154 851 2155
rect 847 2149 851 2150
rect 879 2154 883 2155
rect 879 2149 883 2150
rect 903 2154 907 2155
rect 910 2151 911 2155
rect 915 2151 916 2155
rect 910 2150 916 2151
rect 967 2154 971 2155
rect 903 2149 907 2150
rect 967 2149 971 2150
rect 1095 2154 1099 2155
rect 1174 2154 1180 2155
rect 1186 2155 1192 2156
rect 1095 2149 1099 2150
rect 1134 2152 1140 2153
rect 112 2129 114 2149
rect 232 2137 234 2149
rect 272 2137 274 2149
rect 298 2147 304 2148
rect 298 2143 299 2147
rect 303 2143 304 2147
rect 298 2142 304 2143
rect 230 2136 236 2137
rect 230 2132 231 2136
rect 235 2132 236 2136
rect 230 2131 236 2132
rect 270 2136 276 2137
rect 270 2132 271 2136
rect 275 2132 276 2136
rect 270 2131 276 2132
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 300 2124 302 2142
rect 312 2137 314 2149
rect 338 2147 344 2148
rect 338 2143 339 2147
rect 343 2143 344 2147
rect 338 2142 344 2143
rect 310 2136 316 2137
rect 310 2132 311 2136
rect 315 2132 316 2136
rect 310 2131 316 2132
rect 340 2124 342 2142
rect 360 2137 362 2149
rect 382 2143 388 2144
rect 382 2139 383 2143
rect 387 2139 388 2143
rect 382 2138 388 2139
rect 358 2136 364 2137
rect 358 2132 359 2136
rect 363 2132 364 2136
rect 358 2131 364 2132
rect 384 2124 386 2138
rect 424 2137 426 2149
rect 488 2137 490 2149
rect 560 2137 562 2149
rect 640 2137 642 2149
rect 720 2137 722 2149
rect 726 2147 732 2148
rect 726 2143 727 2147
rect 731 2143 732 2147
rect 726 2142 732 2143
rect 422 2136 428 2137
rect 422 2132 423 2136
rect 427 2132 428 2136
rect 422 2131 428 2132
rect 486 2136 492 2137
rect 486 2132 487 2136
rect 491 2132 492 2136
rect 486 2131 492 2132
rect 558 2136 564 2137
rect 558 2132 559 2136
rect 563 2132 564 2136
rect 558 2131 564 2132
rect 638 2136 644 2137
rect 638 2132 639 2136
rect 643 2132 644 2136
rect 638 2131 644 2132
rect 718 2136 724 2137
rect 718 2132 719 2136
rect 723 2132 724 2136
rect 718 2131 724 2132
rect 110 2123 116 2124
rect 298 2123 304 2124
rect 298 2119 299 2123
rect 303 2119 304 2123
rect 298 2118 304 2119
rect 338 2123 344 2124
rect 338 2119 339 2123
rect 343 2119 344 2123
rect 338 2118 344 2119
rect 382 2123 388 2124
rect 382 2119 383 2123
rect 387 2119 388 2123
rect 382 2118 388 2119
rect 478 2123 484 2124
rect 478 2119 479 2123
rect 483 2119 484 2123
rect 478 2118 484 2119
rect 110 2111 116 2112
rect 110 2107 111 2111
rect 115 2107 116 2111
rect 110 2106 116 2107
rect 230 2108 236 2109
rect 112 2099 114 2106
rect 230 2104 231 2108
rect 235 2104 236 2108
rect 230 2103 236 2104
rect 270 2108 276 2109
rect 270 2104 271 2108
rect 275 2104 276 2108
rect 270 2103 276 2104
rect 310 2108 316 2109
rect 310 2104 311 2108
rect 315 2104 316 2108
rect 310 2103 316 2104
rect 358 2108 364 2109
rect 358 2104 359 2108
rect 363 2104 364 2108
rect 358 2103 364 2104
rect 422 2108 428 2109
rect 422 2104 423 2108
rect 427 2104 428 2108
rect 422 2103 428 2104
rect 232 2099 234 2103
rect 272 2099 274 2103
rect 312 2099 314 2103
rect 360 2099 362 2103
rect 424 2099 426 2103
rect 111 2098 115 2099
rect 111 2093 115 2094
rect 231 2098 235 2099
rect 231 2093 235 2094
rect 271 2098 275 2099
rect 271 2093 275 2094
rect 303 2098 307 2099
rect 303 2093 307 2094
rect 311 2098 315 2099
rect 311 2093 315 2094
rect 351 2098 355 2099
rect 351 2093 355 2094
rect 359 2098 363 2099
rect 359 2093 363 2094
rect 407 2098 411 2099
rect 407 2093 411 2094
rect 423 2098 427 2099
rect 423 2093 427 2094
rect 471 2098 475 2099
rect 471 2093 475 2094
rect 112 2090 114 2093
rect 302 2092 308 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 302 2088 303 2092
rect 307 2088 308 2092
rect 302 2087 308 2088
rect 350 2092 356 2093
rect 350 2088 351 2092
rect 355 2088 356 2092
rect 350 2087 356 2088
rect 406 2092 412 2093
rect 406 2088 407 2092
rect 411 2088 412 2092
rect 406 2087 412 2088
rect 470 2092 476 2093
rect 470 2088 471 2092
rect 475 2088 476 2092
rect 470 2087 476 2088
rect 110 2084 116 2085
rect 286 2075 292 2076
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 286 2071 287 2075
rect 291 2071 292 2075
rect 286 2070 292 2071
rect 398 2075 404 2076
rect 398 2071 399 2075
rect 403 2071 404 2075
rect 398 2070 404 2071
rect 462 2075 468 2076
rect 462 2071 463 2075
rect 467 2071 468 2075
rect 462 2070 468 2071
rect 110 2067 116 2068
rect 112 2043 114 2067
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 183 2042 187 2043
rect 183 2037 187 2038
rect 279 2042 283 2043
rect 279 2037 283 2038
rect 112 2017 114 2037
rect 184 2025 186 2037
rect 254 2035 260 2036
rect 254 2031 255 2035
rect 259 2031 260 2035
rect 254 2030 260 2031
rect 182 2024 188 2025
rect 182 2020 183 2024
rect 187 2020 188 2024
rect 182 2019 188 2020
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 256 2012 258 2030
rect 280 2025 282 2037
rect 288 2036 290 2070
rect 302 2064 308 2065
rect 302 2060 303 2064
rect 307 2060 308 2064
rect 302 2059 308 2060
rect 350 2064 356 2065
rect 350 2060 351 2064
rect 355 2060 356 2064
rect 350 2059 356 2060
rect 304 2043 306 2059
rect 352 2043 354 2059
rect 400 2052 402 2070
rect 406 2064 412 2065
rect 406 2060 407 2064
rect 411 2060 412 2064
rect 406 2059 412 2060
rect 390 2051 396 2052
rect 390 2047 391 2051
rect 395 2047 396 2051
rect 390 2046 396 2047
rect 398 2051 404 2052
rect 398 2047 399 2051
rect 403 2047 404 2051
rect 398 2046 404 2047
rect 303 2042 307 2043
rect 303 2037 307 2038
rect 351 2042 355 2043
rect 351 2037 355 2038
rect 375 2042 379 2043
rect 375 2037 379 2038
rect 286 2035 292 2036
rect 286 2031 287 2035
rect 291 2031 292 2035
rect 286 2030 292 2031
rect 376 2025 378 2037
rect 278 2024 284 2025
rect 278 2020 279 2024
rect 283 2020 284 2024
rect 278 2019 284 2020
rect 374 2024 380 2025
rect 374 2020 375 2024
rect 379 2020 380 2024
rect 374 2019 380 2020
rect 392 2012 394 2046
rect 408 2043 410 2059
rect 464 2052 466 2070
rect 470 2064 476 2065
rect 470 2060 471 2064
rect 475 2060 476 2064
rect 470 2059 476 2060
rect 462 2051 468 2052
rect 462 2047 463 2051
rect 467 2047 468 2051
rect 462 2046 468 2047
rect 472 2043 474 2059
rect 480 2044 482 2118
rect 486 2108 492 2109
rect 486 2104 487 2108
rect 491 2104 492 2108
rect 486 2103 492 2104
rect 558 2108 564 2109
rect 558 2104 559 2108
rect 563 2104 564 2108
rect 558 2103 564 2104
rect 638 2108 644 2109
rect 638 2104 639 2108
rect 643 2104 644 2108
rect 638 2103 644 2104
rect 718 2108 724 2109
rect 718 2104 719 2108
rect 723 2104 724 2108
rect 718 2103 724 2104
rect 488 2099 490 2103
rect 560 2099 562 2103
rect 640 2099 642 2103
rect 720 2099 722 2103
rect 487 2098 491 2099
rect 487 2093 491 2094
rect 543 2098 547 2099
rect 543 2093 547 2094
rect 559 2098 563 2099
rect 559 2093 563 2094
rect 623 2098 627 2099
rect 623 2093 627 2094
rect 639 2098 643 2099
rect 639 2093 643 2094
rect 703 2098 707 2099
rect 703 2093 707 2094
rect 719 2098 723 2099
rect 719 2093 723 2094
rect 542 2092 548 2093
rect 542 2088 543 2092
rect 547 2088 548 2092
rect 542 2087 548 2088
rect 622 2092 628 2093
rect 622 2088 623 2092
rect 627 2088 628 2092
rect 622 2087 628 2088
rect 702 2092 708 2093
rect 702 2088 703 2092
rect 707 2088 708 2092
rect 702 2087 708 2088
rect 728 2076 730 2142
rect 800 2137 802 2149
rect 826 2147 832 2148
rect 826 2143 827 2147
rect 831 2143 832 2147
rect 826 2142 832 2143
rect 798 2136 804 2137
rect 798 2132 799 2136
rect 803 2132 804 2136
rect 798 2131 804 2132
rect 828 2124 830 2142
rect 880 2137 882 2149
rect 968 2137 970 2149
rect 878 2136 884 2137
rect 878 2132 879 2136
rect 883 2132 884 2136
rect 878 2131 884 2132
rect 966 2136 972 2137
rect 966 2132 967 2136
rect 971 2132 972 2136
rect 966 2131 972 2132
rect 1096 2129 1098 2149
rect 1134 2148 1135 2152
rect 1139 2148 1140 2152
rect 1134 2147 1140 2148
rect 1094 2128 1100 2129
rect 1094 2124 1095 2128
rect 1099 2124 1100 2128
rect 1136 2127 1138 2147
rect 1158 2144 1164 2145
rect 1158 2140 1159 2144
rect 1163 2140 1164 2144
rect 1158 2139 1164 2140
rect 1160 2127 1162 2139
rect 1176 2132 1178 2154
rect 1186 2151 1187 2155
rect 1191 2151 1192 2155
rect 1186 2150 1192 2151
rect 1226 2155 1232 2156
rect 1226 2151 1227 2155
rect 1231 2151 1232 2155
rect 1226 2150 1232 2151
rect 1266 2155 1272 2156
rect 1266 2151 1267 2155
rect 1271 2151 1272 2155
rect 1266 2150 1272 2151
rect 1188 2132 1190 2150
rect 1198 2144 1204 2145
rect 1198 2140 1199 2144
rect 1203 2140 1204 2144
rect 1198 2139 1204 2140
rect 1174 2131 1180 2132
rect 1174 2127 1175 2131
rect 1179 2127 1180 2131
rect 826 2123 832 2124
rect 826 2119 827 2123
rect 831 2119 832 2123
rect 826 2118 832 2119
rect 1030 2123 1036 2124
rect 1094 2123 1100 2124
rect 1135 2126 1139 2127
rect 1030 2119 1031 2123
rect 1035 2119 1036 2123
rect 1135 2121 1139 2122
rect 1159 2126 1163 2127
rect 1174 2126 1180 2127
rect 1186 2131 1192 2132
rect 1186 2127 1187 2131
rect 1191 2127 1192 2131
rect 1200 2127 1202 2139
rect 1228 2132 1230 2150
rect 1238 2144 1244 2145
rect 1238 2140 1239 2144
rect 1243 2140 1244 2144
rect 1238 2139 1244 2140
rect 1226 2131 1232 2132
rect 1226 2127 1227 2131
rect 1231 2127 1232 2131
rect 1240 2127 1242 2139
rect 1268 2132 1270 2150
rect 1278 2144 1284 2145
rect 1278 2140 1279 2144
rect 1283 2140 1284 2144
rect 1278 2139 1284 2140
rect 1266 2131 1272 2132
rect 1266 2127 1267 2131
rect 1271 2127 1272 2131
rect 1280 2127 1282 2139
rect 1186 2126 1192 2127
rect 1199 2126 1203 2127
rect 1226 2126 1232 2127
rect 1239 2126 1243 2127
rect 1266 2126 1272 2127
rect 1279 2126 1283 2127
rect 1159 2121 1163 2122
rect 1199 2121 1203 2122
rect 1239 2121 1243 2122
rect 1279 2121 1283 2122
rect 1295 2126 1299 2127
rect 1295 2121 1299 2122
rect 1030 2118 1036 2119
rect 798 2108 804 2109
rect 798 2104 799 2108
rect 803 2104 804 2108
rect 798 2103 804 2104
rect 878 2108 884 2109
rect 878 2104 879 2108
rect 883 2104 884 2108
rect 878 2103 884 2104
rect 966 2108 972 2109
rect 966 2104 967 2108
rect 971 2104 972 2108
rect 966 2103 972 2104
rect 800 2099 802 2103
rect 880 2099 882 2103
rect 968 2099 970 2103
rect 783 2098 787 2099
rect 783 2093 787 2094
rect 799 2098 803 2099
rect 799 2093 803 2094
rect 863 2098 867 2099
rect 863 2093 867 2094
rect 879 2098 883 2099
rect 879 2093 883 2094
rect 951 2098 955 2099
rect 951 2093 955 2094
rect 967 2098 971 2099
rect 967 2093 971 2094
rect 782 2092 788 2093
rect 782 2088 783 2092
rect 787 2088 788 2092
rect 782 2087 788 2088
rect 862 2092 868 2093
rect 862 2088 863 2092
rect 867 2088 868 2092
rect 862 2087 868 2088
rect 950 2092 956 2093
rect 950 2088 951 2092
rect 955 2088 956 2092
rect 950 2087 956 2088
rect 534 2075 540 2076
rect 534 2071 535 2075
rect 539 2071 540 2075
rect 534 2070 540 2071
rect 614 2075 620 2076
rect 614 2071 615 2075
rect 619 2071 620 2075
rect 614 2070 620 2071
rect 630 2075 636 2076
rect 630 2071 631 2075
rect 635 2071 636 2075
rect 630 2070 636 2071
rect 726 2075 732 2076
rect 726 2071 727 2075
rect 731 2071 732 2075
rect 726 2070 732 2071
rect 822 2075 828 2076
rect 822 2071 823 2075
rect 827 2071 828 2075
rect 822 2070 828 2071
rect 536 2052 538 2070
rect 542 2064 548 2065
rect 542 2060 543 2064
rect 547 2060 548 2064
rect 542 2059 548 2060
rect 534 2051 540 2052
rect 534 2047 535 2051
rect 539 2047 540 2051
rect 534 2046 540 2047
rect 478 2043 484 2044
rect 544 2043 546 2059
rect 616 2052 618 2070
rect 622 2064 628 2065
rect 622 2060 623 2064
rect 627 2060 628 2064
rect 622 2059 628 2060
rect 614 2051 620 2052
rect 614 2047 615 2051
rect 619 2047 620 2051
rect 614 2046 620 2047
rect 624 2043 626 2059
rect 632 2044 634 2070
rect 702 2064 708 2065
rect 702 2060 703 2064
rect 707 2060 708 2064
rect 702 2059 708 2060
rect 782 2064 788 2065
rect 782 2060 783 2064
rect 787 2060 788 2064
rect 782 2059 788 2060
rect 630 2043 636 2044
rect 704 2043 706 2059
rect 774 2051 780 2052
rect 774 2047 775 2051
rect 779 2047 780 2051
rect 774 2046 780 2047
rect 407 2042 411 2043
rect 407 2037 411 2038
rect 463 2042 467 2043
rect 463 2037 467 2038
rect 471 2042 475 2043
rect 478 2039 479 2043
rect 483 2039 484 2043
rect 478 2038 484 2039
rect 543 2042 547 2043
rect 471 2037 475 2038
rect 543 2037 547 2038
rect 623 2042 627 2043
rect 630 2039 631 2043
rect 635 2039 636 2043
rect 630 2038 636 2039
rect 695 2042 699 2043
rect 623 2037 627 2038
rect 695 2037 699 2038
rect 703 2042 707 2043
rect 703 2037 707 2038
rect 759 2042 763 2043
rect 759 2037 763 2038
rect 398 2035 404 2036
rect 398 2031 399 2035
rect 403 2031 404 2035
rect 398 2030 404 2031
rect 110 2011 116 2012
rect 166 2011 172 2012
rect 166 2007 167 2011
rect 171 2007 172 2011
rect 166 2006 172 2007
rect 254 2011 260 2012
rect 254 2007 255 2011
rect 259 2007 260 2011
rect 254 2006 260 2007
rect 390 2011 396 2012
rect 390 2007 391 2011
rect 395 2007 396 2011
rect 390 2006 396 2007
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 112 1991 114 1994
rect 111 1990 115 1991
rect 111 1985 115 1986
rect 159 1990 163 1991
rect 159 1985 163 1986
rect 112 1982 114 1985
rect 158 1984 164 1985
rect 110 1981 116 1982
rect 110 1977 111 1981
rect 115 1977 116 1981
rect 158 1980 159 1984
rect 163 1980 164 1984
rect 158 1979 164 1980
rect 110 1976 116 1977
rect 110 1964 116 1965
rect 110 1960 111 1964
rect 115 1960 116 1964
rect 110 1959 116 1960
rect 112 1935 114 1959
rect 158 1956 164 1957
rect 158 1952 159 1956
rect 163 1952 164 1956
rect 158 1951 164 1952
rect 160 1935 162 1951
rect 168 1944 170 2006
rect 182 1996 188 1997
rect 182 1992 183 1996
rect 187 1992 188 1996
rect 182 1991 188 1992
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 374 1996 380 1997
rect 374 1992 375 1996
rect 379 1992 380 1996
rect 374 1991 380 1992
rect 183 1990 187 1991
rect 183 1985 187 1986
rect 231 1990 235 1991
rect 231 1985 235 1986
rect 279 1990 283 1991
rect 279 1985 283 1986
rect 303 1990 307 1991
rect 303 1985 307 1986
rect 375 1990 379 1991
rect 375 1985 379 1986
rect 230 1984 236 1985
rect 230 1980 231 1984
rect 235 1980 236 1984
rect 230 1979 236 1980
rect 302 1984 308 1985
rect 302 1980 303 1984
rect 307 1980 308 1984
rect 302 1979 308 1980
rect 374 1984 380 1985
rect 374 1980 375 1984
rect 379 1980 380 1984
rect 374 1979 380 1980
rect 400 1968 402 2030
rect 464 2025 466 2037
rect 530 2035 536 2036
rect 530 2031 531 2035
rect 535 2031 536 2035
rect 530 2030 536 2031
rect 462 2024 468 2025
rect 462 2020 463 2024
rect 467 2020 468 2024
rect 462 2019 468 2020
rect 532 2012 534 2030
rect 544 2025 546 2037
rect 624 2025 626 2037
rect 642 2035 648 2036
rect 642 2031 643 2035
rect 647 2031 648 2035
rect 642 2030 648 2031
rect 650 2035 656 2036
rect 650 2031 651 2035
rect 655 2031 656 2035
rect 650 2030 656 2031
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 622 2024 628 2025
rect 622 2020 623 2024
rect 627 2020 628 2024
rect 622 2019 628 2020
rect 454 2011 460 2012
rect 454 2007 455 2011
rect 459 2007 460 2011
rect 454 2006 460 2007
rect 530 2011 536 2012
rect 530 2007 531 2011
rect 535 2007 536 2011
rect 530 2006 536 2007
rect 447 1990 451 1991
rect 447 1985 451 1986
rect 446 1984 452 1985
rect 446 1980 447 1984
rect 451 1980 452 1984
rect 446 1979 452 1980
rect 182 1967 188 1968
rect 182 1963 183 1967
rect 187 1963 188 1967
rect 182 1962 188 1963
rect 294 1967 300 1968
rect 294 1963 295 1967
rect 299 1963 300 1967
rect 294 1962 300 1963
rect 366 1967 372 1968
rect 366 1963 367 1967
rect 371 1963 372 1967
rect 366 1962 372 1963
rect 398 1967 404 1968
rect 398 1963 399 1967
rect 403 1963 404 1967
rect 398 1962 404 1963
rect 166 1943 172 1944
rect 166 1939 167 1943
rect 171 1939 172 1943
rect 166 1938 172 1939
rect 111 1934 115 1935
rect 111 1929 115 1930
rect 135 1934 139 1935
rect 135 1929 139 1930
rect 159 1934 163 1935
rect 159 1929 163 1930
rect 175 1934 179 1935
rect 175 1929 179 1930
rect 112 1909 114 1929
rect 136 1917 138 1929
rect 176 1917 178 1929
rect 184 1928 186 1962
rect 230 1956 236 1957
rect 230 1952 231 1956
rect 235 1952 236 1956
rect 230 1951 236 1952
rect 198 1935 204 1936
rect 232 1935 234 1951
rect 296 1944 298 1962
rect 302 1956 308 1957
rect 302 1952 303 1956
rect 307 1952 308 1956
rect 302 1951 308 1952
rect 294 1943 300 1944
rect 294 1939 295 1943
rect 299 1939 300 1943
rect 294 1938 300 1939
rect 304 1935 306 1951
rect 368 1944 370 1962
rect 374 1956 380 1957
rect 374 1952 375 1956
rect 379 1952 380 1956
rect 374 1951 380 1952
rect 446 1956 452 1957
rect 446 1952 447 1956
rect 451 1952 452 1956
rect 446 1951 452 1952
rect 366 1943 372 1944
rect 366 1939 367 1943
rect 371 1939 372 1943
rect 366 1938 372 1939
rect 376 1935 378 1951
rect 448 1935 450 1951
rect 456 1944 458 2006
rect 462 1996 468 1997
rect 462 1992 463 1996
rect 467 1992 468 1996
rect 462 1991 468 1992
rect 542 1996 548 1997
rect 542 1992 543 1996
rect 547 1992 548 1996
rect 542 1991 548 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 463 1990 467 1991
rect 463 1985 467 1986
rect 527 1990 531 1991
rect 527 1985 531 1986
rect 543 1990 547 1991
rect 543 1985 547 1986
rect 607 1990 611 1991
rect 607 1985 611 1986
rect 623 1990 627 1991
rect 623 1985 627 1986
rect 526 1984 532 1985
rect 526 1980 527 1984
rect 531 1980 532 1984
rect 526 1979 532 1980
rect 606 1984 612 1985
rect 606 1980 607 1984
rect 611 1980 612 1984
rect 606 1979 612 1980
rect 644 1976 646 2030
rect 652 2012 654 2030
rect 696 2025 698 2037
rect 722 2035 728 2036
rect 722 2031 723 2035
rect 727 2031 728 2035
rect 722 2030 728 2031
rect 694 2024 700 2025
rect 694 2020 695 2024
rect 699 2020 700 2024
rect 694 2019 700 2020
rect 724 2012 726 2030
rect 760 2025 762 2037
rect 758 2024 764 2025
rect 758 2020 759 2024
rect 763 2020 764 2024
rect 758 2019 764 2020
rect 776 2012 778 2046
rect 784 2043 786 2059
rect 783 2042 787 2043
rect 783 2037 787 2038
rect 815 2042 819 2043
rect 815 2037 819 2038
rect 816 2025 818 2037
rect 824 2036 826 2070
rect 862 2064 868 2065
rect 862 2060 863 2064
rect 867 2060 868 2064
rect 862 2059 868 2060
rect 950 2064 956 2065
rect 950 2060 951 2064
rect 955 2060 956 2064
rect 950 2059 956 2060
rect 864 2043 866 2059
rect 952 2043 954 2059
rect 1032 2052 1034 2118
rect 1094 2111 1100 2112
rect 1094 2107 1095 2111
rect 1099 2107 1100 2111
rect 1094 2106 1100 2107
rect 1096 2099 1098 2106
rect 1136 2101 1138 2121
rect 1160 2109 1162 2121
rect 1178 2119 1184 2120
rect 1178 2115 1179 2119
rect 1183 2115 1184 2119
rect 1178 2114 1184 2115
rect 1186 2119 1192 2120
rect 1186 2115 1187 2119
rect 1191 2115 1192 2119
rect 1186 2114 1192 2115
rect 1158 2108 1164 2109
rect 1158 2104 1159 2108
rect 1163 2104 1164 2108
rect 1158 2103 1164 2104
rect 1134 2100 1140 2101
rect 1039 2098 1043 2099
rect 1039 2093 1043 2094
rect 1095 2098 1099 2099
rect 1134 2096 1135 2100
rect 1139 2096 1140 2100
rect 1134 2095 1140 2096
rect 1095 2093 1099 2094
rect 1038 2092 1044 2093
rect 1038 2088 1039 2092
rect 1043 2088 1044 2092
rect 1096 2090 1098 2093
rect 1038 2087 1044 2088
rect 1094 2089 1100 2090
rect 1094 2085 1095 2089
rect 1099 2085 1100 2089
rect 1094 2084 1100 2085
rect 1134 2083 1140 2084
rect 1134 2079 1135 2083
rect 1139 2079 1140 2083
rect 1134 2078 1140 2079
rect 1158 2080 1164 2081
rect 1136 2075 1138 2078
rect 1158 2076 1159 2080
rect 1163 2076 1164 2080
rect 1158 2075 1164 2076
rect 1135 2074 1139 2075
rect 1094 2072 1100 2073
rect 1094 2068 1095 2072
rect 1099 2068 1100 2072
rect 1135 2069 1139 2070
rect 1159 2074 1163 2075
rect 1159 2069 1163 2070
rect 1094 2067 1100 2068
rect 1038 2064 1044 2065
rect 1038 2060 1039 2064
rect 1043 2060 1044 2064
rect 1038 2059 1044 2060
rect 1030 2051 1036 2052
rect 1030 2047 1031 2051
rect 1035 2047 1036 2051
rect 1030 2046 1036 2047
rect 1040 2043 1042 2059
rect 1096 2043 1098 2067
rect 1136 2066 1138 2069
rect 1158 2068 1164 2069
rect 1134 2065 1140 2066
rect 1134 2061 1135 2065
rect 1139 2061 1140 2065
rect 1158 2064 1159 2068
rect 1163 2064 1164 2068
rect 1158 2063 1164 2064
rect 1134 2060 1140 2061
rect 1180 2052 1182 2114
rect 1188 2096 1190 2114
rect 1200 2109 1202 2121
rect 1226 2119 1232 2120
rect 1226 2115 1227 2119
rect 1231 2115 1232 2119
rect 1226 2114 1232 2115
rect 1198 2108 1204 2109
rect 1198 2104 1199 2108
rect 1203 2104 1204 2108
rect 1198 2103 1204 2104
rect 1228 2096 1230 2114
rect 1240 2109 1242 2121
rect 1266 2119 1272 2120
rect 1266 2115 1267 2119
rect 1271 2115 1272 2119
rect 1266 2114 1272 2115
rect 1238 2108 1244 2109
rect 1238 2104 1239 2108
rect 1243 2104 1244 2108
rect 1238 2103 1244 2104
rect 1268 2096 1270 2114
rect 1296 2109 1298 2121
rect 1294 2108 1300 2109
rect 1294 2104 1295 2108
rect 1299 2104 1300 2108
rect 1294 2103 1300 2104
rect 1320 2096 1322 2158
rect 1680 2156 1682 2218
rect 1688 2213 1690 2225
rect 1714 2223 1720 2224
rect 1714 2219 1715 2223
rect 1719 2219 1720 2223
rect 1714 2218 1720 2219
rect 1686 2212 1692 2213
rect 1686 2208 1687 2212
rect 1691 2208 1692 2212
rect 1686 2207 1692 2208
rect 1716 2200 1718 2218
rect 1728 2213 1730 2225
rect 1750 2223 1756 2224
rect 1750 2219 1751 2223
rect 1755 2219 1756 2223
rect 1750 2218 1756 2219
rect 1726 2212 1732 2213
rect 1726 2208 1727 2212
rect 1731 2208 1732 2212
rect 1726 2207 1732 2208
rect 1752 2200 1754 2218
rect 1768 2213 1770 2225
rect 1794 2223 1800 2224
rect 1794 2219 1795 2223
rect 1799 2219 1800 2223
rect 1794 2218 1800 2219
rect 1766 2212 1772 2213
rect 1766 2208 1767 2212
rect 1771 2208 1772 2212
rect 1766 2207 1772 2208
rect 1796 2200 1798 2218
rect 1808 2213 1810 2225
rect 1806 2212 1812 2213
rect 1806 2208 1807 2212
rect 1811 2208 1812 2212
rect 1806 2207 1812 2208
rect 2120 2205 2122 2225
rect 2118 2204 2124 2205
rect 2118 2200 2119 2204
rect 2123 2200 2124 2204
rect 1714 2199 1720 2200
rect 1714 2195 1715 2199
rect 1719 2195 1720 2199
rect 1714 2194 1720 2195
rect 1750 2199 1756 2200
rect 1750 2195 1751 2199
rect 1755 2195 1756 2199
rect 1750 2194 1756 2195
rect 1794 2199 1800 2200
rect 1794 2195 1795 2199
rect 1799 2195 1800 2199
rect 1794 2194 1800 2195
rect 1814 2199 1820 2200
rect 2118 2199 2124 2200
rect 1814 2195 1815 2199
rect 1819 2195 1820 2199
rect 1814 2194 1820 2195
rect 1686 2184 1692 2185
rect 1686 2180 1687 2184
rect 1691 2180 1692 2184
rect 1686 2179 1692 2180
rect 1726 2184 1732 2185
rect 1726 2180 1727 2184
rect 1731 2180 1732 2184
rect 1726 2179 1732 2180
rect 1766 2184 1772 2185
rect 1766 2180 1767 2184
rect 1771 2180 1772 2184
rect 1766 2179 1772 2180
rect 1806 2184 1812 2185
rect 1806 2180 1807 2184
rect 1811 2180 1812 2184
rect 1806 2179 1812 2180
rect 1687 2178 1691 2179
rect 1687 2173 1691 2174
rect 1727 2178 1731 2179
rect 1727 2173 1731 2174
rect 1735 2178 1739 2179
rect 1735 2173 1739 2174
rect 1767 2178 1771 2179
rect 1767 2173 1771 2174
rect 1807 2178 1811 2179
rect 1807 2173 1811 2174
rect 1734 2172 1740 2173
rect 1734 2168 1735 2172
rect 1739 2168 1740 2172
rect 1734 2167 1740 2168
rect 1806 2172 1812 2173
rect 1806 2168 1807 2172
rect 1811 2168 1812 2172
rect 1806 2167 1812 2168
rect 1766 2163 1772 2164
rect 1766 2159 1767 2163
rect 1771 2159 1772 2163
rect 1766 2158 1772 2159
rect 1326 2155 1332 2156
rect 1326 2151 1327 2155
rect 1331 2151 1332 2155
rect 1326 2150 1332 2151
rect 1382 2155 1388 2156
rect 1382 2151 1383 2155
rect 1387 2151 1388 2155
rect 1382 2150 1388 2151
rect 1446 2155 1452 2156
rect 1446 2151 1447 2155
rect 1451 2151 1452 2155
rect 1446 2150 1452 2151
rect 1498 2155 1504 2156
rect 1498 2151 1499 2155
rect 1503 2151 1504 2155
rect 1498 2150 1504 2151
rect 1534 2155 1540 2156
rect 1534 2151 1535 2155
rect 1539 2151 1540 2155
rect 1534 2150 1540 2151
rect 1654 2155 1660 2156
rect 1654 2151 1655 2155
rect 1659 2151 1660 2155
rect 1654 2150 1660 2151
rect 1678 2155 1684 2156
rect 1678 2151 1679 2155
rect 1683 2151 1684 2155
rect 1678 2150 1684 2151
rect 1758 2155 1764 2156
rect 1758 2151 1759 2155
rect 1763 2151 1764 2155
rect 1758 2150 1764 2151
rect 1328 2132 1330 2150
rect 1334 2144 1340 2145
rect 1334 2140 1335 2144
rect 1339 2140 1340 2144
rect 1334 2139 1340 2140
rect 1326 2131 1332 2132
rect 1326 2127 1327 2131
rect 1331 2127 1332 2131
rect 1336 2127 1338 2139
rect 1384 2132 1386 2150
rect 1390 2144 1396 2145
rect 1390 2140 1391 2144
rect 1395 2140 1396 2144
rect 1390 2139 1396 2140
rect 1382 2131 1388 2132
rect 1382 2127 1383 2131
rect 1387 2127 1388 2131
rect 1392 2127 1394 2139
rect 1448 2132 1450 2150
rect 1454 2144 1460 2145
rect 1454 2140 1455 2144
rect 1459 2140 1460 2144
rect 1454 2139 1460 2140
rect 1446 2131 1452 2132
rect 1446 2127 1447 2131
rect 1451 2127 1452 2131
rect 1456 2127 1458 2139
rect 1500 2132 1502 2150
rect 1526 2144 1532 2145
rect 1526 2140 1527 2144
rect 1531 2140 1532 2144
rect 1526 2139 1532 2140
rect 1498 2131 1504 2132
rect 1498 2127 1499 2131
rect 1503 2127 1504 2131
rect 1528 2127 1530 2139
rect 1326 2126 1332 2127
rect 1335 2126 1339 2127
rect 1335 2121 1339 2122
rect 1367 2126 1371 2127
rect 1382 2126 1388 2127
rect 1391 2126 1395 2127
rect 1367 2121 1371 2122
rect 1391 2121 1395 2122
rect 1439 2126 1443 2127
rect 1446 2126 1452 2127
rect 1455 2126 1459 2127
rect 1498 2126 1504 2127
rect 1519 2126 1523 2127
rect 1439 2121 1443 2122
rect 1455 2121 1459 2122
rect 1519 2121 1523 2122
rect 1527 2126 1531 2127
rect 1527 2121 1531 2122
rect 1368 2109 1370 2121
rect 1402 2119 1408 2120
rect 1402 2115 1403 2119
rect 1407 2115 1408 2119
rect 1402 2114 1408 2115
rect 1366 2108 1372 2109
rect 1366 2104 1367 2108
rect 1371 2104 1372 2108
rect 1366 2103 1372 2104
rect 1404 2096 1406 2114
rect 1440 2109 1442 2121
rect 1520 2109 1522 2121
rect 1536 2120 1538 2150
rect 1590 2144 1596 2145
rect 1590 2140 1591 2144
rect 1595 2140 1596 2144
rect 1590 2139 1596 2140
rect 1592 2127 1594 2139
rect 1656 2132 1658 2150
rect 1662 2144 1668 2145
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1734 2144 1740 2145
rect 1734 2140 1735 2144
rect 1739 2140 1740 2144
rect 1734 2139 1740 2140
rect 1646 2131 1652 2132
rect 1646 2127 1647 2131
rect 1651 2127 1652 2131
rect 1591 2126 1595 2127
rect 1591 2121 1595 2122
rect 1599 2126 1603 2127
rect 1646 2126 1652 2127
rect 1654 2131 1660 2132
rect 1654 2127 1655 2131
rect 1659 2127 1660 2131
rect 1664 2127 1666 2139
rect 1736 2127 1738 2139
rect 1654 2126 1660 2127
rect 1663 2126 1667 2127
rect 1599 2121 1603 2122
rect 1534 2119 1540 2120
rect 1534 2115 1535 2119
rect 1539 2115 1540 2119
rect 1534 2114 1540 2115
rect 1600 2109 1602 2121
rect 1614 2119 1620 2120
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1626 2119 1632 2120
rect 1626 2115 1627 2119
rect 1631 2115 1632 2119
rect 1626 2114 1632 2115
rect 1438 2108 1444 2109
rect 1438 2104 1439 2108
rect 1443 2104 1444 2108
rect 1438 2103 1444 2104
rect 1518 2108 1524 2109
rect 1518 2104 1519 2108
rect 1523 2104 1524 2108
rect 1518 2103 1524 2104
rect 1598 2108 1604 2109
rect 1598 2104 1599 2108
rect 1603 2104 1604 2108
rect 1598 2103 1604 2104
rect 1186 2095 1192 2096
rect 1186 2091 1187 2095
rect 1191 2091 1192 2095
rect 1186 2090 1192 2091
rect 1226 2095 1232 2096
rect 1226 2091 1227 2095
rect 1231 2091 1232 2095
rect 1226 2090 1232 2091
rect 1266 2095 1272 2096
rect 1266 2091 1267 2095
rect 1271 2091 1272 2095
rect 1266 2090 1272 2091
rect 1318 2095 1324 2096
rect 1318 2091 1319 2095
rect 1323 2091 1324 2095
rect 1318 2090 1324 2091
rect 1402 2095 1408 2096
rect 1402 2091 1403 2095
rect 1407 2091 1408 2095
rect 1402 2090 1408 2091
rect 1486 2095 1492 2096
rect 1486 2091 1487 2095
rect 1491 2091 1492 2095
rect 1486 2090 1492 2091
rect 1198 2080 1204 2081
rect 1198 2076 1199 2080
rect 1203 2076 1204 2080
rect 1198 2075 1204 2076
rect 1238 2080 1244 2081
rect 1238 2076 1239 2080
rect 1243 2076 1244 2080
rect 1238 2075 1244 2076
rect 1294 2080 1300 2081
rect 1294 2076 1295 2080
rect 1299 2076 1300 2080
rect 1294 2075 1300 2076
rect 1366 2080 1372 2081
rect 1366 2076 1367 2080
rect 1371 2076 1372 2080
rect 1366 2075 1372 2076
rect 1438 2080 1444 2081
rect 1438 2076 1439 2080
rect 1443 2076 1444 2080
rect 1438 2075 1444 2076
rect 1199 2074 1203 2075
rect 1199 2069 1203 2070
rect 1215 2074 1219 2075
rect 1215 2069 1219 2070
rect 1239 2074 1243 2075
rect 1239 2069 1243 2070
rect 1295 2074 1299 2075
rect 1295 2069 1299 2070
rect 1303 2074 1307 2075
rect 1303 2069 1307 2070
rect 1367 2074 1371 2075
rect 1367 2069 1371 2070
rect 1399 2074 1403 2075
rect 1399 2069 1403 2070
rect 1439 2074 1443 2075
rect 1439 2069 1443 2070
rect 1214 2068 1220 2069
rect 1214 2064 1215 2068
rect 1219 2064 1220 2068
rect 1214 2063 1220 2064
rect 1302 2068 1308 2069
rect 1302 2064 1303 2068
rect 1307 2064 1308 2068
rect 1302 2063 1308 2064
rect 1398 2068 1404 2069
rect 1398 2064 1399 2068
rect 1403 2064 1404 2068
rect 1398 2063 1404 2064
rect 1178 2051 1184 2052
rect 1134 2048 1140 2049
rect 1134 2044 1135 2048
rect 1139 2044 1140 2048
rect 1178 2047 1179 2051
rect 1183 2047 1184 2051
rect 1178 2046 1184 2047
rect 1358 2051 1364 2052
rect 1358 2047 1359 2051
rect 1363 2047 1364 2051
rect 1358 2046 1364 2047
rect 1134 2043 1140 2044
rect 863 2042 867 2043
rect 863 2037 867 2038
rect 911 2042 915 2043
rect 911 2037 915 2038
rect 951 2042 955 2043
rect 951 2037 955 2038
rect 959 2042 963 2043
rect 959 2037 963 2038
rect 1007 2042 1011 2043
rect 1007 2037 1011 2038
rect 1039 2042 1043 2043
rect 1039 2037 1043 2038
rect 1047 2042 1051 2043
rect 1047 2037 1051 2038
rect 1095 2042 1099 2043
rect 1095 2037 1099 2038
rect 822 2035 828 2036
rect 822 2031 823 2035
rect 827 2031 828 2035
rect 822 2030 828 2031
rect 842 2035 848 2036
rect 842 2031 843 2035
rect 847 2031 848 2035
rect 842 2030 848 2031
rect 814 2024 820 2025
rect 814 2020 815 2024
rect 819 2020 820 2024
rect 814 2019 820 2020
rect 844 2012 846 2030
rect 864 2025 866 2037
rect 890 2035 896 2036
rect 890 2031 891 2035
rect 895 2031 896 2035
rect 890 2030 896 2031
rect 862 2024 868 2025
rect 862 2020 863 2024
rect 867 2020 868 2024
rect 862 2019 868 2020
rect 892 2012 894 2030
rect 912 2025 914 2037
rect 938 2035 944 2036
rect 938 2031 939 2035
rect 943 2031 944 2035
rect 938 2030 944 2031
rect 910 2024 916 2025
rect 910 2020 911 2024
rect 915 2020 916 2024
rect 910 2019 916 2020
rect 940 2012 942 2030
rect 960 2025 962 2037
rect 986 2035 992 2036
rect 986 2031 987 2035
rect 991 2031 992 2035
rect 986 2030 992 2031
rect 958 2024 964 2025
rect 958 2020 959 2024
rect 963 2020 964 2024
rect 958 2019 964 2020
rect 988 2012 990 2030
rect 1008 2025 1010 2037
rect 1030 2035 1036 2036
rect 1030 2031 1031 2035
rect 1035 2031 1036 2035
rect 1030 2030 1036 2031
rect 1006 2024 1012 2025
rect 1006 2020 1007 2024
rect 1011 2020 1012 2024
rect 1006 2019 1012 2020
rect 1032 2012 1034 2030
rect 1048 2025 1050 2037
rect 1046 2024 1052 2025
rect 1046 2020 1047 2024
rect 1051 2020 1052 2024
rect 1046 2019 1052 2020
rect 1096 2017 1098 2037
rect 1136 2023 1138 2043
rect 1158 2040 1164 2041
rect 1158 2036 1159 2040
rect 1163 2036 1164 2040
rect 1158 2035 1164 2036
rect 1214 2040 1220 2041
rect 1214 2036 1215 2040
rect 1219 2036 1220 2040
rect 1214 2035 1220 2036
rect 1302 2040 1308 2041
rect 1302 2036 1303 2040
rect 1307 2036 1308 2040
rect 1302 2035 1308 2036
rect 1160 2023 1162 2035
rect 1216 2023 1218 2035
rect 1266 2027 1272 2028
rect 1266 2023 1267 2027
rect 1271 2023 1272 2027
rect 1304 2023 1306 2035
rect 1135 2022 1139 2023
rect 1135 2017 1139 2018
rect 1159 2022 1163 2023
rect 1159 2017 1163 2018
rect 1215 2022 1219 2023
rect 1215 2017 1219 2018
rect 1239 2022 1243 2023
rect 1266 2022 1272 2023
rect 1303 2022 1307 2023
rect 1239 2017 1243 2018
rect 1094 2016 1100 2017
rect 1094 2012 1095 2016
rect 1099 2012 1100 2016
rect 650 2011 656 2012
rect 650 2007 651 2011
rect 655 2007 656 2011
rect 650 2006 656 2007
rect 722 2011 728 2012
rect 722 2007 723 2011
rect 727 2007 728 2011
rect 722 2006 728 2007
rect 774 2011 780 2012
rect 774 2007 775 2011
rect 779 2007 780 2011
rect 774 2006 780 2007
rect 842 2011 848 2012
rect 842 2007 843 2011
rect 847 2007 848 2011
rect 842 2006 848 2007
rect 890 2011 896 2012
rect 890 2007 891 2011
rect 895 2007 896 2011
rect 890 2006 896 2007
rect 938 2011 944 2012
rect 938 2007 939 2011
rect 943 2007 944 2011
rect 938 2006 944 2007
rect 986 2011 992 2012
rect 986 2007 987 2011
rect 991 2007 992 2011
rect 986 2006 992 2007
rect 1030 2011 1036 2012
rect 1094 2011 1100 2012
rect 1030 2007 1031 2011
rect 1035 2007 1036 2011
rect 1030 2006 1036 2007
rect 1094 1999 1100 2000
rect 694 1996 700 1997
rect 694 1992 695 1996
rect 699 1992 700 1996
rect 694 1991 700 1992
rect 758 1996 764 1997
rect 758 1992 759 1996
rect 763 1992 764 1996
rect 758 1991 764 1992
rect 814 1996 820 1997
rect 814 1992 815 1996
rect 819 1992 820 1996
rect 814 1991 820 1992
rect 862 1996 868 1997
rect 862 1992 863 1996
rect 867 1992 868 1996
rect 862 1991 868 1992
rect 910 1996 916 1997
rect 910 1992 911 1996
rect 915 1992 916 1996
rect 910 1991 916 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1006 1996 1012 1997
rect 1006 1992 1007 1996
rect 1011 1992 1012 1996
rect 1006 1991 1012 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1094 1995 1095 1999
rect 1099 1995 1100 1999
rect 1136 1997 1138 2017
rect 1160 2005 1162 2017
rect 1186 2015 1192 2016
rect 1186 2011 1187 2015
rect 1191 2011 1192 2015
rect 1186 2010 1192 2011
rect 1158 2004 1164 2005
rect 1158 2000 1159 2004
rect 1163 2000 1164 2004
rect 1158 1999 1164 2000
rect 1094 1994 1100 1995
rect 1134 1996 1140 1997
rect 1046 1991 1052 1992
rect 1096 1991 1098 1994
rect 1134 1992 1135 1996
rect 1139 1992 1140 1996
rect 1188 1992 1190 2010
rect 1240 2005 1242 2017
rect 1238 2004 1244 2005
rect 1238 2000 1239 2004
rect 1243 2000 1244 2004
rect 1238 1999 1244 2000
rect 1268 1992 1270 2022
rect 1303 2017 1307 2018
rect 1351 2022 1355 2023
rect 1351 2017 1355 2018
rect 1352 2005 1354 2017
rect 1360 2016 1362 2046
rect 1398 2040 1404 2041
rect 1398 2036 1399 2040
rect 1403 2036 1404 2040
rect 1398 2035 1404 2036
rect 1400 2023 1402 2035
rect 1488 2028 1490 2090
rect 1518 2080 1524 2081
rect 1518 2076 1519 2080
rect 1523 2076 1524 2080
rect 1518 2075 1524 2076
rect 1598 2080 1604 2081
rect 1598 2076 1599 2080
rect 1603 2076 1604 2080
rect 1598 2075 1604 2076
rect 1495 2074 1499 2075
rect 1495 2069 1499 2070
rect 1519 2074 1523 2075
rect 1519 2069 1523 2070
rect 1591 2074 1595 2075
rect 1591 2069 1595 2070
rect 1599 2074 1603 2075
rect 1599 2069 1603 2070
rect 1494 2068 1500 2069
rect 1494 2064 1495 2068
rect 1499 2064 1500 2068
rect 1494 2063 1500 2064
rect 1590 2068 1596 2069
rect 1590 2064 1591 2068
rect 1595 2064 1596 2068
rect 1590 2063 1596 2064
rect 1616 2052 1618 2114
rect 1628 2096 1630 2114
rect 1648 2096 1650 2126
rect 1663 2121 1667 2122
rect 1679 2126 1683 2127
rect 1679 2121 1683 2122
rect 1735 2126 1739 2127
rect 1735 2121 1739 2122
rect 1751 2126 1755 2127
rect 1751 2121 1755 2122
rect 1680 2109 1682 2121
rect 1752 2109 1754 2121
rect 1760 2120 1762 2150
rect 1768 2132 1770 2158
rect 1806 2144 1812 2145
rect 1806 2140 1807 2144
rect 1811 2140 1812 2144
rect 1806 2139 1812 2140
rect 1766 2131 1772 2132
rect 1766 2127 1767 2131
rect 1771 2127 1772 2131
rect 1808 2127 1810 2139
rect 1816 2132 1818 2194
rect 2118 2187 2124 2188
rect 2118 2183 2119 2187
rect 2123 2183 2124 2187
rect 2118 2182 2124 2183
rect 2120 2179 2122 2182
rect 1879 2178 1883 2179
rect 1879 2173 1883 2174
rect 2119 2178 2123 2179
rect 2119 2173 2123 2174
rect 1878 2172 1884 2173
rect 1878 2168 1879 2172
rect 1883 2168 1884 2172
rect 2120 2170 2122 2173
rect 1878 2167 1884 2168
rect 2118 2169 2124 2170
rect 2118 2165 2119 2169
rect 2123 2165 2124 2169
rect 2118 2164 2124 2165
rect 1870 2155 1876 2156
rect 1870 2151 1871 2155
rect 1875 2151 1876 2155
rect 1870 2150 1876 2151
rect 2118 2152 2124 2153
rect 1872 2132 1874 2150
rect 2118 2148 2119 2152
rect 2123 2148 2124 2152
rect 2118 2147 2124 2148
rect 1878 2144 1884 2145
rect 1878 2140 1879 2144
rect 1883 2140 1884 2144
rect 1878 2139 1884 2140
rect 1814 2131 1820 2132
rect 1814 2127 1815 2131
rect 1819 2127 1820 2131
rect 1870 2131 1876 2132
rect 1870 2127 1871 2131
rect 1875 2127 1876 2131
rect 1880 2127 1882 2139
rect 2120 2127 2122 2147
rect 1766 2126 1772 2127
rect 1807 2126 1811 2127
rect 1814 2126 1820 2127
rect 1823 2126 1827 2127
rect 1870 2126 1876 2127
rect 1879 2126 1883 2127
rect 1807 2121 1811 2122
rect 1823 2121 1827 2122
rect 1879 2121 1883 2122
rect 1887 2126 1891 2127
rect 1887 2121 1891 2122
rect 1951 2126 1955 2127
rect 1951 2121 1955 2122
rect 2023 2126 2027 2127
rect 2023 2121 2027 2122
rect 2071 2126 2075 2127
rect 2071 2121 2075 2122
rect 2119 2126 2123 2127
rect 2119 2121 2123 2122
rect 1758 2119 1764 2120
rect 1758 2115 1759 2119
rect 1763 2115 1764 2119
rect 1758 2114 1764 2115
rect 1798 2119 1804 2120
rect 1798 2115 1799 2119
rect 1803 2115 1804 2119
rect 1798 2114 1804 2115
rect 1678 2108 1684 2109
rect 1678 2104 1679 2108
rect 1683 2104 1684 2108
rect 1678 2103 1684 2104
rect 1750 2108 1756 2109
rect 1750 2104 1751 2108
rect 1755 2104 1756 2108
rect 1750 2103 1756 2104
rect 1800 2096 1802 2114
rect 1824 2109 1826 2121
rect 1866 2119 1872 2120
rect 1866 2115 1867 2119
rect 1871 2115 1872 2119
rect 1866 2114 1872 2115
rect 1822 2108 1828 2109
rect 1822 2104 1823 2108
rect 1827 2104 1828 2108
rect 1822 2103 1828 2104
rect 1868 2096 1870 2114
rect 1888 2109 1890 2121
rect 1952 2109 1954 2121
rect 1982 2119 1988 2120
rect 1982 2115 1983 2119
rect 1987 2115 1988 2119
rect 1982 2114 1988 2115
rect 1994 2119 2000 2120
rect 1994 2115 1995 2119
rect 1999 2115 2000 2119
rect 1994 2114 2000 2115
rect 1886 2108 1892 2109
rect 1886 2104 1887 2108
rect 1891 2104 1892 2108
rect 1886 2103 1892 2104
rect 1950 2108 1956 2109
rect 1950 2104 1951 2108
rect 1955 2104 1956 2108
rect 1950 2103 1956 2104
rect 1626 2095 1632 2096
rect 1626 2091 1627 2095
rect 1631 2091 1632 2095
rect 1626 2090 1632 2091
rect 1646 2095 1652 2096
rect 1646 2091 1647 2095
rect 1651 2091 1652 2095
rect 1646 2090 1652 2091
rect 1798 2095 1804 2096
rect 1798 2091 1799 2095
rect 1803 2091 1804 2095
rect 1798 2090 1804 2091
rect 1866 2095 1872 2096
rect 1866 2091 1867 2095
rect 1871 2091 1872 2095
rect 1866 2090 1872 2091
rect 1902 2095 1908 2096
rect 1902 2091 1903 2095
rect 1907 2091 1908 2095
rect 1902 2090 1908 2091
rect 1678 2080 1684 2081
rect 1678 2076 1679 2080
rect 1683 2076 1684 2080
rect 1678 2075 1684 2076
rect 1750 2080 1756 2081
rect 1750 2076 1751 2080
rect 1755 2076 1756 2080
rect 1750 2075 1756 2076
rect 1822 2080 1828 2081
rect 1822 2076 1823 2080
rect 1827 2076 1828 2080
rect 1822 2075 1828 2076
rect 1886 2080 1892 2081
rect 1886 2076 1887 2080
rect 1891 2076 1892 2080
rect 1886 2075 1892 2076
rect 1679 2074 1683 2075
rect 1679 2069 1683 2070
rect 1751 2074 1755 2075
rect 1751 2069 1755 2070
rect 1759 2074 1763 2075
rect 1759 2069 1763 2070
rect 1823 2074 1827 2075
rect 1823 2069 1827 2070
rect 1831 2074 1835 2075
rect 1831 2069 1835 2070
rect 1887 2074 1891 2075
rect 1887 2069 1891 2070
rect 1895 2074 1899 2075
rect 1895 2069 1899 2070
rect 1678 2068 1684 2069
rect 1678 2064 1679 2068
rect 1683 2064 1684 2068
rect 1678 2063 1684 2064
rect 1758 2068 1764 2069
rect 1758 2064 1759 2068
rect 1763 2064 1764 2068
rect 1758 2063 1764 2064
rect 1830 2068 1836 2069
rect 1830 2064 1831 2068
rect 1835 2064 1836 2068
rect 1830 2063 1836 2064
rect 1894 2068 1900 2069
rect 1894 2064 1895 2068
rect 1899 2064 1900 2068
rect 1894 2063 1900 2064
rect 1614 2051 1620 2052
rect 1614 2047 1615 2051
rect 1619 2047 1620 2051
rect 1614 2046 1620 2047
rect 1646 2051 1652 2052
rect 1646 2047 1647 2051
rect 1651 2047 1652 2051
rect 1646 2046 1652 2047
rect 1750 2051 1756 2052
rect 1750 2047 1751 2051
rect 1755 2047 1756 2051
rect 1750 2046 1756 2047
rect 1494 2040 1500 2041
rect 1494 2036 1495 2040
rect 1499 2036 1500 2040
rect 1494 2035 1500 2036
rect 1590 2040 1596 2041
rect 1590 2036 1591 2040
rect 1595 2036 1596 2040
rect 1590 2035 1596 2036
rect 1486 2027 1492 2028
rect 1486 2023 1487 2027
rect 1491 2023 1492 2027
rect 1496 2023 1498 2035
rect 1592 2023 1594 2035
rect 1648 2028 1650 2046
rect 1678 2040 1684 2041
rect 1678 2036 1679 2040
rect 1683 2036 1684 2040
rect 1678 2035 1684 2036
rect 1646 2027 1652 2028
rect 1646 2023 1647 2027
rect 1651 2023 1652 2027
rect 1670 2027 1676 2028
rect 1670 2023 1671 2027
rect 1675 2023 1676 2027
rect 1680 2023 1682 2035
rect 1399 2022 1403 2023
rect 1399 2017 1403 2018
rect 1455 2022 1459 2023
rect 1486 2022 1492 2023
rect 1495 2022 1499 2023
rect 1455 2017 1459 2018
rect 1495 2017 1499 2018
rect 1559 2022 1563 2023
rect 1559 2017 1563 2018
rect 1591 2022 1595 2023
rect 1646 2022 1652 2023
rect 1655 2022 1659 2023
rect 1670 2022 1676 2023
rect 1679 2022 1683 2023
rect 1591 2017 1595 2018
rect 1655 2017 1659 2018
rect 1358 2015 1364 2016
rect 1358 2011 1359 2015
rect 1363 2011 1364 2015
rect 1358 2010 1364 2011
rect 1378 2015 1384 2016
rect 1378 2011 1379 2015
rect 1383 2011 1384 2015
rect 1378 2010 1384 2011
rect 1350 2004 1356 2005
rect 1350 2000 1351 2004
rect 1355 2000 1356 2004
rect 1350 1999 1356 2000
rect 1380 1992 1382 2010
rect 1456 2005 1458 2017
rect 1560 2005 1562 2017
rect 1646 2015 1652 2016
rect 1646 2011 1647 2015
rect 1651 2011 1652 2015
rect 1646 2010 1652 2011
rect 1454 2004 1460 2005
rect 1454 2000 1455 2004
rect 1459 2000 1460 2004
rect 1454 1999 1460 2000
rect 1558 2004 1564 2005
rect 1558 2000 1559 2004
rect 1563 2000 1564 2004
rect 1558 1999 1564 2000
rect 1134 1991 1140 1992
rect 1186 1991 1192 1992
rect 687 1990 691 1991
rect 687 1985 691 1986
rect 695 1990 699 1991
rect 695 1985 699 1986
rect 759 1990 763 1991
rect 759 1985 763 1986
rect 815 1990 819 1991
rect 815 1985 819 1986
rect 831 1990 835 1991
rect 831 1985 835 1986
rect 863 1990 867 1991
rect 863 1985 867 1986
rect 911 1990 915 1991
rect 911 1985 915 1986
rect 959 1990 963 1991
rect 959 1985 963 1986
rect 991 1990 995 1991
rect 991 1985 995 1986
rect 1007 1990 1011 1991
rect 1007 1985 1011 1986
rect 1047 1990 1051 1991
rect 1047 1985 1051 1986
rect 1095 1990 1099 1991
rect 1186 1987 1187 1991
rect 1191 1987 1192 1991
rect 1186 1986 1192 1987
rect 1266 1991 1272 1992
rect 1266 1987 1267 1991
rect 1271 1987 1272 1991
rect 1266 1986 1272 1987
rect 1378 1991 1384 1992
rect 1378 1987 1379 1991
rect 1383 1987 1384 1991
rect 1378 1986 1384 1987
rect 1566 1991 1572 1992
rect 1566 1987 1567 1991
rect 1571 1987 1572 1991
rect 1566 1986 1572 1987
rect 1095 1985 1099 1986
rect 686 1984 692 1985
rect 686 1980 687 1984
rect 691 1980 692 1984
rect 686 1979 692 1980
rect 758 1984 764 1985
rect 758 1980 759 1984
rect 763 1980 764 1984
rect 758 1979 764 1980
rect 830 1984 836 1985
rect 830 1980 831 1984
rect 835 1980 836 1984
rect 830 1979 836 1980
rect 910 1984 916 1985
rect 910 1980 911 1984
rect 915 1980 916 1984
rect 910 1979 916 1980
rect 990 1984 996 1985
rect 990 1980 991 1984
rect 995 1980 996 1984
rect 1096 1982 1098 1985
rect 990 1979 996 1980
rect 1094 1981 1100 1982
rect 1094 1977 1095 1981
rect 1099 1977 1100 1981
rect 1094 1976 1100 1977
rect 1134 1979 1140 1980
rect 642 1975 648 1976
rect 642 1971 643 1975
rect 647 1971 648 1975
rect 642 1970 648 1971
rect 858 1975 864 1976
rect 858 1971 859 1975
rect 863 1971 864 1975
rect 1134 1975 1135 1979
rect 1139 1975 1140 1979
rect 1134 1974 1140 1975
rect 1158 1976 1164 1977
rect 858 1970 864 1971
rect 518 1967 524 1968
rect 518 1963 519 1967
rect 523 1963 524 1967
rect 518 1962 524 1963
rect 598 1967 604 1968
rect 598 1963 599 1967
rect 603 1963 604 1967
rect 598 1962 604 1963
rect 678 1967 684 1968
rect 678 1963 679 1967
rect 683 1963 684 1967
rect 678 1962 684 1963
rect 710 1967 716 1968
rect 710 1963 711 1967
rect 715 1963 716 1967
rect 710 1962 716 1963
rect 520 1944 522 1962
rect 526 1956 532 1957
rect 526 1952 527 1956
rect 531 1952 532 1956
rect 526 1951 532 1952
rect 454 1943 460 1944
rect 454 1939 455 1943
rect 459 1939 460 1943
rect 454 1938 460 1939
rect 518 1943 524 1944
rect 518 1939 519 1943
rect 523 1939 524 1943
rect 518 1938 524 1939
rect 470 1935 476 1936
rect 528 1935 530 1951
rect 600 1944 602 1962
rect 606 1956 612 1957
rect 606 1952 607 1956
rect 611 1952 612 1956
rect 606 1951 612 1952
rect 598 1943 604 1944
rect 598 1939 599 1943
rect 603 1939 604 1943
rect 598 1938 604 1939
rect 608 1935 610 1951
rect 680 1944 682 1962
rect 686 1956 692 1957
rect 686 1952 687 1956
rect 691 1952 692 1956
rect 686 1951 692 1952
rect 678 1943 684 1944
rect 678 1939 679 1943
rect 683 1939 684 1943
rect 678 1938 684 1939
rect 688 1935 690 1951
rect 198 1931 199 1935
rect 203 1931 204 1935
rect 198 1930 204 1931
rect 231 1934 235 1935
rect 182 1927 188 1928
rect 182 1923 183 1927
rect 187 1923 188 1927
rect 182 1922 188 1923
rect 134 1916 140 1917
rect 134 1912 135 1916
rect 139 1912 140 1916
rect 134 1911 140 1912
rect 174 1916 180 1917
rect 174 1912 175 1916
rect 179 1912 180 1916
rect 174 1911 180 1912
rect 110 1908 116 1909
rect 110 1904 111 1908
rect 115 1904 116 1908
rect 200 1904 202 1930
rect 231 1929 235 1930
rect 295 1934 299 1935
rect 295 1929 299 1930
rect 303 1934 307 1935
rect 303 1929 307 1930
rect 367 1934 371 1935
rect 367 1929 371 1930
rect 375 1934 379 1935
rect 375 1929 379 1930
rect 447 1934 451 1935
rect 470 1931 471 1935
rect 475 1931 476 1935
rect 470 1930 476 1931
rect 527 1934 531 1935
rect 447 1929 451 1930
rect 232 1917 234 1929
rect 258 1927 264 1928
rect 258 1923 259 1927
rect 263 1923 264 1927
rect 258 1922 264 1923
rect 230 1916 236 1917
rect 230 1912 231 1916
rect 235 1912 236 1916
rect 230 1911 236 1912
rect 260 1904 262 1922
rect 296 1917 298 1929
rect 322 1927 328 1928
rect 322 1923 323 1927
rect 327 1923 328 1927
rect 322 1922 328 1923
rect 294 1916 300 1917
rect 294 1912 295 1916
rect 299 1912 300 1916
rect 294 1911 300 1912
rect 324 1904 326 1922
rect 368 1917 370 1929
rect 394 1927 400 1928
rect 394 1923 395 1927
rect 399 1923 400 1927
rect 394 1922 400 1923
rect 366 1916 372 1917
rect 366 1912 367 1916
rect 371 1912 372 1916
rect 366 1911 372 1912
rect 396 1904 398 1922
rect 448 1917 450 1929
rect 446 1916 452 1917
rect 446 1912 447 1916
rect 451 1912 452 1916
rect 446 1911 452 1912
rect 472 1904 474 1930
rect 527 1929 531 1930
rect 607 1934 611 1935
rect 607 1929 611 1930
rect 615 1934 619 1935
rect 615 1929 619 1930
rect 687 1934 691 1935
rect 687 1929 691 1930
rect 703 1934 707 1935
rect 703 1929 707 1930
rect 528 1917 530 1929
rect 554 1927 560 1928
rect 554 1923 555 1927
rect 559 1923 560 1927
rect 554 1922 560 1923
rect 526 1916 532 1917
rect 526 1912 527 1916
rect 531 1912 532 1916
rect 526 1911 532 1912
rect 556 1904 558 1922
rect 616 1917 618 1929
rect 704 1917 706 1929
rect 712 1928 714 1962
rect 758 1956 764 1957
rect 758 1952 759 1956
rect 763 1952 764 1956
rect 758 1951 764 1952
rect 830 1956 836 1957
rect 830 1952 831 1956
rect 835 1952 836 1956
rect 830 1951 836 1952
rect 726 1935 732 1936
rect 760 1935 762 1951
rect 832 1935 834 1951
rect 860 1944 862 1970
rect 982 1967 988 1968
rect 982 1963 983 1967
rect 987 1963 988 1967
rect 982 1962 988 1963
rect 1094 1964 1100 1965
rect 910 1956 916 1957
rect 910 1952 911 1956
rect 915 1952 916 1956
rect 910 1951 916 1952
rect 858 1943 864 1944
rect 858 1939 859 1943
rect 863 1939 864 1943
rect 858 1938 864 1939
rect 902 1943 908 1944
rect 902 1939 903 1943
rect 907 1939 908 1943
rect 902 1938 908 1939
rect 726 1931 727 1935
rect 731 1931 732 1935
rect 726 1930 732 1931
rect 759 1934 763 1935
rect 710 1927 716 1928
rect 710 1923 711 1927
rect 715 1923 716 1927
rect 710 1922 716 1923
rect 614 1916 620 1917
rect 614 1912 615 1916
rect 619 1912 620 1916
rect 614 1911 620 1912
rect 702 1916 708 1917
rect 702 1912 703 1916
rect 707 1912 708 1916
rect 702 1911 708 1912
rect 728 1904 730 1930
rect 759 1929 763 1930
rect 791 1934 795 1935
rect 791 1929 795 1930
rect 831 1934 835 1935
rect 831 1929 835 1930
rect 879 1934 883 1935
rect 879 1929 883 1930
rect 792 1917 794 1929
rect 810 1927 816 1928
rect 810 1923 811 1927
rect 815 1923 816 1927
rect 810 1922 816 1923
rect 818 1927 824 1928
rect 818 1923 819 1927
rect 823 1923 824 1927
rect 818 1922 824 1923
rect 790 1916 796 1917
rect 790 1912 791 1916
rect 795 1912 796 1916
rect 790 1911 796 1912
rect 110 1903 116 1904
rect 162 1903 168 1904
rect 162 1899 163 1903
rect 167 1899 168 1903
rect 162 1898 168 1899
rect 198 1903 204 1904
rect 198 1899 199 1903
rect 203 1899 204 1903
rect 198 1898 204 1899
rect 258 1903 264 1904
rect 258 1899 259 1903
rect 263 1899 264 1903
rect 258 1898 264 1899
rect 322 1903 328 1904
rect 322 1899 323 1903
rect 327 1899 328 1903
rect 322 1898 328 1899
rect 394 1903 400 1904
rect 394 1899 395 1903
rect 399 1899 400 1903
rect 394 1898 400 1899
rect 470 1903 476 1904
rect 470 1899 471 1903
rect 475 1899 476 1903
rect 470 1898 476 1899
rect 554 1903 560 1904
rect 554 1899 555 1903
rect 559 1899 560 1903
rect 554 1898 560 1899
rect 638 1903 644 1904
rect 638 1899 639 1903
rect 643 1899 644 1903
rect 638 1898 644 1899
rect 726 1903 732 1904
rect 726 1899 727 1903
rect 731 1899 732 1903
rect 726 1898 732 1899
rect 110 1891 116 1892
rect 110 1887 111 1891
rect 115 1887 116 1891
rect 110 1886 116 1887
rect 134 1888 140 1889
rect 112 1879 114 1886
rect 134 1884 135 1888
rect 139 1884 140 1888
rect 134 1883 140 1884
rect 136 1879 138 1883
rect 111 1878 115 1879
rect 111 1873 115 1874
rect 135 1878 139 1879
rect 135 1873 139 1874
rect 112 1870 114 1873
rect 134 1872 140 1873
rect 110 1869 116 1870
rect 110 1865 111 1869
rect 115 1865 116 1869
rect 134 1868 135 1872
rect 139 1868 140 1872
rect 134 1867 140 1868
rect 110 1864 116 1865
rect 142 1855 148 1856
rect 110 1852 116 1853
rect 110 1848 111 1852
rect 115 1848 116 1852
rect 142 1851 143 1855
rect 147 1851 148 1855
rect 142 1850 148 1851
rect 110 1847 116 1848
rect 112 1823 114 1847
rect 134 1844 140 1845
rect 134 1840 135 1844
rect 139 1840 140 1844
rect 134 1839 140 1840
rect 136 1823 138 1839
rect 111 1822 115 1823
rect 111 1817 115 1818
rect 135 1822 139 1823
rect 135 1817 139 1818
rect 112 1797 114 1817
rect 136 1805 138 1817
rect 144 1816 146 1850
rect 164 1832 166 1898
rect 174 1888 180 1889
rect 174 1884 175 1888
rect 179 1884 180 1888
rect 174 1883 180 1884
rect 230 1888 236 1889
rect 230 1884 231 1888
rect 235 1884 236 1888
rect 230 1883 236 1884
rect 294 1888 300 1889
rect 294 1884 295 1888
rect 299 1884 300 1888
rect 294 1883 300 1884
rect 366 1888 372 1889
rect 366 1884 367 1888
rect 371 1884 372 1888
rect 366 1883 372 1884
rect 446 1888 452 1889
rect 446 1884 447 1888
rect 451 1884 452 1888
rect 446 1883 452 1884
rect 526 1888 532 1889
rect 526 1884 527 1888
rect 531 1884 532 1888
rect 526 1883 532 1884
rect 614 1888 620 1889
rect 614 1884 615 1888
rect 619 1884 620 1888
rect 614 1883 620 1884
rect 176 1879 178 1883
rect 232 1879 234 1883
rect 296 1879 298 1883
rect 368 1879 370 1883
rect 448 1879 450 1883
rect 528 1879 530 1883
rect 616 1879 618 1883
rect 175 1878 179 1879
rect 175 1873 179 1874
rect 223 1878 227 1879
rect 223 1873 227 1874
rect 231 1878 235 1879
rect 231 1873 235 1874
rect 287 1878 291 1879
rect 287 1873 291 1874
rect 295 1878 299 1879
rect 295 1873 299 1874
rect 359 1878 363 1879
rect 359 1873 363 1874
rect 367 1878 371 1879
rect 367 1873 371 1874
rect 431 1878 435 1879
rect 431 1873 435 1874
rect 447 1878 451 1879
rect 447 1873 451 1874
rect 503 1878 507 1879
rect 503 1873 507 1874
rect 527 1878 531 1879
rect 527 1873 531 1874
rect 567 1878 571 1879
rect 567 1873 571 1874
rect 615 1878 619 1879
rect 615 1873 619 1874
rect 631 1878 635 1879
rect 631 1873 635 1874
rect 174 1872 180 1873
rect 174 1868 175 1872
rect 179 1868 180 1872
rect 174 1867 180 1868
rect 222 1872 228 1873
rect 222 1868 223 1872
rect 227 1868 228 1872
rect 222 1867 228 1868
rect 286 1872 292 1873
rect 286 1868 287 1872
rect 291 1868 292 1872
rect 286 1867 292 1868
rect 358 1872 364 1873
rect 358 1868 359 1872
rect 363 1868 364 1872
rect 358 1867 364 1868
rect 430 1872 436 1873
rect 430 1868 431 1872
rect 435 1868 436 1872
rect 430 1867 436 1868
rect 502 1872 508 1873
rect 502 1868 503 1872
rect 507 1868 508 1872
rect 502 1867 508 1868
rect 566 1872 572 1873
rect 566 1868 567 1872
rect 571 1868 572 1872
rect 566 1867 572 1868
rect 630 1872 636 1873
rect 630 1868 631 1872
rect 635 1868 636 1872
rect 630 1867 636 1868
rect 310 1863 316 1864
rect 310 1859 311 1863
rect 315 1859 316 1863
rect 310 1858 316 1859
rect 526 1863 532 1864
rect 526 1859 527 1863
rect 531 1859 532 1863
rect 526 1858 532 1859
rect 214 1855 220 1856
rect 214 1851 215 1855
rect 219 1851 220 1855
rect 214 1850 220 1851
rect 230 1855 236 1856
rect 230 1851 231 1855
rect 235 1851 236 1855
rect 230 1850 236 1851
rect 174 1844 180 1845
rect 174 1840 175 1844
rect 179 1840 180 1844
rect 174 1839 180 1840
rect 162 1831 168 1832
rect 162 1827 163 1831
rect 167 1827 168 1831
rect 162 1826 168 1827
rect 176 1823 178 1839
rect 216 1832 218 1850
rect 222 1844 228 1845
rect 222 1840 223 1844
rect 227 1840 228 1844
rect 222 1839 228 1840
rect 214 1831 220 1832
rect 214 1827 215 1831
rect 219 1827 220 1831
rect 214 1826 220 1827
rect 224 1823 226 1839
rect 232 1824 234 1850
rect 286 1844 292 1845
rect 286 1840 287 1844
rect 291 1840 292 1844
rect 286 1839 292 1840
rect 230 1823 236 1824
rect 288 1823 290 1839
rect 312 1832 314 1858
rect 422 1855 428 1856
rect 422 1851 423 1855
rect 427 1851 428 1855
rect 422 1850 428 1851
rect 358 1844 364 1845
rect 358 1840 359 1844
rect 363 1840 364 1844
rect 358 1839 364 1840
rect 310 1831 316 1832
rect 310 1827 311 1831
rect 315 1827 316 1831
rect 310 1826 316 1827
rect 360 1823 362 1839
rect 424 1832 426 1850
rect 430 1844 436 1845
rect 430 1840 431 1844
rect 435 1840 436 1844
rect 430 1839 436 1840
rect 502 1844 508 1845
rect 502 1840 503 1844
rect 507 1840 508 1844
rect 502 1839 508 1840
rect 374 1831 380 1832
rect 374 1827 375 1831
rect 379 1827 380 1831
rect 374 1826 380 1827
rect 422 1831 428 1832
rect 422 1827 423 1831
rect 427 1827 428 1831
rect 422 1826 428 1827
rect 175 1822 179 1823
rect 175 1817 179 1818
rect 183 1822 187 1823
rect 183 1817 187 1818
rect 223 1822 227 1823
rect 230 1819 231 1823
rect 235 1819 236 1823
rect 230 1818 236 1819
rect 263 1822 267 1823
rect 223 1817 227 1818
rect 263 1817 267 1818
rect 287 1822 291 1823
rect 287 1817 291 1818
rect 351 1822 355 1823
rect 351 1817 355 1818
rect 359 1822 363 1823
rect 359 1817 363 1818
rect 142 1815 148 1816
rect 142 1811 143 1815
rect 147 1811 148 1815
rect 142 1810 148 1811
rect 162 1815 168 1816
rect 162 1811 163 1815
rect 167 1811 168 1815
rect 162 1810 168 1811
rect 134 1804 140 1805
rect 134 1800 135 1804
rect 139 1800 140 1804
rect 134 1799 140 1800
rect 110 1796 116 1797
rect 110 1792 111 1796
rect 115 1792 116 1796
rect 164 1792 166 1810
rect 184 1805 186 1817
rect 264 1805 266 1817
rect 298 1815 304 1816
rect 298 1811 299 1815
rect 303 1811 304 1815
rect 298 1810 304 1811
rect 182 1804 188 1805
rect 182 1800 183 1804
rect 187 1800 188 1804
rect 182 1799 188 1800
rect 262 1804 268 1805
rect 262 1800 263 1804
rect 267 1800 268 1804
rect 262 1799 268 1800
rect 300 1792 302 1810
rect 352 1805 354 1817
rect 350 1804 356 1805
rect 350 1800 351 1804
rect 355 1800 356 1804
rect 350 1799 356 1800
rect 376 1792 378 1826
rect 432 1823 434 1839
rect 462 1823 468 1824
rect 504 1823 506 1839
rect 528 1832 530 1858
rect 558 1855 564 1856
rect 558 1851 559 1855
rect 563 1851 564 1855
rect 558 1850 564 1851
rect 594 1855 600 1856
rect 594 1851 595 1855
rect 599 1851 600 1855
rect 594 1850 600 1851
rect 560 1832 562 1850
rect 566 1844 572 1845
rect 566 1840 567 1844
rect 571 1840 572 1844
rect 566 1839 572 1840
rect 526 1831 532 1832
rect 526 1827 527 1831
rect 531 1827 532 1831
rect 526 1826 532 1827
rect 558 1831 564 1832
rect 558 1827 559 1831
rect 563 1827 564 1831
rect 558 1826 564 1827
rect 568 1823 570 1839
rect 431 1822 435 1823
rect 431 1817 435 1818
rect 439 1822 443 1823
rect 462 1819 463 1823
rect 467 1819 468 1823
rect 462 1818 468 1819
rect 503 1822 507 1823
rect 439 1817 443 1818
rect 440 1805 442 1817
rect 438 1804 444 1805
rect 438 1800 439 1804
rect 443 1800 444 1804
rect 438 1799 444 1800
rect 464 1792 466 1818
rect 503 1817 507 1818
rect 527 1822 531 1823
rect 527 1817 531 1818
rect 567 1822 571 1823
rect 567 1817 571 1818
rect 510 1815 516 1816
rect 510 1811 511 1815
rect 515 1811 516 1815
rect 510 1810 516 1811
rect 518 1815 524 1816
rect 518 1811 519 1815
rect 523 1811 524 1815
rect 518 1810 524 1811
rect 512 1792 514 1810
rect 110 1791 116 1792
rect 162 1791 168 1792
rect 162 1787 163 1791
rect 167 1787 168 1791
rect 162 1786 168 1787
rect 170 1791 176 1792
rect 170 1787 171 1791
rect 175 1787 176 1791
rect 170 1786 176 1787
rect 298 1791 304 1792
rect 298 1787 299 1791
rect 303 1787 304 1791
rect 298 1786 304 1787
rect 374 1791 380 1792
rect 374 1787 375 1791
rect 379 1787 380 1791
rect 374 1786 380 1787
rect 462 1791 468 1792
rect 462 1787 463 1791
rect 467 1787 468 1791
rect 462 1786 468 1787
rect 510 1791 516 1792
rect 510 1787 511 1791
rect 515 1787 516 1791
rect 510 1786 516 1787
rect 110 1779 116 1780
rect 110 1775 111 1779
rect 115 1775 116 1779
rect 110 1774 116 1775
rect 134 1776 140 1777
rect 112 1763 114 1774
rect 134 1772 135 1776
rect 139 1772 140 1776
rect 134 1771 140 1772
rect 136 1763 138 1771
rect 111 1762 115 1763
rect 111 1757 115 1758
rect 135 1762 139 1763
rect 135 1757 139 1758
rect 112 1754 114 1757
rect 134 1756 140 1757
rect 110 1753 116 1754
rect 110 1749 111 1753
rect 115 1749 116 1753
rect 134 1752 135 1756
rect 139 1752 140 1756
rect 134 1751 140 1752
rect 110 1748 116 1749
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 112 1707 114 1731
rect 134 1728 140 1729
rect 134 1724 135 1728
rect 139 1724 140 1728
rect 134 1723 140 1724
rect 136 1707 138 1723
rect 172 1716 174 1786
rect 182 1776 188 1777
rect 182 1772 183 1776
rect 187 1772 188 1776
rect 182 1771 188 1772
rect 262 1776 268 1777
rect 262 1772 263 1776
rect 267 1772 268 1776
rect 262 1771 268 1772
rect 350 1776 356 1777
rect 350 1772 351 1776
rect 355 1772 356 1776
rect 350 1771 356 1772
rect 438 1776 444 1777
rect 438 1772 439 1776
rect 443 1772 444 1776
rect 438 1771 444 1772
rect 184 1763 186 1771
rect 264 1763 266 1771
rect 352 1763 354 1771
rect 440 1763 442 1771
rect 183 1762 187 1763
rect 183 1757 187 1758
rect 199 1762 203 1763
rect 199 1757 203 1758
rect 263 1762 267 1763
rect 263 1757 267 1758
rect 295 1762 299 1763
rect 295 1757 299 1758
rect 351 1762 355 1763
rect 351 1757 355 1758
rect 399 1762 403 1763
rect 399 1757 403 1758
rect 439 1762 443 1763
rect 439 1757 443 1758
rect 495 1762 499 1763
rect 495 1757 499 1758
rect 198 1756 204 1757
rect 198 1752 199 1756
rect 203 1752 204 1756
rect 198 1751 204 1752
rect 294 1756 300 1757
rect 294 1752 295 1756
rect 299 1752 300 1756
rect 294 1751 300 1752
rect 398 1756 404 1757
rect 398 1752 399 1756
rect 403 1752 404 1756
rect 398 1751 404 1752
rect 494 1756 500 1757
rect 494 1752 495 1756
rect 499 1752 500 1756
rect 494 1751 500 1752
rect 430 1747 436 1748
rect 430 1743 431 1747
rect 435 1743 436 1747
rect 430 1742 436 1743
rect 182 1739 188 1740
rect 182 1735 183 1739
rect 187 1735 188 1739
rect 182 1734 188 1735
rect 286 1739 292 1740
rect 286 1735 287 1739
rect 291 1735 292 1739
rect 286 1734 292 1735
rect 310 1739 316 1740
rect 310 1735 311 1739
rect 315 1735 316 1739
rect 310 1734 316 1735
rect 184 1716 186 1734
rect 198 1728 204 1729
rect 198 1724 199 1728
rect 203 1724 204 1728
rect 198 1723 204 1724
rect 170 1715 176 1716
rect 170 1711 171 1715
rect 175 1711 176 1715
rect 170 1710 176 1711
rect 182 1715 188 1716
rect 182 1711 183 1715
rect 187 1711 188 1715
rect 182 1710 188 1711
rect 200 1707 202 1723
rect 288 1716 290 1734
rect 294 1728 300 1729
rect 294 1724 295 1728
rect 299 1724 300 1728
rect 294 1723 300 1724
rect 286 1715 292 1716
rect 286 1711 287 1715
rect 291 1711 292 1715
rect 286 1710 292 1711
rect 296 1707 298 1723
rect 312 1708 314 1734
rect 398 1728 404 1729
rect 398 1724 399 1728
rect 403 1724 404 1728
rect 398 1723 404 1724
rect 310 1707 316 1708
rect 400 1707 402 1723
rect 432 1716 434 1742
rect 520 1740 522 1810
rect 528 1805 530 1817
rect 596 1816 598 1850
rect 630 1844 636 1845
rect 630 1840 631 1844
rect 635 1840 636 1844
rect 630 1839 636 1840
rect 632 1823 634 1839
rect 640 1832 642 1898
rect 702 1888 708 1889
rect 702 1884 703 1888
rect 707 1884 708 1888
rect 702 1883 708 1884
rect 790 1888 796 1889
rect 790 1884 791 1888
rect 795 1884 796 1888
rect 790 1883 796 1884
rect 704 1879 706 1883
rect 792 1879 794 1883
rect 695 1878 699 1879
rect 695 1873 699 1874
rect 703 1878 707 1879
rect 703 1873 707 1874
rect 759 1878 763 1879
rect 759 1873 763 1874
rect 791 1878 795 1879
rect 791 1873 795 1874
rect 694 1872 700 1873
rect 694 1868 695 1872
rect 699 1868 700 1872
rect 694 1867 700 1868
rect 758 1872 764 1873
rect 758 1868 759 1872
rect 763 1868 764 1872
rect 758 1867 764 1868
rect 812 1864 814 1922
rect 820 1904 822 1922
rect 880 1917 882 1929
rect 878 1916 884 1917
rect 878 1912 879 1916
rect 883 1912 884 1916
rect 878 1911 884 1912
rect 904 1904 906 1938
rect 912 1935 914 1951
rect 984 1944 986 1962
rect 1094 1960 1095 1964
rect 1099 1960 1100 1964
rect 1094 1959 1100 1960
rect 1136 1959 1138 1974
rect 1158 1972 1159 1976
rect 1163 1972 1164 1976
rect 1158 1971 1164 1972
rect 1238 1976 1244 1977
rect 1238 1972 1239 1976
rect 1243 1972 1244 1976
rect 1238 1971 1244 1972
rect 1350 1976 1356 1977
rect 1350 1972 1351 1976
rect 1355 1972 1356 1976
rect 1350 1971 1356 1972
rect 1454 1976 1460 1977
rect 1454 1972 1455 1976
rect 1459 1972 1460 1976
rect 1454 1971 1460 1972
rect 1558 1976 1564 1977
rect 1558 1972 1559 1976
rect 1563 1972 1564 1976
rect 1558 1971 1564 1972
rect 1160 1959 1162 1971
rect 1240 1959 1242 1971
rect 1352 1959 1354 1971
rect 1456 1959 1458 1971
rect 1560 1959 1562 1971
rect 990 1956 996 1957
rect 990 1952 991 1956
rect 995 1952 996 1956
rect 990 1951 996 1952
rect 982 1943 988 1944
rect 982 1939 983 1943
rect 987 1939 988 1943
rect 982 1938 988 1939
rect 992 1935 994 1951
rect 1096 1935 1098 1959
rect 1135 1958 1139 1959
rect 1135 1953 1139 1954
rect 1159 1958 1163 1959
rect 1159 1953 1163 1954
rect 1239 1958 1243 1959
rect 1239 1953 1243 1954
rect 1351 1958 1355 1959
rect 1351 1953 1355 1954
rect 1359 1958 1363 1959
rect 1359 1953 1363 1954
rect 1423 1958 1427 1959
rect 1423 1953 1427 1954
rect 1455 1958 1459 1959
rect 1455 1953 1459 1954
rect 1487 1958 1491 1959
rect 1487 1953 1491 1954
rect 1559 1958 1563 1959
rect 1559 1953 1563 1954
rect 1136 1950 1138 1953
rect 1358 1952 1364 1953
rect 1134 1949 1140 1950
rect 1134 1945 1135 1949
rect 1139 1945 1140 1949
rect 1358 1948 1359 1952
rect 1363 1948 1364 1952
rect 1358 1947 1364 1948
rect 1422 1952 1428 1953
rect 1422 1948 1423 1952
rect 1427 1948 1428 1952
rect 1422 1947 1428 1948
rect 1486 1952 1492 1953
rect 1486 1948 1487 1952
rect 1491 1948 1492 1952
rect 1486 1947 1492 1948
rect 1558 1952 1564 1953
rect 1558 1948 1559 1952
rect 1563 1948 1564 1952
rect 1558 1947 1564 1948
rect 1134 1944 1140 1945
rect 1382 1943 1388 1944
rect 1382 1939 1383 1943
rect 1387 1939 1388 1943
rect 1382 1938 1388 1939
rect 911 1934 915 1935
rect 911 1929 915 1930
rect 991 1934 995 1935
rect 991 1929 995 1930
rect 1095 1934 1099 1935
rect 1095 1929 1099 1930
rect 1134 1932 1140 1933
rect 1096 1909 1098 1929
rect 1134 1928 1135 1932
rect 1139 1928 1140 1932
rect 1134 1927 1140 1928
rect 1094 1908 1100 1909
rect 1094 1904 1095 1908
rect 1099 1904 1100 1908
rect 1136 1907 1138 1927
rect 1358 1924 1364 1925
rect 1358 1920 1359 1924
rect 1363 1920 1364 1924
rect 1358 1919 1364 1920
rect 1342 1907 1348 1908
rect 1360 1907 1362 1919
rect 1384 1912 1386 1938
rect 1414 1935 1420 1936
rect 1414 1931 1415 1935
rect 1419 1931 1420 1935
rect 1414 1930 1420 1931
rect 1446 1935 1452 1936
rect 1446 1931 1447 1935
rect 1451 1931 1452 1935
rect 1446 1930 1452 1931
rect 1416 1912 1418 1930
rect 1422 1924 1428 1925
rect 1422 1920 1423 1924
rect 1427 1920 1428 1924
rect 1422 1919 1428 1920
rect 1382 1911 1388 1912
rect 1382 1907 1383 1911
rect 1387 1907 1388 1911
rect 818 1903 824 1904
rect 818 1899 819 1903
rect 823 1899 824 1903
rect 818 1898 824 1899
rect 902 1903 908 1904
rect 1094 1903 1100 1904
rect 1135 1906 1139 1907
rect 902 1899 903 1903
rect 907 1899 908 1903
rect 1135 1901 1139 1902
rect 1231 1906 1235 1907
rect 1231 1901 1235 1902
rect 1271 1906 1275 1907
rect 1271 1901 1275 1902
rect 1319 1906 1323 1907
rect 1342 1903 1343 1907
rect 1347 1903 1348 1907
rect 1342 1902 1348 1903
rect 1359 1906 1363 1907
rect 1319 1901 1323 1902
rect 902 1898 908 1899
rect 1094 1891 1100 1892
rect 878 1888 884 1889
rect 878 1884 879 1888
rect 883 1884 884 1888
rect 1094 1887 1095 1891
rect 1099 1887 1100 1891
rect 1094 1886 1100 1887
rect 878 1883 884 1884
rect 880 1879 882 1883
rect 1096 1879 1098 1886
rect 1136 1881 1138 1901
rect 1232 1889 1234 1901
rect 1258 1899 1264 1900
rect 1258 1895 1259 1899
rect 1263 1895 1264 1899
rect 1258 1894 1264 1895
rect 1230 1888 1236 1889
rect 1230 1884 1231 1888
rect 1235 1884 1236 1888
rect 1230 1883 1236 1884
rect 1134 1880 1140 1881
rect 831 1878 835 1879
rect 831 1873 835 1874
rect 879 1878 883 1879
rect 879 1873 883 1874
rect 1095 1878 1099 1879
rect 1134 1876 1135 1880
rect 1139 1876 1140 1880
rect 1260 1876 1262 1894
rect 1272 1889 1274 1901
rect 1320 1889 1322 1901
rect 1270 1888 1276 1889
rect 1270 1884 1271 1888
rect 1275 1884 1276 1888
rect 1270 1883 1276 1884
rect 1318 1888 1324 1889
rect 1318 1884 1319 1888
rect 1323 1884 1324 1888
rect 1318 1883 1324 1884
rect 1344 1876 1346 1902
rect 1359 1901 1363 1902
rect 1375 1906 1379 1907
rect 1382 1906 1388 1907
rect 1414 1911 1420 1912
rect 1414 1907 1415 1911
rect 1419 1907 1420 1911
rect 1424 1907 1426 1919
rect 1414 1906 1420 1907
rect 1423 1906 1427 1907
rect 1375 1901 1379 1902
rect 1423 1901 1427 1902
rect 1439 1906 1443 1907
rect 1439 1901 1443 1902
rect 1376 1889 1378 1901
rect 1440 1889 1442 1901
rect 1448 1900 1450 1930
rect 1486 1924 1492 1925
rect 1486 1920 1487 1924
rect 1491 1920 1492 1924
rect 1486 1919 1492 1920
rect 1558 1924 1564 1925
rect 1558 1920 1559 1924
rect 1563 1920 1564 1924
rect 1558 1919 1564 1920
rect 1474 1907 1480 1908
rect 1488 1907 1490 1919
rect 1560 1907 1562 1919
rect 1568 1912 1570 1986
rect 1631 1958 1635 1959
rect 1631 1953 1635 1954
rect 1630 1952 1636 1953
rect 1630 1948 1631 1952
rect 1635 1948 1636 1952
rect 1630 1947 1636 1948
rect 1648 1936 1650 2010
rect 1656 2005 1658 2017
rect 1654 2004 1660 2005
rect 1654 2000 1655 2004
rect 1659 2000 1660 2004
rect 1654 1999 1660 2000
rect 1672 1992 1674 2022
rect 1679 2017 1683 2018
rect 1743 2022 1747 2023
rect 1743 2017 1747 2018
rect 1744 2005 1746 2017
rect 1752 2016 1754 2046
rect 1758 2040 1764 2041
rect 1758 2036 1759 2040
rect 1763 2036 1764 2040
rect 1758 2035 1764 2036
rect 1830 2040 1836 2041
rect 1830 2036 1831 2040
rect 1835 2036 1836 2040
rect 1830 2035 1836 2036
rect 1894 2040 1900 2041
rect 1894 2036 1895 2040
rect 1899 2036 1900 2040
rect 1894 2035 1900 2036
rect 1760 2023 1762 2035
rect 1832 2023 1834 2035
rect 1896 2023 1898 2035
rect 1904 2028 1906 2090
rect 1950 2080 1956 2081
rect 1950 2076 1951 2080
rect 1955 2076 1956 2080
rect 1950 2075 1956 2076
rect 1951 2074 1955 2075
rect 1951 2069 1955 2070
rect 1959 2074 1963 2075
rect 1959 2069 1963 2070
rect 1958 2068 1964 2069
rect 1958 2064 1959 2068
rect 1963 2064 1964 2068
rect 1958 2063 1964 2064
rect 1984 2052 1986 2114
rect 1996 2096 1998 2114
rect 2024 2109 2026 2121
rect 2050 2119 2056 2120
rect 2050 2115 2051 2119
rect 2055 2115 2056 2119
rect 2050 2114 2056 2115
rect 2022 2108 2028 2109
rect 2022 2104 2023 2108
rect 2027 2104 2028 2108
rect 2022 2103 2028 2104
rect 2052 2096 2054 2114
rect 2072 2109 2074 2121
rect 2070 2108 2076 2109
rect 2070 2104 2071 2108
rect 2075 2104 2076 2108
rect 2070 2103 2076 2104
rect 2120 2101 2122 2121
rect 2118 2100 2124 2101
rect 2118 2096 2119 2100
rect 2123 2096 2124 2100
rect 1994 2095 2000 2096
rect 1994 2091 1995 2095
rect 1999 2091 2000 2095
rect 1994 2090 2000 2091
rect 2050 2095 2056 2096
rect 2050 2091 2051 2095
rect 2055 2091 2056 2095
rect 2050 2090 2056 2091
rect 2058 2095 2064 2096
rect 2118 2095 2124 2096
rect 2058 2091 2059 2095
rect 2063 2091 2064 2095
rect 2058 2090 2064 2091
rect 2022 2080 2028 2081
rect 2022 2076 2023 2080
rect 2027 2076 2028 2080
rect 2022 2075 2028 2076
rect 2023 2074 2027 2075
rect 2023 2069 2027 2070
rect 2022 2068 2028 2069
rect 2022 2064 2023 2068
rect 2027 2064 2028 2068
rect 2022 2063 2028 2064
rect 2060 2059 2062 2090
rect 2118 2083 2124 2084
rect 2070 2080 2076 2081
rect 2070 2076 2071 2080
rect 2075 2076 2076 2080
rect 2118 2079 2119 2083
rect 2123 2079 2124 2083
rect 2118 2078 2124 2079
rect 2070 2075 2076 2076
rect 2120 2075 2122 2078
rect 2071 2074 2075 2075
rect 2071 2069 2075 2070
rect 2119 2074 2123 2075
rect 2119 2069 2123 2070
rect 2070 2068 2076 2069
rect 2070 2064 2071 2068
rect 2075 2064 2076 2068
rect 2120 2066 2122 2069
rect 2070 2063 2076 2064
rect 2118 2065 2124 2066
rect 2118 2061 2119 2065
rect 2123 2061 2124 2065
rect 2118 2060 2124 2061
rect 2056 2057 2062 2059
rect 1982 2051 1988 2052
rect 1982 2047 1983 2051
rect 1987 2047 1988 2051
rect 1982 2046 1988 2047
rect 1958 2040 1964 2041
rect 1958 2036 1959 2040
rect 1963 2036 1964 2040
rect 1958 2035 1964 2036
rect 2022 2040 2028 2041
rect 2022 2036 2023 2040
rect 2027 2036 2028 2040
rect 2022 2035 2028 2036
rect 1902 2027 1908 2028
rect 1902 2023 1903 2027
rect 1907 2023 1908 2027
rect 1960 2023 1962 2035
rect 2024 2023 2026 2035
rect 2056 2028 2058 2057
rect 2062 2051 2068 2052
rect 2062 2047 2063 2051
rect 2067 2047 2068 2051
rect 2062 2046 2068 2047
rect 2078 2051 2084 2052
rect 2078 2047 2079 2051
rect 2083 2047 2084 2051
rect 2078 2046 2084 2047
rect 2118 2048 2124 2049
rect 2064 2028 2066 2046
rect 2070 2040 2076 2041
rect 2070 2036 2071 2040
rect 2075 2036 2076 2040
rect 2070 2035 2076 2036
rect 2054 2027 2060 2028
rect 2054 2023 2055 2027
rect 2059 2023 2060 2027
rect 1759 2022 1763 2023
rect 1759 2017 1763 2018
rect 1823 2022 1827 2023
rect 1823 2017 1827 2018
rect 1831 2022 1835 2023
rect 1831 2017 1835 2018
rect 1895 2022 1899 2023
rect 1902 2022 1908 2023
rect 1959 2022 1963 2023
rect 1895 2017 1899 2018
rect 1959 2017 1963 2018
rect 2023 2022 2027 2023
rect 2054 2022 2060 2023
rect 2062 2027 2068 2028
rect 2062 2023 2063 2027
rect 2067 2023 2068 2027
rect 2072 2023 2074 2035
rect 2062 2022 2068 2023
rect 2071 2022 2075 2023
rect 2023 2017 2027 2018
rect 2071 2017 2075 2018
rect 1750 2015 1756 2016
rect 1750 2011 1751 2015
rect 1755 2011 1756 2015
rect 1750 2010 1756 2011
rect 1770 2015 1776 2016
rect 1770 2011 1771 2015
rect 1775 2011 1776 2015
rect 1770 2010 1776 2011
rect 1742 2004 1748 2005
rect 1742 2000 1743 2004
rect 1747 2000 1748 2004
rect 1742 1999 1748 2000
rect 1772 1992 1774 2010
rect 1824 2005 1826 2017
rect 1850 2015 1856 2016
rect 1850 2011 1851 2015
rect 1855 2011 1856 2015
rect 1850 2010 1856 2011
rect 1822 2004 1828 2005
rect 1822 2000 1823 2004
rect 1827 2000 1828 2004
rect 1822 1999 1828 2000
rect 1852 1992 1854 2010
rect 1896 2005 1898 2017
rect 1938 2015 1944 2016
rect 1938 2011 1939 2015
rect 1943 2011 1944 2015
rect 1938 2010 1944 2011
rect 1894 2004 1900 2005
rect 1894 2000 1895 2004
rect 1899 2000 1900 2004
rect 1894 1999 1900 2000
rect 1940 1992 1942 2010
rect 1960 2005 1962 2017
rect 1986 2015 1992 2016
rect 1986 2011 1987 2015
rect 1991 2011 1992 2015
rect 1986 2010 1992 2011
rect 1958 2004 1964 2005
rect 1958 2000 1959 2004
rect 1963 2000 1964 2004
rect 1958 1999 1964 2000
rect 1988 1992 1990 2010
rect 2024 2005 2026 2017
rect 2072 2005 2074 2017
rect 2080 2016 2082 2046
rect 2118 2044 2119 2048
rect 2123 2044 2124 2048
rect 2118 2043 2124 2044
rect 2120 2023 2122 2043
rect 2119 2022 2123 2023
rect 2119 2017 2123 2018
rect 2078 2015 2084 2016
rect 2078 2011 2079 2015
rect 2083 2011 2084 2015
rect 2078 2010 2084 2011
rect 2022 2004 2028 2005
rect 2022 2000 2023 2004
rect 2027 2000 2028 2004
rect 2022 1999 2028 2000
rect 2070 2004 2076 2005
rect 2070 2000 2071 2004
rect 2075 2000 2076 2004
rect 2070 1999 2076 2000
rect 2120 1997 2122 2017
rect 2118 1996 2124 1997
rect 2118 1992 2119 1996
rect 2123 1992 2124 1996
rect 1670 1991 1676 1992
rect 1670 1987 1671 1991
rect 1675 1987 1676 1991
rect 1670 1986 1676 1987
rect 1770 1991 1776 1992
rect 1770 1987 1771 1991
rect 1775 1987 1776 1991
rect 1770 1986 1776 1987
rect 1850 1991 1856 1992
rect 1850 1987 1851 1991
rect 1855 1987 1856 1991
rect 1850 1986 1856 1987
rect 1938 1991 1944 1992
rect 1938 1987 1939 1991
rect 1943 1987 1944 1991
rect 1938 1986 1944 1987
rect 1986 1991 1992 1992
rect 1986 1987 1987 1991
rect 1991 1987 1992 1991
rect 2058 1991 2064 1992
rect 2118 1991 2124 1992
rect 2058 1990 2059 1991
rect 1986 1986 1992 1987
rect 2056 1987 2059 1990
rect 2063 1987 2064 1991
rect 2056 1986 2064 1987
rect 1654 1976 1660 1977
rect 1654 1972 1655 1976
rect 1659 1972 1660 1976
rect 1654 1971 1660 1972
rect 1742 1976 1748 1977
rect 1742 1972 1743 1976
rect 1747 1972 1748 1976
rect 1742 1971 1748 1972
rect 1822 1976 1828 1977
rect 1822 1972 1823 1976
rect 1827 1972 1828 1976
rect 1822 1971 1828 1972
rect 1894 1976 1900 1977
rect 1894 1972 1895 1976
rect 1899 1972 1900 1976
rect 1894 1971 1900 1972
rect 1958 1976 1964 1977
rect 1958 1972 1959 1976
rect 1963 1972 1964 1976
rect 1958 1971 1964 1972
rect 2022 1976 2028 1977
rect 2022 1972 2023 1976
rect 2027 1972 2028 1976
rect 2022 1971 2028 1972
rect 1656 1959 1658 1971
rect 1744 1959 1746 1971
rect 1824 1959 1826 1971
rect 1896 1959 1898 1971
rect 1960 1959 1962 1971
rect 2024 1959 2026 1971
rect 1655 1958 1659 1959
rect 1655 1953 1659 1954
rect 1703 1958 1707 1959
rect 1703 1953 1707 1954
rect 1743 1958 1747 1959
rect 1743 1953 1747 1954
rect 1775 1958 1779 1959
rect 1775 1953 1779 1954
rect 1823 1958 1827 1959
rect 1823 1953 1827 1954
rect 1847 1958 1851 1959
rect 1847 1953 1851 1954
rect 1895 1958 1899 1959
rect 1895 1953 1899 1954
rect 1927 1958 1931 1959
rect 1927 1953 1931 1954
rect 1959 1958 1963 1959
rect 1959 1953 1963 1954
rect 2007 1958 2011 1959
rect 2007 1953 2011 1954
rect 2023 1958 2027 1959
rect 2023 1953 2027 1954
rect 1702 1952 1708 1953
rect 1702 1948 1703 1952
rect 1707 1948 1708 1952
rect 1702 1947 1708 1948
rect 1774 1952 1780 1953
rect 1774 1948 1775 1952
rect 1779 1948 1780 1952
rect 1774 1947 1780 1948
rect 1846 1952 1852 1953
rect 1846 1948 1847 1952
rect 1851 1948 1852 1952
rect 1846 1947 1852 1948
rect 1926 1952 1932 1953
rect 1926 1948 1927 1952
rect 1931 1948 1932 1952
rect 1926 1947 1932 1948
rect 2006 1952 2012 1953
rect 2006 1948 2007 1952
rect 2011 1948 2012 1952
rect 2006 1947 2012 1948
rect 1646 1935 1652 1936
rect 1646 1931 1647 1935
rect 1651 1931 1652 1935
rect 1646 1930 1652 1931
rect 1630 1924 1636 1925
rect 1630 1920 1631 1924
rect 1635 1920 1636 1924
rect 1630 1919 1636 1920
rect 1702 1924 1708 1925
rect 1702 1920 1703 1924
rect 1707 1920 1708 1924
rect 1702 1919 1708 1920
rect 1774 1924 1780 1925
rect 1774 1920 1775 1924
rect 1779 1920 1780 1924
rect 1774 1919 1780 1920
rect 1846 1924 1852 1925
rect 1846 1920 1847 1924
rect 1851 1920 1852 1924
rect 1846 1919 1852 1920
rect 1926 1924 1932 1925
rect 1926 1920 1927 1924
rect 1931 1920 1932 1924
rect 1926 1919 1932 1920
rect 2006 1924 2012 1925
rect 2006 1920 2007 1924
rect 2011 1920 2012 1924
rect 2006 1919 2012 1920
rect 1566 1911 1572 1912
rect 1566 1907 1567 1911
rect 1571 1907 1572 1911
rect 1632 1907 1634 1919
rect 1704 1907 1706 1919
rect 1776 1907 1778 1919
rect 1848 1907 1850 1919
rect 1928 1907 1930 1919
rect 1986 1911 1992 1912
rect 1986 1907 1987 1911
rect 1991 1907 1992 1911
rect 2008 1907 2010 1919
rect 2056 1912 2058 1986
rect 2118 1979 2124 1980
rect 2070 1976 2076 1977
rect 2070 1972 2071 1976
rect 2075 1972 2076 1976
rect 2118 1975 2119 1979
rect 2123 1975 2124 1979
rect 2118 1974 2124 1975
rect 2070 1971 2076 1972
rect 2072 1959 2074 1971
rect 2120 1959 2122 1974
rect 2071 1958 2075 1959
rect 2071 1953 2075 1954
rect 2119 1958 2123 1959
rect 2119 1953 2123 1954
rect 2070 1952 2076 1953
rect 2070 1948 2071 1952
rect 2075 1948 2076 1952
rect 2120 1950 2122 1953
rect 2070 1947 2076 1948
rect 2118 1949 2124 1950
rect 2118 1945 2119 1949
rect 2123 1945 2124 1949
rect 2118 1944 2124 1945
rect 2062 1935 2068 1936
rect 2062 1931 2063 1935
rect 2067 1931 2068 1935
rect 2062 1930 2068 1931
rect 2078 1935 2084 1936
rect 2078 1931 2079 1935
rect 2083 1931 2084 1935
rect 2078 1930 2084 1931
rect 2118 1932 2124 1933
rect 2064 1912 2066 1930
rect 2070 1924 2076 1925
rect 2070 1920 2071 1924
rect 2075 1920 2076 1924
rect 2070 1919 2076 1920
rect 2054 1911 2060 1912
rect 2054 1907 2055 1911
rect 2059 1907 2060 1911
rect 1474 1903 1475 1907
rect 1479 1903 1480 1907
rect 1474 1902 1480 1903
rect 1487 1906 1491 1907
rect 1446 1899 1452 1900
rect 1446 1895 1447 1899
rect 1451 1895 1452 1899
rect 1446 1894 1452 1895
rect 1466 1899 1472 1900
rect 1466 1895 1467 1899
rect 1471 1895 1472 1899
rect 1466 1894 1472 1895
rect 1374 1888 1380 1889
rect 1374 1884 1375 1888
rect 1379 1884 1380 1888
rect 1374 1883 1380 1884
rect 1438 1888 1444 1889
rect 1438 1884 1439 1888
rect 1443 1884 1444 1888
rect 1438 1883 1444 1884
rect 1468 1876 1470 1894
rect 1476 1876 1478 1902
rect 1487 1901 1491 1902
rect 1503 1906 1507 1907
rect 1503 1901 1507 1902
rect 1559 1906 1563 1907
rect 1566 1906 1572 1907
rect 1575 1906 1579 1907
rect 1559 1901 1563 1902
rect 1575 1901 1579 1902
rect 1631 1906 1635 1907
rect 1631 1901 1635 1902
rect 1655 1906 1659 1907
rect 1655 1901 1659 1902
rect 1703 1906 1707 1907
rect 1703 1901 1707 1902
rect 1751 1906 1755 1907
rect 1751 1901 1755 1902
rect 1775 1906 1779 1907
rect 1775 1901 1779 1902
rect 1847 1906 1851 1907
rect 1847 1901 1851 1902
rect 1863 1906 1867 1907
rect 1863 1901 1867 1902
rect 1927 1906 1931 1907
rect 1927 1901 1931 1902
rect 1975 1906 1979 1907
rect 1986 1906 1992 1907
rect 2007 1906 2011 1907
rect 2054 1906 2060 1907
rect 2062 1911 2068 1912
rect 2062 1907 2063 1911
rect 2067 1907 2068 1911
rect 2072 1907 2074 1919
rect 2062 1906 2068 1907
rect 2071 1906 2075 1907
rect 1975 1901 1979 1902
rect 1504 1889 1506 1901
rect 1566 1899 1572 1900
rect 1566 1895 1567 1899
rect 1571 1895 1572 1899
rect 1566 1894 1572 1895
rect 1502 1888 1508 1889
rect 1502 1884 1503 1888
rect 1507 1884 1508 1888
rect 1502 1883 1508 1884
rect 1134 1875 1140 1876
rect 1258 1875 1264 1876
rect 1095 1873 1099 1874
rect 830 1872 836 1873
rect 830 1868 831 1872
rect 835 1868 836 1872
rect 1096 1870 1098 1873
rect 1258 1871 1259 1875
rect 1263 1871 1264 1875
rect 1258 1870 1264 1871
rect 1294 1875 1300 1876
rect 1294 1871 1295 1875
rect 1299 1871 1300 1875
rect 1294 1870 1300 1871
rect 1342 1875 1348 1876
rect 1342 1871 1343 1875
rect 1347 1871 1348 1875
rect 1342 1870 1348 1871
rect 1466 1875 1472 1876
rect 1466 1871 1467 1875
rect 1471 1871 1472 1875
rect 1466 1870 1472 1871
rect 1474 1875 1480 1876
rect 1474 1871 1475 1875
rect 1479 1871 1480 1875
rect 1474 1870 1480 1871
rect 830 1867 836 1868
rect 1094 1869 1100 1870
rect 1094 1865 1095 1869
rect 1099 1865 1100 1869
rect 1094 1864 1100 1865
rect 810 1863 816 1864
rect 810 1859 811 1863
rect 815 1859 816 1863
rect 810 1858 816 1859
rect 1134 1863 1140 1864
rect 1134 1859 1135 1863
rect 1139 1859 1140 1863
rect 1134 1858 1140 1859
rect 1230 1860 1236 1861
rect 750 1855 756 1856
rect 750 1851 751 1855
rect 755 1851 756 1855
rect 750 1850 756 1851
rect 822 1855 828 1856
rect 822 1851 823 1855
rect 827 1851 828 1855
rect 822 1850 828 1851
rect 1094 1852 1100 1853
rect 694 1844 700 1845
rect 694 1840 695 1844
rect 699 1840 700 1844
rect 694 1839 700 1840
rect 638 1831 644 1832
rect 638 1827 639 1831
rect 643 1827 644 1831
rect 638 1826 644 1827
rect 696 1823 698 1839
rect 752 1832 754 1850
rect 758 1844 764 1845
rect 758 1840 759 1844
rect 763 1840 764 1844
rect 758 1839 764 1840
rect 742 1831 748 1832
rect 742 1827 743 1831
rect 747 1827 748 1831
rect 742 1826 748 1827
rect 750 1831 756 1832
rect 750 1827 751 1831
rect 755 1827 756 1831
rect 750 1826 756 1827
rect 607 1822 611 1823
rect 607 1817 611 1818
rect 631 1822 635 1823
rect 631 1817 635 1818
rect 687 1822 691 1823
rect 687 1817 691 1818
rect 695 1822 699 1823
rect 695 1817 699 1818
rect 594 1815 600 1816
rect 594 1811 595 1815
rect 599 1811 600 1815
rect 594 1810 600 1811
rect 608 1805 610 1817
rect 688 1805 690 1817
rect 714 1815 720 1816
rect 714 1811 715 1815
rect 719 1811 720 1815
rect 714 1810 720 1811
rect 526 1804 532 1805
rect 526 1800 527 1804
rect 531 1800 532 1804
rect 526 1799 532 1800
rect 606 1804 612 1805
rect 606 1800 607 1804
rect 611 1800 612 1804
rect 606 1799 612 1800
rect 686 1804 692 1805
rect 686 1800 687 1804
rect 691 1800 692 1804
rect 686 1799 692 1800
rect 716 1792 718 1810
rect 744 1792 746 1826
rect 760 1823 762 1839
rect 824 1832 826 1850
rect 1094 1848 1095 1852
rect 1099 1848 1100 1852
rect 1136 1851 1138 1858
rect 1230 1856 1231 1860
rect 1235 1856 1236 1860
rect 1230 1855 1236 1856
rect 1270 1860 1276 1861
rect 1270 1856 1271 1860
rect 1275 1856 1276 1860
rect 1270 1855 1276 1856
rect 1232 1851 1234 1855
rect 1272 1851 1274 1855
rect 1094 1847 1100 1848
rect 1135 1850 1139 1851
rect 830 1844 836 1845
rect 830 1840 831 1844
rect 835 1840 836 1844
rect 830 1839 836 1840
rect 822 1831 828 1832
rect 822 1827 823 1831
rect 827 1827 828 1831
rect 822 1826 828 1827
rect 832 1823 834 1839
rect 1014 1823 1020 1824
rect 1096 1823 1098 1847
rect 1135 1845 1139 1846
rect 1159 1850 1163 1851
rect 1159 1845 1163 1846
rect 1199 1850 1203 1851
rect 1199 1845 1203 1846
rect 1231 1850 1235 1851
rect 1231 1845 1235 1846
rect 1239 1850 1243 1851
rect 1239 1845 1243 1846
rect 1271 1850 1275 1851
rect 1271 1845 1275 1846
rect 1136 1842 1138 1845
rect 1158 1844 1164 1845
rect 1134 1841 1140 1842
rect 1134 1837 1135 1841
rect 1139 1837 1140 1841
rect 1158 1840 1159 1844
rect 1163 1840 1164 1844
rect 1158 1839 1164 1840
rect 1198 1844 1204 1845
rect 1198 1840 1199 1844
rect 1203 1840 1204 1844
rect 1198 1839 1204 1840
rect 1238 1844 1244 1845
rect 1238 1840 1239 1844
rect 1243 1840 1244 1844
rect 1238 1839 1244 1840
rect 1134 1836 1140 1837
rect 1134 1824 1140 1825
rect 759 1822 763 1823
rect 759 1817 763 1818
rect 767 1822 771 1823
rect 767 1817 771 1818
rect 831 1822 835 1823
rect 831 1817 835 1818
rect 839 1822 843 1823
rect 839 1817 843 1818
rect 911 1822 915 1823
rect 911 1817 915 1818
rect 991 1822 995 1823
rect 1014 1819 1015 1823
rect 1019 1819 1020 1823
rect 1014 1818 1020 1819
rect 1047 1822 1051 1823
rect 991 1817 995 1818
rect 768 1805 770 1817
rect 840 1805 842 1817
rect 866 1815 872 1816
rect 866 1811 867 1815
rect 871 1811 872 1815
rect 866 1810 872 1811
rect 766 1804 772 1805
rect 766 1800 767 1804
rect 771 1800 772 1804
rect 766 1799 772 1800
rect 838 1804 844 1805
rect 838 1800 839 1804
rect 843 1800 844 1804
rect 838 1799 844 1800
rect 868 1792 870 1810
rect 912 1805 914 1817
rect 992 1805 994 1817
rect 910 1804 916 1805
rect 910 1800 911 1804
rect 915 1800 916 1804
rect 910 1799 916 1800
rect 990 1804 996 1805
rect 990 1800 991 1804
rect 995 1800 996 1804
rect 990 1799 996 1800
rect 1016 1792 1018 1818
rect 1047 1817 1051 1818
rect 1095 1822 1099 1823
rect 1134 1820 1135 1824
rect 1139 1820 1140 1824
rect 1134 1819 1140 1820
rect 1095 1817 1099 1818
rect 1034 1815 1040 1816
rect 1034 1811 1035 1815
rect 1039 1811 1040 1815
rect 1034 1810 1040 1811
rect 1036 1792 1038 1810
rect 1048 1805 1050 1817
rect 1046 1804 1052 1805
rect 1046 1800 1047 1804
rect 1051 1800 1052 1804
rect 1046 1799 1052 1800
rect 1096 1797 1098 1817
rect 1094 1796 1100 1797
rect 1094 1792 1095 1796
rect 1099 1792 1100 1796
rect 714 1791 720 1792
rect 714 1787 715 1791
rect 719 1787 720 1791
rect 714 1786 720 1787
rect 742 1791 748 1792
rect 742 1787 743 1791
rect 747 1787 748 1791
rect 742 1786 748 1787
rect 866 1791 872 1792
rect 866 1787 867 1791
rect 871 1787 872 1791
rect 866 1786 872 1787
rect 950 1791 956 1792
rect 950 1787 951 1791
rect 955 1787 956 1791
rect 950 1786 956 1787
rect 1014 1791 1020 1792
rect 1014 1787 1015 1791
rect 1019 1787 1020 1791
rect 1014 1786 1020 1787
rect 1034 1791 1040 1792
rect 1094 1791 1100 1792
rect 1136 1791 1138 1819
rect 1158 1816 1164 1817
rect 1158 1812 1159 1816
rect 1163 1812 1164 1816
rect 1158 1811 1164 1812
rect 1198 1816 1204 1817
rect 1198 1812 1199 1816
rect 1203 1812 1204 1816
rect 1198 1811 1204 1812
rect 1238 1816 1244 1817
rect 1238 1812 1239 1816
rect 1243 1812 1244 1816
rect 1238 1811 1244 1812
rect 1160 1791 1162 1811
rect 1200 1791 1202 1811
rect 1240 1791 1242 1811
rect 1296 1804 1298 1870
rect 1318 1860 1324 1861
rect 1318 1856 1319 1860
rect 1323 1856 1324 1860
rect 1318 1855 1324 1856
rect 1374 1860 1380 1861
rect 1374 1856 1375 1860
rect 1379 1856 1380 1860
rect 1374 1855 1380 1856
rect 1438 1860 1444 1861
rect 1438 1856 1439 1860
rect 1443 1856 1444 1860
rect 1438 1855 1444 1856
rect 1502 1860 1508 1861
rect 1502 1856 1503 1860
rect 1507 1856 1508 1860
rect 1502 1855 1508 1856
rect 1320 1851 1322 1855
rect 1376 1851 1378 1855
rect 1440 1851 1442 1855
rect 1504 1851 1506 1855
rect 1303 1850 1307 1851
rect 1303 1845 1307 1846
rect 1319 1850 1323 1851
rect 1319 1845 1323 1846
rect 1367 1850 1371 1851
rect 1367 1845 1371 1846
rect 1375 1850 1379 1851
rect 1375 1845 1379 1846
rect 1431 1850 1435 1851
rect 1431 1845 1435 1846
rect 1439 1850 1443 1851
rect 1439 1845 1443 1846
rect 1503 1850 1507 1851
rect 1503 1845 1507 1846
rect 1302 1844 1308 1845
rect 1302 1840 1303 1844
rect 1307 1840 1308 1844
rect 1302 1839 1308 1840
rect 1366 1844 1372 1845
rect 1366 1840 1367 1844
rect 1371 1840 1372 1844
rect 1366 1839 1372 1840
rect 1430 1844 1436 1845
rect 1430 1840 1431 1844
rect 1435 1840 1436 1844
rect 1430 1839 1436 1840
rect 1502 1844 1508 1845
rect 1502 1840 1503 1844
rect 1507 1840 1508 1844
rect 1502 1839 1508 1840
rect 1568 1836 1570 1894
rect 1576 1889 1578 1901
rect 1602 1899 1608 1900
rect 1602 1895 1603 1899
rect 1607 1895 1608 1899
rect 1602 1894 1608 1895
rect 1574 1888 1580 1889
rect 1574 1884 1575 1888
rect 1579 1884 1580 1888
rect 1574 1883 1580 1884
rect 1604 1876 1606 1894
rect 1656 1889 1658 1901
rect 1682 1899 1688 1900
rect 1682 1895 1683 1899
rect 1687 1895 1688 1899
rect 1682 1894 1688 1895
rect 1654 1888 1660 1889
rect 1654 1884 1655 1888
rect 1659 1884 1660 1888
rect 1654 1883 1660 1884
rect 1684 1876 1686 1894
rect 1752 1889 1754 1901
rect 1774 1895 1780 1896
rect 1774 1891 1775 1895
rect 1779 1891 1780 1895
rect 1774 1890 1780 1891
rect 1750 1888 1756 1889
rect 1750 1884 1751 1888
rect 1755 1884 1756 1888
rect 1750 1883 1756 1884
rect 1776 1876 1778 1890
rect 1864 1889 1866 1901
rect 1890 1899 1896 1900
rect 1890 1895 1891 1899
rect 1895 1895 1896 1899
rect 1890 1894 1896 1895
rect 1862 1888 1868 1889
rect 1862 1884 1863 1888
rect 1867 1884 1868 1888
rect 1862 1883 1868 1884
rect 1892 1876 1894 1894
rect 1976 1889 1978 1901
rect 1974 1888 1980 1889
rect 1974 1884 1975 1888
rect 1979 1884 1980 1888
rect 1974 1883 1980 1884
rect 1988 1876 1990 1906
rect 2007 1901 2011 1902
rect 2071 1901 2075 1902
rect 2072 1889 2074 1901
rect 2080 1900 2082 1930
rect 2118 1928 2119 1932
rect 2123 1928 2124 1932
rect 2118 1927 2124 1928
rect 2120 1907 2122 1927
rect 2119 1906 2123 1907
rect 2119 1901 2123 1902
rect 2078 1899 2084 1900
rect 2078 1895 2079 1899
rect 2083 1895 2084 1899
rect 2078 1894 2084 1895
rect 2070 1888 2076 1889
rect 2070 1884 2071 1888
rect 2075 1884 2076 1888
rect 2070 1883 2076 1884
rect 2120 1881 2122 1901
rect 2118 1880 2124 1881
rect 2118 1876 2119 1880
rect 2123 1876 2124 1880
rect 1602 1875 1608 1876
rect 1602 1871 1603 1875
rect 1607 1871 1608 1875
rect 1602 1870 1608 1871
rect 1682 1875 1688 1876
rect 1682 1871 1683 1875
rect 1687 1871 1688 1875
rect 1682 1870 1688 1871
rect 1774 1875 1780 1876
rect 1774 1871 1775 1875
rect 1779 1871 1780 1875
rect 1774 1870 1780 1871
rect 1890 1875 1896 1876
rect 1890 1871 1891 1875
rect 1895 1871 1896 1875
rect 1890 1870 1896 1871
rect 1986 1875 1992 1876
rect 2118 1875 2124 1876
rect 1986 1871 1987 1875
rect 1991 1871 1992 1875
rect 1986 1870 1992 1871
rect 2118 1863 2124 1864
rect 1574 1860 1580 1861
rect 1574 1856 1575 1860
rect 1579 1856 1580 1860
rect 1574 1855 1580 1856
rect 1654 1860 1660 1861
rect 1654 1856 1655 1860
rect 1659 1856 1660 1860
rect 1654 1855 1660 1856
rect 1750 1860 1756 1861
rect 1750 1856 1751 1860
rect 1755 1856 1756 1860
rect 1750 1855 1756 1856
rect 1862 1860 1868 1861
rect 1862 1856 1863 1860
rect 1867 1856 1868 1860
rect 1862 1855 1868 1856
rect 1974 1860 1980 1861
rect 1974 1856 1975 1860
rect 1979 1856 1980 1860
rect 1974 1855 1980 1856
rect 2070 1860 2076 1861
rect 2070 1856 2071 1860
rect 2075 1856 2076 1860
rect 2118 1859 2119 1863
rect 2123 1859 2124 1863
rect 2118 1858 2124 1859
rect 2070 1855 2076 1856
rect 1576 1851 1578 1855
rect 1656 1851 1658 1855
rect 1752 1851 1754 1855
rect 1864 1851 1866 1855
rect 1976 1851 1978 1855
rect 2072 1851 2074 1855
rect 2120 1851 2122 1858
rect 1575 1850 1579 1851
rect 1575 1845 1579 1846
rect 1583 1850 1587 1851
rect 1583 1845 1587 1846
rect 1655 1850 1659 1851
rect 1655 1845 1659 1846
rect 1671 1850 1675 1851
rect 1671 1845 1675 1846
rect 1751 1850 1755 1851
rect 1751 1845 1755 1846
rect 1767 1850 1771 1851
rect 1767 1845 1771 1846
rect 1863 1850 1867 1851
rect 1863 1845 1867 1846
rect 1871 1850 1875 1851
rect 1871 1845 1875 1846
rect 1975 1850 1979 1851
rect 1975 1845 1979 1846
rect 1983 1850 1987 1851
rect 1983 1845 1987 1846
rect 2071 1850 2075 1851
rect 2071 1845 2075 1846
rect 2119 1850 2123 1851
rect 2119 1845 2123 1846
rect 1582 1844 1588 1845
rect 1582 1840 1583 1844
rect 1587 1840 1588 1844
rect 1582 1839 1588 1840
rect 1670 1844 1676 1845
rect 1670 1840 1671 1844
rect 1675 1840 1676 1844
rect 1670 1839 1676 1840
rect 1766 1844 1772 1845
rect 1766 1840 1767 1844
rect 1771 1840 1772 1844
rect 1766 1839 1772 1840
rect 1870 1844 1876 1845
rect 1870 1840 1871 1844
rect 1875 1840 1876 1844
rect 1870 1839 1876 1840
rect 1982 1844 1988 1845
rect 1982 1840 1983 1844
rect 1987 1840 1988 1844
rect 1982 1839 1988 1840
rect 2070 1844 2076 1845
rect 2070 1840 2071 1844
rect 2075 1840 2076 1844
rect 2120 1842 2122 1845
rect 2070 1839 2076 1840
rect 2118 1841 2124 1842
rect 2118 1837 2119 1841
rect 2123 1837 2124 1841
rect 2118 1836 2124 1837
rect 1566 1835 1572 1836
rect 1566 1831 1567 1835
rect 1571 1831 1572 1835
rect 1566 1830 1572 1831
rect 1358 1827 1364 1828
rect 1358 1823 1359 1827
rect 1363 1823 1364 1827
rect 1358 1822 1364 1823
rect 1374 1827 1380 1828
rect 1374 1823 1375 1827
rect 1379 1823 1380 1827
rect 1374 1822 1380 1823
rect 1494 1827 1500 1828
rect 1494 1823 1495 1827
rect 1499 1823 1500 1827
rect 1494 1822 1500 1823
rect 1574 1827 1580 1828
rect 1574 1823 1575 1827
rect 1579 1823 1580 1827
rect 1574 1822 1580 1823
rect 1662 1827 1668 1828
rect 1662 1823 1663 1827
rect 1667 1823 1668 1827
rect 1662 1822 1668 1823
rect 1758 1827 1764 1828
rect 1758 1823 1759 1827
rect 1763 1823 1764 1827
rect 1758 1822 1764 1823
rect 1862 1827 1868 1828
rect 1862 1823 1863 1827
rect 1867 1823 1868 1827
rect 1862 1822 1868 1823
rect 2062 1827 2068 1828
rect 2062 1823 2063 1827
rect 2067 1823 2068 1827
rect 2062 1822 2068 1823
rect 2078 1827 2084 1828
rect 2078 1823 2079 1827
rect 2083 1823 2084 1827
rect 2078 1822 2084 1823
rect 2118 1824 2124 1825
rect 1302 1816 1308 1817
rect 1302 1812 1303 1816
rect 1307 1812 1308 1816
rect 1302 1811 1308 1812
rect 1294 1803 1300 1804
rect 1294 1799 1295 1803
rect 1299 1799 1300 1803
rect 1294 1798 1300 1799
rect 1304 1791 1306 1811
rect 1360 1804 1362 1822
rect 1366 1816 1372 1817
rect 1366 1812 1367 1816
rect 1371 1812 1372 1816
rect 1366 1811 1372 1812
rect 1358 1803 1364 1804
rect 1358 1799 1359 1803
rect 1363 1799 1364 1803
rect 1358 1798 1364 1799
rect 1368 1791 1370 1811
rect 1376 1796 1378 1822
rect 1430 1816 1436 1817
rect 1430 1812 1431 1816
rect 1435 1812 1436 1816
rect 1430 1811 1436 1812
rect 1439 1812 1443 1813
rect 1374 1795 1380 1796
rect 1374 1791 1375 1795
rect 1379 1791 1380 1795
rect 1432 1791 1434 1811
rect 1439 1807 1443 1808
rect 1440 1804 1442 1807
rect 1496 1804 1498 1822
rect 1502 1816 1508 1817
rect 1502 1812 1503 1816
rect 1507 1812 1508 1816
rect 1502 1811 1508 1812
rect 1438 1803 1444 1804
rect 1438 1799 1439 1803
rect 1443 1799 1444 1803
rect 1438 1798 1444 1799
rect 1494 1803 1500 1804
rect 1494 1799 1495 1803
rect 1499 1799 1500 1803
rect 1494 1798 1500 1799
rect 1504 1791 1506 1811
rect 1576 1804 1578 1822
rect 1582 1816 1588 1817
rect 1582 1812 1583 1816
rect 1587 1812 1588 1816
rect 1582 1811 1588 1812
rect 1574 1803 1580 1804
rect 1574 1799 1575 1803
rect 1579 1799 1580 1803
rect 1574 1798 1580 1799
rect 1584 1791 1586 1811
rect 1664 1804 1666 1822
rect 1670 1816 1676 1817
rect 1670 1812 1671 1816
rect 1675 1812 1676 1816
rect 1670 1811 1676 1812
rect 1662 1803 1668 1804
rect 1662 1799 1663 1803
rect 1667 1799 1668 1803
rect 1662 1798 1668 1799
rect 1672 1791 1674 1811
rect 1760 1804 1762 1822
rect 1766 1816 1772 1817
rect 1766 1812 1767 1816
rect 1771 1812 1772 1816
rect 1766 1811 1772 1812
rect 1758 1803 1764 1804
rect 1758 1799 1759 1803
rect 1763 1799 1764 1803
rect 1758 1798 1764 1799
rect 1768 1791 1770 1811
rect 1864 1804 1866 1822
rect 1870 1816 1876 1817
rect 1870 1812 1871 1816
rect 1875 1812 1876 1816
rect 1870 1811 1876 1812
rect 1982 1816 1988 1817
rect 1982 1812 1983 1816
rect 1987 1812 1988 1816
rect 1982 1811 1988 1812
rect 2007 1812 2011 1813
rect 1862 1803 1868 1804
rect 1862 1799 1863 1803
rect 1867 1799 1868 1803
rect 1862 1798 1868 1799
rect 1872 1791 1874 1811
rect 1984 1791 1986 1811
rect 2007 1807 2011 1808
rect 1034 1787 1035 1791
rect 1039 1787 1040 1791
rect 1034 1786 1040 1787
rect 1135 1790 1139 1791
rect 526 1776 532 1777
rect 526 1772 527 1776
rect 531 1772 532 1776
rect 526 1771 532 1772
rect 606 1776 612 1777
rect 606 1772 607 1776
rect 611 1772 612 1776
rect 606 1771 612 1772
rect 686 1776 692 1777
rect 686 1772 687 1776
rect 691 1772 692 1776
rect 686 1771 692 1772
rect 766 1776 772 1777
rect 766 1772 767 1776
rect 771 1772 772 1776
rect 766 1771 772 1772
rect 838 1776 844 1777
rect 838 1772 839 1776
rect 843 1772 844 1776
rect 838 1771 844 1772
rect 910 1776 916 1777
rect 910 1772 911 1776
rect 915 1772 916 1776
rect 910 1771 916 1772
rect 528 1763 530 1771
rect 608 1763 610 1771
rect 688 1763 690 1771
rect 768 1763 770 1771
rect 840 1763 842 1771
rect 912 1763 914 1771
rect 527 1762 531 1763
rect 527 1757 531 1758
rect 591 1762 595 1763
rect 591 1757 595 1758
rect 607 1762 611 1763
rect 607 1757 611 1758
rect 671 1762 675 1763
rect 671 1757 675 1758
rect 687 1762 691 1763
rect 687 1757 691 1758
rect 751 1762 755 1763
rect 751 1757 755 1758
rect 767 1762 771 1763
rect 767 1757 771 1758
rect 823 1762 827 1763
rect 823 1757 827 1758
rect 839 1762 843 1763
rect 839 1757 843 1758
rect 887 1762 891 1763
rect 887 1757 891 1758
rect 911 1762 915 1763
rect 911 1757 915 1758
rect 590 1756 596 1757
rect 590 1752 591 1756
rect 595 1752 596 1756
rect 590 1751 596 1752
rect 670 1756 676 1757
rect 670 1752 671 1756
rect 675 1752 676 1756
rect 670 1751 676 1752
rect 750 1756 756 1757
rect 750 1752 751 1756
rect 755 1752 756 1756
rect 750 1751 756 1752
rect 822 1756 828 1757
rect 822 1752 823 1756
rect 827 1752 828 1756
rect 822 1751 828 1752
rect 886 1756 892 1757
rect 886 1752 887 1756
rect 891 1752 892 1756
rect 886 1751 892 1752
rect 910 1747 916 1748
rect 910 1743 911 1747
rect 915 1743 916 1747
rect 910 1742 916 1743
rect 486 1739 492 1740
rect 486 1735 487 1739
rect 491 1735 492 1739
rect 486 1734 492 1735
rect 518 1739 524 1740
rect 518 1735 519 1739
rect 523 1735 524 1739
rect 518 1734 524 1735
rect 742 1739 748 1740
rect 742 1735 743 1739
rect 747 1735 748 1739
rect 742 1734 748 1735
rect 798 1739 804 1740
rect 798 1735 799 1739
rect 803 1735 804 1739
rect 798 1734 804 1735
rect 488 1716 490 1734
rect 494 1728 500 1729
rect 494 1724 495 1728
rect 499 1724 500 1728
rect 494 1723 500 1724
rect 590 1728 596 1729
rect 590 1724 591 1728
rect 595 1724 596 1728
rect 590 1723 596 1724
rect 670 1728 676 1729
rect 670 1724 671 1728
rect 675 1724 676 1728
rect 670 1723 676 1724
rect 430 1715 436 1716
rect 430 1711 431 1715
rect 435 1711 436 1715
rect 430 1710 436 1711
rect 486 1715 492 1716
rect 486 1711 487 1715
rect 491 1711 492 1715
rect 486 1710 492 1711
rect 496 1707 498 1723
rect 562 1715 568 1716
rect 562 1711 563 1715
rect 567 1711 568 1715
rect 562 1710 568 1711
rect 111 1706 115 1707
rect 111 1701 115 1702
rect 135 1706 139 1707
rect 135 1701 139 1702
rect 151 1706 155 1707
rect 151 1701 155 1702
rect 199 1706 203 1707
rect 199 1701 203 1702
rect 223 1706 227 1707
rect 223 1701 227 1702
rect 295 1706 299 1707
rect 295 1701 299 1702
rect 303 1706 307 1707
rect 310 1703 311 1707
rect 315 1703 316 1707
rect 310 1702 316 1703
rect 383 1706 387 1707
rect 303 1701 307 1702
rect 383 1701 387 1702
rect 399 1706 403 1707
rect 399 1701 403 1702
rect 463 1706 467 1707
rect 463 1701 467 1702
rect 495 1706 499 1707
rect 495 1701 499 1702
rect 535 1706 539 1707
rect 535 1701 539 1702
rect 112 1681 114 1701
rect 152 1689 154 1701
rect 210 1699 216 1700
rect 210 1695 211 1699
rect 215 1695 216 1699
rect 210 1694 216 1695
rect 150 1688 156 1689
rect 150 1684 151 1688
rect 155 1684 156 1688
rect 150 1683 156 1684
rect 110 1680 116 1681
rect 110 1676 111 1680
rect 115 1676 116 1680
rect 212 1676 214 1694
rect 224 1689 226 1701
rect 304 1689 306 1701
rect 322 1699 328 1700
rect 322 1695 323 1699
rect 327 1695 328 1699
rect 322 1694 328 1695
rect 330 1699 336 1700
rect 330 1695 331 1699
rect 335 1695 336 1699
rect 330 1694 336 1695
rect 222 1688 228 1689
rect 222 1684 223 1688
rect 227 1684 228 1688
rect 222 1683 228 1684
rect 302 1688 308 1689
rect 302 1684 303 1688
rect 307 1684 308 1688
rect 302 1683 308 1684
rect 110 1675 116 1676
rect 166 1675 172 1676
rect 166 1671 167 1675
rect 171 1671 172 1675
rect 166 1670 172 1671
rect 210 1675 216 1676
rect 210 1671 211 1675
rect 215 1671 216 1675
rect 210 1670 216 1671
rect 110 1663 116 1664
rect 110 1659 111 1663
rect 115 1659 116 1663
rect 110 1658 116 1659
rect 150 1660 156 1661
rect 112 1651 114 1658
rect 150 1656 151 1660
rect 155 1656 156 1660
rect 150 1655 156 1656
rect 152 1651 154 1655
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 151 1650 155 1651
rect 151 1645 155 1646
rect 112 1642 114 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 110 1636 116 1637
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 112 1591 114 1619
rect 168 1604 170 1670
rect 222 1660 228 1661
rect 222 1656 223 1660
rect 227 1656 228 1660
rect 222 1655 228 1656
rect 302 1660 308 1661
rect 302 1656 303 1660
rect 307 1656 308 1660
rect 302 1655 308 1656
rect 224 1651 226 1655
rect 304 1651 306 1655
rect 175 1650 179 1651
rect 175 1645 179 1646
rect 215 1650 219 1651
rect 215 1645 219 1646
rect 223 1650 227 1651
rect 223 1645 227 1646
rect 255 1650 259 1651
rect 255 1645 259 1646
rect 303 1650 307 1651
rect 303 1645 307 1646
rect 174 1644 180 1645
rect 174 1640 175 1644
rect 179 1640 180 1644
rect 174 1639 180 1640
rect 214 1644 220 1645
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 254 1644 260 1645
rect 254 1640 255 1644
rect 259 1640 260 1644
rect 254 1639 260 1640
rect 302 1644 308 1645
rect 302 1640 303 1644
rect 307 1640 308 1644
rect 302 1639 308 1640
rect 324 1628 326 1694
rect 332 1676 334 1694
rect 384 1689 386 1701
rect 410 1699 416 1700
rect 410 1695 411 1699
rect 415 1695 416 1699
rect 410 1694 416 1695
rect 382 1688 388 1689
rect 382 1684 383 1688
rect 387 1684 388 1688
rect 382 1683 388 1684
rect 412 1676 414 1694
rect 464 1689 466 1701
rect 536 1689 538 1701
rect 462 1688 468 1689
rect 462 1684 463 1688
rect 467 1684 468 1688
rect 462 1683 468 1684
rect 534 1688 540 1689
rect 534 1684 535 1688
rect 539 1684 540 1688
rect 534 1683 540 1684
rect 564 1676 566 1710
rect 592 1707 594 1723
rect 672 1707 674 1723
rect 744 1716 746 1734
rect 750 1728 756 1729
rect 750 1724 751 1728
rect 755 1724 756 1728
rect 750 1723 756 1724
rect 742 1715 748 1716
rect 742 1711 743 1715
rect 747 1711 748 1715
rect 742 1710 748 1711
rect 752 1707 754 1723
rect 591 1706 595 1707
rect 591 1701 595 1702
rect 607 1706 611 1707
rect 607 1701 611 1702
rect 671 1706 675 1707
rect 671 1701 675 1702
rect 735 1706 739 1707
rect 735 1701 739 1702
rect 751 1706 755 1707
rect 751 1701 755 1702
rect 608 1689 610 1701
rect 658 1699 664 1700
rect 658 1695 659 1699
rect 663 1695 664 1699
rect 658 1694 664 1695
rect 606 1688 612 1689
rect 606 1684 607 1688
rect 611 1684 612 1688
rect 606 1683 612 1684
rect 660 1683 662 1694
rect 672 1689 674 1701
rect 736 1689 738 1701
rect 800 1700 802 1734
rect 822 1728 828 1729
rect 822 1724 823 1728
rect 827 1724 828 1728
rect 822 1723 828 1724
rect 886 1728 892 1729
rect 886 1724 887 1728
rect 891 1724 892 1728
rect 886 1723 892 1724
rect 824 1707 826 1723
rect 888 1707 890 1723
rect 912 1716 914 1742
rect 952 1716 954 1786
rect 1135 1785 1139 1786
rect 1159 1790 1163 1791
rect 1159 1785 1163 1786
rect 1199 1790 1203 1791
rect 1199 1785 1203 1786
rect 1239 1790 1243 1791
rect 1239 1785 1243 1786
rect 1303 1790 1307 1791
rect 1303 1785 1307 1786
rect 1311 1790 1315 1791
rect 1311 1785 1315 1786
rect 1351 1790 1355 1791
rect 1351 1785 1355 1786
rect 1367 1790 1371 1791
rect 1374 1790 1380 1791
rect 1391 1790 1395 1791
rect 1367 1785 1371 1786
rect 1391 1785 1395 1786
rect 1431 1790 1435 1791
rect 1431 1785 1435 1786
rect 1471 1790 1475 1791
rect 1471 1785 1475 1786
rect 1503 1790 1507 1791
rect 1503 1785 1507 1786
rect 1511 1790 1515 1791
rect 1511 1785 1515 1786
rect 1551 1790 1555 1791
rect 1551 1785 1555 1786
rect 1583 1790 1587 1791
rect 1583 1785 1587 1786
rect 1607 1790 1611 1791
rect 1607 1785 1611 1786
rect 1671 1790 1675 1791
rect 1671 1785 1675 1786
rect 1679 1790 1683 1791
rect 1679 1785 1683 1786
rect 1767 1790 1771 1791
rect 1767 1785 1771 1786
rect 1871 1790 1875 1791
rect 1871 1785 1875 1786
rect 1983 1790 1987 1791
rect 1983 1785 1987 1786
rect 1094 1779 1100 1780
rect 990 1776 996 1777
rect 990 1772 991 1776
rect 995 1772 996 1776
rect 990 1771 996 1772
rect 1046 1776 1052 1777
rect 1046 1772 1047 1776
rect 1051 1772 1052 1776
rect 1094 1775 1095 1779
rect 1099 1775 1100 1779
rect 1094 1774 1100 1775
rect 1046 1771 1052 1772
rect 992 1763 994 1771
rect 1048 1763 1050 1771
rect 1096 1763 1098 1774
rect 1136 1765 1138 1785
rect 1312 1773 1314 1785
rect 1330 1783 1336 1784
rect 1330 1779 1331 1783
rect 1335 1779 1336 1783
rect 1330 1778 1336 1779
rect 1338 1783 1344 1784
rect 1338 1779 1339 1783
rect 1343 1779 1344 1783
rect 1338 1778 1344 1779
rect 1310 1772 1316 1773
rect 1310 1768 1311 1772
rect 1315 1768 1316 1772
rect 1310 1767 1316 1768
rect 1134 1764 1140 1765
rect 959 1762 963 1763
rect 959 1757 963 1758
rect 991 1762 995 1763
rect 991 1757 995 1758
rect 1031 1762 1035 1763
rect 1031 1757 1035 1758
rect 1047 1762 1051 1763
rect 1047 1757 1051 1758
rect 1095 1762 1099 1763
rect 1134 1760 1135 1764
rect 1139 1760 1140 1764
rect 1134 1759 1140 1760
rect 1095 1757 1099 1758
rect 958 1756 964 1757
rect 958 1752 959 1756
rect 963 1752 964 1756
rect 958 1751 964 1752
rect 1030 1756 1036 1757
rect 1030 1752 1031 1756
rect 1035 1752 1036 1756
rect 1096 1754 1098 1757
rect 1030 1751 1036 1752
rect 1094 1753 1100 1754
rect 1094 1749 1095 1753
rect 1099 1749 1100 1753
rect 1094 1748 1100 1749
rect 1134 1747 1140 1748
rect 1134 1743 1135 1747
rect 1139 1743 1140 1747
rect 1134 1742 1140 1743
rect 1310 1744 1316 1745
rect 1022 1739 1028 1740
rect 1022 1735 1023 1739
rect 1027 1735 1028 1739
rect 1022 1734 1028 1735
rect 1094 1736 1100 1737
rect 958 1728 964 1729
rect 958 1724 959 1728
rect 963 1724 964 1728
rect 958 1723 964 1724
rect 910 1715 916 1716
rect 910 1711 911 1715
rect 915 1711 916 1715
rect 910 1710 916 1711
rect 950 1715 956 1716
rect 950 1711 951 1715
rect 955 1711 956 1715
rect 950 1710 956 1711
rect 960 1707 962 1723
rect 1024 1716 1026 1734
rect 1094 1732 1095 1736
rect 1099 1732 1100 1736
rect 1136 1735 1138 1742
rect 1310 1740 1311 1744
rect 1315 1740 1316 1744
rect 1310 1739 1316 1740
rect 1312 1735 1314 1739
rect 1094 1731 1100 1732
rect 1135 1734 1139 1735
rect 1030 1728 1036 1729
rect 1030 1724 1031 1728
rect 1035 1724 1036 1728
rect 1030 1723 1036 1724
rect 1022 1715 1028 1716
rect 1022 1711 1023 1715
rect 1027 1711 1028 1715
rect 1022 1710 1028 1711
rect 1032 1707 1034 1723
rect 1096 1707 1098 1731
rect 1135 1729 1139 1730
rect 1263 1734 1267 1735
rect 1263 1729 1267 1730
rect 1311 1734 1315 1735
rect 1311 1729 1315 1730
rect 1319 1734 1323 1735
rect 1319 1729 1323 1730
rect 1136 1726 1138 1729
rect 1262 1728 1268 1729
rect 1134 1725 1140 1726
rect 1134 1721 1135 1725
rect 1139 1721 1140 1725
rect 1262 1724 1263 1728
rect 1267 1724 1268 1728
rect 1262 1723 1268 1724
rect 1318 1728 1324 1729
rect 1318 1724 1319 1728
rect 1323 1724 1324 1728
rect 1318 1723 1324 1724
rect 1134 1720 1140 1721
rect 1332 1716 1334 1778
rect 1340 1760 1342 1778
rect 1352 1773 1354 1785
rect 1378 1783 1384 1784
rect 1378 1779 1379 1783
rect 1383 1779 1384 1783
rect 1378 1778 1384 1779
rect 1350 1772 1356 1773
rect 1350 1768 1351 1772
rect 1355 1768 1356 1772
rect 1350 1767 1356 1768
rect 1380 1760 1382 1778
rect 1392 1773 1394 1785
rect 1418 1783 1424 1784
rect 1418 1779 1419 1783
rect 1423 1779 1424 1783
rect 1418 1778 1424 1779
rect 1390 1772 1396 1773
rect 1390 1768 1391 1772
rect 1395 1768 1396 1772
rect 1390 1767 1396 1768
rect 1420 1760 1422 1778
rect 1432 1773 1434 1785
rect 1454 1783 1460 1784
rect 1454 1779 1455 1783
rect 1459 1779 1460 1783
rect 1454 1778 1460 1779
rect 1430 1772 1436 1773
rect 1430 1768 1431 1772
rect 1435 1768 1436 1772
rect 1430 1767 1436 1768
rect 1456 1760 1458 1778
rect 1472 1773 1474 1785
rect 1494 1783 1500 1784
rect 1494 1779 1495 1783
rect 1499 1779 1500 1783
rect 1494 1778 1500 1779
rect 1470 1772 1476 1773
rect 1470 1768 1471 1772
rect 1475 1768 1476 1772
rect 1470 1767 1476 1768
rect 1496 1760 1498 1778
rect 1512 1773 1514 1785
rect 1538 1783 1544 1784
rect 1538 1779 1539 1783
rect 1543 1779 1544 1783
rect 1538 1778 1544 1779
rect 1510 1772 1516 1773
rect 1510 1768 1511 1772
rect 1515 1768 1516 1772
rect 1510 1767 1516 1768
rect 1540 1760 1542 1778
rect 1552 1773 1554 1785
rect 1608 1773 1610 1785
rect 1634 1783 1640 1784
rect 1634 1779 1635 1783
rect 1639 1779 1640 1783
rect 1634 1778 1640 1779
rect 1550 1772 1556 1773
rect 1550 1768 1551 1772
rect 1555 1768 1556 1772
rect 1550 1767 1556 1768
rect 1606 1772 1612 1773
rect 1606 1768 1607 1772
rect 1611 1768 1612 1772
rect 1606 1767 1612 1768
rect 1636 1760 1638 1778
rect 1680 1773 1682 1785
rect 1706 1783 1712 1784
rect 1706 1779 1707 1783
rect 1711 1779 1712 1783
rect 1706 1778 1712 1779
rect 1678 1772 1684 1773
rect 1678 1768 1679 1772
rect 1683 1768 1684 1772
rect 1678 1767 1684 1768
rect 1708 1760 1710 1778
rect 1768 1773 1770 1785
rect 1794 1783 1800 1784
rect 1794 1779 1795 1783
rect 1799 1779 1800 1783
rect 1794 1778 1800 1779
rect 1766 1772 1772 1773
rect 1766 1768 1767 1772
rect 1771 1768 1772 1772
rect 1766 1767 1772 1768
rect 1796 1760 1798 1778
rect 1872 1773 1874 1785
rect 1898 1783 1904 1784
rect 1898 1779 1899 1783
rect 1903 1779 1904 1783
rect 1898 1778 1904 1779
rect 1870 1772 1876 1773
rect 1870 1768 1871 1772
rect 1875 1768 1876 1772
rect 1870 1767 1876 1768
rect 1900 1760 1902 1778
rect 1984 1773 1986 1785
rect 1982 1772 1988 1773
rect 1982 1768 1983 1772
rect 1987 1768 1988 1772
rect 1982 1767 1988 1768
rect 2008 1760 2010 1807
rect 2064 1804 2066 1822
rect 2070 1816 2076 1817
rect 2070 1812 2071 1816
rect 2075 1812 2076 1816
rect 2070 1811 2076 1812
rect 2062 1803 2068 1804
rect 2062 1799 2063 1803
rect 2067 1799 2068 1803
rect 2062 1798 2068 1799
rect 2072 1791 2074 1811
rect 2071 1790 2075 1791
rect 2071 1785 2075 1786
rect 2072 1773 2074 1785
rect 2080 1784 2082 1822
rect 2118 1820 2119 1824
rect 2123 1820 2124 1824
rect 2118 1819 2124 1820
rect 2120 1791 2122 1819
rect 2119 1790 2123 1791
rect 2119 1785 2123 1786
rect 2078 1783 2084 1784
rect 2078 1779 2079 1783
rect 2083 1779 2084 1783
rect 2078 1778 2084 1779
rect 2070 1772 2076 1773
rect 2070 1768 2071 1772
rect 2075 1768 2076 1772
rect 2070 1767 2076 1768
rect 2120 1765 2122 1785
rect 2118 1764 2124 1765
rect 2118 1760 2119 1764
rect 2123 1760 2124 1764
rect 1338 1759 1344 1760
rect 1338 1755 1339 1759
rect 1343 1755 1344 1759
rect 1338 1754 1344 1755
rect 1378 1759 1384 1760
rect 1378 1755 1379 1759
rect 1383 1755 1384 1759
rect 1378 1754 1384 1755
rect 1418 1759 1424 1760
rect 1418 1755 1419 1759
rect 1423 1755 1424 1759
rect 1418 1754 1424 1755
rect 1454 1759 1460 1760
rect 1454 1755 1455 1759
rect 1459 1755 1460 1759
rect 1454 1754 1460 1755
rect 1494 1759 1500 1760
rect 1494 1755 1495 1759
rect 1499 1755 1500 1759
rect 1494 1754 1500 1755
rect 1538 1759 1544 1760
rect 1538 1755 1539 1759
rect 1543 1755 1544 1759
rect 1538 1754 1544 1755
rect 1634 1759 1640 1760
rect 1634 1755 1635 1759
rect 1639 1755 1640 1759
rect 1634 1754 1640 1755
rect 1706 1759 1712 1760
rect 1706 1755 1707 1759
rect 1711 1755 1712 1759
rect 1706 1754 1712 1755
rect 1794 1759 1800 1760
rect 1794 1755 1795 1759
rect 1799 1755 1800 1759
rect 1794 1754 1800 1755
rect 1898 1759 1904 1760
rect 1898 1755 1899 1759
rect 1903 1755 1904 1759
rect 1898 1754 1904 1755
rect 2006 1759 2012 1760
rect 2006 1755 2007 1759
rect 2011 1755 2012 1759
rect 2006 1754 2012 1755
rect 2090 1759 2096 1760
rect 2118 1759 2124 1760
rect 2090 1755 2091 1759
rect 2095 1755 2096 1759
rect 2090 1754 2096 1755
rect 1350 1744 1356 1745
rect 1350 1740 1351 1744
rect 1355 1740 1356 1744
rect 1350 1739 1356 1740
rect 1390 1744 1396 1745
rect 1390 1740 1391 1744
rect 1395 1740 1396 1744
rect 1390 1739 1396 1740
rect 1430 1744 1436 1745
rect 1430 1740 1431 1744
rect 1435 1740 1436 1744
rect 1430 1739 1436 1740
rect 1470 1744 1476 1745
rect 1470 1740 1471 1744
rect 1475 1740 1476 1744
rect 1470 1739 1476 1740
rect 1510 1744 1516 1745
rect 1510 1740 1511 1744
rect 1515 1740 1516 1744
rect 1510 1739 1516 1740
rect 1550 1744 1556 1745
rect 1550 1740 1551 1744
rect 1555 1740 1556 1744
rect 1550 1739 1556 1740
rect 1606 1744 1612 1745
rect 1606 1740 1607 1744
rect 1611 1740 1612 1744
rect 1606 1739 1612 1740
rect 1678 1744 1684 1745
rect 1678 1740 1679 1744
rect 1683 1740 1684 1744
rect 1678 1739 1684 1740
rect 1766 1744 1772 1745
rect 1766 1740 1767 1744
rect 1771 1740 1772 1744
rect 1766 1739 1772 1740
rect 1870 1744 1876 1745
rect 1870 1740 1871 1744
rect 1875 1740 1876 1744
rect 1870 1739 1876 1740
rect 1982 1744 1988 1745
rect 1982 1740 1983 1744
rect 1987 1740 1988 1744
rect 1982 1739 1988 1740
rect 2070 1744 2076 1745
rect 2070 1740 2071 1744
rect 2075 1740 2076 1744
rect 2070 1739 2076 1740
rect 1352 1735 1354 1739
rect 1392 1735 1394 1739
rect 1432 1735 1434 1739
rect 1472 1735 1474 1739
rect 1512 1735 1514 1739
rect 1552 1735 1554 1739
rect 1608 1735 1610 1739
rect 1680 1735 1682 1739
rect 1768 1735 1770 1739
rect 1872 1735 1874 1739
rect 1984 1735 1986 1739
rect 2072 1735 2074 1739
rect 1351 1734 1355 1735
rect 1351 1729 1355 1730
rect 1383 1734 1387 1735
rect 1383 1729 1387 1730
rect 1391 1734 1395 1735
rect 1391 1729 1395 1730
rect 1431 1734 1435 1735
rect 1431 1729 1435 1730
rect 1455 1734 1459 1735
rect 1455 1729 1459 1730
rect 1471 1734 1475 1735
rect 1471 1729 1475 1730
rect 1511 1734 1515 1735
rect 1511 1729 1515 1730
rect 1535 1734 1539 1735
rect 1535 1729 1539 1730
rect 1551 1734 1555 1735
rect 1551 1729 1555 1730
rect 1607 1734 1611 1735
rect 1607 1729 1611 1730
rect 1615 1734 1619 1735
rect 1615 1729 1619 1730
rect 1679 1734 1683 1735
rect 1679 1729 1683 1730
rect 1687 1734 1691 1735
rect 1687 1729 1691 1730
rect 1759 1734 1763 1735
rect 1759 1729 1763 1730
rect 1767 1734 1771 1735
rect 1767 1729 1771 1730
rect 1831 1734 1835 1735
rect 1831 1729 1835 1730
rect 1871 1734 1875 1735
rect 1871 1729 1875 1730
rect 1895 1734 1899 1735
rect 1895 1729 1899 1730
rect 1959 1734 1963 1735
rect 1959 1729 1963 1730
rect 1983 1734 1987 1735
rect 1983 1729 1987 1730
rect 2023 1734 2027 1735
rect 2023 1729 2027 1730
rect 2071 1734 2075 1735
rect 2071 1729 2075 1730
rect 1382 1728 1388 1729
rect 1382 1724 1383 1728
rect 1387 1724 1388 1728
rect 1382 1723 1388 1724
rect 1454 1728 1460 1729
rect 1454 1724 1455 1728
rect 1459 1724 1460 1728
rect 1454 1723 1460 1724
rect 1534 1728 1540 1729
rect 1534 1724 1535 1728
rect 1539 1724 1540 1728
rect 1534 1723 1540 1724
rect 1614 1728 1620 1729
rect 1614 1724 1615 1728
rect 1619 1724 1620 1728
rect 1614 1723 1620 1724
rect 1686 1728 1692 1729
rect 1686 1724 1687 1728
rect 1691 1724 1692 1728
rect 1686 1723 1692 1724
rect 1758 1728 1764 1729
rect 1758 1724 1759 1728
rect 1763 1724 1764 1728
rect 1758 1723 1764 1724
rect 1830 1728 1836 1729
rect 1830 1724 1831 1728
rect 1835 1724 1836 1728
rect 1830 1723 1836 1724
rect 1894 1728 1900 1729
rect 1894 1724 1895 1728
rect 1899 1724 1900 1728
rect 1894 1723 1900 1724
rect 1958 1728 1964 1729
rect 1958 1724 1959 1728
rect 1963 1724 1964 1728
rect 1958 1723 1964 1724
rect 2022 1728 2028 1729
rect 2022 1724 2023 1728
rect 2027 1724 2028 1728
rect 2022 1723 2028 1724
rect 2070 1728 2076 1729
rect 2070 1724 2071 1728
rect 2075 1724 2076 1728
rect 2070 1723 2076 1724
rect 1710 1719 1716 1720
rect 1330 1715 1336 1716
rect 1310 1711 1316 1712
rect 1134 1708 1140 1709
rect 807 1706 811 1707
rect 807 1701 811 1702
rect 823 1706 827 1707
rect 823 1701 827 1702
rect 879 1706 883 1707
rect 879 1701 883 1702
rect 887 1706 891 1707
rect 887 1701 891 1702
rect 959 1706 963 1707
rect 959 1701 963 1702
rect 1031 1706 1035 1707
rect 1031 1701 1035 1702
rect 1095 1706 1099 1707
rect 1134 1704 1135 1708
rect 1139 1704 1140 1708
rect 1310 1707 1311 1711
rect 1315 1707 1316 1711
rect 1330 1711 1331 1715
rect 1335 1711 1336 1715
rect 1710 1715 1711 1719
rect 1715 1715 1716 1719
rect 1710 1714 1716 1715
rect 1330 1710 1336 1711
rect 1374 1711 1380 1712
rect 1310 1706 1316 1707
rect 1374 1707 1375 1711
rect 1379 1707 1380 1711
rect 1374 1706 1380 1707
rect 1446 1711 1452 1712
rect 1446 1707 1447 1711
rect 1451 1707 1452 1711
rect 1446 1706 1452 1707
rect 1526 1711 1532 1712
rect 1526 1707 1527 1711
rect 1531 1707 1532 1711
rect 1526 1706 1532 1707
rect 1606 1711 1612 1712
rect 1606 1707 1607 1711
rect 1611 1707 1612 1711
rect 1606 1706 1612 1707
rect 1134 1703 1140 1704
rect 1095 1701 1099 1702
rect 790 1699 796 1700
rect 790 1695 791 1699
rect 795 1695 796 1699
rect 790 1694 796 1695
rect 798 1699 804 1700
rect 798 1695 799 1699
rect 803 1695 804 1699
rect 798 1694 804 1695
rect 670 1688 676 1689
rect 670 1684 671 1688
rect 675 1684 676 1688
rect 670 1683 676 1684
rect 734 1688 740 1689
rect 734 1684 735 1688
rect 739 1684 740 1688
rect 734 1683 740 1684
rect 660 1681 666 1683
rect 664 1676 666 1681
rect 792 1680 794 1694
rect 808 1689 810 1701
rect 834 1699 840 1700
rect 834 1695 835 1699
rect 839 1695 840 1699
rect 834 1694 840 1695
rect 806 1688 812 1689
rect 806 1684 807 1688
rect 811 1684 812 1688
rect 806 1683 812 1684
rect 790 1679 796 1680
rect 330 1675 336 1676
rect 330 1671 331 1675
rect 335 1671 336 1675
rect 330 1670 336 1671
rect 410 1675 416 1676
rect 410 1671 411 1675
rect 415 1671 416 1675
rect 410 1670 416 1671
rect 562 1675 568 1676
rect 562 1671 563 1675
rect 567 1671 568 1675
rect 562 1670 568 1671
rect 654 1675 660 1676
rect 654 1671 655 1675
rect 659 1671 660 1675
rect 654 1670 660 1671
rect 662 1675 668 1676
rect 662 1671 663 1675
rect 667 1671 668 1675
rect 790 1675 791 1679
rect 795 1675 796 1679
rect 836 1676 838 1694
rect 880 1689 882 1701
rect 878 1688 884 1689
rect 878 1684 879 1688
rect 883 1684 884 1688
rect 878 1683 884 1684
rect 1096 1681 1098 1701
rect 1136 1683 1138 1703
rect 1262 1700 1268 1701
rect 1262 1696 1263 1700
rect 1267 1696 1268 1700
rect 1262 1695 1268 1696
rect 1264 1683 1266 1695
rect 1312 1688 1314 1706
rect 1318 1700 1324 1701
rect 1318 1696 1319 1700
rect 1323 1696 1324 1700
rect 1318 1695 1324 1696
rect 1302 1687 1308 1688
rect 1302 1683 1303 1687
rect 1307 1683 1308 1687
rect 1135 1682 1139 1683
rect 1094 1680 1100 1681
rect 1094 1676 1095 1680
rect 1099 1676 1100 1680
rect 1135 1677 1139 1678
rect 1167 1682 1171 1683
rect 1167 1677 1171 1678
rect 1247 1682 1251 1683
rect 1247 1677 1251 1678
rect 1263 1682 1267 1683
rect 1302 1682 1308 1683
rect 1310 1687 1316 1688
rect 1310 1683 1311 1687
rect 1315 1683 1316 1687
rect 1320 1683 1322 1695
rect 1376 1688 1378 1706
rect 1382 1700 1388 1701
rect 1382 1696 1383 1700
rect 1387 1696 1388 1700
rect 1382 1695 1388 1696
rect 1374 1687 1380 1688
rect 1374 1683 1375 1687
rect 1379 1683 1380 1687
rect 1384 1683 1386 1695
rect 1448 1688 1450 1706
rect 1454 1700 1460 1701
rect 1454 1696 1455 1700
rect 1459 1696 1460 1700
rect 1454 1695 1460 1696
rect 1446 1687 1452 1688
rect 1446 1683 1447 1687
rect 1451 1683 1452 1687
rect 1456 1683 1458 1695
rect 1528 1688 1530 1706
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1526 1687 1532 1688
rect 1526 1683 1527 1687
rect 1531 1683 1532 1687
rect 1536 1683 1538 1695
rect 1608 1688 1610 1706
rect 1614 1700 1620 1701
rect 1614 1696 1615 1700
rect 1619 1696 1620 1700
rect 1614 1695 1620 1696
rect 1686 1700 1692 1701
rect 1686 1696 1687 1700
rect 1691 1696 1692 1700
rect 1686 1695 1692 1696
rect 1606 1687 1612 1688
rect 1606 1683 1607 1687
rect 1611 1683 1612 1687
rect 1616 1683 1618 1695
rect 1688 1683 1690 1695
rect 1712 1688 1714 1714
rect 1742 1711 1748 1712
rect 1742 1707 1743 1711
rect 1747 1707 1748 1711
rect 1742 1706 1748 1707
rect 1806 1711 1812 1712
rect 1806 1707 1807 1711
rect 1811 1707 1812 1711
rect 1806 1706 1812 1707
rect 2082 1711 2088 1712
rect 2082 1707 2083 1711
rect 2087 1707 2088 1711
rect 2082 1706 2088 1707
rect 1744 1688 1746 1706
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1710 1687 1716 1688
rect 1710 1683 1711 1687
rect 1715 1683 1716 1687
rect 1310 1682 1316 1683
rect 1319 1682 1323 1683
rect 1263 1677 1267 1678
rect 790 1674 796 1675
rect 834 1675 840 1676
rect 1094 1675 1100 1676
rect 662 1670 668 1671
rect 834 1671 835 1675
rect 839 1671 840 1675
rect 834 1670 840 1671
rect 382 1660 388 1661
rect 382 1656 383 1660
rect 387 1656 388 1660
rect 382 1655 388 1656
rect 462 1660 468 1661
rect 462 1656 463 1660
rect 467 1656 468 1660
rect 462 1655 468 1656
rect 534 1660 540 1661
rect 534 1656 535 1660
rect 539 1656 540 1660
rect 534 1655 540 1656
rect 606 1660 612 1661
rect 606 1656 607 1660
rect 611 1656 612 1660
rect 606 1655 612 1656
rect 384 1651 386 1655
rect 464 1651 466 1655
rect 470 1651 476 1652
rect 536 1651 538 1655
rect 608 1651 610 1655
rect 359 1650 363 1651
rect 359 1645 363 1646
rect 383 1650 387 1651
rect 383 1645 387 1646
rect 407 1650 411 1651
rect 407 1645 411 1646
rect 455 1650 459 1651
rect 455 1645 459 1646
rect 463 1650 467 1651
rect 470 1647 471 1651
rect 475 1647 476 1651
rect 470 1646 476 1647
rect 503 1650 507 1651
rect 463 1645 467 1646
rect 358 1644 364 1645
rect 358 1640 359 1644
rect 363 1640 364 1644
rect 358 1639 364 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 454 1644 460 1645
rect 454 1640 455 1644
rect 459 1640 460 1644
rect 454 1639 460 1640
rect 330 1635 336 1636
rect 330 1631 331 1635
rect 335 1631 336 1635
rect 330 1630 336 1631
rect 202 1627 208 1628
rect 202 1623 203 1627
rect 207 1623 208 1627
rect 202 1622 208 1623
rect 242 1627 248 1628
rect 242 1623 243 1627
rect 247 1623 248 1627
rect 242 1622 248 1623
rect 278 1627 284 1628
rect 278 1623 279 1627
rect 283 1623 284 1627
rect 278 1622 284 1623
rect 322 1627 328 1628
rect 322 1623 323 1627
rect 327 1623 328 1627
rect 322 1622 328 1623
rect 174 1616 180 1617
rect 174 1612 175 1616
rect 179 1612 180 1616
rect 174 1611 180 1612
rect 166 1603 172 1604
rect 166 1599 167 1603
rect 171 1599 172 1603
rect 166 1598 172 1599
rect 176 1591 178 1611
rect 204 1604 206 1622
rect 214 1616 220 1617
rect 214 1612 215 1616
rect 219 1612 220 1616
rect 214 1611 220 1612
rect 202 1603 208 1604
rect 202 1599 203 1603
rect 207 1599 208 1603
rect 202 1598 208 1599
rect 216 1591 218 1611
rect 244 1604 246 1622
rect 254 1616 260 1617
rect 254 1612 255 1616
rect 259 1612 260 1616
rect 254 1611 260 1612
rect 242 1603 248 1604
rect 242 1599 243 1603
rect 247 1599 248 1603
rect 242 1598 248 1599
rect 256 1591 258 1611
rect 111 1590 115 1591
rect 111 1585 115 1586
rect 143 1590 147 1591
rect 143 1585 147 1586
rect 175 1590 179 1591
rect 175 1585 179 1586
rect 183 1590 187 1591
rect 183 1585 187 1586
rect 215 1590 219 1591
rect 215 1585 219 1586
rect 231 1590 235 1591
rect 231 1585 235 1586
rect 255 1590 259 1591
rect 255 1585 259 1586
rect 112 1565 114 1585
rect 144 1573 146 1585
rect 184 1573 186 1585
rect 232 1573 234 1585
rect 280 1584 282 1622
rect 302 1616 308 1617
rect 302 1612 303 1616
rect 307 1612 308 1616
rect 302 1611 308 1612
rect 304 1591 306 1611
rect 332 1604 334 1630
rect 398 1627 404 1628
rect 398 1623 399 1627
rect 403 1623 404 1627
rect 398 1622 404 1623
rect 358 1616 364 1617
rect 358 1612 359 1616
rect 363 1612 364 1616
rect 358 1611 364 1612
rect 330 1603 336 1604
rect 330 1599 331 1603
rect 335 1599 336 1603
rect 330 1598 336 1599
rect 360 1591 362 1611
rect 400 1604 402 1622
rect 406 1616 412 1617
rect 406 1612 407 1616
rect 411 1612 412 1616
rect 406 1611 412 1612
rect 454 1616 460 1617
rect 454 1612 455 1616
rect 459 1612 460 1616
rect 454 1611 460 1612
rect 374 1603 380 1604
rect 374 1599 375 1603
rect 379 1599 380 1603
rect 374 1598 380 1599
rect 398 1603 404 1604
rect 398 1599 399 1603
rect 403 1599 404 1603
rect 398 1598 404 1599
rect 287 1590 291 1591
rect 287 1585 291 1586
rect 303 1590 307 1591
rect 303 1585 307 1586
rect 351 1590 355 1591
rect 351 1585 355 1586
rect 359 1590 363 1591
rect 359 1585 363 1586
rect 270 1583 276 1584
rect 270 1579 271 1583
rect 275 1579 276 1583
rect 270 1578 276 1579
rect 278 1583 284 1584
rect 278 1579 279 1583
rect 283 1579 284 1583
rect 278 1578 284 1579
rect 142 1572 148 1573
rect 142 1568 143 1572
rect 147 1568 148 1572
rect 142 1567 148 1568
rect 182 1572 188 1573
rect 182 1568 183 1572
rect 187 1568 188 1572
rect 182 1567 188 1568
rect 230 1572 236 1573
rect 230 1568 231 1572
rect 235 1568 236 1572
rect 230 1567 236 1568
rect 110 1564 116 1565
rect 110 1560 111 1564
rect 115 1560 116 1564
rect 272 1560 274 1578
rect 288 1573 290 1585
rect 352 1573 354 1585
rect 286 1572 292 1573
rect 286 1568 287 1572
rect 291 1568 292 1572
rect 286 1567 292 1568
rect 350 1572 356 1573
rect 350 1568 351 1572
rect 355 1568 356 1572
rect 350 1567 356 1568
rect 376 1560 378 1598
rect 408 1591 410 1611
rect 456 1591 458 1611
rect 472 1604 474 1646
rect 503 1645 507 1646
rect 535 1650 539 1651
rect 535 1645 539 1646
rect 551 1650 555 1651
rect 551 1645 555 1646
rect 607 1650 611 1651
rect 607 1645 611 1646
rect 502 1644 508 1645
rect 502 1640 503 1644
rect 507 1640 508 1644
rect 502 1639 508 1640
rect 550 1644 556 1645
rect 550 1640 551 1644
rect 555 1640 556 1644
rect 550 1639 556 1640
rect 606 1644 612 1645
rect 606 1640 607 1644
rect 611 1640 612 1644
rect 606 1639 612 1640
rect 534 1635 540 1636
rect 534 1631 535 1635
rect 539 1631 540 1635
rect 534 1630 540 1631
rect 494 1627 500 1628
rect 494 1623 495 1627
rect 499 1623 500 1627
rect 494 1622 500 1623
rect 496 1604 498 1622
rect 502 1616 508 1617
rect 502 1612 503 1616
rect 507 1612 508 1616
rect 502 1611 508 1612
rect 470 1603 476 1604
rect 470 1599 471 1603
rect 475 1599 476 1603
rect 470 1598 476 1599
rect 494 1603 500 1604
rect 494 1599 495 1603
rect 499 1599 500 1603
rect 494 1598 500 1599
rect 504 1591 506 1611
rect 407 1590 411 1591
rect 407 1585 411 1586
rect 415 1590 419 1591
rect 415 1585 419 1586
rect 455 1590 459 1591
rect 455 1585 459 1586
rect 479 1590 483 1591
rect 479 1585 483 1586
rect 503 1590 507 1591
rect 503 1585 507 1586
rect 416 1573 418 1585
rect 466 1583 472 1584
rect 466 1579 467 1583
rect 471 1579 472 1583
rect 466 1578 472 1579
rect 414 1572 420 1573
rect 414 1568 415 1572
rect 419 1568 420 1572
rect 414 1567 420 1568
rect 468 1560 470 1578
rect 480 1573 482 1585
rect 536 1584 538 1630
rect 542 1627 548 1628
rect 542 1623 543 1627
rect 547 1623 548 1627
rect 542 1622 548 1623
rect 598 1627 604 1628
rect 598 1623 599 1627
rect 603 1623 604 1627
rect 598 1622 604 1623
rect 544 1604 546 1622
rect 550 1616 556 1617
rect 550 1612 551 1616
rect 555 1612 556 1616
rect 550 1611 556 1612
rect 542 1603 548 1604
rect 542 1599 543 1603
rect 547 1599 548 1603
rect 542 1598 548 1599
rect 552 1591 554 1611
rect 600 1604 602 1622
rect 606 1616 612 1617
rect 606 1612 607 1616
rect 611 1612 612 1616
rect 606 1611 612 1612
rect 598 1603 604 1604
rect 598 1599 599 1603
rect 603 1599 604 1603
rect 598 1598 604 1599
rect 558 1591 564 1592
rect 608 1591 610 1611
rect 656 1604 658 1670
rect 1094 1663 1100 1664
rect 670 1660 676 1661
rect 670 1656 671 1660
rect 675 1656 676 1660
rect 670 1655 676 1656
rect 734 1660 740 1661
rect 734 1656 735 1660
rect 739 1656 740 1660
rect 734 1655 740 1656
rect 806 1660 812 1661
rect 806 1656 807 1660
rect 811 1656 812 1660
rect 806 1655 812 1656
rect 878 1660 884 1661
rect 878 1656 879 1660
rect 883 1656 884 1660
rect 1094 1659 1095 1663
rect 1099 1659 1100 1663
rect 1094 1658 1100 1659
rect 878 1655 884 1656
rect 672 1651 674 1655
rect 736 1651 738 1655
rect 808 1651 810 1655
rect 880 1651 882 1655
rect 1096 1651 1098 1658
rect 1136 1657 1138 1677
rect 1168 1665 1170 1677
rect 1186 1675 1192 1676
rect 1186 1671 1187 1675
rect 1191 1671 1192 1675
rect 1186 1670 1192 1671
rect 1194 1675 1200 1676
rect 1194 1671 1195 1675
rect 1199 1671 1200 1675
rect 1194 1670 1200 1671
rect 1166 1664 1172 1665
rect 1166 1660 1167 1664
rect 1171 1660 1172 1664
rect 1166 1659 1172 1660
rect 1134 1656 1140 1657
rect 1134 1652 1135 1656
rect 1139 1652 1140 1656
rect 1134 1651 1140 1652
rect 663 1650 667 1651
rect 663 1645 667 1646
rect 671 1650 675 1651
rect 671 1645 675 1646
rect 719 1650 723 1651
rect 719 1645 723 1646
rect 735 1650 739 1651
rect 735 1645 739 1646
rect 807 1650 811 1651
rect 807 1645 811 1646
rect 879 1650 883 1651
rect 879 1645 883 1646
rect 1095 1650 1099 1651
rect 1095 1645 1099 1646
rect 662 1644 668 1645
rect 662 1640 663 1644
rect 667 1640 668 1644
rect 662 1639 668 1640
rect 718 1644 724 1645
rect 718 1640 719 1644
rect 723 1640 724 1644
rect 1096 1642 1098 1645
rect 718 1639 724 1640
rect 1094 1641 1100 1642
rect 1094 1637 1095 1641
rect 1099 1637 1100 1641
rect 1094 1636 1100 1637
rect 1134 1639 1140 1640
rect 1134 1635 1135 1639
rect 1139 1635 1140 1639
rect 1134 1634 1140 1635
rect 1166 1636 1172 1637
rect 710 1627 716 1628
rect 1136 1627 1138 1634
rect 1166 1632 1167 1636
rect 1171 1632 1172 1636
rect 1166 1631 1172 1632
rect 1168 1627 1170 1631
rect 1178 1627 1184 1628
rect 710 1623 711 1627
rect 715 1623 716 1627
rect 1135 1626 1139 1627
rect 710 1622 716 1623
rect 1094 1624 1100 1625
rect 662 1616 668 1617
rect 662 1612 663 1616
rect 667 1612 668 1616
rect 662 1611 668 1612
rect 654 1603 660 1604
rect 654 1599 655 1603
rect 659 1599 660 1603
rect 654 1598 660 1599
rect 664 1591 666 1611
rect 712 1604 714 1622
rect 1094 1620 1095 1624
rect 1099 1620 1100 1624
rect 1135 1621 1139 1622
rect 1159 1626 1163 1627
rect 1159 1621 1163 1622
rect 1167 1626 1171 1627
rect 1178 1623 1179 1627
rect 1183 1623 1184 1627
rect 1178 1622 1184 1623
rect 1167 1621 1171 1622
rect 1094 1619 1100 1620
rect 718 1616 724 1617
rect 718 1612 719 1616
rect 723 1612 724 1616
rect 718 1611 724 1612
rect 710 1603 716 1604
rect 710 1599 711 1603
rect 715 1599 716 1603
rect 710 1598 716 1599
rect 720 1591 722 1611
rect 1096 1591 1098 1619
rect 1136 1618 1138 1621
rect 1158 1620 1164 1621
rect 1134 1617 1140 1618
rect 1134 1613 1135 1617
rect 1139 1613 1140 1617
rect 1158 1616 1159 1620
rect 1163 1616 1164 1620
rect 1158 1615 1164 1616
rect 1134 1612 1140 1613
rect 1134 1600 1140 1601
rect 1134 1596 1135 1600
rect 1139 1596 1140 1600
rect 1134 1595 1140 1596
rect 543 1590 547 1591
rect 543 1585 547 1586
rect 551 1590 555 1591
rect 558 1587 559 1591
rect 563 1587 564 1591
rect 558 1586 564 1587
rect 607 1590 611 1591
rect 551 1585 555 1586
rect 534 1583 540 1584
rect 534 1579 535 1583
rect 539 1579 540 1583
rect 534 1578 540 1579
rect 544 1573 546 1585
rect 478 1572 484 1573
rect 478 1568 479 1572
rect 483 1568 484 1572
rect 478 1567 484 1568
rect 542 1572 548 1573
rect 542 1568 543 1572
rect 547 1568 548 1572
rect 542 1567 548 1568
rect 110 1559 116 1560
rect 150 1559 156 1560
rect 150 1555 151 1559
rect 155 1555 156 1559
rect 150 1554 156 1555
rect 270 1559 276 1560
rect 270 1555 271 1559
rect 275 1555 276 1559
rect 270 1554 276 1555
rect 374 1559 380 1560
rect 374 1555 375 1559
rect 379 1555 380 1559
rect 374 1554 380 1555
rect 466 1559 472 1560
rect 466 1555 467 1559
rect 471 1555 472 1559
rect 466 1554 472 1555
rect 110 1547 116 1548
rect 110 1543 111 1547
rect 115 1543 116 1547
rect 110 1542 116 1543
rect 142 1544 148 1545
rect 112 1531 114 1542
rect 142 1540 143 1544
rect 147 1540 148 1544
rect 142 1539 148 1540
rect 144 1531 146 1539
rect 111 1530 115 1531
rect 111 1525 115 1526
rect 135 1530 139 1531
rect 135 1525 139 1526
rect 143 1530 147 1531
rect 143 1525 147 1526
rect 112 1522 114 1525
rect 134 1524 140 1525
rect 110 1521 116 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 134 1520 135 1524
rect 139 1520 140 1524
rect 134 1519 140 1520
rect 110 1516 116 1517
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 110 1499 116 1500
rect 112 1471 114 1499
rect 134 1496 140 1497
rect 134 1492 135 1496
rect 139 1492 140 1496
rect 134 1491 140 1492
rect 136 1471 138 1491
rect 152 1484 154 1554
rect 182 1544 188 1545
rect 182 1540 183 1544
rect 187 1540 188 1544
rect 182 1539 188 1540
rect 230 1544 236 1545
rect 230 1540 231 1544
rect 235 1540 236 1544
rect 230 1539 236 1540
rect 286 1544 292 1545
rect 286 1540 287 1544
rect 291 1540 292 1544
rect 286 1539 292 1540
rect 350 1544 356 1545
rect 350 1540 351 1544
rect 355 1540 356 1544
rect 350 1539 356 1540
rect 414 1544 420 1545
rect 414 1540 415 1544
rect 419 1540 420 1544
rect 414 1539 420 1540
rect 478 1544 484 1545
rect 478 1540 479 1544
rect 483 1540 484 1544
rect 478 1539 484 1540
rect 542 1544 548 1545
rect 542 1540 543 1544
rect 547 1540 548 1544
rect 542 1539 548 1540
rect 184 1531 186 1539
rect 232 1531 234 1539
rect 288 1531 290 1539
rect 352 1531 354 1539
rect 416 1531 418 1539
rect 480 1531 482 1539
rect 544 1531 546 1539
rect 175 1530 179 1531
rect 175 1525 179 1526
rect 183 1530 187 1531
rect 183 1525 187 1526
rect 215 1530 219 1531
rect 215 1525 219 1526
rect 231 1530 235 1531
rect 231 1525 235 1526
rect 255 1530 259 1531
rect 255 1525 259 1526
rect 287 1530 291 1531
rect 287 1525 291 1526
rect 295 1530 299 1531
rect 295 1525 299 1526
rect 335 1530 339 1531
rect 335 1525 339 1526
rect 351 1530 355 1531
rect 351 1525 355 1526
rect 375 1530 379 1531
rect 375 1525 379 1526
rect 415 1530 419 1531
rect 415 1525 419 1526
rect 455 1530 459 1531
rect 455 1525 459 1526
rect 479 1530 483 1531
rect 479 1525 483 1526
rect 495 1530 499 1531
rect 495 1525 499 1526
rect 535 1530 539 1531
rect 535 1525 539 1526
rect 543 1530 547 1531
rect 543 1525 547 1526
rect 174 1524 180 1525
rect 174 1520 175 1524
rect 179 1520 180 1524
rect 174 1519 180 1520
rect 214 1524 220 1525
rect 214 1520 215 1524
rect 219 1520 220 1524
rect 214 1519 220 1520
rect 254 1524 260 1525
rect 254 1520 255 1524
rect 259 1520 260 1524
rect 254 1519 260 1520
rect 294 1524 300 1525
rect 294 1520 295 1524
rect 299 1520 300 1524
rect 294 1519 300 1520
rect 334 1524 340 1525
rect 334 1520 335 1524
rect 339 1520 340 1524
rect 334 1519 340 1520
rect 374 1524 380 1525
rect 374 1520 375 1524
rect 379 1520 380 1524
rect 374 1519 380 1520
rect 414 1524 420 1525
rect 414 1520 415 1524
rect 419 1520 420 1524
rect 414 1519 420 1520
rect 454 1524 460 1525
rect 454 1520 455 1524
rect 459 1520 460 1524
rect 454 1519 460 1520
rect 494 1524 500 1525
rect 494 1520 495 1524
rect 499 1520 500 1524
rect 494 1519 500 1520
rect 534 1524 540 1525
rect 534 1520 535 1524
rect 539 1520 540 1524
rect 534 1519 540 1520
rect 560 1508 562 1586
rect 607 1585 611 1586
rect 663 1590 667 1591
rect 663 1585 667 1586
rect 719 1590 723 1591
rect 719 1585 723 1586
rect 727 1590 731 1591
rect 727 1585 731 1586
rect 791 1590 795 1591
rect 791 1585 795 1586
rect 855 1590 859 1591
rect 855 1585 859 1586
rect 1095 1590 1099 1591
rect 1095 1585 1099 1586
rect 570 1583 576 1584
rect 570 1579 571 1583
rect 575 1579 576 1583
rect 570 1578 576 1579
rect 572 1560 574 1578
rect 608 1573 610 1585
rect 634 1583 640 1584
rect 634 1579 635 1583
rect 639 1579 640 1583
rect 634 1578 640 1579
rect 606 1572 612 1573
rect 606 1568 607 1572
rect 611 1568 612 1572
rect 606 1567 612 1568
rect 636 1560 638 1578
rect 664 1573 666 1585
rect 690 1583 696 1584
rect 690 1579 691 1583
rect 695 1579 696 1583
rect 690 1578 696 1579
rect 662 1572 668 1573
rect 662 1568 663 1572
rect 667 1568 668 1572
rect 662 1567 668 1568
rect 692 1560 694 1578
rect 728 1573 730 1585
rect 754 1583 760 1584
rect 754 1579 755 1583
rect 759 1579 760 1583
rect 754 1578 760 1579
rect 726 1572 732 1573
rect 726 1568 727 1572
rect 731 1568 732 1572
rect 726 1567 732 1568
rect 756 1560 758 1578
rect 792 1573 794 1585
rect 818 1583 824 1584
rect 818 1579 819 1583
rect 823 1579 824 1583
rect 818 1578 824 1579
rect 790 1572 796 1573
rect 790 1568 791 1572
rect 795 1568 796 1572
rect 790 1567 796 1568
rect 820 1560 822 1578
rect 856 1573 858 1585
rect 854 1572 860 1573
rect 854 1568 855 1572
rect 859 1568 860 1572
rect 854 1567 860 1568
rect 1096 1565 1098 1585
rect 1136 1575 1138 1595
rect 1158 1592 1164 1593
rect 1158 1588 1159 1592
rect 1163 1588 1164 1592
rect 1158 1587 1164 1588
rect 1160 1575 1162 1587
rect 1180 1580 1182 1622
rect 1188 1612 1190 1670
rect 1196 1652 1198 1670
rect 1248 1665 1250 1677
rect 1274 1675 1280 1676
rect 1274 1671 1275 1675
rect 1279 1671 1280 1675
rect 1274 1670 1280 1671
rect 1246 1664 1252 1665
rect 1246 1660 1247 1664
rect 1251 1660 1252 1664
rect 1246 1659 1252 1660
rect 1276 1652 1278 1670
rect 1304 1656 1306 1682
rect 1319 1677 1323 1678
rect 1335 1682 1339 1683
rect 1374 1682 1380 1683
rect 1383 1682 1387 1683
rect 1335 1677 1339 1678
rect 1383 1677 1387 1678
rect 1423 1682 1427 1683
rect 1446 1682 1452 1683
rect 1455 1682 1459 1683
rect 1423 1677 1427 1678
rect 1455 1677 1459 1678
rect 1511 1682 1515 1683
rect 1526 1682 1532 1683
rect 1535 1682 1539 1683
rect 1511 1677 1515 1678
rect 1535 1677 1539 1678
rect 1599 1682 1603 1683
rect 1606 1682 1612 1683
rect 1615 1682 1619 1683
rect 1599 1677 1603 1678
rect 1615 1677 1619 1678
rect 1679 1682 1683 1683
rect 1679 1677 1683 1678
rect 1687 1682 1691 1683
rect 1710 1682 1716 1683
rect 1742 1687 1748 1688
rect 1742 1683 1743 1687
rect 1747 1683 1748 1687
rect 1760 1683 1762 1695
rect 1742 1682 1748 1683
rect 1751 1682 1755 1683
rect 1687 1677 1691 1678
rect 1751 1677 1755 1678
rect 1759 1682 1763 1683
rect 1759 1677 1763 1678
rect 1336 1665 1338 1677
rect 1362 1675 1368 1676
rect 1362 1671 1363 1675
rect 1367 1671 1368 1675
rect 1362 1670 1368 1671
rect 1334 1664 1340 1665
rect 1334 1660 1335 1664
rect 1339 1660 1340 1664
rect 1334 1659 1340 1660
rect 1302 1655 1308 1656
rect 1194 1651 1200 1652
rect 1194 1647 1195 1651
rect 1199 1647 1200 1651
rect 1194 1646 1200 1647
rect 1274 1651 1280 1652
rect 1274 1647 1275 1651
rect 1279 1647 1280 1651
rect 1302 1651 1303 1655
rect 1307 1651 1308 1655
rect 1364 1652 1366 1670
rect 1424 1665 1426 1677
rect 1512 1665 1514 1677
rect 1600 1665 1602 1677
rect 1626 1675 1632 1676
rect 1618 1671 1624 1672
rect 1618 1667 1619 1671
rect 1623 1667 1624 1671
rect 1626 1671 1627 1675
rect 1631 1671 1632 1675
rect 1626 1670 1632 1671
rect 1618 1666 1624 1667
rect 1422 1664 1428 1665
rect 1422 1660 1423 1664
rect 1427 1660 1428 1664
rect 1422 1659 1428 1660
rect 1510 1664 1516 1665
rect 1510 1660 1511 1664
rect 1515 1660 1516 1664
rect 1510 1659 1516 1660
rect 1598 1664 1604 1665
rect 1598 1660 1599 1664
rect 1603 1660 1604 1664
rect 1598 1659 1604 1660
rect 1302 1650 1308 1651
rect 1362 1651 1368 1652
rect 1274 1646 1280 1647
rect 1362 1647 1363 1651
rect 1367 1647 1368 1651
rect 1362 1646 1368 1647
rect 1246 1636 1252 1637
rect 1246 1632 1247 1636
rect 1251 1632 1252 1636
rect 1246 1631 1252 1632
rect 1334 1636 1340 1637
rect 1334 1632 1335 1636
rect 1339 1632 1340 1636
rect 1334 1631 1340 1632
rect 1422 1636 1428 1637
rect 1422 1632 1423 1636
rect 1427 1632 1428 1636
rect 1422 1631 1428 1632
rect 1510 1636 1516 1637
rect 1510 1632 1511 1636
rect 1515 1632 1516 1636
rect 1510 1631 1516 1632
rect 1598 1636 1604 1637
rect 1598 1632 1599 1636
rect 1603 1632 1604 1636
rect 1598 1631 1604 1632
rect 1248 1627 1250 1631
rect 1336 1627 1338 1631
rect 1424 1627 1426 1631
rect 1470 1627 1476 1628
rect 1512 1627 1514 1631
rect 1600 1627 1602 1631
rect 1620 1628 1622 1666
rect 1628 1652 1630 1670
rect 1680 1665 1682 1677
rect 1752 1665 1754 1677
rect 1808 1676 1810 1706
rect 1830 1700 1836 1701
rect 1830 1696 1831 1700
rect 1835 1696 1836 1700
rect 1830 1695 1836 1696
rect 1894 1700 1900 1701
rect 1894 1696 1895 1700
rect 1899 1696 1900 1700
rect 1894 1695 1900 1696
rect 1958 1700 1964 1701
rect 1958 1696 1959 1700
rect 1963 1696 1964 1700
rect 1958 1695 1964 1696
rect 2022 1700 2028 1701
rect 2022 1696 2023 1700
rect 2027 1696 2028 1700
rect 2022 1695 2028 1696
rect 2070 1700 2076 1701
rect 2070 1696 2071 1700
rect 2075 1696 2076 1700
rect 2070 1695 2076 1696
rect 1832 1683 1834 1695
rect 1896 1683 1898 1695
rect 1960 1683 1962 1695
rect 2010 1687 2016 1688
rect 2010 1683 2011 1687
rect 2015 1683 2016 1687
rect 2024 1683 2026 1695
rect 2072 1683 2074 1695
rect 1815 1682 1819 1683
rect 1815 1677 1819 1678
rect 1831 1682 1835 1683
rect 1831 1677 1835 1678
rect 1871 1682 1875 1683
rect 1871 1677 1875 1678
rect 1895 1682 1899 1683
rect 1895 1677 1899 1678
rect 1927 1682 1931 1683
rect 1927 1677 1931 1678
rect 1959 1682 1963 1683
rect 1959 1677 1963 1678
rect 1983 1682 1987 1683
rect 2010 1682 2016 1683
rect 2023 1682 2027 1683
rect 1983 1677 1987 1678
rect 1798 1675 1804 1676
rect 1798 1671 1799 1675
rect 1803 1671 1804 1675
rect 1798 1670 1804 1671
rect 1806 1675 1812 1676
rect 1806 1671 1807 1675
rect 1811 1671 1812 1675
rect 1806 1670 1812 1671
rect 1678 1664 1684 1665
rect 1678 1660 1679 1664
rect 1683 1660 1684 1664
rect 1678 1659 1684 1660
rect 1750 1664 1756 1665
rect 1750 1660 1751 1664
rect 1755 1660 1756 1664
rect 1750 1659 1756 1660
rect 1800 1652 1802 1670
rect 1816 1665 1818 1677
rect 1872 1665 1874 1677
rect 1906 1675 1912 1676
rect 1906 1671 1907 1675
rect 1911 1671 1912 1675
rect 1906 1670 1912 1671
rect 1814 1664 1820 1665
rect 1814 1660 1815 1664
rect 1819 1660 1820 1664
rect 1814 1659 1820 1660
rect 1870 1664 1876 1665
rect 1870 1660 1871 1664
rect 1875 1660 1876 1664
rect 1870 1659 1876 1660
rect 1908 1652 1910 1670
rect 1928 1665 1930 1677
rect 1984 1665 1986 1677
rect 1926 1664 1932 1665
rect 1926 1660 1927 1664
rect 1931 1660 1932 1664
rect 1926 1659 1932 1660
rect 1982 1664 1988 1665
rect 1982 1660 1983 1664
rect 1987 1660 1988 1664
rect 1982 1659 1988 1660
rect 2012 1652 2014 1682
rect 2023 1677 2027 1678
rect 2031 1682 2035 1683
rect 2031 1677 2035 1678
rect 2071 1682 2075 1683
rect 2071 1677 2075 1678
rect 2032 1665 2034 1677
rect 2072 1665 2074 1677
rect 2084 1676 2086 1706
rect 2092 1688 2094 1754
rect 2118 1747 2124 1748
rect 2118 1743 2119 1747
rect 2123 1743 2124 1747
rect 2118 1742 2124 1743
rect 2120 1735 2122 1742
rect 2119 1734 2123 1735
rect 2119 1729 2123 1730
rect 2120 1726 2122 1729
rect 2118 1725 2124 1726
rect 2118 1721 2119 1725
rect 2123 1721 2124 1725
rect 2118 1720 2124 1721
rect 2118 1708 2124 1709
rect 2118 1704 2119 1708
rect 2123 1704 2124 1708
rect 2118 1703 2124 1704
rect 2090 1687 2096 1688
rect 2090 1683 2091 1687
rect 2095 1683 2096 1687
rect 2120 1683 2122 1703
rect 2090 1682 2096 1683
rect 2119 1682 2123 1683
rect 2119 1677 2123 1678
rect 2082 1675 2088 1676
rect 2082 1671 2083 1675
rect 2087 1671 2088 1675
rect 2082 1670 2088 1671
rect 2030 1664 2036 1665
rect 2030 1660 2031 1664
rect 2035 1660 2036 1664
rect 2030 1659 2036 1660
rect 2070 1664 2076 1665
rect 2070 1660 2071 1664
rect 2075 1660 2076 1664
rect 2070 1659 2076 1660
rect 2120 1657 2122 1677
rect 2118 1656 2124 1657
rect 2118 1652 2119 1656
rect 2123 1652 2124 1656
rect 1626 1651 1632 1652
rect 1626 1647 1627 1651
rect 1631 1647 1632 1651
rect 1626 1646 1632 1647
rect 1742 1651 1748 1652
rect 1742 1647 1743 1651
rect 1747 1647 1748 1651
rect 1742 1646 1748 1647
rect 1774 1651 1780 1652
rect 1774 1647 1775 1651
rect 1779 1647 1780 1651
rect 1774 1646 1780 1647
rect 1798 1651 1804 1652
rect 1798 1647 1799 1651
rect 1803 1647 1804 1651
rect 1798 1646 1804 1647
rect 1906 1651 1912 1652
rect 1906 1647 1907 1651
rect 1911 1647 1912 1651
rect 1906 1646 1912 1647
rect 2010 1651 2016 1652
rect 2118 1651 2124 1652
rect 2010 1647 2011 1651
rect 2015 1647 2016 1651
rect 2010 1646 2016 1647
rect 1678 1636 1684 1637
rect 1678 1632 1679 1636
rect 1683 1632 1684 1636
rect 1678 1631 1684 1632
rect 1618 1627 1624 1628
rect 1680 1627 1682 1631
rect 1199 1626 1203 1627
rect 1199 1621 1203 1622
rect 1247 1626 1251 1627
rect 1247 1621 1251 1622
rect 1319 1626 1323 1627
rect 1319 1621 1323 1622
rect 1335 1626 1339 1627
rect 1335 1621 1339 1622
rect 1391 1626 1395 1627
rect 1391 1621 1395 1622
rect 1423 1626 1427 1627
rect 1423 1621 1427 1622
rect 1463 1626 1467 1627
rect 1470 1623 1471 1627
rect 1475 1623 1476 1627
rect 1470 1622 1476 1623
rect 1511 1626 1515 1627
rect 1463 1621 1467 1622
rect 1198 1620 1204 1621
rect 1198 1616 1199 1620
rect 1203 1616 1204 1620
rect 1198 1615 1204 1616
rect 1246 1620 1252 1621
rect 1246 1616 1247 1620
rect 1251 1616 1252 1620
rect 1246 1615 1252 1616
rect 1318 1620 1324 1621
rect 1318 1616 1319 1620
rect 1323 1616 1324 1620
rect 1318 1615 1324 1616
rect 1390 1620 1396 1621
rect 1390 1616 1391 1620
rect 1395 1616 1396 1620
rect 1390 1615 1396 1616
rect 1462 1620 1468 1621
rect 1462 1616 1463 1620
rect 1467 1616 1468 1620
rect 1462 1615 1468 1616
rect 1186 1611 1192 1612
rect 1186 1607 1187 1611
rect 1191 1607 1192 1611
rect 1186 1606 1192 1607
rect 1472 1604 1474 1622
rect 1511 1621 1515 1622
rect 1535 1626 1539 1627
rect 1535 1621 1539 1622
rect 1599 1626 1603 1627
rect 1599 1621 1603 1622
rect 1607 1626 1611 1627
rect 1618 1623 1619 1627
rect 1623 1623 1624 1627
rect 1618 1622 1624 1623
rect 1679 1626 1683 1627
rect 1607 1621 1611 1622
rect 1679 1621 1683 1622
rect 1534 1620 1540 1621
rect 1534 1616 1535 1620
rect 1539 1616 1540 1620
rect 1534 1615 1540 1616
rect 1606 1620 1612 1621
rect 1606 1616 1607 1620
rect 1611 1616 1612 1620
rect 1606 1615 1612 1616
rect 1678 1620 1684 1621
rect 1678 1616 1679 1620
rect 1683 1616 1684 1620
rect 1678 1615 1684 1616
rect 1558 1611 1564 1612
rect 1558 1607 1559 1611
rect 1563 1607 1564 1611
rect 1558 1606 1564 1607
rect 1702 1611 1708 1612
rect 1702 1607 1703 1611
rect 1707 1607 1708 1611
rect 1702 1606 1708 1607
rect 1186 1603 1192 1604
rect 1186 1599 1187 1603
rect 1191 1599 1192 1603
rect 1186 1598 1192 1599
rect 1310 1603 1316 1604
rect 1310 1599 1311 1603
rect 1315 1599 1316 1603
rect 1310 1598 1316 1599
rect 1454 1603 1460 1604
rect 1454 1599 1455 1603
rect 1459 1599 1460 1603
rect 1454 1598 1460 1599
rect 1470 1603 1476 1604
rect 1470 1599 1471 1603
rect 1475 1599 1476 1603
rect 1470 1598 1476 1599
rect 1188 1580 1190 1598
rect 1198 1592 1204 1593
rect 1198 1588 1199 1592
rect 1203 1588 1204 1592
rect 1198 1587 1204 1588
rect 1246 1592 1252 1593
rect 1246 1588 1247 1592
rect 1251 1588 1252 1592
rect 1246 1587 1252 1588
rect 1178 1579 1184 1580
rect 1178 1575 1179 1579
rect 1183 1575 1184 1579
rect 1135 1574 1139 1575
rect 1135 1569 1139 1570
rect 1159 1574 1163 1575
rect 1178 1574 1184 1575
rect 1186 1579 1192 1580
rect 1186 1575 1187 1579
rect 1191 1575 1192 1579
rect 1200 1575 1202 1587
rect 1248 1575 1250 1587
rect 1312 1580 1314 1598
rect 1318 1592 1324 1593
rect 1318 1588 1319 1592
rect 1323 1588 1324 1592
rect 1318 1587 1324 1588
rect 1390 1592 1396 1593
rect 1390 1588 1391 1592
rect 1395 1588 1396 1592
rect 1390 1587 1396 1588
rect 1310 1579 1316 1580
rect 1310 1575 1311 1579
rect 1315 1575 1316 1579
rect 1320 1575 1322 1587
rect 1354 1579 1360 1580
rect 1354 1575 1355 1579
rect 1359 1575 1360 1579
rect 1392 1575 1394 1587
rect 1456 1580 1458 1598
rect 1462 1592 1468 1593
rect 1462 1588 1463 1592
rect 1467 1588 1468 1592
rect 1462 1587 1468 1588
rect 1534 1592 1540 1593
rect 1534 1588 1535 1592
rect 1539 1588 1540 1592
rect 1534 1587 1540 1588
rect 1454 1579 1460 1580
rect 1454 1575 1455 1579
rect 1459 1575 1460 1579
rect 1464 1575 1466 1587
rect 1536 1575 1538 1587
rect 1560 1580 1562 1606
rect 1598 1603 1604 1604
rect 1598 1599 1599 1603
rect 1603 1599 1604 1603
rect 1598 1598 1604 1599
rect 1630 1603 1636 1604
rect 1630 1599 1631 1603
rect 1635 1599 1636 1603
rect 1630 1598 1636 1599
rect 1600 1580 1602 1598
rect 1606 1592 1612 1593
rect 1606 1588 1607 1592
rect 1611 1588 1612 1592
rect 1606 1587 1612 1588
rect 1558 1579 1564 1580
rect 1558 1575 1559 1579
rect 1563 1575 1564 1579
rect 1598 1579 1604 1580
rect 1598 1575 1599 1579
rect 1603 1575 1604 1579
rect 1608 1575 1610 1587
rect 1186 1574 1192 1575
rect 1199 1574 1203 1575
rect 1159 1569 1163 1570
rect 1199 1569 1203 1570
rect 1239 1574 1243 1575
rect 1239 1569 1243 1570
rect 1247 1574 1251 1575
rect 1247 1569 1251 1570
rect 1279 1574 1283 1575
rect 1310 1574 1316 1575
rect 1319 1574 1323 1575
rect 1279 1569 1283 1570
rect 1319 1569 1323 1570
rect 1327 1574 1331 1575
rect 1354 1574 1360 1575
rect 1375 1574 1379 1575
rect 1327 1569 1331 1570
rect 1094 1564 1100 1565
rect 1094 1560 1095 1564
rect 1099 1560 1100 1564
rect 570 1559 576 1560
rect 570 1555 571 1559
rect 575 1555 576 1559
rect 570 1554 576 1555
rect 634 1559 640 1560
rect 634 1555 635 1559
rect 639 1555 640 1559
rect 634 1554 640 1555
rect 690 1559 696 1560
rect 690 1555 691 1559
rect 695 1555 696 1559
rect 690 1554 696 1555
rect 754 1559 760 1560
rect 754 1555 755 1559
rect 759 1555 760 1559
rect 754 1554 760 1555
rect 818 1559 824 1560
rect 818 1555 819 1559
rect 823 1555 824 1559
rect 818 1554 824 1555
rect 838 1559 844 1560
rect 1094 1559 1100 1560
rect 838 1555 839 1559
rect 843 1555 844 1559
rect 838 1554 844 1555
rect 606 1544 612 1545
rect 606 1540 607 1544
rect 611 1540 612 1544
rect 606 1539 612 1540
rect 662 1544 668 1545
rect 662 1540 663 1544
rect 667 1540 668 1544
rect 662 1539 668 1540
rect 726 1544 732 1545
rect 726 1540 727 1544
rect 731 1540 732 1544
rect 726 1539 732 1540
rect 790 1544 796 1545
rect 790 1540 791 1544
rect 795 1540 796 1544
rect 790 1539 796 1540
rect 608 1531 610 1539
rect 664 1531 666 1539
rect 728 1531 730 1539
rect 792 1531 794 1539
rect 575 1530 579 1531
rect 575 1525 579 1526
rect 607 1530 611 1531
rect 607 1525 611 1526
rect 615 1530 619 1531
rect 615 1525 619 1526
rect 655 1530 659 1531
rect 655 1525 659 1526
rect 663 1530 667 1531
rect 663 1525 667 1526
rect 695 1530 699 1531
rect 695 1525 699 1526
rect 727 1530 731 1531
rect 727 1525 731 1526
rect 735 1530 739 1531
rect 735 1525 739 1526
rect 775 1530 779 1531
rect 775 1525 779 1526
rect 791 1530 795 1531
rect 791 1525 795 1526
rect 831 1530 835 1531
rect 831 1525 835 1526
rect 574 1524 580 1525
rect 574 1520 575 1524
rect 579 1520 580 1524
rect 574 1519 580 1520
rect 614 1524 620 1525
rect 614 1520 615 1524
rect 619 1520 620 1524
rect 614 1519 620 1520
rect 654 1524 660 1525
rect 654 1520 655 1524
rect 659 1520 660 1524
rect 654 1519 660 1520
rect 694 1524 700 1525
rect 694 1520 695 1524
rect 699 1520 700 1524
rect 694 1519 700 1520
rect 734 1524 740 1525
rect 734 1520 735 1524
rect 739 1520 740 1524
rect 734 1519 740 1520
rect 774 1524 780 1525
rect 774 1520 775 1524
rect 779 1520 780 1524
rect 774 1519 780 1520
rect 830 1524 836 1525
rect 830 1520 831 1524
rect 835 1520 836 1524
rect 830 1519 836 1520
rect 162 1507 168 1508
rect 162 1503 163 1507
rect 167 1503 168 1507
rect 162 1502 168 1503
rect 202 1507 208 1508
rect 202 1503 203 1507
rect 207 1503 208 1507
rect 202 1502 208 1503
rect 242 1507 248 1508
rect 242 1503 243 1507
rect 247 1503 248 1507
rect 242 1502 248 1503
rect 282 1507 288 1508
rect 282 1503 283 1507
rect 287 1503 288 1507
rect 282 1502 288 1503
rect 322 1507 328 1508
rect 322 1503 323 1507
rect 327 1503 328 1507
rect 322 1502 328 1503
rect 362 1507 368 1508
rect 362 1503 363 1507
rect 367 1503 368 1507
rect 362 1502 368 1503
rect 402 1507 408 1508
rect 402 1503 403 1507
rect 407 1503 408 1507
rect 402 1502 408 1503
rect 442 1507 448 1508
rect 442 1503 443 1507
rect 447 1503 448 1507
rect 442 1502 448 1503
rect 482 1507 488 1508
rect 482 1503 483 1507
rect 487 1503 488 1507
rect 482 1502 488 1503
rect 522 1507 528 1508
rect 522 1503 523 1507
rect 527 1503 528 1507
rect 522 1502 528 1503
rect 558 1507 564 1508
rect 558 1503 559 1507
rect 563 1503 564 1507
rect 558 1502 564 1503
rect 602 1507 608 1508
rect 602 1503 603 1507
rect 607 1503 608 1507
rect 602 1502 608 1503
rect 642 1507 648 1508
rect 642 1503 643 1507
rect 647 1503 648 1507
rect 642 1502 648 1503
rect 682 1507 688 1508
rect 682 1503 683 1507
rect 687 1503 688 1507
rect 682 1502 688 1503
rect 722 1507 728 1508
rect 722 1503 723 1507
rect 727 1503 728 1507
rect 722 1502 728 1503
rect 762 1507 768 1508
rect 762 1503 763 1507
rect 767 1503 768 1507
rect 762 1502 768 1503
rect 782 1507 788 1508
rect 782 1503 783 1507
rect 787 1503 788 1507
rect 782 1502 788 1503
rect 164 1484 166 1502
rect 174 1496 180 1497
rect 174 1492 175 1496
rect 179 1492 180 1496
rect 174 1491 180 1492
rect 150 1483 156 1484
rect 150 1479 151 1483
rect 155 1479 156 1483
rect 150 1478 156 1479
rect 162 1483 168 1484
rect 162 1479 163 1483
rect 167 1479 168 1483
rect 162 1478 168 1479
rect 176 1471 178 1491
rect 204 1484 206 1502
rect 214 1496 220 1497
rect 214 1492 215 1496
rect 219 1492 220 1496
rect 214 1491 220 1492
rect 202 1483 208 1484
rect 202 1479 203 1483
rect 207 1479 208 1483
rect 202 1478 208 1479
rect 216 1471 218 1491
rect 244 1484 246 1502
rect 254 1496 260 1497
rect 254 1492 255 1496
rect 259 1492 260 1496
rect 254 1491 260 1492
rect 242 1483 248 1484
rect 242 1479 243 1483
rect 247 1479 248 1483
rect 242 1478 248 1479
rect 256 1471 258 1491
rect 284 1484 286 1502
rect 294 1496 300 1497
rect 294 1492 295 1496
rect 299 1492 300 1496
rect 294 1491 300 1492
rect 282 1483 288 1484
rect 282 1479 283 1483
rect 287 1479 288 1483
rect 282 1478 288 1479
rect 296 1471 298 1491
rect 324 1484 326 1502
rect 334 1496 340 1497
rect 334 1492 335 1496
rect 339 1492 340 1496
rect 334 1491 340 1492
rect 322 1483 328 1484
rect 322 1479 323 1483
rect 327 1479 328 1483
rect 322 1478 328 1479
rect 336 1471 338 1491
rect 364 1484 366 1502
rect 374 1496 380 1497
rect 374 1492 375 1496
rect 379 1492 380 1496
rect 374 1491 380 1492
rect 362 1483 368 1484
rect 362 1479 363 1483
rect 367 1479 368 1483
rect 362 1478 368 1479
rect 376 1471 378 1491
rect 404 1484 406 1502
rect 414 1496 420 1497
rect 414 1492 415 1496
rect 419 1492 420 1496
rect 414 1491 420 1492
rect 402 1483 408 1484
rect 402 1479 403 1483
rect 407 1479 408 1483
rect 402 1478 408 1479
rect 416 1471 418 1491
rect 444 1484 446 1502
rect 454 1496 460 1497
rect 454 1492 455 1496
rect 459 1492 460 1496
rect 454 1491 460 1492
rect 442 1483 448 1484
rect 442 1479 443 1483
rect 447 1479 448 1483
rect 442 1478 448 1479
rect 456 1471 458 1491
rect 484 1484 486 1502
rect 494 1496 500 1497
rect 494 1492 495 1496
rect 499 1492 500 1496
rect 494 1491 500 1492
rect 482 1483 488 1484
rect 482 1479 483 1483
rect 487 1479 488 1483
rect 482 1478 488 1479
rect 496 1471 498 1491
rect 524 1484 526 1502
rect 534 1496 540 1497
rect 534 1492 535 1496
rect 539 1492 540 1496
rect 534 1491 540 1492
rect 574 1496 580 1497
rect 574 1492 575 1496
rect 579 1492 580 1496
rect 574 1491 580 1492
rect 522 1483 528 1484
rect 522 1479 523 1483
rect 527 1479 528 1483
rect 522 1478 528 1479
rect 536 1471 538 1491
rect 546 1483 552 1484
rect 546 1479 547 1483
rect 551 1479 552 1483
rect 546 1478 552 1479
rect 111 1470 115 1471
rect 111 1465 115 1466
rect 135 1470 139 1471
rect 135 1465 139 1466
rect 175 1470 179 1471
rect 175 1465 179 1466
rect 215 1470 219 1471
rect 215 1465 219 1466
rect 255 1470 259 1471
rect 255 1465 259 1466
rect 295 1470 299 1471
rect 295 1465 299 1466
rect 335 1470 339 1471
rect 335 1465 339 1466
rect 375 1470 379 1471
rect 375 1465 379 1466
rect 415 1470 419 1471
rect 415 1465 419 1466
rect 455 1470 459 1471
rect 455 1465 459 1466
rect 495 1470 499 1471
rect 495 1465 499 1466
rect 519 1470 523 1471
rect 519 1465 523 1466
rect 535 1470 539 1471
rect 535 1465 539 1466
rect 112 1445 114 1465
rect 520 1453 522 1465
rect 518 1452 524 1453
rect 518 1448 519 1452
rect 523 1448 524 1452
rect 518 1447 524 1448
rect 110 1444 116 1445
rect 110 1440 111 1444
rect 115 1440 116 1444
rect 548 1440 550 1478
rect 576 1471 578 1491
rect 604 1484 606 1502
rect 614 1496 620 1497
rect 614 1492 615 1496
rect 619 1492 620 1496
rect 614 1491 620 1492
rect 602 1483 608 1484
rect 602 1479 603 1483
rect 607 1479 608 1483
rect 602 1478 608 1479
rect 582 1471 588 1472
rect 616 1471 618 1491
rect 644 1484 646 1502
rect 654 1496 660 1497
rect 654 1492 655 1496
rect 659 1492 660 1496
rect 654 1491 660 1492
rect 642 1483 648 1484
rect 642 1479 643 1483
rect 647 1479 648 1483
rect 642 1478 648 1479
rect 656 1471 658 1491
rect 684 1484 686 1502
rect 694 1496 700 1497
rect 694 1492 695 1496
rect 699 1492 700 1496
rect 694 1491 700 1492
rect 682 1483 688 1484
rect 682 1479 683 1483
rect 687 1479 688 1483
rect 682 1478 688 1479
rect 696 1471 698 1491
rect 724 1484 726 1502
rect 734 1496 740 1497
rect 734 1492 735 1496
rect 739 1492 740 1496
rect 734 1491 740 1492
rect 722 1483 728 1484
rect 722 1479 723 1483
rect 727 1479 728 1483
rect 722 1478 728 1479
rect 736 1471 738 1491
rect 764 1484 766 1502
rect 774 1496 780 1497
rect 774 1492 775 1496
rect 779 1492 780 1496
rect 774 1491 780 1492
rect 762 1483 768 1484
rect 762 1479 763 1483
rect 767 1479 768 1483
rect 762 1478 768 1479
rect 776 1471 778 1491
rect 784 1472 786 1502
rect 830 1496 836 1497
rect 830 1492 831 1496
rect 835 1492 836 1496
rect 830 1491 836 1492
rect 782 1471 788 1472
rect 832 1471 834 1491
rect 840 1484 842 1554
rect 1136 1549 1138 1569
rect 1240 1557 1242 1569
rect 1258 1567 1264 1568
rect 1258 1563 1259 1567
rect 1263 1563 1264 1567
rect 1258 1562 1264 1563
rect 1266 1567 1272 1568
rect 1266 1563 1267 1567
rect 1271 1563 1272 1567
rect 1266 1562 1272 1563
rect 1238 1556 1244 1557
rect 1238 1552 1239 1556
rect 1243 1552 1244 1556
rect 1238 1551 1244 1552
rect 1260 1549 1262 1562
rect 1134 1548 1140 1549
rect 1094 1547 1100 1548
rect 854 1544 860 1545
rect 854 1540 855 1544
rect 859 1540 860 1544
rect 1094 1543 1095 1547
rect 1099 1543 1100 1547
rect 1134 1544 1135 1548
rect 1139 1544 1140 1548
rect 1134 1543 1140 1544
rect 1259 1548 1263 1549
rect 1268 1544 1270 1562
rect 1280 1557 1282 1569
rect 1306 1567 1312 1568
rect 1306 1563 1307 1567
rect 1311 1563 1312 1567
rect 1306 1562 1312 1563
rect 1278 1556 1284 1557
rect 1278 1552 1279 1556
rect 1283 1552 1284 1556
rect 1278 1551 1284 1552
rect 1308 1544 1310 1562
rect 1328 1557 1330 1569
rect 1326 1556 1332 1557
rect 1326 1552 1327 1556
rect 1331 1552 1332 1556
rect 1326 1551 1332 1552
rect 1356 1544 1358 1574
rect 1375 1569 1379 1570
rect 1391 1574 1395 1575
rect 1391 1569 1395 1570
rect 1423 1574 1427 1575
rect 1454 1574 1460 1575
rect 1463 1574 1467 1575
rect 1423 1569 1427 1570
rect 1463 1569 1467 1570
rect 1471 1574 1475 1575
rect 1471 1569 1475 1570
rect 1519 1574 1523 1575
rect 1519 1569 1523 1570
rect 1535 1574 1539 1575
rect 1558 1574 1564 1575
rect 1567 1574 1571 1575
rect 1598 1574 1604 1575
rect 1607 1574 1611 1575
rect 1535 1569 1539 1570
rect 1554 1571 1560 1572
rect 1376 1557 1378 1569
rect 1410 1567 1416 1568
rect 1410 1563 1411 1567
rect 1415 1563 1416 1567
rect 1410 1562 1416 1563
rect 1374 1556 1380 1557
rect 1374 1552 1375 1556
rect 1379 1552 1380 1556
rect 1374 1551 1380 1552
rect 1399 1548 1403 1549
rect 1412 1544 1414 1562
rect 1424 1557 1426 1569
rect 1430 1567 1436 1568
rect 1430 1563 1431 1567
rect 1435 1563 1436 1567
rect 1430 1562 1436 1563
rect 1422 1556 1428 1557
rect 1422 1552 1423 1556
rect 1427 1552 1428 1556
rect 1422 1551 1428 1552
rect 1259 1543 1263 1544
rect 1266 1543 1272 1544
rect 1094 1542 1100 1543
rect 854 1539 860 1540
rect 856 1531 858 1539
rect 1096 1531 1098 1542
rect 1266 1539 1267 1543
rect 1271 1539 1272 1543
rect 1266 1538 1272 1539
rect 1306 1543 1312 1544
rect 1306 1539 1307 1543
rect 1311 1539 1312 1543
rect 1306 1538 1312 1539
rect 1354 1543 1360 1544
rect 1354 1539 1355 1543
rect 1359 1539 1360 1543
rect 1354 1538 1360 1539
rect 1398 1543 1404 1544
rect 1398 1539 1399 1543
rect 1403 1539 1404 1543
rect 1398 1538 1404 1539
rect 1410 1543 1416 1544
rect 1410 1539 1411 1543
rect 1415 1539 1416 1543
rect 1410 1538 1416 1539
rect 1134 1531 1140 1532
rect 855 1530 859 1531
rect 855 1525 859 1526
rect 887 1530 891 1531
rect 887 1525 891 1526
rect 1095 1530 1099 1531
rect 1134 1527 1135 1531
rect 1139 1527 1140 1531
rect 1134 1526 1140 1527
rect 1238 1528 1244 1529
rect 1095 1525 1099 1526
rect 886 1524 892 1525
rect 886 1520 887 1524
rect 891 1520 892 1524
rect 1096 1522 1098 1525
rect 886 1519 892 1520
rect 1094 1521 1100 1522
rect 1094 1517 1095 1521
rect 1099 1517 1100 1521
rect 1136 1519 1138 1526
rect 1238 1524 1239 1528
rect 1243 1524 1244 1528
rect 1238 1523 1244 1524
rect 1278 1528 1284 1529
rect 1278 1524 1279 1528
rect 1283 1524 1284 1528
rect 1278 1523 1284 1524
rect 1326 1528 1332 1529
rect 1326 1524 1327 1528
rect 1331 1524 1332 1528
rect 1326 1523 1332 1524
rect 1374 1528 1380 1529
rect 1374 1524 1375 1528
rect 1379 1524 1380 1528
rect 1374 1523 1380 1524
rect 1422 1528 1428 1529
rect 1422 1524 1423 1528
rect 1427 1524 1428 1528
rect 1422 1523 1428 1524
rect 1240 1519 1242 1523
rect 1280 1519 1282 1523
rect 1328 1519 1330 1523
rect 1376 1519 1378 1523
rect 1424 1519 1426 1523
rect 1094 1516 1100 1517
rect 1135 1518 1139 1519
rect 1135 1513 1139 1514
rect 1239 1518 1243 1519
rect 1239 1513 1243 1514
rect 1279 1518 1283 1519
rect 1279 1513 1283 1514
rect 1319 1518 1323 1519
rect 1319 1513 1323 1514
rect 1327 1518 1331 1519
rect 1327 1513 1331 1514
rect 1359 1518 1363 1519
rect 1359 1513 1363 1514
rect 1375 1518 1379 1519
rect 1375 1513 1379 1514
rect 1399 1518 1403 1519
rect 1399 1513 1403 1514
rect 1423 1518 1427 1519
rect 1423 1513 1427 1514
rect 1136 1510 1138 1513
rect 1318 1512 1324 1513
rect 1134 1509 1140 1510
rect 878 1507 884 1508
rect 878 1503 879 1507
rect 883 1503 884 1507
rect 878 1502 884 1503
rect 926 1507 932 1508
rect 926 1503 927 1507
rect 931 1503 932 1507
rect 1134 1505 1135 1509
rect 1139 1505 1140 1509
rect 1318 1508 1319 1512
rect 1323 1508 1324 1512
rect 1318 1507 1324 1508
rect 1358 1512 1364 1513
rect 1358 1508 1359 1512
rect 1363 1508 1364 1512
rect 1358 1507 1364 1508
rect 1398 1512 1404 1513
rect 1398 1508 1399 1512
rect 1403 1508 1404 1512
rect 1398 1507 1404 1508
rect 926 1502 932 1503
rect 1094 1504 1100 1505
rect 1134 1504 1140 1505
rect 1432 1504 1434 1562
rect 1472 1557 1474 1569
rect 1498 1567 1504 1568
rect 1498 1563 1499 1567
rect 1503 1563 1504 1567
rect 1498 1562 1504 1563
rect 1470 1556 1476 1557
rect 1470 1552 1471 1556
rect 1475 1552 1476 1556
rect 1470 1551 1476 1552
rect 1500 1544 1502 1562
rect 1520 1557 1522 1569
rect 1554 1567 1555 1571
rect 1559 1567 1560 1571
rect 1567 1569 1571 1570
rect 1607 1569 1611 1570
rect 1623 1574 1627 1575
rect 1623 1569 1627 1570
rect 1554 1566 1560 1567
rect 1518 1556 1524 1557
rect 1518 1552 1519 1556
rect 1523 1552 1524 1556
rect 1518 1551 1524 1552
rect 1556 1544 1558 1566
rect 1568 1557 1570 1569
rect 1624 1557 1626 1569
rect 1632 1568 1634 1598
rect 1678 1592 1684 1593
rect 1678 1588 1679 1592
rect 1683 1588 1684 1592
rect 1678 1587 1684 1588
rect 1680 1575 1682 1587
rect 1704 1580 1706 1606
rect 1744 1580 1746 1646
rect 1750 1636 1756 1637
rect 1750 1632 1751 1636
rect 1755 1632 1756 1636
rect 1750 1631 1756 1632
rect 1752 1627 1754 1631
rect 1776 1628 1778 1646
rect 2118 1639 2124 1640
rect 1814 1636 1820 1637
rect 1814 1632 1815 1636
rect 1819 1632 1820 1636
rect 1814 1631 1820 1632
rect 1870 1636 1876 1637
rect 1870 1632 1871 1636
rect 1875 1632 1876 1636
rect 1870 1631 1876 1632
rect 1926 1636 1932 1637
rect 1926 1632 1927 1636
rect 1931 1632 1932 1636
rect 1926 1631 1932 1632
rect 1982 1636 1988 1637
rect 1982 1632 1983 1636
rect 1987 1632 1988 1636
rect 1982 1631 1988 1632
rect 2030 1636 2036 1637
rect 2030 1632 2031 1636
rect 2035 1632 2036 1636
rect 2030 1631 2036 1632
rect 2070 1636 2076 1637
rect 2070 1632 2071 1636
rect 2075 1632 2076 1636
rect 2118 1635 2119 1639
rect 2123 1635 2124 1639
rect 2118 1634 2124 1635
rect 2070 1631 2076 1632
rect 1774 1627 1780 1628
rect 1816 1627 1818 1631
rect 1872 1627 1874 1631
rect 1928 1627 1930 1631
rect 1984 1627 1986 1631
rect 2032 1627 2034 1631
rect 2072 1627 2074 1631
rect 2120 1627 2122 1634
rect 1751 1626 1755 1627
rect 1774 1623 1775 1627
rect 1779 1623 1780 1627
rect 1774 1622 1780 1623
rect 1815 1626 1819 1627
rect 1751 1621 1755 1622
rect 1815 1621 1819 1622
rect 1831 1626 1835 1627
rect 1831 1621 1835 1622
rect 1871 1626 1875 1627
rect 1871 1621 1875 1622
rect 1927 1626 1931 1627
rect 1927 1621 1931 1622
rect 1983 1626 1987 1627
rect 1983 1621 1987 1622
rect 2031 1626 2035 1627
rect 2031 1621 2035 1622
rect 2071 1626 2075 1627
rect 2071 1621 2075 1622
rect 2119 1626 2123 1627
rect 2119 1621 2123 1622
rect 1750 1620 1756 1621
rect 1750 1616 1751 1620
rect 1755 1616 1756 1620
rect 1750 1615 1756 1616
rect 1830 1620 1836 1621
rect 1830 1616 1831 1620
rect 1835 1616 1836 1620
rect 2120 1618 2122 1621
rect 1830 1615 1836 1616
rect 2118 1617 2124 1618
rect 2118 1613 2119 1617
rect 2123 1613 2124 1617
rect 2118 1612 2124 1613
rect 1822 1603 1828 1604
rect 1822 1599 1823 1603
rect 1827 1599 1828 1603
rect 1822 1598 1828 1599
rect 2118 1600 2124 1601
rect 1750 1592 1756 1593
rect 1750 1588 1751 1592
rect 1755 1588 1756 1592
rect 1750 1587 1756 1588
rect 1702 1579 1708 1580
rect 1702 1575 1703 1579
rect 1707 1575 1708 1579
rect 1742 1579 1748 1580
rect 1742 1575 1743 1579
rect 1747 1575 1748 1579
rect 1752 1575 1754 1587
rect 1824 1580 1826 1598
rect 2118 1596 2119 1600
rect 2123 1596 2124 1600
rect 2118 1595 2124 1596
rect 1830 1592 1836 1593
rect 1830 1588 1831 1592
rect 1835 1588 1836 1592
rect 1830 1587 1836 1588
rect 1822 1579 1828 1580
rect 1822 1575 1823 1579
rect 1827 1575 1828 1579
rect 1832 1575 1834 1587
rect 2120 1575 2122 1595
rect 1679 1574 1683 1575
rect 1702 1574 1708 1575
rect 1735 1574 1739 1575
rect 1742 1574 1748 1575
rect 1751 1574 1755 1575
rect 1822 1574 1828 1575
rect 1831 1574 1835 1575
rect 1679 1569 1683 1570
rect 1735 1569 1739 1570
rect 1751 1569 1755 1570
rect 1831 1569 1835 1570
rect 2119 1574 2123 1575
rect 2119 1569 2123 1570
rect 1630 1567 1636 1568
rect 1630 1563 1631 1567
rect 1635 1563 1636 1567
rect 1630 1562 1636 1563
rect 1650 1567 1656 1568
rect 1650 1563 1651 1567
rect 1655 1563 1656 1567
rect 1650 1562 1656 1563
rect 1566 1556 1572 1557
rect 1566 1552 1567 1556
rect 1571 1552 1572 1556
rect 1566 1551 1572 1552
rect 1622 1556 1628 1557
rect 1622 1552 1623 1556
rect 1627 1552 1628 1556
rect 1622 1551 1628 1552
rect 1652 1544 1654 1562
rect 1680 1557 1682 1569
rect 1706 1567 1712 1568
rect 1706 1563 1707 1567
rect 1711 1563 1712 1567
rect 1706 1562 1712 1563
rect 1678 1556 1684 1557
rect 1678 1552 1679 1556
rect 1683 1552 1684 1556
rect 1678 1551 1684 1552
rect 1708 1544 1710 1562
rect 1736 1557 1738 1569
rect 1734 1556 1740 1557
rect 1734 1552 1735 1556
rect 1739 1552 1740 1556
rect 1734 1551 1740 1552
rect 2120 1549 2122 1569
rect 2118 1548 2124 1549
rect 2118 1544 2119 1548
rect 2123 1544 2124 1548
rect 1498 1543 1504 1544
rect 1498 1539 1499 1543
rect 1503 1539 1504 1543
rect 1498 1538 1504 1539
rect 1546 1543 1552 1544
rect 1546 1539 1547 1543
rect 1551 1539 1552 1543
rect 1546 1538 1552 1539
rect 1554 1543 1560 1544
rect 1554 1539 1555 1543
rect 1559 1539 1560 1543
rect 1554 1538 1560 1539
rect 1650 1543 1656 1544
rect 1650 1539 1651 1543
rect 1655 1539 1656 1543
rect 1650 1538 1656 1539
rect 1706 1543 1712 1544
rect 2118 1543 2124 1544
rect 1706 1539 1707 1543
rect 1711 1539 1712 1543
rect 1706 1538 1712 1539
rect 1470 1528 1476 1529
rect 1470 1524 1471 1528
rect 1475 1524 1476 1528
rect 1470 1523 1476 1524
rect 1518 1528 1524 1529
rect 1518 1524 1519 1528
rect 1523 1524 1524 1528
rect 1518 1523 1524 1524
rect 1472 1519 1474 1523
rect 1520 1519 1522 1523
rect 1439 1518 1443 1519
rect 1439 1513 1443 1514
rect 1471 1518 1475 1519
rect 1471 1513 1475 1514
rect 1479 1518 1483 1519
rect 1479 1513 1483 1514
rect 1519 1518 1523 1519
rect 1519 1513 1523 1514
rect 1438 1512 1444 1513
rect 1438 1508 1439 1512
rect 1443 1508 1444 1512
rect 1438 1507 1444 1508
rect 1478 1512 1484 1513
rect 1478 1508 1479 1512
rect 1483 1508 1484 1512
rect 1478 1507 1484 1508
rect 1518 1512 1524 1513
rect 1518 1508 1519 1512
rect 1523 1508 1524 1512
rect 1518 1507 1524 1508
rect 880 1484 882 1502
rect 886 1496 892 1497
rect 886 1492 887 1496
rect 891 1492 892 1496
rect 886 1491 892 1492
rect 838 1483 844 1484
rect 838 1479 839 1483
rect 843 1479 844 1483
rect 838 1478 844 1479
rect 878 1483 884 1484
rect 878 1479 879 1483
rect 883 1479 884 1483
rect 878 1478 884 1479
rect 888 1471 890 1491
rect 559 1470 563 1471
rect 559 1465 563 1466
rect 575 1470 579 1471
rect 582 1467 583 1471
rect 587 1467 588 1471
rect 582 1466 588 1467
rect 599 1470 603 1471
rect 575 1465 579 1466
rect 560 1453 562 1465
rect 558 1452 564 1453
rect 558 1448 559 1452
rect 563 1448 564 1452
rect 558 1447 564 1448
rect 584 1440 586 1466
rect 599 1465 603 1466
rect 615 1470 619 1471
rect 615 1465 619 1466
rect 647 1470 651 1471
rect 647 1465 651 1466
rect 655 1470 659 1471
rect 655 1465 659 1466
rect 695 1470 699 1471
rect 695 1465 699 1466
rect 735 1470 739 1471
rect 735 1465 739 1466
rect 751 1470 755 1471
rect 751 1465 755 1466
rect 775 1470 779 1471
rect 782 1467 783 1471
rect 787 1467 788 1471
rect 782 1466 788 1467
rect 807 1470 811 1471
rect 775 1465 779 1466
rect 807 1465 811 1466
rect 831 1470 835 1471
rect 831 1465 835 1466
rect 871 1470 875 1471
rect 871 1465 875 1466
rect 887 1470 891 1471
rect 887 1465 891 1466
rect 600 1453 602 1465
rect 648 1453 650 1465
rect 674 1463 680 1464
rect 654 1459 660 1460
rect 654 1455 655 1459
rect 659 1455 660 1459
rect 674 1459 675 1463
rect 679 1459 680 1463
rect 674 1458 680 1459
rect 654 1454 660 1455
rect 598 1452 604 1453
rect 598 1448 599 1452
rect 603 1448 604 1452
rect 598 1447 604 1448
rect 646 1452 652 1453
rect 646 1448 647 1452
rect 651 1448 652 1452
rect 646 1447 652 1448
rect 110 1439 116 1440
rect 546 1439 552 1440
rect 546 1435 547 1439
rect 551 1435 552 1439
rect 546 1434 552 1435
rect 582 1439 588 1440
rect 582 1435 583 1439
rect 587 1435 588 1439
rect 582 1434 588 1435
rect 110 1427 116 1428
rect 110 1423 111 1427
rect 115 1423 116 1427
rect 110 1422 116 1423
rect 518 1424 524 1425
rect 112 1415 114 1422
rect 518 1420 519 1424
rect 523 1420 524 1424
rect 518 1419 524 1420
rect 558 1424 564 1425
rect 558 1420 559 1424
rect 563 1420 564 1424
rect 558 1419 564 1420
rect 598 1424 604 1425
rect 598 1420 599 1424
rect 603 1420 604 1424
rect 598 1419 604 1420
rect 646 1424 652 1425
rect 646 1420 647 1424
rect 651 1420 652 1424
rect 646 1419 652 1420
rect 520 1415 522 1419
rect 560 1415 562 1419
rect 600 1415 602 1419
rect 648 1415 650 1419
rect 111 1414 115 1415
rect 111 1409 115 1410
rect 431 1414 435 1415
rect 431 1409 435 1410
rect 471 1414 475 1415
rect 471 1409 475 1410
rect 519 1414 523 1415
rect 519 1409 523 1410
rect 559 1414 563 1415
rect 559 1409 563 1410
rect 575 1414 579 1415
rect 575 1409 579 1410
rect 599 1414 603 1415
rect 599 1409 603 1410
rect 631 1414 635 1415
rect 631 1409 635 1410
rect 647 1414 651 1415
rect 647 1409 651 1410
rect 112 1406 114 1409
rect 430 1408 436 1409
rect 110 1405 116 1406
rect 110 1401 111 1405
rect 115 1401 116 1405
rect 430 1404 431 1408
rect 435 1404 436 1408
rect 430 1403 436 1404
rect 470 1408 476 1409
rect 470 1404 471 1408
rect 475 1404 476 1408
rect 470 1403 476 1404
rect 518 1408 524 1409
rect 518 1404 519 1408
rect 523 1404 524 1408
rect 518 1403 524 1404
rect 574 1408 580 1409
rect 574 1404 575 1408
rect 579 1404 580 1408
rect 574 1403 580 1404
rect 630 1408 636 1409
rect 630 1404 631 1408
rect 635 1404 636 1408
rect 630 1403 636 1404
rect 110 1400 116 1401
rect 656 1392 658 1454
rect 676 1440 678 1458
rect 696 1453 698 1465
rect 752 1453 754 1465
rect 786 1463 792 1464
rect 786 1459 787 1463
rect 791 1459 792 1463
rect 786 1458 792 1459
rect 694 1452 700 1453
rect 694 1448 695 1452
rect 699 1448 700 1452
rect 694 1447 700 1448
rect 750 1452 756 1453
rect 750 1448 751 1452
rect 755 1448 756 1452
rect 750 1447 756 1448
rect 788 1444 790 1458
rect 808 1453 810 1465
rect 872 1453 874 1465
rect 928 1464 930 1502
rect 1094 1500 1095 1504
rect 1099 1500 1100 1504
rect 1094 1499 1100 1500
rect 1430 1503 1436 1504
rect 1430 1499 1431 1503
rect 1435 1499 1436 1503
rect 1096 1471 1098 1499
rect 1430 1498 1436 1499
rect 1346 1495 1352 1496
rect 1134 1492 1140 1493
rect 1134 1488 1135 1492
rect 1139 1488 1140 1492
rect 1346 1491 1347 1495
rect 1351 1491 1352 1495
rect 1346 1490 1352 1491
rect 1382 1495 1388 1496
rect 1382 1491 1383 1495
rect 1387 1491 1388 1495
rect 1382 1490 1388 1491
rect 1426 1495 1432 1496
rect 1426 1491 1427 1495
rect 1431 1491 1432 1495
rect 1426 1490 1432 1491
rect 1466 1495 1472 1496
rect 1466 1491 1467 1495
rect 1471 1491 1472 1495
rect 1466 1490 1472 1491
rect 1506 1495 1512 1496
rect 1506 1491 1507 1495
rect 1511 1491 1512 1495
rect 1506 1490 1512 1491
rect 1134 1487 1140 1488
rect 935 1470 939 1471
rect 935 1465 939 1466
rect 1095 1470 1099 1471
rect 1136 1467 1138 1487
rect 1318 1484 1324 1485
rect 1318 1480 1319 1484
rect 1323 1480 1324 1484
rect 1318 1479 1324 1480
rect 1320 1467 1322 1479
rect 1348 1472 1350 1490
rect 1358 1484 1364 1485
rect 1358 1480 1359 1484
rect 1363 1480 1364 1484
rect 1358 1479 1364 1480
rect 1326 1471 1332 1472
rect 1326 1467 1327 1471
rect 1331 1467 1332 1471
rect 1346 1471 1352 1472
rect 1346 1467 1347 1471
rect 1351 1467 1352 1471
rect 1360 1467 1362 1479
rect 1384 1472 1386 1490
rect 1398 1484 1404 1485
rect 1398 1480 1399 1484
rect 1403 1480 1404 1484
rect 1398 1479 1404 1480
rect 1382 1471 1388 1472
rect 1382 1467 1383 1471
rect 1387 1467 1388 1471
rect 1400 1467 1402 1479
rect 1428 1472 1430 1490
rect 1438 1484 1444 1485
rect 1438 1480 1439 1484
rect 1443 1480 1444 1484
rect 1438 1479 1444 1480
rect 1426 1471 1432 1472
rect 1426 1467 1427 1471
rect 1431 1467 1432 1471
rect 1440 1467 1442 1479
rect 1468 1472 1470 1490
rect 1478 1484 1484 1485
rect 1478 1480 1479 1484
rect 1483 1480 1484 1484
rect 1478 1479 1484 1480
rect 1466 1471 1472 1472
rect 1466 1467 1467 1471
rect 1471 1467 1472 1471
rect 1480 1467 1482 1479
rect 1508 1472 1510 1490
rect 1518 1484 1524 1485
rect 1518 1480 1519 1484
rect 1523 1480 1524 1484
rect 1518 1479 1524 1480
rect 1506 1471 1512 1472
rect 1506 1467 1507 1471
rect 1511 1467 1512 1471
rect 1520 1467 1522 1479
rect 1548 1472 1550 1538
rect 2118 1531 2124 1532
rect 1566 1528 1572 1529
rect 1566 1524 1567 1528
rect 1571 1524 1572 1528
rect 1566 1523 1572 1524
rect 1622 1528 1628 1529
rect 1622 1524 1623 1528
rect 1627 1524 1628 1528
rect 1622 1523 1628 1524
rect 1678 1528 1684 1529
rect 1678 1524 1679 1528
rect 1683 1524 1684 1528
rect 1678 1523 1684 1524
rect 1734 1528 1740 1529
rect 1734 1524 1735 1528
rect 1739 1524 1740 1528
rect 2118 1527 2119 1531
rect 2123 1527 2124 1531
rect 2118 1526 2124 1527
rect 1734 1523 1740 1524
rect 1568 1519 1570 1523
rect 1624 1519 1626 1523
rect 1680 1519 1682 1523
rect 1736 1519 1738 1523
rect 2120 1519 2122 1526
rect 1559 1518 1563 1519
rect 1559 1513 1563 1514
rect 1567 1518 1571 1519
rect 1567 1513 1571 1514
rect 1607 1518 1611 1519
rect 1607 1513 1611 1514
rect 1623 1518 1627 1519
rect 1623 1513 1627 1514
rect 1663 1518 1667 1519
rect 1663 1513 1667 1514
rect 1679 1518 1683 1519
rect 1679 1513 1683 1514
rect 1735 1518 1739 1519
rect 1735 1513 1739 1514
rect 1815 1518 1819 1519
rect 1815 1513 1819 1514
rect 1903 1518 1907 1519
rect 1903 1513 1907 1514
rect 1991 1518 1995 1519
rect 1991 1513 1995 1514
rect 2071 1518 2075 1519
rect 2071 1513 2075 1514
rect 2119 1518 2123 1519
rect 2119 1513 2123 1514
rect 1558 1512 1564 1513
rect 1558 1508 1559 1512
rect 1563 1508 1564 1512
rect 1558 1507 1564 1508
rect 1606 1512 1612 1513
rect 1606 1508 1607 1512
rect 1611 1508 1612 1512
rect 1606 1507 1612 1508
rect 1662 1512 1668 1513
rect 1662 1508 1663 1512
rect 1667 1508 1668 1512
rect 1662 1507 1668 1508
rect 1734 1512 1740 1513
rect 1734 1508 1735 1512
rect 1739 1508 1740 1512
rect 1734 1507 1740 1508
rect 1814 1512 1820 1513
rect 1814 1508 1815 1512
rect 1819 1508 1820 1512
rect 1814 1507 1820 1508
rect 1902 1512 1908 1513
rect 1902 1508 1903 1512
rect 1907 1508 1908 1512
rect 1902 1507 1908 1508
rect 1990 1512 1996 1513
rect 1990 1508 1991 1512
rect 1995 1508 1996 1512
rect 1990 1507 1996 1508
rect 2070 1512 2076 1513
rect 2070 1508 2071 1512
rect 2075 1508 2076 1512
rect 2120 1510 2122 1513
rect 2070 1507 2076 1508
rect 2118 1509 2124 1510
rect 2118 1505 2119 1509
rect 2123 1505 2124 1509
rect 2118 1504 2124 1505
rect 1598 1495 1604 1496
rect 1598 1491 1599 1495
rect 1603 1491 1604 1495
rect 1598 1490 1604 1491
rect 1654 1495 1660 1496
rect 1654 1491 1655 1495
rect 1659 1491 1660 1495
rect 1654 1490 1660 1491
rect 1726 1495 1732 1496
rect 1726 1491 1727 1495
rect 1731 1491 1732 1495
rect 1726 1490 1732 1491
rect 1910 1495 1916 1496
rect 1910 1491 1911 1495
rect 1915 1491 1916 1495
rect 1910 1490 1916 1491
rect 2062 1495 2068 1496
rect 2062 1491 2063 1495
rect 2067 1491 2068 1495
rect 2062 1490 2068 1491
rect 2078 1495 2084 1496
rect 2078 1491 2079 1495
rect 2083 1491 2084 1495
rect 2078 1490 2084 1491
rect 2118 1492 2124 1493
rect 1558 1484 1564 1485
rect 1558 1480 1559 1484
rect 1563 1480 1564 1484
rect 1558 1479 1564 1480
rect 1546 1471 1552 1472
rect 1546 1467 1547 1471
rect 1551 1467 1552 1471
rect 1560 1467 1562 1479
rect 1591 1476 1595 1477
rect 1600 1472 1602 1490
rect 1606 1484 1612 1485
rect 1606 1480 1607 1484
rect 1611 1480 1612 1484
rect 1606 1479 1612 1480
rect 1591 1471 1595 1472
rect 1598 1471 1604 1472
rect 1095 1465 1099 1466
rect 1135 1466 1139 1467
rect 918 1463 924 1464
rect 918 1459 919 1463
rect 923 1459 924 1463
rect 918 1458 924 1459
rect 926 1463 932 1464
rect 926 1459 927 1463
rect 931 1459 932 1463
rect 926 1458 932 1459
rect 806 1452 812 1453
rect 806 1448 807 1452
rect 811 1448 812 1452
rect 806 1447 812 1448
rect 870 1452 876 1453
rect 870 1448 871 1452
rect 875 1448 876 1452
rect 870 1447 876 1448
rect 786 1443 792 1444
rect 674 1439 680 1440
rect 674 1435 675 1439
rect 679 1435 680 1439
rect 786 1439 787 1443
rect 791 1439 792 1443
rect 920 1440 922 1458
rect 936 1453 938 1465
rect 934 1452 940 1453
rect 934 1448 935 1452
rect 939 1448 940 1452
rect 934 1447 940 1448
rect 1096 1445 1098 1465
rect 1135 1461 1139 1462
rect 1231 1466 1235 1467
rect 1231 1461 1235 1462
rect 1279 1466 1283 1467
rect 1279 1461 1283 1462
rect 1319 1466 1323 1467
rect 1326 1466 1332 1467
rect 1335 1466 1339 1467
rect 1346 1466 1352 1467
rect 1359 1466 1363 1467
rect 1382 1466 1388 1467
rect 1391 1466 1395 1467
rect 1319 1461 1323 1462
rect 1094 1444 1100 1445
rect 1094 1440 1095 1444
rect 1099 1440 1100 1444
rect 1136 1441 1138 1461
rect 1232 1449 1234 1461
rect 1250 1459 1256 1460
rect 1250 1455 1251 1459
rect 1255 1455 1256 1459
rect 1250 1454 1256 1455
rect 1258 1459 1264 1460
rect 1258 1455 1259 1459
rect 1263 1455 1264 1459
rect 1258 1454 1264 1455
rect 1230 1448 1236 1449
rect 1230 1444 1231 1448
rect 1235 1444 1236 1448
rect 1230 1443 1236 1444
rect 786 1438 792 1439
rect 830 1439 836 1440
rect 674 1434 680 1435
rect 830 1435 831 1439
rect 835 1435 836 1439
rect 830 1434 836 1435
rect 886 1439 892 1440
rect 886 1435 887 1439
rect 891 1435 892 1439
rect 886 1434 892 1435
rect 918 1439 924 1440
rect 1094 1439 1100 1440
rect 1134 1440 1140 1441
rect 918 1435 919 1439
rect 923 1435 924 1439
rect 1134 1436 1135 1440
rect 1139 1436 1140 1440
rect 1134 1435 1140 1436
rect 918 1434 924 1435
rect 694 1424 700 1425
rect 694 1420 695 1424
rect 699 1420 700 1424
rect 694 1419 700 1420
rect 750 1424 756 1425
rect 750 1420 751 1424
rect 755 1420 756 1424
rect 750 1419 756 1420
rect 806 1424 812 1425
rect 806 1420 807 1424
rect 811 1420 812 1424
rect 806 1419 812 1420
rect 696 1415 698 1419
rect 752 1415 754 1419
rect 808 1415 810 1419
rect 695 1414 699 1415
rect 695 1409 699 1410
rect 751 1414 755 1415
rect 751 1409 755 1410
rect 759 1414 763 1415
rect 759 1409 763 1410
rect 807 1414 811 1415
rect 807 1409 811 1410
rect 823 1414 827 1415
rect 823 1409 827 1410
rect 694 1408 700 1409
rect 694 1404 695 1408
rect 699 1404 700 1408
rect 694 1403 700 1404
rect 758 1408 764 1409
rect 758 1404 759 1408
rect 763 1404 764 1408
rect 758 1403 764 1404
rect 822 1408 828 1409
rect 822 1404 823 1408
rect 827 1404 828 1408
rect 822 1403 828 1404
rect 458 1391 464 1392
rect 110 1388 116 1389
rect 110 1384 111 1388
rect 115 1384 116 1388
rect 458 1387 459 1391
rect 463 1387 464 1391
rect 458 1386 464 1387
rect 510 1391 516 1392
rect 510 1387 511 1391
rect 515 1387 516 1391
rect 510 1386 516 1387
rect 566 1391 572 1392
rect 566 1387 567 1391
rect 571 1387 572 1391
rect 566 1386 572 1387
rect 622 1391 628 1392
rect 622 1387 623 1391
rect 627 1387 628 1391
rect 622 1386 628 1387
rect 654 1391 660 1392
rect 654 1387 655 1391
rect 659 1387 660 1391
rect 654 1386 660 1387
rect 702 1391 708 1392
rect 702 1387 703 1391
rect 707 1387 708 1391
rect 702 1386 708 1387
rect 110 1383 116 1384
rect 112 1363 114 1383
rect 430 1380 436 1381
rect 430 1376 431 1380
rect 435 1376 436 1380
rect 430 1375 436 1376
rect 432 1363 434 1375
rect 460 1368 462 1386
rect 470 1380 476 1381
rect 470 1376 471 1380
rect 475 1376 476 1380
rect 470 1375 476 1376
rect 442 1367 448 1368
rect 442 1363 443 1367
rect 447 1363 448 1367
rect 111 1362 115 1363
rect 111 1357 115 1358
rect 375 1362 379 1363
rect 375 1357 379 1358
rect 423 1362 427 1363
rect 423 1357 427 1358
rect 431 1362 435 1363
rect 442 1362 448 1363
rect 458 1367 464 1368
rect 458 1363 459 1367
rect 463 1363 464 1367
rect 472 1363 474 1375
rect 512 1368 514 1386
rect 518 1380 524 1381
rect 518 1376 519 1380
rect 523 1376 524 1380
rect 518 1375 524 1376
rect 510 1367 516 1368
rect 510 1363 511 1367
rect 515 1363 516 1367
rect 520 1363 522 1375
rect 568 1368 570 1386
rect 574 1380 580 1381
rect 574 1376 575 1380
rect 579 1376 580 1380
rect 574 1375 580 1376
rect 566 1367 572 1368
rect 566 1363 567 1367
rect 571 1363 572 1367
rect 576 1363 578 1375
rect 624 1368 626 1386
rect 630 1380 636 1381
rect 630 1376 631 1380
rect 635 1376 636 1380
rect 630 1375 636 1376
rect 694 1380 700 1381
rect 694 1376 695 1380
rect 699 1376 700 1380
rect 694 1375 700 1376
rect 622 1367 628 1368
rect 622 1363 623 1367
rect 627 1363 628 1367
rect 632 1363 634 1375
rect 696 1363 698 1375
rect 458 1362 464 1363
rect 471 1362 475 1363
rect 431 1357 435 1358
rect 112 1337 114 1357
rect 376 1345 378 1357
rect 382 1355 388 1356
rect 382 1351 383 1355
rect 387 1351 388 1355
rect 382 1350 388 1351
rect 402 1355 408 1356
rect 402 1351 403 1355
rect 407 1351 408 1355
rect 402 1350 408 1351
rect 374 1344 380 1345
rect 374 1340 375 1344
rect 379 1340 380 1344
rect 374 1339 380 1340
rect 110 1336 116 1337
rect 110 1332 111 1336
rect 115 1332 116 1336
rect 110 1331 116 1332
rect 110 1319 116 1320
rect 110 1315 111 1319
rect 115 1315 116 1319
rect 110 1314 116 1315
rect 374 1316 380 1317
rect 112 1311 114 1314
rect 374 1312 375 1316
rect 379 1312 380 1316
rect 374 1311 380 1312
rect 111 1310 115 1311
rect 111 1305 115 1306
rect 335 1310 339 1311
rect 335 1305 339 1306
rect 375 1310 379 1311
rect 375 1305 379 1306
rect 112 1302 114 1305
rect 334 1304 340 1305
rect 110 1301 116 1302
rect 110 1297 111 1301
rect 115 1297 116 1301
rect 334 1300 335 1304
rect 339 1300 340 1304
rect 334 1299 340 1300
rect 110 1296 116 1297
rect 384 1296 386 1350
rect 404 1332 406 1350
rect 424 1345 426 1357
rect 422 1344 428 1345
rect 422 1340 423 1344
rect 427 1340 428 1344
rect 444 1340 446 1362
rect 471 1357 475 1358
rect 479 1362 483 1363
rect 510 1362 516 1363
rect 519 1362 523 1363
rect 479 1357 483 1358
rect 519 1357 523 1358
rect 543 1362 547 1363
rect 566 1362 572 1363
rect 575 1362 579 1363
rect 543 1357 547 1358
rect 575 1357 579 1358
rect 607 1362 611 1363
rect 622 1362 628 1363
rect 631 1362 635 1363
rect 607 1357 611 1358
rect 631 1357 635 1358
rect 671 1362 675 1363
rect 671 1357 675 1358
rect 695 1362 699 1363
rect 695 1357 699 1358
rect 450 1355 456 1356
rect 450 1351 451 1355
rect 455 1351 456 1355
rect 450 1350 456 1351
rect 422 1339 428 1340
rect 442 1339 448 1340
rect 442 1335 443 1339
rect 447 1335 448 1339
rect 442 1334 448 1335
rect 452 1332 454 1350
rect 480 1345 482 1357
rect 506 1355 512 1356
rect 506 1351 507 1355
rect 511 1351 512 1355
rect 506 1350 512 1351
rect 478 1344 484 1345
rect 478 1340 479 1344
rect 483 1340 484 1344
rect 478 1339 484 1340
rect 508 1332 510 1350
rect 544 1345 546 1357
rect 586 1355 592 1356
rect 586 1351 587 1355
rect 591 1351 592 1355
rect 586 1350 592 1351
rect 542 1344 548 1345
rect 542 1340 543 1344
rect 547 1340 548 1344
rect 542 1339 548 1340
rect 588 1332 590 1350
rect 608 1345 610 1357
rect 672 1345 674 1357
rect 704 1356 706 1386
rect 758 1380 764 1381
rect 758 1376 759 1380
rect 763 1376 764 1380
rect 758 1375 764 1376
rect 822 1380 828 1381
rect 822 1376 823 1380
rect 827 1376 828 1380
rect 822 1375 828 1376
rect 760 1363 762 1375
rect 824 1363 826 1375
rect 832 1368 834 1434
rect 870 1424 876 1425
rect 870 1420 871 1424
rect 875 1420 876 1424
rect 870 1419 876 1420
rect 872 1415 874 1419
rect 871 1414 875 1415
rect 871 1409 875 1410
rect 888 1368 890 1434
rect 1094 1427 1100 1428
rect 934 1424 940 1425
rect 934 1420 935 1424
rect 939 1420 940 1424
rect 1094 1423 1095 1427
rect 1099 1423 1100 1427
rect 1094 1422 1100 1423
rect 1134 1423 1140 1424
rect 934 1419 940 1420
rect 936 1415 938 1419
rect 1096 1415 1098 1422
rect 1134 1419 1135 1423
rect 1139 1419 1140 1423
rect 1134 1418 1140 1419
rect 1230 1420 1236 1421
rect 895 1414 899 1415
rect 895 1409 899 1410
rect 935 1414 939 1415
rect 935 1409 939 1410
rect 967 1414 971 1415
rect 967 1409 971 1410
rect 1095 1414 1099 1415
rect 1136 1411 1138 1418
rect 1230 1416 1231 1420
rect 1235 1416 1236 1420
rect 1230 1415 1236 1416
rect 1232 1411 1234 1415
rect 1095 1409 1099 1410
rect 1135 1410 1139 1411
rect 894 1408 900 1409
rect 894 1404 895 1408
rect 899 1404 900 1408
rect 894 1403 900 1404
rect 966 1408 972 1409
rect 966 1404 967 1408
rect 971 1404 972 1408
rect 1096 1406 1098 1409
rect 966 1403 972 1404
rect 1094 1405 1100 1406
rect 1135 1405 1139 1406
rect 1159 1410 1163 1411
rect 1159 1405 1163 1406
rect 1199 1410 1203 1411
rect 1199 1405 1203 1406
rect 1231 1410 1235 1411
rect 1231 1405 1235 1406
rect 1094 1401 1095 1405
rect 1099 1401 1100 1405
rect 1136 1402 1138 1405
rect 1158 1404 1164 1405
rect 1094 1400 1100 1401
rect 1134 1401 1140 1402
rect 1134 1397 1135 1401
rect 1139 1397 1140 1401
rect 1158 1400 1159 1404
rect 1163 1400 1164 1404
rect 1158 1399 1164 1400
rect 1198 1404 1204 1405
rect 1198 1400 1199 1404
rect 1203 1400 1204 1404
rect 1198 1399 1204 1400
rect 1134 1396 1140 1397
rect 1252 1396 1254 1454
rect 1260 1436 1262 1454
rect 1280 1449 1282 1461
rect 1306 1459 1312 1460
rect 1306 1455 1307 1459
rect 1311 1455 1312 1459
rect 1306 1454 1312 1455
rect 1278 1448 1284 1449
rect 1278 1444 1279 1448
rect 1283 1444 1284 1448
rect 1278 1443 1284 1444
rect 1308 1436 1310 1454
rect 1328 1445 1330 1466
rect 1335 1461 1339 1462
rect 1359 1461 1363 1462
rect 1391 1461 1395 1462
rect 1399 1466 1403 1467
rect 1426 1466 1432 1467
rect 1439 1466 1443 1467
rect 1399 1461 1403 1462
rect 1439 1461 1443 1462
rect 1455 1466 1459 1467
rect 1466 1466 1472 1467
rect 1479 1466 1483 1467
rect 1506 1466 1512 1467
rect 1519 1466 1523 1467
rect 1546 1466 1552 1467
rect 1559 1466 1563 1467
rect 1455 1461 1459 1462
rect 1479 1461 1483 1462
rect 1519 1461 1523 1462
rect 1559 1461 1563 1462
rect 1583 1466 1587 1467
rect 1583 1461 1587 1462
rect 1336 1449 1338 1461
rect 1362 1455 1368 1456
rect 1362 1451 1363 1455
rect 1367 1451 1368 1455
rect 1362 1450 1368 1451
rect 1334 1448 1340 1449
rect 1327 1444 1331 1445
rect 1334 1444 1335 1448
rect 1339 1444 1340 1448
rect 1334 1443 1340 1444
rect 1327 1439 1331 1440
rect 1364 1436 1366 1450
rect 1392 1449 1394 1461
rect 1418 1459 1424 1460
rect 1418 1455 1419 1459
rect 1423 1455 1424 1459
rect 1418 1454 1424 1455
rect 1390 1448 1396 1449
rect 1390 1444 1391 1448
rect 1395 1444 1396 1448
rect 1390 1443 1396 1444
rect 1420 1436 1422 1454
rect 1456 1449 1458 1461
rect 1486 1459 1492 1460
rect 1486 1455 1487 1459
rect 1491 1455 1492 1459
rect 1486 1454 1492 1455
rect 1454 1448 1460 1449
rect 1454 1444 1455 1448
rect 1459 1444 1460 1448
rect 1454 1443 1460 1444
rect 1488 1436 1490 1454
rect 1520 1449 1522 1461
rect 1584 1449 1586 1461
rect 1592 1460 1594 1471
rect 1598 1467 1599 1471
rect 1603 1467 1604 1471
rect 1608 1467 1610 1479
rect 1656 1472 1658 1490
rect 1662 1484 1668 1485
rect 1662 1480 1663 1484
rect 1667 1480 1668 1484
rect 1662 1479 1668 1480
rect 1654 1471 1660 1472
rect 1654 1467 1655 1471
rect 1659 1467 1660 1471
rect 1664 1467 1666 1479
rect 1728 1472 1730 1490
rect 1734 1484 1740 1485
rect 1734 1480 1735 1484
rect 1739 1480 1740 1484
rect 1734 1479 1740 1480
rect 1814 1484 1820 1485
rect 1814 1480 1815 1484
rect 1819 1480 1820 1484
rect 1814 1479 1820 1480
rect 1902 1484 1908 1485
rect 1902 1480 1903 1484
rect 1907 1480 1908 1484
rect 1902 1479 1908 1480
rect 1726 1471 1732 1472
rect 1726 1467 1727 1471
rect 1731 1467 1732 1471
rect 1736 1467 1738 1479
rect 1816 1467 1818 1479
rect 1904 1467 1906 1479
rect 1912 1477 1914 1490
rect 1990 1484 1996 1485
rect 1990 1480 1991 1484
rect 1995 1480 1996 1484
rect 1990 1479 1996 1480
rect 1911 1476 1915 1477
rect 1911 1471 1915 1472
rect 1992 1467 1994 1479
rect 2064 1472 2066 1490
rect 2070 1484 2076 1485
rect 2070 1480 2071 1484
rect 2075 1480 2076 1484
rect 2070 1479 2076 1480
rect 2038 1471 2044 1472
rect 2038 1467 2039 1471
rect 2043 1467 2044 1471
rect 1598 1466 1604 1467
rect 1607 1466 1611 1467
rect 1607 1461 1611 1462
rect 1647 1466 1651 1467
rect 1654 1466 1660 1467
rect 1663 1466 1667 1467
rect 1647 1461 1651 1462
rect 1663 1461 1667 1462
rect 1719 1466 1723 1467
rect 1726 1466 1732 1467
rect 1735 1466 1739 1467
rect 1719 1461 1723 1462
rect 1735 1461 1739 1462
rect 1807 1466 1811 1467
rect 1807 1461 1811 1462
rect 1815 1466 1819 1467
rect 1815 1461 1819 1462
rect 1895 1466 1899 1467
rect 1895 1461 1899 1462
rect 1903 1466 1907 1467
rect 1903 1461 1907 1462
rect 1991 1466 1995 1467
rect 2038 1466 2044 1467
rect 2062 1471 2068 1472
rect 2062 1467 2063 1471
rect 2067 1467 2068 1471
rect 2072 1467 2074 1479
rect 2062 1466 2068 1467
rect 2071 1466 2075 1467
rect 1991 1461 1995 1462
rect 1590 1459 1596 1460
rect 1590 1455 1591 1459
rect 1595 1455 1596 1459
rect 1590 1454 1596 1455
rect 1614 1459 1620 1460
rect 1614 1455 1615 1459
rect 1619 1455 1620 1459
rect 1614 1454 1620 1455
rect 1518 1448 1524 1449
rect 1518 1444 1519 1448
rect 1523 1444 1524 1448
rect 1582 1448 1588 1449
rect 1518 1443 1524 1444
rect 1543 1444 1547 1445
rect 1582 1444 1583 1448
rect 1587 1444 1588 1448
rect 1582 1443 1588 1444
rect 1543 1439 1547 1440
rect 1544 1436 1546 1439
rect 1616 1436 1618 1454
rect 1648 1449 1650 1461
rect 1674 1459 1680 1460
rect 1674 1455 1675 1459
rect 1679 1455 1680 1459
rect 1674 1454 1680 1455
rect 1646 1448 1652 1449
rect 1646 1444 1647 1448
rect 1651 1444 1652 1448
rect 1646 1443 1652 1444
rect 1676 1436 1678 1454
rect 1720 1449 1722 1461
rect 1746 1459 1752 1460
rect 1746 1455 1747 1459
rect 1751 1455 1752 1459
rect 1746 1454 1752 1455
rect 1718 1448 1724 1449
rect 1718 1444 1719 1448
rect 1723 1444 1724 1448
rect 1718 1443 1724 1444
rect 1748 1436 1750 1454
rect 1808 1449 1810 1461
rect 1834 1459 1840 1460
rect 1834 1455 1835 1459
rect 1839 1455 1840 1459
rect 1834 1454 1840 1455
rect 1806 1448 1812 1449
rect 1806 1444 1807 1448
rect 1811 1444 1812 1448
rect 1806 1443 1812 1444
rect 1836 1436 1838 1454
rect 1896 1449 1898 1461
rect 1922 1459 1928 1460
rect 1922 1455 1923 1459
rect 1927 1455 1928 1459
rect 1922 1454 1928 1455
rect 1894 1448 1900 1449
rect 1894 1444 1895 1448
rect 1899 1444 1900 1448
rect 1894 1443 1900 1444
rect 1924 1436 1926 1454
rect 1992 1449 1994 1461
rect 1990 1448 1996 1449
rect 1990 1444 1991 1448
rect 1995 1444 1996 1448
rect 1990 1443 1996 1444
rect 1258 1435 1264 1436
rect 1258 1431 1259 1435
rect 1263 1431 1264 1435
rect 1258 1430 1264 1431
rect 1306 1435 1312 1436
rect 1306 1431 1307 1435
rect 1311 1431 1312 1435
rect 1306 1430 1312 1431
rect 1362 1435 1368 1436
rect 1362 1431 1363 1435
rect 1367 1431 1368 1435
rect 1362 1430 1368 1431
rect 1418 1435 1424 1436
rect 1418 1431 1419 1435
rect 1423 1431 1424 1435
rect 1418 1430 1424 1431
rect 1482 1435 1490 1436
rect 1482 1431 1483 1435
rect 1487 1432 1490 1435
rect 1542 1435 1548 1436
rect 1487 1431 1488 1432
rect 1482 1430 1488 1431
rect 1542 1431 1543 1435
rect 1547 1431 1548 1435
rect 1542 1430 1548 1431
rect 1610 1435 1618 1436
rect 1610 1431 1611 1435
rect 1615 1432 1618 1435
rect 1674 1435 1680 1436
rect 1615 1431 1616 1432
rect 1610 1430 1616 1431
rect 1674 1431 1675 1435
rect 1679 1431 1680 1435
rect 1674 1430 1680 1431
rect 1746 1435 1752 1436
rect 1746 1431 1747 1435
rect 1751 1431 1752 1435
rect 1746 1430 1752 1431
rect 1834 1435 1840 1436
rect 1834 1431 1835 1435
rect 1839 1431 1840 1435
rect 1834 1430 1840 1431
rect 1922 1435 1928 1436
rect 1922 1431 1923 1435
rect 1927 1431 1928 1435
rect 1922 1430 1928 1431
rect 1930 1435 1936 1436
rect 1930 1431 1931 1435
rect 1935 1431 1936 1435
rect 1930 1430 1936 1431
rect 1278 1420 1284 1421
rect 1278 1416 1279 1420
rect 1283 1416 1284 1420
rect 1278 1415 1284 1416
rect 1334 1420 1340 1421
rect 1334 1416 1335 1420
rect 1339 1416 1340 1420
rect 1334 1415 1340 1416
rect 1390 1420 1396 1421
rect 1390 1416 1391 1420
rect 1395 1416 1396 1420
rect 1390 1415 1396 1416
rect 1454 1420 1460 1421
rect 1454 1416 1455 1420
rect 1459 1416 1460 1420
rect 1454 1415 1460 1416
rect 1518 1420 1524 1421
rect 1518 1416 1519 1420
rect 1523 1416 1524 1420
rect 1518 1415 1524 1416
rect 1582 1420 1588 1421
rect 1582 1416 1583 1420
rect 1587 1416 1588 1420
rect 1582 1415 1588 1416
rect 1646 1420 1652 1421
rect 1646 1416 1647 1420
rect 1651 1416 1652 1420
rect 1646 1415 1652 1416
rect 1718 1420 1724 1421
rect 1718 1416 1719 1420
rect 1723 1416 1724 1420
rect 1718 1415 1724 1416
rect 1806 1420 1812 1421
rect 1806 1416 1807 1420
rect 1811 1416 1812 1420
rect 1806 1415 1812 1416
rect 1894 1420 1900 1421
rect 1894 1416 1895 1420
rect 1899 1416 1900 1420
rect 1894 1415 1900 1416
rect 1280 1411 1282 1415
rect 1336 1411 1338 1415
rect 1392 1411 1394 1415
rect 1456 1411 1458 1415
rect 1520 1411 1522 1415
rect 1584 1411 1586 1415
rect 1648 1411 1650 1415
rect 1720 1411 1722 1415
rect 1808 1411 1810 1415
rect 1896 1411 1898 1415
rect 1263 1410 1267 1411
rect 1263 1405 1267 1406
rect 1279 1410 1283 1411
rect 1279 1405 1283 1406
rect 1335 1410 1339 1411
rect 1335 1405 1339 1406
rect 1351 1410 1355 1411
rect 1351 1405 1355 1406
rect 1391 1410 1395 1411
rect 1391 1405 1395 1406
rect 1447 1410 1451 1411
rect 1447 1405 1451 1406
rect 1455 1410 1459 1411
rect 1455 1405 1459 1406
rect 1519 1410 1523 1411
rect 1519 1405 1523 1406
rect 1543 1410 1547 1411
rect 1543 1405 1547 1406
rect 1583 1410 1587 1411
rect 1583 1405 1587 1406
rect 1631 1410 1635 1411
rect 1631 1405 1635 1406
rect 1647 1410 1651 1411
rect 1647 1405 1651 1406
rect 1719 1410 1723 1411
rect 1719 1405 1723 1406
rect 1799 1410 1803 1411
rect 1799 1405 1803 1406
rect 1807 1410 1811 1411
rect 1807 1405 1811 1406
rect 1871 1410 1875 1411
rect 1871 1405 1875 1406
rect 1895 1410 1899 1411
rect 1895 1405 1899 1406
rect 1262 1404 1268 1405
rect 1262 1400 1263 1404
rect 1267 1400 1268 1404
rect 1262 1399 1268 1400
rect 1350 1404 1356 1405
rect 1350 1400 1351 1404
rect 1355 1400 1356 1404
rect 1350 1399 1356 1400
rect 1446 1404 1452 1405
rect 1446 1400 1447 1404
rect 1451 1400 1452 1404
rect 1446 1399 1452 1400
rect 1542 1404 1548 1405
rect 1542 1400 1543 1404
rect 1547 1400 1548 1404
rect 1542 1399 1548 1400
rect 1630 1404 1636 1405
rect 1630 1400 1631 1404
rect 1635 1400 1636 1404
rect 1630 1399 1636 1400
rect 1718 1404 1724 1405
rect 1718 1400 1719 1404
rect 1723 1400 1724 1404
rect 1718 1399 1724 1400
rect 1798 1404 1804 1405
rect 1798 1400 1799 1404
rect 1803 1400 1804 1404
rect 1798 1399 1804 1400
rect 1870 1404 1876 1405
rect 1870 1400 1871 1404
rect 1875 1400 1876 1404
rect 1870 1399 1876 1400
rect 1250 1395 1256 1396
rect 958 1391 964 1392
rect 958 1387 959 1391
rect 963 1387 964 1391
rect 958 1386 964 1387
rect 990 1391 996 1392
rect 990 1387 991 1391
rect 995 1387 996 1391
rect 1250 1391 1251 1395
rect 1255 1391 1256 1395
rect 1250 1390 1256 1391
rect 990 1386 996 1387
rect 1094 1388 1100 1389
rect 894 1380 900 1381
rect 894 1376 895 1380
rect 899 1376 900 1380
rect 894 1375 900 1376
rect 830 1367 836 1368
rect 830 1363 831 1367
rect 835 1363 836 1367
rect 886 1367 892 1368
rect 886 1363 887 1367
rect 891 1363 892 1367
rect 896 1363 898 1375
rect 960 1368 962 1386
rect 966 1380 972 1381
rect 966 1376 967 1380
rect 971 1376 972 1380
rect 966 1375 972 1376
rect 958 1367 964 1368
rect 958 1363 959 1367
rect 963 1363 964 1367
rect 968 1363 970 1375
rect 735 1362 739 1363
rect 735 1357 739 1358
rect 759 1362 763 1363
rect 759 1357 763 1358
rect 799 1362 803 1363
rect 799 1357 803 1358
rect 823 1362 827 1363
rect 830 1362 836 1363
rect 863 1362 867 1363
rect 886 1362 892 1363
rect 895 1362 899 1363
rect 823 1357 827 1358
rect 863 1357 867 1358
rect 895 1357 899 1358
rect 927 1362 931 1363
rect 958 1362 964 1363
rect 967 1362 971 1363
rect 927 1357 931 1358
rect 967 1357 971 1358
rect 702 1355 708 1356
rect 702 1351 703 1355
rect 707 1351 708 1355
rect 702 1350 708 1351
rect 736 1345 738 1357
rect 758 1351 764 1352
rect 758 1347 759 1351
rect 763 1347 764 1351
rect 758 1346 764 1347
rect 606 1344 612 1345
rect 606 1340 607 1344
rect 611 1340 612 1344
rect 606 1339 612 1340
rect 670 1344 676 1345
rect 670 1340 671 1344
rect 675 1340 676 1344
rect 670 1339 676 1340
rect 734 1344 740 1345
rect 734 1340 735 1344
rect 739 1340 740 1344
rect 734 1339 740 1340
rect 760 1332 762 1346
rect 800 1345 802 1357
rect 834 1355 840 1356
rect 834 1351 835 1355
rect 839 1351 840 1355
rect 834 1350 840 1351
rect 798 1344 804 1345
rect 798 1340 799 1344
rect 803 1340 804 1344
rect 798 1339 804 1340
rect 836 1332 838 1350
rect 864 1345 866 1357
rect 928 1345 930 1357
rect 992 1356 994 1386
rect 1094 1384 1095 1388
rect 1099 1384 1100 1388
rect 1186 1387 1192 1388
rect 1094 1383 1100 1384
rect 1134 1384 1140 1385
rect 1096 1363 1098 1383
rect 1134 1380 1135 1384
rect 1139 1380 1140 1384
rect 1186 1383 1187 1387
rect 1191 1383 1192 1387
rect 1186 1382 1192 1383
rect 1254 1387 1260 1388
rect 1254 1383 1255 1387
rect 1259 1383 1260 1387
rect 1254 1382 1260 1383
rect 1342 1387 1348 1388
rect 1342 1383 1343 1387
rect 1347 1383 1348 1387
rect 1342 1382 1348 1383
rect 1438 1387 1444 1388
rect 1438 1383 1439 1387
rect 1443 1383 1444 1387
rect 1438 1382 1444 1383
rect 1534 1387 1540 1388
rect 1534 1383 1535 1387
rect 1539 1383 1540 1387
rect 1534 1382 1540 1383
rect 1710 1387 1716 1388
rect 1710 1383 1711 1387
rect 1715 1383 1716 1387
rect 1710 1382 1716 1383
rect 1790 1387 1796 1388
rect 1790 1383 1791 1387
rect 1795 1383 1796 1387
rect 1790 1382 1796 1383
rect 1862 1387 1868 1388
rect 1862 1383 1863 1387
rect 1867 1383 1868 1387
rect 1862 1382 1868 1383
rect 1886 1387 1892 1388
rect 1886 1383 1887 1387
rect 1891 1383 1892 1387
rect 1886 1382 1892 1383
rect 1134 1379 1140 1380
rect 999 1362 1003 1363
rect 999 1357 1003 1358
rect 1047 1362 1051 1363
rect 1047 1357 1051 1358
rect 1095 1362 1099 1363
rect 1095 1357 1099 1358
rect 982 1355 988 1356
rect 982 1351 983 1355
rect 987 1351 988 1355
rect 982 1350 988 1351
rect 990 1355 996 1356
rect 990 1351 991 1355
rect 995 1351 996 1355
rect 990 1350 996 1351
rect 862 1344 868 1345
rect 862 1340 863 1344
rect 867 1340 868 1344
rect 862 1339 868 1340
rect 926 1344 932 1345
rect 926 1340 927 1344
rect 931 1340 932 1344
rect 926 1339 932 1340
rect 984 1332 986 1350
rect 1000 1345 1002 1357
rect 1048 1345 1050 1357
rect 1070 1355 1076 1356
rect 1070 1351 1071 1355
rect 1075 1351 1076 1355
rect 1070 1350 1076 1351
rect 998 1344 1004 1345
rect 998 1340 999 1344
rect 1003 1340 1004 1344
rect 998 1339 1004 1340
rect 1046 1344 1052 1345
rect 1046 1340 1047 1344
rect 1051 1340 1052 1344
rect 1046 1339 1052 1340
rect 402 1331 408 1332
rect 402 1327 403 1331
rect 407 1327 408 1331
rect 402 1326 408 1327
rect 450 1331 456 1332
rect 450 1327 451 1331
rect 455 1327 456 1331
rect 450 1326 456 1327
rect 506 1331 512 1332
rect 506 1327 507 1331
rect 511 1327 512 1331
rect 506 1326 512 1327
rect 586 1331 592 1332
rect 586 1327 587 1331
rect 591 1327 592 1331
rect 586 1326 592 1327
rect 758 1331 764 1332
rect 758 1327 759 1331
rect 763 1327 764 1331
rect 758 1326 764 1327
rect 834 1331 840 1332
rect 834 1327 835 1331
rect 839 1327 840 1331
rect 834 1326 840 1327
rect 842 1331 848 1332
rect 842 1327 843 1331
rect 847 1327 848 1331
rect 842 1326 848 1327
rect 974 1331 980 1332
rect 974 1327 975 1331
rect 979 1327 980 1331
rect 974 1326 980 1327
rect 982 1331 988 1332
rect 982 1327 983 1331
rect 987 1327 988 1331
rect 982 1326 988 1327
rect 422 1316 428 1317
rect 422 1312 423 1316
rect 427 1312 428 1316
rect 422 1311 428 1312
rect 478 1316 484 1317
rect 478 1312 479 1316
rect 483 1312 484 1316
rect 478 1311 484 1312
rect 542 1316 548 1317
rect 542 1312 543 1316
rect 547 1312 548 1316
rect 542 1311 548 1312
rect 606 1316 612 1317
rect 606 1312 607 1316
rect 611 1312 612 1316
rect 606 1311 612 1312
rect 670 1316 676 1317
rect 670 1312 671 1316
rect 675 1312 676 1316
rect 670 1311 676 1312
rect 734 1316 740 1317
rect 734 1312 735 1316
rect 739 1312 740 1316
rect 734 1311 740 1312
rect 798 1316 804 1317
rect 798 1312 799 1316
rect 803 1312 804 1316
rect 798 1311 804 1312
rect 391 1310 395 1311
rect 391 1305 395 1306
rect 423 1310 427 1311
rect 423 1305 427 1306
rect 455 1310 459 1311
rect 455 1305 459 1306
rect 479 1310 483 1311
rect 479 1305 483 1306
rect 527 1310 531 1311
rect 527 1305 531 1306
rect 543 1310 547 1311
rect 543 1305 547 1306
rect 599 1310 603 1311
rect 599 1305 603 1306
rect 607 1310 611 1311
rect 607 1305 611 1306
rect 671 1310 675 1311
rect 671 1305 675 1306
rect 735 1310 739 1311
rect 735 1305 739 1306
rect 743 1310 747 1311
rect 743 1305 747 1306
rect 799 1310 803 1311
rect 799 1305 803 1306
rect 823 1310 827 1311
rect 823 1305 827 1306
rect 390 1304 396 1305
rect 390 1300 391 1304
rect 395 1300 396 1304
rect 390 1299 396 1300
rect 454 1304 460 1305
rect 454 1300 455 1304
rect 459 1300 460 1304
rect 454 1299 460 1300
rect 526 1304 532 1305
rect 526 1300 527 1304
rect 531 1300 532 1304
rect 526 1299 532 1300
rect 598 1304 604 1305
rect 598 1300 599 1304
rect 603 1300 604 1304
rect 598 1299 604 1300
rect 670 1304 676 1305
rect 670 1300 671 1304
rect 675 1300 676 1304
rect 670 1299 676 1300
rect 742 1304 748 1305
rect 742 1300 743 1304
rect 747 1300 748 1304
rect 742 1299 748 1300
rect 822 1304 828 1305
rect 822 1300 823 1304
rect 827 1300 828 1304
rect 822 1299 828 1300
rect 382 1295 388 1296
rect 382 1291 383 1295
rect 387 1291 388 1295
rect 382 1290 388 1291
rect 382 1287 388 1288
rect 110 1284 116 1285
rect 110 1280 111 1284
rect 115 1280 116 1284
rect 382 1283 383 1287
rect 387 1283 388 1287
rect 382 1282 388 1283
rect 446 1287 452 1288
rect 446 1283 447 1287
rect 451 1283 452 1287
rect 446 1282 452 1283
rect 518 1287 524 1288
rect 518 1283 519 1287
rect 523 1283 524 1287
rect 518 1282 524 1283
rect 590 1287 596 1288
rect 590 1283 591 1287
rect 595 1283 596 1287
rect 590 1282 596 1283
rect 734 1287 740 1288
rect 734 1283 735 1287
rect 739 1283 740 1287
rect 734 1282 740 1283
rect 790 1287 796 1288
rect 790 1283 791 1287
rect 795 1283 796 1287
rect 790 1282 796 1283
rect 110 1279 116 1280
rect 112 1255 114 1279
rect 334 1276 340 1277
rect 334 1272 335 1276
rect 339 1272 340 1276
rect 334 1271 340 1272
rect 336 1255 338 1271
rect 384 1264 386 1282
rect 390 1276 396 1277
rect 390 1272 391 1276
rect 395 1272 396 1276
rect 390 1271 396 1272
rect 382 1263 388 1264
rect 382 1259 383 1263
rect 387 1259 388 1263
rect 382 1258 388 1259
rect 392 1255 394 1271
rect 448 1264 450 1282
rect 454 1276 460 1277
rect 454 1272 455 1276
rect 459 1272 460 1276
rect 454 1271 460 1272
rect 446 1263 452 1264
rect 446 1259 447 1263
rect 451 1259 452 1263
rect 446 1258 452 1259
rect 456 1255 458 1271
rect 520 1264 522 1282
rect 526 1276 532 1277
rect 526 1272 527 1276
rect 531 1272 532 1276
rect 526 1271 532 1272
rect 518 1263 524 1264
rect 518 1259 519 1263
rect 523 1259 524 1263
rect 518 1258 524 1259
rect 528 1255 530 1271
rect 592 1264 594 1282
rect 598 1276 604 1277
rect 598 1272 599 1276
rect 603 1272 604 1276
rect 598 1271 604 1272
rect 670 1276 676 1277
rect 670 1272 671 1276
rect 675 1272 676 1276
rect 670 1271 676 1272
rect 590 1263 596 1264
rect 590 1259 591 1263
rect 595 1259 596 1263
rect 590 1258 596 1259
rect 566 1255 572 1256
rect 600 1255 602 1271
rect 672 1255 674 1271
rect 736 1264 738 1282
rect 742 1276 748 1277
rect 742 1272 743 1276
rect 747 1272 748 1276
rect 742 1271 748 1272
rect 734 1263 740 1264
rect 734 1259 735 1263
rect 739 1259 740 1263
rect 734 1258 740 1259
rect 744 1255 746 1271
rect 111 1254 115 1255
rect 111 1249 115 1250
rect 263 1254 267 1255
rect 263 1249 267 1250
rect 311 1254 315 1255
rect 311 1249 315 1250
rect 335 1254 339 1255
rect 335 1249 339 1250
rect 359 1254 363 1255
rect 359 1249 363 1250
rect 391 1254 395 1255
rect 391 1249 395 1250
rect 415 1254 419 1255
rect 415 1249 419 1250
rect 455 1254 459 1255
rect 455 1249 459 1250
rect 479 1254 483 1255
rect 479 1249 483 1250
rect 527 1254 531 1255
rect 527 1249 531 1250
rect 543 1254 547 1255
rect 566 1251 567 1255
rect 571 1251 572 1255
rect 566 1250 572 1251
rect 599 1254 603 1255
rect 543 1249 547 1250
rect 112 1229 114 1249
rect 264 1237 266 1249
rect 270 1247 276 1248
rect 270 1243 271 1247
rect 275 1243 276 1247
rect 270 1242 276 1243
rect 290 1247 296 1248
rect 290 1243 291 1247
rect 295 1243 296 1247
rect 290 1242 296 1243
rect 262 1236 268 1237
rect 262 1232 263 1236
rect 267 1232 268 1236
rect 262 1231 268 1232
rect 110 1228 116 1229
rect 110 1224 111 1228
rect 115 1224 116 1228
rect 110 1223 116 1224
rect 110 1211 116 1212
rect 110 1207 111 1211
rect 115 1207 116 1211
rect 110 1206 116 1207
rect 262 1208 268 1209
rect 112 1203 114 1206
rect 262 1204 263 1208
rect 267 1204 268 1208
rect 262 1203 268 1204
rect 111 1202 115 1203
rect 111 1197 115 1198
rect 223 1202 227 1203
rect 223 1197 227 1198
rect 263 1202 267 1203
rect 263 1197 267 1198
rect 112 1194 114 1197
rect 222 1196 228 1197
rect 110 1193 116 1194
rect 110 1189 111 1193
rect 115 1189 116 1193
rect 222 1192 223 1196
rect 227 1192 228 1196
rect 222 1191 228 1192
rect 110 1188 116 1189
rect 272 1188 274 1242
rect 292 1224 294 1242
rect 312 1237 314 1249
rect 360 1237 362 1249
rect 416 1237 418 1249
rect 442 1247 448 1248
rect 442 1243 443 1247
rect 447 1243 448 1247
rect 442 1242 448 1243
rect 310 1236 316 1237
rect 310 1232 311 1236
rect 315 1232 316 1236
rect 310 1231 316 1232
rect 358 1236 364 1237
rect 358 1232 359 1236
rect 363 1232 364 1236
rect 358 1231 364 1232
rect 414 1236 420 1237
rect 414 1232 415 1236
rect 419 1232 420 1236
rect 414 1231 420 1232
rect 444 1224 446 1242
rect 480 1237 482 1249
rect 518 1247 524 1248
rect 518 1243 519 1247
rect 523 1243 524 1247
rect 518 1242 524 1243
rect 478 1236 484 1237
rect 478 1232 479 1236
rect 483 1232 484 1236
rect 478 1231 484 1232
rect 520 1224 522 1242
rect 544 1237 546 1249
rect 542 1236 548 1237
rect 542 1232 543 1236
rect 547 1232 548 1236
rect 542 1231 548 1232
rect 568 1224 570 1250
rect 599 1249 603 1250
rect 607 1254 611 1255
rect 607 1249 611 1250
rect 671 1254 675 1255
rect 671 1249 675 1250
rect 735 1254 739 1255
rect 735 1249 739 1250
rect 743 1254 747 1255
rect 743 1249 747 1250
rect 608 1237 610 1249
rect 672 1237 674 1249
rect 722 1247 728 1248
rect 722 1243 723 1247
rect 727 1243 728 1247
rect 722 1242 728 1243
rect 606 1236 612 1237
rect 606 1232 607 1236
rect 611 1232 612 1236
rect 606 1231 612 1232
rect 670 1236 676 1237
rect 670 1232 671 1236
rect 675 1232 676 1236
rect 670 1231 676 1232
rect 724 1224 726 1242
rect 736 1237 738 1249
rect 792 1248 794 1282
rect 822 1276 828 1277
rect 822 1272 823 1276
rect 827 1272 828 1276
rect 822 1271 828 1272
rect 824 1255 826 1271
rect 844 1264 846 1326
rect 862 1316 868 1317
rect 862 1312 863 1316
rect 867 1312 868 1316
rect 862 1311 868 1312
rect 926 1316 932 1317
rect 926 1312 927 1316
rect 931 1312 932 1316
rect 926 1311 932 1312
rect 863 1310 867 1311
rect 863 1305 867 1306
rect 903 1310 907 1311
rect 903 1305 907 1306
rect 927 1310 931 1311
rect 927 1305 931 1306
rect 902 1304 908 1305
rect 902 1300 903 1304
rect 907 1300 908 1304
rect 902 1299 908 1300
rect 918 1287 924 1288
rect 918 1283 919 1287
rect 923 1283 924 1287
rect 918 1282 924 1283
rect 902 1276 908 1277
rect 902 1272 903 1276
rect 907 1272 908 1276
rect 902 1271 908 1272
rect 842 1263 848 1264
rect 842 1259 843 1263
rect 847 1259 848 1263
rect 842 1258 848 1259
rect 904 1255 906 1271
rect 799 1254 803 1255
rect 799 1249 803 1250
rect 823 1254 827 1255
rect 823 1249 827 1250
rect 863 1254 867 1255
rect 863 1249 867 1250
rect 903 1254 907 1255
rect 903 1249 907 1250
rect 782 1247 788 1248
rect 782 1243 783 1247
rect 787 1243 788 1247
rect 782 1242 788 1243
rect 790 1247 796 1248
rect 790 1243 791 1247
rect 795 1243 796 1247
rect 790 1242 796 1243
rect 734 1236 740 1237
rect 734 1232 735 1236
rect 739 1232 740 1236
rect 734 1231 740 1232
rect 784 1224 786 1242
rect 800 1237 802 1249
rect 864 1237 866 1249
rect 920 1248 922 1282
rect 976 1264 978 1326
rect 998 1316 1004 1317
rect 998 1312 999 1316
rect 1003 1312 1004 1316
rect 998 1311 1004 1312
rect 1046 1316 1052 1317
rect 1046 1312 1047 1316
rect 1051 1312 1052 1316
rect 1046 1311 1052 1312
rect 983 1310 987 1311
rect 983 1305 987 1306
rect 999 1310 1003 1311
rect 999 1305 1003 1306
rect 1047 1310 1051 1311
rect 1047 1305 1051 1306
rect 982 1304 988 1305
rect 982 1300 983 1304
rect 987 1300 988 1304
rect 982 1299 988 1300
rect 1046 1304 1052 1305
rect 1046 1300 1047 1304
rect 1051 1300 1052 1304
rect 1046 1299 1052 1300
rect 1072 1288 1074 1350
rect 1096 1337 1098 1357
rect 1136 1355 1138 1379
rect 1158 1376 1164 1377
rect 1158 1372 1159 1376
rect 1163 1372 1164 1376
rect 1158 1371 1164 1372
rect 1160 1355 1162 1371
rect 1188 1364 1190 1382
rect 1198 1376 1204 1377
rect 1198 1372 1199 1376
rect 1203 1372 1204 1376
rect 1198 1371 1204 1372
rect 1186 1363 1192 1364
rect 1186 1359 1187 1363
rect 1191 1359 1192 1363
rect 1186 1358 1192 1359
rect 1200 1355 1202 1371
rect 1256 1364 1258 1382
rect 1262 1376 1268 1377
rect 1262 1372 1263 1376
rect 1267 1372 1268 1376
rect 1262 1371 1268 1372
rect 1254 1363 1260 1364
rect 1254 1359 1255 1363
rect 1259 1359 1260 1363
rect 1254 1358 1260 1359
rect 1264 1355 1266 1371
rect 1344 1364 1346 1382
rect 1350 1376 1356 1377
rect 1350 1372 1351 1376
rect 1355 1372 1356 1376
rect 1350 1371 1356 1372
rect 1342 1363 1348 1364
rect 1342 1359 1343 1363
rect 1347 1359 1348 1363
rect 1342 1358 1348 1359
rect 1352 1355 1354 1371
rect 1440 1364 1442 1382
rect 1446 1376 1452 1377
rect 1446 1372 1447 1376
rect 1451 1372 1452 1376
rect 1446 1371 1452 1372
rect 1438 1363 1444 1364
rect 1438 1359 1439 1363
rect 1443 1359 1444 1363
rect 1438 1358 1444 1359
rect 1448 1355 1450 1371
rect 1536 1364 1538 1382
rect 1542 1376 1548 1377
rect 1542 1372 1543 1376
rect 1547 1372 1548 1376
rect 1542 1371 1548 1372
rect 1630 1376 1636 1377
rect 1630 1372 1631 1376
rect 1635 1372 1636 1376
rect 1630 1371 1636 1372
rect 1671 1372 1675 1373
rect 1534 1363 1540 1364
rect 1534 1359 1535 1363
rect 1539 1359 1540 1363
rect 1534 1358 1540 1359
rect 1510 1355 1516 1356
rect 1544 1355 1546 1371
rect 1632 1355 1634 1371
rect 1671 1367 1675 1368
rect 1672 1364 1674 1367
rect 1712 1364 1714 1382
rect 1718 1376 1724 1377
rect 1718 1372 1719 1376
rect 1723 1372 1724 1376
rect 1718 1371 1724 1372
rect 1670 1363 1676 1364
rect 1670 1359 1671 1363
rect 1675 1359 1676 1363
rect 1670 1358 1676 1359
rect 1710 1363 1716 1364
rect 1710 1359 1711 1363
rect 1715 1359 1716 1363
rect 1710 1358 1716 1359
rect 1720 1355 1722 1371
rect 1792 1364 1794 1382
rect 1798 1376 1804 1377
rect 1798 1372 1799 1376
rect 1803 1372 1804 1376
rect 1798 1371 1804 1372
rect 1790 1363 1796 1364
rect 1790 1359 1791 1363
rect 1795 1359 1796 1363
rect 1790 1358 1796 1359
rect 1800 1355 1802 1371
rect 1864 1364 1866 1382
rect 1870 1376 1876 1377
rect 1870 1372 1871 1376
rect 1875 1372 1876 1376
rect 1870 1371 1876 1372
rect 1862 1363 1868 1364
rect 1862 1359 1863 1363
rect 1867 1359 1868 1363
rect 1862 1358 1868 1359
rect 1872 1355 1874 1371
rect 1878 1363 1884 1364
rect 1878 1359 1879 1363
rect 1883 1359 1884 1363
rect 1878 1358 1884 1359
rect 1135 1354 1139 1355
rect 1135 1349 1139 1350
rect 1159 1354 1163 1355
rect 1159 1349 1163 1350
rect 1199 1354 1203 1355
rect 1199 1349 1203 1350
rect 1255 1354 1259 1355
rect 1255 1349 1259 1350
rect 1263 1354 1267 1355
rect 1263 1349 1267 1350
rect 1351 1354 1355 1355
rect 1351 1349 1355 1350
rect 1375 1354 1379 1355
rect 1375 1349 1379 1350
rect 1447 1354 1451 1355
rect 1447 1349 1451 1350
rect 1487 1354 1491 1355
rect 1510 1351 1511 1355
rect 1515 1351 1516 1355
rect 1510 1350 1516 1351
rect 1543 1354 1547 1355
rect 1487 1349 1491 1350
rect 1094 1336 1100 1337
rect 1094 1332 1095 1336
rect 1099 1332 1100 1336
rect 1094 1331 1100 1332
rect 1136 1329 1138 1349
rect 1160 1337 1162 1349
rect 1186 1347 1192 1348
rect 1186 1343 1187 1347
rect 1191 1343 1192 1347
rect 1186 1342 1192 1343
rect 1158 1336 1164 1337
rect 1158 1332 1159 1336
rect 1163 1332 1164 1336
rect 1158 1331 1164 1332
rect 1134 1328 1140 1329
rect 1134 1324 1135 1328
rect 1139 1324 1140 1328
rect 1188 1324 1190 1342
rect 1256 1337 1258 1349
rect 1282 1347 1288 1348
rect 1282 1343 1283 1347
rect 1287 1343 1288 1347
rect 1282 1342 1288 1343
rect 1254 1336 1260 1337
rect 1254 1332 1255 1336
rect 1259 1332 1260 1336
rect 1254 1331 1260 1332
rect 1284 1324 1286 1342
rect 1376 1337 1378 1349
rect 1402 1347 1408 1348
rect 1402 1343 1403 1347
rect 1407 1343 1408 1347
rect 1402 1342 1408 1343
rect 1374 1336 1380 1337
rect 1374 1332 1375 1336
rect 1379 1332 1380 1336
rect 1374 1331 1380 1332
rect 1404 1324 1406 1342
rect 1488 1337 1490 1349
rect 1486 1336 1492 1337
rect 1486 1332 1487 1336
rect 1491 1332 1492 1336
rect 1486 1331 1492 1332
rect 1512 1324 1514 1350
rect 1543 1349 1547 1350
rect 1591 1354 1595 1355
rect 1591 1349 1595 1350
rect 1631 1354 1635 1355
rect 1631 1349 1635 1350
rect 1679 1354 1683 1355
rect 1679 1349 1683 1350
rect 1719 1354 1723 1355
rect 1719 1349 1723 1350
rect 1759 1354 1763 1355
rect 1759 1349 1763 1350
rect 1799 1354 1803 1355
rect 1799 1349 1803 1350
rect 1831 1354 1835 1355
rect 1831 1349 1835 1350
rect 1871 1354 1875 1355
rect 1871 1349 1875 1350
rect 1592 1337 1594 1349
rect 1618 1347 1624 1348
rect 1618 1343 1619 1347
rect 1623 1343 1624 1347
rect 1618 1342 1624 1343
rect 1590 1336 1596 1337
rect 1590 1332 1591 1336
rect 1595 1332 1596 1336
rect 1590 1331 1596 1332
rect 1620 1324 1622 1342
rect 1680 1337 1682 1349
rect 1706 1347 1712 1348
rect 1706 1343 1707 1347
rect 1711 1343 1712 1347
rect 1706 1342 1712 1343
rect 1678 1336 1684 1337
rect 1678 1332 1679 1336
rect 1683 1332 1684 1336
rect 1678 1331 1684 1332
rect 1708 1324 1710 1342
rect 1760 1337 1762 1349
rect 1786 1347 1792 1348
rect 1786 1343 1787 1347
rect 1791 1343 1792 1347
rect 1786 1342 1792 1343
rect 1758 1336 1764 1337
rect 1758 1332 1759 1336
rect 1763 1332 1764 1336
rect 1758 1331 1764 1332
rect 1788 1324 1790 1342
rect 1832 1337 1834 1349
rect 1830 1336 1836 1337
rect 1830 1332 1831 1336
rect 1835 1332 1836 1336
rect 1830 1331 1836 1332
rect 1880 1324 1882 1358
rect 1888 1356 1890 1382
rect 1932 1373 1934 1430
rect 1990 1420 1996 1421
rect 1990 1416 1991 1420
rect 1995 1416 1996 1420
rect 1990 1415 1996 1416
rect 1992 1411 1994 1415
rect 1943 1410 1947 1411
rect 1943 1405 1947 1406
rect 1991 1410 1995 1411
rect 1991 1405 1995 1406
rect 2015 1410 2019 1411
rect 2015 1405 2019 1406
rect 1942 1404 1948 1405
rect 1942 1400 1943 1404
rect 1947 1400 1948 1404
rect 1942 1399 1948 1400
rect 2014 1404 2020 1405
rect 2014 1400 2015 1404
rect 2019 1400 2020 1404
rect 2014 1399 2020 1400
rect 2040 1388 2042 1466
rect 2071 1461 2075 1462
rect 2072 1449 2074 1461
rect 2080 1460 2082 1490
rect 2118 1488 2119 1492
rect 2123 1488 2124 1492
rect 2118 1487 2124 1488
rect 2120 1467 2122 1487
rect 2119 1466 2123 1467
rect 2119 1461 2123 1462
rect 2078 1459 2084 1460
rect 2078 1455 2079 1459
rect 2083 1455 2084 1459
rect 2078 1454 2084 1455
rect 2070 1448 2076 1449
rect 2070 1444 2071 1448
rect 2075 1444 2076 1448
rect 2070 1443 2076 1444
rect 2120 1441 2122 1461
rect 2118 1440 2124 1441
rect 2118 1436 2119 1440
rect 2123 1436 2124 1440
rect 2090 1435 2096 1436
rect 2118 1435 2124 1436
rect 2090 1431 2091 1435
rect 2095 1431 2096 1435
rect 2090 1430 2096 1431
rect 2070 1420 2076 1421
rect 2070 1416 2071 1420
rect 2075 1416 2076 1420
rect 2070 1415 2076 1416
rect 2072 1411 2074 1415
rect 2071 1410 2075 1411
rect 2071 1405 2075 1406
rect 2070 1404 2076 1405
rect 2070 1400 2071 1404
rect 2075 1400 2076 1404
rect 2070 1399 2076 1400
rect 2006 1387 2012 1388
rect 2006 1383 2007 1387
rect 2011 1383 2012 1387
rect 2006 1382 2012 1383
rect 2038 1387 2044 1388
rect 2038 1383 2039 1387
rect 2043 1383 2044 1387
rect 2038 1382 2044 1383
rect 2082 1387 2088 1388
rect 2082 1383 2083 1387
rect 2087 1383 2088 1387
rect 2082 1382 2088 1383
rect 1942 1376 1948 1377
rect 1931 1372 1935 1373
rect 1942 1372 1943 1376
rect 1947 1372 1948 1376
rect 1942 1371 1948 1372
rect 1931 1367 1935 1368
rect 1886 1355 1892 1356
rect 1944 1355 1946 1371
rect 2008 1364 2010 1382
rect 2014 1376 2020 1377
rect 2014 1372 2015 1376
rect 2019 1372 2020 1376
rect 2014 1371 2020 1372
rect 2070 1376 2076 1377
rect 2070 1372 2071 1376
rect 2075 1372 2076 1376
rect 2070 1371 2076 1372
rect 2006 1363 2012 1364
rect 2006 1359 2007 1363
rect 2011 1359 2012 1363
rect 2006 1358 2012 1359
rect 1990 1355 1996 1356
rect 2016 1355 2018 1371
rect 2072 1355 2074 1371
rect 1886 1351 1887 1355
rect 1891 1351 1892 1355
rect 1886 1350 1892 1351
rect 1903 1354 1907 1355
rect 1903 1349 1907 1350
rect 1943 1354 1947 1355
rect 1943 1349 1947 1350
rect 1967 1354 1971 1355
rect 1990 1351 1991 1355
rect 1995 1351 1996 1355
rect 1990 1350 1996 1351
rect 2015 1354 2019 1355
rect 1967 1349 1971 1350
rect 1904 1337 1906 1349
rect 1968 1337 1970 1349
rect 1902 1336 1908 1337
rect 1902 1332 1903 1336
rect 1907 1332 1908 1336
rect 1902 1331 1908 1332
rect 1966 1336 1972 1337
rect 1966 1332 1967 1336
rect 1971 1332 1972 1336
rect 1966 1331 1972 1332
rect 1992 1324 1994 1350
rect 2015 1349 2019 1350
rect 2031 1354 2035 1355
rect 2031 1349 2035 1350
rect 2071 1354 2075 1355
rect 2071 1349 2075 1350
rect 2032 1337 2034 1349
rect 2046 1347 2052 1348
rect 2046 1343 2047 1347
rect 2051 1343 2052 1347
rect 2046 1342 2052 1343
rect 2030 1336 2036 1337
rect 2030 1332 2031 1336
rect 2035 1332 2036 1336
rect 2030 1331 2036 1332
rect 1134 1323 1140 1324
rect 1186 1323 1192 1324
rect 1094 1319 1100 1320
rect 1094 1315 1095 1319
rect 1099 1315 1100 1319
rect 1186 1319 1187 1323
rect 1191 1319 1192 1323
rect 1186 1318 1192 1319
rect 1282 1323 1288 1324
rect 1282 1319 1283 1323
rect 1287 1319 1288 1323
rect 1282 1318 1288 1319
rect 1402 1323 1408 1324
rect 1402 1319 1403 1323
rect 1407 1319 1408 1323
rect 1402 1318 1408 1319
rect 1510 1323 1516 1324
rect 1510 1319 1511 1323
rect 1515 1319 1516 1323
rect 1510 1318 1516 1319
rect 1618 1323 1624 1324
rect 1618 1319 1619 1323
rect 1623 1319 1624 1323
rect 1618 1318 1624 1319
rect 1706 1323 1712 1324
rect 1706 1319 1707 1323
rect 1711 1319 1712 1323
rect 1706 1318 1712 1319
rect 1786 1323 1792 1324
rect 1786 1319 1787 1323
rect 1791 1319 1792 1323
rect 1786 1318 1792 1319
rect 1878 1323 1884 1324
rect 1878 1319 1879 1323
rect 1883 1319 1884 1323
rect 1878 1318 1884 1319
rect 1958 1323 1964 1324
rect 1958 1319 1959 1323
rect 1963 1319 1964 1323
rect 1958 1318 1964 1319
rect 1990 1323 1996 1324
rect 1990 1319 1991 1323
rect 1995 1319 1996 1323
rect 1990 1318 1996 1319
rect 1094 1314 1100 1315
rect 1096 1311 1098 1314
rect 1134 1311 1140 1312
rect 1095 1310 1099 1311
rect 1134 1307 1135 1311
rect 1139 1307 1140 1311
rect 1134 1306 1140 1307
rect 1158 1308 1164 1309
rect 1095 1305 1099 1306
rect 1096 1302 1098 1305
rect 1094 1301 1100 1302
rect 1094 1297 1095 1301
rect 1099 1297 1100 1301
rect 1136 1299 1138 1306
rect 1158 1304 1159 1308
rect 1163 1304 1164 1308
rect 1158 1303 1164 1304
rect 1254 1308 1260 1309
rect 1254 1304 1255 1308
rect 1259 1304 1260 1308
rect 1254 1303 1260 1304
rect 1374 1308 1380 1309
rect 1374 1304 1375 1308
rect 1379 1304 1380 1308
rect 1374 1303 1380 1304
rect 1486 1308 1492 1309
rect 1486 1304 1487 1308
rect 1491 1304 1492 1308
rect 1486 1303 1492 1304
rect 1590 1308 1596 1309
rect 1590 1304 1591 1308
rect 1595 1304 1596 1308
rect 1590 1303 1596 1304
rect 1678 1308 1684 1309
rect 1678 1304 1679 1308
rect 1683 1304 1684 1308
rect 1678 1303 1684 1304
rect 1758 1308 1764 1309
rect 1758 1304 1759 1308
rect 1763 1304 1764 1308
rect 1758 1303 1764 1304
rect 1830 1308 1836 1309
rect 1830 1304 1831 1308
rect 1835 1304 1836 1308
rect 1830 1303 1836 1304
rect 1902 1308 1908 1309
rect 1902 1304 1903 1308
rect 1907 1304 1908 1308
rect 1902 1303 1908 1304
rect 1160 1299 1162 1303
rect 1256 1299 1258 1303
rect 1376 1299 1378 1303
rect 1488 1299 1490 1303
rect 1592 1299 1594 1303
rect 1680 1299 1682 1303
rect 1760 1299 1762 1303
rect 1832 1299 1834 1303
rect 1904 1299 1906 1303
rect 1094 1296 1100 1297
rect 1135 1298 1139 1299
rect 1135 1293 1139 1294
rect 1159 1298 1163 1299
rect 1159 1293 1163 1294
rect 1199 1298 1203 1299
rect 1199 1293 1203 1294
rect 1247 1298 1251 1299
rect 1247 1293 1251 1294
rect 1255 1298 1259 1299
rect 1255 1293 1259 1294
rect 1319 1298 1323 1299
rect 1319 1293 1323 1294
rect 1375 1298 1379 1299
rect 1375 1293 1379 1294
rect 1399 1298 1403 1299
rect 1399 1293 1403 1294
rect 1479 1298 1483 1299
rect 1479 1293 1483 1294
rect 1487 1298 1491 1299
rect 1487 1293 1491 1294
rect 1559 1298 1563 1299
rect 1559 1293 1563 1294
rect 1591 1298 1595 1299
rect 1591 1293 1595 1294
rect 1639 1298 1643 1299
rect 1639 1293 1643 1294
rect 1679 1298 1683 1299
rect 1679 1293 1683 1294
rect 1719 1298 1723 1299
rect 1719 1293 1723 1294
rect 1759 1298 1763 1299
rect 1759 1293 1763 1294
rect 1799 1298 1803 1299
rect 1799 1293 1803 1294
rect 1831 1298 1835 1299
rect 1831 1293 1835 1294
rect 1879 1298 1883 1299
rect 1879 1293 1883 1294
rect 1903 1298 1907 1299
rect 1903 1293 1907 1294
rect 1136 1290 1138 1293
rect 1158 1292 1164 1293
rect 1134 1289 1140 1290
rect 1070 1287 1076 1288
rect 1070 1283 1071 1287
rect 1075 1283 1076 1287
rect 1134 1285 1135 1289
rect 1139 1285 1140 1289
rect 1158 1288 1159 1292
rect 1163 1288 1164 1292
rect 1158 1287 1164 1288
rect 1198 1292 1204 1293
rect 1198 1288 1199 1292
rect 1203 1288 1204 1292
rect 1198 1287 1204 1288
rect 1246 1292 1252 1293
rect 1246 1288 1247 1292
rect 1251 1288 1252 1292
rect 1246 1287 1252 1288
rect 1318 1292 1324 1293
rect 1318 1288 1319 1292
rect 1323 1288 1324 1292
rect 1318 1287 1324 1288
rect 1398 1292 1404 1293
rect 1398 1288 1399 1292
rect 1403 1288 1404 1292
rect 1398 1287 1404 1288
rect 1478 1292 1484 1293
rect 1478 1288 1479 1292
rect 1483 1288 1484 1292
rect 1478 1287 1484 1288
rect 1558 1292 1564 1293
rect 1558 1288 1559 1292
rect 1563 1288 1564 1292
rect 1558 1287 1564 1288
rect 1638 1292 1644 1293
rect 1638 1288 1639 1292
rect 1643 1288 1644 1292
rect 1638 1287 1644 1288
rect 1718 1292 1724 1293
rect 1718 1288 1719 1292
rect 1723 1288 1724 1292
rect 1718 1287 1724 1288
rect 1798 1292 1804 1293
rect 1798 1288 1799 1292
rect 1803 1288 1804 1292
rect 1798 1287 1804 1288
rect 1878 1292 1884 1293
rect 1878 1288 1879 1292
rect 1883 1288 1884 1292
rect 1878 1287 1884 1288
rect 1070 1282 1076 1283
rect 1094 1284 1100 1285
rect 1134 1284 1140 1285
rect 1094 1280 1095 1284
rect 1099 1280 1100 1284
rect 1094 1279 1100 1280
rect 1270 1283 1276 1284
rect 1270 1279 1271 1283
rect 1275 1279 1276 1283
rect 982 1276 988 1277
rect 982 1272 983 1276
rect 987 1272 988 1276
rect 982 1271 988 1272
rect 1046 1276 1052 1277
rect 1046 1272 1047 1276
rect 1051 1272 1052 1276
rect 1046 1271 1052 1272
rect 974 1263 980 1264
rect 974 1259 975 1263
rect 979 1259 980 1263
rect 974 1258 980 1259
rect 984 1255 986 1271
rect 1048 1255 1050 1271
rect 1096 1255 1098 1279
rect 1270 1278 1276 1279
rect 1134 1272 1140 1273
rect 1134 1268 1135 1272
rect 1139 1268 1140 1272
rect 1134 1267 1140 1268
rect 927 1254 931 1255
rect 927 1249 931 1250
rect 983 1254 987 1255
rect 983 1249 987 1250
rect 1047 1254 1051 1255
rect 1047 1249 1051 1250
rect 1095 1254 1099 1255
rect 1095 1249 1099 1250
rect 910 1247 916 1248
rect 910 1243 911 1247
rect 915 1243 916 1247
rect 910 1242 916 1243
rect 918 1247 924 1248
rect 918 1243 919 1247
rect 923 1243 924 1247
rect 918 1242 924 1243
rect 798 1236 804 1237
rect 798 1232 799 1236
rect 803 1232 804 1236
rect 798 1231 804 1232
rect 862 1236 868 1237
rect 862 1232 863 1236
rect 867 1232 868 1236
rect 862 1231 868 1232
rect 912 1224 914 1242
rect 928 1237 930 1249
rect 926 1236 932 1237
rect 926 1232 927 1236
rect 931 1232 932 1236
rect 926 1231 932 1232
rect 1096 1229 1098 1249
rect 1136 1243 1138 1267
rect 1158 1264 1164 1265
rect 1158 1260 1159 1264
rect 1163 1260 1164 1264
rect 1158 1259 1164 1260
rect 1198 1264 1204 1265
rect 1198 1260 1199 1264
rect 1203 1260 1204 1264
rect 1198 1259 1204 1260
rect 1246 1264 1252 1265
rect 1246 1260 1247 1264
rect 1251 1260 1252 1264
rect 1272 1260 1274 1278
rect 1390 1275 1396 1276
rect 1390 1271 1391 1275
rect 1395 1271 1396 1275
rect 1390 1270 1396 1271
rect 1470 1275 1476 1276
rect 1470 1271 1471 1275
rect 1475 1271 1476 1275
rect 1470 1270 1476 1271
rect 1630 1275 1636 1276
rect 1630 1271 1631 1275
rect 1635 1271 1636 1275
rect 1630 1270 1636 1271
rect 1710 1275 1716 1276
rect 1710 1271 1711 1275
rect 1715 1271 1716 1275
rect 1710 1270 1716 1271
rect 1814 1275 1820 1276
rect 1814 1271 1815 1275
rect 1819 1271 1820 1275
rect 1814 1270 1820 1271
rect 1822 1275 1828 1276
rect 1822 1271 1823 1275
rect 1827 1271 1828 1275
rect 1822 1270 1828 1271
rect 1834 1275 1840 1276
rect 1834 1271 1835 1275
rect 1839 1271 1840 1275
rect 1834 1270 1840 1271
rect 1318 1264 1324 1265
rect 1318 1260 1319 1264
rect 1323 1260 1324 1264
rect 1246 1259 1252 1260
rect 1270 1259 1276 1260
rect 1318 1259 1324 1260
rect 1160 1243 1162 1259
rect 1200 1243 1202 1259
rect 1248 1243 1250 1259
rect 1270 1255 1271 1259
rect 1275 1255 1276 1259
rect 1270 1254 1276 1255
rect 1266 1251 1272 1252
rect 1266 1247 1267 1251
rect 1271 1247 1272 1251
rect 1266 1246 1272 1247
rect 1135 1242 1139 1243
rect 1135 1237 1139 1238
rect 1159 1242 1163 1243
rect 1159 1237 1163 1238
rect 1199 1242 1203 1243
rect 1199 1237 1203 1238
rect 1239 1242 1243 1243
rect 1239 1237 1243 1238
rect 1247 1242 1251 1243
rect 1247 1237 1251 1238
rect 1094 1228 1100 1229
rect 1094 1224 1095 1228
rect 1099 1224 1100 1228
rect 290 1223 296 1224
rect 290 1219 291 1223
rect 295 1219 296 1223
rect 290 1218 296 1219
rect 442 1223 448 1224
rect 442 1219 443 1223
rect 447 1219 448 1223
rect 442 1218 448 1219
rect 518 1223 524 1224
rect 518 1219 519 1223
rect 523 1219 524 1223
rect 518 1218 524 1219
rect 566 1223 572 1224
rect 566 1219 567 1223
rect 571 1219 572 1223
rect 566 1218 572 1219
rect 578 1223 584 1224
rect 578 1219 579 1223
rect 583 1219 584 1223
rect 578 1218 584 1219
rect 722 1223 728 1224
rect 722 1219 723 1223
rect 727 1219 728 1223
rect 722 1218 728 1219
rect 782 1223 788 1224
rect 782 1219 783 1223
rect 787 1219 788 1223
rect 782 1218 788 1219
rect 886 1223 892 1224
rect 886 1219 887 1223
rect 891 1219 892 1223
rect 886 1218 892 1219
rect 910 1223 916 1224
rect 1094 1223 1100 1224
rect 910 1219 911 1223
rect 915 1219 916 1223
rect 910 1218 916 1219
rect 310 1208 316 1209
rect 310 1204 311 1208
rect 315 1204 316 1208
rect 310 1203 316 1204
rect 358 1208 364 1209
rect 358 1204 359 1208
rect 363 1204 364 1208
rect 358 1203 364 1204
rect 414 1208 420 1209
rect 414 1204 415 1208
rect 419 1204 420 1208
rect 414 1203 420 1204
rect 478 1208 484 1209
rect 478 1204 479 1208
rect 483 1204 484 1208
rect 478 1203 484 1204
rect 542 1208 548 1209
rect 542 1204 543 1208
rect 547 1204 548 1208
rect 542 1203 548 1204
rect 279 1202 283 1203
rect 279 1197 283 1198
rect 311 1202 315 1203
rect 311 1197 315 1198
rect 343 1202 347 1203
rect 343 1197 347 1198
rect 359 1202 363 1203
rect 359 1197 363 1198
rect 407 1202 411 1203
rect 407 1197 411 1198
rect 415 1202 419 1203
rect 415 1197 419 1198
rect 479 1202 483 1203
rect 479 1197 483 1198
rect 543 1202 547 1203
rect 543 1197 547 1198
rect 551 1202 555 1203
rect 551 1197 555 1198
rect 278 1196 284 1197
rect 278 1192 279 1196
rect 283 1192 284 1196
rect 278 1191 284 1192
rect 342 1196 348 1197
rect 342 1192 343 1196
rect 347 1192 348 1196
rect 342 1191 348 1192
rect 406 1196 412 1197
rect 406 1192 407 1196
rect 411 1192 412 1196
rect 406 1191 412 1192
rect 478 1196 484 1197
rect 478 1192 479 1196
rect 483 1192 484 1196
rect 478 1191 484 1192
rect 550 1196 556 1197
rect 550 1192 551 1196
rect 555 1192 556 1196
rect 550 1191 556 1192
rect 270 1187 276 1188
rect 270 1183 271 1187
rect 275 1183 276 1187
rect 270 1182 276 1183
rect 270 1179 276 1180
rect 110 1176 116 1177
rect 110 1172 111 1176
rect 115 1172 116 1176
rect 270 1175 271 1179
rect 275 1175 276 1179
rect 270 1174 276 1175
rect 334 1179 340 1180
rect 334 1175 335 1179
rect 339 1175 340 1179
rect 334 1174 340 1175
rect 398 1179 404 1180
rect 398 1175 399 1179
rect 403 1175 404 1179
rect 398 1174 404 1175
rect 470 1179 476 1180
rect 470 1175 471 1179
rect 475 1175 476 1179
rect 470 1174 476 1175
rect 110 1171 116 1172
rect 112 1151 114 1171
rect 222 1168 228 1169
rect 222 1164 223 1168
rect 227 1164 228 1168
rect 222 1163 228 1164
rect 224 1151 226 1163
rect 272 1156 274 1174
rect 278 1168 284 1169
rect 278 1164 279 1168
rect 283 1164 284 1168
rect 278 1163 284 1164
rect 262 1155 268 1156
rect 262 1151 263 1155
rect 267 1151 268 1155
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 159 1150 163 1151
rect 159 1145 163 1146
rect 199 1150 203 1151
rect 199 1145 203 1146
rect 223 1150 227 1151
rect 223 1145 227 1146
rect 247 1150 251 1151
rect 262 1150 268 1151
rect 270 1155 276 1156
rect 270 1151 271 1155
rect 275 1151 276 1155
rect 280 1151 282 1163
rect 336 1156 338 1174
rect 342 1168 348 1169
rect 342 1164 343 1168
rect 347 1164 348 1168
rect 342 1163 348 1164
rect 334 1155 340 1156
rect 334 1151 335 1155
rect 339 1151 340 1155
rect 344 1151 346 1163
rect 400 1156 402 1174
rect 406 1168 412 1169
rect 406 1164 407 1168
rect 411 1164 412 1168
rect 406 1163 412 1164
rect 398 1155 404 1156
rect 398 1151 399 1155
rect 403 1151 404 1155
rect 408 1151 410 1163
rect 472 1156 474 1174
rect 478 1168 484 1169
rect 478 1164 479 1168
rect 483 1164 484 1168
rect 478 1163 484 1164
rect 550 1168 556 1169
rect 550 1164 551 1168
rect 555 1164 556 1168
rect 550 1163 556 1164
rect 470 1155 476 1156
rect 470 1151 471 1155
rect 475 1151 476 1155
rect 480 1151 482 1163
rect 552 1151 554 1163
rect 580 1156 582 1218
rect 606 1208 612 1209
rect 606 1204 607 1208
rect 611 1204 612 1208
rect 606 1203 612 1204
rect 670 1208 676 1209
rect 670 1204 671 1208
rect 675 1204 676 1208
rect 670 1203 676 1204
rect 734 1208 740 1209
rect 734 1204 735 1208
rect 739 1204 740 1208
rect 734 1203 740 1204
rect 798 1208 804 1209
rect 798 1204 799 1208
rect 803 1204 804 1208
rect 798 1203 804 1204
rect 862 1208 868 1209
rect 862 1204 863 1208
rect 867 1204 868 1208
rect 862 1203 868 1204
rect 607 1202 611 1203
rect 607 1197 611 1198
rect 631 1202 635 1203
rect 631 1197 635 1198
rect 671 1202 675 1203
rect 671 1197 675 1198
rect 711 1202 715 1203
rect 711 1197 715 1198
rect 735 1202 739 1203
rect 735 1197 739 1198
rect 791 1202 795 1203
rect 791 1197 795 1198
rect 799 1202 803 1203
rect 799 1197 803 1198
rect 863 1202 867 1203
rect 863 1197 867 1198
rect 871 1202 875 1203
rect 871 1197 875 1198
rect 630 1196 636 1197
rect 630 1192 631 1196
rect 635 1192 636 1196
rect 630 1191 636 1192
rect 710 1196 716 1197
rect 710 1192 711 1196
rect 715 1192 716 1196
rect 710 1191 716 1192
rect 790 1196 796 1197
rect 790 1192 791 1196
rect 795 1192 796 1196
rect 790 1191 796 1192
rect 870 1196 876 1197
rect 870 1192 871 1196
rect 875 1192 876 1196
rect 870 1191 876 1192
rect 622 1179 628 1180
rect 622 1175 623 1179
rect 627 1175 628 1179
rect 622 1174 628 1175
rect 702 1179 708 1180
rect 702 1175 703 1179
rect 707 1175 708 1179
rect 702 1174 708 1175
rect 782 1179 788 1180
rect 782 1175 783 1179
rect 787 1175 788 1179
rect 782 1174 788 1175
rect 798 1179 804 1180
rect 798 1175 799 1179
rect 803 1175 804 1179
rect 798 1174 804 1175
rect 624 1156 626 1174
rect 630 1168 636 1169
rect 630 1164 631 1168
rect 635 1164 636 1168
rect 630 1163 636 1164
rect 578 1155 584 1156
rect 578 1151 579 1155
rect 583 1151 584 1155
rect 622 1155 628 1156
rect 622 1151 623 1155
rect 627 1151 628 1155
rect 632 1151 634 1163
rect 704 1156 706 1174
rect 710 1168 716 1169
rect 710 1164 711 1168
rect 715 1164 716 1168
rect 710 1163 716 1164
rect 702 1155 708 1156
rect 702 1151 703 1155
rect 707 1151 708 1155
rect 712 1151 714 1163
rect 784 1156 786 1174
rect 790 1168 796 1169
rect 790 1164 791 1168
rect 795 1164 796 1168
rect 790 1163 796 1164
rect 782 1155 788 1156
rect 782 1151 783 1155
rect 787 1151 788 1155
rect 792 1151 794 1163
rect 270 1150 276 1151
rect 279 1150 283 1151
rect 247 1145 251 1146
rect 112 1125 114 1145
rect 160 1133 162 1145
rect 174 1143 180 1144
rect 174 1139 175 1143
rect 179 1139 180 1143
rect 174 1138 180 1139
rect 182 1143 188 1144
rect 182 1139 183 1143
rect 187 1139 188 1143
rect 182 1138 188 1139
rect 158 1132 164 1133
rect 158 1128 159 1132
rect 163 1128 164 1132
rect 158 1127 164 1128
rect 110 1124 116 1125
rect 110 1120 111 1124
rect 115 1120 116 1124
rect 110 1119 116 1120
rect 110 1107 116 1108
rect 110 1103 111 1107
rect 115 1103 116 1107
rect 110 1102 116 1103
rect 158 1104 164 1105
rect 112 1091 114 1102
rect 158 1100 159 1104
rect 163 1100 164 1104
rect 158 1099 164 1100
rect 160 1091 162 1099
rect 111 1090 115 1091
rect 111 1085 115 1086
rect 159 1090 163 1091
rect 159 1085 163 1086
rect 112 1082 114 1085
rect 110 1081 116 1082
rect 110 1077 111 1081
rect 115 1077 116 1081
rect 110 1076 116 1077
rect 176 1068 178 1138
rect 184 1120 186 1138
rect 200 1133 202 1145
rect 230 1143 236 1144
rect 230 1139 231 1143
rect 235 1139 236 1143
rect 230 1138 236 1139
rect 198 1132 204 1133
rect 198 1128 199 1132
rect 203 1128 204 1132
rect 198 1127 204 1128
rect 232 1120 234 1138
rect 248 1133 250 1145
rect 246 1132 252 1133
rect 246 1128 247 1132
rect 251 1128 252 1132
rect 264 1128 266 1150
rect 279 1145 283 1146
rect 303 1150 307 1151
rect 334 1150 340 1151
rect 343 1150 347 1151
rect 303 1145 307 1146
rect 343 1145 347 1146
rect 367 1150 371 1151
rect 398 1150 404 1151
rect 407 1150 411 1151
rect 367 1145 371 1146
rect 407 1145 411 1146
rect 439 1150 443 1151
rect 470 1150 476 1151
rect 479 1150 483 1151
rect 439 1145 443 1146
rect 479 1145 483 1146
rect 511 1150 515 1151
rect 511 1145 515 1146
rect 551 1150 555 1151
rect 578 1150 584 1151
rect 591 1150 595 1151
rect 622 1150 628 1151
rect 631 1150 635 1151
rect 551 1145 555 1146
rect 591 1145 595 1146
rect 631 1145 635 1146
rect 679 1150 683 1151
rect 702 1150 708 1151
rect 711 1150 715 1151
rect 679 1145 683 1146
rect 711 1145 715 1146
rect 775 1150 779 1151
rect 782 1150 788 1151
rect 791 1150 795 1151
rect 775 1145 779 1146
rect 791 1145 795 1146
rect 286 1143 292 1144
rect 286 1139 287 1143
rect 291 1139 292 1143
rect 286 1138 292 1139
rect 246 1127 252 1128
rect 262 1127 268 1128
rect 262 1123 263 1127
rect 267 1123 268 1127
rect 262 1122 268 1123
rect 288 1120 290 1138
rect 304 1133 306 1145
rect 368 1133 370 1145
rect 394 1143 400 1144
rect 394 1139 395 1143
rect 399 1139 400 1143
rect 394 1138 400 1139
rect 302 1132 308 1133
rect 302 1128 303 1132
rect 307 1128 308 1132
rect 302 1127 308 1128
rect 366 1132 372 1133
rect 366 1128 367 1132
rect 371 1128 372 1132
rect 366 1127 372 1128
rect 396 1120 398 1138
rect 440 1133 442 1145
rect 512 1133 514 1145
rect 578 1143 584 1144
rect 578 1139 579 1143
rect 583 1139 584 1143
rect 578 1138 584 1139
rect 438 1132 444 1133
rect 438 1128 439 1132
rect 443 1128 444 1132
rect 438 1127 444 1128
rect 510 1132 516 1133
rect 510 1128 511 1132
rect 515 1128 516 1132
rect 510 1127 516 1128
rect 580 1120 582 1138
rect 592 1133 594 1145
rect 666 1143 672 1144
rect 666 1139 667 1143
rect 671 1139 672 1143
rect 666 1138 672 1139
rect 590 1132 596 1133
rect 590 1128 591 1132
rect 595 1128 596 1132
rect 590 1127 596 1128
rect 668 1120 670 1138
rect 680 1133 682 1145
rect 762 1143 768 1144
rect 762 1139 763 1143
rect 767 1139 768 1143
rect 762 1138 768 1139
rect 678 1132 684 1133
rect 678 1128 679 1132
rect 683 1128 684 1132
rect 678 1127 684 1128
rect 764 1120 766 1138
rect 776 1133 778 1145
rect 800 1144 802 1174
rect 870 1168 876 1169
rect 870 1164 871 1168
rect 875 1164 876 1168
rect 870 1163 876 1164
rect 872 1151 874 1163
rect 888 1156 890 1218
rect 1136 1217 1138 1237
rect 1160 1225 1162 1237
rect 1186 1235 1192 1236
rect 1186 1231 1187 1235
rect 1191 1231 1192 1235
rect 1186 1230 1192 1231
rect 1158 1224 1164 1225
rect 1158 1220 1159 1224
rect 1163 1220 1164 1224
rect 1158 1219 1164 1220
rect 1134 1216 1140 1217
rect 1134 1212 1135 1216
rect 1139 1212 1140 1216
rect 1188 1212 1190 1230
rect 1200 1225 1202 1237
rect 1226 1235 1232 1236
rect 1226 1231 1227 1235
rect 1231 1231 1232 1235
rect 1226 1230 1232 1231
rect 1198 1224 1204 1225
rect 1198 1220 1199 1224
rect 1203 1220 1204 1224
rect 1198 1219 1204 1220
rect 1228 1212 1230 1230
rect 1240 1225 1242 1237
rect 1238 1224 1244 1225
rect 1238 1220 1239 1224
rect 1243 1220 1244 1224
rect 1238 1219 1244 1220
rect 1268 1212 1270 1246
rect 1302 1243 1308 1244
rect 1320 1243 1322 1259
rect 1392 1252 1394 1270
rect 1398 1264 1404 1265
rect 1398 1260 1399 1264
rect 1403 1260 1404 1264
rect 1398 1259 1404 1260
rect 1390 1251 1396 1252
rect 1390 1247 1391 1251
rect 1395 1247 1396 1251
rect 1390 1246 1396 1247
rect 1400 1243 1402 1259
rect 1472 1252 1474 1270
rect 1478 1264 1484 1265
rect 1478 1260 1479 1264
rect 1483 1260 1484 1264
rect 1478 1259 1484 1260
rect 1558 1264 1564 1265
rect 1558 1260 1559 1264
rect 1563 1260 1564 1264
rect 1558 1259 1564 1260
rect 1470 1251 1476 1252
rect 1470 1247 1471 1251
rect 1475 1247 1476 1251
rect 1470 1246 1476 1247
rect 1446 1243 1452 1244
rect 1480 1243 1482 1259
rect 1546 1243 1552 1244
rect 1560 1243 1562 1259
rect 1632 1252 1634 1270
rect 1638 1264 1644 1265
rect 1638 1260 1639 1264
rect 1643 1260 1644 1264
rect 1638 1259 1644 1260
rect 1630 1251 1636 1252
rect 1630 1247 1631 1251
rect 1635 1247 1636 1251
rect 1630 1246 1636 1247
rect 1640 1243 1642 1259
rect 1712 1252 1714 1270
rect 1718 1264 1724 1265
rect 1718 1260 1719 1264
rect 1723 1260 1724 1264
rect 1718 1259 1724 1260
rect 1798 1264 1804 1265
rect 1798 1260 1799 1264
rect 1803 1260 1804 1264
rect 1798 1259 1804 1260
rect 1710 1251 1716 1252
rect 1710 1247 1711 1251
rect 1715 1247 1716 1251
rect 1710 1246 1716 1247
rect 1720 1243 1722 1259
rect 1800 1243 1802 1259
rect 1279 1242 1283 1243
rect 1302 1239 1303 1243
rect 1307 1239 1308 1243
rect 1302 1238 1308 1239
rect 1319 1242 1323 1243
rect 1279 1237 1283 1238
rect 1280 1225 1282 1237
rect 1278 1224 1284 1225
rect 1278 1220 1279 1224
rect 1283 1220 1284 1224
rect 1278 1219 1284 1220
rect 1304 1212 1306 1238
rect 1319 1237 1323 1238
rect 1327 1242 1331 1243
rect 1327 1237 1331 1238
rect 1375 1242 1379 1243
rect 1375 1237 1379 1238
rect 1399 1242 1403 1243
rect 1399 1237 1403 1238
rect 1423 1242 1427 1243
rect 1446 1239 1447 1243
rect 1451 1239 1452 1243
rect 1446 1238 1452 1239
rect 1471 1242 1475 1243
rect 1423 1237 1427 1238
rect 1328 1225 1330 1237
rect 1376 1225 1378 1237
rect 1390 1235 1396 1236
rect 1390 1231 1391 1235
rect 1395 1231 1396 1235
rect 1390 1230 1396 1231
rect 1326 1224 1332 1225
rect 1326 1220 1327 1224
rect 1331 1220 1332 1224
rect 1326 1219 1332 1220
rect 1374 1224 1380 1225
rect 1374 1220 1375 1224
rect 1379 1220 1380 1224
rect 1374 1219 1380 1220
rect 1094 1211 1100 1212
rect 1134 1211 1140 1212
rect 1186 1211 1192 1212
rect 926 1208 932 1209
rect 926 1204 927 1208
rect 931 1204 932 1208
rect 1094 1207 1095 1211
rect 1099 1207 1100 1211
rect 1094 1206 1100 1207
rect 1186 1207 1187 1211
rect 1191 1207 1192 1211
rect 1186 1206 1192 1207
rect 1226 1211 1232 1212
rect 1226 1207 1227 1211
rect 1231 1207 1232 1211
rect 1226 1206 1232 1207
rect 1266 1211 1272 1212
rect 1266 1207 1267 1211
rect 1271 1207 1272 1211
rect 1266 1206 1272 1207
rect 1302 1211 1308 1212
rect 1302 1207 1303 1211
rect 1307 1207 1308 1211
rect 1302 1206 1308 1207
rect 926 1203 932 1204
rect 1096 1203 1098 1206
rect 927 1202 931 1203
rect 927 1197 931 1198
rect 959 1202 963 1203
rect 959 1197 963 1198
rect 1095 1202 1099 1203
rect 1095 1197 1099 1198
rect 1134 1199 1140 1200
rect 958 1196 964 1197
rect 958 1192 959 1196
rect 963 1192 964 1196
rect 1096 1194 1098 1197
rect 1134 1195 1135 1199
rect 1139 1195 1140 1199
rect 1134 1194 1140 1195
rect 1158 1196 1164 1197
rect 958 1191 964 1192
rect 1094 1193 1100 1194
rect 1094 1189 1095 1193
rect 1099 1189 1100 1193
rect 1136 1191 1138 1194
rect 1158 1192 1159 1196
rect 1163 1192 1164 1196
rect 1158 1191 1164 1192
rect 1198 1196 1204 1197
rect 1198 1192 1199 1196
rect 1203 1192 1204 1196
rect 1198 1191 1204 1192
rect 1238 1196 1244 1197
rect 1238 1192 1239 1196
rect 1243 1192 1244 1196
rect 1238 1191 1244 1192
rect 1278 1196 1284 1197
rect 1278 1192 1279 1196
rect 1283 1192 1284 1196
rect 1278 1191 1284 1192
rect 1326 1196 1332 1197
rect 1326 1192 1327 1196
rect 1331 1192 1332 1196
rect 1326 1191 1332 1192
rect 1374 1196 1380 1197
rect 1374 1192 1375 1196
rect 1379 1192 1380 1196
rect 1374 1191 1380 1192
rect 1094 1188 1100 1189
rect 1135 1190 1139 1191
rect 1135 1185 1139 1186
rect 1159 1190 1163 1191
rect 1159 1185 1163 1186
rect 1199 1190 1203 1191
rect 1199 1185 1203 1186
rect 1239 1190 1243 1191
rect 1239 1185 1243 1186
rect 1279 1190 1283 1191
rect 1279 1185 1283 1186
rect 1287 1190 1291 1191
rect 1287 1185 1291 1186
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1375 1190 1379 1191
rect 1375 1185 1379 1186
rect 1136 1182 1138 1185
rect 1286 1184 1292 1185
rect 1134 1181 1140 1182
rect 950 1179 956 1180
rect 950 1175 951 1179
rect 955 1175 956 1179
rect 950 1174 956 1175
rect 982 1179 988 1180
rect 982 1175 983 1179
rect 987 1175 988 1179
rect 1134 1177 1135 1181
rect 1139 1177 1140 1181
rect 1286 1180 1287 1184
rect 1291 1180 1292 1184
rect 1286 1179 1292 1180
rect 1326 1184 1332 1185
rect 1326 1180 1327 1184
rect 1331 1180 1332 1184
rect 1326 1179 1332 1180
rect 1366 1184 1372 1185
rect 1366 1180 1367 1184
rect 1371 1180 1372 1184
rect 1366 1179 1372 1180
rect 982 1174 988 1175
rect 1094 1176 1100 1177
rect 1134 1176 1140 1177
rect 952 1156 954 1174
rect 958 1168 964 1169
rect 958 1164 959 1168
rect 963 1164 964 1168
rect 958 1163 964 1164
rect 886 1155 892 1156
rect 886 1151 887 1155
rect 891 1151 892 1155
rect 871 1150 875 1151
rect 871 1145 875 1146
rect 879 1150 883 1151
rect 886 1150 892 1151
rect 950 1155 956 1156
rect 950 1151 951 1155
rect 955 1151 956 1155
rect 960 1151 962 1163
rect 950 1150 956 1151
rect 959 1150 963 1151
rect 879 1145 883 1146
rect 959 1145 963 1146
rect 798 1143 804 1144
rect 798 1139 799 1143
rect 803 1139 804 1143
rect 798 1138 804 1139
rect 880 1133 882 1145
rect 984 1144 986 1174
rect 1094 1172 1095 1176
rect 1099 1172 1100 1176
rect 1094 1171 1100 1172
rect 1096 1151 1098 1171
rect 1392 1168 1394 1230
rect 1424 1225 1426 1237
rect 1422 1224 1428 1225
rect 1422 1220 1423 1224
rect 1427 1220 1428 1224
rect 1422 1219 1428 1220
rect 1448 1212 1450 1238
rect 1471 1237 1475 1238
rect 1479 1242 1483 1243
rect 1479 1237 1483 1238
rect 1535 1242 1539 1243
rect 1546 1239 1547 1243
rect 1551 1239 1552 1243
rect 1546 1238 1552 1239
rect 1559 1242 1563 1243
rect 1535 1237 1539 1238
rect 1472 1225 1474 1237
rect 1498 1235 1504 1236
rect 1498 1231 1499 1235
rect 1503 1231 1504 1235
rect 1498 1230 1504 1231
rect 1470 1224 1476 1225
rect 1470 1220 1471 1224
rect 1475 1220 1476 1224
rect 1470 1219 1476 1220
rect 1500 1212 1502 1230
rect 1536 1225 1538 1237
rect 1534 1224 1540 1225
rect 1534 1220 1535 1224
rect 1539 1220 1540 1224
rect 1534 1219 1540 1220
rect 1446 1211 1452 1212
rect 1446 1207 1447 1211
rect 1451 1207 1452 1211
rect 1446 1206 1452 1207
rect 1498 1211 1504 1212
rect 1498 1207 1499 1211
rect 1503 1207 1504 1211
rect 1498 1206 1504 1207
rect 1422 1196 1428 1197
rect 1422 1192 1423 1196
rect 1427 1192 1428 1196
rect 1422 1191 1428 1192
rect 1470 1196 1476 1197
rect 1470 1192 1471 1196
rect 1475 1192 1476 1196
rect 1470 1191 1476 1192
rect 1534 1196 1540 1197
rect 1534 1192 1535 1196
rect 1539 1192 1540 1196
rect 1534 1191 1540 1192
rect 1415 1190 1419 1191
rect 1415 1185 1419 1186
rect 1423 1190 1427 1191
rect 1423 1185 1427 1186
rect 1471 1190 1475 1191
rect 1471 1185 1475 1186
rect 1527 1190 1531 1191
rect 1527 1185 1531 1186
rect 1535 1190 1539 1191
rect 1535 1185 1539 1186
rect 1548 1187 1550 1238
rect 1559 1237 1563 1238
rect 1615 1242 1619 1243
rect 1615 1237 1619 1238
rect 1639 1242 1643 1243
rect 1639 1237 1643 1238
rect 1719 1242 1723 1243
rect 1719 1237 1723 1238
rect 1799 1242 1803 1243
rect 1799 1237 1803 1238
rect 1570 1235 1576 1236
rect 1570 1231 1571 1235
rect 1575 1231 1576 1235
rect 1570 1230 1576 1231
rect 1572 1212 1574 1230
rect 1616 1225 1618 1237
rect 1720 1225 1722 1237
rect 1816 1236 1818 1270
rect 1824 1244 1826 1270
rect 1836 1252 1838 1270
rect 1878 1264 1884 1265
rect 1878 1260 1879 1264
rect 1883 1260 1884 1264
rect 1878 1259 1884 1260
rect 1834 1251 1840 1252
rect 1834 1247 1835 1251
rect 1839 1247 1840 1251
rect 1834 1246 1840 1247
rect 1822 1243 1828 1244
rect 1880 1243 1882 1259
rect 1960 1252 1962 1318
rect 1966 1308 1972 1309
rect 1966 1304 1967 1308
rect 1971 1304 1972 1308
rect 1966 1303 1972 1304
rect 2030 1308 2036 1309
rect 2030 1304 2031 1308
rect 2035 1304 2036 1308
rect 2030 1303 2036 1304
rect 1968 1299 1970 1303
rect 2032 1299 2034 1303
rect 1967 1298 1971 1299
rect 1967 1293 1971 1294
rect 2031 1298 2035 1299
rect 2031 1293 2035 1294
rect 1966 1292 1972 1293
rect 1966 1288 1967 1292
rect 1971 1288 1972 1292
rect 1966 1287 1972 1288
rect 2048 1276 2050 1342
rect 2072 1337 2074 1349
rect 2084 1348 2086 1382
rect 2092 1364 2094 1430
rect 2118 1423 2124 1424
rect 2118 1419 2119 1423
rect 2123 1419 2124 1423
rect 2118 1418 2124 1419
rect 2120 1411 2122 1418
rect 2119 1410 2123 1411
rect 2119 1405 2123 1406
rect 2120 1402 2122 1405
rect 2118 1401 2124 1402
rect 2118 1397 2119 1401
rect 2123 1397 2124 1401
rect 2118 1396 2124 1397
rect 2118 1384 2124 1385
rect 2118 1380 2119 1384
rect 2123 1380 2124 1384
rect 2118 1379 2124 1380
rect 2090 1363 2096 1364
rect 2090 1359 2091 1363
rect 2095 1359 2096 1363
rect 2090 1358 2096 1359
rect 2120 1355 2122 1379
rect 2119 1354 2123 1355
rect 2119 1349 2123 1350
rect 2082 1347 2088 1348
rect 2082 1343 2083 1347
rect 2087 1343 2088 1347
rect 2082 1342 2088 1343
rect 2070 1336 2076 1337
rect 2070 1332 2071 1336
rect 2075 1332 2076 1336
rect 2070 1331 2076 1332
rect 2120 1329 2122 1349
rect 2118 1328 2124 1329
rect 2118 1324 2119 1328
rect 2123 1324 2124 1328
rect 2082 1323 2088 1324
rect 2118 1323 2124 1324
rect 2082 1319 2083 1323
rect 2087 1319 2088 1323
rect 2082 1318 2088 1319
rect 2070 1308 2076 1309
rect 2070 1304 2071 1308
rect 2075 1304 2076 1308
rect 2070 1303 2076 1304
rect 2072 1299 2074 1303
rect 2055 1298 2059 1299
rect 2055 1293 2059 1294
rect 2071 1298 2075 1299
rect 2071 1293 2075 1294
rect 2054 1292 2060 1293
rect 2054 1288 2055 1292
rect 2059 1288 2060 1292
rect 2054 1287 2060 1288
rect 2046 1275 2052 1276
rect 2046 1271 2047 1275
rect 2051 1271 2052 1275
rect 2046 1270 2052 1271
rect 1966 1264 1972 1265
rect 1966 1260 1967 1264
rect 1971 1260 1972 1264
rect 1966 1259 1972 1260
rect 2054 1264 2060 1265
rect 2054 1260 2055 1264
rect 2059 1260 2060 1264
rect 2054 1259 2060 1260
rect 1958 1251 1964 1252
rect 1958 1247 1959 1251
rect 1963 1247 1964 1251
rect 1958 1246 1964 1247
rect 1968 1243 1970 1259
rect 2034 1251 2040 1252
rect 2034 1247 2035 1251
rect 2039 1247 2040 1251
rect 2034 1246 2040 1247
rect 1822 1239 1823 1243
rect 1827 1239 1828 1243
rect 1822 1238 1828 1239
rect 1839 1242 1843 1243
rect 1839 1237 1843 1238
rect 1879 1242 1883 1243
rect 1879 1237 1883 1238
rect 1967 1242 1971 1243
rect 1967 1237 1971 1238
rect 1814 1235 1820 1236
rect 1814 1231 1815 1235
rect 1819 1231 1820 1235
rect 1814 1230 1820 1231
rect 1840 1225 1842 1237
rect 1866 1235 1872 1236
rect 1866 1231 1867 1235
rect 1871 1231 1872 1235
rect 1866 1230 1872 1231
rect 1614 1224 1620 1225
rect 1614 1220 1615 1224
rect 1619 1220 1620 1224
rect 1614 1219 1620 1220
rect 1718 1224 1724 1225
rect 1718 1220 1719 1224
rect 1723 1220 1724 1224
rect 1718 1219 1724 1220
rect 1838 1224 1844 1225
rect 1838 1220 1839 1224
rect 1843 1220 1844 1224
rect 1838 1219 1844 1220
rect 1868 1212 1870 1230
rect 1968 1225 1970 1237
rect 1966 1224 1972 1225
rect 1966 1220 1967 1224
rect 1971 1220 1972 1224
rect 1966 1219 1972 1220
rect 1570 1211 1576 1212
rect 1570 1207 1571 1211
rect 1575 1207 1576 1211
rect 1570 1206 1576 1207
rect 1866 1211 1872 1212
rect 1866 1207 1867 1211
rect 1871 1207 1872 1211
rect 1866 1206 1872 1207
rect 1990 1211 1996 1212
rect 1990 1207 1991 1211
rect 1995 1207 1996 1211
rect 1990 1206 1996 1207
rect 1614 1196 1620 1197
rect 1614 1192 1615 1196
rect 1619 1192 1620 1196
rect 1718 1196 1724 1197
rect 1718 1192 1719 1196
rect 1723 1192 1724 1196
rect 1614 1191 1620 1192
rect 1622 1191 1628 1192
rect 1718 1191 1724 1192
rect 1838 1196 1844 1197
rect 1838 1192 1839 1196
rect 1843 1192 1844 1196
rect 1838 1191 1844 1192
rect 1966 1196 1972 1197
rect 1966 1192 1967 1196
rect 1971 1192 1972 1196
rect 1966 1191 1972 1192
rect 1583 1190 1587 1191
rect 1548 1185 1558 1187
rect 1583 1185 1587 1186
rect 1615 1190 1619 1191
rect 1622 1187 1623 1191
rect 1627 1187 1628 1191
rect 1622 1186 1628 1187
rect 1639 1190 1643 1191
rect 1615 1185 1619 1186
rect 1414 1184 1420 1185
rect 1414 1180 1415 1184
rect 1419 1180 1420 1184
rect 1414 1179 1420 1180
rect 1470 1184 1476 1185
rect 1470 1180 1471 1184
rect 1475 1180 1476 1184
rect 1470 1179 1476 1180
rect 1526 1184 1532 1185
rect 1526 1180 1527 1184
rect 1531 1180 1532 1184
rect 1526 1179 1532 1180
rect 1556 1176 1558 1185
rect 1582 1184 1588 1185
rect 1582 1180 1583 1184
rect 1587 1180 1588 1184
rect 1582 1179 1588 1180
rect 1438 1175 1444 1176
rect 1438 1171 1439 1175
rect 1443 1171 1444 1175
rect 1438 1170 1444 1171
rect 1554 1175 1560 1176
rect 1554 1171 1555 1175
rect 1559 1171 1560 1175
rect 1554 1170 1560 1171
rect 1314 1167 1320 1168
rect 1134 1164 1140 1165
rect 1134 1160 1135 1164
rect 1139 1160 1140 1164
rect 1314 1163 1315 1167
rect 1319 1163 1320 1167
rect 1314 1162 1320 1163
rect 1354 1167 1360 1168
rect 1354 1163 1355 1167
rect 1359 1163 1360 1167
rect 1354 1162 1360 1163
rect 1390 1167 1396 1168
rect 1390 1163 1391 1167
rect 1395 1163 1396 1167
rect 1390 1162 1396 1163
rect 1134 1159 1140 1160
rect 991 1150 995 1151
rect 991 1145 995 1146
rect 1095 1150 1099 1151
rect 1095 1145 1099 1146
rect 974 1143 980 1144
rect 974 1139 975 1143
rect 979 1139 980 1143
rect 974 1138 980 1139
rect 982 1143 988 1144
rect 982 1139 983 1143
rect 987 1139 988 1143
rect 982 1138 988 1139
rect 774 1132 780 1133
rect 774 1128 775 1132
rect 779 1128 780 1132
rect 774 1127 780 1128
rect 878 1132 884 1133
rect 878 1128 879 1132
rect 883 1128 884 1132
rect 878 1127 884 1128
rect 976 1120 978 1138
rect 992 1133 994 1145
rect 990 1132 996 1133
rect 990 1128 991 1132
rect 995 1128 996 1132
rect 990 1127 996 1128
rect 1096 1125 1098 1145
rect 1136 1131 1138 1159
rect 1286 1156 1292 1157
rect 1286 1152 1287 1156
rect 1291 1152 1292 1156
rect 1286 1151 1292 1152
rect 1288 1131 1290 1151
rect 1316 1144 1318 1162
rect 1326 1156 1332 1157
rect 1326 1152 1327 1156
rect 1331 1152 1332 1156
rect 1326 1151 1332 1152
rect 1314 1143 1320 1144
rect 1314 1139 1315 1143
rect 1319 1139 1320 1143
rect 1314 1138 1320 1139
rect 1328 1131 1330 1151
rect 1356 1144 1358 1162
rect 1366 1156 1372 1157
rect 1366 1152 1367 1156
rect 1371 1152 1372 1156
rect 1366 1151 1372 1152
rect 1414 1156 1420 1157
rect 1414 1152 1415 1156
rect 1419 1152 1420 1156
rect 1414 1151 1420 1152
rect 1354 1143 1360 1144
rect 1354 1139 1355 1143
rect 1359 1139 1360 1143
rect 1354 1138 1360 1139
rect 1368 1131 1370 1151
rect 1416 1131 1418 1151
rect 1440 1144 1442 1170
rect 1518 1167 1524 1168
rect 1518 1163 1519 1167
rect 1523 1163 1524 1167
rect 1518 1162 1524 1163
rect 1470 1156 1476 1157
rect 1470 1152 1471 1156
rect 1475 1152 1476 1156
rect 1470 1151 1476 1152
rect 1438 1143 1444 1144
rect 1438 1139 1439 1143
rect 1443 1139 1444 1143
rect 1438 1138 1444 1139
rect 1472 1131 1474 1151
rect 1520 1144 1522 1162
rect 1526 1156 1532 1157
rect 1526 1152 1527 1156
rect 1531 1152 1532 1156
rect 1526 1151 1532 1152
rect 1582 1156 1588 1157
rect 1582 1152 1583 1156
rect 1587 1152 1588 1156
rect 1582 1151 1588 1152
rect 1494 1143 1500 1144
rect 1494 1139 1495 1143
rect 1499 1139 1500 1143
rect 1494 1138 1500 1139
rect 1518 1143 1524 1144
rect 1518 1139 1519 1143
rect 1523 1139 1524 1143
rect 1518 1138 1524 1139
rect 1135 1130 1139 1131
rect 1135 1125 1139 1126
rect 1287 1130 1291 1131
rect 1287 1125 1291 1126
rect 1327 1130 1331 1131
rect 1327 1125 1331 1126
rect 1367 1130 1371 1131
rect 1367 1125 1371 1126
rect 1383 1130 1387 1131
rect 1383 1125 1387 1126
rect 1415 1130 1419 1131
rect 1415 1125 1419 1126
rect 1423 1130 1427 1131
rect 1423 1125 1427 1126
rect 1471 1130 1475 1131
rect 1471 1125 1475 1126
rect 1094 1124 1100 1125
rect 1094 1120 1095 1124
rect 1099 1120 1100 1124
rect 182 1119 188 1120
rect 182 1115 183 1119
rect 187 1115 188 1119
rect 182 1114 188 1115
rect 226 1119 234 1120
rect 226 1115 227 1119
rect 231 1116 234 1119
rect 286 1119 292 1120
rect 231 1115 232 1116
rect 226 1114 232 1115
rect 286 1115 287 1119
rect 291 1115 292 1119
rect 286 1114 292 1115
rect 394 1119 400 1120
rect 394 1115 395 1119
rect 399 1115 400 1119
rect 394 1114 400 1115
rect 518 1119 524 1120
rect 518 1115 519 1119
rect 523 1115 524 1119
rect 518 1114 524 1115
rect 578 1119 584 1120
rect 578 1115 579 1119
rect 583 1115 584 1119
rect 578 1114 584 1115
rect 666 1119 672 1120
rect 666 1115 667 1119
rect 671 1115 672 1119
rect 666 1114 672 1115
rect 762 1119 768 1120
rect 762 1115 763 1119
rect 767 1115 768 1119
rect 762 1114 768 1115
rect 810 1119 816 1120
rect 810 1115 811 1119
rect 815 1115 816 1119
rect 810 1114 816 1115
rect 974 1119 980 1120
rect 1094 1119 1100 1120
rect 974 1115 975 1119
rect 979 1115 980 1119
rect 974 1114 980 1115
rect 198 1104 204 1105
rect 198 1100 199 1104
rect 203 1100 204 1104
rect 198 1099 204 1100
rect 246 1104 252 1105
rect 246 1100 247 1104
rect 251 1100 252 1104
rect 246 1099 252 1100
rect 302 1104 308 1105
rect 302 1100 303 1104
rect 307 1100 308 1104
rect 302 1099 308 1100
rect 366 1104 372 1105
rect 366 1100 367 1104
rect 371 1100 372 1104
rect 366 1099 372 1100
rect 438 1104 444 1105
rect 438 1100 439 1104
rect 443 1100 444 1104
rect 438 1099 444 1100
rect 510 1104 516 1105
rect 510 1100 511 1104
rect 515 1100 516 1104
rect 510 1099 516 1100
rect 200 1091 202 1099
rect 248 1091 250 1099
rect 304 1091 306 1099
rect 368 1091 370 1099
rect 440 1091 442 1099
rect 512 1091 514 1099
rect 199 1090 203 1091
rect 199 1085 203 1086
rect 247 1090 251 1091
rect 247 1085 251 1086
rect 303 1090 307 1091
rect 303 1085 307 1086
rect 367 1090 371 1091
rect 367 1085 371 1086
rect 431 1090 435 1091
rect 431 1085 435 1086
rect 439 1090 443 1091
rect 439 1085 443 1086
rect 503 1090 507 1091
rect 503 1085 507 1086
rect 511 1090 515 1091
rect 511 1085 515 1086
rect 198 1084 204 1085
rect 198 1080 199 1084
rect 203 1080 204 1084
rect 198 1079 204 1080
rect 246 1084 252 1085
rect 246 1080 247 1084
rect 251 1080 252 1084
rect 246 1079 252 1080
rect 302 1084 308 1085
rect 302 1080 303 1084
rect 307 1080 308 1084
rect 302 1079 308 1080
rect 366 1084 372 1085
rect 366 1080 367 1084
rect 371 1080 372 1084
rect 366 1079 372 1080
rect 430 1084 436 1085
rect 430 1080 431 1084
rect 435 1080 436 1084
rect 430 1079 436 1080
rect 502 1084 508 1085
rect 502 1080 503 1084
rect 507 1080 508 1084
rect 502 1079 508 1080
rect 174 1067 180 1068
rect 110 1064 116 1065
rect 110 1060 111 1064
rect 115 1060 116 1064
rect 174 1063 175 1067
rect 179 1063 180 1067
rect 174 1062 180 1063
rect 346 1067 352 1068
rect 346 1063 347 1067
rect 351 1063 352 1067
rect 346 1062 352 1063
rect 110 1059 116 1060
rect 112 1035 114 1059
rect 198 1056 204 1057
rect 198 1052 199 1056
rect 203 1052 204 1056
rect 198 1051 204 1052
rect 246 1056 252 1057
rect 246 1052 247 1056
rect 251 1052 252 1056
rect 246 1051 252 1052
rect 302 1056 308 1057
rect 302 1052 303 1056
rect 307 1052 308 1056
rect 302 1051 308 1052
rect 200 1035 202 1051
rect 248 1035 250 1051
rect 304 1035 306 1051
rect 348 1044 350 1062
rect 366 1056 372 1057
rect 366 1052 367 1056
rect 371 1052 372 1056
rect 366 1051 372 1052
rect 430 1056 436 1057
rect 430 1052 431 1056
rect 435 1052 436 1056
rect 430 1051 436 1052
rect 502 1056 508 1057
rect 502 1052 503 1056
rect 507 1052 508 1056
rect 502 1051 508 1052
rect 346 1043 352 1044
rect 346 1039 347 1043
rect 351 1039 352 1043
rect 346 1038 352 1039
rect 368 1035 370 1051
rect 422 1043 428 1044
rect 422 1039 423 1043
rect 427 1039 428 1043
rect 422 1038 428 1039
rect 111 1034 115 1035
rect 111 1029 115 1030
rect 199 1034 203 1035
rect 199 1029 203 1030
rect 223 1034 227 1035
rect 223 1029 227 1030
rect 247 1034 251 1035
rect 247 1029 251 1030
rect 271 1034 275 1035
rect 271 1029 275 1030
rect 303 1034 307 1035
rect 303 1029 307 1030
rect 335 1034 339 1035
rect 335 1029 339 1030
rect 367 1034 371 1035
rect 367 1029 371 1030
rect 407 1034 411 1035
rect 407 1029 411 1030
rect 112 1009 114 1029
rect 224 1017 226 1029
rect 238 1027 244 1028
rect 238 1023 239 1027
rect 243 1023 244 1027
rect 238 1022 244 1023
rect 254 1027 260 1028
rect 254 1023 255 1027
rect 259 1023 260 1027
rect 254 1022 260 1023
rect 222 1016 228 1017
rect 222 1012 223 1016
rect 227 1012 228 1016
rect 222 1011 228 1012
rect 110 1008 116 1009
rect 110 1004 111 1008
rect 115 1004 116 1008
rect 110 1003 116 1004
rect 110 991 116 992
rect 110 987 111 991
rect 115 987 116 991
rect 110 986 116 987
rect 222 988 228 989
rect 112 979 114 986
rect 222 984 223 988
rect 227 984 228 988
rect 222 983 228 984
rect 224 979 226 983
rect 111 978 115 979
rect 111 973 115 974
rect 151 978 155 979
rect 151 973 155 974
rect 215 978 219 979
rect 215 973 219 974
rect 223 978 227 979
rect 223 973 227 974
rect 112 970 114 973
rect 150 972 156 973
rect 110 969 116 970
rect 110 965 111 969
rect 115 965 116 969
rect 150 968 151 972
rect 155 968 156 972
rect 150 967 156 968
rect 214 972 220 973
rect 214 968 215 972
rect 219 968 220 972
rect 214 967 220 968
rect 110 964 116 965
rect 240 964 242 1022
rect 256 1004 258 1022
rect 272 1017 274 1029
rect 336 1017 338 1029
rect 378 1027 384 1028
rect 378 1023 379 1027
rect 383 1023 384 1027
rect 378 1022 384 1023
rect 270 1016 276 1017
rect 270 1012 271 1016
rect 275 1012 276 1016
rect 270 1011 276 1012
rect 334 1016 340 1017
rect 334 1012 335 1016
rect 339 1012 340 1016
rect 334 1011 340 1012
rect 380 1004 382 1022
rect 408 1017 410 1029
rect 406 1016 412 1017
rect 406 1012 407 1016
rect 411 1012 412 1016
rect 406 1011 412 1012
rect 424 1004 426 1038
rect 432 1035 434 1051
rect 504 1035 506 1051
rect 520 1044 522 1114
rect 590 1104 596 1105
rect 590 1100 591 1104
rect 595 1100 596 1104
rect 590 1099 596 1100
rect 678 1104 684 1105
rect 678 1100 679 1104
rect 683 1100 684 1104
rect 678 1099 684 1100
rect 774 1104 780 1105
rect 774 1100 775 1104
rect 779 1100 780 1104
rect 774 1099 780 1100
rect 592 1091 594 1099
rect 680 1091 682 1099
rect 776 1091 778 1099
rect 575 1090 579 1091
rect 575 1085 579 1086
rect 591 1090 595 1091
rect 591 1085 595 1086
rect 647 1090 651 1091
rect 647 1085 651 1086
rect 679 1090 683 1091
rect 679 1085 683 1086
rect 719 1090 723 1091
rect 719 1085 723 1086
rect 775 1090 779 1091
rect 775 1085 779 1086
rect 783 1090 787 1091
rect 783 1085 787 1086
rect 574 1084 580 1085
rect 574 1080 575 1084
rect 579 1080 580 1084
rect 574 1079 580 1080
rect 646 1084 652 1085
rect 646 1080 647 1084
rect 651 1080 652 1084
rect 646 1079 652 1080
rect 718 1084 724 1085
rect 718 1080 719 1084
rect 723 1080 724 1084
rect 718 1079 724 1080
rect 782 1084 788 1085
rect 782 1080 783 1084
rect 787 1080 788 1084
rect 782 1079 788 1080
rect 566 1067 572 1068
rect 566 1063 567 1067
rect 571 1063 572 1067
rect 566 1062 572 1063
rect 638 1067 644 1068
rect 638 1063 639 1067
rect 643 1063 644 1067
rect 638 1062 644 1063
rect 654 1067 660 1068
rect 654 1063 655 1067
rect 659 1063 660 1067
rect 654 1062 660 1063
rect 774 1067 780 1068
rect 774 1063 775 1067
rect 779 1063 780 1067
rect 774 1062 780 1063
rect 568 1044 570 1062
rect 574 1056 580 1057
rect 574 1052 575 1056
rect 579 1052 580 1056
rect 574 1051 580 1052
rect 518 1043 524 1044
rect 518 1039 519 1043
rect 523 1039 524 1043
rect 518 1038 524 1039
rect 566 1043 572 1044
rect 566 1039 567 1043
rect 571 1039 572 1043
rect 566 1038 572 1039
rect 576 1035 578 1051
rect 640 1044 642 1062
rect 646 1056 652 1057
rect 646 1052 647 1056
rect 651 1052 652 1056
rect 646 1051 652 1052
rect 638 1043 644 1044
rect 638 1039 639 1043
rect 643 1039 644 1043
rect 638 1038 644 1039
rect 648 1035 650 1051
rect 431 1034 435 1035
rect 431 1029 435 1030
rect 479 1034 483 1035
rect 479 1029 483 1030
rect 503 1034 507 1035
rect 503 1029 507 1030
rect 559 1034 563 1035
rect 559 1029 563 1030
rect 575 1034 579 1035
rect 575 1029 579 1030
rect 631 1034 635 1035
rect 631 1029 635 1030
rect 647 1034 651 1035
rect 647 1029 651 1030
rect 480 1017 482 1029
rect 546 1027 552 1028
rect 546 1023 547 1027
rect 551 1023 552 1027
rect 546 1022 552 1023
rect 478 1016 484 1017
rect 478 1012 479 1016
rect 483 1012 484 1016
rect 478 1011 484 1012
rect 548 1004 550 1022
rect 560 1017 562 1029
rect 618 1027 624 1028
rect 618 1023 619 1027
rect 623 1023 624 1027
rect 618 1022 624 1023
rect 558 1016 564 1017
rect 558 1012 559 1016
rect 563 1012 564 1016
rect 558 1011 564 1012
rect 620 1004 622 1022
rect 632 1017 634 1029
rect 656 1028 658 1062
rect 718 1056 724 1057
rect 718 1052 719 1056
rect 723 1052 724 1056
rect 718 1051 724 1052
rect 720 1035 722 1051
rect 776 1044 778 1062
rect 782 1056 788 1057
rect 782 1052 783 1056
rect 787 1052 788 1056
rect 782 1051 788 1052
rect 774 1043 780 1044
rect 774 1039 775 1043
rect 779 1039 780 1043
rect 774 1038 780 1039
rect 784 1035 786 1051
rect 812 1036 814 1114
rect 1094 1107 1100 1108
rect 878 1104 884 1105
rect 878 1100 879 1104
rect 883 1100 884 1104
rect 878 1099 884 1100
rect 990 1104 996 1105
rect 990 1100 991 1104
rect 995 1100 996 1104
rect 1094 1103 1095 1107
rect 1099 1103 1100 1107
rect 1136 1105 1138 1125
rect 1384 1113 1386 1125
rect 1398 1123 1404 1124
rect 1398 1119 1399 1123
rect 1403 1119 1404 1123
rect 1398 1118 1404 1119
rect 1406 1123 1412 1124
rect 1406 1119 1407 1123
rect 1411 1119 1412 1123
rect 1406 1118 1412 1119
rect 1382 1112 1388 1113
rect 1382 1108 1383 1112
rect 1387 1108 1388 1112
rect 1382 1107 1388 1108
rect 1094 1102 1100 1103
rect 1134 1104 1140 1105
rect 990 1099 996 1100
rect 880 1091 882 1099
rect 992 1091 994 1099
rect 1096 1091 1098 1102
rect 1134 1100 1135 1104
rect 1139 1100 1140 1104
rect 1400 1101 1402 1118
rect 1134 1099 1140 1100
rect 1399 1100 1403 1101
rect 1408 1100 1410 1118
rect 1424 1113 1426 1125
rect 1450 1123 1456 1124
rect 1450 1119 1451 1123
rect 1455 1119 1456 1123
rect 1450 1118 1456 1119
rect 1422 1112 1428 1113
rect 1422 1108 1423 1112
rect 1427 1108 1428 1112
rect 1422 1107 1428 1108
rect 1452 1100 1454 1118
rect 1472 1113 1474 1125
rect 1470 1112 1476 1113
rect 1470 1108 1471 1112
rect 1475 1108 1476 1112
rect 1470 1107 1476 1108
rect 1496 1100 1498 1138
rect 1528 1131 1530 1151
rect 1584 1131 1586 1151
rect 1624 1144 1626 1186
rect 1639 1185 1643 1186
rect 1703 1190 1707 1191
rect 1703 1185 1707 1186
rect 1719 1190 1723 1191
rect 1719 1185 1723 1186
rect 1767 1190 1771 1191
rect 1767 1185 1771 1186
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1919 1190 1923 1191
rect 1919 1185 1923 1186
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 1638 1184 1644 1185
rect 1638 1180 1639 1184
rect 1643 1180 1644 1184
rect 1638 1179 1644 1180
rect 1702 1184 1708 1185
rect 1702 1180 1703 1184
rect 1707 1180 1708 1184
rect 1702 1179 1708 1180
rect 1766 1184 1772 1185
rect 1766 1180 1767 1184
rect 1771 1180 1772 1184
rect 1766 1179 1772 1180
rect 1838 1184 1844 1185
rect 1838 1180 1839 1184
rect 1843 1180 1844 1184
rect 1838 1179 1844 1180
rect 1918 1184 1924 1185
rect 1918 1180 1919 1184
rect 1923 1180 1924 1184
rect 1918 1179 1924 1180
rect 1992 1176 1994 1206
rect 2007 1190 2011 1191
rect 2007 1185 2011 1186
rect 2006 1184 2012 1185
rect 2006 1180 2007 1184
rect 2011 1180 2012 1184
rect 2006 1179 2012 1180
rect 1990 1175 1996 1176
rect 1990 1171 1991 1175
rect 1995 1171 1996 1175
rect 1990 1170 1996 1171
rect 2036 1168 2038 1246
rect 2056 1243 2058 1259
rect 2055 1242 2059 1243
rect 2055 1237 2059 1238
rect 2071 1242 2075 1243
rect 2071 1237 2075 1238
rect 2072 1225 2074 1237
rect 2084 1236 2086 1318
rect 2118 1311 2124 1312
rect 2118 1307 2119 1311
rect 2123 1307 2124 1311
rect 2118 1306 2124 1307
rect 2120 1299 2122 1306
rect 2119 1298 2123 1299
rect 2119 1293 2123 1294
rect 2120 1290 2122 1293
rect 2118 1289 2124 1290
rect 2118 1285 2119 1289
rect 2123 1285 2124 1289
rect 2118 1284 2124 1285
rect 2118 1272 2124 1273
rect 2118 1268 2119 1272
rect 2123 1268 2124 1272
rect 2118 1267 2124 1268
rect 2120 1243 2122 1267
rect 2119 1242 2123 1243
rect 2119 1237 2123 1238
rect 2082 1235 2088 1236
rect 2082 1231 2083 1235
rect 2087 1231 2088 1235
rect 2082 1230 2088 1231
rect 2070 1224 2076 1225
rect 2070 1220 2071 1224
rect 2075 1220 2076 1224
rect 2070 1219 2076 1220
rect 2120 1217 2122 1237
rect 2118 1216 2124 1217
rect 2118 1212 2119 1216
rect 2123 1212 2124 1216
rect 2086 1211 2092 1212
rect 2118 1211 2124 1212
rect 2086 1207 2087 1211
rect 2091 1207 2092 1211
rect 2086 1206 2092 1207
rect 2070 1196 2076 1197
rect 2070 1192 2071 1196
rect 2075 1192 2076 1196
rect 2070 1191 2076 1192
rect 2071 1190 2075 1191
rect 2071 1185 2075 1186
rect 2070 1184 2076 1185
rect 2070 1180 2071 1184
rect 2075 1180 2076 1184
rect 2070 1179 2076 1180
rect 1630 1167 1636 1168
rect 1630 1163 1631 1167
rect 1635 1163 1636 1167
rect 1630 1162 1636 1163
rect 1694 1167 1700 1168
rect 1694 1163 1695 1167
rect 1699 1163 1700 1167
rect 1694 1162 1700 1163
rect 1758 1167 1764 1168
rect 1758 1163 1759 1167
rect 1763 1163 1764 1167
rect 1758 1162 1764 1163
rect 1830 1167 1836 1168
rect 1830 1163 1831 1167
rect 1835 1163 1836 1167
rect 1830 1162 1836 1163
rect 1910 1167 1916 1168
rect 1910 1163 1911 1167
rect 1915 1163 1916 1167
rect 1910 1162 1916 1163
rect 1934 1167 1940 1168
rect 1934 1163 1935 1167
rect 1939 1163 1940 1167
rect 1934 1162 1940 1163
rect 2034 1167 2040 1168
rect 2034 1163 2035 1167
rect 2039 1163 2040 1167
rect 2034 1162 2040 1163
rect 2078 1167 2084 1168
rect 2078 1163 2079 1167
rect 2083 1163 2084 1167
rect 2078 1162 2084 1163
rect 1632 1144 1634 1162
rect 1638 1156 1644 1157
rect 1638 1152 1639 1156
rect 1643 1152 1644 1156
rect 1638 1151 1644 1152
rect 1622 1143 1628 1144
rect 1622 1139 1623 1143
rect 1627 1139 1628 1143
rect 1622 1138 1628 1139
rect 1630 1143 1636 1144
rect 1630 1139 1631 1143
rect 1635 1139 1636 1143
rect 1630 1138 1636 1139
rect 1640 1131 1642 1151
rect 1696 1144 1698 1162
rect 1702 1156 1708 1157
rect 1702 1152 1703 1156
rect 1707 1152 1708 1156
rect 1702 1151 1708 1152
rect 1694 1143 1700 1144
rect 1694 1139 1695 1143
rect 1699 1139 1700 1143
rect 1694 1138 1700 1139
rect 1678 1131 1684 1132
rect 1704 1131 1706 1151
rect 1760 1144 1762 1162
rect 1766 1156 1772 1157
rect 1766 1152 1767 1156
rect 1771 1152 1772 1156
rect 1766 1151 1772 1152
rect 1758 1143 1764 1144
rect 1758 1139 1759 1143
rect 1763 1139 1764 1143
rect 1758 1138 1764 1139
rect 1768 1131 1770 1151
rect 1832 1144 1834 1162
rect 1838 1156 1844 1157
rect 1838 1152 1839 1156
rect 1843 1152 1844 1156
rect 1838 1151 1844 1152
rect 1830 1143 1836 1144
rect 1830 1139 1831 1143
rect 1835 1139 1836 1143
rect 1830 1138 1836 1139
rect 1840 1131 1842 1151
rect 1912 1144 1914 1162
rect 1918 1156 1924 1157
rect 1918 1152 1919 1156
rect 1923 1152 1924 1156
rect 1918 1151 1924 1152
rect 1910 1143 1916 1144
rect 1910 1139 1911 1143
rect 1915 1139 1916 1143
rect 1910 1138 1916 1139
rect 1920 1131 1922 1151
rect 1936 1132 1938 1162
rect 2006 1156 2012 1157
rect 2006 1152 2007 1156
rect 2011 1152 2012 1156
rect 2006 1151 2012 1152
rect 2070 1156 2076 1157
rect 2070 1152 2071 1156
rect 2075 1152 2076 1156
rect 2070 1151 2076 1152
rect 1934 1131 1940 1132
rect 2008 1131 2010 1151
rect 2054 1143 2060 1144
rect 2054 1139 2055 1143
rect 2059 1139 2060 1143
rect 2054 1138 2060 1139
rect 1527 1130 1531 1131
rect 1527 1125 1531 1126
rect 1583 1130 1587 1131
rect 1583 1125 1587 1126
rect 1591 1130 1595 1131
rect 1591 1125 1595 1126
rect 1639 1130 1643 1131
rect 1639 1125 1643 1126
rect 1655 1130 1659 1131
rect 1678 1127 1679 1131
rect 1683 1127 1684 1131
rect 1678 1126 1684 1127
rect 1703 1130 1707 1131
rect 1655 1125 1659 1126
rect 1528 1113 1530 1125
rect 1592 1113 1594 1125
rect 1598 1123 1604 1124
rect 1598 1119 1599 1123
rect 1603 1119 1604 1123
rect 1598 1118 1604 1119
rect 1618 1123 1624 1124
rect 1618 1119 1619 1123
rect 1623 1119 1624 1123
rect 1618 1118 1624 1119
rect 1526 1112 1532 1113
rect 1526 1108 1527 1112
rect 1531 1108 1532 1112
rect 1526 1107 1532 1108
rect 1590 1112 1596 1113
rect 1590 1108 1591 1112
rect 1595 1108 1596 1112
rect 1590 1107 1596 1108
rect 1551 1100 1555 1101
rect 1399 1095 1403 1096
rect 1406 1099 1412 1100
rect 1406 1095 1407 1099
rect 1411 1095 1412 1099
rect 1406 1094 1412 1095
rect 1450 1099 1456 1100
rect 1450 1095 1451 1099
rect 1455 1095 1456 1099
rect 1450 1094 1456 1095
rect 1494 1099 1500 1100
rect 1494 1095 1495 1099
rect 1499 1095 1500 1099
rect 1494 1094 1500 1095
rect 1550 1095 1551 1100
rect 1555 1095 1556 1100
rect 1550 1094 1556 1095
rect 839 1090 843 1091
rect 839 1085 843 1086
rect 879 1090 883 1091
rect 879 1085 883 1086
rect 895 1090 899 1091
rect 895 1085 899 1086
rect 951 1090 955 1091
rect 951 1085 955 1086
rect 991 1090 995 1091
rect 991 1085 995 1086
rect 1007 1090 1011 1091
rect 1007 1085 1011 1086
rect 1047 1090 1051 1091
rect 1047 1085 1051 1086
rect 1095 1090 1099 1091
rect 1095 1085 1099 1086
rect 1134 1087 1140 1088
rect 838 1084 844 1085
rect 838 1080 839 1084
rect 843 1080 844 1084
rect 838 1079 844 1080
rect 894 1084 900 1085
rect 894 1080 895 1084
rect 899 1080 900 1084
rect 894 1079 900 1080
rect 950 1084 956 1085
rect 950 1080 951 1084
rect 955 1080 956 1084
rect 950 1079 956 1080
rect 1006 1084 1012 1085
rect 1006 1080 1007 1084
rect 1011 1080 1012 1084
rect 1006 1079 1012 1080
rect 1046 1084 1052 1085
rect 1046 1080 1047 1084
rect 1051 1080 1052 1084
rect 1096 1082 1098 1085
rect 1134 1083 1135 1087
rect 1139 1083 1140 1087
rect 1134 1082 1140 1083
rect 1382 1084 1388 1085
rect 1046 1079 1052 1080
rect 1094 1081 1100 1082
rect 1094 1077 1095 1081
rect 1099 1077 1100 1081
rect 1136 1079 1138 1082
rect 1382 1080 1383 1084
rect 1387 1080 1388 1084
rect 1382 1079 1388 1080
rect 1422 1084 1428 1085
rect 1422 1080 1423 1084
rect 1427 1080 1428 1084
rect 1422 1079 1428 1080
rect 1470 1084 1476 1085
rect 1470 1080 1471 1084
rect 1475 1080 1476 1084
rect 1470 1079 1476 1080
rect 1526 1084 1532 1085
rect 1526 1080 1527 1084
rect 1531 1080 1532 1084
rect 1526 1079 1532 1080
rect 1590 1084 1596 1085
rect 1590 1080 1591 1084
rect 1595 1080 1596 1084
rect 1590 1079 1596 1080
rect 1094 1076 1100 1077
rect 1135 1078 1139 1079
rect 1135 1073 1139 1074
rect 1159 1078 1163 1079
rect 1159 1073 1163 1074
rect 1247 1078 1251 1079
rect 1247 1073 1251 1074
rect 1359 1078 1363 1079
rect 1359 1073 1363 1074
rect 1383 1078 1387 1079
rect 1383 1073 1387 1074
rect 1423 1078 1427 1079
rect 1423 1073 1427 1074
rect 1471 1078 1475 1079
rect 1471 1073 1475 1074
rect 1527 1078 1531 1079
rect 1527 1073 1531 1074
rect 1575 1078 1579 1079
rect 1575 1073 1579 1074
rect 1591 1078 1595 1079
rect 1591 1073 1595 1074
rect 1136 1070 1138 1073
rect 1158 1072 1164 1073
rect 1134 1069 1140 1070
rect 830 1067 836 1068
rect 830 1063 831 1067
rect 835 1063 836 1067
rect 830 1062 836 1063
rect 910 1067 916 1068
rect 910 1063 911 1067
rect 915 1063 916 1067
rect 910 1062 916 1063
rect 942 1067 948 1068
rect 942 1063 943 1067
rect 947 1063 948 1067
rect 942 1062 948 1063
rect 998 1067 1004 1068
rect 998 1063 999 1067
rect 1003 1063 1004 1067
rect 998 1062 1004 1063
rect 1034 1067 1040 1068
rect 1034 1063 1035 1067
rect 1039 1063 1040 1067
rect 1034 1062 1040 1063
rect 1086 1067 1092 1068
rect 1086 1063 1087 1067
rect 1091 1063 1092 1067
rect 1134 1065 1135 1069
rect 1139 1065 1140 1069
rect 1158 1068 1159 1072
rect 1163 1068 1164 1072
rect 1158 1067 1164 1068
rect 1246 1072 1252 1073
rect 1246 1068 1247 1072
rect 1251 1068 1252 1072
rect 1246 1067 1252 1068
rect 1358 1072 1364 1073
rect 1358 1068 1359 1072
rect 1363 1068 1364 1072
rect 1358 1067 1364 1068
rect 1470 1072 1476 1073
rect 1470 1068 1471 1072
rect 1475 1068 1476 1072
rect 1470 1067 1476 1068
rect 1574 1072 1580 1073
rect 1574 1068 1575 1072
rect 1579 1068 1580 1072
rect 1574 1067 1580 1068
rect 1086 1062 1092 1063
rect 1094 1064 1100 1065
rect 1134 1064 1140 1065
rect 832 1044 834 1062
rect 838 1056 844 1057
rect 838 1052 839 1056
rect 843 1052 844 1056
rect 838 1051 844 1052
rect 894 1056 900 1057
rect 894 1052 895 1056
rect 899 1052 900 1056
rect 894 1051 900 1052
rect 830 1043 836 1044
rect 830 1039 831 1043
rect 835 1039 836 1043
rect 830 1038 836 1039
rect 810 1035 816 1036
rect 840 1035 842 1051
rect 896 1035 898 1051
rect 703 1034 707 1035
rect 703 1029 707 1030
rect 719 1034 723 1035
rect 719 1029 723 1030
rect 775 1034 779 1035
rect 775 1029 779 1030
rect 783 1034 787 1035
rect 810 1031 811 1035
rect 815 1031 816 1035
rect 810 1030 816 1031
rect 839 1034 843 1035
rect 783 1029 787 1030
rect 839 1029 843 1030
rect 895 1034 899 1035
rect 895 1029 899 1030
rect 903 1034 907 1035
rect 903 1029 907 1030
rect 654 1027 660 1028
rect 654 1023 655 1027
rect 659 1023 660 1027
rect 654 1022 660 1023
rect 704 1017 706 1029
rect 710 1027 716 1028
rect 710 1023 711 1027
rect 715 1023 716 1027
rect 710 1022 716 1023
rect 730 1027 736 1028
rect 730 1023 731 1027
rect 735 1023 736 1027
rect 730 1022 736 1023
rect 630 1016 636 1017
rect 630 1012 631 1016
rect 635 1012 636 1016
rect 630 1011 636 1012
rect 702 1016 708 1017
rect 702 1012 703 1016
rect 707 1012 708 1016
rect 702 1011 708 1012
rect 250 1003 258 1004
rect 250 999 251 1003
rect 255 1000 258 1003
rect 378 1003 384 1004
rect 255 999 256 1000
rect 250 998 256 999
rect 378 999 379 1003
rect 383 999 384 1003
rect 378 998 384 999
rect 422 1003 428 1004
rect 422 999 423 1003
rect 427 999 428 1003
rect 422 998 428 999
rect 518 1003 524 1004
rect 518 999 519 1003
rect 523 999 524 1003
rect 518 998 524 999
rect 546 1003 552 1004
rect 546 999 547 1003
rect 551 999 552 1003
rect 546 998 552 999
rect 618 1003 624 1004
rect 618 999 619 1003
rect 623 999 624 1003
rect 618 998 624 999
rect 270 988 276 989
rect 270 984 271 988
rect 275 984 276 988
rect 270 983 276 984
rect 334 988 340 989
rect 334 984 335 988
rect 339 984 340 988
rect 334 983 340 984
rect 406 988 412 989
rect 406 984 407 988
rect 411 984 412 988
rect 406 983 412 984
rect 478 988 484 989
rect 478 984 479 988
rect 483 984 484 988
rect 478 983 484 984
rect 272 979 274 983
rect 336 979 338 983
rect 408 979 410 983
rect 480 979 482 983
rect 271 978 275 979
rect 271 973 275 974
rect 287 978 291 979
rect 287 973 291 974
rect 335 978 339 979
rect 335 973 339 974
rect 367 978 371 979
rect 367 973 371 974
rect 407 978 411 979
rect 407 973 411 974
rect 447 978 451 979
rect 447 973 451 974
rect 479 978 483 979
rect 479 973 483 974
rect 286 972 292 973
rect 286 968 287 972
rect 291 968 292 972
rect 286 967 292 968
rect 366 972 372 973
rect 366 968 367 972
rect 371 968 372 972
rect 366 967 372 968
rect 446 972 452 973
rect 446 968 447 972
rect 451 968 452 972
rect 446 967 452 968
rect 238 963 244 964
rect 238 959 239 963
rect 243 959 244 963
rect 238 958 244 959
rect 206 955 212 956
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 206 951 207 955
rect 211 951 212 955
rect 206 950 212 951
rect 278 955 284 956
rect 278 951 279 955
rect 283 951 284 955
rect 278 950 284 951
rect 358 955 364 956
rect 358 951 359 955
rect 363 951 364 955
rect 358 950 364 951
rect 470 955 476 956
rect 470 951 471 955
rect 475 951 476 955
rect 470 950 476 951
rect 482 955 488 956
rect 482 951 483 955
rect 487 951 488 955
rect 482 950 488 951
rect 110 947 116 948
rect 112 927 114 947
rect 150 944 156 945
rect 150 940 151 944
rect 155 940 156 944
rect 150 939 156 940
rect 152 927 154 939
rect 208 932 210 950
rect 214 944 220 945
rect 214 940 215 944
rect 219 940 220 944
rect 214 939 220 940
rect 158 931 164 932
rect 158 927 159 931
rect 163 927 164 931
rect 206 931 212 932
rect 206 927 207 931
rect 211 927 212 931
rect 216 927 218 939
rect 280 932 282 950
rect 286 944 292 945
rect 286 940 287 944
rect 291 940 292 944
rect 286 939 292 940
rect 278 931 284 932
rect 278 927 279 931
rect 283 927 284 931
rect 288 927 290 939
rect 360 932 362 950
rect 366 944 372 945
rect 366 940 367 944
rect 371 940 372 944
rect 366 939 372 940
rect 446 944 452 945
rect 446 940 447 944
rect 451 940 452 944
rect 446 939 452 940
rect 358 931 364 932
rect 358 927 359 931
rect 363 927 364 931
rect 368 927 370 939
rect 448 927 450 939
rect 111 926 115 927
rect 111 921 115 922
rect 135 926 139 927
rect 135 921 139 922
rect 151 926 155 927
rect 158 926 164 927
rect 183 926 187 927
rect 206 926 212 927
rect 215 926 219 927
rect 151 921 155 922
rect 112 901 114 921
rect 136 909 138 921
rect 134 908 140 909
rect 134 904 135 908
rect 139 904 140 908
rect 134 903 140 904
rect 110 900 116 901
rect 110 896 111 900
rect 115 896 116 900
rect 160 896 162 926
rect 183 921 187 922
rect 215 921 219 922
rect 255 926 259 927
rect 278 926 284 927
rect 287 926 291 927
rect 255 921 259 922
rect 287 921 291 922
rect 327 926 331 927
rect 358 926 364 927
rect 367 926 371 927
rect 327 921 331 922
rect 367 921 371 922
rect 399 926 403 927
rect 399 921 403 922
rect 447 926 451 927
rect 447 921 451 922
rect 463 926 467 927
rect 463 921 467 922
rect 170 919 176 920
rect 170 915 171 919
rect 175 915 176 919
rect 170 914 176 915
rect 172 896 174 914
rect 184 909 186 921
rect 242 919 248 920
rect 242 915 243 919
rect 247 915 248 919
rect 242 914 248 915
rect 182 908 188 909
rect 182 904 183 908
rect 187 904 188 908
rect 182 903 188 904
rect 244 896 246 914
rect 256 909 258 921
rect 302 919 308 920
rect 302 915 303 919
rect 307 915 308 919
rect 302 914 308 915
rect 254 908 260 909
rect 254 904 255 908
rect 259 904 260 908
rect 254 903 260 904
rect 110 895 116 896
rect 158 895 164 896
rect 158 891 159 895
rect 163 891 164 895
rect 158 890 164 891
rect 170 895 176 896
rect 170 891 171 895
rect 175 891 176 895
rect 170 890 176 891
rect 242 895 248 896
rect 242 891 243 895
rect 247 891 248 895
rect 242 890 248 891
rect 110 883 116 884
rect 110 879 111 883
rect 115 879 116 883
rect 110 878 116 879
rect 134 880 140 881
rect 112 871 114 878
rect 134 876 135 880
rect 139 876 140 880
rect 134 875 140 876
rect 182 880 188 881
rect 182 876 183 880
rect 187 876 188 880
rect 182 875 188 876
rect 254 880 260 881
rect 254 876 255 880
rect 259 876 260 880
rect 254 875 260 876
rect 136 871 138 875
rect 184 871 186 875
rect 256 871 258 875
rect 111 870 115 871
rect 111 865 115 866
rect 135 870 139 871
rect 135 865 139 866
rect 175 870 179 871
rect 175 865 179 866
rect 183 870 187 871
rect 183 865 187 866
rect 215 870 219 871
rect 215 865 219 866
rect 255 870 259 871
rect 255 865 259 866
rect 279 870 283 871
rect 279 865 283 866
rect 112 862 114 865
rect 134 864 140 865
rect 110 861 116 862
rect 110 857 111 861
rect 115 857 116 861
rect 134 860 135 864
rect 139 860 140 864
rect 134 859 140 860
rect 174 864 180 865
rect 174 860 175 864
rect 179 860 180 864
rect 174 859 180 860
rect 214 864 220 865
rect 214 860 215 864
rect 219 860 220 864
rect 214 859 220 860
rect 278 864 284 865
rect 278 860 279 864
rect 283 860 284 864
rect 278 859 284 860
rect 110 856 116 857
rect 304 848 306 914
rect 328 909 330 921
rect 386 919 392 920
rect 386 915 387 919
rect 391 915 392 919
rect 386 914 392 915
rect 326 908 332 909
rect 326 904 327 908
rect 331 904 332 908
rect 326 903 332 904
rect 388 896 390 914
rect 400 909 402 921
rect 464 909 466 921
rect 472 920 474 950
rect 484 932 486 950
rect 520 932 522 998
rect 558 988 564 989
rect 558 984 559 988
rect 563 984 564 988
rect 558 983 564 984
rect 630 988 636 989
rect 630 984 631 988
rect 635 984 636 988
rect 630 983 636 984
rect 702 988 708 989
rect 702 984 703 988
rect 707 984 708 988
rect 702 983 708 984
rect 560 979 562 983
rect 632 979 634 983
rect 704 979 706 983
rect 527 978 531 979
rect 527 973 531 974
rect 559 978 563 979
rect 559 973 563 974
rect 599 978 603 979
rect 599 973 603 974
rect 631 978 635 979
rect 631 973 635 974
rect 671 978 675 979
rect 671 973 675 974
rect 703 978 707 979
rect 703 973 707 974
rect 526 972 532 973
rect 526 968 527 972
rect 531 968 532 972
rect 526 967 532 968
rect 598 972 604 973
rect 598 968 599 972
rect 603 968 604 972
rect 598 967 604 968
rect 670 972 676 973
rect 670 968 671 972
rect 675 968 676 972
rect 670 967 676 968
rect 712 964 714 1022
rect 732 1004 734 1022
rect 776 1017 778 1029
rect 802 1027 808 1028
rect 802 1023 803 1027
rect 807 1023 808 1027
rect 802 1022 808 1023
rect 774 1016 780 1017
rect 774 1012 775 1016
rect 779 1012 780 1016
rect 774 1011 780 1012
rect 804 1004 806 1022
rect 840 1017 842 1029
rect 866 1027 872 1028
rect 866 1023 867 1027
rect 871 1023 872 1027
rect 866 1022 872 1023
rect 838 1016 844 1017
rect 838 1012 839 1016
rect 843 1012 844 1016
rect 838 1011 844 1012
rect 868 1004 870 1022
rect 904 1017 906 1029
rect 912 1028 914 1062
rect 944 1044 946 1062
rect 950 1056 956 1057
rect 950 1052 951 1056
rect 955 1052 956 1056
rect 950 1051 956 1052
rect 926 1043 932 1044
rect 926 1039 927 1043
rect 931 1039 932 1043
rect 926 1038 932 1039
rect 942 1043 948 1044
rect 942 1039 943 1043
rect 947 1039 948 1043
rect 942 1038 948 1039
rect 910 1027 916 1028
rect 910 1023 911 1027
rect 915 1023 916 1027
rect 910 1022 916 1023
rect 902 1016 908 1017
rect 902 1012 903 1016
rect 907 1012 908 1016
rect 902 1011 908 1012
rect 928 1004 930 1038
rect 952 1035 954 1051
rect 1000 1044 1002 1062
rect 1006 1056 1012 1057
rect 1006 1052 1007 1056
rect 1011 1052 1012 1056
rect 1006 1051 1012 1052
rect 998 1043 1004 1044
rect 998 1039 999 1043
rect 1003 1039 1004 1043
rect 998 1038 1004 1039
rect 1008 1035 1010 1051
rect 1036 1044 1038 1062
rect 1046 1056 1052 1057
rect 1046 1052 1047 1056
rect 1051 1052 1052 1056
rect 1046 1051 1052 1052
rect 1034 1043 1040 1044
rect 1034 1039 1035 1043
rect 1039 1039 1040 1043
rect 1034 1038 1040 1039
rect 1048 1035 1050 1051
rect 951 1034 955 1035
rect 951 1029 955 1030
rect 967 1034 971 1035
rect 967 1029 971 1030
rect 1007 1034 1011 1035
rect 1007 1029 1011 1030
rect 1039 1034 1043 1035
rect 1039 1029 1043 1030
rect 1047 1034 1051 1035
rect 1088 1032 1090 1062
rect 1094 1060 1095 1064
rect 1099 1060 1100 1064
rect 1094 1059 1100 1060
rect 1174 1059 1180 1060
rect 1096 1035 1098 1059
rect 1174 1055 1175 1059
rect 1179 1055 1180 1059
rect 1600 1056 1602 1118
rect 1620 1100 1622 1118
rect 1656 1113 1658 1125
rect 1654 1112 1660 1113
rect 1654 1108 1655 1112
rect 1659 1108 1660 1112
rect 1654 1107 1660 1108
rect 1680 1100 1682 1126
rect 1703 1125 1707 1126
rect 1711 1130 1715 1131
rect 1711 1125 1715 1126
rect 1767 1130 1771 1131
rect 1767 1125 1771 1126
rect 1823 1130 1827 1131
rect 1823 1125 1827 1126
rect 1839 1130 1843 1131
rect 1839 1125 1843 1126
rect 1871 1130 1875 1131
rect 1871 1125 1875 1126
rect 1919 1130 1923 1131
rect 1919 1125 1923 1126
rect 1927 1130 1931 1131
rect 1934 1127 1935 1131
rect 1939 1127 1940 1131
rect 1934 1126 1940 1127
rect 1983 1130 1987 1131
rect 1927 1125 1931 1126
rect 1983 1125 1987 1126
rect 2007 1130 2011 1131
rect 2007 1125 2011 1126
rect 2031 1130 2035 1131
rect 2031 1125 2035 1126
rect 1712 1113 1714 1125
rect 1738 1123 1744 1124
rect 1738 1119 1739 1123
rect 1743 1119 1744 1123
rect 1738 1118 1744 1119
rect 1710 1112 1716 1113
rect 1710 1108 1711 1112
rect 1715 1108 1716 1112
rect 1710 1107 1716 1108
rect 1740 1100 1742 1118
rect 1768 1113 1770 1125
rect 1794 1123 1800 1124
rect 1794 1119 1795 1123
rect 1799 1119 1800 1123
rect 1794 1118 1800 1119
rect 1766 1112 1772 1113
rect 1766 1108 1767 1112
rect 1771 1108 1772 1112
rect 1766 1107 1772 1108
rect 1796 1100 1798 1118
rect 1824 1113 1826 1125
rect 1850 1123 1856 1124
rect 1850 1119 1851 1123
rect 1855 1119 1856 1123
rect 1850 1118 1856 1119
rect 1822 1112 1828 1113
rect 1822 1108 1823 1112
rect 1827 1108 1828 1112
rect 1822 1107 1828 1108
rect 1852 1100 1854 1118
rect 1872 1113 1874 1125
rect 1898 1123 1904 1124
rect 1898 1119 1899 1123
rect 1903 1119 1904 1123
rect 1898 1118 1904 1119
rect 1870 1112 1876 1113
rect 1870 1108 1871 1112
rect 1875 1108 1876 1112
rect 1870 1107 1876 1108
rect 1900 1100 1902 1118
rect 1928 1113 1930 1125
rect 1954 1123 1960 1124
rect 1954 1119 1955 1123
rect 1959 1119 1960 1123
rect 1954 1118 1960 1119
rect 1926 1112 1932 1113
rect 1926 1108 1927 1112
rect 1931 1108 1932 1112
rect 1926 1107 1932 1108
rect 1956 1100 1958 1118
rect 1984 1113 1986 1125
rect 2032 1113 2034 1125
rect 2046 1123 2052 1124
rect 2046 1119 2047 1123
rect 2051 1119 2052 1123
rect 2046 1118 2052 1119
rect 1982 1112 1988 1113
rect 1982 1108 1983 1112
rect 1987 1108 1988 1112
rect 1982 1107 1988 1108
rect 2030 1112 2036 1113
rect 2030 1108 2031 1112
rect 2035 1108 2036 1112
rect 2030 1107 2036 1108
rect 1618 1099 1624 1100
rect 1618 1095 1619 1099
rect 1623 1095 1624 1099
rect 1618 1094 1624 1095
rect 1678 1099 1684 1100
rect 1678 1095 1679 1099
rect 1683 1095 1684 1099
rect 1678 1094 1684 1095
rect 1738 1099 1744 1100
rect 1738 1095 1739 1099
rect 1743 1095 1744 1099
rect 1738 1094 1744 1095
rect 1794 1099 1800 1100
rect 1794 1095 1795 1099
rect 1799 1095 1800 1099
rect 1794 1094 1800 1095
rect 1850 1099 1856 1100
rect 1850 1095 1851 1099
rect 1855 1095 1856 1099
rect 1850 1094 1856 1095
rect 1898 1099 1904 1100
rect 1898 1095 1899 1099
rect 1903 1095 1904 1099
rect 1898 1094 1904 1095
rect 1954 1099 1960 1100
rect 1954 1095 1955 1099
rect 1959 1095 1960 1099
rect 1954 1094 1960 1095
rect 1998 1099 2004 1100
rect 1998 1095 1999 1099
rect 2003 1095 2004 1099
rect 1998 1094 2004 1095
rect 1654 1084 1660 1085
rect 1654 1080 1655 1084
rect 1659 1080 1660 1084
rect 1654 1079 1660 1080
rect 1710 1084 1716 1085
rect 1710 1080 1711 1084
rect 1715 1080 1716 1084
rect 1710 1079 1716 1080
rect 1766 1084 1772 1085
rect 1766 1080 1767 1084
rect 1771 1080 1772 1084
rect 1766 1079 1772 1080
rect 1822 1084 1828 1085
rect 1822 1080 1823 1084
rect 1827 1080 1828 1084
rect 1822 1079 1828 1080
rect 1870 1084 1876 1085
rect 1870 1080 1871 1084
rect 1875 1080 1876 1084
rect 1870 1079 1876 1080
rect 1926 1084 1932 1085
rect 1926 1080 1927 1084
rect 1931 1080 1932 1084
rect 1926 1079 1932 1080
rect 1982 1084 1988 1085
rect 1982 1080 1983 1084
rect 1987 1080 1988 1084
rect 1982 1079 1988 1080
rect 1655 1078 1659 1079
rect 1655 1073 1659 1074
rect 1671 1078 1675 1079
rect 1671 1073 1675 1074
rect 1711 1078 1715 1079
rect 1711 1073 1715 1074
rect 1759 1078 1763 1079
rect 1759 1073 1763 1074
rect 1767 1078 1771 1079
rect 1767 1073 1771 1074
rect 1823 1078 1827 1079
rect 1823 1073 1827 1074
rect 1847 1078 1851 1079
rect 1847 1073 1851 1074
rect 1871 1078 1875 1079
rect 1871 1073 1875 1074
rect 1927 1078 1931 1079
rect 1927 1073 1931 1074
rect 1983 1078 1987 1079
rect 1983 1073 1987 1074
rect 1670 1072 1676 1073
rect 1670 1068 1671 1072
rect 1675 1068 1676 1072
rect 1670 1067 1676 1068
rect 1758 1072 1764 1073
rect 1758 1068 1759 1072
rect 1763 1068 1764 1072
rect 1758 1067 1764 1068
rect 1846 1072 1852 1073
rect 1846 1068 1847 1072
rect 1851 1068 1852 1072
rect 1846 1067 1852 1068
rect 1926 1072 1932 1073
rect 1926 1068 1927 1072
rect 1931 1068 1932 1072
rect 1926 1067 1932 1068
rect 1702 1063 1708 1064
rect 1702 1059 1703 1063
rect 1707 1059 1708 1063
rect 1702 1058 1708 1059
rect 1174 1054 1180 1055
rect 1238 1055 1244 1056
rect 1134 1052 1140 1053
rect 1134 1048 1135 1052
rect 1139 1048 1140 1052
rect 1134 1047 1140 1048
rect 1095 1034 1099 1035
rect 1047 1029 1051 1030
rect 1086 1031 1092 1032
rect 968 1017 970 1029
rect 994 1027 1000 1028
rect 994 1023 995 1027
rect 999 1023 1000 1027
rect 994 1022 1000 1023
rect 966 1016 972 1017
rect 966 1012 967 1016
rect 971 1012 972 1016
rect 966 1011 972 1012
rect 996 1004 998 1022
rect 1040 1017 1042 1029
rect 1086 1027 1087 1031
rect 1091 1027 1092 1031
rect 1095 1029 1099 1030
rect 1086 1026 1092 1027
rect 1038 1016 1044 1017
rect 1038 1012 1039 1016
rect 1043 1012 1044 1016
rect 1038 1011 1044 1012
rect 1096 1009 1098 1029
rect 1136 1027 1138 1047
rect 1158 1044 1164 1045
rect 1158 1040 1159 1044
rect 1163 1040 1164 1044
rect 1158 1039 1164 1040
rect 1160 1027 1162 1039
rect 1135 1026 1139 1027
rect 1135 1021 1139 1022
rect 1159 1026 1163 1027
rect 1159 1021 1163 1022
rect 1094 1008 1100 1009
rect 1094 1004 1095 1008
rect 1099 1004 1100 1008
rect 730 1003 736 1004
rect 730 999 731 1003
rect 735 999 736 1003
rect 730 998 736 999
rect 802 1003 808 1004
rect 802 999 803 1003
rect 807 999 808 1003
rect 802 998 808 999
rect 866 1003 872 1004
rect 866 999 867 1003
rect 871 999 872 1003
rect 866 998 872 999
rect 926 1003 932 1004
rect 926 999 927 1003
rect 931 999 932 1003
rect 926 998 932 999
rect 994 1003 1000 1004
rect 994 999 995 1003
rect 999 999 1000 1003
rect 994 998 1000 999
rect 1054 1003 1060 1004
rect 1094 1003 1100 1004
rect 1054 999 1055 1003
rect 1059 999 1060 1003
rect 1136 1001 1138 1021
rect 1160 1009 1162 1021
rect 1176 1020 1178 1054
rect 1238 1051 1239 1055
rect 1243 1051 1244 1055
rect 1238 1050 1244 1051
rect 1350 1055 1356 1056
rect 1350 1051 1351 1055
rect 1355 1051 1356 1055
rect 1350 1050 1356 1051
rect 1566 1055 1572 1056
rect 1566 1051 1567 1055
rect 1571 1051 1572 1055
rect 1566 1050 1572 1051
rect 1598 1055 1604 1056
rect 1598 1051 1599 1055
rect 1603 1051 1604 1055
rect 1598 1050 1604 1051
rect 1240 1032 1242 1050
rect 1246 1044 1252 1045
rect 1246 1040 1247 1044
rect 1251 1040 1252 1044
rect 1246 1039 1252 1040
rect 1238 1031 1244 1032
rect 1238 1027 1239 1031
rect 1243 1027 1244 1031
rect 1248 1027 1250 1039
rect 1352 1032 1354 1050
rect 1358 1044 1364 1045
rect 1358 1040 1359 1044
rect 1363 1040 1364 1044
rect 1358 1039 1364 1040
rect 1470 1044 1476 1045
rect 1470 1040 1471 1044
rect 1475 1040 1476 1044
rect 1470 1039 1476 1040
rect 1350 1031 1356 1032
rect 1350 1027 1351 1031
rect 1355 1027 1356 1031
rect 1360 1027 1362 1039
rect 1472 1027 1474 1039
rect 1568 1032 1570 1050
rect 1574 1044 1580 1045
rect 1574 1040 1575 1044
rect 1579 1040 1580 1044
rect 1574 1039 1580 1040
rect 1670 1044 1676 1045
rect 1670 1040 1671 1044
rect 1675 1040 1676 1044
rect 1670 1039 1676 1040
rect 1486 1031 1492 1032
rect 1486 1027 1487 1031
rect 1491 1027 1492 1031
rect 1566 1031 1572 1032
rect 1566 1027 1567 1031
rect 1571 1027 1572 1031
rect 1576 1027 1578 1039
rect 1672 1027 1674 1039
rect 1704 1032 1706 1058
rect 1750 1055 1756 1056
rect 1750 1051 1751 1055
rect 1755 1051 1756 1055
rect 1750 1050 1756 1051
rect 1814 1055 1820 1056
rect 1814 1051 1815 1055
rect 1819 1051 1820 1055
rect 1814 1050 1820 1051
rect 1752 1032 1754 1050
rect 1758 1044 1764 1045
rect 1758 1040 1759 1044
rect 1763 1040 1764 1044
rect 1758 1039 1764 1040
rect 1702 1031 1708 1032
rect 1702 1027 1703 1031
rect 1707 1027 1708 1031
rect 1231 1026 1235 1027
rect 1238 1026 1244 1027
rect 1247 1026 1251 1027
rect 1231 1021 1235 1022
rect 1247 1021 1251 1022
rect 1303 1026 1307 1027
rect 1350 1026 1356 1027
rect 1359 1026 1363 1027
rect 1303 1021 1307 1022
rect 1359 1021 1363 1022
rect 1383 1026 1387 1027
rect 1383 1021 1387 1022
rect 1463 1026 1467 1027
rect 1463 1021 1467 1022
rect 1471 1026 1475 1027
rect 1486 1026 1492 1027
rect 1543 1026 1547 1027
rect 1566 1026 1572 1027
rect 1575 1026 1579 1027
rect 1471 1021 1475 1022
rect 1174 1019 1180 1020
rect 1174 1015 1175 1019
rect 1179 1015 1180 1019
rect 1174 1014 1180 1015
rect 1186 1019 1192 1020
rect 1186 1015 1187 1019
rect 1191 1015 1192 1019
rect 1186 1014 1192 1015
rect 1158 1008 1164 1009
rect 1158 1004 1159 1008
rect 1163 1004 1164 1008
rect 1158 1003 1164 1004
rect 1054 998 1060 999
rect 1134 1000 1140 1001
rect 774 988 780 989
rect 774 984 775 988
rect 779 984 780 988
rect 774 983 780 984
rect 838 988 844 989
rect 838 984 839 988
rect 843 984 844 988
rect 838 983 844 984
rect 902 988 908 989
rect 902 984 903 988
rect 907 984 908 988
rect 902 983 908 984
rect 966 988 972 989
rect 966 984 967 988
rect 971 984 972 988
rect 966 983 972 984
rect 1038 988 1044 989
rect 1038 984 1039 988
rect 1043 984 1044 988
rect 1038 983 1044 984
rect 776 979 778 983
rect 840 979 842 983
rect 904 979 906 983
rect 968 979 970 983
rect 1040 979 1042 983
rect 735 978 739 979
rect 735 973 739 974
rect 775 978 779 979
rect 775 973 779 974
rect 799 978 803 979
rect 799 973 803 974
rect 839 978 843 979
rect 839 973 843 974
rect 863 978 867 979
rect 863 973 867 974
rect 903 978 907 979
rect 903 973 907 974
rect 927 978 931 979
rect 927 973 931 974
rect 967 978 971 979
rect 967 973 971 974
rect 991 978 995 979
rect 991 973 995 974
rect 1039 978 1043 979
rect 1039 973 1043 974
rect 1047 978 1051 979
rect 1047 973 1051 974
rect 734 972 740 973
rect 734 968 735 972
rect 739 968 740 972
rect 734 967 740 968
rect 798 972 804 973
rect 798 968 799 972
rect 803 968 804 972
rect 798 967 804 968
rect 862 972 868 973
rect 862 968 863 972
rect 867 968 868 972
rect 862 967 868 968
rect 926 972 932 973
rect 926 968 927 972
rect 931 968 932 972
rect 926 967 932 968
rect 990 972 996 973
rect 990 968 991 972
rect 995 968 996 972
rect 990 967 996 968
rect 1046 972 1052 973
rect 1046 968 1047 972
rect 1051 968 1052 972
rect 1046 967 1052 968
rect 710 963 716 964
rect 710 959 711 963
rect 715 959 716 963
rect 710 958 716 959
rect 662 955 668 956
rect 662 951 663 955
rect 667 951 668 955
rect 662 950 668 951
rect 726 955 732 956
rect 726 951 727 955
rect 731 951 732 955
rect 726 950 732 951
rect 790 955 796 956
rect 790 951 791 955
rect 795 951 796 955
rect 790 950 796 951
rect 854 955 860 956
rect 854 951 855 955
rect 859 951 860 955
rect 854 950 860 951
rect 918 955 924 956
rect 918 951 919 955
rect 923 951 924 955
rect 918 950 924 951
rect 998 955 1004 956
rect 998 951 999 955
rect 1003 951 1004 955
rect 998 950 1004 951
rect 1026 955 1032 956
rect 1026 951 1027 955
rect 1031 951 1032 955
rect 1026 950 1032 951
rect 526 944 532 945
rect 526 940 527 944
rect 531 940 532 944
rect 526 939 532 940
rect 598 944 604 945
rect 598 940 599 944
rect 603 940 604 944
rect 598 939 604 940
rect 482 931 488 932
rect 482 927 483 931
rect 487 927 488 931
rect 482 926 488 927
rect 518 931 524 932
rect 518 927 519 931
rect 523 927 524 931
rect 528 927 530 939
rect 600 927 602 939
rect 664 932 666 950
rect 670 944 676 945
rect 670 940 671 944
rect 675 940 676 944
rect 670 939 676 940
rect 654 931 660 932
rect 654 927 655 931
rect 659 927 660 931
rect 518 926 524 927
rect 527 926 531 927
rect 527 921 531 922
rect 599 926 603 927
rect 654 926 660 927
rect 662 931 668 932
rect 662 927 663 931
rect 667 927 668 931
rect 672 927 674 939
rect 728 932 730 950
rect 734 944 740 945
rect 734 940 735 944
rect 739 940 740 944
rect 734 939 740 940
rect 726 931 732 932
rect 726 927 727 931
rect 731 927 732 931
rect 736 927 738 939
rect 792 932 794 950
rect 798 944 804 945
rect 798 940 799 944
rect 803 940 804 944
rect 798 939 804 940
rect 790 931 796 932
rect 790 927 791 931
rect 795 927 796 931
rect 800 927 802 939
rect 856 932 858 950
rect 862 944 868 945
rect 862 940 863 944
rect 867 940 868 944
rect 862 939 868 940
rect 854 931 860 932
rect 854 927 855 931
rect 859 927 860 931
rect 864 927 866 939
rect 920 932 922 950
rect 926 944 932 945
rect 926 940 927 944
rect 931 940 932 944
rect 926 939 932 940
rect 990 944 996 945
rect 990 940 991 944
rect 995 940 996 944
rect 990 939 996 940
rect 918 931 924 932
rect 918 927 919 931
rect 923 927 924 931
rect 928 927 930 939
rect 992 927 994 939
rect 662 926 668 927
rect 671 926 675 927
rect 726 926 732 927
rect 735 926 739 927
rect 599 921 603 922
rect 470 919 476 920
rect 470 915 471 919
rect 475 915 476 919
rect 470 914 476 915
rect 528 909 530 921
rect 546 919 552 920
rect 546 915 547 919
rect 551 915 552 919
rect 546 914 552 915
rect 554 919 560 920
rect 554 915 555 919
rect 559 915 560 919
rect 554 914 560 915
rect 398 908 404 909
rect 398 904 399 908
rect 403 904 404 908
rect 398 903 404 904
rect 462 908 468 909
rect 462 904 463 908
rect 467 904 468 908
rect 462 903 468 904
rect 526 908 532 909
rect 526 904 527 908
rect 531 904 532 908
rect 526 903 532 904
rect 350 895 356 896
rect 350 891 351 895
rect 355 891 356 895
rect 350 890 356 891
rect 386 895 392 896
rect 386 891 387 895
rect 391 891 392 895
rect 386 890 392 891
rect 326 880 332 881
rect 326 876 327 880
rect 331 876 332 880
rect 326 875 332 876
rect 328 871 330 875
rect 327 870 331 871
rect 327 865 331 866
rect 343 870 347 871
rect 343 865 347 866
rect 342 864 348 865
rect 342 860 343 864
rect 347 860 348 864
rect 342 859 348 860
rect 162 847 168 848
rect 110 844 116 845
rect 110 840 111 844
rect 115 840 116 844
rect 162 843 163 847
rect 167 843 168 847
rect 162 842 168 843
rect 202 847 208 848
rect 202 843 203 847
rect 207 843 208 847
rect 202 842 208 843
rect 270 847 276 848
rect 270 843 271 847
rect 275 843 276 847
rect 270 842 276 843
rect 302 847 308 848
rect 302 843 303 847
rect 307 843 308 847
rect 302 842 308 843
rect 110 839 116 840
rect 112 819 114 839
rect 134 836 140 837
rect 134 832 135 836
rect 139 832 140 836
rect 134 831 140 832
rect 136 819 138 831
rect 164 824 166 842
rect 174 836 180 837
rect 174 832 175 836
rect 179 832 180 836
rect 174 831 180 832
rect 154 823 160 824
rect 154 819 155 823
rect 159 819 160 823
rect 111 818 115 819
rect 111 813 115 814
rect 135 818 139 819
rect 154 818 160 819
rect 162 823 168 824
rect 162 819 163 823
rect 167 819 168 823
rect 176 819 178 831
rect 204 824 206 842
rect 214 836 220 837
rect 214 832 215 836
rect 219 832 220 836
rect 214 831 220 832
rect 202 823 208 824
rect 202 819 203 823
rect 207 819 208 823
rect 216 819 218 831
rect 272 824 274 842
rect 278 836 284 837
rect 278 832 279 836
rect 283 832 284 836
rect 278 831 284 832
rect 342 836 348 837
rect 342 832 343 836
rect 347 832 348 836
rect 342 831 348 832
rect 270 823 276 824
rect 270 819 271 823
rect 275 819 276 823
rect 280 819 282 831
rect 344 819 346 831
rect 352 824 354 890
rect 398 880 404 881
rect 398 876 399 880
rect 403 876 404 880
rect 398 875 404 876
rect 462 880 468 881
rect 462 876 463 880
rect 467 876 468 880
rect 462 875 468 876
rect 526 880 532 881
rect 526 876 527 880
rect 531 876 532 880
rect 526 875 532 876
rect 400 871 402 875
rect 464 871 466 875
rect 528 871 530 875
rect 399 870 403 871
rect 399 865 403 866
rect 463 870 467 871
rect 463 865 467 866
rect 527 870 531 871
rect 527 865 531 866
rect 535 870 539 871
rect 535 865 539 866
rect 398 864 404 865
rect 398 860 399 864
rect 403 860 404 864
rect 398 859 404 860
rect 462 864 468 865
rect 462 860 463 864
rect 467 860 468 864
rect 462 859 468 860
rect 534 864 540 865
rect 534 860 535 864
rect 539 860 540 864
rect 534 859 540 860
rect 548 853 550 914
rect 556 896 558 914
rect 600 909 602 921
rect 626 919 632 920
rect 626 915 627 919
rect 631 915 632 919
rect 626 914 632 915
rect 598 908 604 909
rect 598 904 599 908
rect 603 904 604 908
rect 598 903 604 904
rect 628 896 630 914
rect 554 895 560 896
rect 554 891 555 895
rect 559 891 560 895
rect 554 890 560 891
rect 626 895 632 896
rect 626 891 627 895
rect 631 891 632 895
rect 626 890 632 891
rect 598 880 604 881
rect 598 876 599 880
rect 603 876 604 880
rect 598 875 604 876
rect 600 871 602 875
rect 656 872 658 926
rect 671 921 675 922
rect 735 921 739 922
rect 743 926 747 927
rect 790 926 796 927
rect 799 926 803 927
rect 743 921 747 922
rect 799 921 803 922
rect 815 926 819 927
rect 854 926 860 927
rect 863 926 867 927
rect 815 921 819 922
rect 863 921 867 922
rect 895 926 899 927
rect 918 926 924 927
rect 927 926 931 927
rect 895 921 899 922
rect 927 921 931 922
rect 983 926 987 927
rect 983 921 987 922
rect 991 926 995 927
rect 991 921 995 922
rect 672 909 674 921
rect 698 919 704 920
rect 698 915 699 919
rect 703 915 704 919
rect 698 914 704 915
rect 670 908 676 909
rect 670 904 671 908
rect 675 904 676 908
rect 670 903 676 904
rect 700 896 702 914
rect 744 909 746 921
rect 770 919 776 920
rect 770 915 771 919
rect 775 915 776 919
rect 770 914 776 915
rect 742 908 748 909
rect 742 904 743 908
rect 747 904 748 908
rect 742 903 748 904
rect 772 896 774 914
rect 816 909 818 921
rect 842 919 848 920
rect 842 915 843 919
rect 847 915 848 919
rect 842 914 848 915
rect 814 908 820 909
rect 814 904 815 908
rect 819 904 820 908
rect 814 903 820 904
rect 844 896 846 914
rect 896 909 898 921
rect 984 909 986 921
rect 1000 920 1002 950
rect 1028 932 1030 950
rect 1046 944 1052 945
rect 1046 940 1047 944
rect 1051 940 1052 944
rect 1046 939 1052 940
rect 1026 931 1032 932
rect 1026 927 1027 931
rect 1031 927 1032 931
rect 1048 927 1050 939
rect 1056 932 1058 998
rect 1134 996 1135 1000
rect 1139 996 1140 1000
rect 1188 996 1190 1014
rect 1232 1009 1234 1021
rect 1258 1019 1264 1020
rect 1258 1015 1259 1019
rect 1263 1015 1264 1019
rect 1258 1014 1264 1015
rect 1230 1008 1236 1009
rect 1230 1004 1231 1008
rect 1235 1004 1236 1008
rect 1230 1003 1236 1004
rect 1260 996 1262 1014
rect 1304 1009 1306 1021
rect 1330 1019 1336 1020
rect 1330 1015 1331 1019
rect 1335 1015 1336 1019
rect 1330 1014 1336 1015
rect 1302 1008 1308 1009
rect 1302 1004 1303 1008
rect 1307 1004 1308 1008
rect 1302 1003 1308 1004
rect 1332 996 1334 1014
rect 1384 1009 1386 1021
rect 1464 1009 1466 1021
rect 1382 1008 1388 1009
rect 1382 1004 1383 1008
rect 1387 1004 1388 1008
rect 1382 1003 1388 1004
rect 1462 1008 1468 1009
rect 1462 1004 1463 1008
rect 1467 1004 1468 1008
rect 1462 1003 1468 1004
rect 1488 996 1490 1026
rect 1543 1021 1547 1022
rect 1575 1021 1579 1022
rect 1623 1026 1627 1027
rect 1623 1021 1627 1022
rect 1671 1026 1675 1027
rect 1671 1021 1675 1022
rect 1695 1026 1699 1027
rect 1702 1026 1708 1027
rect 1750 1031 1756 1032
rect 1750 1027 1751 1031
rect 1755 1027 1756 1031
rect 1760 1027 1762 1039
rect 1750 1026 1756 1027
rect 1759 1026 1763 1027
rect 1695 1021 1699 1022
rect 1759 1021 1763 1022
rect 1526 1019 1532 1020
rect 1526 1015 1527 1019
rect 1531 1015 1532 1019
rect 1526 1014 1532 1015
rect 1534 1019 1540 1020
rect 1534 1015 1535 1019
rect 1539 1015 1540 1019
rect 1534 1014 1540 1015
rect 1528 996 1530 1014
rect 1134 995 1140 996
rect 1186 995 1192 996
rect 1094 991 1100 992
rect 1094 987 1095 991
rect 1099 987 1100 991
rect 1186 991 1187 995
rect 1191 991 1192 995
rect 1186 990 1192 991
rect 1258 995 1264 996
rect 1258 991 1259 995
rect 1263 991 1264 995
rect 1258 990 1264 991
rect 1330 995 1336 996
rect 1330 991 1331 995
rect 1335 991 1336 995
rect 1330 990 1336 991
rect 1338 995 1344 996
rect 1338 991 1339 995
rect 1343 991 1344 995
rect 1338 990 1344 991
rect 1486 995 1492 996
rect 1486 991 1487 995
rect 1491 991 1492 995
rect 1486 990 1492 991
rect 1526 995 1532 996
rect 1526 991 1527 995
rect 1531 991 1532 995
rect 1526 990 1532 991
rect 1094 986 1100 987
rect 1096 979 1098 986
rect 1134 983 1140 984
rect 1134 979 1135 983
rect 1139 979 1140 983
rect 1095 978 1099 979
rect 1134 978 1140 979
rect 1158 980 1164 981
rect 1136 975 1138 978
rect 1158 976 1159 980
rect 1163 976 1164 980
rect 1158 975 1164 976
rect 1230 980 1236 981
rect 1230 976 1231 980
rect 1235 976 1236 980
rect 1230 975 1236 976
rect 1302 980 1308 981
rect 1302 976 1303 980
rect 1307 976 1308 980
rect 1302 975 1308 976
rect 1095 973 1099 974
rect 1135 974 1139 975
rect 1096 970 1098 973
rect 1094 969 1100 970
rect 1135 969 1139 970
rect 1159 974 1163 975
rect 1159 969 1163 970
rect 1231 974 1235 975
rect 1231 969 1235 970
rect 1239 974 1243 975
rect 1239 969 1243 970
rect 1303 974 1307 975
rect 1303 969 1307 970
rect 1094 965 1095 969
rect 1099 965 1100 969
rect 1136 966 1138 969
rect 1238 968 1244 969
rect 1094 964 1100 965
rect 1134 965 1140 966
rect 1134 961 1135 965
rect 1139 961 1140 965
rect 1238 964 1239 968
rect 1243 964 1244 968
rect 1238 963 1244 964
rect 1302 968 1308 969
rect 1302 964 1303 968
rect 1307 964 1308 968
rect 1302 963 1308 964
rect 1134 960 1140 961
rect 1094 952 1100 953
rect 1094 948 1095 952
rect 1099 948 1100 952
rect 1294 951 1300 952
rect 1094 947 1100 948
rect 1134 948 1140 949
rect 1054 931 1060 932
rect 1054 927 1055 931
rect 1059 927 1060 931
rect 1096 927 1098 947
rect 1134 944 1135 948
rect 1139 944 1140 948
rect 1294 947 1295 951
rect 1299 947 1300 951
rect 1294 946 1300 947
rect 1134 943 1140 944
rect 1026 926 1032 927
rect 1047 926 1051 927
rect 1054 926 1060 927
rect 1095 926 1099 927
rect 1047 921 1051 922
rect 1095 921 1099 922
rect 998 919 1004 920
rect 998 915 999 919
rect 1003 915 1004 919
rect 998 914 1004 915
rect 1026 919 1032 920
rect 1026 915 1027 919
rect 1031 915 1032 919
rect 1026 914 1032 915
rect 894 908 900 909
rect 894 904 895 908
rect 899 904 900 908
rect 894 903 900 904
rect 982 908 988 909
rect 982 904 983 908
rect 987 904 988 908
rect 982 903 988 904
rect 1028 896 1030 914
rect 1048 909 1050 921
rect 1046 908 1052 909
rect 1046 904 1047 908
rect 1051 904 1052 908
rect 1046 903 1052 904
rect 1096 901 1098 921
rect 1136 919 1138 943
rect 1238 940 1244 941
rect 1238 936 1239 940
rect 1243 936 1244 940
rect 1238 935 1244 936
rect 1240 919 1242 935
rect 1296 928 1298 946
rect 1302 940 1308 941
rect 1302 936 1303 940
rect 1307 936 1308 940
rect 1302 935 1308 936
rect 1294 927 1300 928
rect 1294 923 1295 927
rect 1299 923 1300 927
rect 1294 922 1300 923
rect 1304 919 1306 935
rect 1340 920 1342 990
rect 1382 980 1388 981
rect 1382 976 1383 980
rect 1387 976 1388 980
rect 1382 975 1388 976
rect 1462 980 1468 981
rect 1462 976 1463 980
rect 1467 976 1468 980
rect 1462 975 1468 976
rect 1375 974 1379 975
rect 1375 969 1379 970
rect 1383 974 1387 975
rect 1383 969 1387 970
rect 1439 974 1443 975
rect 1439 969 1443 970
rect 1463 974 1467 975
rect 1463 969 1467 970
rect 1511 974 1515 975
rect 1511 969 1515 970
rect 1374 968 1380 969
rect 1374 964 1375 968
rect 1379 964 1380 968
rect 1374 963 1380 964
rect 1438 968 1444 969
rect 1438 964 1439 968
rect 1443 964 1444 968
rect 1438 963 1444 964
rect 1510 968 1516 969
rect 1510 964 1511 968
rect 1515 964 1516 968
rect 1510 963 1516 964
rect 1536 952 1538 1014
rect 1544 1009 1546 1021
rect 1624 1009 1626 1021
rect 1650 1019 1656 1020
rect 1650 1015 1651 1019
rect 1655 1015 1656 1019
rect 1650 1014 1656 1015
rect 1542 1008 1548 1009
rect 1542 1004 1543 1008
rect 1547 1004 1548 1008
rect 1542 1003 1548 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1652 996 1654 1014
rect 1696 1009 1698 1021
rect 1722 1019 1728 1020
rect 1722 1015 1723 1019
rect 1727 1015 1728 1019
rect 1722 1014 1728 1015
rect 1694 1008 1700 1009
rect 1694 1004 1695 1008
rect 1699 1004 1700 1008
rect 1694 1003 1700 1004
rect 1724 996 1726 1014
rect 1760 1009 1762 1021
rect 1816 1020 1818 1050
rect 1846 1044 1852 1045
rect 1846 1040 1847 1044
rect 1851 1040 1852 1044
rect 1846 1039 1852 1040
rect 1926 1044 1932 1045
rect 1926 1040 1927 1044
rect 1931 1040 1932 1044
rect 1926 1039 1932 1040
rect 1848 1027 1850 1039
rect 1928 1027 1930 1039
rect 2000 1032 2002 1094
rect 2030 1084 2036 1085
rect 2030 1080 2031 1084
rect 2035 1080 2036 1084
rect 2030 1079 2036 1080
rect 2007 1078 2011 1079
rect 2007 1073 2011 1074
rect 2031 1078 2035 1079
rect 2031 1073 2035 1074
rect 2006 1072 2012 1073
rect 2006 1068 2007 1072
rect 2011 1068 2012 1072
rect 2006 1067 2012 1068
rect 2048 1056 2050 1118
rect 2056 1100 2058 1138
rect 2072 1131 2074 1151
rect 2071 1130 2075 1131
rect 2071 1125 2075 1126
rect 2072 1113 2074 1125
rect 2080 1124 2082 1162
rect 2088 1144 2090 1206
rect 2118 1199 2124 1200
rect 2118 1195 2119 1199
rect 2123 1195 2124 1199
rect 2118 1194 2124 1195
rect 2120 1191 2122 1194
rect 2119 1190 2123 1191
rect 2119 1185 2123 1186
rect 2120 1182 2122 1185
rect 2118 1181 2124 1182
rect 2118 1177 2119 1181
rect 2123 1177 2124 1181
rect 2118 1176 2124 1177
rect 2118 1164 2124 1165
rect 2118 1160 2119 1164
rect 2123 1160 2124 1164
rect 2118 1159 2124 1160
rect 2086 1143 2092 1144
rect 2086 1139 2087 1143
rect 2091 1139 2092 1143
rect 2086 1138 2092 1139
rect 2120 1131 2122 1159
rect 2119 1130 2123 1131
rect 2119 1125 2123 1126
rect 2078 1123 2084 1124
rect 2078 1119 2079 1123
rect 2083 1119 2084 1123
rect 2078 1118 2084 1119
rect 2070 1112 2076 1113
rect 2070 1108 2071 1112
rect 2075 1108 2076 1112
rect 2070 1107 2076 1108
rect 2120 1105 2122 1125
rect 2118 1104 2124 1105
rect 2118 1100 2119 1104
rect 2123 1100 2124 1104
rect 2054 1099 2060 1100
rect 2054 1095 2055 1099
rect 2059 1095 2060 1099
rect 2054 1094 2060 1095
rect 2078 1099 2084 1100
rect 2118 1099 2124 1100
rect 2078 1095 2079 1099
rect 2083 1095 2084 1099
rect 2078 1094 2084 1095
rect 2070 1084 2076 1085
rect 2070 1080 2071 1084
rect 2075 1080 2076 1084
rect 2070 1079 2076 1080
rect 2071 1078 2075 1079
rect 2071 1073 2075 1074
rect 2070 1072 2076 1073
rect 2070 1068 2071 1072
rect 2075 1068 2076 1072
rect 2070 1067 2076 1068
rect 2046 1055 2052 1056
rect 2046 1051 2047 1055
rect 2051 1051 2052 1055
rect 2046 1050 2052 1051
rect 2006 1044 2012 1045
rect 2006 1040 2007 1044
rect 2011 1040 2012 1044
rect 2006 1039 2012 1040
rect 2070 1044 2076 1045
rect 2070 1040 2071 1044
rect 2075 1040 2076 1044
rect 2070 1039 2076 1040
rect 1998 1031 2004 1032
rect 1998 1027 1999 1031
rect 2003 1027 2004 1031
rect 2008 1027 2010 1039
rect 2072 1027 2074 1039
rect 2080 1032 2082 1094
rect 2118 1087 2124 1088
rect 2118 1083 2119 1087
rect 2123 1083 2124 1087
rect 2118 1082 2124 1083
rect 2120 1079 2122 1082
rect 2119 1078 2123 1079
rect 2119 1073 2123 1074
rect 2120 1070 2122 1073
rect 2118 1069 2124 1070
rect 2118 1065 2119 1069
rect 2123 1065 2124 1069
rect 2118 1064 2124 1065
rect 2118 1052 2124 1053
rect 2118 1048 2119 1052
rect 2123 1048 2124 1052
rect 2118 1047 2124 1048
rect 2078 1031 2084 1032
rect 2078 1027 2079 1031
rect 2083 1027 2084 1031
rect 2120 1027 2122 1047
rect 1823 1026 1827 1027
rect 1823 1021 1827 1022
rect 1847 1026 1851 1027
rect 1847 1021 1851 1022
rect 1887 1026 1891 1027
rect 1887 1021 1891 1022
rect 1927 1026 1931 1027
rect 1927 1021 1931 1022
rect 1951 1026 1955 1027
rect 1998 1026 2004 1027
rect 2007 1026 2011 1027
rect 1951 1021 1955 1022
rect 2007 1021 2011 1022
rect 2071 1026 2075 1027
rect 2078 1026 2084 1027
rect 2119 1026 2123 1027
rect 2071 1021 2075 1022
rect 2119 1021 2123 1022
rect 1814 1019 1820 1020
rect 1814 1015 1815 1019
rect 1819 1015 1820 1019
rect 1814 1014 1820 1015
rect 1824 1009 1826 1021
rect 1866 1019 1872 1020
rect 1866 1015 1867 1019
rect 1871 1015 1872 1019
rect 1866 1014 1872 1015
rect 1758 1008 1764 1009
rect 1758 1004 1759 1008
rect 1763 1004 1764 1008
rect 1758 1003 1764 1004
rect 1822 1008 1828 1009
rect 1822 1004 1823 1008
rect 1827 1004 1828 1008
rect 1822 1003 1828 1004
rect 1868 1000 1870 1014
rect 1888 1009 1890 1021
rect 1914 1019 1920 1020
rect 1914 1015 1915 1019
rect 1919 1015 1920 1019
rect 1914 1014 1920 1015
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1866 999 1872 1000
rect 1650 995 1656 996
rect 1650 991 1651 995
rect 1655 991 1656 995
rect 1650 990 1656 991
rect 1722 995 1728 996
rect 1722 991 1723 995
rect 1727 991 1728 995
rect 1722 990 1728 991
rect 1786 995 1792 996
rect 1786 991 1787 995
rect 1791 991 1792 995
rect 1866 995 1867 999
rect 1871 995 1872 999
rect 1916 996 1918 1014
rect 1952 1009 1954 1021
rect 1950 1008 1956 1009
rect 1950 1004 1951 1008
rect 1955 1004 1956 1008
rect 1950 1003 1956 1004
rect 2120 1001 2122 1021
rect 2118 1000 2124 1001
rect 2118 996 2119 1000
rect 2123 996 2124 1000
rect 1866 994 1872 995
rect 1914 995 1920 996
rect 2118 995 2124 996
rect 1786 990 1792 991
rect 1914 991 1915 995
rect 1919 991 1920 995
rect 1914 990 1920 991
rect 1542 980 1548 981
rect 1542 976 1543 980
rect 1547 976 1548 980
rect 1542 975 1548 976
rect 1622 980 1628 981
rect 1622 976 1623 980
rect 1627 976 1628 980
rect 1622 975 1628 976
rect 1694 980 1700 981
rect 1694 976 1695 980
rect 1699 976 1700 980
rect 1694 975 1700 976
rect 1758 980 1764 981
rect 1758 976 1759 980
rect 1763 976 1764 980
rect 1758 975 1764 976
rect 1543 974 1547 975
rect 1543 969 1547 970
rect 1583 974 1587 975
rect 1583 969 1587 970
rect 1623 974 1627 975
rect 1623 969 1627 970
rect 1655 974 1659 975
rect 1655 969 1659 970
rect 1695 974 1699 975
rect 1695 969 1699 970
rect 1727 974 1731 975
rect 1727 969 1731 970
rect 1759 974 1763 975
rect 1759 969 1763 970
rect 1582 968 1588 969
rect 1582 964 1583 968
rect 1587 964 1588 968
rect 1582 963 1588 964
rect 1654 968 1660 969
rect 1654 964 1655 968
rect 1659 964 1660 968
rect 1654 963 1660 964
rect 1726 968 1732 969
rect 1726 964 1727 968
rect 1731 964 1732 968
rect 1726 963 1732 964
rect 1610 959 1616 960
rect 1610 955 1611 959
rect 1615 955 1616 959
rect 1610 954 1616 955
rect 1366 951 1372 952
rect 1366 947 1367 951
rect 1371 947 1372 951
rect 1366 946 1372 947
rect 1382 951 1388 952
rect 1382 947 1383 951
rect 1387 947 1388 951
rect 1382 946 1388 947
rect 1502 951 1508 952
rect 1502 947 1503 951
rect 1507 947 1508 951
rect 1502 946 1508 947
rect 1534 951 1540 952
rect 1534 947 1535 951
rect 1539 947 1540 951
rect 1534 946 1540 947
rect 1368 928 1370 946
rect 1374 940 1380 941
rect 1374 936 1375 940
rect 1379 936 1380 940
rect 1374 935 1380 936
rect 1366 927 1372 928
rect 1366 923 1367 927
rect 1371 923 1372 927
rect 1366 922 1372 923
rect 1338 919 1344 920
rect 1376 919 1378 935
rect 1135 918 1139 919
rect 1135 913 1139 914
rect 1239 918 1243 919
rect 1239 913 1243 914
rect 1287 918 1291 919
rect 1287 913 1291 914
rect 1303 918 1307 919
rect 1303 913 1307 914
rect 1327 918 1331 919
rect 1338 915 1339 919
rect 1343 915 1344 919
rect 1338 914 1344 915
rect 1375 918 1379 919
rect 1327 913 1331 914
rect 1375 913 1379 914
rect 1094 900 1100 901
rect 1094 896 1095 900
rect 1099 896 1100 900
rect 698 895 704 896
rect 698 891 699 895
rect 703 891 704 895
rect 698 890 704 891
rect 770 895 776 896
rect 770 891 771 895
rect 775 891 776 895
rect 770 890 776 891
rect 842 895 848 896
rect 842 891 843 895
rect 847 891 848 895
rect 842 890 848 891
rect 918 895 924 896
rect 918 891 919 895
rect 923 891 924 895
rect 918 890 924 891
rect 1026 895 1032 896
rect 1026 891 1027 895
rect 1031 891 1032 895
rect 1026 890 1032 891
rect 1086 895 1092 896
rect 1094 895 1100 896
rect 1086 891 1087 895
rect 1091 891 1092 895
rect 1136 893 1138 913
rect 1288 901 1290 913
rect 1328 901 1330 913
rect 1362 911 1368 912
rect 1362 907 1363 911
rect 1367 907 1368 911
rect 1362 906 1368 907
rect 1286 900 1292 901
rect 1286 896 1287 900
rect 1291 896 1292 900
rect 1286 895 1292 896
rect 1326 900 1332 901
rect 1326 896 1327 900
rect 1331 896 1332 900
rect 1326 895 1332 896
rect 1086 890 1092 891
rect 1134 892 1140 893
rect 670 880 676 881
rect 670 876 671 880
rect 675 876 676 880
rect 670 875 676 876
rect 742 880 748 881
rect 742 876 743 880
rect 747 876 748 880
rect 742 875 748 876
rect 814 880 820 881
rect 814 876 815 880
rect 819 876 820 880
rect 814 875 820 876
rect 894 880 900 881
rect 894 876 895 880
rect 899 876 900 880
rect 894 875 900 876
rect 654 871 660 872
rect 672 871 674 875
rect 744 871 746 875
rect 816 871 818 875
rect 896 871 898 875
rect 920 872 922 890
rect 982 880 988 881
rect 982 876 983 880
rect 987 876 988 880
rect 982 875 988 876
rect 1046 880 1052 881
rect 1046 876 1047 880
rect 1051 876 1052 880
rect 1046 875 1052 876
rect 918 871 924 872
rect 984 871 986 875
rect 1048 871 1050 875
rect 599 870 603 871
rect 599 865 603 866
rect 615 870 619 871
rect 654 867 655 871
rect 659 867 660 871
rect 654 866 660 867
rect 671 870 675 871
rect 615 865 619 866
rect 671 865 675 866
rect 711 870 715 871
rect 711 865 715 866
rect 743 870 747 871
rect 743 865 747 866
rect 815 870 819 871
rect 815 865 819 866
rect 823 870 827 871
rect 823 865 827 866
rect 895 870 899 871
rect 918 867 919 871
rect 923 867 924 871
rect 918 866 924 867
rect 943 870 947 871
rect 895 865 899 866
rect 943 865 947 866
rect 983 870 987 871
rect 983 865 987 866
rect 1047 870 1051 871
rect 1047 865 1051 866
rect 614 864 620 865
rect 614 860 615 864
rect 619 860 620 864
rect 614 859 620 860
rect 710 864 716 865
rect 710 860 711 864
rect 715 860 716 864
rect 710 859 716 860
rect 822 864 828 865
rect 822 860 823 864
rect 827 860 828 864
rect 822 859 828 860
rect 942 864 948 865
rect 942 860 943 864
rect 947 860 948 864
rect 942 859 948 860
rect 1046 864 1052 865
rect 1046 860 1047 864
rect 1051 860 1052 864
rect 1046 859 1052 860
rect 902 855 908 856
rect 547 852 551 853
rect 847 852 851 853
rect 902 851 903 855
rect 907 851 908 855
rect 902 850 908 851
rect 406 847 412 848
rect 406 843 407 847
rect 411 843 412 847
rect 406 842 412 843
rect 470 847 476 848
rect 547 847 551 848
rect 606 847 612 848
rect 470 843 471 847
rect 475 843 476 847
rect 470 842 476 843
rect 606 843 607 847
rect 611 843 612 847
rect 606 842 612 843
rect 702 847 708 848
rect 702 843 703 847
rect 707 843 708 847
rect 702 842 708 843
rect 846 847 852 848
rect 846 843 847 847
rect 851 843 852 847
rect 846 842 852 843
rect 858 847 864 848
rect 858 843 859 847
rect 863 843 864 847
rect 858 842 864 843
rect 398 836 404 837
rect 398 832 399 836
rect 403 832 404 836
rect 398 831 404 832
rect 350 823 356 824
rect 350 819 351 823
rect 355 819 356 823
rect 400 819 402 831
rect 162 818 168 819
rect 175 818 179 819
rect 202 818 208 819
rect 215 818 219 819
rect 270 818 276 819
rect 279 818 283 819
rect 135 813 139 814
rect 112 793 114 813
rect 136 801 138 813
rect 134 800 140 801
rect 134 796 135 800
rect 139 796 140 800
rect 134 795 140 796
rect 110 792 116 793
rect 110 788 111 792
rect 115 788 116 792
rect 156 788 158 818
rect 175 813 179 814
rect 215 813 219 814
rect 279 813 283 814
rect 335 818 339 819
rect 335 813 339 814
rect 343 818 347 819
rect 350 818 356 819
rect 391 818 395 819
rect 343 813 347 814
rect 391 813 395 814
rect 399 818 403 819
rect 399 813 403 814
rect 162 811 168 812
rect 162 807 163 811
rect 167 807 168 811
rect 162 806 168 807
rect 110 787 116 788
rect 154 787 160 788
rect 154 783 155 787
rect 159 783 160 787
rect 154 782 160 783
rect 110 775 116 776
rect 110 771 111 775
rect 115 771 116 775
rect 110 770 116 771
rect 134 772 140 773
rect 112 767 114 770
rect 134 768 135 772
rect 139 768 140 772
rect 134 767 140 768
rect 111 766 115 767
rect 111 761 115 762
rect 135 766 139 767
rect 135 761 139 762
rect 112 758 114 761
rect 134 760 140 761
rect 110 757 116 758
rect 110 753 111 757
rect 115 753 116 757
rect 134 756 135 760
rect 139 756 140 760
rect 134 755 140 756
rect 110 752 116 753
rect 164 744 166 806
rect 176 801 178 813
rect 202 811 208 812
rect 202 807 203 811
rect 207 807 208 811
rect 202 806 208 807
rect 174 800 180 801
rect 174 796 175 800
rect 179 796 180 800
rect 174 795 180 796
rect 204 788 206 806
rect 216 801 218 813
rect 280 801 282 813
rect 322 811 328 812
rect 322 807 323 811
rect 327 807 328 811
rect 322 806 328 807
rect 214 800 220 801
rect 214 796 215 800
rect 219 796 220 800
rect 214 795 220 796
rect 278 800 284 801
rect 278 796 279 800
rect 283 796 284 800
rect 278 795 284 796
rect 324 788 326 806
rect 336 801 338 813
rect 378 811 384 812
rect 378 807 379 811
rect 383 807 384 811
rect 378 806 384 807
rect 334 800 340 801
rect 334 796 335 800
rect 339 796 340 800
rect 334 795 340 796
rect 380 788 382 806
rect 392 801 394 813
rect 408 812 410 842
rect 462 836 468 837
rect 462 832 463 836
rect 467 832 468 836
rect 462 831 468 832
rect 464 819 466 831
rect 455 818 459 819
rect 455 813 459 814
rect 463 818 467 819
rect 463 813 467 814
rect 406 811 412 812
rect 406 807 407 811
rect 411 807 412 811
rect 406 806 412 807
rect 456 801 458 813
rect 472 812 474 842
rect 534 836 540 837
rect 534 832 535 836
rect 539 832 540 836
rect 534 831 540 832
rect 479 828 483 829
rect 478 823 484 824
rect 478 819 479 823
rect 483 819 484 823
rect 536 819 538 831
rect 608 824 610 842
rect 614 836 620 837
rect 614 832 615 836
rect 619 832 620 836
rect 614 831 620 832
rect 598 823 604 824
rect 598 819 599 823
rect 603 819 604 823
rect 478 818 484 819
rect 519 818 523 819
rect 519 813 523 814
rect 535 818 539 819
rect 535 813 539 814
rect 583 818 587 819
rect 598 818 604 819
rect 606 823 612 824
rect 606 819 607 823
rect 611 819 612 823
rect 616 819 618 831
rect 704 824 706 842
rect 710 836 716 837
rect 710 832 711 836
rect 715 832 716 836
rect 710 831 716 832
rect 822 836 828 837
rect 822 832 823 836
rect 827 832 828 836
rect 822 831 828 832
rect 702 823 708 824
rect 702 819 703 823
rect 707 819 708 823
rect 712 819 714 831
rect 824 819 826 831
rect 860 829 862 842
rect 859 828 863 829
rect 842 823 848 824
rect 859 823 863 824
rect 842 819 843 823
rect 847 819 848 823
rect 606 818 612 819
rect 615 818 619 819
rect 583 813 587 814
rect 470 811 476 812
rect 470 807 471 811
rect 475 807 476 811
rect 470 806 476 807
rect 482 811 488 812
rect 482 807 483 811
rect 487 807 488 811
rect 482 806 488 807
rect 390 800 396 801
rect 390 796 391 800
rect 395 796 396 800
rect 390 795 396 796
rect 454 800 460 801
rect 454 796 455 800
rect 459 796 460 800
rect 454 795 460 796
rect 484 788 486 806
rect 520 801 522 813
rect 546 811 552 812
rect 546 807 547 811
rect 551 807 552 811
rect 546 806 552 807
rect 518 800 524 801
rect 518 796 519 800
rect 523 796 524 800
rect 518 795 524 796
rect 548 788 550 806
rect 584 801 586 813
rect 582 800 588 801
rect 582 796 583 800
rect 587 796 588 800
rect 600 796 602 818
rect 615 813 619 814
rect 655 818 659 819
rect 702 818 708 819
rect 711 818 715 819
rect 655 813 659 814
rect 711 813 715 814
rect 735 818 739 819
rect 735 813 739 814
rect 815 818 819 819
rect 815 813 819 814
rect 823 818 827 819
rect 842 818 848 819
rect 895 818 899 819
rect 823 813 827 814
rect 656 801 658 813
rect 718 811 724 812
rect 718 807 719 811
rect 723 807 724 811
rect 718 806 724 807
rect 654 800 660 801
rect 654 796 655 800
rect 659 796 660 800
rect 582 795 588 796
rect 598 795 604 796
rect 654 795 660 796
rect 598 791 599 795
rect 603 791 604 795
rect 598 790 604 791
rect 202 787 208 788
rect 202 783 203 787
rect 207 783 208 787
rect 202 782 208 783
rect 322 787 328 788
rect 322 783 323 787
rect 327 783 328 787
rect 322 782 328 783
rect 378 787 384 788
rect 378 783 379 787
rect 383 783 384 787
rect 378 782 384 783
rect 482 787 488 788
rect 482 783 483 787
rect 487 783 488 787
rect 482 782 488 783
rect 546 787 552 788
rect 546 783 547 787
rect 551 783 552 787
rect 546 782 552 783
rect 554 787 560 788
rect 554 783 555 787
rect 559 783 560 787
rect 554 782 560 783
rect 174 772 180 773
rect 174 768 175 772
rect 179 768 180 772
rect 174 767 180 768
rect 214 772 220 773
rect 214 768 215 772
rect 219 768 220 772
rect 214 767 220 768
rect 278 772 284 773
rect 278 768 279 772
rect 283 768 284 772
rect 278 767 284 768
rect 334 772 340 773
rect 334 768 335 772
rect 339 768 340 772
rect 334 767 340 768
rect 390 772 396 773
rect 390 768 391 772
rect 395 768 396 772
rect 390 767 396 768
rect 454 772 460 773
rect 454 768 455 772
rect 459 768 460 772
rect 454 767 460 768
rect 518 772 524 773
rect 518 768 519 772
rect 523 768 524 772
rect 518 767 524 768
rect 175 766 179 767
rect 175 761 179 762
rect 207 766 211 767
rect 207 761 211 762
rect 215 766 219 767
rect 215 761 219 762
rect 279 766 283 767
rect 279 761 283 762
rect 295 766 299 767
rect 295 761 299 762
rect 335 766 339 767
rect 335 761 339 762
rect 375 766 379 767
rect 375 761 379 762
rect 391 766 395 767
rect 391 761 395 762
rect 447 766 451 767
rect 447 761 451 762
rect 455 766 459 767
rect 455 761 459 762
rect 519 766 523 767
rect 519 761 523 762
rect 206 760 212 761
rect 206 756 207 760
rect 211 756 212 760
rect 206 755 212 756
rect 294 760 300 761
rect 294 756 295 760
rect 299 756 300 760
rect 294 755 300 756
rect 374 760 380 761
rect 374 756 375 760
rect 379 756 380 760
rect 374 755 380 756
rect 446 760 452 761
rect 446 756 447 760
rect 451 756 452 760
rect 446 755 452 756
rect 518 760 524 761
rect 518 756 519 760
rect 523 756 524 760
rect 518 755 524 756
rect 162 743 168 744
rect 110 740 116 741
rect 110 736 111 740
rect 115 736 116 740
rect 162 739 163 743
rect 167 739 168 743
rect 162 738 168 739
rect 286 743 292 744
rect 286 739 287 743
rect 291 739 292 743
rect 286 738 292 739
rect 318 743 324 744
rect 318 739 319 743
rect 323 739 324 743
rect 318 738 324 739
rect 390 743 396 744
rect 390 739 391 743
rect 395 739 396 743
rect 390 738 396 739
rect 418 743 424 744
rect 418 739 419 743
rect 423 739 424 743
rect 418 738 424 739
rect 110 735 116 736
rect 112 711 114 735
rect 134 732 140 733
rect 134 728 135 732
rect 139 728 140 732
rect 134 727 140 728
rect 206 732 212 733
rect 206 728 207 732
rect 211 728 212 732
rect 206 727 212 728
rect 136 711 138 727
rect 158 719 164 720
rect 158 715 159 719
rect 163 715 164 719
rect 158 714 164 715
rect 111 710 115 711
rect 111 705 115 706
rect 135 710 139 711
rect 135 705 139 706
rect 112 685 114 705
rect 136 693 138 705
rect 134 692 140 693
rect 134 688 135 692
rect 139 688 140 692
rect 134 687 140 688
rect 110 684 116 685
rect 110 680 111 684
rect 115 680 116 684
rect 160 680 162 714
rect 208 711 210 727
rect 288 720 290 738
rect 294 732 300 733
rect 294 728 295 732
rect 299 728 300 732
rect 294 727 300 728
rect 286 719 292 720
rect 286 715 287 719
rect 291 715 292 719
rect 286 714 292 715
rect 296 711 298 727
rect 183 710 187 711
rect 183 705 187 706
rect 207 710 211 711
rect 207 705 211 706
rect 247 710 251 711
rect 247 705 251 706
rect 295 710 299 711
rect 295 705 299 706
rect 311 710 315 711
rect 311 705 315 706
rect 170 703 176 704
rect 170 699 171 703
rect 175 699 176 703
rect 170 698 176 699
rect 172 680 174 698
rect 184 693 186 705
rect 234 703 240 704
rect 234 699 235 703
rect 239 699 240 703
rect 234 698 240 699
rect 182 692 188 693
rect 182 688 183 692
rect 187 688 188 692
rect 182 687 188 688
rect 110 679 116 680
rect 158 679 164 680
rect 158 675 159 679
rect 163 675 164 679
rect 158 674 164 675
rect 170 679 176 680
rect 170 675 171 679
rect 175 675 176 679
rect 170 674 176 675
rect 110 667 116 668
rect 110 663 111 667
rect 115 663 116 667
rect 110 662 116 663
rect 134 664 140 665
rect 112 651 114 662
rect 134 660 135 664
rect 139 660 140 664
rect 134 659 140 660
rect 182 664 188 665
rect 182 660 183 664
rect 187 660 188 664
rect 182 659 188 660
rect 136 651 138 659
rect 184 651 186 659
rect 111 650 115 651
rect 111 645 115 646
rect 135 650 139 651
rect 135 645 139 646
rect 159 650 163 651
rect 159 645 163 646
rect 183 650 187 651
rect 183 645 187 646
rect 215 650 219 651
rect 215 645 219 646
rect 112 642 114 645
rect 158 644 164 645
rect 110 641 116 642
rect 110 637 111 641
rect 115 637 116 641
rect 158 640 159 644
rect 163 640 164 644
rect 158 639 164 640
rect 214 644 220 645
rect 214 640 215 644
rect 219 640 220 644
rect 214 639 220 640
rect 110 636 116 637
rect 236 628 238 698
rect 248 693 250 705
rect 282 703 288 704
rect 282 699 283 703
rect 287 699 288 703
rect 282 698 288 699
rect 246 692 252 693
rect 246 688 247 692
rect 251 688 252 692
rect 246 687 252 688
rect 284 680 286 698
rect 312 693 314 705
rect 320 704 322 738
rect 374 732 380 733
rect 374 728 375 732
rect 379 728 380 732
rect 374 727 380 728
rect 376 711 378 727
rect 375 710 379 711
rect 375 705 379 706
rect 383 710 387 711
rect 383 705 387 706
rect 318 703 324 704
rect 318 699 319 703
rect 323 699 324 703
rect 318 698 324 699
rect 384 693 386 705
rect 392 704 394 738
rect 420 720 422 738
rect 446 732 452 733
rect 446 728 447 732
rect 451 728 452 732
rect 446 727 452 728
rect 518 732 524 733
rect 518 728 519 732
rect 523 728 524 732
rect 518 727 524 728
rect 418 719 424 720
rect 418 715 419 719
rect 423 715 424 719
rect 418 714 424 715
rect 448 711 450 727
rect 520 711 522 727
rect 556 720 558 782
rect 582 772 588 773
rect 582 768 583 772
rect 587 768 588 772
rect 582 767 588 768
rect 654 772 660 773
rect 654 768 655 772
rect 659 768 660 772
rect 654 767 660 768
rect 583 766 587 767
rect 583 761 587 762
rect 639 766 643 767
rect 639 761 643 762
rect 655 766 659 767
rect 655 761 659 762
rect 687 766 691 767
rect 687 761 691 762
rect 582 760 588 761
rect 582 756 583 760
rect 587 756 588 760
rect 582 755 588 756
rect 638 760 644 761
rect 638 756 639 760
rect 643 756 644 760
rect 638 755 644 756
rect 686 760 692 761
rect 686 756 687 760
rect 691 756 692 760
rect 686 755 692 756
rect 720 744 722 806
rect 736 801 738 813
rect 762 811 768 812
rect 762 807 763 811
rect 767 807 768 811
rect 762 806 768 807
rect 734 800 740 801
rect 734 796 735 800
rect 739 796 740 800
rect 734 795 740 796
rect 764 788 766 806
rect 816 801 818 813
rect 814 800 820 801
rect 814 796 815 800
rect 819 796 820 800
rect 814 795 820 796
rect 844 788 846 818
rect 895 813 899 814
rect 896 801 898 813
rect 904 812 906 850
rect 942 836 948 837
rect 942 832 943 836
rect 947 832 948 836
rect 942 831 948 832
rect 1046 836 1052 837
rect 1046 832 1047 836
rect 1051 832 1052 836
rect 1088 832 1090 890
rect 1134 888 1135 892
rect 1139 888 1140 892
rect 1364 888 1366 906
rect 1376 901 1378 913
rect 1384 912 1386 946
rect 1438 940 1444 941
rect 1438 936 1439 940
rect 1443 936 1444 940
rect 1438 935 1444 936
rect 1440 919 1442 935
rect 1504 928 1506 946
rect 1510 940 1516 941
rect 1510 936 1511 940
rect 1515 936 1516 940
rect 1510 935 1516 936
rect 1582 940 1588 941
rect 1582 936 1583 940
rect 1587 936 1588 940
rect 1582 935 1588 936
rect 1446 927 1452 928
rect 1446 923 1447 927
rect 1451 923 1452 927
rect 1446 922 1452 923
rect 1502 927 1508 928
rect 1502 923 1503 927
rect 1507 923 1508 927
rect 1502 922 1508 923
rect 1423 918 1427 919
rect 1423 913 1427 914
rect 1439 918 1443 919
rect 1439 913 1443 914
rect 1382 911 1388 912
rect 1382 907 1383 911
rect 1387 907 1388 911
rect 1382 906 1388 907
rect 1424 901 1426 913
rect 1374 900 1380 901
rect 1374 896 1375 900
rect 1379 896 1380 900
rect 1374 895 1380 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1448 888 1450 922
rect 1512 919 1514 935
rect 1584 919 1586 935
rect 1612 928 1614 954
rect 1646 951 1652 952
rect 1646 947 1647 951
rect 1651 947 1652 951
rect 1646 946 1652 947
rect 1718 951 1724 952
rect 1718 947 1719 951
rect 1723 947 1724 951
rect 1718 946 1724 947
rect 1778 951 1784 952
rect 1778 947 1779 951
rect 1783 947 1784 951
rect 1778 946 1784 947
rect 1648 928 1650 946
rect 1654 940 1660 941
rect 1654 936 1655 940
rect 1659 936 1660 940
rect 1654 935 1660 936
rect 1610 927 1616 928
rect 1610 923 1611 927
rect 1615 923 1616 927
rect 1610 922 1616 923
rect 1646 927 1652 928
rect 1646 923 1647 927
rect 1651 923 1652 927
rect 1646 922 1652 923
rect 1656 919 1658 935
rect 1720 928 1722 946
rect 1726 940 1732 941
rect 1726 936 1727 940
rect 1731 936 1732 940
rect 1726 935 1732 936
rect 1718 927 1724 928
rect 1718 923 1719 927
rect 1723 923 1724 927
rect 1718 922 1724 923
rect 1728 919 1730 935
rect 1479 918 1483 919
rect 1479 913 1483 914
rect 1511 918 1515 919
rect 1511 913 1515 914
rect 1551 918 1555 919
rect 1551 913 1555 914
rect 1583 918 1587 919
rect 1583 913 1587 914
rect 1623 918 1627 919
rect 1623 913 1627 914
rect 1655 918 1659 919
rect 1655 913 1659 914
rect 1703 918 1707 919
rect 1703 913 1707 914
rect 1727 918 1731 919
rect 1727 913 1731 914
rect 1466 911 1472 912
rect 1466 907 1467 911
rect 1471 907 1472 911
rect 1466 906 1472 907
rect 1468 888 1470 906
rect 1480 901 1482 913
rect 1494 911 1500 912
rect 1494 907 1495 911
rect 1499 907 1500 911
rect 1494 906 1500 907
rect 1478 900 1484 901
rect 1478 896 1479 900
rect 1483 896 1484 900
rect 1478 895 1484 896
rect 1134 887 1140 888
rect 1206 887 1212 888
rect 1094 883 1100 884
rect 1094 879 1095 883
rect 1099 879 1100 883
rect 1206 883 1207 887
rect 1211 883 1212 887
rect 1206 882 1212 883
rect 1362 887 1368 888
rect 1362 883 1363 887
rect 1367 883 1368 887
rect 1362 882 1368 883
rect 1446 887 1452 888
rect 1446 883 1447 887
rect 1451 883 1452 887
rect 1446 882 1452 883
rect 1466 887 1472 888
rect 1466 883 1467 887
rect 1471 883 1472 887
rect 1466 882 1472 883
rect 1094 878 1100 879
rect 1096 871 1098 878
rect 1134 875 1140 876
rect 1134 871 1135 875
rect 1139 871 1140 875
rect 1095 870 1099 871
rect 1134 870 1140 871
rect 1136 867 1138 870
rect 1095 865 1099 866
rect 1135 866 1139 867
rect 1096 862 1098 865
rect 1094 861 1100 862
rect 1135 861 1139 862
rect 1159 866 1163 867
rect 1159 861 1163 862
rect 1199 866 1203 867
rect 1199 861 1203 862
rect 1094 857 1095 861
rect 1099 857 1100 861
rect 1136 858 1138 861
rect 1158 860 1164 861
rect 1094 856 1100 857
rect 1134 857 1140 858
rect 1134 853 1135 857
rect 1139 853 1140 857
rect 1158 856 1159 860
rect 1163 856 1164 860
rect 1158 855 1164 856
rect 1198 860 1204 861
rect 1198 856 1199 860
rect 1203 856 1204 860
rect 1198 855 1204 856
rect 1134 852 1140 853
rect 1094 844 1100 845
rect 1094 840 1095 844
rect 1099 840 1100 844
rect 1142 843 1148 844
rect 1094 839 1100 840
rect 1134 840 1140 841
rect 1046 831 1052 832
rect 1086 831 1092 832
rect 944 819 946 831
rect 1048 819 1050 831
rect 1086 827 1087 831
rect 1091 827 1092 831
rect 1086 826 1092 827
rect 1096 819 1098 839
rect 1134 836 1135 840
rect 1139 836 1140 840
rect 1142 839 1143 843
rect 1147 839 1148 843
rect 1142 838 1148 839
rect 1134 835 1140 836
rect 943 818 947 819
rect 943 813 947 814
rect 983 818 987 819
rect 983 813 987 814
rect 1047 818 1051 819
rect 1047 813 1051 814
rect 1095 818 1099 819
rect 1095 813 1099 814
rect 902 811 908 812
rect 902 807 903 811
rect 907 807 908 811
rect 902 806 908 807
rect 922 811 928 812
rect 922 807 923 811
rect 927 807 928 811
rect 922 806 928 807
rect 894 800 900 801
rect 894 796 895 800
rect 899 796 900 800
rect 894 795 900 796
rect 924 788 926 806
rect 984 801 986 813
rect 1010 811 1016 812
rect 1010 807 1011 811
rect 1015 807 1016 811
rect 1010 806 1016 807
rect 982 800 988 801
rect 982 796 983 800
rect 987 796 988 800
rect 982 795 988 796
rect 1012 788 1014 806
rect 1048 801 1050 813
rect 1046 800 1052 801
rect 1046 796 1047 800
rect 1051 796 1052 800
rect 1046 795 1052 796
rect 1096 793 1098 813
rect 1136 807 1138 835
rect 1144 824 1146 838
rect 1158 832 1164 833
rect 1158 828 1159 832
rect 1163 828 1164 832
rect 1158 827 1164 828
rect 1198 832 1204 833
rect 1198 828 1199 832
rect 1203 828 1204 832
rect 1198 827 1204 828
rect 1142 823 1148 824
rect 1142 819 1143 823
rect 1147 819 1148 823
rect 1142 818 1148 819
rect 1160 807 1162 827
rect 1200 807 1202 827
rect 1208 820 1210 882
rect 1286 872 1292 873
rect 1286 868 1287 872
rect 1291 868 1292 872
rect 1286 867 1292 868
rect 1326 872 1332 873
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 1326 867 1332 868
rect 1374 872 1380 873
rect 1374 868 1375 872
rect 1379 868 1380 872
rect 1374 867 1380 868
rect 1422 872 1428 873
rect 1422 868 1423 872
rect 1427 868 1428 872
rect 1422 867 1428 868
rect 1478 872 1484 873
rect 1478 868 1479 872
rect 1483 868 1484 872
rect 1478 867 1484 868
rect 1263 866 1267 867
rect 1263 861 1267 862
rect 1287 866 1291 867
rect 1287 861 1291 862
rect 1327 866 1331 867
rect 1327 861 1331 862
rect 1375 866 1379 867
rect 1375 861 1379 862
rect 1399 866 1403 867
rect 1399 861 1403 862
rect 1423 866 1427 867
rect 1423 861 1427 862
rect 1471 866 1475 867
rect 1471 861 1475 862
rect 1479 866 1483 867
rect 1479 861 1483 862
rect 1262 860 1268 861
rect 1262 856 1263 860
rect 1267 856 1268 860
rect 1262 855 1268 856
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1398 860 1404 861
rect 1398 856 1399 860
rect 1403 856 1404 860
rect 1398 855 1404 856
rect 1470 860 1476 861
rect 1470 856 1471 860
rect 1475 856 1476 860
rect 1470 855 1476 856
rect 1496 844 1498 906
rect 1552 901 1554 913
rect 1610 911 1616 912
rect 1610 907 1611 911
rect 1615 907 1616 911
rect 1610 906 1616 907
rect 1550 900 1556 901
rect 1550 896 1551 900
rect 1555 896 1556 900
rect 1550 895 1556 896
rect 1612 888 1614 906
rect 1624 901 1626 913
rect 1690 911 1696 912
rect 1690 907 1691 911
rect 1695 907 1696 911
rect 1690 906 1696 907
rect 1622 900 1628 901
rect 1622 896 1623 900
rect 1627 896 1628 900
rect 1622 895 1628 896
rect 1692 888 1694 906
rect 1704 901 1706 913
rect 1780 912 1782 946
rect 1788 928 1790 990
rect 2118 983 2124 984
rect 1822 980 1828 981
rect 1822 976 1823 980
rect 1827 976 1828 980
rect 1822 975 1828 976
rect 1886 980 1892 981
rect 1886 976 1887 980
rect 1891 976 1892 980
rect 1886 975 1892 976
rect 1950 980 1956 981
rect 1950 976 1951 980
rect 1955 976 1956 980
rect 2118 979 2119 983
rect 2123 979 2124 983
rect 2118 978 2124 979
rect 1950 975 1956 976
rect 2120 975 2122 978
rect 1799 974 1803 975
rect 1799 969 1803 970
rect 1823 974 1827 975
rect 1823 969 1827 970
rect 1871 974 1875 975
rect 1871 969 1875 970
rect 1887 974 1891 975
rect 1887 969 1891 970
rect 1943 974 1947 975
rect 1943 969 1947 970
rect 1951 974 1955 975
rect 1951 969 1955 970
rect 2015 974 2019 975
rect 2015 969 2019 970
rect 2071 974 2075 975
rect 2071 969 2075 970
rect 2119 974 2123 975
rect 2119 969 2123 970
rect 1798 968 1804 969
rect 1798 964 1799 968
rect 1803 964 1804 968
rect 1798 963 1804 964
rect 1870 968 1876 969
rect 1870 964 1871 968
rect 1875 964 1876 968
rect 1870 963 1876 964
rect 1942 968 1948 969
rect 1942 964 1943 968
rect 1947 964 1948 968
rect 1942 963 1948 964
rect 2014 968 2020 969
rect 2014 964 2015 968
rect 2019 964 2020 968
rect 2014 963 2020 964
rect 2070 968 2076 969
rect 2070 964 2071 968
rect 2075 964 2076 968
rect 2120 966 2122 969
rect 2070 963 2076 964
rect 2118 965 2124 966
rect 2118 961 2119 965
rect 2123 961 2124 965
rect 2118 960 2124 961
rect 1862 951 1868 952
rect 1862 947 1863 951
rect 1867 947 1868 951
rect 1862 946 1868 947
rect 1990 951 1996 952
rect 1990 947 1991 951
rect 1995 947 1996 951
rect 1990 946 1996 947
rect 2118 948 2124 949
rect 1798 940 1804 941
rect 1798 936 1799 940
rect 1803 936 1804 940
rect 1798 935 1804 936
rect 1786 927 1792 928
rect 1786 923 1787 927
rect 1791 923 1792 927
rect 1786 922 1792 923
rect 1800 919 1802 935
rect 1864 928 1866 946
rect 1870 940 1876 941
rect 1870 936 1871 940
rect 1875 936 1876 940
rect 1870 935 1876 936
rect 1942 940 1948 941
rect 1942 936 1943 940
rect 1947 936 1948 940
rect 1942 935 1948 936
rect 1862 927 1868 928
rect 1862 923 1863 927
rect 1867 923 1868 927
rect 1862 922 1868 923
rect 1872 919 1874 935
rect 1944 919 1946 935
rect 1992 928 1994 946
rect 2118 944 2119 948
rect 2123 944 2124 948
rect 2006 943 2012 944
rect 2118 943 2124 944
rect 2006 939 2007 943
rect 2011 939 2012 943
rect 2006 938 2012 939
rect 2014 940 2020 941
rect 1990 927 1996 928
rect 1990 923 1991 927
rect 1995 923 1996 927
rect 1990 922 1996 923
rect 1791 918 1795 919
rect 1791 913 1795 914
rect 1799 918 1803 919
rect 1799 913 1803 914
rect 1871 918 1875 919
rect 1871 913 1875 914
rect 1879 918 1883 919
rect 1879 913 1883 914
rect 1943 918 1947 919
rect 1943 913 1947 914
rect 1967 918 1971 919
rect 1967 913 1971 914
rect 1770 911 1776 912
rect 1770 907 1771 911
rect 1775 907 1776 911
rect 1770 906 1776 907
rect 1778 911 1784 912
rect 1778 907 1779 911
rect 1783 907 1784 911
rect 1778 906 1784 907
rect 1702 900 1708 901
rect 1702 896 1703 900
rect 1707 896 1708 900
rect 1702 895 1708 896
rect 1772 888 1774 906
rect 1792 901 1794 913
rect 1870 907 1876 908
rect 1870 903 1871 907
rect 1875 903 1876 907
rect 1870 902 1876 903
rect 1790 900 1796 901
rect 1790 896 1791 900
rect 1795 896 1796 900
rect 1790 895 1796 896
rect 1558 887 1564 888
rect 1558 883 1559 887
rect 1563 883 1564 887
rect 1558 882 1564 883
rect 1610 887 1616 888
rect 1610 883 1611 887
rect 1615 883 1616 887
rect 1610 882 1616 883
rect 1690 887 1696 888
rect 1690 883 1691 887
rect 1695 883 1696 887
rect 1690 882 1696 883
rect 1770 887 1776 888
rect 1770 883 1771 887
rect 1775 883 1776 887
rect 1770 882 1776 883
rect 1550 872 1556 873
rect 1550 868 1551 872
rect 1555 868 1556 872
rect 1550 867 1556 868
rect 1543 866 1547 867
rect 1543 861 1547 862
rect 1551 866 1555 867
rect 1551 861 1555 862
rect 1542 860 1548 861
rect 1542 856 1543 860
rect 1547 856 1548 860
rect 1542 855 1548 856
rect 1254 843 1260 844
rect 1254 839 1255 843
rect 1259 839 1260 843
rect 1254 838 1260 839
rect 1318 843 1324 844
rect 1318 839 1319 843
rect 1323 839 1324 843
rect 1318 838 1324 839
rect 1390 843 1396 844
rect 1390 839 1391 843
rect 1395 839 1396 843
rect 1390 838 1396 839
rect 1462 843 1468 844
rect 1462 839 1463 843
rect 1467 839 1468 843
rect 1462 838 1468 839
rect 1494 843 1500 844
rect 1494 839 1495 843
rect 1499 839 1500 843
rect 1494 838 1500 839
rect 1256 820 1258 838
rect 1262 832 1268 833
rect 1262 828 1263 832
rect 1267 828 1268 832
rect 1262 827 1268 828
rect 1206 819 1212 820
rect 1206 815 1207 819
rect 1211 815 1212 819
rect 1206 814 1212 815
rect 1254 819 1260 820
rect 1254 815 1255 819
rect 1259 815 1260 819
rect 1254 814 1260 815
rect 1264 807 1266 827
rect 1320 820 1322 838
rect 1326 832 1332 833
rect 1326 828 1327 832
rect 1331 828 1332 832
rect 1326 827 1332 828
rect 1318 819 1324 820
rect 1318 815 1319 819
rect 1323 815 1324 819
rect 1318 814 1324 815
rect 1328 807 1330 827
rect 1392 820 1394 838
rect 1398 832 1404 833
rect 1398 828 1399 832
rect 1403 828 1404 832
rect 1398 827 1404 828
rect 1390 819 1396 820
rect 1390 815 1391 819
rect 1395 815 1396 819
rect 1390 814 1396 815
rect 1400 807 1402 827
rect 1464 820 1466 838
rect 1470 832 1476 833
rect 1470 828 1471 832
rect 1475 828 1476 832
rect 1470 827 1476 828
rect 1542 832 1548 833
rect 1542 828 1543 832
rect 1547 828 1548 832
rect 1542 827 1548 828
rect 1462 819 1468 820
rect 1462 815 1463 819
rect 1467 815 1468 819
rect 1462 814 1468 815
rect 1472 807 1474 827
rect 1544 807 1546 827
rect 1560 820 1562 882
rect 1622 872 1628 873
rect 1622 868 1623 872
rect 1627 868 1628 872
rect 1622 867 1628 868
rect 1702 872 1708 873
rect 1702 868 1703 872
rect 1707 868 1708 872
rect 1702 867 1708 868
rect 1790 872 1796 873
rect 1790 868 1791 872
rect 1795 868 1796 872
rect 1790 867 1796 868
rect 1623 866 1627 867
rect 1623 861 1627 862
rect 1703 866 1707 867
rect 1703 861 1707 862
rect 1775 866 1779 867
rect 1775 861 1779 862
rect 1791 866 1795 867
rect 1791 861 1795 862
rect 1855 866 1859 867
rect 1855 861 1859 862
rect 1622 860 1628 861
rect 1622 856 1623 860
rect 1627 856 1628 860
rect 1622 855 1628 856
rect 1702 860 1708 861
rect 1702 856 1703 860
rect 1707 856 1708 860
rect 1702 855 1708 856
rect 1774 860 1780 861
rect 1774 856 1775 860
rect 1779 856 1780 860
rect 1774 855 1780 856
rect 1854 860 1860 861
rect 1854 856 1855 860
rect 1859 856 1860 860
rect 1854 855 1860 856
rect 1872 844 1874 902
rect 1880 901 1882 913
rect 1906 911 1912 912
rect 1906 907 1907 911
rect 1911 907 1912 911
rect 1906 906 1912 907
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1908 888 1910 906
rect 1968 901 1970 913
rect 1994 911 2000 912
rect 1994 907 1995 911
rect 1999 907 2000 911
rect 1994 906 2000 907
rect 1966 900 1972 901
rect 1966 896 1967 900
rect 1971 896 1972 900
rect 1966 895 1972 896
rect 1996 888 1998 906
rect 1906 887 1912 888
rect 1906 883 1907 887
rect 1911 883 1912 887
rect 1906 882 1912 883
rect 1994 887 2000 888
rect 1994 883 1995 887
rect 1999 883 2000 887
rect 1994 882 2000 883
rect 1878 872 1884 873
rect 1878 868 1879 872
rect 1883 868 1884 872
rect 1878 867 1884 868
rect 1966 872 1972 873
rect 1966 868 1967 872
rect 1971 868 1972 872
rect 1966 867 1972 868
rect 1879 866 1883 867
rect 1879 861 1883 862
rect 1935 866 1939 867
rect 1935 861 1939 862
rect 1967 866 1971 867
rect 1967 861 1971 862
rect 1934 860 1940 861
rect 1934 856 1935 860
rect 1939 856 1940 860
rect 1934 855 1940 856
rect 1614 843 1620 844
rect 1614 839 1615 843
rect 1619 839 1620 843
rect 1614 838 1620 839
rect 1694 843 1700 844
rect 1694 839 1695 843
rect 1699 839 1700 843
rect 1694 838 1700 839
rect 1766 843 1772 844
rect 1766 839 1767 843
rect 1771 839 1772 843
rect 1766 838 1772 839
rect 1782 843 1788 844
rect 1782 839 1783 843
rect 1787 839 1788 843
rect 1782 838 1788 839
rect 1870 843 1876 844
rect 1870 839 1871 843
rect 1875 839 1876 843
rect 1870 838 1876 839
rect 1898 843 1904 844
rect 1898 839 1899 843
rect 1903 839 1904 843
rect 1898 838 1904 839
rect 1616 820 1618 838
rect 1622 832 1628 833
rect 1622 828 1623 832
rect 1627 828 1628 832
rect 1622 827 1628 828
rect 1558 819 1564 820
rect 1558 815 1559 819
rect 1563 815 1564 819
rect 1558 814 1564 815
rect 1614 819 1620 820
rect 1614 815 1615 819
rect 1619 815 1620 819
rect 1614 814 1620 815
rect 1624 807 1626 827
rect 1696 820 1698 838
rect 1702 832 1708 833
rect 1702 828 1703 832
rect 1707 828 1708 832
rect 1702 827 1708 828
rect 1694 819 1700 820
rect 1694 815 1695 819
rect 1699 815 1700 819
rect 1694 814 1700 815
rect 1704 807 1706 827
rect 1768 820 1770 838
rect 1774 832 1780 833
rect 1774 828 1775 832
rect 1779 828 1780 832
rect 1774 827 1780 828
rect 1766 819 1772 820
rect 1766 815 1767 819
rect 1771 815 1772 819
rect 1766 814 1772 815
rect 1776 807 1778 827
rect 1135 806 1139 807
rect 1135 801 1139 802
rect 1159 806 1163 807
rect 1159 801 1163 802
rect 1199 806 1203 807
rect 1199 801 1203 802
rect 1239 806 1243 807
rect 1239 801 1243 802
rect 1263 806 1267 807
rect 1263 801 1267 802
rect 1327 806 1331 807
rect 1327 801 1331 802
rect 1343 806 1347 807
rect 1343 801 1347 802
rect 1399 806 1403 807
rect 1399 801 1403 802
rect 1447 806 1451 807
rect 1447 801 1451 802
rect 1471 806 1475 807
rect 1471 801 1475 802
rect 1543 806 1547 807
rect 1543 801 1547 802
rect 1551 806 1555 807
rect 1551 801 1555 802
rect 1623 806 1627 807
rect 1623 801 1627 802
rect 1655 806 1659 807
rect 1655 801 1659 802
rect 1703 806 1707 807
rect 1703 801 1707 802
rect 1751 806 1755 807
rect 1751 801 1755 802
rect 1775 806 1779 807
rect 1775 801 1779 802
rect 1094 792 1100 793
rect 1094 788 1095 792
rect 1099 788 1100 792
rect 762 787 768 788
rect 762 783 763 787
rect 767 783 768 787
rect 762 782 768 783
rect 842 787 848 788
rect 842 783 843 787
rect 847 783 848 787
rect 842 782 848 783
rect 922 787 928 788
rect 922 783 923 787
rect 927 783 928 787
rect 922 782 928 783
rect 1010 787 1016 788
rect 1094 787 1100 788
rect 1010 783 1011 787
rect 1015 783 1016 787
rect 1010 782 1016 783
rect 1136 781 1138 801
rect 1160 789 1162 801
rect 1186 799 1192 800
rect 1186 795 1187 799
rect 1191 795 1192 799
rect 1186 794 1192 795
rect 1158 788 1164 789
rect 1158 784 1159 788
rect 1163 784 1164 788
rect 1158 783 1164 784
rect 1134 780 1140 781
rect 1134 776 1135 780
rect 1139 776 1140 780
rect 1188 776 1190 794
rect 1240 789 1242 801
rect 1302 799 1308 800
rect 1302 795 1303 799
rect 1307 795 1308 799
rect 1302 794 1308 795
rect 1238 788 1244 789
rect 1238 784 1239 788
rect 1243 784 1244 788
rect 1238 783 1244 784
rect 1304 780 1306 794
rect 1344 789 1346 801
rect 1448 789 1450 801
rect 1552 789 1554 801
rect 1642 799 1648 800
rect 1642 795 1643 799
rect 1647 795 1648 799
rect 1642 794 1648 795
rect 1342 788 1348 789
rect 1342 784 1343 788
rect 1347 784 1348 788
rect 1342 783 1348 784
rect 1446 788 1452 789
rect 1446 784 1447 788
rect 1451 784 1452 788
rect 1446 783 1452 784
rect 1550 788 1556 789
rect 1550 784 1551 788
rect 1555 784 1556 788
rect 1550 783 1556 784
rect 1302 779 1308 780
rect 1094 775 1100 776
rect 1134 775 1140 776
rect 1186 775 1192 776
rect 734 772 740 773
rect 734 768 735 772
rect 739 768 740 772
rect 734 767 740 768
rect 814 772 820 773
rect 814 768 815 772
rect 819 768 820 772
rect 814 767 820 768
rect 894 772 900 773
rect 894 768 895 772
rect 899 768 900 772
rect 894 767 900 768
rect 982 772 988 773
rect 982 768 983 772
rect 987 768 988 772
rect 982 767 988 768
rect 1046 772 1052 773
rect 1046 768 1047 772
rect 1051 768 1052 772
rect 1094 771 1095 775
rect 1099 771 1100 775
rect 1094 770 1100 771
rect 1186 771 1187 775
rect 1191 771 1192 775
rect 1302 775 1303 779
rect 1307 775 1308 779
rect 1644 776 1646 794
rect 1656 789 1658 801
rect 1738 799 1744 800
rect 1738 795 1739 799
rect 1743 795 1744 799
rect 1738 794 1744 795
rect 1654 788 1660 789
rect 1654 784 1655 788
rect 1659 784 1660 788
rect 1654 783 1660 784
rect 1740 776 1742 794
rect 1752 789 1754 801
rect 1784 800 1786 838
rect 1854 832 1860 833
rect 1854 828 1855 832
rect 1859 828 1860 832
rect 1854 827 1860 828
rect 1856 807 1858 827
rect 1900 820 1902 838
rect 1934 832 1940 833
rect 1934 828 1935 832
rect 1939 828 1940 832
rect 1934 827 1940 828
rect 1898 819 1904 820
rect 1898 815 1899 819
rect 1903 815 1904 819
rect 1898 814 1904 815
rect 1936 807 1938 827
rect 2008 820 2010 938
rect 2014 936 2015 940
rect 2019 936 2020 940
rect 2014 935 2020 936
rect 2070 940 2076 941
rect 2070 936 2071 940
rect 2075 936 2076 940
rect 2070 935 2076 936
rect 2016 919 2018 935
rect 2072 919 2074 935
rect 2086 927 2092 928
rect 2086 923 2087 927
rect 2091 923 2092 927
rect 2086 922 2092 923
rect 2015 918 2019 919
rect 2015 913 2019 914
rect 2063 918 2067 919
rect 2063 913 2067 914
rect 2071 918 2075 919
rect 2071 913 2075 914
rect 2064 901 2066 913
rect 2062 900 2068 901
rect 2062 896 2063 900
rect 2067 896 2068 900
rect 2062 895 2068 896
rect 2088 888 2090 922
rect 2120 919 2122 943
rect 2119 918 2123 919
rect 2119 913 2123 914
rect 2120 893 2122 913
rect 2118 892 2124 893
rect 2118 888 2119 892
rect 2123 888 2124 892
rect 2086 887 2092 888
rect 2118 887 2124 888
rect 2086 883 2087 887
rect 2091 883 2092 887
rect 2086 882 2092 883
rect 2118 875 2124 876
rect 2062 872 2068 873
rect 2062 868 2063 872
rect 2067 868 2068 872
rect 2118 871 2119 875
rect 2123 871 2124 875
rect 2118 870 2124 871
rect 2062 867 2068 868
rect 2120 867 2122 870
rect 2015 866 2019 867
rect 2015 861 2019 862
rect 2063 866 2067 867
rect 2063 861 2067 862
rect 2071 866 2075 867
rect 2071 861 2075 862
rect 2119 866 2123 867
rect 2119 861 2123 862
rect 2014 860 2020 861
rect 2014 856 2015 860
rect 2019 856 2020 860
rect 2014 855 2020 856
rect 2070 860 2076 861
rect 2070 856 2071 860
rect 2075 856 2076 860
rect 2120 858 2122 861
rect 2070 855 2076 856
rect 2118 857 2124 858
rect 2118 853 2119 857
rect 2123 853 2124 857
rect 2118 852 2124 853
rect 2062 843 2068 844
rect 2062 839 2063 843
rect 2067 839 2068 843
rect 2062 838 2068 839
rect 2078 843 2084 844
rect 2078 839 2079 843
rect 2083 839 2084 843
rect 2078 838 2084 839
rect 2118 840 2124 841
rect 2014 832 2020 833
rect 2014 828 2015 832
rect 2019 828 2020 832
rect 2014 827 2020 828
rect 1998 819 2004 820
rect 1998 815 1999 819
rect 2003 815 2004 819
rect 1998 814 2004 815
rect 2006 819 2012 820
rect 2006 815 2007 819
rect 2011 815 2012 819
rect 2006 814 2012 815
rect 1839 806 1843 807
rect 1839 801 1843 802
rect 1855 806 1859 807
rect 1855 801 1859 802
rect 1919 806 1923 807
rect 1919 801 1923 802
rect 1935 806 1939 807
rect 1935 801 1939 802
rect 1782 799 1788 800
rect 1782 795 1783 799
rect 1787 795 1788 799
rect 1782 794 1788 795
rect 1830 799 1836 800
rect 1830 795 1831 799
rect 1835 795 1836 799
rect 1830 794 1836 795
rect 1750 788 1756 789
rect 1750 784 1751 788
rect 1755 784 1756 788
rect 1750 783 1756 784
rect 1302 774 1308 775
rect 1310 775 1316 776
rect 1186 770 1192 771
rect 1310 771 1311 775
rect 1315 771 1316 775
rect 1310 770 1316 771
rect 1518 775 1524 776
rect 1518 771 1519 775
rect 1523 771 1524 775
rect 1518 770 1524 771
rect 1642 775 1648 776
rect 1642 771 1643 775
rect 1647 771 1648 775
rect 1642 770 1648 771
rect 1738 775 1744 776
rect 1738 771 1739 775
rect 1743 771 1744 775
rect 1738 770 1744 771
rect 1046 767 1052 768
rect 1096 767 1098 770
rect 735 766 739 767
rect 735 761 739 762
rect 743 766 747 767
rect 743 761 747 762
rect 799 766 803 767
rect 799 761 803 762
rect 815 766 819 767
rect 815 761 819 762
rect 855 766 859 767
rect 855 761 859 762
rect 895 766 899 767
rect 895 761 899 762
rect 983 766 987 767
rect 983 761 987 762
rect 1047 766 1051 767
rect 1047 761 1051 762
rect 1095 766 1099 767
rect 1095 761 1099 762
rect 1134 763 1140 764
rect 742 760 748 761
rect 742 756 743 760
rect 747 756 748 760
rect 742 755 748 756
rect 798 760 804 761
rect 798 756 799 760
rect 803 756 804 760
rect 798 755 804 756
rect 854 760 860 761
rect 854 756 855 760
rect 859 756 860 760
rect 1096 758 1098 761
rect 1134 759 1135 763
rect 1139 759 1140 763
rect 1134 758 1140 759
rect 1158 760 1164 761
rect 854 755 860 756
rect 1094 757 1100 758
rect 1094 753 1095 757
rect 1099 753 1100 757
rect 1136 755 1138 758
rect 1158 756 1159 760
rect 1163 756 1164 760
rect 1158 755 1164 756
rect 1238 760 1244 761
rect 1238 756 1239 760
rect 1243 756 1244 760
rect 1238 755 1244 756
rect 1094 752 1100 753
rect 1135 754 1139 755
rect 1135 749 1139 750
rect 1159 754 1163 755
rect 1159 749 1163 750
rect 1199 754 1203 755
rect 1199 749 1203 750
rect 1239 754 1243 755
rect 1239 749 1243 750
rect 1287 754 1291 755
rect 1287 749 1291 750
rect 1136 746 1138 749
rect 1158 748 1164 749
rect 1134 745 1140 746
rect 678 743 684 744
rect 678 739 679 743
rect 683 739 684 743
rect 678 738 684 739
rect 714 743 722 744
rect 714 739 715 743
rect 719 740 722 743
rect 726 743 732 744
rect 719 739 720 740
rect 714 738 720 739
rect 726 739 727 743
rect 731 739 732 743
rect 726 738 732 739
rect 846 743 852 744
rect 846 739 847 743
rect 851 739 852 743
rect 846 738 852 739
rect 862 743 868 744
rect 862 739 863 743
rect 867 739 868 743
rect 1134 741 1135 745
rect 1139 741 1140 745
rect 1158 744 1159 748
rect 1163 744 1164 748
rect 1158 743 1164 744
rect 1198 748 1204 749
rect 1198 744 1199 748
rect 1203 744 1204 748
rect 1198 743 1204 744
rect 1238 748 1244 749
rect 1238 744 1239 748
rect 1243 744 1244 748
rect 1238 743 1244 744
rect 1286 748 1292 749
rect 1286 744 1287 748
rect 1291 744 1292 748
rect 1286 743 1292 744
rect 862 738 868 739
rect 1094 740 1100 741
rect 1134 740 1140 741
rect 582 732 588 733
rect 582 728 583 732
rect 587 728 588 732
rect 582 727 588 728
rect 638 732 644 733
rect 638 728 639 732
rect 643 728 644 732
rect 638 727 644 728
rect 554 719 560 720
rect 554 715 555 719
rect 559 715 560 719
rect 554 714 560 715
rect 584 711 586 727
rect 606 719 612 720
rect 606 715 607 719
rect 611 715 612 719
rect 606 714 612 715
rect 447 710 451 711
rect 447 705 451 706
rect 455 710 459 711
rect 455 705 459 706
rect 519 710 523 711
rect 519 705 523 706
rect 583 710 587 711
rect 583 705 587 706
rect 390 703 396 704
rect 390 699 391 703
rect 395 699 396 703
rect 390 698 396 699
rect 410 703 416 704
rect 410 699 411 703
rect 415 699 416 703
rect 410 698 416 699
rect 310 692 316 693
rect 310 688 311 692
rect 315 688 316 692
rect 310 687 316 688
rect 382 692 388 693
rect 382 688 383 692
rect 387 688 388 692
rect 382 687 388 688
rect 412 680 414 698
rect 456 693 458 705
rect 482 703 488 704
rect 482 699 483 703
rect 487 699 488 703
rect 482 698 488 699
rect 454 692 460 693
rect 454 688 455 692
rect 459 688 460 692
rect 454 687 460 688
rect 484 680 486 698
rect 520 693 522 705
rect 584 693 586 705
rect 518 692 524 693
rect 518 688 519 692
rect 523 688 524 692
rect 518 687 524 688
rect 582 692 588 693
rect 582 688 583 692
rect 587 688 588 692
rect 582 687 588 688
rect 608 680 610 714
rect 640 711 642 727
rect 680 720 682 738
rect 686 732 692 733
rect 686 728 687 732
rect 691 728 692 732
rect 686 727 692 728
rect 678 719 684 720
rect 678 715 679 719
rect 683 715 684 719
rect 678 714 684 715
rect 688 711 690 727
rect 728 712 730 738
rect 742 732 748 733
rect 742 728 743 732
rect 747 728 748 732
rect 742 727 748 728
rect 798 732 804 733
rect 798 728 799 732
rect 803 728 804 732
rect 798 727 804 728
rect 726 711 732 712
rect 744 711 746 727
rect 790 719 796 720
rect 790 715 791 719
rect 795 715 796 719
rect 790 714 796 715
rect 639 710 643 711
rect 639 705 643 706
rect 647 710 651 711
rect 647 705 651 706
rect 687 710 691 711
rect 687 705 691 706
rect 711 710 715 711
rect 726 707 727 711
rect 731 707 732 711
rect 726 706 732 707
rect 743 710 747 711
rect 711 705 715 706
rect 743 705 747 706
rect 767 710 771 711
rect 767 705 771 706
rect 630 703 636 704
rect 630 699 631 703
rect 635 699 636 703
rect 630 698 636 699
rect 632 680 634 698
rect 648 693 650 705
rect 654 703 660 704
rect 654 699 655 703
rect 659 699 660 703
rect 654 698 660 699
rect 646 692 652 693
rect 646 688 647 692
rect 651 688 652 692
rect 646 687 652 688
rect 274 679 280 680
rect 274 675 275 679
rect 279 675 280 679
rect 274 674 280 675
rect 282 679 288 680
rect 282 675 283 679
rect 287 675 288 679
rect 282 674 288 675
rect 410 679 416 680
rect 410 675 411 679
rect 415 675 416 679
rect 410 674 416 675
rect 482 679 488 680
rect 482 675 483 679
rect 487 675 488 679
rect 482 674 488 675
rect 534 679 540 680
rect 534 675 535 679
rect 539 675 540 679
rect 534 674 540 675
rect 606 679 612 680
rect 606 675 607 679
rect 611 675 612 679
rect 606 674 612 675
rect 630 679 636 680
rect 630 675 631 679
rect 635 675 636 679
rect 630 674 636 675
rect 246 664 252 665
rect 246 660 247 664
rect 251 660 252 664
rect 246 659 252 660
rect 248 651 250 659
rect 247 650 251 651
rect 247 645 251 646
rect 206 627 212 628
rect 110 624 116 625
rect 110 620 111 624
rect 115 620 116 624
rect 206 623 207 627
rect 211 623 212 627
rect 206 622 212 623
rect 234 627 240 628
rect 234 623 235 627
rect 239 623 240 627
rect 234 622 240 623
rect 262 627 268 628
rect 262 623 263 627
rect 267 623 268 627
rect 262 622 268 623
rect 110 619 116 620
rect 112 595 114 619
rect 158 616 164 617
rect 158 612 159 616
rect 163 612 164 616
rect 158 611 164 612
rect 160 595 162 611
rect 208 604 210 622
rect 214 616 220 617
rect 214 612 215 616
rect 219 612 220 616
rect 214 611 220 612
rect 182 603 188 604
rect 182 599 183 603
rect 187 599 188 603
rect 182 598 188 599
rect 206 603 212 604
rect 206 599 207 603
rect 211 599 212 603
rect 206 598 212 599
rect 111 594 115 595
rect 111 589 115 590
rect 159 594 163 595
rect 159 589 163 590
rect 112 569 114 589
rect 160 577 162 589
rect 158 576 164 577
rect 158 572 159 576
rect 163 572 164 576
rect 158 571 164 572
rect 110 568 116 569
rect 110 564 111 568
rect 115 564 116 568
rect 184 564 186 598
rect 216 595 218 611
rect 207 594 211 595
rect 207 589 211 590
rect 215 594 219 595
rect 215 589 219 590
rect 255 594 259 595
rect 255 589 259 590
rect 208 577 210 589
rect 242 587 248 588
rect 242 583 243 587
rect 247 583 248 587
rect 242 582 248 583
rect 206 576 212 577
rect 206 572 207 576
rect 211 572 212 576
rect 206 571 212 572
rect 244 564 246 582
rect 256 577 258 589
rect 264 588 266 622
rect 276 604 278 674
rect 310 664 316 665
rect 310 660 311 664
rect 315 660 316 664
rect 310 659 316 660
rect 382 664 388 665
rect 382 660 383 664
rect 387 660 388 664
rect 382 659 388 660
rect 454 664 460 665
rect 454 660 455 664
rect 459 660 460 664
rect 454 659 460 660
rect 518 664 524 665
rect 518 660 519 664
rect 523 660 524 664
rect 518 659 524 660
rect 312 651 314 659
rect 384 651 386 659
rect 456 651 458 659
rect 520 651 522 659
rect 287 650 291 651
rect 287 645 291 646
rect 311 650 315 651
rect 311 645 315 646
rect 367 650 371 651
rect 367 645 371 646
rect 383 650 387 651
rect 383 645 387 646
rect 455 650 459 651
rect 455 645 459 646
rect 519 650 523 651
rect 519 645 523 646
rect 286 644 292 645
rect 286 640 287 644
rect 291 640 292 644
rect 286 639 292 640
rect 366 644 372 645
rect 366 640 367 644
rect 371 640 372 644
rect 366 639 372 640
rect 454 644 460 645
rect 454 640 455 644
rect 459 640 460 644
rect 454 639 460 640
rect 390 627 396 628
rect 390 623 391 627
rect 395 623 396 627
rect 390 622 396 623
rect 402 627 408 628
rect 402 623 403 627
rect 407 623 408 627
rect 402 622 408 623
rect 286 616 292 617
rect 286 612 287 616
rect 291 612 292 616
rect 286 611 292 612
rect 366 616 372 617
rect 366 612 367 616
rect 371 612 372 616
rect 366 611 372 612
rect 274 603 280 604
rect 274 599 275 603
rect 279 599 280 603
rect 274 598 280 599
rect 288 595 290 611
rect 334 595 340 596
rect 368 595 370 611
rect 287 594 291 595
rect 287 589 291 590
rect 311 594 315 595
rect 334 591 335 595
rect 339 591 340 595
rect 334 590 340 591
rect 367 594 371 595
rect 311 589 315 590
rect 262 587 268 588
rect 262 583 263 587
rect 267 583 268 587
rect 262 582 268 583
rect 312 577 314 589
rect 254 576 260 577
rect 254 572 255 576
rect 259 572 260 576
rect 254 571 260 572
rect 310 576 316 577
rect 310 572 311 576
rect 315 572 316 576
rect 310 571 316 572
rect 336 564 338 590
rect 367 589 371 590
rect 383 594 387 595
rect 383 589 387 590
rect 370 583 376 584
rect 370 579 371 583
rect 375 579 376 583
rect 370 578 376 579
rect 110 563 116 564
rect 182 563 188 564
rect 182 559 183 563
rect 187 559 188 563
rect 182 558 188 559
rect 230 563 236 564
rect 230 559 231 563
rect 235 559 236 563
rect 230 558 236 559
rect 242 563 248 564
rect 242 559 243 563
rect 247 559 248 563
rect 242 558 248 559
rect 334 563 340 564
rect 334 559 335 563
rect 339 559 340 563
rect 334 558 340 559
rect 110 551 116 552
rect 110 547 111 551
rect 115 547 116 551
rect 110 546 116 547
rect 158 548 164 549
rect 112 535 114 546
rect 158 544 159 548
rect 163 544 164 548
rect 158 543 164 544
rect 206 548 212 549
rect 206 544 207 548
rect 211 544 212 548
rect 206 543 212 544
rect 160 535 162 543
rect 208 535 210 543
rect 111 534 115 535
rect 111 529 115 530
rect 159 534 163 535
rect 159 529 163 530
rect 167 534 171 535
rect 167 529 171 530
rect 207 534 211 535
rect 207 529 211 530
rect 223 534 227 535
rect 223 529 227 530
rect 112 526 114 529
rect 166 528 172 529
rect 110 525 116 526
rect 110 521 111 525
rect 115 521 116 525
rect 166 524 167 528
rect 171 524 172 528
rect 166 523 172 524
rect 222 528 228 529
rect 222 524 223 528
rect 227 524 228 528
rect 222 523 228 524
rect 110 520 116 521
rect 174 511 180 512
rect 110 508 116 509
rect 110 504 111 508
rect 115 504 116 508
rect 174 507 175 511
rect 179 507 180 511
rect 174 506 180 507
rect 110 503 116 504
rect 112 483 114 503
rect 166 500 172 501
rect 166 496 167 500
rect 171 496 172 500
rect 166 495 172 496
rect 168 483 170 495
rect 111 482 115 483
rect 111 477 115 478
rect 167 482 171 483
rect 167 477 171 478
rect 112 457 114 477
rect 168 465 170 477
rect 176 476 178 506
rect 222 500 228 501
rect 222 496 223 500
rect 227 496 228 500
rect 222 495 228 496
rect 224 483 226 495
rect 232 492 234 558
rect 254 548 260 549
rect 254 544 255 548
rect 259 544 260 548
rect 254 543 260 544
rect 310 548 316 549
rect 310 544 311 548
rect 315 544 316 548
rect 310 543 316 544
rect 256 535 258 543
rect 312 535 314 543
rect 255 534 259 535
rect 255 529 259 530
rect 287 534 291 535
rect 287 529 291 530
rect 311 534 315 535
rect 311 529 315 530
rect 359 534 363 535
rect 359 529 363 530
rect 286 528 292 529
rect 286 524 287 528
rect 291 524 292 528
rect 286 523 292 524
rect 358 528 364 529
rect 358 524 359 528
rect 363 524 364 528
rect 358 523 364 524
rect 372 512 374 578
rect 384 577 386 589
rect 392 588 394 622
rect 404 604 406 622
rect 454 616 460 617
rect 454 612 455 616
rect 459 612 460 616
rect 454 611 460 612
rect 402 603 408 604
rect 402 599 403 603
rect 407 599 408 603
rect 402 598 408 599
rect 456 595 458 611
rect 536 604 538 674
rect 582 664 588 665
rect 582 660 583 664
rect 587 660 588 664
rect 582 659 588 660
rect 646 664 652 665
rect 646 660 647 664
rect 651 660 652 664
rect 646 659 652 660
rect 584 651 586 659
rect 648 651 650 659
rect 543 650 547 651
rect 543 645 547 646
rect 583 650 587 651
rect 583 645 587 646
rect 631 650 635 651
rect 631 645 635 646
rect 647 650 651 651
rect 647 645 651 646
rect 542 644 548 645
rect 542 640 543 644
rect 547 640 548 644
rect 542 639 548 640
rect 630 644 636 645
rect 630 640 631 644
rect 635 640 636 644
rect 630 639 636 640
rect 656 628 658 698
rect 712 693 714 705
rect 734 703 740 704
rect 734 699 735 703
rect 739 699 740 703
rect 734 698 740 699
rect 710 692 716 693
rect 710 688 711 692
rect 715 688 716 692
rect 710 687 716 688
rect 736 685 738 698
rect 768 693 770 705
rect 766 692 772 693
rect 766 688 767 692
rect 771 688 772 692
rect 766 687 772 688
rect 735 684 739 685
rect 792 680 794 714
rect 800 711 802 727
rect 848 720 850 738
rect 854 732 860 733
rect 854 728 855 732
rect 859 728 860 732
rect 854 727 860 728
rect 846 719 852 720
rect 846 715 847 719
rect 851 715 852 719
rect 846 714 852 715
rect 856 711 858 727
rect 864 712 866 738
rect 1094 736 1095 740
rect 1099 736 1100 740
rect 1094 735 1100 736
rect 862 711 868 712
rect 1096 711 1098 735
rect 1186 731 1192 732
rect 1134 728 1140 729
rect 1134 724 1135 728
rect 1139 724 1140 728
rect 1186 727 1187 731
rect 1191 727 1192 731
rect 1186 726 1192 727
rect 1226 731 1232 732
rect 1226 727 1227 731
rect 1231 727 1232 731
rect 1226 726 1232 727
rect 1278 731 1284 732
rect 1278 727 1279 731
rect 1283 727 1284 731
rect 1278 726 1284 727
rect 1134 723 1140 724
rect 799 710 803 711
rect 799 705 803 706
rect 823 710 827 711
rect 823 705 827 706
rect 855 710 859 711
rect 862 707 863 711
rect 867 707 868 711
rect 862 706 868 707
rect 879 710 883 711
rect 855 705 859 706
rect 879 705 883 706
rect 943 710 947 711
rect 943 705 947 706
rect 1095 710 1099 711
rect 1095 705 1099 706
rect 814 703 820 704
rect 814 699 815 703
rect 819 699 820 703
rect 814 698 820 699
rect 735 679 739 680
rect 790 679 796 680
rect 790 675 791 679
rect 795 675 796 679
rect 790 674 796 675
rect 710 664 716 665
rect 710 660 711 664
rect 715 660 716 664
rect 710 659 716 660
rect 766 664 772 665
rect 766 660 767 664
rect 771 660 772 664
rect 766 659 772 660
rect 712 651 714 659
rect 768 651 770 659
rect 711 650 715 651
rect 711 645 715 646
rect 719 650 723 651
rect 719 645 723 646
rect 767 650 771 651
rect 767 645 771 646
rect 799 650 803 651
rect 799 645 803 646
rect 718 644 724 645
rect 718 640 719 644
rect 723 640 724 644
rect 718 639 724 640
rect 798 644 804 645
rect 798 640 799 644
rect 803 640 804 644
rect 798 639 804 640
rect 816 628 818 698
rect 824 693 826 705
rect 880 693 882 705
rect 906 703 912 704
rect 906 699 907 703
rect 911 699 912 703
rect 906 698 912 699
rect 822 692 828 693
rect 822 688 823 692
rect 827 688 828 692
rect 822 687 828 688
rect 878 692 884 693
rect 878 688 879 692
rect 883 688 884 692
rect 878 687 884 688
rect 908 680 910 698
rect 944 693 946 705
rect 942 692 948 693
rect 942 688 943 692
rect 947 688 948 692
rect 942 687 948 688
rect 1096 685 1098 705
rect 1136 699 1138 723
rect 1158 720 1164 721
rect 1158 716 1159 720
rect 1163 716 1164 720
rect 1158 715 1164 716
rect 1160 699 1162 715
rect 1188 708 1190 726
rect 1198 720 1204 721
rect 1198 716 1199 720
rect 1203 716 1204 720
rect 1198 715 1204 716
rect 1186 707 1192 708
rect 1186 703 1187 707
rect 1191 703 1192 707
rect 1186 702 1192 703
rect 1200 699 1202 715
rect 1228 708 1230 726
rect 1238 720 1244 721
rect 1238 716 1239 720
rect 1243 716 1244 720
rect 1238 715 1244 716
rect 1226 707 1232 708
rect 1226 703 1227 707
rect 1231 703 1232 707
rect 1226 702 1232 703
rect 1240 699 1242 715
rect 1280 708 1282 726
rect 1286 720 1292 721
rect 1286 716 1287 720
rect 1291 716 1292 720
rect 1286 715 1292 716
rect 1278 707 1284 708
rect 1278 703 1279 707
rect 1283 703 1284 707
rect 1278 702 1284 703
rect 1288 699 1290 715
rect 1312 700 1314 770
rect 1342 760 1348 761
rect 1342 756 1343 760
rect 1347 756 1348 760
rect 1342 755 1348 756
rect 1446 760 1452 761
rect 1446 756 1447 760
rect 1451 756 1452 760
rect 1446 755 1452 756
rect 1343 754 1347 755
rect 1343 749 1347 750
rect 1359 754 1363 755
rect 1359 749 1363 750
rect 1439 754 1443 755
rect 1439 749 1443 750
rect 1447 754 1451 755
rect 1447 749 1451 750
rect 1358 748 1364 749
rect 1358 744 1359 748
rect 1363 744 1364 748
rect 1358 743 1364 744
rect 1438 748 1444 749
rect 1438 744 1439 748
rect 1443 744 1444 748
rect 1438 743 1444 744
rect 1342 739 1348 740
rect 1342 735 1343 739
rect 1347 735 1348 739
rect 1342 734 1348 735
rect 1310 699 1316 700
rect 1135 698 1139 699
rect 1135 693 1139 694
rect 1159 698 1163 699
rect 1159 693 1163 694
rect 1199 698 1203 699
rect 1199 693 1203 694
rect 1239 698 1243 699
rect 1239 693 1243 694
rect 1287 698 1291 699
rect 1310 695 1311 699
rect 1315 695 1316 699
rect 1310 694 1316 695
rect 1335 698 1339 699
rect 1287 693 1291 694
rect 1335 693 1339 694
rect 967 684 971 685
rect 1094 684 1100 685
rect 1094 680 1095 684
rect 1099 680 1100 684
rect 906 679 912 680
rect 906 675 907 679
rect 911 675 912 679
rect 906 674 912 675
rect 966 679 972 680
rect 1094 679 1100 680
rect 966 675 967 679
rect 971 675 972 679
rect 966 674 972 675
rect 1136 673 1138 693
rect 1240 681 1242 693
rect 1274 691 1280 692
rect 1274 687 1275 691
rect 1279 687 1280 691
rect 1274 686 1280 687
rect 1238 680 1244 681
rect 1238 676 1239 680
rect 1243 676 1244 680
rect 1238 675 1244 676
rect 1134 672 1140 673
rect 1134 668 1135 672
rect 1139 668 1140 672
rect 1276 668 1278 686
rect 1288 681 1290 693
rect 1322 691 1328 692
rect 1322 687 1323 691
rect 1327 687 1328 691
rect 1322 686 1328 687
rect 1286 680 1292 681
rect 1286 676 1287 680
rect 1291 676 1292 680
rect 1286 675 1292 676
rect 1324 668 1326 686
rect 1336 681 1338 693
rect 1344 692 1346 734
rect 1350 731 1356 732
rect 1350 727 1351 731
rect 1355 727 1356 731
rect 1350 726 1356 727
rect 1430 731 1436 732
rect 1430 727 1431 731
rect 1435 727 1436 731
rect 1430 726 1436 727
rect 1352 708 1354 726
rect 1358 720 1364 721
rect 1358 716 1359 720
rect 1363 716 1364 720
rect 1358 715 1364 716
rect 1350 707 1356 708
rect 1350 703 1351 707
rect 1355 703 1356 707
rect 1350 702 1356 703
rect 1360 699 1362 715
rect 1432 708 1434 726
rect 1438 720 1444 721
rect 1438 716 1439 720
rect 1443 716 1444 720
rect 1438 715 1444 716
rect 1430 707 1436 708
rect 1430 703 1431 707
rect 1435 703 1436 707
rect 1430 702 1436 703
rect 1440 699 1442 715
rect 1520 708 1522 770
rect 1550 760 1556 761
rect 1550 756 1551 760
rect 1555 756 1556 760
rect 1550 755 1556 756
rect 1654 760 1660 761
rect 1654 756 1655 760
rect 1659 756 1660 760
rect 1654 755 1660 756
rect 1750 760 1756 761
rect 1750 756 1751 760
rect 1755 756 1756 760
rect 1750 755 1756 756
rect 1527 754 1531 755
rect 1527 749 1531 750
rect 1551 754 1555 755
rect 1551 749 1555 750
rect 1615 754 1619 755
rect 1615 749 1619 750
rect 1655 754 1659 755
rect 1655 749 1659 750
rect 1711 754 1715 755
rect 1711 749 1715 750
rect 1751 754 1755 755
rect 1751 749 1755 750
rect 1807 754 1811 755
rect 1807 749 1811 750
rect 1526 748 1532 749
rect 1526 744 1527 748
rect 1531 744 1532 748
rect 1526 743 1532 744
rect 1614 748 1620 749
rect 1614 744 1615 748
rect 1619 744 1620 748
rect 1614 743 1620 744
rect 1710 748 1716 749
rect 1710 744 1711 748
rect 1715 744 1716 748
rect 1710 743 1716 744
rect 1806 748 1812 749
rect 1806 744 1807 748
rect 1811 744 1812 748
rect 1806 743 1812 744
rect 1832 732 1834 794
rect 1840 789 1842 801
rect 1866 799 1872 800
rect 1866 795 1867 799
rect 1871 795 1872 799
rect 1866 794 1872 795
rect 1838 788 1844 789
rect 1838 784 1839 788
rect 1843 784 1844 788
rect 1838 783 1844 784
rect 1868 776 1870 794
rect 1920 789 1922 801
rect 1946 799 1952 800
rect 1946 795 1947 799
rect 1951 795 1952 799
rect 1946 794 1952 795
rect 1918 788 1924 789
rect 1918 784 1919 788
rect 1923 784 1924 788
rect 1918 783 1924 784
rect 1948 776 1950 794
rect 2000 776 2002 814
rect 2016 807 2018 827
rect 2064 820 2066 838
rect 2070 832 2076 833
rect 2070 828 2071 832
rect 2075 828 2076 832
rect 2070 827 2076 828
rect 2062 819 2068 820
rect 2062 815 2063 819
rect 2067 815 2068 819
rect 2062 814 2068 815
rect 2072 807 2074 827
rect 2007 806 2011 807
rect 2007 801 2011 802
rect 2015 806 2019 807
rect 2015 801 2019 802
rect 2071 806 2075 807
rect 2071 801 2075 802
rect 2008 789 2010 801
rect 2072 789 2074 801
rect 2080 800 2082 838
rect 2118 836 2119 840
rect 2123 836 2124 840
rect 2118 835 2124 836
rect 2120 807 2122 835
rect 2119 806 2123 807
rect 2119 801 2123 802
rect 2078 799 2084 800
rect 2078 795 2079 799
rect 2083 795 2084 799
rect 2078 794 2084 795
rect 2006 788 2012 789
rect 2006 784 2007 788
rect 2011 784 2012 788
rect 2006 783 2012 784
rect 2070 788 2076 789
rect 2070 784 2071 788
rect 2075 784 2076 788
rect 2070 783 2076 784
rect 2120 781 2122 801
rect 2118 780 2124 781
rect 2118 776 2119 780
rect 2123 776 2124 780
rect 1866 775 1872 776
rect 1866 771 1867 775
rect 1871 771 1872 775
rect 1866 770 1872 771
rect 1946 775 1952 776
rect 1946 771 1947 775
rect 1951 771 1952 775
rect 1946 770 1952 771
rect 1998 775 2004 776
rect 1998 771 1999 775
rect 2003 771 2004 775
rect 1998 770 2004 771
rect 2086 775 2092 776
rect 2118 775 2124 776
rect 2086 771 2087 775
rect 2091 771 2092 775
rect 2086 770 2092 771
rect 1838 760 1844 761
rect 1838 756 1839 760
rect 1843 756 1844 760
rect 1838 755 1844 756
rect 1918 760 1924 761
rect 1918 756 1919 760
rect 1923 756 1924 760
rect 1918 755 1924 756
rect 2006 760 2012 761
rect 2006 756 2007 760
rect 2011 756 2012 760
rect 2006 755 2012 756
rect 2070 760 2076 761
rect 2070 756 2071 760
rect 2075 756 2076 760
rect 2070 755 2076 756
rect 1839 754 1843 755
rect 1839 749 1843 750
rect 1903 754 1907 755
rect 1903 749 1907 750
rect 1919 754 1923 755
rect 1919 749 1923 750
rect 1999 754 2003 755
rect 1999 749 2003 750
rect 2007 754 2011 755
rect 2007 749 2011 750
rect 2071 754 2075 755
rect 2071 749 2075 750
rect 1902 748 1908 749
rect 1902 744 1903 748
rect 1907 744 1908 748
rect 1902 743 1908 744
rect 1998 748 2004 749
rect 1998 744 1999 748
rect 2003 744 2004 748
rect 1998 743 2004 744
rect 2070 748 2076 749
rect 2070 744 2071 748
rect 2075 744 2076 748
rect 2070 743 2076 744
rect 1606 731 1612 732
rect 1606 727 1607 731
rect 1611 727 1612 731
rect 1606 726 1612 727
rect 1702 731 1708 732
rect 1702 727 1703 731
rect 1707 727 1708 731
rect 1702 726 1708 727
rect 1718 731 1724 732
rect 1718 727 1719 731
rect 1723 727 1724 731
rect 1718 726 1724 727
rect 1830 731 1836 732
rect 1830 727 1831 731
rect 1835 727 1836 731
rect 1830 726 1836 727
rect 2078 731 2084 732
rect 2078 727 2079 731
rect 2083 727 2084 731
rect 2078 726 2084 727
rect 1526 720 1532 721
rect 1526 716 1527 720
rect 1531 716 1532 720
rect 1526 715 1532 716
rect 1518 707 1524 708
rect 1518 703 1519 707
rect 1523 703 1524 707
rect 1518 702 1524 703
rect 1528 699 1530 715
rect 1608 708 1610 726
rect 1614 720 1620 721
rect 1614 716 1615 720
rect 1619 716 1620 720
rect 1614 715 1620 716
rect 1606 707 1612 708
rect 1606 703 1607 707
rect 1611 703 1612 707
rect 1606 702 1612 703
rect 1534 699 1540 700
rect 1616 699 1618 715
rect 1704 708 1706 726
rect 1710 720 1716 721
rect 1710 716 1711 720
rect 1715 716 1716 720
rect 1710 715 1716 716
rect 1702 707 1708 708
rect 1702 703 1703 707
rect 1707 703 1708 707
rect 1702 702 1708 703
rect 1712 699 1714 715
rect 1720 700 1722 726
rect 1806 720 1812 721
rect 1806 716 1807 720
rect 1811 716 1812 720
rect 1806 715 1812 716
rect 1902 720 1908 721
rect 1902 716 1903 720
rect 1907 716 1908 720
rect 1902 715 1908 716
rect 1998 720 2004 721
rect 1998 716 1999 720
rect 2003 716 2004 720
rect 1998 715 2004 716
rect 2070 720 2076 721
rect 2070 716 2071 720
rect 2075 716 2076 720
rect 2070 715 2076 716
rect 1718 699 1724 700
rect 1808 699 1810 715
rect 1904 699 1906 715
rect 1986 707 1992 708
rect 1986 703 1987 707
rect 1991 703 1992 707
rect 1986 702 1992 703
rect 1359 698 1363 699
rect 1359 693 1363 694
rect 1391 698 1395 699
rect 1391 693 1395 694
rect 1439 698 1443 699
rect 1439 693 1443 694
rect 1447 698 1451 699
rect 1447 693 1451 694
rect 1511 698 1515 699
rect 1511 693 1515 694
rect 1527 698 1531 699
rect 1534 695 1535 699
rect 1539 695 1540 699
rect 1534 694 1540 695
rect 1575 698 1579 699
rect 1527 693 1531 694
rect 1342 691 1348 692
rect 1342 687 1343 691
rect 1347 687 1348 691
rect 1342 686 1348 687
rect 1392 681 1394 693
rect 1448 681 1450 693
rect 1512 681 1514 693
rect 1334 680 1340 681
rect 1334 676 1335 680
rect 1339 676 1340 680
rect 1334 675 1340 676
rect 1390 680 1396 681
rect 1390 676 1391 680
rect 1395 676 1396 680
rect 1390 675 1396 676
rect 1446 680 1452 681
rect 1446 676 1447 680
rect 1451 676 1452 680
rect 1446 675 1452 676
rect 1510 680 1516 681
rect 1510 676 1511 680
rect 1515 676 1516 680
rect 1510 675 1516 676
rect 1536 668 1538 694
rect 1575 693 1579 694
rect 1615 698 1619 699
rect 1615 693 1619 694
rect 1639 698 1643 699
rect 1639 693 1643 694
rect 1703 698 1707 699
rect 1703 693 1707 694
rect 1711 698 1715 699
rect 1718 695 1719 699
rect 1723 695 1724 699
rect 1718 694 1724 695
rect 1767 698 1771 699
rect 1711 693 1715 694
rect 1767 693 1771 694
rect 1807 698 1811 699
rect 1807 693 1811 694
rect 1831 698 1835 699
rect 1831 693 1835 694
rect 1895 698 1899 699
rect 1895 693 1899 694
rect 1903 698 1907 699
rect 1903 693 1907 694
rect 1959 698 1963 699
rect 1959 693 1963 694
rect 1562 691 1568 692
rect 1562 687 1563 691
rect 1567 687 1568 691
rect 1562 686 1568 687
rect 1564 668 1566 686
rect 1576 681 1578 693
rect 1626 691 1632 692
rect 1626 687 1627 691
rect 1631 687 1632 691
rect 1626 686 1632 687
rect 1574 680 1580 681
rect 1574 676 1575 680
rect 1579 676 1580 680
rect 1574 675 1580 676
rect 1628 668 1630 686
rect 1640 681 1642 693
rect 1704 681 1706 693
rect 1730 691 1736 692
rect 1710 687 1716 688
rect 1710 683 1711 687
rect 1715 683 1716 687
rect 1730 687 1731 691
rect 1735 687 1736 691
rect 1730 686 1736 687
rect 1710 682 1716 683
rect 1638 680 1644 681
rect 1638 676 1639 680
rect 1643 676 1644 680
rect 1638 675 1644 676
rect 1702 680 1708 681
rect 1702 676 1703 680
rect 1707 676 1708 680
rect 1702 675 1708 676
rect 1094 667 1100 668
rect 1134 667 1140 668
rect 1266 667 1272 668
rect 822 664 828 665
rect 822 660 823 664
rect 827 660 828 664
rect 822 659 828 660
rect 878 664 884 665
rect 878 660 879 664
rect 883 660 884 664
rect 878 659 884 660
rect 942 664 948 665
rect 942 660 943 664
rect 947 660 948 664
rect 1094 663 1095 667
rect 1099 663 1100 667
rect 1094 662 1100 663
rect 1266 663 1267 667
rect 1271 663 1272 667
rect 1266 662 1272 663
rect 1274 667 1280 668
rect 1274 663 1275 667
rect 1279 663 1280 667
rect 1274 662 1280 663
rect 1322 667 1328 668
rect 1322 663 1323 667
rect 1327 663 1328 667
rect 1322 662 1328 663
rect 1470 667 1476 668
rect 1470 663 1471 667
rect 1475 663 1476 667
rect 1470 662 1476 663
rect 1534 667 1540 668
rect 1534 663 1535 667
rect 1539 663 1540 667
rect 1534 662 1540 663
rect 1562 667 1568 668
rect 1562 663 1563 667
rect 1567 663 1568 667
rect 1562 662 1568 663
rect 1626 667 1632 668
rect 1626 663 1627 667
rect 1631 663 1632 667
rect 1626 662 1632 663
rect 942 659 948 660
rect 824 651 826 659
rect 880 651 882 659
rect 944 651 946 659
rect 1096 651 1098 662
rect 1134 655 1140 656
rect 1134 651 1135 655
rect 1139 651 1140 655
rect 823 650 827 651
rect 823 645 827 646
rect 871 650 875 651
rect 871 645 875 646
rect 879 650 883 651
rect 879 645 883 646
rect 943 650 947 651
rect 943 645 947 646
rect 951 650 955 651
rect 951 645 955 646
rect 1031 650 1035 651
rect 1031 645 1035 646
rect 1095 650 1099 651
rect 1134 650 1140 651
rect 1238 652 1244 653
rect 1136 647 1138 650
rect 1238 648 1239 652
rect 1243 648 1244 652
rect 1238 647 1244 648
rect 1095 645 1099 646
rect 1135 646 1139 647
rect 870 644 876 645
rect 870 640 871 644
rect 875 640 876 644
rect 870 639 876 640
rect 950 644 956 645
rect 950 640 951 644
rect 955 640 956 644
rect 950 639 956 640
rect 1030 644 1036 645
rect 1030 640 1031 644
rect 1035 640 1036 644
rect 1096 642 1098 645
rect 1030 639 1036 640
rect 1094 641 1100 642
rect 1135 641 1139 642
rect 1239 646 1243 647
rect 1239 641 1243 642
rect 1094 637 1095 641
rect 1099 637 1100 641
rect 1136 638 1138 641
rect 1094 636 1100 637
rect 1134 637 1140 638
rect 1134 633 1135 637
rect 1139 633 1140 637
rect 1134 632 1140 633
rect 654 627 660 628
rect 654 623 655 627
rect 659 623 660 627
rect 654 622 660 623
rect 790 627 796 628
rect 790 623 791 627
rect 795 623 796 627
rect 790 622 796 623
rect 814 627 820 628
rect 814 623 815 627
rect 819 623 820 627
rect 814 622 820 623
rect 942 627 948 628
rect 942 623 943 627
rect 947 623 948 627
rect 942 622 948 623
rect 1022 627 1028 628
rect 1022 623 1023 627
rect 1027 623 1028 627
rect 1022 622 1028 623
rect 1038 627 1044 628
rect 1038 623 1039 627
rect 1043 623 1044 627
rect 1038 622 1044 623
rect 1094 624 1100 625
rect 542 616 548 617
rect 542 612 543 616
rect 547 612 548 616
rect 542 611 548 612
rect 630 616 636 617
rect 630 612 631 616
rect 635 612 636 616
rect 630 611 636 612
rect 718 616 724 617
rect 718 612 719 616
rect 723 612 724 616
rect 718 611 724 612
rect 727 612 731 613
rect 534 603 540 604
rect 534 599 535 603
rect 539 599 540 603
rect 534 598 540 599
rect 544 595 546 611
rect 632 595 634 611
rect 646 603 652 604
rect 646 599 647 603
rect 651 599 652 603
rect 646 598 652 599
rect 455 594 459 595
rect 455 589 459 590
rect 463 594 467 595
rect 463 589 467 590
rect 543 594 547 595
rect 543 589 547 590
rect 623 594 627 595
rect 623 589 627 590
rect 631 594 635 595
rect 631 589 635 590
rect 390 587 396 588
rect 390 583 391 587
rect 395 583 396 587
rect 390 582 396 583
rect 410 587 416 588
rect 410 583 411 587
rect 415 583 416 587
rect 410 582 416 583
rect 382 576 388 577
rect 382 572 383 576
rect 387 572 388 576
rect 382 571 388 572
rect 412 564 414 582
rect 464 577 466 589
rect 490 587 496 588
rect 490 583 491 587
rect 495 583 496 587
rect 490 582 496 583
rect 462 576 468 577
rect 462 572 463 576
rect 467 572 468 576
rect 462 571 468 572
rect 492 564 494 582
rect 544 577 546 589
rect 624 577 626 589
rect 542 576 548 577
rect 542 572 543 576
rect 547 572 548 576
rect 542 571 548 572
rect 622 576 628 577
rect 622 572 623 576
rect 627 572 628 576
rect 622 571 628 572
rect 648 564 650 598
rect 720 595 722 611
rect 727 607 731 608
rect 728 604 730 607
rect 792 604 794 622
rect 798 616 804 617
rect 798 612 799 616
rect 803 612 804 616
rect 798 611 804 612
rect 870 616 876 617
rect 870 612 871 616
rect 875 612 876 616
rect 870 611 876 612
rect 726 603 732 604
rect 726 599 727 603
rect 731 599 732 603
rect 726 598 732 599
rect 790 603 796 604
rect 790 599 791 603
rect 795 599 796 603
rect 790 598 796 599
rect 800 595 802 611
rect 872 595 874 611
rect 944 604 946 622
rect 950 616 956 617
rect 950 612 951 616
rect 955 612 956 616
rect 950 611 956 612
rect 878 603 884 604
rect 878 599 879 603
rect 883 599 884 603
rect 878 598 884 599
rect 942 603 948 604
rect 942 599 943 603
rect 947 599 948 603
rect 942 598 948 599
rect 703 594 707 595
rect 703 589 707 590
rect 719 594 723 595
rect 719 589 723 590
rect 783 594 787 595
rect 783 589 787 590
rect 799 594 803 595
rect 799 589 803 590
rect 855 594 859 595
rect 855 589 859 590
rect 871 594 875 595
rect 871 589 875 590
rect 682 587 688 588
rect 682 583 683 587
rect 687 583 688 587
rect 682 582 688 583
rect 690 587 696 588
rect 690 583 691 587
rect 695 583 696 587
rect 690 582 696 583
rect 684 564 686 582
rect 410 563 416 564
rect 410 559 411 563
rect 415 559 416 563
rect 410 558 416 559
rect 490 563 496 564
rect 490 559 491 563
rect 495 559 496 563
rect 490 558 496 559
rect 582 563 588 564
rect 582 559 583 563
rect 587 559 588 563
rect 582 558 588 559
rect 646 563 652 564
rect 646 559 647 563
rect 651 559 652 563
rect 646 558 652 559
rect 682 563 688 564
rect 682 559 683 563
rect 687 559 688 563
rect 682 558 688 559
rect 382 548 388 549
rect 382 544 383 548
rect 387 544 388 548
rect 382 543 388 544
rect 462 548 468 549
rect 462 544 463 548
rect 467 544 468 548
rect 462 543 468 544
rect 542 548 548 549
rect 542 544 543 548
rect 547 544 548 548
rect 542 543 548 544
rect 384 535 386 543
rect 464 535 466 543
rect 544 535 546 543
rect 383 534 387 535
rect 383 529 387 530
rect 431 534 435 535
rect 431 529 435 530
rect 463 534 467 535
rect 463 529 467 530
rect 511 534 515 535
rect 511 529 515 530
rect 543 534 547 535
rect 543 529 547 530
rect 430 528 436 529
rect 430 524 431 528
rect 435 524 436 528
rect 430 523 436 524
rect 510 528 516 529
rect 510 524 511 528
rect 515 524 516 528
rect 510 523 516 524
rect 350 511 356 512
rect 350 507 351 511
rect 355 507 356 511
rect 350 506 356 507
rect 370 511 376 512
rect 370 507 371 511
rect 375 507 376 511
rect 370 506 376 507
rect 394 511 400 512
rect 394 507 395 511
rect 399 507 400 511
rect 394 506 400 507
rect 546 511 552 512
rect 546 507 547 511
rect 551 507 552 511
rect 546 506 552 507
rect 286 500 292 501
rect 286 496 287 500
rect 291 496 292 500
rect 286 495 292 496
rect 230 491 236 492
rect 230 487 231 491
rect 235 487 236 491
rect 230 486 236 487
rect 258 487 264 488
rect 258 483 259 487
rect 263 483 264 487
rect 288 483 290 495
rect 352 488 354 506
rect 358 500 364 501
rect 358 496 359 500
rect 363 496 364 500
rect 358 495 364 496
rect 350 487 356 488
rect 350 483 351 487
rect 355 483 356 487
rect 360 483 362 495
rect 223 482 227 483
rect 223 477 227 478
rect 231 482 235 483
rect 258 482 264 483
rect 287 482 291 483
rect 231 477 235 478
rect 174 475 180 476
rect 174 471 175 475
rect 179 471 180 475
rect 174 470 180 471
rect 232 465 234 477
rect 166 464 172 465
rect 166 460 167 464
rect 171 460 172 464
rect 166 459 172 460
rect 230 464 236 465
rect 230 460 231 464
rect 235 460 236 464
rect 230 459 236 460
rect 110 456 116 457
rect 110 452 111 456
rect 115 452 116 456
rect 260 452 262 482
rect 287 477 291 478
rect 303 482 307 483
rect 350 482 356 483
rect 359 482 363 483
rect 303 477 307 478
rect 359 477 363 478
rect 375 482 379 483
rect 375 477 379 478
rect 294 475 300 476
rect 294 471 295 475
rect 299 471 300 475
rect 294 470 300 471
rect 110 451 116 452
rect 158 451 164 452
rect 158 447 159 451
rect 163 447 164 451
rect 158 446 164 447
rect 258 451 264 452
rect 258 447 259 451
rect 263 447 264 451
rect 258 446 264 447
rect 110 439 116 440
rect 110 435 111 439
rect 115 435 116 439
rect 110 434 116 435
rect 112 431 114 434
rect 111 430 115 431
rect 111 425 115 426
rect 151 430 155 431
rect 151 425 155 426
rect 112 422 114 425
rect 150 424 156 425
rect 110 421 116 422
rect 110 417 111 421
rect 115 417 116 421
rect 150 420 151 424
rect 155 420 156 424
rect 150 419 156 420
rect 110 416 116 417
rect 110 404 116 405
rect 110 400 111 404
rect 115 400 116 404
rect 110 399 116 400
rect 112 379 114 399
rect 150 396 156 397
rect 150 392 151 396
rect 155 392 156 396
rect 150 391 156 392
rect 152 379 154 391
rect 160 384 162 446
rect 166 436 172 437
rect 166 432 167 436
rect 171 432 172 436
rect 166 431 172 432
rect 230 436 236 437
rect 230 432 231 436
rect 235 432 236 436
rect 230 431 236 432
rect 167 430 171 431
rect 167 425 171 426
rect 215 430 219 431
rect 215 425 219 426
rect 231 430 235 431
rect 231 425 235 426
rect 279 430 283 431
rect 279 425 283 426
rect 214 424 220 425
rect 214 420 215 424
rect 219 420 220 424
rect 214 419 220 420
rect 278 424 284 425
rect 278 420 279 424
rect 283 420 284 424
rect 278 419 284 420
rect 296 408 298 470
rect 304 465 306 477
rect 376 465 378 477
rect 396 476 398 506
rect 430 500 436 501
rect 430 496 431 500
rect 435 496 436 500
rect 430 495 436 496
rect 510 500 516 501
rect 510 496 511 500
rect 515 496 516 500
rect 510 495 516 496
rect 432 483 434 495
rect 512 483 514 495
rect 548 488 550 506
rect 584 488 586 558
rect 622 548 628 549
rect 622 544 623 548
rect 627 544 628 548
rect 622 543 628 544
rect 624 535 626 543
rect 591 534 595 535
rect 591 529 595 530
rect 623 534 627 535
rect 623 529 627 530
rect 663 534 667 535
rect 663 529 667 530
rect 590 528 596 529
rect 590 524 591 528
rect 595 524 596 528
rect 590 523 596 524
rect 662 528 668 529
rect 662 524 663 528
rect 667 524 668 528
rect 662 523 668 524
rect 692 512 694 582
rect 704 577 706 589
rect 784 577 786 589
rect 810 587 816 588
rect 810 583 811 587
rect 815 583 816 587
rect 810 582 816 583
rect 702 576 708 577
rect 702 572 703 576
rect 707 572 708 576
rect 702 571 708 572
rect 782 576 788 577
rect 782 572 783 576
rect 787 572 788 576
rect 782 571 788 572
rect 812 564 814 582
rect 856 577 858 589
rect 854 576 860 577
rect 854 572 855 576
rect 859 572 860 576
rect 854 571 860 572
rect 880 564 882 598
rect 942 595 948 596
rect 952 595 954 611
rect 1024 604 1026 622
rect 1030 616 1036 617
rect 1030 612 1031 616
rect 1035 612 1036 616
rect 1040 613 1042 622
rect 1094 620 1095 624
rect 1099 620 1100 624
rect 1094 619 1100 620
rect 1134 620 1140 621
rect 1030 611 1036 612
rect 1039 612 1043 613
rect 1022 603 1028 604
rect 1022 599 1023 603
rect 1027 599 1028 603
rect 1022 598 1028 599
rect 1032 595 1034 611
rect 1039 607 1043 608
rect 1096 595 1098 619
rect 1134 616 1135 620
rect 1139 616 1140 620
rect 1134 615 1140 616
rect 1136 595 1138 615
rect 1268 600 1270 662
rect 1286 652 1292 653
rect 1286 648 1287 652
rect 1291 648 1292 652
rect 1286 647 1292 648
rect 1334 652 1340 653
rect 1334 648 1335 652
rect 1339 648 1340 652
rect 1334 647 1340 648
rect 1390 652 1396 653
rect 1390 648 1391 652
rect 1395 648 1396 652
rect 1390 647 1396 648
rect 1446 652 1452 653
rect 1446 648 1447 652
rect 1451 648 1452 652
rect 1446 647 1452 648
rect 1279 646 1283 647
rect 1279 641 1283 642
rect 1287 646 1291 647
rect 1287 641 1291 642
rect 1319 646 1323 647
rect 1319 641 1323 642
rect 1335 646 1339 647
rect 1335 641 1339 642
rect 1367 646 1371 647
rect 1367 641 1371 642
rect 1391 646 1395 647
rect 1391 641 1395 642
rect 1423 646 1427 647
rect 1423 641 1427 642
rect 1447 646 1451 647
rect 1447 641 1451 642
rect 1278 640 1284 641
rect 1278 636 1279 640
rect 1283 636 1284 640
rect 1278 635 1284 636
rect 1318 640 1324 641
rect 1318 636 1319 640
rect 1323 636 1324 640
rect 1318 635 1324 636
rect 1366 640 1372 641
rect 1366 636 1367 640
rect 1371 636 1372 640
rect 1366 635 1372 636
rect 1422 640 1428 641
rect 1422 636 1423 640
rect 1427 636 1428 640
rect 1422 635 1428 636
rect 1342 631 1348 632
rect 1342 627 1343 631
rect 1347 627 1348 631
rect 1342 626 1348 627
rect 1306 623 1312 624
rect 1306 619 1307 623
rect 1311 619 1312 623
rect 1306 618 1312 619
rect 1278 612 1284 613
rect 1278 608 1279 612
rect 1283 608 1284 612
rect 1278 607 1284 608
rect 1266 599 1272 600
rect 1266 595 1267 599
rect 1271 595 1272 599
rect 1280 595 1282 607
rect 1308 600 1310 618
rect 1318 612 1324 613
rect 1318 608 1319 612
rect 1323 608 1324 612
rect 1318 607 1324 608
rect 1306 599 1312 600
rect 1306 595 1307 599
rect 1311 595 1312 599
rect 1320 595 1322 607
rect 927 594 931 595
rect 942 591 943 595
rect 947 591 948 595
rect 942 590 948 591
rect 951 594 955 595
rect 927 589 931 590
rect 928 577 930 589
rect 926 576 932 577
rect 926 572 927 576
rect 931 572 932 576
rect 926 571 932 572
rect 944 564 946 590
rect 951 589 955 590
rect 999 594 1003 595
rect 999 589 1003 590
rect 1031 594 1035 595
rect 1031 589 1035 590
rect 1047 594 1051 595
rect 1047 589 1051 590
rect 1095 594 1099 595
rect 1095 589 1099 590
rect 1135 594 1139 595
rect 1266 594 1272 595
rect 1279 594 1283 595
rect 1306 594 1312 595
rect 1319 594 1323 595
rect 1135 589 1139 590
rect 1279 589 1283 590
rect 1319 589 1323 590
rect 1335 594 1339 595
rect 1335 589 1339 590
rect 986 587 992 588
rect 986 583 987 587
rect 991 583 992 587
rect 986 582 992 583
rect 988 564 990 582
rect 1000 577 1002 589
rect 1048 577 1050 589
rect 1070 587 1076 588
rect 1070 583 1071 587
rect 1075 583 1076 587
rect 1070 582 1076 583
rect 998 576 1004 577
rect 998 572 999 576
rect 1003 572 1004 576
rect 998 571 1004 572
rect 1046 576 1052 577
rect 1046 572 1047 576
rect 1051 572 1052 576
rect 1046 571 1052 572
rect 810 563 816 564
rect 810 559 811 563
rect 815 559 816 563
rect 810 558 816 559
rect 878 563 884 564
rect 878 559 879 563
rect 883 559 884 563
rect 878 558 884 559
rect 942 563 948 564
rect 942 559 943 563
rect 947 559 948 563
rect 942 558 948 559
rect 986 563 992 564
rect 986 559 987 563
rect 991 559 992 563
rect 986 558 992 559
rect 702 548 708 549
rect 702 544 703 548
rect 707 544 708 548
rect 702 543 708 544
rect 782 548 788 549
rect 782 544 783 548
rect 787 544 788 548
rect 782 543 788 544
rect 854 548 860 549
rect 854 544 855 548
rect 859 544 860 548
rect 854 543 860 544
rect 926 548 932 549
rect 926 544 927 548
rect 931 544 932 548
rect 926 543 932 544
rect 998 548 1004 549
rect 998 544 999 548
rect 1003 544 1004 548
rect 998 543 1004 544
rect 1046 548 1052 549
rect 1046 544 1047 548
rect 1051 544 1052 548
rect 1046 543 1052 544
rect 704 535 706 543
rect 784 535 786 543
rect 856 535 858 543
rect 928 535 930 543
rect 1000 535 1002 543
rect 1048 535 1050 543
rect 703 534 707 535
rect 703 529 707 530
rect 735 534 739 535
rect 735 529 739 530
rect 783 534 787 535
rect 783 529 787 530
rect 807 534 811 535
rect 807 529 811 530
rect 855 534 859 535
rect 855 529 859 530
rect 871 534 875 535
rect 871 529 875 530
rect 927 534 931 535
rect 927 529 931 530
rect 935 534 939 535
rect 935 529 939 530
rect 999 534 1003 535
rect 999 529 1003 530
rect 1047 534 1051 535
rect 1047 529 1051 530
rect 734 528 740 529
rect 734 524 735 528
rect 739 524 740 528
rect 734 523 740 524
rect 806 528 812 529
rect 806 524 807 528
rect 811 524 812 528
rect 806 523 812 524
rect 870 528 876 529
rect 870 524 871 528
rect 875 524 876 528
rect 870 523 876 524
rect 934 528 940 529
rect 934 524 935 528
rect 939 524 940 528
rect 934 523 940 524
rect 998 528 1004 529
rect 998 524 999 528
rect 1003 524 1004 528
rect 998 523 1004 524
rect 1046 528 1052 529
rect 1046 524 1047 528
rect 1051 524 1052 528
rect 1046 523 1052 524
rect 966 519 972 520
rect 966 515 967 519
rect 971 515 972 519
rect 966 514 972 515
rect 690 511 696 512
rect 690 507 691 511
rect 695 507 696 511
rect 690 506 696 507
rect 862 511 868 512
rect 862 507 863 511
rect 867 507 868 511
rect 862 506 868 507
rect 926 511 932 512
rect 926 507 927 511
rect 931 507 932 511
rect 926 506 932 507
rect 590 500 596 501
rect 590 496 591 500
rect 595 496 596 500
rect 590 495 596 496
rect 662 500 668 501
rect 662 496 663 500
rect 667 496 668 500
rect 662 495 668 496
rect 734 500 740 501
rect 734 496 735 500
rect 739 496 740 500
rect 734 495 740 496
rect 806 500 812 501
rect 806 496 807 500
rect 811 496 812 500
rect 806 495 812 496
rect 546 487 552 488
rect 546 483 547 487
rect 551 483 552 487
rect 431 482 435 483
rect 431 477 435 478
rect 455 482 459 483
rect 455 477 459 478
rect 511 482 515 483
rect 511 477 515 478
rect 535 482 539 483
rect 546 482 552 483
rect 582 487 588 488
rect 582 483 583 487
rect 587 483 588 487
rect 592 483 594 495
rect 634 487 640 488
rect 634 483 635 487
rect 639 483 640 487
rect 664 483 666 495
rect 736 483 738 495
rect 808 483 810 495
rect 864 488 866 506
rect 870 500 876 501
rect 870 496 871 500
rect 875 496 876 500
rect 870 495 876 496
rect 862 487 868 488
rect 862 483 863 487
rect 867 483 868 487
rect 872 483 874 495
rect 928 488 930 506
rect 934 500 940 501
rect 934 496 935 500
rect 939 496 940 500
rect 934 495 940 496
rect 926 487 932 488
rect 926 483 927 487
rect 931 483 932 487
rect 936 483 938 495
rect 582 482 588 483
rect 591 482 595 483
rect 535 477 539 478
rect 591 477 595 478
rect 607 482 611 483
rect 634 482 640 483
rect 663 482 667 483
rect 607 477 611 478
rect 394 475 400 476
rect 394 471 395 475
rect 399 471 400 475
rect 394 470 400 471
rect 402 475 408 476
rect 402 471 403 475
rect 407 471 408 475
rect 402 470 408 471
rect 302 464 308 465
rect 302 460 303 464
rect 307 460 308 464
rect 302 459 308 460
rect 374 464 380 465
rect 374 460 375 464
rect 379 460 380 464
rect 374 459 380 460
rect 404 452 406 470
rect 456 465 458 477
rect 482 475 488 476
rect 482 471 483 475
rect 487 471 488 475
rect 482 470 488 471
rect 454 464 460 465
rect 454 460 455 464
rect 459 460 460 464
rect 454 459 460 460
rect 484 452 486 470
rect 536 465 538 477
rect 578 475 584 476
rect 578 471 579 475
rect 583 471 584 475
rect 578 470 584 471
rect 534 464 540 465
rect 534 460 535 464
rect 539 460 540 464
rect 534 459 540 460
rect 402 451 408 452
rect 402 447 403 451
rect 407 447 408 451
rect 402 446 408 447
rect 482 451 488 452
rect 482 447 483 451
rect 487 447 488 451
rect 482 446 488 447
rect 494 451 500 452
rect 494 447 495 451
rect 499 447 500 451
rect 494 446 500 447
rect 302 436 308 437
rect 302 432 303 436
rect 307 432 308 436
rect 302 431 308 432
rect 374 436 380 437
rect 374 432 375 436
rect 379 432 380 436
rect 374 431 380 432
rect 454 436 460 437
rect 454 432 455 436
rect 459 432 460 436
rect 454 431 460 432
rect 303 430 307 431
rect 303 425 307 426
rect 351 430 355 431
rect 351 425 355 426
rect 375 430 379 431
rect 375 425 379 426
rect 423 430 427 431
rect 423 425 427 426
rect 455 430 459 431
rect 455 425 459 426
rect 487 430 491 431
rect 487 425 491 426
rect 350 424 356 425
rect 350 420 351 424
rect 355 420 356 424
rect 350 419 356 420
rect 422 424 428 425
rect 422 420 423 424
rect 427 420 428 424
rect 422 419 428 420
rect 486 424 492 425
rect 486 420 487 424
rect 491 420 492 424
rect 486 419 492 420
rect 206 407 212 408
rect 206 403 207 407
rect 211 403 212 407
rect 206 402 212 403
rect 294 407 300 408
rect 294 403 295 407
rect 299 403 300 407
rect 294 402 300 403
rect 390 407 396 408
rect 390 403 391 407
rect 395 403 396 407
rect 390 402 396 403
rect 158 383 164 384
rect 158 379 159 383
rect 163 379 164 383
rect 111 378 115 379
rect 111 373 115 374
rect 135 378 139 379
rect 135 373 139 374
rect 151 378 155 379
rect 158 378 164 379
rect 175 378 179 379
rect 151 373 155 374
rect 175 373 179 374
rect 112 353 114 373
rect 136 361 138 373
rect 176 361 178 373
rect 208 372 210 402
rect 214 396 220 397
rect 214 392 215 396
rect 219 392 220 396
rect 214 391 220 392
rect 278 396 284 397
rect 278 392 279 396
rect 283 392 284 396
rect 278 391 284 392
rect 350 396 356 397
rect 350 392 351 396
rect 355 392 356 396
rect 350 391 356 392
rect 216 379 218 391
rect 280 379 282 391
rect 352 379 354 391
rect 215 378 219 379
rect 215 373 219 374
rect 271 378 275 379
rect 271 373 275 374
rect 279 378 283 379
rect 279 373 283 374
rect 335 378 339 379
rect 335 373 339 374
rect 351 378 355 379
rect 351 373 355 374
rect 206 371 212 372
rect 206 367 207 371
rect 211 367 212 371
rect 206 366 212 367
rect 216 361 218 373
rect 242 371 248 372
rect 242 367 243 371
rect 247 367 248 371
rect 242 366 248 367
rect 134 360 140 361
rect 134 356 135 360
rect 139 356 140 360
rect 134 355 140 356
rect 174 360 180 361
rect 174 356 175 360
rect 179 356 180 360
rect 174 355 180 356
rect 214 360 220 361
rect 214 356 215 360
rect 219 356 220 360
rect 214 355 220 356
rect 110 352 116 353
rect 110 348 111 352
rect 115 348 116 352
rect 244 348 246 366
rect 272 361 274 373
rect 298 371 304 372
rect 298 367 299 371
rect 303 367 304 371
rect 298 366 304 367
rect 270 360 276 361
rect 270 356 271 360
rect 275 356 276 360
rect 270 355 276 356
rect 300 348 302 366
rect 336 361 338 373
rect 392 372 394 402
rect 422 396 428 397
rect 422 392 423 396
rect 427 392 428 396
rect 422 391 428 392
rect 486 396 492 397
rect 486 392 487 396
rect 491 392 492 396
rect 486 391 492 392
rect 424 379 426 391
rect 488 379 490 391
rect 496 384 498 446
rect 534 436 540 437
rect 534 432 535 436
rect 539 432 540 436
rect 534 431 540 432
rect 535 430 539 431
rect 535 425 539 426
rect 551 430 555 431
rect 551 425 555 426
rect 550 424 556 425
rect 550 420 551 424
rect 555 420 556 424
rect 550 419 556 420
rect 580 408 582 470
rect 608 465 610 477
rect 606 464 612 465
rect 606 460 607 464
rect 611 460 612 464
rect 606 459 612 460
rect 636 452 638 482
rect 663 477 667 478
rect 679 482 683 483
rect 679 477 683 478
rect 735 482 739 483
rect 735 477 739 478
rect 743 482 747 483
rect 743 477 747 478
rect 799 482 803 483
rect 799 477 803 478
rect 807 482 811 483
rect 807 477 811 478
rect 855 482 859 483
rect 862 482 868 483
rect 871 482 875 483
rect 855 477 859 478
rect 871 477 875 478
rect 903 482 907 483
rect 926 482 932 483
rect 935 482 939 483
rect 903 477 907 478
rect 935 477 939 478
rect 959 482 963 483
rect 959 477 963 478
rect 680 465 682 477
rect 698 475 704 476
rect 698 471 699 475
rect 703 471 704 475
rect 698 470 704 471
rect 706 475 712 476
rect 706 471 707 475
rect 711 471 712 475
rect 706 470 712 471
rect 678 464 684 465
rect 678 460 679 464
rect 683 460 684 464
rect 678 459 684 460
rect 634 451 640 452
rect 634 447 635 451
rect 639 447 640 451
rect 634 446 640 447
rect 606 436 612 437
rect 606 432 607 436
rect 611 432 612 436
rect 606 431 612 432
rect 678 436 684 437
rect 678 432 679 436
rect 683 432 684 436
rect 678 431 684 432
rect 607 430 611 431
rect 607 425 611 426
rect 615 430 619 431
rect 615 425 619 426
rect 671 430 675 431
rect 671 425 675 426
rect 679 430 683 431
rect 679 425 683 426
rect 614 424 620 425
rect 614 420 615 424
rect 619 420 620 424
rect 614 419 620 420
rect 670 424 676 425
rect 670 420 671 424
rect 675 420 676 424
rect 670 419 676 420
rect 700 416 702 470
rect 708 452 710 470
rect 744 465 746 477
rect 770 475 776 476
rect 770 471 771 475
rect 775 471 776 475
rect 770 470 776 471
rect 742 464 748 465
rect 742 460 743 464
rect 747 460 748 464
rect 742 459 748 460
rect 772 452 774 470
rect 800 465 802 477
rect 826 475 832 476
rect 826 471 827 475
rect 831 471 832 475
rect 826 470 832 471
rect 798 464 804 465
rect 798 460 799 464
rect 803 460 804 464
rect 798 459 804 460
rect 828 452 830 470
rect 856 465 858 477
rect 882 475 888 476
rect 882 471 883 475
rect 887 471 888 475
rect 882 470 888 471
rect 854 464 860 465
rect 854 460 855 464
rect 859 460 860 464
rect 854 459 860 460
rect 884 452 886 470
rect 904 465 906 477
rect 960 465 962 477
rect 968 476 970 514
rect 1072 512 1074 582
rect 1096 569 1098 589
rect 1136 569 1138 589
rect 1336 577 1338 589
rect 1344 588 1346 626
rect 1358 623 1364 624
rect 1358 619 1359 623
rect 1363 619 1364 623
rect 1358 618 1364 619
rect 1406 623 1412 624
rect 1406 619 1407 623
rect 1411 619 1412 623
rect 1406 618 1412 619
rect 1360 600 1362 618
rect 1366 612 1372 613
rect 1366 608 1367 612
rect 1371 608 1372 612
rect 1366 607 1372 608
rect 1358 599 1364 600
rect 1358 595 1359 599
rect 1363 595 1364 599
rect 1368 595 1370 607
rect 1408 600 1410 618
rect 1422 612 1428 613
rect 1422 608 1423 612
rect 1427 608 1428 612
rect 1422 607 1428 608
rect 1406 599 1412 600
rect 1406 595 1407 599
rect 1411 595 1412 599
rect 1424 595 1426 607
rect 1472 600 1474 662
rect 1510 652 1516 653
rect 1510 648 1511 652
rect 1515 648 1516 652
rect 1510 647 1516 648
rect 1574 652 1580 653
rect 1574 648 1575 652
rect 1579 648 1580 652
rect 1574 647 1580 648
rect 1638 652 1644 653
rect 1638 648 1639 652
rect 1643 648 1644 652
rect 1638 647 1644 648
rect 1702 652 1708 653
rect 1702 648 1703 652
rect 1707 648 1708 652
rect 1702 647 1708 648
rect 1479 646 1483 647
rect 1479 641 1483 642
rect 1511 646 1515 647
rect 1511 641 1515 642
rect 1535 646 1539 647
rect 1535 641 1539 642
rect 1575 646 1579 647
rect 1575 641 1579 642
rect 1591 646 1595 647
rect 1591 641 1595 642
rect 1639 646 1643 647
rect 1639 641 1643 642
rect 1647 646 1651 647
rect 1647 641 1651 642
rect 1703 646 1707 647
rect 1703 641 1707 642
rect 1478 640 1484 641
rect 1478 636 1479 640
rect 1483 636 1484 640
rect 1478 635 1484 636
rect 1534 640 1540 641
rect 1534 636 1535 640
rect 1539 636 1540 640
rect 1534 635 1540 636
rect 1590 640 1596 641
rect 1590 636 1591 640
rect 1595 636 1596 640
rect 1590 635 1596 636
rect 1646 640 1652 641
rect 1646 636 1647 640
rect 1651 636 1652 640
rect 1646 635 1652 636
rect 1712 632 1714 682
rect 1732 668 1734 686
rect 1768 681 1770 693
rect 1832 681 1834 693
rect 1858 691 1864 692
rect 1858 687 1859 691
rect 1863 687 1864 691
rect 1858 686 1864 687
rect 1766 680 1772 681
rect 1766 676 1767 680
rect 1771 676 1772 680
rect 1766 675 1772 676
rect 1830 680 1836 681
rect 1830 676 1831 680
rect 1835 676 1836 680
rect 1830 675 1836 676
rect 1860 668 1862 686
rect 1896 681 1898 693
rect 1930 691 1936 692
rect 1930 687 1931 691
rect 1935 687 1936 691
rect 1930 686 1936 687
rect 1894 680 1900 681
rect 1894 676 1895 680
rect 1899 676 1900 680
rect 1894 675 1900 676
rect 1932 668 1934 686
rect 1960 681 1962 693
rect 1958 680 1964 681
rect 1958 676 1959 680
rect 1963 676 1964 680
rect 1958 675 1964 676
rect 1988 668 1990 702
rect 2000 699 2002 715
rect 2072 699 2074 715
rect 1999 698 2003 699
rect 1999 693 2003 694
rect 2023 698 2027 699
rect 2023 693 2027 694
rect 2071 698 2075 699
rect 2071 693 2075 694
rect 2024 681 2026 693
rect 2058 691 2064 692
rect 2058 687 2059 691
rect 2063 687 2064 691
rect 2058 686 2064 687
rect 2022 680 2028 681
rect 2022 676 2023 680
rect 2027 676 2028 680
rect 2022 675 2028 676
rect 2060 668 2062 686
rect 2072 681 2074 693
rect 2080 692 2082 726
rect 2088 708 2090 770
rect 2118 763 2124 764
rect 2118 759 2119 763
rect 2123 759 2124 763
rect 2118 758 2124 759
rect 2120 755 2122 758
rect 2119 754 2123 755
rect 2119 749 2123 750
rect 2120 746 2122 749
rect 2118 745 2124 746
rect 2118 741 2119 745
rect 2123 741 2124 745
rect 2118 740 2124 741
rect 2118 728 2124 729
rect 2118 724 2119 728
rect 2123 724 2124 728
rect 2118 723 2124 724
rect 2086 707 2092 708
rect 2086 703 2087 707
rect 2091 703 2092 707
rect 2086 702 2092 703
rect 2120 699 2122 723
rect 2119 698 2123 699
rect 2119 693 2123 694
rect 2078 691 2084 692
rect 2078 687 2079 691
rect 2083 687 2084 691
rect 2078 686 2084 687
rect 2070 680 2076 681
rect 2070 676 2071 680
rect 2075 676 2076 680
rect 2070 675 2076 676
rect 2120 673 2122 693
rect 2118 672 2124 673
rect 2118 668 2119 672
rect 2123 668 2124 672
rect 1730 667 1736 668
rect 1730 663 1731 667
rect 1735 663 1736 667
rect 1730 662 1736 663
rect 1858 667 1864 668
rect 1858 663 1859 667
rect 1863 663 1864 667
rect 1858 662 1864 663
rect 1930 667 1936 668
rect 1930 663 1931 667
rect 1935 663 1936 667
rect 1930 662 1936 663
rect 1986 667 1992 668
rect 1986 663 1987 667
rect 1991 663 1992 667
rect 1986 662 1992 663
rect 2050 667 2056 668
rect 2050 663 2051 667
rect 2055 663 2056 667
rect 2050 662 2056 663
rect 2058 667 2064 668
rect 2118 667 2124 668
rect 2058 663 2059 667
rect 2063 663 2064 667
rect 2058 662 2064 663
rect 1766 652 1772 653
rect 1766 648 1767 652
rect 1771 648 1772 652
rect 1766 647 1772 648
rect 1830 652 1836 653
rect 1830 648 1831 652
rect 1835 648 1836 652
rect 1830 647 1836 648
rect 1894 652 1900 653
rect 1894 648 1895 652
rect 1899 648 1900 652
rect 1894 647 1900 648
rect 1958 652 1964 653
rect 1958 648 1959 652
rect 1963 648 1964 652
rect 1958 647 1964 648
rect 2022 652 2028 653
rect 2022 648 2023 652
rect 2027 648 2028 652
rect 2022 647 2028 648
rect 1719 646 1723 647
rect 1719 641 1723 642
rect 1767 646 1771 647
rect 1767 641 1771 642
rect 1799 646 1803 647
rect 1799 641 1803 642
rect 1831 646 1835 647
rect 1831 641 1835 642
rect 1879 646 1883 647
rect 1879 641 1883 642
rect 1895 646 1899 647
rect 1895 641 1899 642
rect 1959 646 1963 647
rect 1959 641 1963 642
rect 1967 646 1971 647
rect 1967 641 1971 642
rect 2023 646 2027 647
rect 2023 641 2027 642
rect 1718 640 1724 641
rect 1718 636 1719 640
rect 1723 636 1724 640
rect 1718 635 1724 636
rect 1798 640 1804 641
rect 1798 636 1799 640
rect 1803 636 1804 640
rect 1798 635 1804 636
rect 1878 640 1884 641
rect 1878 636 1879 640
rect 1883 636 1884 640
rect 1878 635 1884 636
rect 1966 640 1972 641
rect 1966 636 1967 640
rect 1971 636 1972 640
rect 1966 635 1972 636
rect 1710 631 1716 632
rect 1710 627 1711 631
rect 1715 627 1716 631
rect 1710 626 1716 627
rect 1526 623 1532 624
rect 1526 619 1527 623
rect 1531 619 1532 623
rect 1526 618 1532 619
rect 1574 623 1580 624
rect 1574 619 1575 623
rect 1579 619 1580 623
rect 1574 618 1580 619
rect 1638 623 1644 624
rect 1638 619 1639 623
rect 1643 619 1644 623
rect 1638 618 1644 619
rect 1710 623 1716 624
rect 1710 619 1711 623
rect 1715 619 1716 623
rect 1710 618 1716 619
rect 1790 623 1796 624
rect 1790 619 1791 623
rect 1795 619 1796 623
rect 1790 618 1796 619
rect 1870 623 1876 624
rect 1870 619 1871 623
rect 1875 619 1876 623
rect 1870 618 1876 619
rect 1958 623 1964 624
rect 1958 619 1959 623
rect 1963 619 1964 623
rect 1958 618 1964 619
rect 1478 612 1484 613
rect 1478 608 1479 612
rect 1483 608 1484 612
rect 1478 607 1484 608
rect 1470 599 1476 600
rect 1470 595 1471 599
rect 1475 595 1476 599
rect 1480 595 1482 607
rect 1528 600 1530 618
rect 1534 612 1540 613
rect 1534 608 1535 612
rect 1539 608 1540 612
rect 1534 607 1540 608
rect 1526 599 1532 600
rect 1526 595 1527 599
rect 1531 595 1532 599
rect 1536 595 1538 607
rect 1358 594 1364 595
rect 1367 594 1371 595
rect 1367 589 1371 590
rect 1375 594 1379 595
rect 1406 594 1412 595
rect 1415 594 1419 595
rect 1375 589 1379 590
rect 1415 589 1419 590
rect 1423 594 1427 595
rect 1423 589 1427 590
rect 1463 594 1467 595
rect 1470 594 1476 595
rect 1479 594 1483 595
rect 1463 589 1467 590
rect 1479 589 1483 590
rect 1519 594 1523 595
rect 1526 594 1532 595
rect 1535 594 1539 595
rect 1519 589 1523 590
rect 1535 589 1539 590
rect 1342 587 1348 588
rect 1342 583 1343 587
rect 1347 583 1348 587
rect 1342 582 1348 583
rect 1358 587 1364 588
rect 1358 583 1359 587
rect 1363 583 1364 587
rect 1358 582 1364 583
rect 1334 576 1340 577
rect 1334 572 1335 576
rect 1339 572 1340 576
rect 1334 571 1340 572
rect 1094 568 1100 569
rect 1094 564 1095 568
rect 1099 564 1100 568
rect 1094 563 1100 564
rect 1134 568 1140 569
rect 1134 564 1135 568
rect 1139 564 1140 568
rect 1360 564 1362 582
rect 1376 577 1378 589
rect 1402 587 1408 588
rect 1402 583 1403 587
rect 1407 583 1408 587
rect 1402 582 1408 583
rect 1374 576 1380 577
rect 1374 572 1375 576
rect 1379 572 1380 576
rect 1374 571 1380 572
rect 1404 564 1406 582
rect 1416 577 1418 589
rect 1442 587 1448 588
rect 1442 583 1443 587
rect 1447 583 1448 587
rect 1442 582 1448 583
rect 1414 576 1420 577
rect 1414 572 1415 576
rect 1419 572 1420 576
rect 1414 571 1420 572
rect 1444 564 1446 582
rect 1464 577 1466 589
rect 1490 587 1496 588
rect 1490 583 1491 587
rect 1495 583 1496 587
rect 1490 582 1496 583
rect 1462 576 1468 577
rect 1462 572 1463 576
rect 1467 572 1468 576
rect 1462 571 1468 572
rect 1492 564 1494 582
rect 1520 577 1522 589
rect 1576 588 1578 618
rect 1590 612 1596 613
rect 1590 608 1591 612
rect 1595 608 1596 612
rect 1590 607 1596 608
rect 1592 595 1594 607
rect 1640 600 1642 618
rect 1646 612 1652 613
rect 1646 608 1647 612
rect 1651 608 1652 612
rect 1646 607 1652 608
rect 1630 599 1636 600
rect 1630 595 1631 599
rect 1635 595 1636 599
rect 1583 594 1587 595
rect 1583 589 1587 590
rect 1591 594 1595 595
rect 1630 594 1636 595
rect 1638 599 1644 600
rect 1638 595 1639 599
rect 1643 595 1644 599
rect 1648 595 1650 607
rect 1712 600 1714 618
rect 1718 612 1724 613
rect 1718 608 1719 612
rect 1723 608 1724 612
rect 1718 607 1724 608
rect 1710 599 1716 600
rect 1710 595 1711 599
rect 1715 595 1716 599
rect 1720 595 1722 607
rect 1792 600 1794 618
rect 1798 612 1804 613
rect 1798 608 1799 612
rect 1803 608 1804 612
rect 1798 607 1804 608
rect 1790 599 1796 600
rect 1790 595 1791 599
rect 1795 595 1796 599
rect 1800 595 1802 607
rect 1872 600 1874 618
rect 1878 612 1884 613
rect 1878 608 1879 612
rect 1883 608 1884 612
rect 1878 607 1884 608
rect 1870 599 1876 600
rect 1870 595 1871 599
rect 1875 595 1876 599
rect 1880 595 1882 607
rect 1960 600 1962 618
rect 1966 612 1972 613
rect 1966 608 1967 612
rect 1971 608 1972 612
rect 1966 607 1972 608
rect 1958 599 1964 600
rect 1958 595 1959 599
rect 1963 595 1964 599
rect 1968 595 1970 607
rect 2052 600 2054 662
rect 2118 655 2124 656
rect 2070 652 2076 653
rect 2070 648 2071 652
rect 2075 648 2076 652
rect 2118 651 2119 655
rect 2123 651 2124 655
rect 2118 650 2124 651
rect 2070 647 2076 648
rect 2120 647 2122 650
rect 2063 646 2067 647
rect 2063 641 2067 642
rect 2071 646 2075 647
rect 2071 641 2075 642
rect 2119 646 2123 647
rect 2119 641 2123 642
rect 2062 640 2068 641
rect 2062 636 2063 640
rect 2067 636 2068 640
rect 2120 638 2122 641
rect 2062 635 2068 636
rect 2118 637 2124 638
rect 2118 633 2119 637
rect 2123 633 2124 637
rect 2118 632 2124 633
rect 2070 623 2076 624
rect 2070 619 2071 623
rect 2075 619 2076 623
rect 2070 618 2076 619
rect 2118 620 2124 621
rect 2062 612 2068 613
rect 2062 608 2063 612
rect 2067 608 2068 612
rect 2062 607 2068 608
rect 2050 599 2056 600
rect 2050 595 2051 599
rect 2055 595 2056 599
rect 2064 595 2066 607
rect 1638 594 1644 595
rect 1647 594 1651 595
rect 1591 589 1595 590
rect 1574 587 1580 588
rect 1574 583 1575 587
rect 1579 583 1580 587
rect 1574 582 1580 583
rect 1584 577 1586 589
rect 1610 587 1616 588
rect 1610 583 1611 587
rect 1615 583 1616 587
rect 1610 582 1616 583
rect 1518 576 1524 577
rect 1518 572 1519 576
rect 1523 572 1524 576
rect 1518 571 1524 572
rect 1582 576 1588 577
rect 1582 572 1583 576
rect 1587 572 1588 576
rect 1582 571 1588 572
rect 1612 564 1614 582
rect 1632 568 1634 594
rect 1647 589 1651 590
rect 1655 594 1659 595
rect 1710 594 1716 595
rect 1719 594 1723 595
rect 1655 589 1659 590
rect 1719 589 1723 590
rect 1727 594 1731 595
rect 1790 594 1796 595
rect 1799 594 1803 595
rect 1727 589 1731 590
rect 1799 589 1803 590
rect 1807 594 1811 595
rect 1870 594 1876 595
rect 1879 594 1883 595
rect 1807 589 1811 590
rect 1879 589 1883 590
rect 1887 594 1891 595
rect 1958 594 1964 595
rect 1967 594 1971 595
rect 1887 589 1891 590
rect 1967 589 1971 590
rect 1975 594 1979 595
rect 2050 594 2056 595
rect 2063 594 2067 595
rect 1975 589 1979 590
rect 2063 589 2067 590
rect 1656 577 1658 589
rect 1728 577 1730 589
rect 1790 587 1796 588
rect 1790 583 1791 587
rect 1795 583 1796 587
rect 1790 582 1796 583
rect 1654 576 1660 577
rect 1654 572 1655 576
rect 1659 572 1660 576
rect 1654 571 1660 572
rect 1726 576 1732 577
rect 1726 572 1727 576
rect 1731 572 1732 576
rect 1726 571 1732 572
rect 1630 567 1636 568
rect 1134 563 1140 564
rect 1358 563 1364 564
rect 1358 559 1359 563
rect 1363 559 1364 563
rect 1358 558 1364 559
rect 1402 563 1408 564
rect 1402 559 1403 563
rect 1407 559 1408 563
rect 1402 558 1408 559
rect 1442 563 1448 564
rect 1442 559 1443 563
rect 1447 559 1448 563
rect 1442 558 1448 559
rect 1490 563 1496 564
rect 1490 559 1491 563
rect 1495 559 1496 563
rect 1490 558 1496 559
rect 1502 563 1508 564
rect 1502 559 1503 563
rect 1507 559 1508 563
rect 1502 558 1508 559
rect 1610 563 1616 564
rect 1610 559 1611 563
rect 1615 559 1616 563
rect 1630 563 1631 567
rect 1635 563 1636 567
rect 1792 564 1794 582
rect 1808 577 1810 589
rect 1870 587 1876 588
rect 1870 583 1871 587
rect 1875 583 1876 587
rect 1870 582 1876 583
rect 1878 583 1884 584
rect 1806 576 1812 577
rect 1806 572 1807 576
rect 1811 572 1812 576
rect 1806 571 1812 572
rect 1872 564 1874 582
rect 1878 579 1879 583
rect 1883 579 1884 583
rect 1878 578 1884 579
rect 1630 562 1636 563
rect 1678 563 1684 564
rect 1610 558 1616 559
rect 1678 559 1679 563
rect 1683 559 1684 563
rect 1678 558 1684 559
rect 1790 563 1796 564
rect 1790 559 1791 563
rect 1795 559 1796 563
rect 1790 558 1796 559
rect 1870 563 1876 564
rect 1870 559 1871 563
rect 1875 559 1876 563
rect 1870 558 1876 559
rect 1094 551 1100 552
rect 1094 547 1095 551
rect 1099 547 1100 551
rect 1094 546 1100 547
rect 1134 551 1140 552
rect 1134 547 1135 551
rect 1139 547 1140 551
rect 1134 546 1140 547
rect 1334 548 1340 549
rect 1096 535 1098 546
rect 1136 539 1138 546
rect 1334 544 1335 548
rect 1339 544 1340 548
rect 1334 543 1340 544
rect 1374 548 1380 549
rect 1374 544 1375 548
rect 1379 544 1380 548
rect 1374 543 1380 544
rect 1414 548 1420 549
rect 1414 544 1415 548
rect 1419 544 1420 548
rect 1414 543 1420 544
rect 1462 548 1468 549
rect 1462 544 1463 548
rect 1467 544 1468 548
rect 1462 543 1468 544
rect 1336 539 1338 543
rect 1376 539 1378 543
rect 1416 539 1418 543
rect 1464 539 1466 543
rect 1135 538 1139 539
rect 1095 534 1099 535
rect 1135 533 1139 534
rect 1191 538 1195 539
rect 1191 533 1195 534
rect 1239 538 1243 539
rect 1239 533 1243 534
rect 1287 538 1291 539
rect 1287 533 1291 534
rect 1335 538 1339 539
rect 1335 533 1339 534
rect 1343 538 1347 539
rect 1343 533 1347 534
rect 1375 538 1379 539
rect 1375 533 1379 534
rect 1407 538 1411 539
rect 1407 533 1411 534
rect 1415 538 1419 539
rect 1415 533 1419 534
rect 1463 538 1467 539
rect 1463 533 1467 534
rect 1479 538 1483 539
rect 1479 533 1483 534
rect 1136 530 1138 533
rect 1190 532 1196 533
rect 1095 529 1099 530
rect 1134 529 1140 530
rect 1096 526 1098 529
rect 1094 525 1100 526
rect 1094 521 1095 525
rect 1099 521 1100 525
rect 1134 525 1135 529
rect 1139 525 1140 529
rect 1190 528 1191 532
rect 1195 528 1196 532
rect 1190 527 1196 528
rect 1238 532 1244 533
rect 1238 528 1239 532
rect 1243 528 1244 532
rect 1238 527 1244 528
rect 1286 532 1292 533
rect 1286 528 1287 532
rect 1291 528 1292 532
rect 1286 527 1292 528
rect 1342 532 1348 533
rect 1342 528 1343 532
rect 1347 528 1348 532
rect 1342 527 1348 528
rect 1406 532 1412 533
rect 1406 528 1407 532
rect 1411 528 1412 532
rect 1406 527 1412 528
rect 1478 532 1484 533
rect 1478 528 1479 532
rect 1483 528 1484 532
rect 1478 527 1484 528
rect 1134 524 1140 525
rect 1094 520 1100 521
rect 1214 523 1220 524
rect 1206 519 1212 520
rect 1206 515 1207 519
rect 1211 515 1212 519
rect 1214 519 1215 523
rect 1219 519 1220 523
rect 1214 518 1220 519
rect 1206 514 1212 515
rect 1134 512 1140 513
rect 990 511 996 512
rect 990 507 991 511
rect 995 507 996 511
rect 990 506 996 507
rect 1038 511 1044 512
rect 1038 507 1039 511
rect 1043 507 1044 511
rect 1038 506 1044 507
rect 1070 511 1076 512
rect 1070 507 1071 511
rect 1075 507 1076 511
rect 1070 506 1076 507
rect 1094 508 1100 509
rect 992 488 994 506
rect 998 500 1004 501
rect 998 496 999 500
rect 1003 496 1004 500
rect 998 495 1004 496
rect 990 487 996 488
rect 990 483 991 487
rect 995 483 996 487
rect 1000 483 1002 495
rect 1040 488 1042 506
rect 1094 504 1095 508
rect 1099 504 1100 508
rect 1134 508 1135 512
rect 1139 508 1140 512
rect 1134 507 1140 508
rect 1094 503 1100 504
rect 1046 500 1052 501
rect 1046 496 1047 500
rect 1051 496 1052 500
rect 1046 495 1052 496
rect 1038 487 1044 488
rect 1038 483 1039 487
rect 1043 483 1044 487
rect 1048 483 1050 495
rect 1096 483 1098 503
rect 1136 487 1138 507
rect 1190 504 1196 505
rect 1190 500 1191 504
rect 1195 500 1196 504
rect 1190 499 1196 500
rect 1192 487 1194 499
rect 1135 486 1139 487
rect 990 482 996 483
rect 999 482 1003 483
rect 999 477 1003 478
rect 1007 482 1011 483
rect 1038 482 1044 483
rect 1047 482 1051 483
rect 1007 477 1011 478
rect 1095 482 1099 483
rect 1047 477 1051 478
rect 1074 479 1080 480
rect 966 475 972 476
rect 966 471 967 475
rect 971 471 972 475
rect 966 470 972 471
rect 986 475 992 476
rect 986 471 987 475
rect 991 471 992 475
rect 986 470 992 471
rect 902 464 908 465
rect 902 460 903 464
rect 907 460 908 464
rect 902 459 908 460
rect 958 464 964 465
rect 958 460 959 464
rect 963 460 964 464
rect 958 459 964 460
rect 988 452 990 470
rect 1008 465 1010 477
rect 1034 475 1040 476
rect 1034 471 1035 475
rect 1039 471 1040 475
rect 1034 470 1040 471
rect 1006 464 1012 465
rect 1006 460 1007 464
rect 1011 460 1012 464
rect 1006 459 1012 460
rect 1036 452 1038 470
rect 1048 465 1050 477
rect 1074 475 1075 479
rect 1079 475 1080 479
rect 1135 481 1139 482
rect 1159 486 1163 487
rect 1159 481 1163 482
rect 1191 486 1195 487
rect 1191 481 1195 482
rect 1095 477 1099 478
rect 1074 474 1080 475
rect 1046 464 1052 465
rect 1046 460 1047 464
rect 1051 460 1052 464
rect 1046 459 1052 460
rect 1076 452 1078 474
rect 1096 457 1098 477
rect 1136 461 1138 481
rect 1160 469 1162 481
rect 1158 468 1164 469
rect 1158 464 1159 468
rect 1163 464 1164 468
rect 1158 463 1164 464
rect 1134 460 1140 461
rect 1094 456 1100 457
rect 1094 452 1095 456
rect 1099 452 1100 456
rect 1134 456 1135 460
rect 1139 456 1140 460
rect 1208 456 1210 514
rect 1216 492 1218 518
rect 1230 515 1236 516
rect 1230 511 1231 515
rect 1235 511 1236 515
rect 1230 510 1236 511
rect 1278 515 1284 516
rect 1278 511 1279 515
rect 1283 511 1284 515
rect 1278 510 1284 511
rect 1358 515 1364 516
rect 1358 511 1359 515
rect 1363 511 1364 515
rect 1358 510 1364 511
rect 1442 515 1448 516
rect 1442 511 1443 515
rect 1447 511 1448 515
rect 1442 510 1448 511
rect 1232 492 1234 510
rect 1238 504 1244 505
rect 1238 500 1239 504
rect 1243 500 1244 504
rect 1238 499 1244 500
rect 1214 491 1220 492
rect 1214 487 1215 491
rect 1219 487 1220 491
rect 1214 486 1220 487
rect 1230 491 1236 492
rect 1230 487 1231 491
rect 1235 487 1236 491
rect 1240 487 1242 499
rect 1280 492 1282 510
rect 1286 504 1292 505
rect 1286 500 1287 504
rect 1291 500 1292 504
rect 1286 499 1292 500
rect 1342 504 1348 505
rect 1342 500 1343 504
rect 1347 500 1348 504
rect 1342 499 1348 500
rect 1278 491 1284 492
rect 1278 487 1279 491
rect 1283 487 1284 491
rect 1288 487 1290 499
rect 1344 487 1346 499
rect 1230 486 1236 487
rect 1239 486 1243 487
rect 1239 481 1243 482
rect 1263 486 1267 487
rect 1278 486 1284 487
rect 1287 486 1291 487
rect 1263 481 1267 482
rect 1287 481 1291 482
rect 1343 486 1347 487
rect 1343 481 1347 482
rect 1264 469 1266 481
rect 1360 480 1362 510
rect 1406 504 1412 505
rect 1406 500 1407 504
rect 1411 500 1412 504
rect 1406 499 1412 500
rect 1408 487 1410 499
rect 1444 492 1446 510
rect 1478 504 1484 505
rect 1478 500 1479 504
rect 1483 500 1484 504
rect 1478 499 1484 500
rect 1442 491 1448 492
rect 1442 487 1443 491
rect 1447 487 1448 491
rect 1480 487 1482 499
rect 1504 492 1506 558
rect 1518 548 1524 549
rect 1518 544 1519 548
rect 1523 544 1524 548
rect 1518 543 1524 544
rect 1582 548 1588 549
rect 1582 544 1583 548
rect 1587 544 1588 548
rect 1582 543 1588 544
rect 1654 548 1660 549
rect 1654 544 1655 548
rect 1659 544 1660 548
rect 1654 543 1660 544
rect 1520 539 1522 543
rect 1550 539 1556 540
rect 1584 539 1586 543
rect 1656 539 1658 543
rect 1680 540 1682 558
rect 1726 548 1732 549
rect 1726 544 1727 548
rect 1731 544 1732 548
rect 1726 543 1732 544
rect 1806 548 1812 549
rect 1806 544 1807 548
rect 1811 544 1812 548
rect 1806 543 1812 544
rect 1678 539 1684 540
rect 1728 539 1730 543
rect 1808 539 1810 543
rect 1519 538 1523 539
rect 1519 533 1523 534
rect 1543 538 1547 539
rect 1550 535 1551 539
rect 1555 535 1556 539
rect 1550 534 1556 535
rect 1583 538 1587 539
rect 1543 533 1547 534
rect 1542 532 1548 533
rect 1542 528 1543 532
rect 1547 528 1548 532
rect 1542 527 1548 528
rect 1542 504 1548 505
rect 1542 500 1543 504
rect 1547 500 1548 504
rect 1542 499 1548 500
rect 1502 491 1508 492
rect 1502 487 1503 491
rect 1507 487 1508 491
rect 1544 487 1546 499
rect 1552 492 1554 534
rect 1583 533 1587 534
rect 1607 538 1611 539
rect 1607 533 1611 534
rect 1655 538 1659 539
rect 1655 533 1659 534
rect 1671 538 1675 539
rect 1678 535 1679 539
rect 1683 535 1684 539
rect 1678 534 1684 535
rect 1727 538 1731 539
rect 1671 533 1675 534
rect 1727 533 1731 534
rect 1735 538 1739 539
rect 1735 533 1739 534
rect 1799 538 1803 539
rect 1799 533 1803 534
rect 1807 538 1811 539
rect 1807 533 1811 534
rect 1863 538 1867 539
rect 1863 533 1867 534
rect 1606 532 1612 533
rect 1606 528 1607 532
rect 1611 528 1612 532
rect 1606 527 1612 528
rect 1670 532 1676 533
rect 1670 528 1671 532
rect 1675 528 1676 532
rect 1670 527 1676 528
rect 1734 532 1740 533
rect 1734 528 1735 532
rect 1739 528 1740 532
rect 1734 527 1740 528
rect 1798 532 1804 533
rect 1798 528 1799 532
rect 1803 528 1804 532
rect 1798 527 1804 528
rect 1862 532 1868 533
rect 1862 528 1863 532
rect 1867 528 1868 532
rect 1862 527 1868 528
rect 1758 523 1764 524
rect 1758 519 1759 523
rect 1763 519 1764 523
rect 1758 518 1764 519
rect 1590 515 1596 516
rect 1590 511 1591 515
rect 1595 511 1596 515
rect 1590 510 1596 511
rect 1662 515 1668 516
rect 1662 511 1663 515
rect 1667 511 1668 515
rect 1662 510 1668 511
rect 1694 515 1700 516
rect 1694 511 1695 515
rect 1699 511 1700 515
rect 1694 510 1700 511
rect 1592 492 1594 510
rect 1606 504 1612 505
rect 1606 500 1607 504
rect 1611 500 1612 504
rect 1606 499 1612 500
rect 1550 491 1556 492
rect 1550 487 1551 491
rect 1555 487 1556 491
rect 1383 486 1387 487
rect 1383 481 1387 482
rect 1407 486 1411 487
rect 1442 486 1448 487
rect 1479 486 1483 487
rect 1407 481 1411 482
rect 1479 481 1483 482
rect 1495 486 1499 487
rect 1502 486 1508 487
rect 1543 486 1547 487
rect 1550 486 1556 487
rect 1590 491 1596 492
rect 1590 487 1591 491
rect 1595 487 1596 491
rect 1608 487 1610 499
rect 1664 492 1666 510
rect 1670 504 1676 505
rect 1670 500 1671 504
rect 1675 500 1676 504
rect 1670 499 1676 500
rect 1662 491 1668 492
rect 1662 487 1663 491
rect 1667 487 1668 491
rect 1672 487 1674 499
rect 1590 486 1596 487
rect 1599 486 1603 487
rect 1495 481 1499 482
rect 1543 481 1547 482
rect 1599 481 1603 482
rect 1607 486 1611 487
rect 1662 486 1668 487
rect 1671 486 1675 487
rect 1607 481 1611 482
rect 1671 481 1675 482
rect 1350 479 1356 480
rect 1350 475 1351 479
rect 1355 475 1356 479
rect 1350 474 1356 475
rect 1358 479 1364 480
rect 1358 475 1359 479
rect 1363 475 1364 479
rect 1358 474 1364 475
rect 1262 468 1268 469
rect 1262 464 1263 468
rect 1267 464 1268 468
rect 1262 463 1268 464
rect 1352 456 1354 474
rect 1384 469 1386 481
rect 1496 469 1498 481
rect 1586 479 1592 480
rect 1586 475 1587 479
rect 1591 475 1592 479
rect 1586 474 1592 475
rect 1382 468 1388 469
rect 1382 464 1383 468
rect 1387 464 1388 468
rect 1382 463 1388 464
rect 1494 468 1500 469
rect 1494 464 1495 468
rect 1499 464 1500 468
rect 1588 467 1590 474
rect 1600 469 1602 481
rect 1696 480 1698 510
rect 1734 504 1740 505
rect 1734 500 1735 504
rect 1739 500 1740 504
rect 1734 499 1740 500
rect 1736 487 1738 499
rect 1760 492 1762 518
rect 1880 516 1882 578
rect 1888 577 1890 589
rect 1976 577 1978 589
rect 2050 587 2056 588
rect 2050 583 2051 587
rect 2055 583 2056 587
rect 2050 582 2056 583
rect 1886 576 1892 577
rect 1886 572 1887 576
rect 1891 572 1892 576
rect 1886 571 1892 572
rect 1974 576 1980 577
rect 1974 572 1975 576
rect 1979 572 1980 576
rect 1974 571 1980 572
rect 2052 564 2054 582
rect 2064 577 2066 589
rect 2072 588 2074 618
rect 2118 616 2119 620
rect 2123 616 2124 620
rect 2118 615 2124 616
rect 2120 595 2122 615
rect 2119 594 2123 595
rect 2119 589 2123 590
rect 2070 587 2076 588
rect 2070 583 2071 587
rect 2075 583 2076 587
rect 2070 582 2076 583
rect 2062 576 2068 577
rect 2062 572 2063 576
rect 2067 572 2068 576
rect 2062 571 2068 572
rect 2120 569 2122 589
rect 2118 568 2124 569
rect 2118 564 2119 568
rect 2123 564 2124 568
rect 1998 563 2004 564
rect 1998 559 1999 563
rect 2003 559 2004 563
rect 1998 558 2004 559
rect 2050 563 2056 564
rect 2118 563 2124 564
rect 2050 559 2051 563
rect 2055 559 2056 563
rect 2050 558 2056 559
rect 1886 548 1892 549
rect 1886 544 1887 548
rect 1891 544 1892 548
rect 1886 543 1892 544
rect 1974 548 1980 549
rect 1974 544 1975 548
rect 1979 544 1980 548
rect 1974 543 1980 544
rect 1888 539 1890 543
rect 1976 539 1978 543
rect 1887 538 1891 539
rect 1887 533 1891 534
rect 1935 538 1939 539
rect 1935 533 1939 534
rect 1975 538 1979 539
rect 1975 533 1979 534
rect 1934 532 1940 533
rect 1934 528 1935 532
rect 1939 528 1940 532
rect 1934 527 1940 528
rect 1790 515 1796 516
rect 1790 511 1791 515
rect 1795 511 1796 515
rect 1790 510 1796 511
rect 1854 515 1860 516
rect 1854 511 1855 515
rect 1859 511 1860 515
rect 1854 510 1860 511
rect 1878 515 1884 516
rect 1878 511 1879 515
rect 1883 511 1884 515
rect 1878 510 1884 511
rect 1792 492 1794 510
rect 1798 504 1804 505
rect 1798 500 1799 504
rect 1803 500 1804 504
rect 1798 499 1804 500
rect 1758 491 1764 492
rect 1758 487 1759 491
rect 1763 487 1764 491
rect 1703 486 1707 487
rect 1703 481 1707 482
rect 1735 486 1739 487
rect 1758 486 1764 487
rect 1790 491 1796 492
rect 1790 487 1791 491
rect 1795 487 1796 491
rect 1800 487 1802 499
rect 1856 492 1858 510
rect 1862 504 1868 505
rect 1862 500 1863 504
rect 1867 500 1868 504
rect 1862 499 1868 500
rect 1934 504 1940 505
rect 1934 500 1935 504
rect 1939 500 1940 504
rect 1934 499 1940 500
rect 1854 491 1860 492
rect 1854 487 1855 491
rect 1859 487 1860 491
rect 1864 487 1866 499
rect 1936 487 1938 499
rect 2000 492 2002 558
rect 2118 551 2124 552
rect 2062 548 2068 549
rect 2062 544 2063 548
rect 2067 544 2068 548
rect 2118 547 2119 551
rect 2123 547 2124 551
rect 2118 546 2124 547
rect 2062 543 2068 544
rect 2064 539 2066 543
rect 2120 539 2122 546
rect 2007 538 2011 539
rect 2007 533 2011 534
rect 2063 538 2067 539
rect 2063 533 2067 534
rect 2071 538 2075 539
rect 2071 533 2075 534
rect 2119 538 2123 539
rect 2119 533 2123 534
rect 2006 532 2012 533
rect 2006 528 2007 532
rect 2011 528 2012 532
rect 2006 527 2012 528
rect 2070 532 2076 533
rect 2070 528 2071 532
rect 2075 528 2076 532
rect 2120 530 2122 533
rect 2070 527 2076 528
rect 2118 529 2124 530
rect 2118 525 2119 529
rect 2123 525 2124 529
rect 2118 524 2124 525
rect 2062 515 2068 516
rect 2062 511 2063 515
rect 2067 511 2068 515
rect 2062 510 2068 511
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2118 512 2124 513
rect 2006 504 2012 505
rect 2006 500 2007 504
rect 2011 500 2012 504
rect 2006 499 2012 500
rect 1966 491 1972 492
rect 1966 487 1967 491
rect 1971 487 1972 491
rect 1998 491 2004 492
rect 1998 487 1999 491
rect 2003 487 2004 491
rect 2008 487 2010 499
rect 2064 492 2066 510
rect 2070 504 2076 505
rect 2070 500 2071 504
rect 2075 500 2076 504
rect 2070 499 2076 500
rect 2062 491 2068 492
rect 2062 487 2063 491
rect 2067 487 2068 491
rect 2072 487 2074 499
rect 1790 486 1796 487
rect 1799 486 1803 487
rect 1854 486 1860 487
rect 1863 486 1867 487
rect 1735 481 1739 482
rect 1799 481 1803 482
rect 1863 481 1867 482
rect 1887 486 1891 487
rect 1887 481 1891 482
rect 1935 486 1939 487
rect 1966 486 1972 487
rect 1983 486 1987 487
rect 1998 486 2004 487
rect 2007 486 2011 487
rect 2062 486 2068 487
rect 2071 486 2075 487
rect 1935 481 1939 482
rect 1686 479 1692 480
rect 1686 475 1687 479
rect 1691 475 1692 479
rect 1686 474 1692 475
rect 1694 479 1700 480
rect 1694 475 1695 479
rect 1699 475 1700 479
rect 1694 474 1700 475
rect 1598 468 1604 469
rect 1588 465 1594 467
rect 1494 463 1500 464
rect 1592 456 1594 465
rect 1598 464 1599 468
rect 1603 464 1604 468
rect 1598 463 1604 464
rect 1688 456 1690 474
rect 1704 469 1706 481
rect 1800 469 1802 481
rect 1826 479 1832 480
rect 1826 475 1827 479
rect 1831 475 1832 479
rect 1826 474 1832 475
rect 1702 468 1708 469
rect 1702 464 1703 468
rect 1707 464 1708 468
rect 1702 463 1708 464
rect 1798 468 1804 469
rect 1798 464 1799 468
rect 1803 464 1804 468
rect 1798 463 1804 464
rect 1828 456 1830 474
rect 1846 471 1852 472
rect 1846 467 1847 471
rect 1851 467 1852 471
rect 1888 469 1890 481
rect 1914 479 1920 480
rect 1914 475 1915 479
rect 1919 475 1920 479
rect 1914 474 1920 475
rect 1846 466 1852 467
rect 1886 468 1892 469
rect 1134 455 1140 456
rect 1166 455 1172 456
rect 706 451 712 452
rect 706 447 707 451
rect 711 447 712 451
rect 706 446 712 447
rect 770 451 776 452
rect 770 447 771 451
rect 775 447 776 451
rect 770 446 776 447
rect 826 451 832 452
rect 826 447 827 451
rect 831 447 832 451
rect 826 446 832 447
rect 882 451 888 452
rect 882 447 883 451
rect 887 447 888 451
rect 882 446 888 447
rect 986 451 992 452
rect 986 447 987 451
rect 991 447 992 451
rect 986 446 992 447
rect 1034 451 1040 452
rect 1034 447 1035 451
rect 1039 447 1040 451
rect 1034 446 1040 447
rect 1074 451 1080 452
rect 1094 451 1100 452
rect 1166 451 1167 455
rect 1171 451 1172 455
rect 1074 447 1075 451
rect 1079 447 1080 451
rect 1166 450 1172 451
rect 1206 455 1212 456
rect 1206 451 1207 455
rect 1211 451 1212 455
rect 1206 450 1212 451
rect 1350 455 1356 456
rect 1350 451 1351 455
rect 1355 451 1356 455
rect 1350 450 1356 451
rect 1582 455 1588 456
rect 1582 451 1583 455
rect 1587 451 1588 455
rect 1582 450 1588 451
rect 1590 455 1596 456
rect 1590 451 1591 455
rect 1595 451 1596 455
rect 1590 450 1596 451
rect 1686 455 1692 456
rect 1686 451 1687 455
rect 1691 451 1692 455
rect 1686 450 1692 451
rect 1826 455 1832 456
rect 1826 451 1827 455
rect 1831 451 1832 455
rect 1826 450 1832 451
rect 1074 446 1080 447
rect 1134 443 1140 444
rect 1094 439 1100 440
rect 742 436 748 437
rect 742 432 743 436
rect 747 432 748 436
rect 742 431 748 432
rect 798 436 804 437
rect 798 432 799 436
rect 803 432 804 436
rect 798 431 804 432
rect 854 436 860 437
rect 854 432 855 436
rect 859 432 860 436
rect 854 431 860 432
rect 902 436 908 437
rect 902 432 903 436
rect 907 432 908 436
rect 902 431 908 432
rect 958 436 964 437
rect 958 432 959 436
rect 963 432 964 436
rect 958 431 964 432
rect 1006 436 1012 437
rect 1006 432 1007 436
rect 1011 432 1012 436
rect 1006 431 1012 432
rect 1046 436 1052 437
rect 1046 432 1047 436
rect 1051 432 1052 436
rect 1094 435 1095 439
rect 1099 435 1100 439
rect 1134 439 1135 443
rect 1139 439 1140 443
rect 1134 438 1140 439
rect 1158 440 1164 441
rect 1136 435 1138 438
rect 1158 436 1159 440
rect 1163 436 1164 440
rect 1158 435 1164 436
rect 1094 434 1100 435
rect 1135 434 1139 435
rect 1046 431 1052 432
rect 1096 431 1098 434
rect 727 430 731 431
rect 727 425 731 426
rect 743 430 747 431
rect 743 425 747 426
rect 791 430 795 431
rect 791 425 795 426
rect 799 430 803 431
rect 799 425 803 426
rect 855 430 859 431
rect 855 425 859 426
rect 903 430 907 431
rect 903 425 907 426
rect 959 430 963 431
rect 959 425 963 426
rect 1007 430 1011 431
rect 1007 425 1011 426
rect 1047 430 1051 431
rect 1047 425 1051 426
rect 1095 430 1099 431
rect 1135 429 1139 430
rect 1159 434 1163 435
rect 1159 429 1163 430
rect 1136 426 1138 429
rect 1158 428 1164 429
rect 1095 425 1099 426
rect 1134 425 1140 426
rect 726 424 732 425
rect 726 420 727 424
rect 731 420 732 424
rect 726 419 732 420
rect 790 424 796 425
rect 790 420 791 424
rect 795 420 796 424
rect 790 419 796 420
rect 854 424 860 425
rect 854 420 855 424
rect 859 420 860 424
rect 1096 422 1098 425
rect 854 419 860 420
rect 1094 421 1100 422
rect 1094 417 1095 421
rect 1099 417 1100 421
rect 1134 421 1135 425
rect 1139 421 1140 425
rect 1158 424 1159 428
rect 1163 424 1164 428
rect 1158 423 1164 424
rect 1134 420 1140 421
rect 1094 416 1100 417
rect 698 415 704 416
rect 698 411 699 415
rect 703 411 704 415
rect 698 410 704 411
rect 1134 408 1140 409
rect 578 407 584 408
rect 578 403 579 407
rect 583 403 584 407
rect 578 402 584 403
rect 662 407 668 408
rect 662 403 663 407
rect 667 403 668 407
rect 662 402 668 403
rect 718 407 724 408
rect 718 403 719 407
rect 723 403 724 407
rect 718 402 724 403
rect 782 407 788 408
rect 782 403 783 407
rect 787 403 788 407
rect 782 402 788 403
rect 846 407 852 408
rect 846 403 847 407
rect 851 403 852 407
rect 846 402 852 403
rect 1094 404 1100 405
rect 550 396 556 397
rect 550 392 551 396
rect 555 392 556 396
rect 550 391 556 392
rect 614 396 620 397
rect 614 392 615 396
rect 619 392 620 396
rect 614 391 620 392
rect 494 383 500 384
rect 494 379 495 383
rect 499 379 500 383
rect 542 383 548 384
rect 542 379 543 383
rect 547 379 548 383
rect 552 379 554 391
rect 602 383 608 384
rect 602 379 603 383
rect 607 379 608 383
rect 616 379 618 391
rect 664 384 666 402
rect 670 396 676 397
rect 670 392 671 396
rect 675 392 676 396
rect 670 391 676 392
rect 662 383 668 384
rect 662 379 663 383
rect 667 379 668 383
rect 672 379 674 391
rect 720 384 722 402
rect 726 396 732 397
rect 726 392 727 396
rect 731 392 732 396
rect 726 391 732 392
rect 718 383 724 384
rect 718 379 719 383
rect 723 379 724 383
rect 728 379 730 391
rect 784 384 786 402
rect 790 396 796 397
rect 790 392 791 396
rect 795 392 796 396
rect 790 391 796 392
rect 782 383 788 384
rect 782 379 783 383
rect 787 379 788 383
rect 792 379 794 391
rect 848 384 850 402
rect 1094 400 1095 404
rect 1099 400 1100 404
rect 1134 404 1135 408
rect 1139 404 1140 408
rect 1134 403 1140 404
rect 1094 399 1100 400
rect 854 396 860 397
rect 854 392 855 396
rect 859 392 860 396
rect 854 391 860 392
rect 846 383 852 384
rect 846 379 847 383
rect 851 379 852 383
rect 856 379 858 391
rect 1096 379 1098 399
rect 1136 379 1138 403
rect 1158 400 1164 401
rect 1158 396 1159 400
rect 1163 396 1164 400
rect 1158 395 1164 396
rect 1160 379 1162 395
rect 1168 388 1170 450
rect 1262 440 1268 441
rect 1262 436 1263 440
rect 1267 436 1268 440
rect 1262 435 1268 436
rect 1382 440 1388 441
rect 1382 436 1383 440
rect 1387 436 1388 440
rect 1382 435 1388 436
rect 1494 440 1500 441
rect 1494 436 1495 440
rect 1499 436 1500 440
rect 1494 435 1500 436
rect 1199 434 1203 435
rect 1199 429 1203 430
rect 1255 434 1259 435
rect 1255 429 1259 430
rect 1263 434 1267 435
rect 1263 429 1267 430
rect 1335 434 1339 435
rect 1335 429 1339 430
rect 1383 434 1387 435
rect 1383 429 1387 430
rect 1415 434 1419 435
rect 1415 429 1419 430
rect 1495 434 1499 435
rect 1495 429 1499 430
rect 1503 434 1507 435
rect 1503 429 1507 430
rect 1198 428 1204 429
rect 1198 424 1199 428
rect 1203 424 1204 428
rect 1198 423 1204 424
rect 1254 428 1260 429
rect 1254 424 1255 428
rect 1259 424 1260 428
rect 1254 423 1260 424
rect 1334 428 1340 429
rect 1334 424 1335 428
rect 1339 424 1340 428
rect 1334 423 1340 424
rect 1414 428 1420 429
rect 1414 424 1415 428
rect 1419 424 1420 428
rect 1414 423 1420 424
rect 1502 428 1508 429
rect 1502 424 1503 428
rect 1507 424 1508 428
rect 1502 423 1508 424
rect 1186 411 1192 412
rect 1186 407 1187 411
rect 1191 407 1192 411
rect 1186 406 1192 407
rect 1246 411 1252 412
rect 1246 407 1247 411
rect 1251 407 1252 411
rect 1246 406 1252 407
rect 1326 411 1332 412
rect 1326 407 1327 411
rect 1331 407 1332 411
rect 1326 406 1332 407
rect 1406 411 1412 412
rect 1406 407 1407 411
rect 1411 407 1412 411
rect 1406 406 1412 407
rect 1494 411 1500 412
rect 1494 407 1495 411
rect 1499 407 1500 411
rect 1494 406 1500 407
rect 1510 411 1516 412
rect 1510 407 1511 411
rect 1515 407 1516 411
rect 1510 406 1516 407
rect 1188 388 1190 406
rect 1198 400 1204 401
rect 1198 396 1199 400
rect 1203 396 1204 400
rect 1198 395 1204 396
rect 1166 387 1172 388
rect 1166 383 1167 387
rect 1171 383 1172 387
rect 1166 382 1172 383
rect 1186 387 1192 388
rect 1186 383 1187 387
rect 1191 383 1192 387
rect 1186 382 1192 383
rect 1200 379 1202 395
rect 1248 388 1250 406
rect 1254 400 1260 401
rect 1254 396 1255 400
rect 1259 396 1260 400
rect 1254 395 1260 396
rect 1246 387 1252 388
rect 1246 383 1247 387
rect 1251 383 1252 387
rect 1246 382 1252 383
rect 1256 379 1258 395
rect 1328 388 1330 406
rect 1334 400 1340 401
rect 1334 396 1335 400
rect 1339 396 1340 400
rect 1334 395 1340 396
rect 1326 387 1332 388
rect 1326 383 1327 387
rect 1331 383 1332 387
rect 1326 382 1332 383
rect 1336 379 1338 395
rect 1408 388 1410 406
rect 1414 400 1420 401
rect 1414 396 1415 400
rect 1419 396 1420 400
rect 1414 395 1420 396
rect 1406 387 1412 388
rect 1406 383 1407 387
rect 1411 383 1412 387
rect 1406 382 1412 383
rect 1416 379 1418 395
rect 1496 388 1498 406
rect 1502 400 1508 401
rect 1502 396 1503 400
rect 1507 396 1508 400
rect 1502 395 1508 396
rect 1494 387 1500 388
rect 1494 383 1495 387
rect 1499 383 1500 387
rect 1494 382 1500 383
rect 1504 379 1506 395
rect 1512 380 1514 406
rect 1584 388 1586 450
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1702 440 1708 441
rect 1702 436 1703 440
rect 1707 436 1708 440
rect 1702 435 1708 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1591 434 1595 435
rect 1591 429 1595 430
rect 1599 434 1603 435
rect 1599 429 1603 430
rect 1671 434 1675 435
rect 1671 429 1675 430
rect 1703 434 1707 435
rect 1703 429 1707 430
rect 1751 434 1755 435
rect 1751 429 1755 430
rect 1799 434 1803 435
rect 1799 429 1803 430
rect 1823 434 1827 435
rect 1823 429 1827 430
rect 1590 428 1596 429
rect 1590 424 1591 428
rect 1595 424 1596 428
rect 1590 423 1596 424
rect 1670 428 1676 429
rect 1670 424 1671 428
rect 1675 424 1676 428
rect 1670 423 1676 424
rect 1750 428 1756 429
rect 1750 424 1751 428
rect 1755 424 1756 428
rect 1750 423 1756 424
rect 1822 428 1828 429
rect 1822 424 1823 428
rect 1827 424 1828 428
rect 1822 423 1828 424
rect 1848 412 1850 466
rect 1886 464 1887 468
rect 1891 464 1892 468
rect 1886 463 1892 464
rect 1916 456 1918 474
rect 1968 456 1970 486
rect 1983 481 1987 482
rect 2007 481 2011 482
rect 2071 481 2075 482
rect 1984 469 1986 481
rect 2072 469 2074 481
rect 2080 480 2082 510
rect 2118 508 2119 512
rect 2123 508 2124 512
rect 2118 507 2124 508
rect 2120 487 2122 507
rect 2119 486 2123 487
rect 2119 481 2123 482
rect 2078 479 2084 480
rect 2078 475 2079 479
rect 2083 475 2084 479
rect 2078 474 2084 475
rect 1982 468 1988 469
rect 1982 464 1983 468
rect 1987 464 1988 468
rect 1982 463 1988 464
rect 2070 468 2076 469
rect 2070 464 2071 468
rect 2075 464 2076 468
rect 2070 463 2076 464
rect 2120 461 2122 481
rect 2118 460 2124 461
rect 2118 456 2119 460
rect 2123 456 2124 460
rect 1914 455 1920 456
rect 1914 451 1915 455
rect 1919 451 1920 455
rect 1914 450 1920 451
rect 1966 455 1972 456
rect 1966 451 1967 455
rect 1971 451 1972 455
rect 1966 450 1972 451
rect 2030 455 2036 456
rect 2118 455 2124 456
rect 2030 451 2031 455
rect 2035 451 2036 455
rect 2030 450 2036 451
rect 1886 440 1892 441
rect 1886 436 1887 440
rect 1891 436 1892 440
rect 1886 435 1892 436
rect 1982 440 1988 441
rect 1982 436 1983 440
rect 1987 436 1988 440
rect 1982 435 1988 436
rect 1887 434 1891 435
rect 1887 429 1891 430
rect 1951 434 1955 435
rect 1951 429 1955 430
rect 1983 434 1987 435
rect 1983 429 1987 430
rect 2023 434 2027 435
rect 2023 429 2027 430
rect 1886 428 1892 429
rect 1886 424 1887 428
rect 1891 424 1892 428
rect 1886 423 1892 424
rect 1950 428 1956 429
rect 1950 424 1951 428
rect 1955 424 1956 428
rect 1950 423 1956 424
rect 2022 428 2028 429
rect 2022 424 2023 428
rect 2027 424 2028 428
rect 2022 423 2028 424
rect 1662 411 1668 412
rect 1662 407 1663 411
rect 1667 407 1668 411
rect 1662 406 1668 407
rect 1742 411 1748 412
rect 1742 407 1743 411
rect 1747 407 1748 411
rect 1742 406 1748 407
rect 1814 411 1820 412
rect 1814 407 1815 411
rect 1819 407 1820 411
rect 1814 406 1820 407
rect 1846 411 1852 412
rect 1846 407 1847 411
rect 1851 407 1852 411
rect 1846 406 1852 407
rect 1922 411 1928 412
rect 1922 407 1923 411
rect 1927 407 1928 411
rect 1922 406 1928 407
rect 1590 400 1596 401
rect 1590 396 1591 400
rect 1595 396 1596 400
rect 1590 395 1596 396
rect 1582 387 1588 388
rect 1582 383 1583 387
rect 1587 383 1588 387
rect 1582 382 1588 383
rect 1510 379 1516 380
rect 1592 379 1594 395
rect 1664 388 1666 406
rect 1670 400 1676 401
rect 1670 396 1671 400
rect 1675 396 1676 400
rect 1670 395 1676 396
rect 1662 387 1668 388
rect 1662 383 1663 387
rect 1667 383 1668 387
rect 1662 382 1668 383
rect 1672 379 1674 395
rect 1744 388 1746 406
rect 1750 400 1756 401
rect 1750 396 1751 400
rect 1755 396 1756 400
rect 1750 395 1756 396
rect 1742 387 1748 388
rect 1742 383 1743 387
rect 1747 383 1748 387
rect 1742 382 1748 383
rect 1752 379 1754 395
rect 399 378 403 379
rect 399 373 403 374
rect 423 378 427 379
rect 423 373 427 374
rect 463 378 467 379
rect 463 373 467 374
rect 487 378 491 379
rect 494 378 500 379
rect 519 378 523 379
rect 542 378 548 379
rect 551 378 555 379
rect 487 373 491 374
rect 519 373 523 374
rect 390 371 396 372
rect 390 367 391 371
rect 395 367 396 371
rect 390 366 396 367
rect 400 361 402 373
rect 410 371 416 372
rect 410 367 411 371
rect 415 367 416 371
rect 410 366 416 367
rect 334 360 340 361
rect 334 356 335 360
rect 339 356 340 360
rect 334 355 340 356
rect 398 360 404 361
rect 398 356 399 360
rect 403 356 404 360
rect 398 355 404 356
rect 110 347 116 348
rect 142 347 148 348
rect 142 343 143 347
rect 147 343 148 347
rect 142 342 148 343
rect 242 347 248 348
rect 242 343 243 347
rect 247 343 248 347
rect 242 342 248 343
rect 298 347 304 348
rect 298 343 299 347
rect 303 343 304 347
rect 298 342 304 343
rect 370 347 376 348
rect 370 343 371 347
rect 375 343 376 347
rect 370 342 376 343
rect 110 335 116 336
rect 110 331 111 335
rect 115 331 116 335
rect 110 330 116 331
rect 134 332 140 333
rect 112 323 114 330
rect 134 328 135 332
rect 139 328 140 332
rect 134 327 140 328
rect 136 323 138 327
rect 111 322 115 323
rect 111 317 115 318
rect 135 322 139 323
rect 135 317 139 318
rect 112 314 114 317
rect 134 316 140 317
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 134 312 135 316
rect 139 312 140 316
rect 134 311 140 312
rect 110 308 116 309
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 112 271 114 291
rect 134 288 140 289
rect 134 284 135 288
rect 139 284 140 288
rect 134 283 140 284
rect 136 271 138 283
rect 144 276 146 342
rect 174 332 180 333
rect 174 328 175 332
rect 179 328 180 332
rect 174 327 180 328
rect 214 332 220 333
rect 214 328 215 332
rect 219 328 220 332
rect 214 327 220 328
rect 270 332 276 333
rect 270 328 271 332
rect 275 328 276 332
rect 270 327 276 328
rect 334 332 340 333
rect 334 328 335 332
rect 339 328 340 332
rect 334 327 340 328
rect 176 323 178 327
rect 216 323 218 327
rect 272 323 274 327
rect 336 323 338 327
rect 372 324 374 342
rect 398 332 404 333
rect 398 328 399 332
rect 403 328 404 332
rect 398 327 404 328
rect 370 323 376 324
rect 400 323 402 327
rect 175 322 179 323
rect 175 317 179 318
rect 207 322 211 323
rect 207 317 211 318
rect 215 322 219 323
rect 215 317 219 318
rect 271 322 275 323
rect 271 317 275 318
rect 295 322 299 323
rect 295 317 299 318
rect 335 322 339 323
rect 370 319 371 323
rect 375 319 376 323
rect 370 318 376 319
rect 383 322 387 323
rect 335 317 339 318
rect 383 317 387 318
rect 399 322 403 323
rect 399 317 403 318
rect 206 316 212 317
rect 206 312 207 316
rect 211 312 212 316
rect 206 311 212 312
rect 294 316 300 317
rect 294 312 295 316
rect 299 312 300 316
rect 294 311 300 312
rect 382 316 388 317
rect 382 312 383 316
rect 387 312 388 316
rect 382 311 388 312
rect 412 300 414 366
rect 464 361 466 373
rect 498 371 504 372
rect 498 367 499 371
rect 503 367 504 371
rect 498 366 504 367
rect 462 360 468 361
rect 462 356 463 360
rect 467 356 468 360
rect 462 355 468 356
rect 500 348 502 366
rect 520 361 522 373
rect 518 360 524 361
rect 518 356 519 360
rect 523 356 524 360
rect 518 355 524 356
rect 544 348 546 378
rect 551 373 555 374
rect 575 378 579 379
rect 602 378 608 379
rect 615 378 619 379
rect 575 373 579 374
rect 576 361 578 373
rect 574 360 580 361
rect 574 356 575 360
rect 579 356 580 360
rect 574 355 580 356
rect 604 348 606 378
rect 615 373 619 374
rect 631 378 635 379
rect 662 378 668 379
rect 671 378 675 379
rect 631 373 635 374
rect 671 373 675 374
rect 687 378 691 379
rect 718 378 724 379
rect 727 378 731 379
rect 687 373 691 374
rect 727 373 731 374
rect 751 378 755 379
rect 782 378 788 379
rect 791 378 795 379
rect 846 378 852 379
rect 855 378 859 379
rect 751 373 755 374
rect 791 373 795 374
rect 855 373 859 374
rect 1095 378 1099 379
rect 1095 373 1099 374
rect 1135 378 1139 379
rect 1135 373 1139 374
rect 1159 378 1163 379
rect 1159 373 1163 374
rect 1199 378 1203 379
rect 1199 373 1203 374
rect 1255 378 1259 379
rect 1255 373 1259 374
rect 1303 378 1307 379
rect 1303 373 1307 374
rect 1335 378 1339 379
rect 1335 373 1339 374
rect 1343 378 1347 379
rect 1343 373 1347 374
rect 1383 378 1387 379
rect 1383 373 1387 374
rect 1415 378 1419 379
rect 1415 373 1419 374
rect 1423 378 1427 379
rect 1423 373 1427 374
rect 1463 378 1467 379
rect 1463 373 1467 374
rect 1503 378 1507 379
rect 1510 375 1511 379
rect 1515 375 1516 379
rect 1510 374 1516 375
rect 1551 378 1555 379
rect 1503 373 1507 374
rect 1551 373 1555 374
rect 1591 378 1595 379
rect 1591 373 1595 374
rect 1615 378 1619 379
rect 1615 373 1619 374
rect 1671 378 1675 379
rect 1671 373 1675 374
rect 1679 378 1683 379
rect 1679 373 1683 374
rect 1751 378 1755 379
rect 1751 373 1755 374
rect 632 361 634 373
rect 646 371 652 372
rect 646 367 647 371
rect 651 367 652 371
rect 646 366 652 367
rect 658 371 664 372
rect 658 367 659 371
rect 663 367 664 371
rect 658 366 664 367
rect 630 360 636 361
rect 630 356 631 360
rect 635 356 636 360
rect 630 355 636 356
rect 498 347 504 348
rect 498 343 499 347
rect 503 343 504 347
rect 498 342 504 343
rect 542 347 548 348
rect 542 343 543 347
rect 547 343 548 347
rect 542 342 548 343
rect 602 347 608 348
rect 602 343 603 347
rect 607 343 608 347
rect 602 342 608 343
rect 462 332 468 333
rect 462 328 463 332
rect 467 328 468 332
rect 462 327 468 328
rect 518 332 524 333
rect 518 328 519 332
rect 523 328 524 332
rect 518 327 524 328
rect 574 332 580 333
rect 574 328 575 332
rect 579 328 580 332
rect 574 327 580 328
rect 630 332 636 333
rect 630 328 631 332
rect 635 328 636 332
rect 630 327 636 328
rect 464 323 466 327
rect 520 323 522 327
rect 576 323 578 327
rect 632 323 634 327
rect 463 322 467 323
rect 463 317 467 318
rect 471 322 475 323
rect 471 317 475 318
rect 519 322 523 323
rect 519 317 523 318
rect 551 322 555 323
rect 551 317 555 318
rect 575 322 579 323
rect 575 317 579 318
rect 623 322 627 323
rect 623 317 627 318
rect 631 322 635 323
rect 631 317 635 318
rect 470 316 476 317
rect 470 312 471 316
rect 475 312 476 316
rect 470 311 476 312
rect 550 316 556 317
rect 550 312 551 316
rect 555 312 556 316
rect 550 311 556 312
rect 622 316 628 317
rect 622 312 623 316
rect 627 312 628 316
rect 622 311 628 312
rect 648 300 650 366
rect 660 348 662 366
rect 688 361 690 373
rect 714 371 720 372
rect 714 367 715 371
rect 719 367 720 371
rect 714 366 720 367
rect 686 360 692 361
rect 686 356 687 360
rect 691 356 692 360
rect 686 355 692 356
rect 716 348 718 366
rect 752 361 754 373
rect 750 360 756 361
rect 750 356 751 360
rect 755 356 756 360
rect 750 355 756 356
rect 1096 353 1098 373
rect 1136 353 1138 373
rect 1304 361 1306 373
rect 1326 371 1332 372
rect 1326 367 1327 371
rect 1331 367 1332 371
rect 1326 366 1332 367
rect 1302 360 1308 361
rect 1302 356 1303 360
rect 1307 356 1308 360
rect 1302 355 1308 356
rect 1094 352 1100 353
rect 1094 348 1095 352
rect 1099 348 1100 352
rect 658 347 664 348
rect 658 343 659 347
rect 663 343 664 347
rect 658 342 664 343
rect 714 347 720 348
rect 1094 347 1100 348
rect 1134 352 1140 353
rect 1134 348 1135 352
rect 1139 348 1140 352
rect 1328 348 1330 366
rect 1344 361 1346 373
rect 1370 371 1376 372
rect 1370 367 1371 371
rect 1375 367 1376 371
rect 1370 366 1376 367
rect 1342 360 1348 361
rect 1342 356 1343 360
rect 1347 356 1348 360
rect 1342 355 1348 356
rect 1372 348 1374 366
rect 1384 361 1386 373
rect 1406 371 1412 372
rect 1406 367 1407 371
rect 1411 367 1412 371
rect 1406 366 1412 367
rect 1382 360 1388 361
rect 1382 356 1383 360
rect 1387 356 1388 360
rect 1382 355 1388 356
rect 1408 348 1410 366
rect 1424 361 1426 373
rect 1450 371 1456 372
rect 1450 367 1451 371
rect 1455 367 1456 371
rect 1450 366 1456 367
rect 1422 360 1428 361
rect 1422 356 1423 360
rect 1427 356 1428 360
rect 1422 355 1428 356
rect 1452 348 1454 366
rect 1464 361 1466 373
rect 1490 371 1496 372
rect 1490 367 1491 371
rect 1495 367 1496 371
rect 1490 366 1496 367
rect 1462 360 1468 361
rect 1462 356 1463 360
rect 1467 356 1468 360
rect 1462 355 1468 356
rect 1492 348 1494 366
rect 1504 361 1506 373
rect 1552 361 1554 373
rect 1570 371 1576 372
rect 1570 367 1571 371
rect 1575 367 1576 371
rect 1570 366 1576 367
rect 1578 371 1584 372
rect 1578 367 1579 371
rect 1583 367 1584 371
rect 1578 366 1584 367
rect 1502 360 1508 361
rect 1502 356 1503 360
rect 1507 356 1508 360
rect 1502 355 1508 356
rect 1550 360 1556 361
rect 1550 356 1551 360
rect 1555 356 1556 360
rect 1550 355 1556 356
rect 1134 347 1140 348
rect 1326 347 1332 348
rect 714 343 715 347
rect 719 343 720 347
rect 714 342 720 343
rect 1326 343 1327 347
rect 1331 343 1332 347
rect 1326 342 1332 343
rect 1370 347 1376 348
rect 1370 343 1371 347
rect 1375 343 1376 347
rect 1370 342 1376 343
rect 1406 347 1412 348
rect 1406 343 1407 347
rect 1411 343 1412 347
rect 1406 342 1412 343
rect 1450 347 1456 348
rect 1450 343 1451 347
rect 1455 343 1456 347
rect 1450 342 1456 343
rect 1490 347 1496 348
rect 1490 343 1491 347
rect 1495 343 1496 347
rect 1490 342 1496 343
rect 1542 347 1548 348
rect 1542 343 1543 347
rect 1547 343 1548 347
rect 1542 342 1548 343
rect 1094 335 1100 336
rect 686 332 692 333
rect 686 328 687 332
rect 691 328 692 332
rect 686 327 692 328
rect 750 332 756 333
rect 750 328 751 332
rect 755 328 756 332
rect 1094 331 1095 335
rect 1099 331 1100 335
rect 1094 330 1100 331
rect 1134 335 1140 336
rect 1134 331 1135 335
rect 1139 331 1140 335
rect 1134 330 1140 331
rect 1302 332 1308 333
rect 750 327 756 328
rect 688 323 690 327
rect 752 323 754 327
rect 1096 323 1098 330
rect 1136 323 1138 330
rect 1302 328 1303 332
rect 1307 328 1308 332
rect 1302 327 1308 328
rect 1342 332 1348 333
rect 1342 328 1343 332
rect 1347 328 1348 332
rect 1342 327 1348 328
rect 1382 332 1388 333
rect 1382 328 1383 332
rect 1387 328 1388 332
rect 1382 327 1388 328
rect 1422 332 1428 333
rect 1422 328 1423 332
rect 1427 328 1428 332
rect 1422 327 1428 328
rect 1462 332 1468 333
rect 1462 328 1463 332
rect 1467 328 1468 332
rect 1462 327 1468 328
rect 1502 332 1508 333
rect 1502 328 1503 332
rect 1507 328 1508 332
rect 1502 327 1508 328
rect 1304 323 1306 327
rect 1344 323 1346 327
rect 1384 323 1386 327
rect 1424 323 1426 327
rect 1464 323 1466 327
rect 1504 323 1506 327
rect 687 322 691 323
rect 687 317 691 318
rect 751 322 755 323
rect 751 317 755 318
rect 807 322 811 323
rect 807 317 811 318
rect 871 322 875 323
rect 871 317 875 318
rect 935 322 939 323
rect 935 317 939 318
rect 1095 322 1099 323
rect 1095 317 1099 318
rect 1135 322 1139 323
rect 1135 317 1139 318
rect 1167 322 1171 323
rect 1167 317 1171 318
rect 1207 322 1211 323
rect 1207 317 1211 318
rect 1247 322 1251 323
rect 1247 317 1251 318
rect 1295 322 1299 323
rect 1295 317 1299 318
rect 1303 322 1307 323
rect 1303 317 1307 318
rect 1343 322 1347 323
rect 1343 317 1347 318
rect 1383 322 1387 323
rect 1383 317 1387 318
rect 1391 322 1395 323
rect 1391 317 1395 318
rect 1423 322 1427 323
rect 1423 317 1427 318
rect 1439 322 1443 323
rect 1439 317 1443 318
rect 1463 322 1467 323
rect 1463 317 1467 318
rect 1495 322 1499 323
rect 1495 317 1499 318
rect 1503 322 1507 323
rect 1503 317 1507 318
rect 686 316 692 317
rect 686 312 687 316
rect 691 312 692 316
rect 686 311 692 312
rect 750 316 756 317
rect 750 312 751 316
rect 755 312 756 316
rect 750 311 756 312
rect 806 316 812 317
rect 806 312 807 316
rect 811 312 812 316
rect 806 311 812 312
rect 870 316 876 317
rect 870 312 871 316
rect 875 312 876 316
rect 870 311 876 312
rect 934 316 940 317
rect 934 312 935 316
rect 939 312 940 316
rect 1096 314 1098 317
rect 1136 314 1138 317
rect 1166 316 1172 317
rect 934 311 940 312
rect 1094 313 1100 314
rect 1094 309 1095 313
rect 1099 309 1100 313
rect 1094 308 1100 309
rect 1134 313 1140 314
rect 1134 309 1135 313
rect 1139 309 1140 313
rect 1166 312 1167 316
rect 1171 312 1172 316
rect 1166 311 1172 312
rect 1206 316 1212 317
rect 1206 312 1207 316
rect 1211 312 1212 316
rect 1206 311 1212 312
rect 1246 316 1252 317
rect 1246 312 1247 316
rect 1251 312 1252 316
rect 1246 311 1252 312
rect 1294 316 1300 317
rect 1294 312 1295 316
rect 1299 312 1300 316
rect 1294 311 1300 312
rect 1342 316 1348 317
rect 1342 312 1343 316
rect 1347 312 1348 316
rect 1342 311 1348 312
rect 1390 316 1396 317
rect 1390 312 1391 316
rect 1395 312 1396 316
rect 1390 311 1396 312
rect 1438 316 1444 317
rect 1438 312 1439 316
rect 1443 312 1444 316
rect 1438 311 1444 312
rect 1494 316 1500 317
rect 1494 312 1495 316
rect 1499 312 1500 316
rect 1494 311 1500 312
rect 1134 308 1140 309
rect 1318 307 1324 308
rect 1318 303 1319 307
rect 1323 303 1324 307
rect 1318 302 1324 303
rect 1462 307 1468 308
rect 1462 303 1463 307
rect 1467 303 1468 307
rect 1462 302 1468 303
rect 286 299 292 300
rect 286 295 287 299
rect 291 295 292 299
rect 286 294 292 295
rect 302 299 308 300
rect 302 295 303 299
rect 307 295 308 299
rect 302 294 308 295
rect 410 299 416 300
rect 410 295 411 299
rect 415 295 416 299
rect 410 294 416 295
rect 418 299 424 300
rect 418 295 419 299
rect 423 295 424 299
rect 418 294 424 295
rect 646 299 652 300
rect 646 295 647 299
rect 651 295 652 299
rect 646 294 652 295
rect 722 299 728 300
rect 722 295 723 299
rect 727 295 728 299
rect 1174 299 1180 300
rect 722 294 728 295
rect 1094 296 1100 297
rect 206 288 212 289
rect 206 284 207 288
rect 211 284 212 288
rect 206 283 212 284
rect 142 275 148 276
rect 142 271 143 275
rect 147 271 148 275
rect 208 271 210 283
rect 288 276 290 294
rect 294 288 300 289
rect 294 284 295 288
rect 299 284 300 288
rect 294 283 300 284
rect 286 275 292 276
rect 286 271 287 275
rect 291 271 292 275
rect 296 271 298 283
rect 111 270 115 271
rect 111 265 115 266
rect 135 270 139 271
rect 142 270 148 271
rect 199 270 203 271
rect 135 265 139 266
rect 199 265 203 266
rect 207 270 211 271
rect 207 265 211 266
rect 279 270 283 271
rect 286 270 292 271
rect 295 270 299 271
rect 279 265 283 266
rect 295 265 299 266
rect 112 245 114 265
rect 136 253 138 265
rect 186 263 192 264
rect 186 259 187 263
rect 191 259 192 263
rect 186 258 192 259
rect 134 252 140 253
rect 134 248 135 252
rect 139 248 140 252
rect 134 247 140 248
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 188 240 190 258
rect 200 253 202 265
rect 266 263 272 264
rect 266 259 267 263
rect 271 259 272 263
rect 266 258 272 259
rect 198 252 204 253
rect 198 248 199 252
rect 203 248 204 252
rect 198 247 204 248
rect 268 240 270 258
rect 280 253 282 265
rect 304 264 306 294
rect 382 288 388 289
rect 382 284 383 288
rect 387 284 388 288
rect 382 283 388 284
rect 384 271 386 283
rect 420 276 422 294
rect 470 288 476 289
rect 470 284 471 288
rect 475 284 476 288
rect 470 283 476 284
rect 550 288 556 289
rect 550 284 551 288
rect 555 284 556 288
rect 550 283 556 284
rect 622 288 628 289
rect 622 284 623 288
rect 627 284 628 288
rect 622 283 628 284
rect 686 288 692 289
rect 686 284 687 288
rect 691 284 692 288
rect 686 283 692 284
rect 418 275 424 276
rect 418 271 419 275
rect 423 271 424 275
rect 472 271 474 283
rect 538 275 544 276
rect 538 271 539 275
rect 543 271 544 275
rect 552 271 554 283
rect 624 271 626 283
rect 688 271 690 283
rect 724 276 726 294
rect 1094 292 1095 296
rect 1099 292 1100 296
rect 1094 291 1100 292
rect 1134 296 1140 297
rect 1134 292 1135 296
rect 1139 292 1140 296
rect 1174 295 1175 299
rect 1179 295 1180 299
rect 1174 294 1180 295
rect 1134 291 1140 292
rect 750 288 756 289
rect 750 284 751 288
rect 755 284 756 288
rect 750 283 756 284
rect 806 288 812 289
rect 806 284 807 288
rect 811 284 812 288
rect 806 283 812 284
rect 870 288 876 289
rect 870 284 871 288
rect 875 284 876 288
rect 870 283 876 284
rect 934 288 940 289
rect 934 284 935 288
rect 939 284 940 288
rect 934 283 940 284
rect 722 275 728 276
rect 722 271 723 275
rect 727 271 728 275
rect 752 271 754 283
rect 808 271 810 283
rect 872 271 874 283
rect 906 275 912 276
rect 906 271 907 275
rect 911 271 912 275
rect 936 271 938 283
rect 1096 271 1098 291
rect 359 270 363 271
rect 359 265 363 266
rect 383 270 387 271
rect 418 270 424 271
rect 439 270 443 271
rect 383 265 387 266
rect 439 265 443 266
rect 471 270 475 271
rect 471 265 475 266
rect 511 270 515 271
rect 538 270 544 271
rect 551 270 555 271
rect 511 265 515 266
rect 302 263 308 264
rect 302 259 303 263
rect 307 259 308 263
rect 302 258 308 259
rect 350 263 356 264
rect 350 259 351 263
rect 355 259 356 263
rect 350 258 356 259
rect 278 252 284 253
rect 278 248 279 252
rect 283 248 284 252
rect 278 247 284 248
rect 110 239 116 240
rect 142 239 148 240
rect 142 235 143 239
rect 147 235 148 239
rect 142 234 148 235
rect 186 239 192 240
rect 186 235 187 239
rect 191 235 192 239
rect 186 234 192 235
rect 266 239 272 240
rect 266 235 267 239
rect 271 235 272 239
rect 266 234 272 235
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 134 224 140 225
rect 112 215 114 222
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 136 215 138 219
rect 111 214 115 215
rect 111 209 115 210
rect 135 214 139 215
rect 135 209 139 210
rect 112 206 114 209
rect 134 208 140 209
rect 110 205 116 206
rect 110 201 111 205
rect 115 201 116 205
rect 134 204 135 208
rect 139 204 140 208
rect 134 203 140 204
rect 110 200 116 201
rect 110 188 116 189
rect 110 184 111 188
rect 115 184 116 188
rect 110 183 116 184
rect 112 139 114 183
rect 134 180 140 181
rect 134 176 135 180
rect 139 176 140 180
rect 134 175 140 176
rect 136 139 138 175
rect 144 168 146 234
rect 198 224 204 225
rect 198 220 199 224
rect 203 220 204 224
rect 198 219 204 220
rect 278 224 284 225
rect 278 220 279 224
rect 283 220 284 224
rect 278 219 284 220
rect 200 215 202 219
rect 280 215 282 219
rect 183 214 187 215
rect 183 209 187 210
rect 199 214 203 215
rect 199 209 203 210
rect 231 214 235 215
rect 231 209 235 210
rect 279 214 283 215
rect 279 209 283 210
rect 327 214 331 215
rect 327 209 331 210
rect 182 208 188 209
rect 182 204 183 208
rect 187 204 188 208
rect 182 203 188 204
rect 230 208 236 209
rect 230 204 231 208
rect 235 204 236 208
rect 230 203 236 204
rect 278 208 284 209
rect 278 204 279 208
rect 283 204 284 208
rect 278 203 284 204
rect 326 208 332 209
rect 326 204 327 208
rect 331 204 332 208
rect 326 203 332 204
rect 352 192 354 258
rect 360 253 362 265
rect 390 263 396 264
rect 390 259 391 263
rect 395 259 396 263
rect 390 258 396 259
rect 358 252 364 253
rect 358 248 359 252
rect 363 248 364 252
rect 358 247 364 248
rect 392 240 394 258
rect 440 253 442 265
rect 512 253 514 265
rect 438 252 444 253
rect 438 248 439 252
rect 443 248 444 252
rect 438 247 444 248
rect 510 252 516 253
rect 510 248 511 252
rect 515 248 516 252
rect 510 247 516 248
rect 540 240 542 270
rect 551 265 555 266
rect 583 270 587 271
rect 583 265 587 266
rect 623 270 627 271
rect 623 265 627 266
rect 647 270 651 271
rect 647 265 651 266
rect 687 270 691 271
rect 687 265 691 266
rect 703 270 707 271
rect 722 270 728 271
rect 751 270 755 271
rect 703 265 707 266
rect 751 265 755 266
rect 759 270 763 271
rect 759 265 763 266
rect 807 270 811 271
rect 807 265 811 266
rect 815 270 819 271
rect 815 265 819 266
rect 871 270 875 271
rect 871 265 875 266
rect 879 270 883 271
rect 906 270 912 271
rect 935 270 939 271
rect 879 265 883 266
rect 584 253 586 265
rect 590 263 596 264
rect 590 259 591 263
rect 595 259 596 263
rect 590 258 596 259
rect 610 263 616 264
rect 610 259 611 263
rect 615 259 616 263
rect 610 258 616 259
rect 582 252 588 253
rect 582 248 583 252
rect 587 248 588 252
rect 582 247 588 248
rect 386 239 394 240
rect 386 235 387 239
rect 391 236 394 239
rect 538 239 544 240
rect 391 235 392 236
rect 386 234 392 235
rect 538 235 539 239
rect 543 235 544 239
rect 538 234 544 235
rect 358 224 364 225
rect 358 220 359 224
rect 363 220 364 224
rect 358 219 364 220
rect 438 224 444 225
rect 438 220 439 224
rect 443 220 444 224
rect 438 219 444 220
rect 510 224 516 225
rect 510 220 511 224
rect 515 220 516 224
rect 510 219 516 220
rect 582 224 588 225
rect 582 220 583 224
rect 587 220 588 224
rect 582 219 588 220
rect 360 215 362 219
rect 440 215 442 219
rect 512 215 514 219
rect 584 215 586 219
rect 359 214 363 215
rect 359 209 363 210
rect 375 214 379 215
rect 375 209 379 210
rect 415 214 419 215
rect 415 209 419 210
rect 439 214 443 215
rect 439 209 443 210
rect 455 214 459 215
rect 455 209 459 210
rect 503 214 507 215
rect 503 209 507 210
rect 511 214 515 215
rect 511 209 515 210
rect 551 214 555 215
rect 551 209 555 210
rect 583 214 587 215
rect 583 209 587 210
rect 374 208 380 209
rect 374 204 375 208
rect 379 204 380 208
rect 374 203 380 204
rect 414 208 420 209
rect 414 204 415 208
rect 419 204 420 208
rect 414 203 420 204
rect 454 208 460 209
rect 454 204 455 208
rect 459 204 460 208
rect 454 203 460 204
rect 502 208 508 209
rect 502 204 503 208
rect 507 204 508 208
rect 502 203 508 204
rect 550 208 556 209
rect 550 204 551 208
rect 555 204 556 208
rect 550 203 556 204
rect 592 200 594 258
rect 612 240 614 258
rect 648 253 650 265
rect 704 253 706 265
rect 730 263 736 264
rect 730 259 731 263
rect 735 259 736 263
rect 730 258 736 259
rect 646 252 652 253
rect 646 248 647 252
rect 651 248 652 252
rect 646 247 652 248
rect 702 252 708 253
rect 702 248 703 252
rect 707 248 708 252
rect 702 247 708 248
rect 732 240 734 258
rect 760 253 762 265
rect 786 263 792 264
rect 786 259 787 263
rect 791 259 792 263
rect 786 258 792 259
rect 758 252 764 253
rect 758 248 759 252
rect 763 248 764 252
rect 758 247 764 248
rect 788 240 790 258
rect 816 253 818 265
rect 842 263 848 264
rect 842 259 843 263
rect 847 259 848 263
rect 842 258 848 259
rect 814 252 820 253
rect 814 248 815 252
rect 819 248 820 252
rect 814 247 820 248
rect 844 240 846 258
rect 880 253 882 265
rect 878 252 884 253
rect 878 248 879 252
rect 883 248 884 252
rect 878 247 884 248
rect 908 240 910 270
rect 935 265 939 266
rect 1095 270 1099 271
rect 1095 265 1099 266
rect 1096 245 1098 265
rect 1136 263 1138 291
rect 1166 288 1172 289
rect 1166 284 1167 288
rect 1171 284 1172 288
rect 1166 283 1172 284
rect 1168 263 1170 283
rect 1135 262 1139 263
rect 1135 257 1139 258
rect 1159 262 1163 263
rect 1159 257 1163 258
rect 1167 262 1171 263
rect 1167 257 1171 258
rect 1094 244 1100 245
rect 1094 240 1095 244
rect 1099 240 1100 244
rect 610 239 616 240
rect 610 235 611 239
rect 615 235 616 239
rect 610 234 616 235
rect 730 239 736 240
rect 730 235 731 239
rect 735 235 736 239
rect 730 234 736 235
rect 786 239 792 240
rect 786 235 787 239
rect 791 235 792 239
rect 786 234 792 235
rect 842 239 848 240
rect 842 235 843 239
rect 847 235 848 239
rect 842 234 848 235
rect 906 239 912 240
rect 1094 239 1100 240
rect 906 235 907 239
rect 911 235 912 239
rect 1136 237 1138 257
rect 1160 245 1162 257
rect 1176 256 1178 294
rect 1206 288 1212 289
rect 1206 284 1207 288
rect 1211 284 1212 288
rect 1206 283 1212 284
rect 1246 288 1252 289
rect 1246 284 1247 288
rect 1251 284 1252 288
rect 1246 283 1252 284
rect 1294 288 1300 289
rect 1294 284 1295 288
rect 1299 284 1300 288
rect 1294 283 1300 284
rect 1208 263 1210 283
rect 1248 263 1250 283
rect 1296 263 1298 283
rect 1320 276 1322 302
rect 1382 299 1388 300
rect 1382 295 1383 299
rect 1387 295 1388 299
rect 1382 294 1388 295
rect 1342 288 1348 289
rect 1342 284 1343 288
rect 1347 284 1348 288
rect 1342 283 1348 284
rect 1318 275 1324 276
rect 1318 271 1319 275
rect 1323 271 1324 275
rect 1318 270 1324 271
rect 1344 263 1346 283
rect 1384 276 1386 294
rect 1390 288 1396 289
rect 1390 284 1391 288
rect 1395 284 1396 288
rect 1390 283 1396 284
rect 1438 288 1444 289
rect 1438 284 1439 288
rect 1443 284 1444 288
rect 1438 283 1444 284
rect 1350 275 1356 276
rect 1350 271 1351 275
rect 1355 271 1356 275
rect 1350 270 1356 271
rect 1382 275 1388 276
rect 1382 271 1383 275
rect 1387 271 1388 275
rect 1382 270 1388 271
rect 1207 262 1211 263
rect 1207 257 1211 258
rect 1247 262 1251 263
rect 1247 257 1251 258
rect 1271 262 1275 263
rect 1271 257 1275 258
rect 1295 262 1299 263
rect 1295 257 1299 258
rect 1327 262 1331 263
rect 1327 257 1331 258
rect 1343 262 1347 263
rect 1343 257 1347 258
rect 1174 255 1180 256
rect 1174 251 1175 255
rect 1179 251 1180 255
rect 1174 250 1180 251
rect 1186 255 1192 256
rect 1186 251 1187 255
rect 1191 251 1192 255
rect 1186 250 1192 251
rect 1158 244 1164 245
rect 1158 240 1159 244
rect 1163 240 1164 244
rect 1158 239 1164 240
rect 906 234 912 235
rect 1134 236 1140 237
rect 1134 232 1135 236
rect 1139 232 1140 236
rect 1188 232 1190 250
rect 1208 245 1210 257
rect 1234 255 1240 256
rect 1234 251 1235 255
rect 1239 251 1240 255
rect 1234 250 1240 251
rect 1206 244 1212 245
rect 1206 240 1207 244
rect 1211 240 1212 244
rect 1206 239 1212 240
rect 1236 232 1238 250
rect 1272 245 1274 257
rect 1328 245 1330 257
rect 1270 244 1276 245
rect 1270 240 1271 244
rect 1275 240 1276 244
rect 1270 239 1276 240
rect 1326 244 1332 245
rect 1326 240 1327 244
rect 1331 240 1332 244
rect 1326 239 1332 240
rect 1352 232 1354 270
rect 1392 263 1394 283
rect 1440 263 1442 283
rect 1464 276 1466 302
rect 1486 299 1492 300
rect 1486 295 1487 299
rect 1491 295 1492 299
rect 1486 294 1492 295
rect 1518 299 1524 300
rect 1518 295 1519 299
rect 1523 295 1524 299
rect 1518 294 1524 295
rect 1488 276 1490 294
rect 1494 288 1500 289
rect 1494 284 1495 288
rect 1499 284 1500 288
rect 1494 283 1500 284
rect 1462 275 1468 276
rect 1462 271 1463 275
rect 1467 271 1468 275
rect 1462 270 1468 271
rect 1486 275 1492 276
rect 1486 271 1487 275
rect 1491 271 1492 275
rect 1486 270 1492 271
rect 1496 263 1498 283
rect 1391 262 1395 263
rect 1391 257 1395 258
rect 1439 262 1443 263
rect 1439 257 1443 258
rect 1455 262 1459 263
rect 1455 257 1459 258
rect 1495 262 1499 263
rect 1495 257 1499 258
rect 1378 255 1384 256
rect 1378 251 1379 255
rect 1383 251 1384 255
rect 1378 250 1384 251
rect 1380 232 1382 250
rect 1392 245 1394 257
rect 1422 255 1428 256
rect 1422 251 1423 255
rect 1427 251 1428 255
rect 1422 250 1428 251
rect 1390 244 1396 245
rect 1390 240 1391 244
rect 1395 240 1396 244
rect 1390 239 1396 240
rect 1134 231 1140 232
rect 1186 231 1192 232
rect 1094 227 1100 228
rect 646 224 652 225
rect 646 220 647 224
rect 651 220 652 224
rect 646 219 652 220
rect 702 224 708 225
rect 702 220 703 224
rect 707 220 708 224
rect 702 219 708 220
rect 758 224 764 225
rect 758 220 759 224
rect 763 220 764 224
rect 758 219 764 220
rect 814 224 820 225
rect 814 220 815 224
rect 819 220 820 224
rect 814 219 820 220
rect 878 224 884 225
rect 878 220 879 224
rect 883 220 884 224
rect 1094 223 1095 227
rect 1099 223 1100 227
rect 1186 227 1187 231
rect 1191 227 1192 231
rect 1186 226 1192 227
rect 1234 231 1240 232
rect 1234 227 1235 231
rect 1239 227 1240 231
rect 1234 226 1240 227
rect 1278 231 1284 232
rect 1278 227 1279 231
rect 1283 227 1284 231
rect 1278 226 1284 227
rect 1350 231 1356 232
rect 1350 227 1351 231
rect 1355 227 1356 231
rect 1350 226 1356 227
rect 1378 231 1384 232
rect 1378 227 1379 231
rect 1383 227 1384 231
rect 1378 226 1384 227
rect 1094 222 1100 223
rect 878 219 884 220
rect 648 215 650 219
rect 704 215 706 219
rect 760 215 762 219
rect 816 215 818 219
rect 880 215 882 219
rect 1096 215 1098 222
rect 1134 219 1140 220
rect 1134 215 1135 219
rect 1139 215 1140 219
rect 599 214 603 215
rect 599 209 603 210
rect 647 214 651 215
rect 647 209 651 210
rect 695 214 699 215
rect 695 209 699 210
rect 703 214 707 215
rect 703 209 707 210
rect 743 214 747 215
rect 743 209 747 210
rect 759 214 763 215
rect 759 209 763 210
rect 815 214 819 215
rect 815 209 819 210
rect 879 214 883 215
rect 879 209 883 210
rect 1095 214 1099 215
rect 1134 214 1140 215
rect 1158 216 1164 217
rect 1136 211 1138 214
rect 1158 212 1159 216
rect 1163 212 1164 216
rect 1158 211 1164 212
rect 1206 216 1212 217
rect 1206 212 1207 216
rect 1211 212 1212 216
rect 1206 211 1212 212
rect 1270 216 1276 217
rect 1270 212 1271 216
rect 1275 212 1276 216
rect 1270 211 1276 212
rect 1095 209 1099 210
rect 1135 210 1139 211
rect 598 208 604 209
rect 598 204 599 208
rect 603 204 604 208
rect 598 203 604 204
rect 646 208 652 209
rect 646 204 647 208
rect 651 204 652 208
rect 646 203 652 204
rect 694 208 700 209
rect 694 204 695 208
rect 699 204 700 208
rect 694 203 700 204
rect 742 208 748 209
rect 742 204 743 208
rect 747 204 748 208
rect 1096 206 1098 209
rect 742 203 748 204
rect 1094 205 1100 206
rect 1135 205 1139 206
rect 1159 210 1163 211
rect 1159 205 1163 206
rect 1199 210 1203 211
rect 1199 205 1203 206
rect 1207 210 1211 211
rect 1207 205 1211 206
rect 1263 210 1267 211
rect 1263 205 1267 206
rect 1271 210 1275 211
rect 1271 205 1275 206
rect 1094 201 1095 205
rect 1099 201 1100 205
rect 1136 202 1138 205
rect 1158 204 1164 205
rect 1094 200 1100 201
rect 1134 201 1140 202
rect 590 199 596 200
rect 590 195 591 199
rect 595 195 596 199
rect 1134 197 1135 201
rect 1139 197 1140 201
rect 1158 200 1159 204
rect 1163 200 1164 204
rect 1158 199 1164 200
rect 1198 204 1204 205
rect 1198 200 1199 204
rect 1203 200 1204 204
rect 1198 199 1204 200
rect 1262 204 1268 205
rect 1262 200 1263 204
rect 1267 200 1268 204
rect 1262 199 1268 200
rect 1134 196 1140 197
rect 590 194 596 195
rect 174 191 180 192
rect 174 187 175 191
rect 179 187 180 191
rect 174 186 180 187
rect 222 191 228 192
rect 222 187 223 191
rect 227 187 228 191
rect 222 186 228 187
rect 270 191 276 192
rect 270 187 271 191
rect 275 187 276 191
rect 270 186 276 187
rect 286 191 292 192
rect 286 187 287 191
rect 291 187 292 191
rect 286 186 292 187
rect 350 191 356 192
rect 350 187 351 191
rect 355 187 356 191
rect 350 186 356 187
rect 494 191 500 192
rect 494 187 495 191
rect 499 187 500 191
rect 494 186 500 187
rect 542 191 548 192
rect 542 187 543 191
rect 547 187 548 191
rect 542 186 548 187
rect 590 191 596 192
rect 590 187 591 191
rect 595 187 596 191
rect 590 186 596 187
rect 638 191 644 192
rect 638 187 639 191
rect 643 187 644 191
rect 638 186 644 187
rect 686 191 692 192
rect 686 187 687 191
rect 691 187 692 191
rect 686 186 692 187
rect 734 191 740 192
rect 734 187 735 191
rect 739 187 740 191
rect 734 186 740 187
rect 1094 188 1100 189
rect 176 168 178 186
rect 182 180 188 181
rect 182 176 183 180
rect 187 176 188 180
rect 182 175 188 176
rect 142 167 148 168
rect 142 163 143 167
rect 147 163 148 167
rect 142 162 148 163
rect 174 167 180 168
rect 174 163 175 167
rect 179 163 180 167
rect 174 162 180 163
rect 184 139 186 175
rect 224 168 226 186
rect 230 180 236 181
rect 230 176 231 180
rect 235 176 236 180
rect 230 175 236 176
rect 222 167 228 168
rect 222 163 223 167
rect 227 163 228 167
rect 222 162 228 163
rect 232 139 234 175
rect 272 168 274 186
rect 278 180 284 181
rect 278 176 279 180
rect 283 176 284 180
rect 278 175 284 176
rect 270 167 276 168
rect 270 163 271 167
rect 275 163 276 167
rect 270 162 276 163
rect 280 139 282 175
rect 288 140 290 186
rect 326 180 332 181
rect 326 176 327 180
rect 331 176 332 180
rect 326 175 332 176
rect 374 180 380 181
rect 374 176 375 180
rect 379 176 380 180
rect 374 175 380 176
rect 414 180 420 181
rect 414 176 415 180
rect 419 176 420 180
rect 414 175 420 176
rect 454 180 460 181
rect 454 176 455 180
rect 459 176 460 180
rect 454 175 460 176
rect 286 139 292 140
rect 328 139 330 175
rect 376 139 378 175
rect 416 139 418 175
rect 456 139 458 175
rect 496 168 498 186
rect 502 180 508 181
rect 502 176 503 180
rect 507 176 508 180
rect 502 175 508 176
rect 494 167 500 168
rect 494 163 495 167
rect 499 163 500 167
rect 494 162 500 163
rect 504 139 506 175
rect 544 168 546 186
rect 550 180 556 181
rect 550 176 551 180
rect 555 176 556 180
rect 550 175 556 176
rect 542 167 548 168
rect 542 163 543 167
rect 547 163 548 167
rect 542 162 548 163
rect 526 151 532 152
rect 526 147 527 151
rect 531 147 532 151
rect 526 146 532 147
rect 111 138 115 139
rect 111 133 115 134
rect 135 138 139 139
rect 135 133 139 134
rect 143 138 147 139
rect 143 133 147 134
rect 183 138 187 139
rect 183 133 187 134
rect 223 138 227 139
rect 223 133 227 134
rect 231 138 235 139
rect 231 133 235 134
rect 263 138 267 139
rect 263 133 267 134
rect 279 138 283 139
rect 286 135 287 139
rect 291 135 292 139
rect 286 134 292 135
rect 303 138 307 139
rect 279 133 283 134
rect 303 133 307 134
rect 327 138 331 139
rect 327 133 331 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 383 138 387 139
rect 383 133 387 134
rect 415 138 419 139
rect 415 133 419 134
rect 423 138 427 139
rect 423 133 427 134
rect 455 138 459 139
rect 455 133 459 134
rect 463 138 467 139
rect 463 133 467 134
rect 503 138 507 139
rect 503 133 507 134
rect 112 113 114 133
rect 144 121 146 133
rect 170 131 176 132
rect 170 127 171 131
rect 175 127 176 131
rect 170 126 176 127
rect 142 120 148 121
rect 142 116 143 120
rect 147 116 148 120
rect 142 115 148 116
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 172 108 174 126
rect 184 121 186 133
rect 210 131 216 132
rect 210 127 211 131
rect 215 127 216 131
rect 210 126 216 127
rect 182 120 188 121
rect 182 116 183 120
rect 187 116 188 120
rect 182 115 188 116
rect 212 108 214 126
rect 224 121 226 133
rect 246 131 252 132
rect 246 127 247 131
rect 251 127 252 131
rect 246 126 252 127
rect 222 120 228 121
rect 222 116 223 120
rect 227 116 228 120
rect 222 115 228 116
rect 248 108 250 126
rect 264 121 266 133
rect 290 131 296 132
rect 290 127 291 131
rect 295 127 296 131
rect 290 126 296 127
rect 262 120 268 121
rect 262 116 263 120
rect 267 116 268 120
rect 262 115 268 116
rect 292 108 294 126
rect 304 121 306 133
rect 334 131 340 132
rect 334 127 335 131
rect 339 127 340 131
rect 334 126 340 127
rect 302 120 308 121
rect 302 116 303 120
rect 307 116 308 120
rect 302 115 308 116
rect 336 108 338 126
rect 344 121 346 133
rect 366 131 372 132
rect 366 127 367 131
rect 371 127 372 131
rect 366 126 372 127
rect 342 120 348 121
rect 342 116 343 120
rect 347 116 348 120
rect 342 115 348 116
rect 368 108 370 126
rect 384 121 386 133
rect 406 131 412 132
rect 406 127 407 131
rect 411 127 412 131
rect 406 126 412 127
rect 382 120 388 121
rect 382 116 383 120
rect 387 116 388 120
rect 382 115 388 116
rect 408 108 410 126
rect 424 121 426 133
rect 446 131 452 132
rect 446 127 447 131
rect 451 127 452 131
rect 446 126 452 127
rect 422 120 428 121
rect 422 116 423 120
rect 427 116 428 120
rect 422 115 428 116
rect 448 108 450 126
rect 464 121 466 133
rect 490 131 496 132
rect 490 127 491 131
rect 495 127 496 131
rect 490 126 496 127
rect 462 120 468 121
rect 462 116 463 120
rect 467 116 468 120
rect 462 115 468 116
rect 492 108 494 126
rect 504 121 506 133
rect 502 120 508 121
rect 502 116 503 120
rect 507 116 508 120
rect 502 115 508 116
rect 528 108 530 146
rect 552 139 554 175
rect 592 168 594 186
rect 598 180 604 181
rect 598 176 599 180
rect 603 176 604 180
rect 598 175 604 176
rect 590 167 596 168
rect 590 163 591 167
rect 595 163 596 167
rect 590 162 596 163
rect 566 159 572 160
rect 566 155 567 159
rect 571 155 572 159
rect 566 154 572 155
rect 543 138 547 139
rect 543 133 547 134
rect 551 138 555 139
rect 551 133 555 134
rect 544 121 546 133
rect 542 120 548 121
rect 542 116 543 120
rect 547 116 548 120
rect 542 115 548 116
rect 568 108 570 154
rect 600 139 602 175
rect 640 168 642 186
rect 646 180 652 181
rect 646 176 647 180
rect 651 176 652 180
rect 646 175 652 176
rect 638 167 644 168
rect 638 163 639 167
rect 643 163 644 167
rect 638 162 644 163
rect 648 139 650 175
rect 688 168 690 186
rect 694 180 700 181
rect 694 176 695 180
rect 699 176 700 180
rect 694 175 700 176
rect 686 167 692 168
rect 686 163 687 167
rect 691 163 692 167
rect 686 162 692 163
rect 696 139 698 175
rect 736 168 738 186
rect 1094 184 1095 188
rect 1099 184 1100 188
rect 1170 187 1176 188
rect 1094 183 1100 184
rect 1134 184 1140 185
rect 742 180 748 181
rect 742 176 743 180
rect 747 176 748 180
rect 742 175 748 176
rect 734 167 740 168
rect 734 163 735 167
rect 739 163 740 167
rect 734 162 740 163
rect 744 139 746 175
rect 1096 139 1098 183
rect 1134 180 1135 184
rect 1139 180 1140 184
rect 1170 183 1171 187
rect 1175 183 1176 187
rect 1170 182 1176 183
rect 1134 179 1140 180
rect 1136 139 1138 179
rect 1158 176 1164 177
rect 1158 172 1159 176
rect 1163 172 1164 176
rect 1158 171 1164 172
rect 1160 139 1162 171
rect 583 138 587 139
rect 583 133 587 134
rect 599 138 603 139
rect 599 133 603 134
rect 623 138 627 139
rect 623 133 627 134
rect 647 138 651 139
rect 647 133 651 134
rect 663 138 667 139
rect 663 133 667 134
rect 695 138 699 139
rect 695 133 699 134
rect 703 138 707 139
rect 703 133 707 134
rect 743 138 747 139
rect 743 133 747 134
rect 783 138 787 139
rect 783 133 787 134
rect 831 138 835 139
rect 831 133 835 134
rect 879 138 883 139
rect 879 133 883 134
rect 927 138 931 139
rect 927 133 931 134
rect 967 138 971 139
rect 967 133 971 134
rect 1007 138 1011 139
rect 1007 133 1011 134
rect 1047 138 1051 139
rect 1047 133 1051 134
rect 1095 138 1099 139
rect 1095 133 1099 134
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1159 138 1163 139
rect 1159 133 1163 134
rect 584 121 586 133
rect 624 121 626 133
rect 664 121 666 133
rect 704 121 706 133
rect 744 121 746 133
rect 784 121 786 133
rect 818 131 824 132
rect 818 127 819 131
rect 823 127 824 131
rect 818 126 824 127
rect 582 120 588 121
rect 582 116 583 120
rect 587 116 588 120
rect 582 115 588 116
rect 622 120 628 121
rect 622 116 623 120
rect 627 116 628 120
rect 622 115 628 116
rect 662 120 668 121
rect 662 116 663 120
rect 667 116 668 120
rect 662 115 668 116
rect 702 120 708 121
rect 702 116 703 120
rect 707 116 708 120
rect 702 115 708 116
rect 742 120 748 121
rect 742 116 743 120
rect 747 116 748 120
rect 742 115 748 116
rect 782 120 788 121
rect 782 116 783 120
rect 787 116 788 120
rect 782 115 788 116
rect 820 108 822 126
rect 832 121 834 133
rect 866 131 872 132
rect 866 127 867 131
rect 871 127 872 131
rect 866 126 872 127
rect 830 120 836 121
rect 830 116 831 120
rect 835 116 836 120
rect 830 115 836 116
rect 868 108 870 126
rect 880 121 882 133
rect 928 121 930 133
rect 968 121 970 133
rect 1008 121 1010 133
rect 1048 121 1050 133
rect 878 120 884 121
rect 878 116 879 120
rect 883 116 884 120
rect 878 115 884 116
rect 926 120 932 121
rect 926 116 927 120
rect 931 116 932 120
rect 926 115 932 116
rect 966 120 972 121
rect 966 116 967 120
rect 971 116 972 120
rect 966 115 972 116
rect 1006 120 1012 121
rect 1006 116 1007 120
rect 1011 116 1012 120
rect 1006 115 1012 116
rect 1046 120 1052 121
rect 1046 116 1047 120
rect 1051 116 1052 120
rect 1046 115 1052 116
rect 1096 113 1098 133
rect 1136 113 1138 133
rect 1142 131 1148 132
rect 1142 127 1143 131
rect 1147 127 1148 131
rect 1142 126 1148 127
rect 1094 112 1100 113
rect 1094 108 1095 112
rect 1099 108 1100 112
rect 110 107 116 108
rect 170 107 176 108
rect 170 103 171 107
rect 175 103 176 107
rect 170 102 176 103
rect 210 107 216 108
rect 210 103 211 107
rect 215 103 216 107
rect 210 102 216 103
rect 246 107 252 108
rect 246 103 247 107
rect 251 103 252 107
rect 246 102 252 103
rect 290 107 296 108
rect 290 103 291 107
rect 295 103 296 107
rect 290 102 296 103
rect 330 107 338 108
rect 330 103 331 107
rect 335 104 338 107
rect 366 107 372 108
rect 335 103 336 104
rect 330 102 336 103
rect 366 103 367 107
rect 371 103 372 107
rect 366 102 372 103
rect 406 107 412 108
rect 406 103 407 107
rect 411 103 412 107
rect 406 102 412 103
rect 446 107 452 108
rect 446 103 447 107
rect 451 103 452 107
rect 446 102 452 103
rect 490 107 496 108
rect 490 103 491 107
rect 495 103 496 107
rect 490 102 496 103
rect 526 107 532 108
rect 526 103 527 107
rect 531 103 532 107
rect 526 102 532 103
rect 566 107 572 108
rect 566 103 567 107
rect 571 103 572 107
rect 566 102 572 103
rect 818 107 824 108
rect 818 103 819 107
rect 823 103 824 107
rect 818 102 824 103
rect 866 107 872 108
rect 1094 107 1100 108
rect 1134 112 1140 113
rect 1134 108 1135 112
rect 1139 108 1140 112
rect 1144 108 1146 126
rect 1160 121 1162 133
rect 1172 132 1174 182
rect 1198 176 1204 177
rect 1198 172 1199 176
rect 1203 172 1204 176
rect 1198 171 1204 172
rect 1262 176 1268 177
rect 1262 172 1263 176
rect 1267 172 1268 176
rect 1262 171 1268 172
rect 1200 139 1202 171
rect 1264 139 1266 171
rect 1280 164 1282 226
rect 1326 216 1332 217
rect 1326 212 1327 216
rect 1331 212 1332 216
rect 1326 211 1332 212
rect 1390 216 1396 217
rect 1390 212 1391 216
rect 1395 212 1396 216
rect 1390 211 1396 212
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1391 210 1395 211
rect 1391 205 1395 206
rect 1399 210 1403 211
rect 1399 205 1403 206
rect 1326 204 1332 205
rect 1326 200 1327 204
rect 1331 200 1332 204
rect 1326 199 1332 200
rect 1398 204 1404 205
rect 1398 200 1399 204
rect 1403 200 1404 204
rect 1398 199 1404 200
rect 1424 188 1426 250
rect 1456 245 1458 257
rect 1520 256 1522 294
rect 1544 276 1546 342
rect 1550 332 1556 333
rect 1550 328 1551 332
rect 1555 328 1556 332
rect 1550 327 1556 328
rect 1552 323 1554 327
rect 1551 322 1555 323
rect 1551 317 1555 318
rect 1559 322 1563 323
rect 1559 317 1563 318
rect 1558 316 1564 317
rect 1558 312 1559 316
rect 1563 312 1564 316
rect 1558 311 1564 312
rect 1572 300 1574 366
rect 1580 348 1582 366
rect 1616 361 1618 373
rect 1642 371 1648 372
rect 1642 367 1643 371
rect 1647 367 1648 371
rect 1642 366 1648 367
rect 1614 360 1620 361
rect 1614 356 1615 360
rect 1619 356 1620 360
rect 1614 355 1620 356
rect 1644 348 1646 366
rect 1680 361 1682 373
rect 1706 371 1712 372
rect 1706 367 1707 371
rect 1711 367 1712 371
rect 1706 366 1712 367
rect 1678 360 1684 361
rect 1678 356 1679 360
rect 1683 356 1684 360
rect 1678 355 1684 356
rect 1708 348 1710 366
rect 1752 361 1754 373
rect 1816 372 1818 406
rect 1822 400 1828 401
rect 1822 396 1823 400
rect 1827 396 1828 400
rect 1822 395 1828 396
rect 1886 400 1892 401
rect 1886 396 1887 400
rect 1891 396 1892 400
rect 1886 395 1892 396
rect 1824 379 1826 395
rect 1888 379 1890 395
rect 1924 388 1926 406
rect 1950 400 1956 401
rect 1950 396 1951 400
rect 1955 396 1956 400
rect 1950 395 1956 396
rect 2022 400 2028 401
rect 2022 396 2023 400
rect 2027 396 2028 400
rect 2022 395 2028 396
rect 1922 387 1928 388
rect 1922 383 1923 387
rect 1927 383 1928 387
rect 1922 382 1928 383
rect 1952 379 1954 395
rect 1998 387 2004 388
rect 1998 383 1999 387
rect 2003 383 2004 387
rect 1998 382 2004 383
rect 1823 378 1827 379
rect 1823 373 1827 374
rect 1831 378 1835 379
rect 1831 373 1835 374
rect 1887 378 1891 379
rect 1887 373 1891 374
rect 1919 378 1923 379
rect 1919 373 1923 374
rect 1951 378 1955 379
rect 1951 373 1955 374
rect 1814 371 1820 372
rect 1814 367 1815 371
rect 1819 367 1820 371
rect 1814 366 1820 367
rect 1832 361 1834 373
rect 1920 361 1922 373
rect 1942 371 1948 372
rect 1942 367 1943 371
rect 1947 367 1948 371
rect 1942 366 1948 367
rect 1750 360 1756 361
rect 1750 356 1751 360
rect 1755 356 1756 360
rect 1750 355 1756 356
rect 1830 360 1836 361
rect 1830 356 1831 360
rect 1835 356 1836 360
rect 1830 355 1836 356
rect 1918 360 1924 361
rect 1918 356 1919 360
rect 1923 356 1924 360
rect 1918 355 1924 356
rect 1578 347 1584 348
rect 1578 343 1579 347
rect 1583 343 1584 347
rect 1578 342 1584 343
rect 1642 347 1648 348
rect 1642 343 1643 347
rect 1647 343 1648 347
rect 1642 342 1648 343
rect 1706 347 1712 348
rect 1706 343 1707 347
rect 1711 343 1712 347
rect 1706 342 1712 343
rect 1714 347 1720 348
rect 1714 343 1715 347
rect 1719 343 1720 347
rect 1714 342 1720 343
rect 1786 347 1792 348
rect 1786 343 1787 347
rect 1791 343 1792 347
rect 1786 342 1792 343
rect 1614 332 1620 333
rect 1614 328 1615 332
rect 1619 328 1620 332
rect 1614 327 1620 328
rect 1678 332 1684 333
rect 1678 328 1679 332
rect 1683 328 1684 332
rect 1678 327 1684 328
rect 1616 323 1618 327
rect 1680 323 1682 327
rect 1615 322 1619 323
rect 1615 317 1619 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1679 322 1683 323
rect 1679 317 1683 318
rect 1695 322 1699 323
rect 1695 317 1699 318
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1694 316 1700 317
rect 1694 312 1695 316
rect 1699 312 1700 316
rect 1694 311 1700 312
rect 1570 299 1576 300
rect 1570 295 1571 299
rect 1575 295 1576 299
rect 1570 294 1576 295
rect 1558 288 1564 289
rect 1558 284 1559 288
rect 1563 284 1564 288
rect 1558 283 1564 284
rect 1622 288 1628 289
rect 1622 284 1623 288
rect 1627 284 1628 288
rect 1622 283 1628 284
rect 1694 288 1700 289
rect 1694 284 1695 288
rect 1699 284 1700 288
rect 1694 283 1700 284
rect 1542 275 1548 276
rect 1542 271 1543 275
rect 1547 271 1548 275
rect 1542 270 1548 271
rect 1560 263 1562 283
rect 1624 263 1626 283
rect 1696 263 1698 283
rect 1716 268 1718 342
rect 1750 332 1756 333
rect 1750 328 1751 332
rect 1755 328 1756 332
rect 1750 327 1756 328
rect 1752 323 1754 327
rect 1751 322 1755 323
rect 1751 317 1755 318
rect 1775 322 1779 323
rect 1775 317 1779 318
rect 1774 316 1780 317
rect 1774 312 1775 316
rect 1779 312 1780 316
rect 1774 311 1780 312
rect 1730 299 1736 300
rect 1730 295 1731 299
rect 1735 295 1736 299
rect 1730 294 1736 295
rect 1732 276 1734 294
rect 1774 288 1780 289
rect 1774 284 1775 288
rect 1779 284 1780 288
rect 1774 283 1780 284
rect 1730 275 1736 276
rect 1730 271 1731 275
rect 1735 271 1736 275
rect 1730 270 1736 271
rect 1714 267 1720 268
rect 1714 263 1715 267
rect 1719 263 1720 267
rect 1776 263 1778 283
rect 1788 276 1790 342
rect 1830 332 1836 333
rect 1830 328 1831 332
rect 1835 328 1836 332
rect 1830 327 1836 328
rect 1918 332 1924 333
rect 1918 328 1919 332
rect 1923 328 1924 332
rect 1918 327 1924 328
rect 1832 323 1834 327
rect 1920 323 1922 327
rect 1831 322 1835 323
rect 1831 317 1835 318
rect 1855 322 1859 323
rect 1855 317 1859 318
rect 1919 322 1923 323
rect 1919 317 1923 318
rect 1935 322 1939 323
rect 1935 317 1939 318
rect 1854 316 1860 317
rect 1854 312 1855 316
rect 1859 312 1860 316
rect 1854 311 1860 312
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 1934 311 1940 312
rect 1944 300 1946 366
rect 2000 348 2002 382
rect 2024 379 2026 395
rect 2032 388 2034 450
rect 2118 443 2124 444
rect 2070 440 2076 441
rect 2070 436 2071 440
rect 2075 436 2076 440
rect 2118 439 2119 443
rect 2123 439 2124 443
rect 2118 438 2124 439
rect 2070 435 2076 436
rect 2120 435 2122 438
rect 2071 434 2075 435
rect 2071 429 2075 430
rect 2119 434 2123 435
rect 2119 429 2123 430
rect 2070 428 2076 429
rect 2070 424 2071 428
rect 2075 424 2076 428
rect 2120 426 2122 429
rect 2070 423 2076 424
rect 2118 425 2124 426
rect 2118 421 2119 425
rect 2123 421 2124 425
rect 2118 420 2124 421
rect 2062 411 2068 412
rect 2062 407 2063 411
rect 2067 407 2068 411
rect 2062 406 2068 407
rect 2082 411 2088 412
rect 2082 407 2083 411
rect 2087 407 2088 411
rect 2082 406 2088 407
rect 2118 408 2124 409
rect 2064 388 2066 406
rect 2070 400 2076 401
rect 2070 396 2071 400
rect 2075 396 2076 400
rect 2070 395 2076 396
rect 2030 387 2036 388
rect 2030 383 2031 387
rect 2035 383 2036 387
rect 2030 382 2036 383
rect 2062 387 2068 388
rect 2062 383 2063 387
rect 2067 383 2068 387
rect 2062 382 2068 383
rect 2072 379 2074 395
rect 2007 378 2011 379
rect 2007 373 2011 374
rect 2023 378 2027 379
rect 2023 373 2027 374
rect 2071 378 2075 379
rect 2071 373 2075 374
rect 2008 361 2010 373
rect 2072 361 2074 373
rect 2084 372 2086 406
rect 2118 404 2119 408
rect 2123 404 2124 408
rect 2118 403 2124 404
rect 2120 379 2122 403
rect 2119 378 2123 379
rect 2119 373 2123 374
rect 2082 371 2088 372
rect 2082 367 2083 371
rect 2087 367 2088 371
rect 2082 366 2088 367
rect 2006 360 2012 361
rect 2006 356 2007 360
rect 2011 356 2012 360
rect 2006 355 2012 356
rect 2070 360 2076 361
rect 2070 356 2071 360
rect 2075 356 2076 360
rect 2070 355 2076 356
rect 2120 353 2122 373
rect 2118 352 2124 353
rect 2118 348 2119 352
rect 2123 348 2124 352
rect 1998 347 2004 348
rect 1998 343 1999 347
rect 2003 343 2004 347
rect 1998 342 2004 343
rect 2078 347 2084 348
rect 2118 347 2124 348
rect 2078 343 2079 347
rect 2083 343 2084 347
rect 2078 342 2084 343
rect 2006 332 2012 333
rect 2006 328 2007 332
rect 2011 328 2012 332
rect 2006 327 2012 328
rect 2070 332 2076 333
rect 2070 328 2071 332
rect 2075 328 2076 332
rect 2070 327 2076 328
rect 2008 323 2010 327
rect 2072 323 2074 327
rect 2007 322 2011 323
rect 2007 317 2011 318
rect 2015 322 2019 323
rect 2015 317 2019 318
rect 2071 322 2075 323
rect 2071 317 2075 318
rect 2014 316 2020 317
rect 2014 312 2015 316
rect 2019 312 2020 316
rect 2014 311 2020 312
rect 2070 316 2076 317
rect 2070 312 2071 316
rect 2075 312 2076 316
rect 2070 311 2076 312
rect 1926 299 1932 300
rect 1926 295 1927 299
rect 1931 295 1932 299
rect 1926 294 1932 295
rect 1942 299 1948 300
rect 1942 295 1943 299
rect 1947 295 1948 299
rect 1942 294 1948 295
rect 2006 299 2012 300
rect 2006 295 2007 299
rect 2011 295 2012 299
rect 2006 294 2012 295
rect 1854 288 1860 289
rect 1854 284 1855 288
rect 1859 284 1860 288
rect 1854 283 1860 284
rect 1786 275 1792 276
rect 1786 271 1787 275
rect 1791 271 1792 275
rect 1786 270 1792 271
rect 1856 263 1858 283
rect 1928 276 1930 294
rect 1934 288 1940 289
rect 1934 284 1935 288
rect 1939 284 1940 288
rect 1934 283 1940 284
rect 1862 275 1868 276
rect 1862 271 1863 275
rect 1867 271 1868 275
rect 1862 270 1868 271
rect 1926 275 1932 276
rect 1926 271 1927 275
rect 1931 271 1932 275
rect 1926 270 1932 271
rect 1527 262 1531 263
rect 1527 257 1531 258
rect 1559 262 1563 263
rect 1559 257 1563 258
rect 1607 262 1611 263
rect 1607 257 1611 258
rect 1623 262 1627 263
rect 1623 257 1627 258
rect 1687 262 1691 263
rect 1687 257 1691 258
rect 1695 262 1699 263
rect 1714 262 1720 263
rect 1767 262 1771 263
rect 1695 257 1699 258
rect 1767 257 1771 258
rect 1775 262 1779 263
rect 1775 257 1779 258
rect 1839 262 1843 263
rect 1839 257 1843 258
rect 1855 262 1859 263
rect 1855 257 1859 258
rect 1510 255 1516 256
rect 1510 251 1511 255
rect 1515 251 1516 255
rect 1510 250 1516 251
rect 1518 255 1524 256
rect 1518 251 1519 255
rect 1523 251 1524 255
rect 1518 250 1524 251
rect 1454 244 1460 245
rect 1454 240 1455 244
rect 1459 240 1460 244
rect 1454 239 1460 240
rect 1512 232 1514 250
rect 1528 245 1530 257
rect 1608 245 1610 257
rect 1634 255 1640 256
rect 1634 251 1635 255
rect 1639 251 1640 255
rect 1634 250 1640 251
rect 1526 244 1532 245
rect 1526 240 1527 244
rect 1531 240 1532 244
rect 1526 239 1532 240
rect 1606 244 1612 245
rect 1606 240 1607 244
rect 1611 240 1612 244
rect 1606 239 1612 240
rect 1636 232 1638 250
rect 1688 245 1690 257
rect 1714 255 1720 256
rect 1714 251 1715 255
rect 1719 251 1720 255
rect 1714 250 1720 251
rect 1686 244 1692 245
rect 1686 240 1687 244
rect 1691 240 1692 244
rect 1686 239 1692 240
rect 1716 232 1718 250
rect 1768 245 1770 257
rect 1840 245 1842 257
rect 1766 244 1772 245
rect 1766 240 1767 244
rect 1771 240 1772 244
rect 1766 239 1772 240
rect 1838 244 1844 245
rect 1838 240 1839 244
rect 1843 240 1844 244
rect 1838 239 1844 240
rect 1864 232 1866 270
rect 1936 263 1938 283
rect 1919 262 1923 263
rect 1919 257 1923 258
rect 1935 262 1939 263
rect 1935 257 1939 258
rect 1999 262 2003 263
rect 1999 257 2003 258
rect 1906 255 1912 256
rect 1906 251 1907 255
rect 1911 251 1912 255
rect 1906 250 1912 251
rect 1908 232 1910 250
rect 1920 245 1922 257
rect 1974 255 1980 256
rect 1974 251 1975 255
rect 1979 251 1980 255
rect 1974 250 1980 251
rect 1918 244 1924 245
rect 1918 240 1919 244
rect 1923 240 1924 244
rect 1918 239 1924 240
rect 1478 231 1484 232
rect 1478 227 1479 231
rect 1483 227 1484 231
rect 1478 226 1484 227
rect 1510 231 1516 232
rect 1510 227 1511 231
rect 1515 227 1516 231
rect 1510 226 1516 227
rect 1634 231 1640 232
rect 1634 227 1635 231
rect 1639 227 1640 231
rect 1634 226 1640 227
rect 1714 231 1720 232
rect 1714 227 1715 231
rect 1719 227 1720 231
rect 1714 226 1720 227
rect 1742 231 1748 232
rect 1742 227 1743 231
rect 1747 227 1748 231
rect 1742 226 1748 227
rect 1862 231 1868 232
rect 1862 227 1863 231
rect 1867 227 1868 231
rect 1862 226 1868 227
rect 1906 231 1912 232
rect 1906 227 1907 231
rect 1911 227 1912 231
rect 1906 226 1912 227
rect 1454 216 1460 217
rect 1454 212 1455 216
rect 1459 212 1460 216
rect 1454 211 1460 212
rect 1455 210 1459 211
rect 1455 205 1459 206
rect 1471 210 1475 211
rect 1471 205 1475 206
rect 1470 204 1476 205
rect 1470 200 1471 204
rect 1475 200 1476 204
rect 1470 199 1476 200
rect 1390 187 1396 188
rect 1390 183 1391 187
rect 1395 183 1396 187
rect 1390 182 1396 183
rect 1422 187 1428 188
rect 1422 183 1423 187
rect 1427 183 1428 187
rect 1422 182 1428 183
rect 1326 176 1332 177
rect 1326 172 1327 176
rect 1331 172 1332 176
rect 1326 171 1332 172
rect 1278 163 1284 164
rect 1278 159 1279 163
rect 1283 159 1284 163
rect 1278 158 1284 159
rect 1298 163 1304 164
rect 1298 159 1299 163
rect 1303 159 1304 163
rect 1298 158 1304 159
rect 1199 138 1203 139
rect 1199 133 1203 134
rect 1207 138 1211 139
rect 1207 133 1211 134
rect 1263 138 1267 139
rect 1263 133 1267 134
rect 1271 138 1275 139
rect 1271 133 1275 134
rect 1170 131 1176 132
rect 1170 127 1171 131
rect 1175 127 1176 131
rect 1170 126 1176 127
rect 1208 121 1210 133
rect 1234 131 1240 132
rect 1234 127 1235 131
rect 1239 127 1240 131
rect 1234 126 1240 127
rect 1158 120 1164 121
rect 1158 116 1159 120
rect 1163 116 1164 120
rect 1158 115 1164 116
rect 1206 120 1212 121
rect 1206 116 1207 120
rect 1211 116 1212 120
rect 1206 115 1212 116
rect 1236 108 1238 126
rect 1272 121 1274 133
rect 1270 120 1276 121
rect 1270 116 1271 120
rect 1275 116 1276 120
rect 1270 115 1276 116
rect 1300 108 1302 158
rect 1328 139 1330 171
rect 1392 164 1394 182
rect 1398 176 1404 177
rect 1398 172 1399 176
rect 1403 172 1404 176
rect 1398 171 1404 172
rect 1470 176 1476 177
rect 1470 172 1471 176
rect 1475 172 1476 176
rect 1470 171 1476 172
rect 1390 163 1396 164
rect 1390 159 1391 163
rect 1395 159 1396 163
rect 1390 158 1396 159
rect 1358 139 1364 140
rect 1400 139 1402 171
rect 1472 139 1474 171
rect 1480 164 1482 226
rect 1526 216 1532 217
rect 1526 212 1527 216
rect 1531 212 1532 216
rect 1526 211 1532 212
rect 1606 216 1612 217
rect 1606 212 1607 216
rect 1611 212 1612 216
rect 1606 211 1612 212
rect 1686 216 1692 217
rect 1686 212 1687 216
rect 1691 212 1692 216
rect 1686 211 1692 212
rect 1527 210 1531 211
rect 1527 205 1531 206
rect 1543 210 1547 211
rect 1543 205 1547 206
rect 1607 210 1611 211
rect 1607 205 1611 206
rect 1671 210 1675 211
rect 1671 205 1675 206
rect 1687 210 1691 211
rect 1687 205 1691 206
rect 1735 210 1739 211
rect 1735 205 1739 206
rect 1542 204 1548 205
rect 1542 200 1543 204
rect 1547 200 1548 204
rect 1542 199 1548 200
rect 1606 204 1612 205
rect 1606 200 1607 204
rect 1611 200 1612 204
rect 1606 199 1612 200
rect 1670 204 1676 205
rect 1670 200 1671 204
rect 1675 200 1676 204
rect 1670 199 1676 200
rect 1734 204 1740 205
rect 1734 200 1735 204
rect 1739 200 1740 204
rect 1734 199 1740 200
rect 1534 187 1540 188
rect 1534 183 1535 187
rect 1539 183 1540 187
rect 1534 182 1540 183
rect 1550 187 1556 188
rect 1550 183 1551 187
rect 1555 183 1556 187
rect 1550 182 1556 183
rect 1578 187 1584 188
rect 1578 183 1579 187
rect 1583 183 1584 187
rect 1578 182 1584 183
rect 1536 164 1538 182
rect 1542 176 1548 177
rect 1542 172 1543 176
rect 1547 172 1548 176
rect 1542 171 1548 172
rect 1478 163 1484 164
rect 1478 159 1479 163
rect 1483 159 1484 163
rect 1478 158 1484 159
rect 1534 163 1540 164
rect 1534 159 1535 163
rect 1539 159 1540 163
rect 1534 158 1540 159
rect 1544 139 1546 171
rect 1552 140 1554 182
rect 1550 139 1556 140
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1335 138 1339 139
rect 1358 135 1359 139
rect 1363 135 1364 139
rect 1358 134 1364 135
rect 1399 138 1403 139
rect 1335 133 1339 134
rect 1336 121 1338 133
rect 1334 120 1340 121
rect 1334 116 1335 120
rect 1339 116 1340 120
rect 1334 115 1340 116
rect 1360 108 1362 134
rect 1399 133 1403 134
rect 1455 138 1459 139
rect 1455 133 1459 134
rect 1471 138 1475 139
rect 1471 133 1475 134
rect 1511 138 1515 139
rect 1511 133 1515 134
rect 1543 138 1547 139
rect 1550 135 1551 139
rect 1555 135 1556 139
rect 1550 134 1556 135
rect 1559 138 1563 139
rect 1543 133 1547 134
rect 1559 133 1563 134
rect 1386 131 1392 132
rect 1386 127 1387 131
rect 1391 127 1392 131
rect 1386 126 1392 127
rect 1388 108 1390 126
rect 1400 121 1402 133
rect 1438 131 1444 132
rect 1438 127 1439 131
rect 1443 127 1444 131
rect 1438 126 1444 127
rect 1398 120 1404 121
rect 1398 116 1399 120
rect 1403 116 1404 120
rect 1398 115 1404 116
rect 1440 108 1442 126
rect 1456 121 1458 133
rect 1498 131 1504 132
rect 1498 127 1499 131
rect 1503 127 1504 131
rect 1498 126 1504 127
rect 1454 120 1460 121
rect 1454 116 1455 120
rect 1459 116 1460 120
rect 1454 115 1460 116
rect 1500 108 1502 126
rect 1512 121 1514 133
rect 1560 121 1562 133
rect 1580 132 1582 182
rect 1606 176 1612 177
rect 1606 172 1607 176
rect 1611 172 1612 176
rect 1606 171 1612 172
rect 1670 176 1676 177
rect 1670 172 1671 176
rect 1675 172 1676 176
rect 1670 171 1676 172
rect 1734 176 1740 177
rect 1734 172 1735 176
rect 1739 172 1740 176
rect 1734 171 1740 172
rect 1608 139 1610 171
rect 1672 139 1674 171
rect 1736 139 1738 171
rect 1744 164 1746 226
rect 1766 216 1772 217
rect 1766 212 1767 216
rect 1771 212 1772 216
rect 1766 211 1772 212
rect 1838 216 1844 217
rect 1838 212 1839 216
rect 1843 212 1844 216
rect 1838 211 1844 212
rect 1918 216 1924 217
rect 1918 212 1919 216
rect 1923 212 1924 216
rect 1918 211 1924 212
rect 1767 210 1771 211
rect 1767 205 1771 206
rect 1807 210 1811 211
rect 1807 205 1811 206
rect 1839 210 1843 211
rect 1839 205 1843 206
rect 1879 210 1883 211
rect 1879 205 1883 206
rect 1919 210 1923 211
rect 1919 205 1923 206
rect 1951 210 1955 211
rect 1951 205 1955 206
rect 1806 204 1812 205
rect 1806 200 1807 204
rect 1811 200 1812 204
rect 1806 199 1812 200
rect 1878 204 1884 205
rect 1878 200 1879 204
rect 1883 200 1884 204
rect 1878 199 1884 200
rect 1950 204 1956 205
rect 1950 200 1951 204
rect 1955 200 1956 204
rect 1950 199 1956 200
rect 1976 196 1978 250
rect 2000 245 2002 257
rect 2008 256 2010 294
rect 2014 288 2020 289
rect 2014 284 2015 288
rect 2019 284 2020 288
rect 2014 283 2020 284
rect 2070 288 2076 289
rect 2070 284 2071 288
rect 2075 284 2076 288
rect 2070 283 2076 284
rect 2016 263 2018 283
rect 2072 263 2074 283
rect 2080 276 2082 342
rect 2118 335 2124 336
rect 2118 331 2119 335
rect 2123 331 2124 335
rect 2118 330 2124 331
rect 2120 323 2122 330
rect 2119 322 2123 323
rect 2119 317 2123 318
rect 2120 314 2122 317
rect 2118 313 2124 314
rect 2118 309 2119 313
rect 2123 309 2124 313
rect 2118 308 2124 309
rect 2118 296 2124 297
rect 2118 292 2119 296
rect 2123 292 2124 296
rect 2118 291 2124 292
rect 2078 275 2084 276
rect 2078 271 2079 275
rect 2083 271 2084 275
rect 2078 270 2084 271
rect 2120 263 2122 291
rect 2015 262 2019 263
rect 2015 257 2019 258
rect 2071 262 2075 263
rect 2071 257 2075 258
rect 2119 262 2123 263
rect 2119 257 2123 258
rect 2006 255 2012 256
rect 2006 251 2007 255
rect 2011 251 2012 255
rect 2006 250 2012 251
rect 2026 255 2032 256
rect 2026 251 2027 255
rect 2031 251 2032 255
rect 2026 250 2032 251
rect 1998 244 2004 245
rect 1998 240 1999 244
rect 2003 240 2004 244
rect 1998 239 2004 240
rect 2028 232 2030 250
rect 2072 245 2074 257
rect 2070 244 2076 245
rect 2070 240 2071 244
rect 2075 240 2076 244
rect 2070 239 2076 240
rect 2120 237 2122 257
rect 2118 236 2124 237
rect 2118 232 2119 236
rect 2123 232 2124 236
rect 2026 231 2032 232
rect 2026 227 2027 231
rect 2031 227 2032 231
rect 2026 226 2032 227
rect 2086 231 2092 232
rect 2118 231 2124 232
rect 2086 227 2087 231
rect 2091 227 2092 231
rect 2086 226 2092 227
rect 1998 216 2004 217
rect 1998 212 1999 216
rect 2003 212 2004 216
rect 1998 211 2004 212
rect 2070 216 2076 217
rect 2070 212 2071 216
rect 2075 212 2076 216
rect 2070 211 2076 212
rect 1999 210 2003 211
rect 1999 205 2003 206
rect 2023 210 2027 211
rect 2023 205 2027 206
rect 2071 210 2075 211
rect 2071 205 2075 206
rect 2022 204 2028 205
rect 2022 200 2023 204
rect 2027 200 2028 204
rect 2022 199 2028 200
rect 2070 204 2076 205
rect 2070 200 2071 204
rect 2075 200 2076 204
rect 2070 199 2076 200
rect 1974 195 1980 196
rect 1974 191 1975 195
rect 1979 191 1980 195
rect 1974 190 1980 191
rect 1870 187 1876 188
rect 1870 183 1871 187
rect 1875 183 1876 187
rect 1870 182 1876 183
rect 1942 187 1948 188
rect 1942 183 1943 187
rect 1947 183 1948 187
rect 1942 182 1948 183
rect 2014 187 2020 188
rect 2014 183 2015 187
rect 2019 183 2020 187
rect 2014 182 2020 183
rect 2078 187 2084 188
rect 2078 183 2079 187
rect 2083 183 2084 187
rect 2078 182 2084 183
rect 1806 176 1812 177
rect 1806 172 1807 176
rect 1811 172 1812 176
rect 1806 171 1812 172
rect 1742 163 1748 164
rect 1742 159 1743 163
rect 1747 159 1748 163
rect 1742 158 1748 159
rect 1808 139 1810 171
rect 1872 164 1874 182
rect 1878 176 1884 177
rect 1878 172 1879 176
rect 1883 172 1884 176
rect 1878 171 1884 172
rect 1870 163 1876 164
rect 1870 159 1871 163
rect 1875 159 1876 163
rect 1870 158 1876 159
rect 1880 139 1882 171
rect 1944 164 1946 182
rect 1950 176 1956 177
rect 1950 172 1951 176
rect 1955 172 1956 176
rect 1950 171 1956 172
rect 1942 163 1948 164
rect 1942 159 1943 163
rect 1947 159 1948 163
rect 1942 158 1948 159
rect 1952 139 1954 171
rect 2016 164 2018 182
rect 2022 176 2028 177
rect 2022 172 2023 176
rect 2027 172 2028 176
rect 2022 171 2028 172
rect 2070 176 2076 177
rect 2070 172 2071 176
rect 2075 172 2076 176
rect 2070 171 2076 172
rect 2014 163 2020 164
rect 2014 159 2015 163
rect 2019 159 2020 163
rect 2014 158 2020 159
rect 1974 155 1980 156
rect 1974 151 1975 155
rect 1979 151 1980 155
rect 1974 150 1980 151
rect 1607 138 1611 139
rect 1607 133 1611 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1671 138 1675 139
rect 1671 133 1675 134
rect 1687 138 1691 139
rect 1687 133 1691 134
rect 1727 138 1731 139
rect 1727 133 1731 134
rect 1735 138 1739 139
rect 1735 133 1739 134
rect 1767 138 1771 139
rect 1767 133 1771 134
rect 1807 138 1811 139
rect 1807 133 1811 134
rect 1855 138 1859 139
rect 1855 133 1859 134
rect 1879 138 1883 139
rect 1879 133 1883 134
rect 1903 138 1907 139
rect 1903 133 1907 134
rect 1951 138 1955 139
rect 1951 133 1955 134
rect 1578 131 1584 132
rect 1578 127 1579 131
rect 1583 127 1584 131
rect 1578 126 1584 127
rect 1586 131 1592 132
rect 1586 127 1587 131
rect 1591 127 1592 131
rect 1586 126 1592 127
rect 1510 120 1516 121
rect 1510 116 1511 120
rect 1515 116 1516 120
rect 1510 115 1516 116
rect 1558 120 1564 121
rect 1558 116 1559 120
rect 1563 116 1564 120
rect 1558 115 1564 116
rect 1588 108 1590 126
rect 1608 121 1610 133
rect 1634 131 1640 132
rect 1634 127 1635 131
rect 1639 127 1640 131
rect 1634 126 1640 127
rect 1606 120 1612 121
rect 1606 116 1607 120
rect 1611 116 1612 120
rect 1606 115 1612 116
rect 1636 108 1638 126
rect 1648 121 1650 133
rect 1678 131 1684 132
rect 1678 127 1679 131
rect 1683 127 1684 131
rect 1678 126 1684 127
rect 1646 120 1652 121
rect 1646 116 1647 120
rect 1651 116 1652 120
rect 1646 115 1652 116
rect 1680 108 1682 126
rect 1688 121 1690 133
rect 1714 131 1720 132
rect 1714 127 1715 131
rect 1719 127 1720 131
rect 1714 126 1720 127
rect 1686 120 1692 121
rect 1686 116 1687 120
rect 1691 116 1692 120
rect 1686 115 1692 116
rect 1716 108 1718 126
rect 1728 121 1730 133
rect 1754 131 1760 132
rect 1754 127 1755 131
rect 1759 127 1760 131
rect 1754 126 1760 127
rect 1726 120 1732 121
rect 1726 116 1727 120
rect 1731 116 1732 120
rect 1726 115 1732 116
rect 1756 108 1758 126
rect 1768 121 1770 133
rect 1794 131 1800 132
rect 1794 127 1795 131
rect 1799 127 1800 131
rect 1794 126 1800 127
rect 1766 120 1772 121
rect 1766 116 1767 120
rect 1771 116 1772 120
rect 1766 115 1772 116
rect 1796 108 1798 126
rect 1808 121 1810 133
rect 1834 131 1840 132
rect 1834 127 1835 131
rect 1839 127 1840 131
rect 1834 126 1840 127
rect 1806 120 1812 121
rect 1806 116 1807 120
rect 1811 116 1812 120
rect 1806 115 1812 116
rect 1836 108 1838 126
rect 1856 121 1858 133
rect 1904 121 1906 133
rect 1930 131 1936 132
rect 1930 127 1931 131
rect 1935 127 1936 131
rect 1930 126 1936 127
rect 1854 120 1860 121
rect 1854 116 1855 120
rect 1859 116 1860 120
rect 1854 115 1860 116
rect 1902 120 1908 121
rect 1902 116 1903 120
rect 1907 116 1908 120
rect 1902 115 1908 116
rect 1932 108 1934 126
rect 1952 121 1954 133
rect 1950 120 1956 121
rect 1950 116 1951 120
rect 1955 116 1956 120
rect 1950 115 1956 116
rect 1976 108 1978 150
rect 2024 139 2026 171
rect 2072 139 2074 171
rect 1991 138 1995 139
rect 1991 133 1995 134
rect 2023 138 2027 139
rect 2023 133 2027 134
rect 2031 138 2035 139
rect 2031 133 2035 134
rect 2071 138 2075 139
rect 2071 133 2075 134
rect 1992 121 1994 133
rect 2014 131 2020 132
rect 2014 127 2015 131
rect 2019 127 2020 131
rect 2014 126 2020 127
rect 1990 120 1996 121
rect 1990 116 1991 120
rect 1995 116 1996 120
rect 1990 115 1996 116
rect 2016 108 2018 126
rect 2032 121 2034 133
rect 2072 121 2074 133
rect 2080 132 2082 182
rect 2088 164 2090 226
rect 2118 219 2124 220
rect 2118 215 2119 219
rect 2123 215 2124 219
rect 2118 214 2124 215
rect 2120 211 2122 214
rect 2119 210 2123 211
rect 2119 205 2123 206
rect 2120 202 2122 205
rect 2118 201 2124 202
rect 2118 197 2119 201
rect 2123 197 2124 201
rect 2118 196 2124 197
rect 2118 184 2124 185
rect 2118 180 2119 184
rect 2123 180 2124 184
rect 2118 179 2124 180
rect 2086 163 2092 164
rect 2086 159 2087 163
rect 2091 159 2092 163
rect 2086 158 2092 159
rect 2120 139 2122 179
rect 2119 138 2123 139
rect 2119 133 2123 134
rect 2078 131 2084 132
rect 2078 127 2079 131
rect 2083 127 2084 131
rect 2078 126 2084 127
rect 2030 120 2036 121
rect 2030 116 2031 120
rect 2035 116 2036 120
rect 2030 115 2036 116
rect 2070 120 2076 121
rect 2070 116 2071 120
rect 2075 116 2076 120
rect 2070 115 2076 116
rect 2120 113 2122 133
rect 2118 112 2124 113
rect 2118 108 2119 112
rect 2123 108 2124 112
rect 1134 107 1140 108
rect 1142 107 1148 108
rect 866 103 867 107
rect 871 103 872 107
rect 866 102 872 103
rect 1142 103 1143 107
rect 1147 103 1148 107
rect 1142 102 1148 103
rect 1234 107 1240 108
rect 1234 103 1235 107
rect 1239 103 1240 107
rect 1234 102 1240 103
rect 1298 107 1304 108
rect 1298 103 1299 107
rect 1303 103 1304 107
rect 1298 102 1304 103
rect 1358 107 1364 108
rect 1358 103 1359 107
rect 1363 103 1364 107
rect 1358 102 1364 103
rect 1386 107 1392 108
rect 1386 103 1387 107
rect 1391 103 1392 107
rect 1386 102 1392 103
rect 1438 107 1444 108
rect 1438 103 1439 107
rect 1443 103 1444 107
rect 1438 102 1444 103
rect 1498 107 1504 108
rect 1498 103 1499 107
rect 1503 103 1504 107
rect 1498 102 1504 103
rect 1586 107 1592 108
rect 1586 103 1587 107
rect 1591 103 1592 107
rect 1586 102 1592 103
rect 1634 107 1640 108
rect 1634 103 1635 107
rect 1639 103 1640 107
rect 1634 102 1640 103
rect 1674 107 1682 108
rect 1674 103 1675 107
rect 1679 104 1682 107
rect 1714 107 1720 108
rect 1679 103 1680 104
rect 1674 102 1680 103
rect 1714 103 1715 107
rect 1719 103 1720 107
rect 1714 102 1720 103
rect 1754 107 1760 108
rect 1754 103 1755 107
rect 1759 103 1760 107
rect 1754 102 1760 103
rect 1794 107 1800 108
rect 1794 103 1795 107
rect 1799 103 1800 107
rect 1794 102 1800 103
rect 1834 107 1840 108
rect 1834 103 1835 107
rect 1839 103 1840 107
rect 1834 102 1840 103
rect 1930 107 1936 108
rect 1930 103 1931 107
rect 1935 103 1936 107
rect 1930 102 1936 103
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 1974 102 1980 103
rect 2014 107 2020 108
rect 2118 107 2124 108
rect 2014 103 2015 107
rect 2019 103 2020 107
rect 2014 102 2020 103
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1094 95 1100 96
rect 110 90 116 91
rect 142 92 148 93
rect 112 87 114 90
rect 142 88 143 92
rect 147 88 148 92
rect 142 87 148 88
rect 182 92 188 93
rect 182 88 183 92
rect 187 88 188 92
rect 182 87 188 88
rect 222 92 228 93
rect 222 88 223 92
rect 227 88 228 92
rect 222 87 228 88
rect 262 92 268 93
rect 262 88 263 92
rect 267 88 268 92
rect 262 87 268 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 342 92 348 93
rect 342 88 343 92
rect 347 88 348 92
rect 342 87 348 88
rect 382 92 388 93
rect 382 88 383 92
rect 387 88 388 92
rect 382 87 388 88
rect 422 92 428 93
rect 422 88 423 92
rect 427 88 428 92
rect 422 87 428 88
rect 462 92 468 93
rect 462 88 463 92
rect 467 88 468 92
rect 462 87 468 88
rect 502 92 508 93
rect 502 88 503 92
rect 507 88 508 92
rect 502 87 508 88
rect 542 92 548 93
rect 542 88 543 92
rect 547 88 548 92
rect 542 87 548 88
rect 582 92 588 93
rect 582 88 583 92
rect 587 88 588 92
rect 582 87 588 88
rect 622 92 628 93
rect 622 88 623 92
rect 627 88 628 92
rect 622 87 628 88
rect 662 92 668 93
rect 662 88 663 92
rect 667 88 668 92
rect 662 87 668 88
rect 702 92 708 93
rect 702 88 703 92
rect 707 88 708 92
rect 702 87 708 88
rect 742 92 748 93
rect 742 88 743 92
rect 747 88 748 92
rect 742 87 748 88
rect 782 92 788 93
rect 782 88 783 92
rect 787 88 788 92
rect 782 87 788 88
rect 830 92 836 93
rect 830 88 831 92
rect 835 88 836 92
rect 830 87 836 88
rect 878 92 884 93
rect 878 88 879 92
rect 883 88 884 92
rect 878 87 884 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 966 92 972 93
rect 966 88 967 92
rect 971 88 972 92
rect 966 87 972 88
rect 1006 92 1012 93
rect 1006 88 1007 92
rect 1011 88 1012 92
rect 1006 87 1012 88
rect 1046 92 1052 93
rect 1046 88 1047 92
rect 1051 88 1052 92
rect 1094 91 1095 95
rect 1099 91 1100 95
rect 1094 90 1100 91
rect 1134 95 1140 96
rect 1134 91 1135 95
rect 1139 91 1140 95
rect 2118 95 2124 96
rect 1134 90 1140 91
rect 1158 92 1164 93
rect 1046 87 1052 88
rect 1096 87 1098 90
rect 1136 87 1138 90
rect 1158 88 1159 92
rect 1163 88 1164 92
rect 1158 87 1164 88
rect 1206 92 1212 93
rect 1206 88 1207 92
rect 1211 88 1212 92
rect 1206 87 1212 88
rect 1270 92 1276 93
rect 1270 88 1271 92
rect 1275 88 1276 92
rect 1270 87 1276 88
rect 1334 92 1340 93
rect 1334 88 1335 92
rect 1339 88 1340 92
rect 1334 87 1340 88
rect 1398 92 1404 93
rect 1398 88 1399 92
rect 1403 88 1404 92
rect 1398 87 1404 88
rect 1454 92 1460 93
rect 1454 88 1455 92
rect 1459 88 1460 92
rect 1454 87 1460 88
rect 1510 92 1516 93
rect 1510 88 1511 92
rect 1515 88 1516 92
rect 1510 87 1516 88
rect 1558 92 1564 93
rect 1558 88 1559 92
rect 1563 88 1564 92
rect 1558 87 1564 88
rect 1606 92 1612 93
rect 1606 88 1607 92
rect 1611 88 1612 92
rect 1606 87 1612 88
rect 1646 92 1652 93
rect 1646 88 1647 92
rect 1651 88 1652 92
rect 1646 87 1652 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1726 92 1732 93
rect 1726 88 1727 92
rect 1731 88 1732 92
rect 1726 87 1732 88
rect 1766 92 1772 93
rect 1766 88 1767 92
rect 1771 88 1772 92
rect 1766 87 1772 88
rect 1806 92 1812 93
rect 1806 88 1807 92
rect 1811 88 1812 92
rect 1806 87 1812 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1902 92 1908 93
rect 1902 88 1903 92
rect 1907 88 1908 92
rect 1902 87 1908 88
rect 1950 92 1956 93
rect 1950 88 1951 92
rect 1955 88 1956 92
rect 1950 87 1956 88
rect 1990 92 1996 93
rect 1990 88 1991 92
rect 1995 88 1996 92
rect 1990 87 1996 88
rect 2030 92 2036 93
rect 2030 88 2031 92
rect 2035 88 2036 92
rect 2030 87 2036 88
rect 2070 92 2076 93
rect 2070 88 2071 92
rect 2075 88 2076 92
rect 2118 91 2119 95
rect 2123 91 2124 95
rect 2118 90 2124 91
rect 2070 87 2076 88
rect 2120 87 2122 90
rect 111 86 115 87
rect 111 81 115 82
rect 143 86 147 87
rect 143 81 147 82
rect 183 86 187 87
rect 183 81 187 82
rect 223 86 227 87
rect 223 81 227 82
rect 263 86 267 87
rect 263 81 267 82
rect 303 86 307 87
rect 303 81 307 82
rect 343 86 347 87
rect 343 81 347 82
rect 383 86 387 87
rect 383 81 387 82
rect 423 86 427 87
rect 423 81 427 82
rect 463 86 467 87
rect 463 81 467 82
rect 503 86 507 87
rect 503 81 507 82
rect 543 86 547 87
rect 543 81 547 82
rect 583 86 587 87
rect 583 81 587 82
rect 623 86 627 87
rect 623 81 627 82
rect 663 86 667 87
rect 663 81 667 82
rect 703 86 707 87
rect 703 81 707 82
rect 743 86 747 87
rect 743 81 747 82
rect 783 86 787 87
rect 783 81 787 82
rect 831 86 835 87
rect 831 81 835 82
rect 879 86 883 87
rect 879 81 883 82
rect 927 86 931 87
rect 927 81 931 82
rect 967 86 971 87
rect 967 81 971 82
rect 1007 86 1011 87
rect 1007 81 1011 82
rect 1047 86 1051 87
rect 1047 81 1051 82
rect 1095 86 1099 87
rect 1095 81 1099 82
rect 1135 86 1139 87
rect 1135 81 1139 82
rect 1159 86 1163 87
rect 1159 81 1163 82
rect 1207 86 1211 87
rect 1207 81 1211 82
rect 1271 86 1275 87
rect 1271 81 1275 82
rect 1335 86 1339 87
rect 1335 81 1339 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1455 86 1459 87
rect 1455 81 1459 82
rect 1511 86 1515 87
rect 1511 81 1515 82
rect 1559 86 1563 87
rect 1559 81 1563 82
rect 1607 86 1611 87
rect 1607 81 1611 82
rect 1647 86 1651 87
rect 1647 81 1651 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1727 86 1731 87
rect 1727 81 1731 82
rect 1767 86 1771 87
rect 1767 81 1771 82
rect 1807 86 1811 87
rect 1807 81 1811 82
rect 1855 86 1859 87
rect 1855 81 1859 82
rect 1903 86 1907 87
rect 1903 81 1907 82
rect 1951 86 1955 87
rect 1951 81 1955 82
rect 1991 86 1995 87
rect 1991 81 1995 82
rect 2031 86 2035 87
rect 2031 81 2035 82
rect 2071 86 2075 87
rect 2071 81 2075 82
rect 2119 86 2123 87
rect 2119 81 2123 82
<< m4c >>
rect 1135 2226 1139 2230
rect 1687 2226 1691 2230
rect 1727 2226 1731 2230
rect 1767 2226 1771 2230
rect 1807 2226 1811 2230
rect 2119 2226 2123 2230
rect 111 2210 115 2214
rect 135 2210 139 2214
rect 175 2210 179 2214
rect 215 2210 219 2214
rect 255 2210 259 2214
rect 319 2210 323 2214
rect 383 2210 387 2214
rect 447 2210 451 2214
rect 511 2210 515 2214
rect 575 2210 579 2214
rect 631 2210 635 2214
rect 687 2210 691 2214
rect 735 2210 739 2214
rect 791 2210 795 2214
rect 847 2210 851 2214
rect 903 2210 907 2214
rect 1095 2210 1099 2214
rect 1135 2174 1139 2178
rect 1159 2174 1163 2178
rect 1199 2174 1203 2178
rect 1239 2174 1243 2178
rect 1279 2174 1283 2178
rect 1335 2174 1339 2178
rect 1391 2174 1395 2178
rect 1455 2174 1459 2178
rect 1527 2174 1531 2178
rect 1591 2174 1595 2178
rect 1663 2174 1667 2178
rect 111 2150 115 2154
rect 135 2150 139 2154
rect 175 2150 179 2154
rect 215 2150 219 2154
rect 231 2150 235 2154
rect 255 2150 259 2154
rect 271 2150 275 2154
rect 311 2150 315 2154
rect 319 2150 323 2154
rect 359 2150 363 2154
rect 383 2150 387 2154
rect 423 2150 427 2154
rect 447 2150 451 2154
rect 487 2150 491 2154
rect 511 2150 515 2154
rect 559 2150 563 2154
rect 575 2150 579 2154
rect 631 2150 635 2154
rect 639 2150 643 2154
rect 687 2150 691 2154
rect 719 2150 723 2154
rect 735 2150 739 2154
rect 791 2150 795 2154
rect 799 2150 803 2154
rect 847 2150 851 2154
rect 879 2150 883 2154
rect 903 2150 907 2154
rect 967 2150 971 2154
rect 1095 2150 1099 2154
rect 111 2094 115 2098
rect 231 2094 235 2098
rect 271 2094 275 2098
rect 303 2094 307 2098
rect 311 2094 315 2098
rect 351 2094 355 2098
rect 359 2094 363 2098
rect 407 2094 411 2098
rect 423 2094 427 2098
rect 471 2094 475 2098
rect 111 2038 115 2042
rect 183 2038 187 2042
rect 279 2038 283 2042
rect 303 2038 307 2042
rect 351 2038 355 2042
rect 375 2038 379 2042
rect 487 2094 491 2098
rect 543 2094 547 2098
rect 559 2094 563 2098
rect 623 2094 627 2098
rect 639 2094 643 2098
rect 703 2094 707 2098
rect 719 2094 723 2098
rect 1135 2122 1139 2126
rect 1159 2122 1163 2126
rect 1199 2122 1203 2126
rect 1239 2122 1243 2126
rect 1279 2122 1283 2126
rect 1295 2122 1299 2126
rect 783 2094 787 2098
rect 799 2094 803 2098
rect 863 2094 867 2098
rect 879 2094 883 2098
rect 951 2094 955 2098
rect 967 2094 971 2098
rect 407 2038 411 2042
rect 463 2038 467 2042
rect 471 2038 475 2042
rect 543 2038 547 2042
rect 623 2038 627 2042
rect 695 2038 699 2042
rect 703 2038 707 2042
rect 759 2038 763 2042
rect 111 1986 115 1990
rect 159 1986 163 1990
rect 183 1986 187 1990
rect 231 1986 235 1990
rect 279 1986 283 1990
rect 303 1986 307 1990
rect 375 1986 379 1990
rect 447 1986 451 1990
rect 111 1930 115 1934
rect 135 1930 139 1934
rect 159 1930 163 1934
rect 175 1930 179 1934
rect 463 1986 467 1990
rect 527 1986 531 1990
rect 543 1986 547 1990
rect 607 1986 611 1990
rect 623 1986 627 1990
rect 783 2038 787 2042
rect 815 2038 819 2042
rect 1039 2094 1043 2098
rect 1095 2094 1099 2098
rect 1135 2070 1139 2074
rect 1159 2070 1163 2074
rect 1687 2174 1691 2178
rect 1727 2174 1731 2178
rect 1735 2174 1739 2178
rect 1767 2174 1771 2178
rect 1807 2174 1811 2178
rect 1335 2122 1339 2126
rect 1367 2122 1371 2126
rect 1391 2122 1395 2126
rect 1439 2122 1443 2126
rect 1455 2122 1459 2126
rect 1519 2122 1523 2126
rect 1527 2122 1531 2126
rect 1591 2122 1595 2126
rect 1599 2122 1603 2126
rect 1199 2070 1203 2074
rect 1215 2070 1219 2074
rect 1239 2070 1243 2074
rect 1295 2070 1299 2074
rect 1303 2070 1307 2074
rect 1367 2070 1371 2074
rect 1399 2070 1403 2074
rect 1439 2070 1443 2074
rect 863 2038 867 2042
rect 911 2038 915 2042
rect 951 2038 955 2042
rect 959 2038 963 2042
rect 1007 2038 1011 2042
rect 1039 2038 1043 2042
rect 1047 2038 1051 2042
rect 1095 2038 1099 2042
rect 1135 2018 1139 2022
rect 1159 2018 1163 2022
rect 1215 2018 1219 2022
rect 1239 2018 1243 2022
rect 1303 2018 1307 2022
rect 1351 2018 1355 2022
rect 1495 2070 1499 2074
rect 1519 2070 1523 2074
rect 1591 2070 1595 2074
rect 1599 2070 1603 2074
rect 1663 2122 1667 2126
rect 1679 2122 1683 2126
rect 1735 2122 1739 2126
rect 1751 2122 1755 2126
rect 1879 2174 1883 2178
rect 2119 2174 2123 2178
rect 1807 2122 1811 2126
rect 1823 2122 1827 2126
rect 1879 2122 1883 2126
rect 1887 2122 1891 2126
rect 1951 2122 1955 2126
rect 2023 2122 2027 2126
rect 2071 2122 2075 2126
rect 2119 2122 2123 2126
rect 1679 2070 1683 2074
rect 1751 2070 1755 2074
rect 1759 2070 1763 2074
rect 1823 2070 1827 2074
rect 1831 2070 1835 2074
rect 1887 2070 1891 2074
rect 1895 2070 1899 2074
rect 1399 2018 1403 2022
rect 1455 2018 1459 2022
rect 1495 2018 1499 2022
rect 1559 2018 1563 2022
rect 1591 2018 1595 2022
rect 1655 2018 1659 2022
rect 687 1986 691 1990
rect 695 1986 699 1990
rect 759 1986 763 1990
rect 815 1986 819 1990
rect 831 1986 835 1990
rect 863 1986 867 1990
rect 911 1986 915 1990
rect 959 1986 963 1990
rect 991 1986 995 1990
rect 1007 1986 1011 1990
rect 1047 1986 1051 1990
rect 1095 1986 1099 1990
rect 231 1930 235 1934
rect 295 1930 299 1934
rect 303 1930 307 1934
rect 367 1930 371 1934
rect 375 1930 379 1934
rect 447 1930 451 1934
rect 527 1930 531 1934
rect 607 1930 611 1934
rect 615 1930 619 1934
rect 687 1930 691 1934
rect 703 1930 707 1934
rect 759 1930 763 1934
rect 791 1930 795 1934
rect 831 1930 835 1934
rect 879 1930 883 1934
rect 111 1874 115 1878
rect 135 1874 139 1878
rect 111 1818 115 1822
rect 135 1818 139 1822
rect 175 1874 179 1878
rect 223 1874 227 1878
rect 231 1874 235 1878
rect 287 1874 291 1878
rect 295 1874 299 1878
rect 359 1874 363 1878
rect 367 1874 371 1878
rect 431 1874 435 1878
rect 447 1874 451 1878
rect 503 1874 507 1878
rect 527 1874 531 1878
rect 567 1874 571 1878
rect 615 1874 619 1878
rect 631 1874 635 1878
rect 175 1818 179 1822
rect 183 1818 187 1822
rect 223 1818 227 1822
rect 263 1818 267 1822
rect 287 1818 291 1822
rect 351 1818 355 1822
rect 359 1818 363 1822
rect 431 1818 435 1822
rect 439 1818 443 1822
rect 503 1818 507 1822
rect 527 1818 531 1822
rect 567 1818 571 1822
rect 111 1758 115 1762
rect 135 1758 139 1762
rect 183 1758 187 1762
rect 199 1758 203 1762
rect 263 1758 267 1762
rect 295 1758 299 1762
rect 351 1758 355 1762
rect 399 1758 403 1762
rect 439 1758 443 1762
rect 495 1758 499 1762
rect 695 1874 699 1878
rect 703 1874 707 1878
rect 759 1874 763 1878
rect 791 1874 795 1878
rect 1135 1954 1139 1958
rect 1159 1954 1163 1958
rect 1239 1954 1243 1958
rect 1351 1954 1355 1958
rect 1359 1954 1363 1958
rect 1423 1954 1427 1958
rect 1455 1954 1459 1958
rect 1487 1954 1491 1958
rect 1559 1954 1563 1958
rect 911 1930 915 1934
rect 991 1930 995 1934
rect 1095 1930 1099 1934
rect 1135 1902 1139 1906
rect 1231 1902 1235 1906
rect 1271 1902 1275 1906
rect 1319 1902 1323 1906
rect 1359 1902 1363 1906
rect 831 1874 835 1878
rect 879 1874 883 1878
rect 1095 1874 1099 1878
rect 1375 1902 1379 1906
rect 1423 1902 1427 1906
rect 1439 1902 1443 1906
rect 1631 1954 1635 1958
rect 1679 2018 1683 2022
rect 1743 2018 1747 2022
rect 1951 2070 1955 2074
rect 1959 2070 1963 2074
rect 2023 2070 2027 2074
rect 2071 2070 2075 2074
rect 2119 2070 2123 2074
rect 1759 2018 1763 2022
rect 1823 2018 1827 2022
rect 1831 2018 1835 2022
rect 1895 2018 1899 2022
rect 1959 2018 1963 2022
rect 2023 2018 2027 2022
rect 2071 2018 2075 2022
rect 2119 2018 2123 2022
rect 1655 1954 1659 1958
rect 1703 1954 1707 1958
rect 1743 1954 1747 1958
rect 1775 1954 1779 1958
rect 1823 1954 1827 1958
rect 1847 1954 1851 1958
rect 1895 1954 1899 1958
rect 1927 1954 1931 1958
rect 1959 1954 1963 1958
rect 2007 1954 2011 1958
rect 2023 1954 2027 1958
rect 2071 1954 2075 1958
rect 2119 1954 2123 1958
rect 1487 1902 1491 1906
rect 1503 1902 1507 1906
rect 1559 1902 1563 1906
rect 1575 1902 1579 1906
rect 1631 1902 1635 1906
rect 1655 1902 1659 1906
rect 1703 1902 1707 1906
rect 1751 1902 1755 1906
rect 1775 1902 1779 1906
rect 1847 1902 1851 1906
rect 1863 1902 1867 1906
rect 1927 1902 1931 1906
rect 1975 1902 1979 1906
rect 607 1818 611 1822
rect 631 1818 635 1822
rect 687 1818 691 1822
rect 695 1818 699 1822
rect 1135 1846 1139 1850
rect 1159 1846 1163 1850
rect 1199 1846 1203 1850
rect 1231 1846 1235 1850
rect 1239 1846 1243 1850
rect 1271 1846 1275 1850
rect 759 1818 763 1822
rect 767 1818 771 1822
rect 831 1818 835 1822
rect 839 1818 843 1822
rect 911 1818 915 1822
rect 991 1818 995 1822
rect 1047 1818 1051 1822
rect 1095 1818 1099 1822
rect 1303 1846 1307 1850
rect 1319 1846 1323 1850
rect 1367 1846 1371 1850
rect 1375 1846 1379 1850
rect 1431 1846 1435 1850
rect 1439 1846 1443 1850
rect 1503 1846 1507 1850
rect 2007 1902 2011 1906
rect 2071 1902 2075 1906
rect 2119 1902 2123 1906
rect 1575 1846 1579 1850
rect 1583 1846 1587 1850
rect 1655 1846 1659 1850
rect 1671 1846 1675 1850
rect 1751 1846 1755 1850
rect 1767 1846 1771 1850
rect 1863 1846 1867 1850
rect 1871 1846 1875 1850
rect 1975 1846 1979 1850
rect 1983 1846 1987 1850
rect 2071 1846 2075 1850
rect 2119 1846 2123 1850
rect 1439 1808 1443 1812
rect 2007 1808 2011 1812
rect 1135 1786 1139 1790
rect 527 1758 531 1762
rect 591 1758 595 1762
rect 607 1758 611 1762
rect 671 1758 675 1762
rect 687 1758 691 1762
rect 751 1758 755 1762
rect 767 1758 771 1762
rect 823 1758 827 1762
rect 839 1758 843 1762
rect 887 1758 891 1762
rect 911 1758 915 1762
rect 111 1702 115 1706
rect 135 1702 139 1706
rect 151 1702 155 1706
rect 199 1702 203 1706
rect 223 1702 227 1706
rect 295 1702 299 1706
rect 303 1702 307 1706
rect 383 1702 387 1706
rect 399 1702 403 1706
rect 463 1702 467 1706
rect 495 1702 499 1706
rect 535 1702 539 1706
rect 111 1646 115 1650
rect 151 1646 155 1650
rect 175 1646 179 1650
rect 215 1646 219 1650
rect 223 1646 227 1650
rect 255 1646 259 1650
rect 303 1646 307 1650
rect 591 1702 595 1706
rect 607 1702 611 1706
rect 671 1702 675 1706
rect 735 1702 739 1706
rect 751 1702 755 1706
rect 1159 1786 1163 1790
rect 1199 1786 1203 1790
rect 1239 1786 1243 1790
rect 1303 1786 1307 1790
rect 1311 1786 1315 1790
rect 1351 1786 1355 1790
rect 1367 1786 1371 1790
rect 1391 1786 1395 1790
rect 1431 1786 1435 1790
rect 1471 1786 1475 1790
rect 1503 1786 1507 1790
rect 1511 1786 1515 1790
rect 1551 1786 1555 1790
rect 1583 1786 1587 1790
rect 1607 1786 1611 1790
rect 1671 1786 1675 1790
rect 1679 1786 1683 1790
rect 1767 1786 1771 1790
rect 1871 1786 1875 1790
rect 1983 1786 1987 1790
rect 959 1758 963 1762
rect 991 1758 995 1762
rect 1031 1758 1035 1762
rect 1047 1758 1051 1762
rect 1095 1758 1099 1762
rect 1135 1730 1139 1734
rect 1263 1730 1267 1734
rect 1311 1730 1315 1734
rect 1319 1730 1323 1734
rect 2071 1786 2075 1790
rect 2119 1786 2123 1790
rect 1351 1730 1355 1734
rect 1383 1730 1387 1734
rect 1391 1730 1395 1734
rect 1431 1730 1435 1734
rect 1455 1730 1459 1734
rect 1471 1730 1475 1734
rect 1511 1730 1515 1734
rect 1535 1730 1539 1734
rect 1551 1730 1555 1734
rect 1607 1730 1611 1734
rect 1615 1730 1619 1734
rect 1679 1730 1683 1734
rect 1687 1730 1691 1734
rect 1759 1730 1763 1734
rect 1767 1730 1771 1734
rect 1831 1730 1835 1734
rect 1871 1730 1875 1734
rect 1895 1730 1899 1734
rect 1959 1730 1963 1734
rect 1983 1730 1987 1734
rect 2023 1730 2027 1734
rect 2071 1730 2075 1734
rect 807 1702 811 1706
rect 823 1702 827 1706
rect 879 1702 883 1706
rect 887 1702 891 1706
rect 959 1702 963 1706
rect 1031 1702 1035 1706
rect 1095 1702 1099 1706
rect 1135 1678 1139 1682
rect 1167 1678 1171 1682
rect 1247 1678 1251 1682
rect 1263 1678 1267 1682
rect 359 1646 363 1650
rect 383 1646 387 1650
rect 407 1646 411 1650
rect 455 1646 459 1650
rect 463 1646 467 1650
rect 503 1646 507 1650
rect 111 1586 115 1590
rect 143 1586 147 1590
rect 175 1586 179 1590
rect 183 1586 187 1590
rect 215 1586 219 1590
rect 231 1586 235 1590
rect 255 1586 259 1590
rect 287 1586 291 1590
rect 303 1586 307 1590
rect 351 1586 355 1590
rect 359 1586 363 1590
rect 535 1646 539 1650
rect 551 1646 555 1650
rect 607 1646 611 1650
rect 407 1586 411 1590
rect 415 1586 419 1590
rect 455 1586 459 1590
rect 479 1586 483 1590
rect 503 1586 507 1590
rect 663 1646 667 1650
rect 671 1646 675 1650
rect 719 1646 723 1650
rect 735 1646 739 1650
rect 807 1646 811 1650
rect 879 1646 883 1650
rect 1095 1646 1099 1650
rect 1135 1622 1139 1626
rect 1159 1622 1163 1626
rect 1167 1622 1171 1626
rect 543 1586 547 1590
rect 551 1586 555 1590
rect 607 1586 611 1590
rect 111 1526 115 1530
rect 135 1526 139 1530
rect 143 1526 147 1530
rect 175 1526 179 1530
rect 183 1526 187 1530
rect 215 1526 219 1530
rect 231 1526 235 1530
rect 255 1526 259 1530
rect 287 1526 291 1530
rect 295 1526 299 1530
rect 335 1526 339 1530
rect 351 1526 355 1530
rect 375 1526 379 1530
rect 415 1526 419 1530
rect 455 1526 459 1530
rect 479 1526 483 1530
rect 495 1526 499 1530
rect 535 1526 539 1530
rect 543 1526 547 1530
rect 663 1586 667 1590
rect 719 1586 723 1590
rect 727 1586 731 1590
rect 791 1586 795 1590
rect 855 1586 859 1590
rect 1095 1586 1099 1590
rect 1319 1678 1323 1682
rect 1335 1678 1339 1682
rect 1383 1678 1387 1682
rect 1423 1678 1427 1682
rect 1455 1678 1459 1682
rect 1511 1678 1515 1682
rect 1535 1678 1539 1682
rect 1599 1678 1603 1682
rect 1615 1678 1619 1682
rect 1679 1678 1683 1682
rect 1687 1678 1691 1682
rect 1751 1678 1755 1682
rect 1759 1678 1763 1682
rect 1815 1678 1819 1682
rect 1831 1678 1835 1682
rect 1871 1678 1875 1682
rect 1895 1678 1899 1682
rect 1927 1678 1931 1682
rect 1959 1678 1963 1682
rect 1983 1678 1987 1682
rect 2023 1678 2027 1682
rect 2031 1678 2035 1682
rect 2071 1678 2075 1682
rect 2119 1730 2123 1734
rect 2119 1678 2123 1682
rect 1199 1622 1203 1626
rect 1247 1622 1251 1626
rect 1319 1622 1323 1626
rect 1335 1622 1339 1626
rect 1391 1622 1395 1626
rect 1423 1622 1427 1626
rect 1463 1622 1467 1626
rect 1511 1622 1515 1626
rect 1535 1622 1539 1626
rect 1599 1622 1603 1626
rect 1607 1622 1611 1626
rect 1679 1622 1683 1626
rect 1135 1570 1139 1574
rect 1159 1570 1163 1574
rect 1199 1570 1203 1574
rect 1239 1570 1243 1574
rect 1247 1570 1251 1574
rect 1279 1570 1283 1574
rect 1319 1570 1323 1574
rect 1327 1570 1331 1574
rect 575 1526 579 1530
rect 607 1526 611 1530
rect 615 1526 619 1530
rect 655 1526 659 1530
rect 663 1526 667 1530
rect 695 1526 699 1530
rect 727 1526 731 1530
rect 735 1526 739 1530
rect 775 1526 779 1530
rect 791 1526 795 1530
rect 831 1526 835 1530
rect 111 1466 115 1470
rect 135 1466 139 1470
rect 175 1466 179 1470
rect 215 1466 219 1470
rect 255 1466 259 1470
rect 295 1466 299 1470
rect 335 1466 339 1470
rect 375 1466 379 1470
rect 415 1466 419 1470
rect 455 1466 459 1470
rect 495 1466 499 1470
rect 519 1466 523 1470
rect 535 1466 539 1470
rect 1259 1544 1263 1548
rect 1375 1570 1379 1574
rect 1391 1570 1395 1574
rect 1423 1570 1427 1574
rect 1463 1570 1467 1574
rect 1471 1570 1475 1574
rect 1519 1570 1523 1574
rect 1535 1570 1539 1574
rect 1399 1544 1403 1548
rect 855 1526 859 1530
rect 887 1526 891 1530
rect 1095 1526 1099 1530
rect 1135 1514 1139 1518
rect 1239 1514 1243 1518
rect 1279 1514 1283 1518
rect 1319 1514 1323 1518
rect 1327 1514 1331 1518
rect 1359 1514 1363 1518
rect 1375 1514 1379 1518
rect 1399 1514 1403 1518
rect 1423 1514 1427 1518
rect 1567 1570 1571 1574
rect 1607 1570 1611 1574
rect 1623 1570 1627 1574
rect 1751 1622 1755 1626
rect 1815 1622 1819 1626
rect 1831 1622 1835 1626
rect 1871 1622 1875 1626
rect 1927 1622 1931 1626
rect 1983 1622 1987 1626
rect 2031 1622 2035 1626
rect 2071 1622 2075 1626
rect 2119 1622 2123 1626
rect 1679 1570 1683 1574
rect 1735 1570 1739 1574
rect 1751 1570 1755 1574
rect 1831 1570 1835 1574
rect 2119 1570 2123 1574
rect 1439 1514 1443 1518
rect 1471 1514 1475 1518
rect 1479 1514 1483 1518
rect 1519 1514 1523 1518
rect 559 1466 563 1470
rect 575 1466 579 1470
rect 599 1466 603 1470
rect 615 1466 619 1470
rect 647 1466 651 1470
rect 655 1466 659 1470
rect 695 1466 699 1470
rect 735 1466 739 1470
rect 751 1466 755 1470
rect 775 1466 779 1470
rect 807 1466 811 1470
rect 831 1466 835 1470
rect 871 1466 875 1470
rect 887 1466 891 1470
rect 111 1410 115 1414
rect 431 1410 435 1414
rect 471 1410 475 1414
rect 519 1410 523 1414
rect 559 1410 563 1414
rect 575 1410 579 1414
rect 599 1410 603 1414
rect 631 1410 635 1414
rect 647 1410 651 1414
rect 935 1466 939 1470
rect 1095 1466 1099 1470
rect 1559 1514 1563 1518
rect 1567 1514 1571 1518
rect 1607 1514 1611 1518
rect 1623 1514 1627 1518
rect 1663 1514 1667 1518
rect 1679 1514 1683 1518
rect 1735 1514 1739 1518
rect 1815 1514 1819 1518
rect 1903 1514 1907 1518
rect 1991 1514 1995 1518
rect 2071 1514 2075 1518
rect 2119 1514 2123 1518
rect 1591 1472 1595 1476
rect 1135 1462 1139 1466
rect 1231 1462 1235 1466
rect 1279 1462 1283 1466
rect 1319 1462 1323 1466
rect 695 1410 699 1414
rect 751 1410 755 1414
rect 759 1410 763 1414
rect 807 1410 811 1414
rect 823 1410 827 1414
rect 111 1358 115 1362
rect 375 1358 379 1362
rect 423 1358 427 1362
rect 431 1358 435 1362
rect 111 1306 115 1310
rect 335 1306 339 1310
rect 375 1306 379 1310
rect 471 1358 475 1362
rect 479 1358 483 1362
rect 519 1358 523 1362
rect 543 1358 547 1362
rect 575 1358 579 1362
rect 607 1358 611 1362
rect 631 1358 635 1362
rect 671 1358 675 1362
rect 695 1358 699 1362
rect 871 1410 875 1414
rect 895 1410 899 1414
rect 935 1410 939 1414
rect 967 1410 971 1414
rect 1095 1410 1099 1414
rect 1135 1406 1139 1410
rect 1159 1406 1163 1410
rect 1199 1406 1203 1410
rect 1231 1406 1235 1410
rect 1335 1462 1339 1466
rect 1359 1462 1363 1466
rect 1391 1462 1395 1466
rect 1399 1462 1403 1466
rect 1439 1462 1443 1466
rect 1455 1462 1459 1466
rect 1479 1462 1483 1466
rect 1519 1462 1523 1466
rect 1559 1462 1563 1466
rect 1583 1462 1587 1466
rect 1327 1440 1331 1444
rect 1911 1472 1915 1476
rect 1607 1462 1611 1466
rect 1647 1462 1651 1466
rect 1663 1462 1667 1466
rect 1719 1462 1723 1466
rect 1735 1462 1739 1466
rect 1807 1462 1811 1466
rect 1815 1462 1819 1466
rect 1895 1462 1899 1466
rect 1903 1462 1907 1466
rect 1991 1462 1995 1466
rect 1543 1440 1547 1444
rect 1263 1406 1267 1410
rect 1279 1406 1283 1410
rect 1335 1406 1339 1410
rect 1351 1406 1355 1410
rect 1391 1406 1395 1410
rect 1447 1406 1451 1410
rect 1455 1406 1459 1410
rect 1519 1406 1523 1410
rect 1543 1406 1547 1410
rect 1583 1406 1587 1410
rect 1631 1406 1635 1410
rect 1647 1406 1651 1410
rect 1719 1406 1723 1410
rect 1799 1406 1803 1410
rect 1807 1406 1811 1410
rect 1871 1406 1875 1410
rect 1895 1406 1899 1410
rect 735 1358 739 1362
rect 759 1358 763 1362
rect 799 1358 803 1362
rect 823 1358 827 1362
rect 863 1358 867 1362
rect 895 1358 899 1362
rect 927 1358 931 1362
rect 967 1358 971 1362
rect 999 1358 1003 1362
rect 1047 1358 1051 1362
rect 1095 1358 1099 1362
rect 391 1306 395 1310
rect 423 1306 427 1310
rect 455 1306 459 1310
rect 479 1306 483 1310
rect 527 1306 531 1310
rect 543 1306 547 1310
rect 599 1306 603 1310
rect 607 1306 611 1310
rect 671 1306 675 1310
rect 735 1306 739 1310
rect 743 1306 747 1310
rect 799 1306 803 1310
rect 823 1306 827 1310
rect 111 1250 115 1254
rect 263 1250 267 1254
rect 311 1250 315 1254
rect 335 1250 339 1254
rect 359 1250 363 1254
rect 391 1250 395 1254
rect 415 1250 419 1254
rect 455 1250 459 1254
rect 479 1250 483 1254
rect 527 1250 531 1254
rect 543 1250 547 1254
rect 599 1250 603 1254
rect 111 1198 115 1202
rect 223 1198 227 1202
rect 263 1198 267 1202
rect 607 1250 611 1254
rect 671 1250 675 1254
rect 735 1250 739 1254
rect 743 1250 747 1254
rect 863 1306 867 1310
rect 903 1306 907 1310
rect 927 1306 931 1310
rect 799 1250 803 1254
rect 823 1250 827 1254
rect 863 1250 867 1254
rect 903 1250 907 1254
rect 983 1306 987 1310
rect 999 1306 1003 1310
rect 1047 1306 1051 1310
rect 1671 1368 1675 1372
rect 1135 1350 1139 1354
rect 1159 1350 1163 1354
rect 1199 1350 1203 1354
rect 1255 1350 1259 1354
rect 1263 1350 1267 1354
rect 1351 1350 1355 1354
rect 1375 1350 1379 1354
rect 1447 1350 1451 1354
rect 1487 1350 1491 1354
rect 1543 1350 1547 1354
rect 1591 1350 1595 1354
rect 1631 1350 1635 1354
rect 1679 1350 1683 1354
rect 1719 1350 1723 1354
rect 1759 1350 1763 1354
rect 1799 1350 1803 1354
rect 1831 1350 1835 1354
rect 1871 1350 1875 1354
rect 1943 1406 1947 1410
rect 1991 1406 1995 1410
rect 2015 1406 2019 1410
rect 2071 1462 2075 1466
rect 2119 1462 2123 1466
rect 2071 1406 2075 1410
rect 1931 1368 1935 1372
rect 1903 1350 1907 1354
rect 1943 1350 1947 1354
rect 1967 1350 1971 1354
rect 2015 1350 2019 1354
rect 2031 1350 2035 1354
rect 2071 1350 2075 1354
rect 1095 1306 1099 1310
rect 1135 1294 1139 1298
rect 1159 1294 1163 1298
rect 1199 1294 1203 1298
rect 1247 1294 1251 1298
rect 1255 1294 1259 1298
rect 1319 1294 1323 1298
rect 1375 1294 1379 1298
rect 1399 1294 1403 1298
rect 1479 1294 1483 1298
rect 1487 1294 1491 1298
rect 1559 1294 1563 1298
rect 1591 1294 1595 1298
rect 1639 1294 1643 1298
rect 1679 1294 1683 1298
rect 1719 1294 1723 1298
rect 1759 1294 1763 1298
rect 1799 1294 1803 1298
rect 1831 1294 1835 1298
rect 1879 1294 1883 1298
rect 1903 1294 1907 1298
rect 927 1250 931 1254
rect 983 1250 987 1254
rect 1047 1250 1051 1254
rect 1095 1250 1099 1254
rect 1135 1238 1139 1242
rect 1159 1238 1163 1242
rect 1199 1238 1203 1242
rect 1239 1238 1243 1242
rect 1247 1238 1251 1242
rect 279 1198 283 1202
rect 311 1198 315 1202
rect 343 1198 347 1202
rect 359 1198 363 1202
rect 407 1198 411 1202
rect 415 1198 419 1202
rect 479 1198 483 1202
rect 543 1198 547 1202
rect 551 1198 555 1202
rect 111 1146 115 1150
rect 159 1146 163 1150
rect 199 1146 203 1150
rect 223 1146 227 1150
rect 607 1198 611 1202
rect 631 1198 635 1202
rect 671 1198 675 1202
rect 711 1198 715 1202
rect 735 1198 739 1202
rect 791 1198 795 1202
rect 799 1198 803 1202
rect 863 1198 867 1202
rect 871 1198 875 1202
rect 247 1146 251 1150
rect 111 1086 115 1090
rect 159 1086 163 1090
rect 279 1146 283 1150
rect 303 1146 307 1150
rect 343 1146 347 1150
rect 367 1146 371 1150
rect 407 1146 411 1150
rect 439 1146 443 1150
rect 479 1146 483 1150
rect 511 1146 515 1150
rect 551 1146 555 1150
rect 591 1146 595 1150
rect 631 1146 635 1150
rect 679 1146 683 1150
rect 711 1146 715 1150
rect 775 1146 779 1150
rect 791 1146 795 1150
rect 1279 1238 1283 1242
rect 1319 1238 1323 1242
rect 1327 1238 1331 1242
rect 1375 1238 1379 1242
rect 1399 1238 1403 1242
rect 1423 1238 1427 1242
rect 1471 1238 1475 1242
rect 927 1198 931 1202
rect 959 1198 963 1202
rect 1095 1198 1099 1202
rect 1135 1186 1139 1190
rect 1159 1186 1163 1190
rect 1199 1186 1203 1190
rect 1239 1186 1243 1190
rect 1279 1186 1283 1190
rect 1287 1186 1291 1190
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1375 1186 1379 1190
rect 871 1146 875 1150
rect 879 1146 883 1150
rect 959 1146 963 1150
rect 1479 1238 1483 1242
rect 1535 1238 1539 1242
rect 1559 1238 1563 1242
rect 1415 1186 1419 1190
rect 1423 1186 1427 1190
rect 1471 1186 1475 1190
rect 1527 1186 1531 1190
rect 1535 1186 1539 1190
rect 1615 1238 1619 1242
rect 1639 1238 1643 1242
rect 1719 1238 1723 1242
rect 1799 1238 1803 1242
rect 1967 1294 1971 1298
rect 2031 1294 2035 1298
rect 2119 1406 2123 1410
rect 2119 1350 2123 1354
rect 2055 1294 2059 1298
rect 2071 1294 2075 1298
rect 1839 1238 1843 1242
rect 1879 1238 1883 1242
rect 1967 1238 1971 1242
rect 1583 1186 1587 1190
rect 1615 1186 1619 1190
rect 1639 1186 1643 1190
rect 991 1146 995 1150
rect 1095 1146 1099 1150
rect 1135 1126 1139 1130
rect 1287 1126 1291 1130
rect 1327 1126 1331 1130
rect 1367 1126 1371 1130
rect 1383 1126 1387 1130
rect 1415 1126 1419 1130
rect 1423 1126 1427 1130
rect 1471 1126 1475 1130
rect 199 1086 203 1090
rect 247 1086 251 1090
rect 303 1086 307 1090
rect 367 1086 371 1090
rect 431 1086 435 1090
rect 439 1086 443 1090
rect 503 1086 507 1090
rect 511 1086 515 1090
rect 111 1030 115 1034
rect 199 1030 203 1034
rect 223 1030 227 1034
rect 247 1030 251 1034
rect 271 1030 275 1034
rect 303 1030 307 1034
rect 335 1030 339 1034
rect 367 1030 371 1034
rect 407 1030 411 1034
rect 111 974 115 978
rect 151 974 155 978
rect 215 974 219 978
rect 223 974 227 978
rect 575 1086 579 1090
rect 591 1086 595 1090
rect 647 1086 651 1090
rect 679 1086 683 1090
rect 719 1086 723 1090
rect 775 1086 779 1090
rect 783 1086 787 1090
rect 431 1030 435 1034
rect 479 1030 483 1034
rect 503 1030 507 1034
rect 559 1030 563 1034
rect 575 1030 579 1034
rect 631 1030 635 1034
rect 647 1030 651 1034
rect 1703 1186 1707 1190
rect 1719 1186 1723 1190
rect 1767 1186 1771 1190
rect 1839 1186 1843 1190
rect 1919 1186 1923 1190
rect 1967 1186 1971 1190
rect 2007 1186 2011 1190
rect 2055 1238 2059 1242
rect 2071 1238 2075 1242
rect 2119 1294 2123 1298
rect 2119 1238 2123 1242
rect 2071 1186 2075 1190
rect 1527 1126 1531 1130
rect 1583 1126 1587 1130
rect 1591 1126 1595 1130
rect 1639 1126 1643 1130
rect 1655 1126 1659 1130
rect 1703 1126 1707 1130
rect 1399 1096 1403 1100
rect 1551 1099 1555 1100
rect 1551 1096 1555 1099
rect 839 1086 843 1090
rect 879 1086 883 1090
rect 895 1086 899 1090
rect 951 1086 955 1090
rect 991 1086 995 1090
rect 1007 1086 1011 1090
rect 1047 1086 1051 1090
rect 1095 1086 1099 1090
rect 1135 1074 1139 1078
rect 1159 1074 1163 1078
rect 1247 1074 1251 1078
rect 1359 1074 1363 1078
rect 1383 1074 1387 1078
rect 1423 1074 1427 1078
rect 1471 1074 1475 1078
rect 1527 1074 1531 1078
rect 1575 1074 1579 1078
rect 1591 1074 1595 1078
rect 703 1030 707 1034
rect 719 1030 723 1034
rect 775 1030 779 1034
rect 783 1030 787 1034
rect 839 1030 843 1034
rect 895 1030 899 1034
rect 903 1030 907 1034
rect 271 974 275 978
rect 287 974 291 978
rect 335 974 339 978
rect 367 974 371 978
rect 407 974 411 978
rect 447 974 451 978
rect 479 974 483 978
rect 111 922 115 926
rect 135 922 139 926
rect 151 922 155 926
rect 183 922 187 926
rect 215 922 219 926
rect 255 922 259 926
rect 287 922 291 926
rect 327 922 331 926
rect 367 922 371 926
rect 399 922 403 926
rect 447 922 451 926
rect 463 922 467 926
rect 111 866 115 870
rect 135 866 139 870
rect 175 866 179 870
rect 183 866 187 870
rect 215 866 219 870
rect 255 866 259 870
rect 279 866 283 870
rect 527 974 531 978
rect 559 974 563 978
rect 599 974 603 978
rect 631 974 635 978
rect 671 974 675 978
rect 703 974 707 978
rect 951 1030 955 1034
rect 967 1030 971 1034
rect 1007 1030 1011 1034
rect 1039 1030 1043 1034
rect 1047 1030 1051 1034
rect 1711 1126 1715 1130
rect 1767 1126 1771 1130
rect 1823 1126 1827 1130
rect 1839 1126 1843 1130
rect 1871 1126 1875 1130
rect 1919 1126 1923 1130
rect 1927 1126 1931 1130
rect 1983 1126 1987 1130
rect 2007 1126 2011 1130
rect 2031 1126 2035 1130
rect 1655 1074 1659 1078
rect 1671 1074 1675 1078
rect 1711 1074 1715 1078
rect 1759 1074 1763 1078
rect 1767 1074 1771 1078
rect 1823 1074 1827 1078
rect 1847 1074 1851 1078
rect 1871 1074 1875 1078
rect 1927 1074 1931 1078
rect 1983 1074 1987 1078
rect 1095 1030 1099 1034
rect 1135 1022 1139 1026
rect 1159 1022 1163 1026
rect 1231 1022 1235 1026
rect 1247 1022 1251 1026
rect 1303 1022 1307 1026
rect 1359 1022 1363 1026
rect 1383 1022 1387 1026
rect 1463 1022 1467 1026
rect 1471 1022 1475 1026
rect 735 974 739 978
rect 775 974 779 978
rect 799 974 803 978
rect 839 974 843 978
rect 863 974 867 978
rect 903 974 907 978
rect 927 974 931 978
rect 967 974 971 978
rect 991 974 995 978
rect 1039 974 1043 978
rect 1047 974 1051 978
rect 527 922 531 926
rect 599 922 603 926
rect 327 866 331 870
rect 343 866 347 870
rect 111 814 115 818
rect 399 866 403 870
rect 463 866 467 870
rect 527 866 531 870
rect 535 866 539 870
rect 671 922 675 926
rect 735 922 739 926
rect 743 922 747 926
rect 799 922 803 926
rect 815 922 819 926
rect 863 922 867 926
rect 895 922 899 926
rect 927 922 931 926
rect 983 922 987 926
rect 991 922 995 926
rect 1543 1022 1547 1026
rect 1575 1022 1579 1026
rect 1623 1022 1627 1026
rect 1671 1022 1675 1026
rect 1695 1022 1699 1026
rect 1759 1022 1763 1026
rect 1095 974 1099 978
rect 1135 970 1139 974
rect 1159 970 1163 974
rect 1231 970 1235 974
rect 1239 970 1243 974
rect 1303 970 1307 974
rect 1047 922 1051 926
rect 1095 922 1099 926
rect 1375 970 1379 974
rect 1383 970 1387 974
rect 1439 970 1443 974
rect 1463 970 1467 974
rect 1511 970 1515 974
rect 2007 1074 2011 1078
rect 2031 1074 2035 1078
rect 2071 1126 2075 1130
rect 2119 1186 2123 1190
rect 2119 1126 2123 1130
rect 2071 1074 2075 1078
rect 2119 1074 2123 1078
rect 1823 1022 1827 1026
rect 1847 1022 1851 1026
rect 1887 1022 1891 1026
rect 1927 1022 1931 1026
rect 1951 1022 1955 1026
rect 2007 1022 2011 1026
rect 2071 1022 2075 1026
rect 2119 1022 2123 1026
rect 1543 970 1547 974
rect 1583 970 1587 974
rect 1623 970 1627 974
rect 1655 970 1659 974
rect 1695 970 1699 974
rect 1727 970 1731 974
rect 1759 970 1763 974
rect 1135 914 1139 918
rect 1239 914 1243 918
rect 1287 914 1291 918
rect 1303 914 1307 918
rect 1327 914 1331 918
rect 1375 914 1379 918
rect 599 866 603 870
rect 615 866 619 870
rect 671 866 675 870
rect 711 866 715 870
rect 743 866 747 870
rect 815 866 819 870
rect 823 866 827 870
rect 895 866 899 870
rect 943 866 947 870
rect 983 866 987 870
rect 1047 866 1051 870
rect 547 848 551 852
rect 847 848 851 852
rect 135 814 139 818
rect 175 814 179 818
rect 215 814 219 818
rect 279 814 283 818
rect 335 814 339 818
rect 343 814 347 818
rect 391 814 395 818
rect 399 814 403 818
rect 111 762 115 766
rect 135 762 139 766
rect 455 814 459 818
rect 463 814 467 818
rect 479 824 483 828
rect 519 814 523 818
rect 535 814 539 818
rect 859 824 863 828
rect 583 814 587 818
rect 615 814 619 818
rect 655 814 659 818
rect 711 814 715 818
rect 735 814 739 818
rect 815 814 819 818
rect 823 814 827 818
rect 175 762 179 766
rect 207 762 211 766
rect 215 762 219 766
rect 279 762 283 766
rect 295 762 299 766
rect 335 762 339 766
rect 375 762 379 766
rect 391 762 395 766
rect 447 762 451 766
rect 455 762 459 766
rect 519 762 523 766
rect 111 706 115 710
rect 135 706 139 710
rect 183 706 187 710
rect 207 706 211 710
rect 247 706 251 710
rect 295 706 299 710
rect 311 706 315 710
rect 111 646 115 650
rect 135 646 139 650
rect 159 646 163 650
rect 183 646 187 650
rect 215 646 219 650
rect 375 706 379 710
rect 383 706 387 710
rect 583 762 587 766
rect 639 762 643 766
rect 655 762 659 766
rect 687 762 691 766
rect 895 814 899 818
rect 1423 914 1427 918
rect 1439 914 1443 918
rect 1479 914 1483 918
rect 1511 914 1515 918
rect 1551 914 1555 918
rect 1583 914 1587 918
rect 1623 914 1627 918
rect 1655 914 1659 918
rect 1703 914 1707 918
rect 1727 914 1731 918
rect 1095 866 1099 870
rect 1135 862 1139 866
rect 1159 862 1163 866
rect 1199 862 1203 866
rect 943 814 947 818
rect 983 814 987 818
rect 1047 814 1051 818
rect 1095 814 1099 818
rect 1263 862 1267 866
rect 1287 862 1291 866
rect 1327 862 1331 866
rect 1375 862 1379 866
rect 1399 862 1403 866
rect 1423 862 1427 866
rect 1471 862 1475 866
rect 1479 862 1483 866
rect 1799 970 1803 974
rect 1823 970 1827 974
rect 1871 970 1875 974
rect 1887 970 1891 974
rect 1943 970 1947 974
rect 1951 970 1955 974
rect 2015 970 2019 974
rect 2071 970 2075 974
rect 2119 970 2123 974
rect 1791 914 1795 918
rect 1799 914 1803 918
rect 1871 914 1875 918
rect 1879 914 1883 918
rect 1943 914 1947 918
rect 1967 914 1971 918
rect 1543 862 1547 866
rect 1551 862 1555 866
rect 1623 862 1627 866
rect 1703 862 1707 866
rect 1775 862 1779 866
rect 1791 862 1795 866
rect 1855 862 1859 866
rect 1879 862 1883 866
rect 1935 862 1939 866
rect 1967 862 1971 866
rect 1135 802 1139 806
rect 1159 802 1163 806
rect 1199 802 1203 806
rect 1239 802 1243 806
rect 1263 802 1267 806
rect 1327 802 1331 806
rect 1343 802 1347 806
rect 1399 802 1403 806
rect 1447 802 1451 806
rect 1471 802 1475 806
rect 1543 802 1547 806
rect 1551 802 1555 806
rect 1623 802 1627 806
rect 1655 802 1659 806
rect 1703 802 1707 806
rect 1751 802 1755 806
rect 1775 802 1779 806
rect 2015 914 2019 918
rect 2063 914 2067 918
rect 2071 914 2075 918
rect 2119 914 2123 918
rect 2015 862 2019 866
rect 2063 862 2067 866
rect 2071 862 2075 866
rect 2119 862 2123 866
rect 1839 802 1843 806
rect 1855 802 1859 806
rect 1919 802 1923 806
rect 1935 802 1939 806
rect 735 762 739 766
rect 743 762 747 766
rect 799 762 803 766
rect 815 762 819 766
rect 855 762 859 766
rect 895 762 899 766
rect 983 762 987 766
rect 1047 762 1051 766
rect 1095 762 1099 766
rect 1135 750 1139 754
rect 1159 750 1163 754
rect 1199 750 1203 754
rect 1239 750 1243 754
rect 1287 750 1291 754
rect 447 706 451 710
rect 455 706 459 710
rect 519 706 523 710
rect 583 706 587 710
rect 639 706 643 710
rect 647 706 651 710
rect 687 706 691 710
rect 711 706 715 710
rect 743 706 747 710
rect 767 706 771 710
rect 247 646 251 650
rect 111 590 115 594
rect 159 590 163 594
rect 207 590 211 594
rect 215 590 219 594
rect 255 590 259 594
rect 287 646 291 650
rect 311 646 315 650
rect 367 646 371 650
rect 383 646 387 650
rect 455 646 459 650
rect 519 646 523 650
rect 287 590 291 594
rect 311 590 315 594
rect 367 590 371 594
rect 383 590 387 594
rect 111 530 115 534
rect 159 530 163 534
rect 167 530 171 534
rect 207 530 211 534
rect 223 530 227 534
rect 111 478 115 482
rect 167 478 171 482
rect 255 530 259 534
rect 287 530 291 534
rect 311 530 315 534
rect 359 530 363 534
rect 543 646 547 650
rect 583 646 587 650
rect 631 646 635 650
rect 647 646 651 650
rect 735 680 739 684
rect 799 706 803 710
rect 823 706 827 710
rect 855 706 859 710
rect 879 706 883 710
rect 943 706 947 710
rect 1095 706 1099 710
rect 711 646 715 650
rect 719 646 723 650
rect 767 646 771 650
rect 799 646 803 650
rect 1343 750 1347 754
rect 1359 750 1363 754
rect 1439 750 1443 754
rect 1447 750 1451 754
rect 1135 694 1139 698
rect 1159 694 1163 698
rect 1199 694 1203 698
rect 1239 694 1243 698
rect 1287 694 1291 698
rect 1335 694 1339 698
rect 967 680 971 684
rect 1527 750 1531 754
rect 1551 750 1555 754
rect 1615 750 1619 754
rect 1655 750 1659 754
rect 1711 750 1715 754
rect 1751 750 1755 754
rect 1807 750 1811 754
rect 2007 802 2011 806
rect 2015 802 2019 806
rect 2071 802 2075 806
rect 2119 802 2123 806
rect 1839 750 1843 754
rect 1903 750 1907 754
rect 1919 750 1923 754
rect 1999 750 2003 754
rect 2007 750 2011 754
rect 2071 750 2075 754
rect 1359 694 1363 698
rect 1391 694 1395 698
rect 1439 694 1443 698
rect 1447 694 1451 698
rect 1511 694 1515 698
rect 1527 694 1531 698
rect 1575 694 1579 698
rect 1615 694 1619 698
rect 1639 694 1643 698
rect 1703 694 1707 698
rect 1711 694 1715 698
rect 1767 694 1771 698
rect 1807 694 1811 698
rect 1831 694 1835 698
rect 1895 694 1899 698
rect 1903 694 1907 698
rect 1959 694 1963 698
rect 823 646 827 650
rect 871 646 875 650
rect 879 646 883 650
rect 943 646 947 650
rect 951 646 955 650
rect 1031 646 1035 650
rect 1095 646 1099 650
rect 1135 642 1139 646
rect 1239 642 1243 646
rect 455 590 459 594
rect 463 590 467 594
rect 543 590 547 594
rect 623 590 627 594
rect 631 590 635 594
rect 727 608 731 612
rect 703 590 707 594
rect 719 590 723 594
rect 783 590 787 594
rect 799 590 803 594
rect 855 590 859 594
rect 871 590 875 594
rect 383 530 387 534
rect 431 530 435 534
rect 463 530 467 534
rect 511 530 515 534
rect 543 530 547 534
rect 223 478 227 482
rect 231 478 235 482
rect 287 478 291 482
rect 303 478 307 482
rect 359 478 363 482
rect 375 478 379 482
rect 111 426 115 430
rect 151 426 155 430
rect 167 426 171 430
rect 215 426 219 430
rect 231 426 235 430
rect 279 426 283 430
rect 591 530 595 534
rect 623 530 627 534
rect 663 530 667 534
rect 1039 608 1043 612
rect 1279 642 1283 646
rect 1287 642 1291 646
rect 1319 642 1323 646
rect 1335 642 1339 646
rect 1367 642 1371 646
rect 1391 642 1395 646
rect 1423 642 1427 646
rect 1447 642 1451 646
rect 927 590 931 594
rect 951 590 955 594
rect 999 590 1003 594
rect 1031 590 1035 594
rect 1047 590 1051 594
rect 1095 590 1099 594
rect 1135 590 1139 594
rect 1279 590 1283 594
rect 1319 590 1323 594
rect 1335 590 1339 594
rect 703 530 707 534
rect 735 530 739 534
rect 783 530 787 534
rect 807 530 811 534
rect 855 530 859 534
rect 871 530 875 534
rect 927 530 931 534
rect 935 530 939 534
rect 999 530 1003 534
rect 1047 530 1051 534
rect 431 478 435 482
rect 455 478 459 482
rect 511 478 515 482
rect 535 478 539 482
rect 591 478 595 482
rect 607 478 611 482
rect 303 426 307 430
rect 351 426 355 430
rect 375 426 379 430
rect 423 426 427 430
rect 455 426 459 430
rect 487 426 491 430
rect 111 374 115 378
rect 135 374 139 378
rect 151 374 155 378
rect 175 374 179 378
rect 215 374 219 378
rect 271 374 275 378
rect 279 374 283 378
rect 335 374 339 378
rect 351 374 355 378
rect 535 426 539 430
rect 551 426 555 430
rect 663 478 667 482
rect 679 478 683 482
rect 735 478 739 482
rect 743 478 747 482
rect 799 478 803 482
rect 807 478 811 482
rect 855 478 859 482
rect 871 478 875 482
rect 903 478 907 482
rect 935 478 939 482
rect 959 478 963 482
rect 607 426 611 430
rect 615 426 619 430
rect 671 426 675 430
rect 679 426 683 430
rect 1479 642 1483 646
rect 1511 642 1515 646
rect 1535 642 1539 646
rect 1575 642 1579 646
rect 1591 642 1595 646
rect 1639 642 1643 646
rect 1647 642 1651 646
rect 1703 642 1707 646
rect 1999 694 2003 698
rect 2023 694 2027 698
rect 2071 694 2075 698
rect 2119 750 2123 754
rect 2119 694 2123 698
rect 1719 642 1723 646
rect 1767 642 1771 646
rect 1799 642 1803 646
rect 1831 642 1835 646
rect 1879 642 1883 646
rect 1895 642 1899 646
rect 1959 642 1963 646
rect 1967 642 1971 646
rect 2023 642 2027 646
rect 1367 590 1371 594
rect 1375 590 1379 594
rect 1415 590 1419 594
rect 1423 590 1427 594
rect 1463 590 1467 594
rect 1479 590 1483 594
rect 1519 590 1523 594
rect 1535 590 1539 594
rect 1583 590 1587 594
rect 2063 642 2067 646
rect 2071 642 2075 646
rect 2119 642 2123 646
rect 1591 590 1595 594
rect 1647 590 1651 594
rect 1655 590 1659 594
rect 1719 590 1723 594
rect 1727 590 1731 594
rect 1799 590 1803 594
rect 1807 590 1811 594
rect 1879 590 1883 594
rect 1887 590 1891 594
rect 1967 590 1971 594
rect 1975 590 1979 594
rect 2063 590 2067 594
rect 1095 530 1099 534
rect 1135 534 1139 538
rect 1191 534 1195 538
rect 1239 534 1243 538
rect 1287 534 1291 538
rect 1335 534 1339 538
rect 1343 534 1347 538
rect 1375 534 1379 538
rect 1407 534 1411 538
rect 1415 534 1419 538
rect 1463 534 1467 538
rect 1479 534 1483 538
rect 999 478 1003 482
rect 1007 478 1011 482
rect 1047 478 1051 482
rect 1095 478 1099 482
rect 1135 482 1139 486
rect 1159 482 1163 486
rect 1191 482 1195 486
rect 1239 482 1243 486
rect 1263 482 1267 486
rect 1287 482 1291 486
rect 1343 482 1347 486
rect 1519 534 1523 538
rect 1543 534 1547 538
rect 1583 534 1587 538
rect 1607 534 1611 538
rect 1655 534 1659 538
rect 1671 534 1675 538
rect 1727 534 1731 538
rect 1735 534 1739 538
rect 1799 534 1803 538
rect 1807 534 1811 538
rect 1863 534 1867 538
rect 1383 482 1387 486
rect 1407 482 1411 486
rect 1479 482 1483 486
rect 1495 482 1499 486
rect 1543 482 1547 486
rect 1599 482 1603 486
rect 1607 482 1611 486
rect 1671 482 1675 486
rect 2119 590 2123 594
rect 1887 534 1891 538
rect 1935 534 1939 538
rect 1975 534 1979 538
rect 1703 482 1707 486
rect 2007 534 2011 538
rect 2063 534 2067 538
rect 2071 534 2075 538
rect 2119 534 2123 538
rect 1735 482 1739 486
rect 1799 482 1803 486
rect 1863 482 1867 486
rect 1887 482 1891 486
rect 1935 482 1939 486
rect 727 426 731 430
rect 743 426 747 430
rect 791 426 795 430
rect 799 426 803 430
rect 855 426 859 430
rect 903 426 907 430
rect 959 426 963 430
rect 1007 426 1011 430
rect 1047 426 1051 430
rect 1095 426 1099 430
rect 1135 430 1139 434
rect 1159 430 1163 434
rect 1199 430 1203 434
rect 1255 430 1259 434
rect 1263 430 1267 434
rect 1335 430 1339 434
rect 1383 430 1387 434
rect 1415 430 1419 434
rect 1495 430 1499 434
rect 1503 430 1507 434
rect 1591 430 1595 434
rect 1599 430 1603 434
rect 1671 430 1675 434
rect 1703 430 1707 434
rect 1751 430 1755 434
rect 1799 430 1803 434
rect 1823 430 1827 434
rect 1983 482 1987 486
rect 2007 482 2011 486
rect 2071 482 2075 486
rect 2119 482 2123 486
rect 1887 430 1891 434
rect 1951 430 1955 434
rect 1983 430 1987 434
rect 2023 430 2027 434
rect 399 374 403 378
rect 423 374 427 378
rect 463 374 467 378
rect 487 374 491 378
rect 519 374 523 378
rect 111 318 115 322
rect 135 318 139 322
rect 175 318 179 322
rect 207 318 211 322
rect 215 318 219 322
rect 271 318 275 322
rect 295 318 299 322
rect 335 318 339 322
rect 383 318 387 322
rect 399 318 403 322
rect 551 374 555 378
rect 575 374 579 378
rect 615 374 619 378
rect 631 374 635 378
rect 671 374 675 378
rect 687 374 691 378
rect 727 374 731 378
rect 751 374 755 378
rect 791 374 795 378
rect 855 374 859 378
rect 1095 374 1099 378
rect 1135 374 1139 378
rect 1159 374 1163 378
rect 1199 374 1203 378
rect 1255 374 1259 378
rect 1303 374 1307 378
rect 1335 374 1339 378
rect 1343 374 1347 378
rect 1383 374 1387 378
rect 1415 374 1419 378
rect 1423 374 1427 378
rect 1463 374 1467 378
rect 1503 374 1507 378
rect 1551 374 1555 378
rect 1591 374 1595 378
rect 1615 374 1619 378
rect 1671 374 1675 378
rect 1679 374 1683 378
rect 1751 374 1755 378
rect 463 318 467 322
rect 471 318 475 322
rect 519 318 523 322
rect 551 318 555 322
rect 575 318 579 322
rect 623 318 627 322
rect 631 318 635 322
rect 687 318 691 322
rect 751 318 755 322
rect 807 318 811 322
rect 871 318 875 322
rect 935 318 939 322
rect 1095 318 1099 322
rect 1135 318 1139 322
rect 1167 318 1171 322
rect 1207 318 1211 322
rect 1247 318 1251 322
rect 1295 318 1299 322
rect 1303 318 1307 322
rect 1343 318 1347 322
rect 1383 318 1387 322
rect 1391 318 1395 322
rect 1423 318 1427 322
rect 1439 318 1443 322
rect 1463 318 1467 322
rect 1495 318 1499 322
rect 1503 318 1507 322
rect 111 266 115 270
rect 135 266 139 270
rect 199 266 203 270
rect 207 266 211 270
rect 279 266 283 270
rect 295 266 299 270
rect 359 266 363 270
rect 383 266 387 270
rect 439 266 443 270
rect 471 266 475 270
rect 511 266 515 270
rect 111 210 115 214
rect 135 210 139 214
rect 183 210 187 214
rect 199 210 203 214
rect 231 210 235 214
rect 279 210 283 214
rect 327 210 331 214
rect 551 266 555 270
rect 583 266 587 270
rect 623 266 627 270
rect 647 266 651 270
rect 687 266 691 270
rect 703 266 707 270
rect 751 266 755 270
rect 759 266 763 270
rect 807 266 811 270
rect 815 266 819 270
rect 871 266 875 270
rect 879 266 883 270
rect 359 210 363 214
rect 375 210 379 214
rect 415 210 419 214
rect 439 210 443 214
rect 455 210 459 214
rect 503 210 507 214
rect 511 210 515 214
rect 551 210 555 214
rect 583 210 587 214
rect 935 266 939 270
rect 1095 266 1099 270
rect 1135 258 1139 262
rect 1159 258 1163 262
rect 1167 258 1171 262
rect 1207 258 1211 262
rect 1247 258 1251 262
rect 1271 258 1275 262
rect 1295 258 1299 262
rect 1327 258 1331 262
rect 1343 258 1347 262
rect 1391 258 1395 262
rect 1439 258 1443 262
rect 1455 258 1459 262
rect 1495 258 1499 262
rect 599 210 603 214
rect 647 210 651 214
rect 695 210 699 214
rect 703 210 707 214
rect 743 210 747 214
rect 759 210 763 214
rect 815 210 819 214
rect 879 210 883 214
rect 1095 210 1099 214
rect 1135 206 1139 210
rect 1159 206 1163 210
rect 1199 206 1203 210
rect 1207 206 1211 210
rect 1263 206 1267 210
rect 1271 206 1275 210
rect 111 134 115 138
rect 135 134 139 138
rect 143 134 147 138
rect 183 134 187 138
rect 223 134 227 138
rect 231 134 235 138
rect 263 134 267 138
rect 279 134 283 138
rect 303 134 307 138
rect 327 134 331 138
rect 343 134 347 138
rect 375 134 379 138
rect 383 134 387 138
rect 415 134 419 138
rect 423 134 427 138
rect 455 134 459 138
rect 463 134 467 138
rect 503 134 507 138
rect 543 134 547 138
rect 551 134 555 138
rect 583 134 587 138
rect 599 134 603 138
rect 623 134 627 138
rect 647 134 651 138
rect 663 134 667 138
rect 695 134 699 138
rect 703 134 707 138
rect 743 134 747 138
rect 783 134 787 138
rect 831 134 835 138
rect 879 134 883 138
rect 927 134 931 138
rect 967 134 971 138
rect 1007 134 1011 138
rect 1047 134 1051 138
rect 1095 134 1099 138
rect 1135 134 1139 138
rect 1159 134 1163 138
rect 1327 206 1331 210
rect 1391 206 1395 210
rect 1399 206 1403 210
rect 1551 318 1555 322
rect 1559 318 1563 322
rect 1823 374 1827 378
rect 1831 374 1835 378
rect 1887 374 1891 378
rect 1919 374 1923 378
rect 1951 374 1955 378
rect 1615 318 1619 322
rect 1623 318 1627 322
rect 1679 318 1683 322
rect 1695 318 1699 322
rect 1751 318 1755 322
rect 1775 318 1779 322
rect 1831 318 1835 322
rect 1855 318 1859 322
rect 1919 318 1923 322
rect 1935 318 1939 322
rect 2071 430 2075 434
rect 2119 430 2123 434
rect 2007 374 2011 378
rect 2023 374 2027 378
rect 2071 374 2075 378
rect 2119 374 2123 378
rect 2007 318 2011 322
rect 2015 318 2019 322
rect 2071 318 2075 322
rect 1527 258 1531 262
rect 1559 258 1563 262
rect 1607 258 1611 262
rect 1623 258 1627 262
rect 1687 258 1691 262
rect 1695 258 1699 262
rect 1767 258 1771 262
rect 1775 258 1779 262
rect 1839 258 1843 262
rect 1855 258 1859 262
rect 1919 258 1923 262
rect 1935 258 1939 262
rect 1999 258 2003 262
rect 1455 206 1459 210
rect 1471 206 1475 210
rect 1199 134 1203 138
rect 1207 134 1211 138
rect 1263 134 1267 138
rect 1271 134 1275 138
rect 1527 206 1531 210
rect 1543 206 1547 210
rect 1607 206 1611 210
rect 1671 206 1675 210
rect 1687 206 1691 210
rect 1735 206 1739 210
rect 1327 134 1331 138
rect 1335 134 1339 138
rect 1399 134 1403 138
rect 1455 134 1459 138
rect 1471 134 1475 138
rect 1511 134 1515 138
rect 1543 134 1547 138
rect 1559 134 1563 138
rect 1767 206 1771 210
rect 1807 206 1811 210
rect 1839 206 1843 210
rect 1879 206 1883 210
rect 1919 206 1923 210
rect 1951 206 1955 210
rect 2119 318 2123 322
rect 2015 258 2019 262
rect 2071 258 2075 262
rect 2119 258 2123 262
rect 1999 206 2003 210
rect 2023 206 2027 210
rect 2071 206 2075 210
rect 1607 134 1611 138
rect 1647 134 1651 138
rect 1671 134 1675 138
rect 1687 134 1691 138
rect 1727 134 1731 138
rect 1735 134 1739 138
rect 1767 134 1771 138
rect 1807 134 1811 138
rect 1855 134 1859 138
rect 1879 134 1883 138
rect 1903 134 1907 138
rect 1951 134 1955 138
rect 1991 134 1995 138
rect 2023 134 2027 138
rect 2031 134 2035 138
rect 2071 134 2075 138
rect 2119 206 2123 210
rect 2119 134 2123 138
rect 111 82 115 86
rect 143 82 147 86
rect 183 82 187 86
rect 223 82 227 86
rect 263 82 267 86
rect 303 82 307 86
rect 343 82 347 86
rect 383 82 387 86
rect 423 82 427 86
rect 463 82 467 86
rect 503 82 507 86
rect 543 82 547 86
rect 583 82 587 86
rect 623 82 627 86
rect 663 82 667 86
rect 703 82 707 86
rect 743 82 747 86
rect 783 82 787 86
rect 831 82 835 86
rect 879 82 883 86
rect 927 82 931 86
rect 967 82 971 86
rect 1007 82 1011 86
rect 1047 82 1051 86
rect 1095 82 1099 86
rect 1135 82 1139 86
rect 1159 82 1163 86
rect 1207 82 1211 86
rect 1271 82 1275 86
rect 1335 82 1339 86
rect 1399 82 1403 86
rect 1455 82 1459 86
rect 1511 82 1515 86
rect 1559 82 1563 86
rect 1607 82 1611 86
rect 1647 82 1651 86
rect 1687 82 1691 86
rect 1727 82 1731 86
rect 1767 82 1771 86
rect 1807 82 1811 86
rect 1855 82 1859 86
rect 1903 82 1907 86
rect 1951 82 1955 86
rect 1991 82 1995 86
rect 2031 82 2035 86
rect 2071 82 2075 86
rect 2119 82 2123 86
<< m4 >>
rect 1118 2225 1119 2231
rect 1125 2230 2155 2231
rect 1125 2226 1135 2230
rect 1139 2226 1687 2230
rect 1691 2226 1727 2230
rect 1731 2226 1767 2230
rect 1771 2226 1807 2230
rect 1811 2226 2119 2230
rect 2123 2226 2155 2230
rect 1125 2225 2155 2226
rect 2161 2225 2162 2231
rect 84 2209 85 2215
rect 91 2214 1107 2215
rect 91 2210 111 2214
rect 115 2210 135 2214
rect 139 2210 175 2214
rect 179 2210 215 2214
rect 219 2210 255 2214
rect 259 2210 319 2214
rect 323 2210 383 2214
rect 387 2210 447 2214
rect 451 2210 511 2214
rect 515 2210 575 2214
rect 579 2210 631 2214
rect 635 2210 687 2214
rect 691 2210 735 2214
rect 739 2210 791 2214
rect 795 2210 847 2214
rect 851 2210 903 2214
rect 907 2210 1095 2214
rect 1099 2210 1107 2214
rect 91 2209 1107 2210
rect 1113 2209 1114 2215
rect 1106 2173 1107 2179
rect 1113 2178 2143 2179
rect 1113 2174 1135 2178
rect 1139 2174 1159 2178
rect 1163 2174 1199 2178
rect 1203 2174 1239 2178
rect 1243 2174 1279 2178
rect 1283 2174 1335 2178
rect 1339 2174 1391 2178
rect 1395 2174 1455 2178
rect 1459 2174 1527 2178
rect 1531 2174 1591 2178
rect 1595 2174 1663 2178
rect 1667 2174 1687 2178
rect 1691 2174 1727 2178
rect 1731 2174 1735 2178
rect 1739 2174 1767 2178
rect 1771 2174 1807 2178
rect 1811 2174 1879 2178
rect 1883 2174 2119 2178
rect 2123 2174 2143 2178
rect 1113 2173 2143 2174
rect 2149 2173 2150 2179
rect 96 2149 97 2155
rect 103 2154 1119 2155
rect 103 2150 111 2154
rect 115 2150 135 2154
rect 139 2150 175 2154
rect 179 2150 215 2154
rect 219 2150 231 2154
rect 235 2150 255 2154
rect 259 2150 271 2154
rect 275 2150 311 2154
rect 315 2150 319 2154
rect 323 2150 359 2154
rect 363 2150 383 2154
rect 387 2150 423 2154
rect 427 2150 447 2154
rect 451 2150 487 2154
rect 491 2150 511 2154
rect 515 2150 559 2154
rect 563 2150 575 2154
rect 579 2150 631 2154
rect 635 2150 639 2154
rect 643 2150 687 2154
rect 691 2150 719 2154
rect 723 2150 735 2154
rect 739 2150 791 2154
rect 795 2150 799 2154
rect 803 2150 847 2154
rect 851 2150 879 2154
rect 883 2150 903 2154
rect 907 2150 967 2154
rect 971 2150 1095 2154
rect 1099 2150 1119 2154
rect 103 2149 1119 2150
rect 1125 2149 1126 2155
rect 1118 2121 1119 2127
rect 1125 2126 2155 2127
rect 1125 2122 1135 2126
rect 1139 2122 1159 2126
rect 1163 2122 1199 2126
rect 1203 2122 1239 2126
rect 1243 2122 1279 2126
rect 1283 2122 1295 2126
rect 1299 2122 1335 2126
rect 1339 2122 1367 2126
rect 1371 2122 1391 2126
rect 1395 2122 1439 2126
rect 1443 2122 1455 2126
rect 1459 2122 1519 2126
rect 1523 2122 1527 2126
rect 1531 2122 1591 2126
rect 1595 2122 1599 2126
rect 1603 2122 1663 2126
rect 1667 2122 1679 2126
rect 1683 2122 1735 2126
rect 1739 2122 1751 2126
rect 1755 2122 1807 2126
rect 1811 2122 1823 2126
rect 1827 2122 1879 2126
rect 1883 2122 1887 2126
rect 1891 2122 1951 2126
rect 1955 2122 2023 2126
rect 2027 2122 2071 2126
rect 2075 2122 2119 2126
rect 2123 2122 2155 2126
rect 1125 2121 2155 2122
rect 2161 2121 2162 2127
rect 84 2093 85 2099
rect 91 2098 1107 2099
rect 91 2094 111 2098
rect 115 2094 231 2098
rect 235 2094 271 2098
rect 275 2094 303 2098
rect 307 2094 311 2098
rect 315 2094 351 2098
rect 355 2094 359 2098
rect 363 2094 407 2098
rect 411 2094 423 2098
rect 427 2094 471 2098
rect 475 2094 487 2098
rect 491 2094 543 2098
rect 547 2094 559 2098
rect 563 2094 623 2098
rect 627 2094 639 2098
rect 643 2094 703 2098
rect 707 2094 719 2098
rect 723 2094 783 2098
rect 787 2094 799 2098
rect 803 2094 863 2098
rect 867 2094 879 2098
rect 883 2094 951 2098
rect 955 2094 967 2098
rect 971 2094 1039 2098
rect 1043 2094 1095 2098
rect 1099 2094 1107 2098
rect 91 2093 1107 2094
rect 1113 2093 1114 2099
rect 1106 2069 1107 2075
rect 1113 2074 2143 2075
rect 1113 2070 1135 2074
rect 1139 2070 1159 2074
rect 1163 2070 1199 2074
rect 1203 2070 1215 2074
rect 1219 2070 1239 2074
rect 1243 2070 1295 2074
rect 1299 2070 1303 2074
rect 1307 2070 1367 2074
rect 1371 2070 1399 2074
rect 1403 2070 1439 2074
rect 1443 2070 1495 2074
rect 1499 2070 1519 2074
rect 1523 2070 1591 2074
rect 1595 2070 1599 2074
rect 1603 2070 1679 2074
rect 1683 2070 1751 2074
rect 1755 2070 1759 2074
rect 1763 2070 1823 2074
rect 1827 2070 1831 2074
rect 1835 2070 1887 2074
rect 1891 2070 1895 2074
rect 1899 2070 1951 2074
rect 1955 2070 1959 2074
rect 1963 2070 2023 2074
rect 2027 2070 2071 2074
rect 2075 2070 2119 2074
rect 2123 2070 2143 2074
rect 1113 2069 2143 2070
rect 2149 2069 2150 2075
rect 96 2037 97 2043
rect 103 2042 1119 2043
rect 103 2038 111 2042
rect 115 2038 183 2042
rect 187 2038 279 2042
rect 283 2038 303 2042
rect 307 2038 351 2042
rect 355 2038 375 2042
rect 379 2038 407 2042
rect 411 2038 463 2042
rect 467 2038 471 2042
rect 475 2038 543 2042
rect 547 2038 623 2042
rect 627 2038 695 2042
rect 699 2038 703 2042
rect 707 2038 759 2042
rect 763 2038 783 2042
rect 787 2038 815 2042
rect 819 2038 863 2042
rect 867 2038 911 2042
rect 915 2038 951 2042
rect 955 2038 959 2042
rect 963 2038 1007 2042
rect 1011 2038 1039 2042
rect 1043 2038 1047 2042
rect 1051 2038 1095 2042
rect 1099 2038 1119 2042
rect 103 2037 1119 2038
rect 1125 2037 1126 2043
rect 1118 2017 1119 2023
rect 1125 2022 2155 2023
rect 1125 2018 1135 2022
rect 1139 2018 1159 2022
rect 1163 2018 1215 2022
rect 1219 2018 1239 2022
rect 1243 2018 1303 2022
rect 1307 2018 1351 2022
rect 1355 2018 1399 2022
rect 1403 2018 1455 2022
rect 1459 2018 1495 2022
rect 1499 2018 1559 2022
rect 1563 2018 1591 2022
rect 1595 2018 1655 2022
rect 1659 2018 1679 2022
rect 1683 2018 1743 2022
rect 1747 2018 1759 2022
rect 1763 2018 1823 2022
rect 1827 2018 1831 2022
rect 1835 2018 1895 2022
rect 1899 2018 1959 2022
rect 1963 2018 2023 2022
rect 2027 2018 2071 2022
rect 2075 2018 2119 2022
rect 2123 2018 2155 2022
rect 1125 2017 2155 2018
rect 2161 2017 2162 2023
rect 84 1985 85 1991
rect 91 1990 1107 1991
rect 91 1986 111 1990
rect 115 1986 159 1990
rect 163 1986 183 1990
rect 187 1986 231 1990
rect 235 1986 279 1990
rect 283 1986 303 1990
rect 307 1986 375 1990
rect 379 1986 447 1990
rect 451 1986 463 1990
rect 467 1986 527 1990
rect 531 1986 543 1990
rect 547 1986 607 1990
rect 611 1986 623 1990
rect 627 1986 687 1990
rect 691 1986 695 1990
rect 699 1986 759 1990
rect 763 1986 815 1990
rect 819 1986 831 1990
rect 835 1986 863 1990
rect 867 1986 911 1990
rect 915 1986 959 1990
rect 963 1986 991 1990
rect 995 1986 1007 1990
rect 1011 1986 1047 1990
rect 1051 1986 1095 1990
rect 1099 1986 1107 1990
rect 91 1985 1107 1986
rect 1113 1985 1114 1991
rect 1106 1953 1107 1959
rect 1113 1958 2143 1959
rect 1113 1954 1135 1958
rect 1139 1954 1159 1958
rect 1163 1954 1239 1958
rect 1243 1954 1351 1958
rect 1355 1954 1359 1958
rect 1363 1954 1423 1958
rect 1427 1954 1455 1958
rect 1459 1954 1487 1958
rect 1491 1954 1559 1958
rect 1563 1954 1631 1958
rect 1635 1954 1655 1958
rect 1659 1954 1703 1958
rect 1707 1954 1743 1958
rect 1747 1954 1775 1958
rect 1779 1954 1823 1958
rect 1827 1954 1847 1958
rect 1851 1954 1895 1958
rect 1899 1954 1927 1958
rect 1931 1954 1959 1958
rect 1963 1954 2007 1958
rect 2011 1954 2023 1958
rect 2027 1954 2071 1958
rect 2075 1954 2119 1958
rect 2123 1954 2143 1958
rect 1113 1953 2143 1954
rect 2149 1953 2150 1959
rect 96 1929 97 1935
rect 103 1934 1119 1935
rect 103 1930 111 1934
rect 115 1930 135 1934
rect 139 1930 159 1934
rect 163 1930 175 1934
rect 179 1930 231 1934
rect 235 1930 295 1934
rect 299 1930 303 1934
rect 307 1930 367 1934
rect 371 1930 375 1934
rect 379 1930 447 1934
rect 451 1930 527 1934
rect 531 1930 607 1934
rect 611 1930 615 1934
rect 619 1930 687 1934
rect 691 1930 703 1934
rect 707 1930 759 1934
rect 763 1930 791 1934
rect 795 1930 831 1934
rect 835 1930 879 1934
rect 883 1930 911 1934
rect 915 1930 991 1934
rect 995 1930 1095 1934
rect 1099 1930 1119 1934
rect 103 1929 1119 1930
rect 1125 1929 1126 1935
rect 1118 1901 1119 1907
rect 1125 1906 2155 1907
rect 1125 1902 1135 1906
rect 1139 1902 1231 1906
rect 1235 1902 1271 1906
rect 1275 1902 1319 1906
rect 1323 1902 1359 1906
rect 1363 1902 1375 1906
rect 1379 1902 1423 1906
rect 1427 1902 1439 1906
rect 1443 1902 1487 1906
rect 1491 1902 1503 1906
rect 1507 1902 1559 1906
rect 1563 1902 1575 1906
rect 1579 1902 1631 1906
rect 1635 1902 1655 1906
rect 1659 1902 1703 1906
rect 1707 1902 1751 1906
rect 1755 1902 1775 1906
rect 1779 1902 1847 1906
rect 1851 1902 1863 1906
rect 1867 1902 1927 1906
rect 1931 1902 1975 1906
rect 1979 1902 2007 1906
rect 2011 1902 2071 1906
rect 2075 1902 2119 1906
rect 2123 1902 2155 1906
rect 1125 1901 2155 1902
rect 2161 1901 2162 1907
rect 84 1873 85 1879
rect 91 1878 1107 1879
rect 91 1874 111 1878
rect 115 1874 135 1878
rect 139 1874 175 1878
rect 179 1874 223 1878
rect 227 1874 231 1878
rect 235 1874 287 1878
rect 291 1874 295 1878
rect 299 1874 359 1878
rect 363 1874 367 1878
rect 371 1874 431 1878
rect 435 1874 447 1878
rect 451 1874 503 1878
rect 507 1874 527 1878
rect 531 1874 567 1878
rect 571 1874 615 1878
rect 619 1874 631 1878
rect 635 1874 695 1878
rect 699 1874 703 1878
rect 707 1874 759 1878
rect 763 1874 791 1878
rect 795 1874 831 1878
rect 835 1874 879 1878
rect 883 1874 1095 1878
rect 1099 1874 1107 1878
rect 91 1873 1107 1874
rect 1113 1873 1114 1879
rect 1106 1845 1107 1851
rect 1113 1850 2143 1851
rect 1113 1846 1135 1850
rect 1139 1846 1159 1850
rect 1163 1846 1199 1850
rect 1203 1846 1231 1850
rect 1235 1846 1239 1850
rect 1243 1846 1271 1850
rect 1275 1846 1303 1850
rect 1307 1846 1319 1850
rect 1323 1846 1367 1850
rect 1371 1846 1375 1850
rect 1379 1846 1431 1850
rect 1435 1846 1439 1850
rect 1443 1846 1503 1850
rect 1507 1846 1575 1850
rect 1579 1846 1583 1850
rect 1587 1846 1655 1850
rect 1659 1846 1671 1850
rect 1675 1846 1751 1850
rect 1755 1846 1767 1850
rect 1771 1846 1863 1850
rect 1867 1846 1871 1850
rect 1875 1846 1975 1850
rect 1979 1846 1983 1850
rect 1987 1846 2071 1850
rect 2075 1846 2119 1850
rect 2123 1846 2143 1850
rect 1113 1845 2143 1846
rect 2149 1845 2150 1851
rect 96 1817 97 1823
rect 103 1822 1119 1823
rect 103 1818 111 1822
rect 115 1818 135 1822
rect 139 1818 175 1822
rect 179 1818 183 1822
rect 187 1818 223 1822
rect 227 1818 263 1822
rect 267 1818 287 1822
rect 291 1818 351 1822
rect 355 1818 359 1822
rect 363 1818 431 1822
rect 435 1818 439 1822
rect 443 1818 503 1822
rect 507 1818 527 1822
rect 531 1818 567 1822
rect 571 1818 607 1822
rect 611 1818 631 1822
rect 635 1818 687 1822
rect 691 1818 695 1822
rect 699 1818 759 1822
rect 763 1818 767 1822
rect 771 1818 831 1822
rect 835 1818 839 1822
rect 843 1818 911 1822
rect 915 1818 991 1822
rect 995 1818 1047 1822
rect 1051 1818 1095 1822
rect 1099 1818 1119 1822
rect 103 1817 1119 1818
rect 1125 1817 1126 1823
rect 1438 1812 1444 1813
rect 2006 1812 2012 1813
rect 1438 1808 1439 1812
rect 1443 1808 2007 1812
rect 2011 1808 2012 1812
rect 1438 1807 1444 1808
rect 2006 1807 2012 1808
rect 1118 1785 1119 1791
rect 1125 1790 2155 1791
rect 1125 1786 1135 1790
rect 1139 1786 1159 1790
rect 1163 1786 1199 1790
rect 1203 1786 1239 1790
rect 1243 1786 1303 1790
rect 1307 1786 1311 1790
rect 1315 1786 1351 1790
rect 1355 1786 1367 1790
rect 1371 1786 1391 1790
rect 1395 1786 1431 1790
rect 1435 1786 1471 1790
rect 1475 1786 1503 1790
rect 1507 1786 1511 1790
rect 1515 1786 1551 1790
rect 1555 1786 1583 1790
rect 1587 1786 1607 1790
rect 1611 1786 1671 1790
rect 1675 1786 1679 1790
rect 1683 1786 1767 1790
rect 1771 1786 1871 1790
rect 1875 1786 1983 1790
rect 1987 1786 2071 1790
rect 2075 1786 2119 1790
rect 2123 1786 2155 1790
rect 1125 1785 2155 1786
rect 2161 1785 2162 1791
rect 84 1757 85 1763
rect 91 1762 1107 1763
rect 91 1758 111 1762
rect 115 1758 135 1762
rect 139 1758 183 1762
rect 187 1758 199 1762
rect 203 1758 263 1762
rect 267 1758 295 1762
rect 299 1758 351 1762
rect 355 1758 399 1762
rect 403 1758 439 1762
rect 443 1758 495 1762
rect 499 1758 527 1762
rect 531 1758 591 1762
rect 595 1758 607 1762
rect 611 1758 671 1762
rect 675 1758 687 1762
rect 691 1758 751 1762
rect 755 1758 767 1762
rect 771 1758 823 1762
rect 827 1758 839 1762
rect 843 1758 887 1762
rect 891 1758 911 1762
rect 915 1758 959 1762
rect 963 1758 991 1762
rect 995 1758 1031 1762
rect 1035 1758 1047 1762
rect 1051 1758 1095 1762
rect 1099 1758 1107 1762
rect 91 1757 1107 1758
rect 1113 1757 1114 1763
rect 1106 1729 1107 1735
rect 1113 1734 2143 1735
rect 1113 1730 1135 1734
rect 1139 1730 1263 1734
rect 1267 1730 1311 1734
rect 1315 1730 1319 1734
rect 1323 1730 1351 1734
rect 1355 1730 1383 1734
rect 1387 1730 1391 1734
rect 1395 1730 1431 1734
rect 1435 1730 1455 1734
rect 1459 1730 1471 1734
rect 1475 1730 1511 1734
rect 1515 1730 1535 1734
rect 1539 1730 1551 1734
rect 1555 1730 1607 1734
rect 1611 1730 1615 1734
rect 1619 1730 1679 1734
rect 1683 1730 1687 1734
rect 1691 1730 1759 1734
rect 1763 1730 1767 1734
rect 1771 1730 1831 1734
rect 1835 1730 1871 1734
rect 1875 1730 1895 1734
rect 1899 1730 1959 1734
rect 1963 1730 1983 1734
rect 1987 1730 2023 1734
rect 2027 1730 2071 1734
rect 2075 1730 2119 1734
rect 2123 1730 2143 1734
rect 1113 1729 2143 1730
rect 2149 1729 2150 1735
rect 96 1701 97 1707
rect 103 1706 1119 1707
rect 103 1702 111 1706
rect 115 1702 135 1706
rect 139 1702 151 1706
rect 155 1702 199 1706
rect 203 1702 223 1706
rect 227 1702 295 1706
rect 299 1702 303 1706
rect 307 1702 383 1706
rect 387 1702 399 1706
rect 403 1702 463 1706
rect 467 1702 495 1706
rect 499 1702 535 1706
rect 539 1702 591 1706
rect 595 1702 607 1706
rect 611 1702 671 1706
rect 675 1702 735 1706
rect 739 1702 751 1706
rect 755 1702 807 1706
rect 811 1702 823 1706
rect 827 1702 879 1706
rect 883 1702 887 1706
rect 891 1702 959 1706
rect 963 1702 1031 1706
rect 1035 1702 1095 1706
rect 1099 1702 1119 1706
rect 103 1701 1119 1702
rect 1125 1701 1126 1707
rect 1118 1677 1119 1683
rect 1125 1682 2155 1683
rect 1125 1678 1135 1682
rect 1139 1678 1167 1682
rect 1171 1678 1247 1682
rect 1251 1678 1263 1682
rect 1267 1678 1319 1682
rect 1323 1678 1335 1682
rect 1339 1678 1383 1682
rect 1387 1678 1423 1682
rect 1427 1678 1455 1682
rect 1459 1678 1511 1682
rect 1515 1678 1535 1682
rect 1539 1678 1599 1682
rect 1603 1678 1615 1682
rect 1619 1678 1679 1682
rect 1683 1678 1687 1682
rect 1691 1678 1751 1682
rect 1755 1678 1759 1682
rect 1763 1678 1815 1682
rect 1819 1678 1831 1682
rect 1835 1678 1871 1682
rect 1875 1678 1895 1682
rect 1899 1678 1927 1682
rect 1931 1678 1959 1682
rect 1963 1678 1983 1682
rect 1987 1678 2023 1682
rect 2027 1678 2031 1682
rect 2035 1678 2071 1682
rect 2075 1678 2119 1682
rect 2123 1678 2155 1682
rect 1125 1677 2155 1678
rect 2161 1677 2162 1683
rect 84 1645 85 1651
rect 91 1650 1107 1651
rect 91 1646 111 1650
rect 115 1646 151 1650
rect 155 1646 175 1650
rect 179 1646 215 1650
rect 219 1646 223 1650
rect 227 1646 255 1650
rect 259 1646 303 1650
rect 307 1646 359 1650
rect 363 1646 383 1650
rect 387 1646 407 1650
rect 411 1646 455 1650
rect 459 1646 463 1650
rect 467 1646 503 1650
rect 507 1646 535 1650
rect 539 1646 551 1650
rect 555 1646 607 1650
rect 611 1646 663 1650
rect 667 1646 671 1650
rect 675 1646 719 1650
rect 723 1646 735 1650
rect 739 1646 807 1650
rect 811 1646 879 1650
rect 883 1646 1095 1650
rect 1099 1646 1107 1650
rect 91 1645 1107 1646
rect 1113 1645 1114 1651
rect 1106 1621 1107 1627
rect 1113 1626 2143 1627
rect 1113 1622 1135 1626
rect 1139 1622 1159 1626
rect 1163 1622 1167 1626
rect 1171 1622 1199 1626
rect 1203 1622 1247 1626
rect 1251 1622 1319 1626
rect 1323 1622 1335 1626
rect 1339 1622 1391 1626
rect 1395 1622 1423 1626
rect 1427 1622 1463 1626
rect 1467 1622 1511 1626
rect 1515 1622 1535 1626
rect 1539 1622 1599 1626
rect 1603 1622 1607 1626
rect 1611 1622 1679 1626
rect 1683 1622 1751 1626
rect 1755 1622 1815 1626
rect 1819 1622 1831 1626
rect 1835 1622 1871 1626
rect 1875 1622 1927 1626
rect 1931 1622 1983 1626
rect 1987 1622 2031 1626
rect 2035 1622 2071 1626
rect 2075 1622 2119 1626
rect 2123 1622 2143 1626
rect 1113 1621 2143 1622
rect 2149 1621 2150 1627
rect 96 1585 97 1591
rect 103 1590 1119 1591
rect 103 1586 111 1590
rect 115 1586 143 1590
rect 147 1586 175 1590
rect 179 1586 183 1590
rect 187 1586 215 1590
rect 219 1586 231 1590
rect 235 1586 255 1590
rect 259 1586 287 1590
rect 291 1586 303 1590
rect 307 1586 351 1590
rect 355 1586 359 1590
rect 363 1586 407 1590
rect 411 1586 415 1590
rect 419 1586 455 1590
rect 459 1586 479 1590
rect 483 1586 503 1590
rect 507 1586 543 1590
rect 547 1586 551 1590
rect 555 1586 607 1590
rect 611 1586 663 1590
rect 667 1586 719 1590
rect 723 1586 727 1590
rect 731 1586 791 1590
rect 795 1586 855 1590
rect 859 1586 1095 1590
rect 1099 1586 1119 1590
rect 103 1585 1119 1586
rect 1125 1585 1126 1591
rect 1118 1569 1119 1575
rect 1125 1574 2155 1575
rect 1125 1570 1135 1574
rect 1139 1570 1159 1574
rect 1163 1570 1199 1574
rect 1203 1570 1239 1574
rect 1243 1570 1247 1574
rect 1251 1570 1279 1574
rect 1283 1570 1319 1574
rect 1323 1570 1327 1574
rect 1331 1570 1375 1574
rect 1379 1570 1391 1574
rect 1395 1570 1423 1574
rect 1427 1570 1463 1574
rect 1467 1570 1471 1574
rect 1475 1570 1519 1574
rect 1523 1570 1535 1574
rect 1539 1570 1567 1574
rect 1571 1570 1607 1574
rect 1611 1570 1623 1574
rect 1627 1570 1679 1574
rect 1683 1570 1735 1574
rect 1739 1570 1751 1574
rect 1755 1570 1831 1574
rect 1835 1570 2119 1574
rect 2123 1570 2155 1574
rect 1125 1569 2155 1570
rect 2161 1569 2162 1575
rect 1258 1548 1264 1549
rect 1398 1548 1404 1549
rect 1258 1544 1259 1548
rect 1263 1544 1399 1548
rect 1403 1544 1404 1548
rect 1258 1543 1264 1544
rect 1398 1543 1404 1544
rect 84 1525 85 1531
rect 91 1530 1107 1531
rect 91 1526 111 1530
rect 115 1526 135 1530
rect 139 1526 143 1530
rect 147 1526 175 1530
rect 179 1526 183 1530
rect 187 1526 215 1530
rect 219 1526 231 1530
rect 235 1526 255 1530
rect 259 1526 287 1530
rect 291 1526 295 1530
rect 299 1526 335 1530
rect 339 1526 351 1530
rect 355 1526 375 1530
rect 379 1526 415 1530
rect 419 1526 455 1530
rect 459 1526 479 1530
rect 483 1526 495 1530
rect 499 1526 535 1530
rect 539 1526 543 1530
rect 547 1526 575 1530
rect 579 1526 607 1530
rect 611 1526 615 1530
rect 619 1526 655 1530
rect 659 1526 663 1530
rect 667 1526 695 1530
rect 699 1526 727 1530
rect 731 1526 735 1530
rect 739 1526 775 1530
rect 779 1526 791 1530
rect 795 1526 831 1530
rect 835 1526 855 1530
rect 859 1526 887 1530
rect 891 1526 1095 1530
rect 1099 1526 1107 1530
rect 91 1525 1107 1526
rect 1113 1525 1114 1531
rect 1106 1513 1107 1519
rect 1113 1518 2143 1519
rect 1113 1514 1135 1518
rect 1139 1514 1239 1518
rect 1243 1514 1279 1518
rect 1283 1514 1319 1518
rect 1323 1514 1327 1518
rect 1331 1514 1359 1518
rect 1363 1514 1375 1518
rect 1379 1514 1399 1518
rect 1403 1514 1423 1518
rect 1427 1514 1439 1518
rect 1443 1514 1471 1518
rect 1475 1514 1479 1518
rect 1483 1514 1519 1518
rect 1523 1514 1559 1518
rect 1563 1514 1567 1518
rect 1571 1514 1607 1518
rect 1611 1514 1623 1518
rect 1627 1514 1663 1518
rect 1667 1514 1679 1518
rect 1683 1514 1735 1518
rect 1739 1514 1815 1518
rect 1819 1514 1903 1518
rect 1907 1514 1991 1518
rect 1995 1514 2071 1518
rect 2075 1514 2119 1518
rect 2123 1514 2143 1518
rect 1113 1513 2143 1514
rect 2149 1513 2150 1519
rect 1590 1476 1596 1477
rect 1910 1476 1916 1477
rect 1590 1472 1591 1476
rect 1595 1472 1911 1476
rect 1915 1472 1916 1476
rect 1590 1471 1596 1472
rect 1910 1471 1916 1472
rect 96 1465 97 1471
rect 103 1470 1119 1471
rect 103 1466 111 1470
rect 115 1466 135 1470
rect 139 1466 175 1470
rect 179 1466 215 1470
rect 219 1466 255 1470
rect 259 1466 295 1470
rect 299 1466 335 1470
rect 339 1466 375 1470
rect 379 1466 415 1470
rect 419 1466 455 1470
rect 459 1466 495 1470
rect 499 1466 519 1470
rect 523 1466 535 1470
rect 539 1466 559 1470
rect 563 1466 575 1470
rect 579 1466 599 1470
rect 603 1466 615 1470
rect 619 1466 647 1470
rect 651 1466 655 1470
rect 659 1466 695 1470
rect 699 1466 735 1470
rect 739 1466 751 1470
rect 755 1466 775 1470
rect 779 1466 807 1470
rect 811 1466 831 1470
rect 835 1466 871 1470
rect 875 1466 887 1470
rect 891 1466 935 1470
rect 939 1466 1095 1470
rect 1099 1466 1119 1470
rect 103 1465 1119 1466
rect 1125 1467 1126 1471
rect 1125 1466 2162 1467
rect 1125 1465 1135 1466
rect 1118 1462 1135 1465
rect 1139 1462 1231 1466
rect 1235 1462 1279 1466
rect 1283 1462 1319 1466
rect 1323 1462 1335 1466
rect 1339 1462 1359 1466
rect 1363 1462 1391 1466
rect 1395 1462 1399 1466
rect 1403 1462 1439 1466
rect 1443 1462 1455 1466
rect 1459 1462 1479 1466
rect 1483 1462 1519 1466
rect 1523 1462 1559 1466
rect 1563 1462 1583 1466
rect 1587 1462 1607 1466
rect 1611 1462 1647 1466
rect 1651 1462 1663 1466
rect 1667 1462 1719 1466
rect 1723 1462 1735 1466
rect 1739 1462 1807 1466
rect 1811 1462 1815 1466
rect 1819 1462 1895 1466
rect 1899 1462 1903 1466
rect 1907 1462 1991 1466
rect 1995 1462 2071 1466
rect 2075 1462 2119 1466
rect 2123 1462 2162 1466
rect 1118 1461 2162 1462
rect 1326 1444 1332 1445
rect 1542 1444 1548 1445
rect 1326 1440 1327 1444
rect 1331 1440 1543 1444
rect 1547 1440 1548 1444
rect 1326 1439 1332 1440
rect 1542 1439 1548 1440
rect 84 1409 85 1415
rect 91 1414 1107 1415
rect 91 1410 111 1414
rect 115 1410 431 1414
rect 435 1410 471 1414
rect 475 1410 519 1414
rect 523 1410 559 1414
rect 563 1410 575 1414
rect 579 1410 599 1414
rect 603 1410 631 1414
rect 635 1410 647 1414
rect 651 1410 695 1414
rect 699 1410 751 1414
rect 755 1410 759 1414
rect 763 1410 807 1414
rect 811 1410 823 1414
rect 827 1410 871 1414
rect 875 1410 895 1414
rect 899 1410 935 1414
rect 939 1410 967 1414
rect 971 1410 1095 1414
rect 1099 1410 1107 1414
rect 91 1409 1107 1410
rect 1113 1411 1114 1415
rect 1113 1410 2150 1411
rect 1113 1409 1135 1410
rect 1106 1406 1135 1409
rect 1139 1406 1159 1410
rect 1163 1406 1199 1410
rect 1203 1406 1231 1410
rect 1235 1406 1263 1410
rect 1267 1406 1279 1410
rect 1283 1406 1335 1410
rect 1339 1406 1351 1410
rect 1355 1406 1391 1410
rect 1395 1406 1447 1410
rect 1451 1406 1455 1410
rect 1459 1406 1519 1410
rect 1523 1406 1543 1410
rect 1547 1406 1583 1410
rect 1587 1406 1631 1410
rect 1635 1406 1647 1410
rect 1651 1406 1719 1410
rect 1723 1406 1799 1410
rect 1803 1406 1807 1410
rect 1811 1406 1871 1410
rect 1875 1406 1895 1410
rect 1899 1406 1943 1410
rect 1947 1406 1991 1410
rect 1995 1406 2015 1410
rect 2019 1406 2071 1410
rect 2075 1406 2119 1410
rect 2123 1406 2150 1410
rect 1106 1405 2150 1406
rect 1670 1372 1676 1373
rect 1930 1372 1936 1373
rect 1670 1368 1671 1372
rect 1675 1368 1931 1372
rect 1935 1368 1936 1372
rect 1670 1367 1676 1368
rect 1930 1367 1936 1368
rect 96 1357 97 1363
rect 103 1362 1119 1363
rect 103 1358 111 1362
rect 115 1358 375 1362
rect 379 1358 423 1362
rect 427 1358 431 1362
rect 435 1358 471 1362
rect 475 1358 479 1362
rect 483 1358 519 1362
rect 523 1358 543 1362
rect 547 1358 575 1362
rect 579 1358 607 1362
rect 611 1358 631 1362
rect 635 1358 671 1362
rect 675 1358 695 1362
rect 699 1358 735 1362
rect 739 1358 759 1362
rect 763 1358 799 1362
rect 803 1358 823 1362
rect 827 1358 863 1362
rect 867 1358 895 1362
rect 899 1358 927 1362
rect 931 1358 967 1362
rect 971 1358 999 1362
rect 1003 1358 1047 1362
rect 1051 1358 1095 1362
rect 1099 1358 1119 1362
rect 103 1357 1119 1358
rect 1125 1357 1126 1363
rect 1118 1355 1126 1357
rect 1118 1349 1119 1355
rect 1125 1354 2155 1355
rect 1125 1350 1135 1354
rect 1139 1350 1159 1354
rect 1163 1350 1199 1354
rect 1203 1350 1255 1354
rect 1259 1350 1263 1354
rect 1267 1350 1351 1354
rect 1355 1350 1375 1354
rect 1379 1350 1447 1354
rect 1451 1350 1487 1354
rect 1491 1350 1543 1354
rect 1547 1350 1591 1354
rect 1595 1350 1631 1354
rect 1635 1350 1679 1354
rect 1683 1350 1719 1354
rect 1723 1350 1759 1354
rect 1763 1350 1799 1354
rect 1803 1350 1831 1354
rect 1835 1350 1871 1354
rect 1875 1350 1903 1354
rect 1907 1350 1943 1354
rect 1947 1350 1967 1354
rect 1971 1350 2015 1354
rect 2019 1350 2031 1354
rect 2035 1350 2071 1354
rect 2075 1350 2119 1354
rect 2123 1350 2155 1354
rect 1125 1349 2155 1350
rect 2161 1349 2162 1355
rect 84 1305 85 1311
rect 91 1310 1107 1311
rect 91 1306 111 1310
rect 115 1306 335 1310
rect 339 1306 375 1310
rect 379 1306 391 1310
rect 395 1306 423 1310
rect 427 1306 455 1310
rect 459 1306 479 1310
rect 483 1306 527 1310
rect 531 1306 543 1310
rect 547 1306 599 1310
rect 603 1306 607 1310
rect 611 1306 671 1310
rect 675 1306 735 1310
rect 739 1306 743 1310
rect 747 1306 799 1310
rect 803 1306 823 1310
rect 827 1306 863 1310
rect 867 1306 903 1310
rect 907 1306 927 1310
rect 931 1306 983 1310
rect 987 1306 999 1310
rect 1003 1306 1047 1310
rect 1051 1306 1095 1310
rect 1099 1306 1107 1310
rect 91 1305 1107 1306
rect 1113 1305 1114 1311
rect 1106 1293 1107 1299
rect 1113 1298 2143 1299
rect 1113 1294 1135 1298
rect 1139 1294 1159 1298
rect 1163 1294 1199 1298
rect 1203 1294 1247 1298
rect 1251 1294 1255 1298
rect 1259 1294 1319 1298
rect 1323 1294 1375 1298
rect 1379 1294 1399 1298
rect 1403 1294 1479 1298
rect 1483 1294 1487 1298
rect 1491 1294 1559 1298
rect 1563 1294 1591 1298
rect 1595 1294 1639 1298
rect 1643 1294 1679 1298
rect 1683 1294 1719 1298
rect 1723 1294 1759 1298
rect 1763 1294 1799 1298
rect 1803 1294 1831 1298
rect 1835 1294 1879 1298
rect 1883 1294 1903 1298
rect 1907 1294 1967 1298
rect 1971 1294 2031 1298
rect 2035 1294 2055 1298
rect 2059 1294 2071 1298
rect 2075 1294 2119 1298
rect 2123 1294 2143 1298
rect 1113 1293 2143 1294
rect 2149 1293 2150 1299
rect 96 1249 97 1255
rect 103 1254 1119 1255
rect 103 1250 111 1254
rect 115 1250 263 1254
rect 267 1250 311 1254
rect 315 1250 335 1254
rect 339 1250 359 1254
rect 363 1250 391 1254
rect 395 1250 415 1254
rect 419 1250 455 1254
rect 459 1250 479 1254
rect 483 1250 527 1254
rect 531 1250 543 1254
rect 547 1250 599 1254
rect 603 1250 607 1254
rect 611 1250 671 1254
rect 675 1250 735 1254
rect 739 1250 743 1254
rect 747 1250 799 1254
rect 803 1250 823 1254
rect 827 1250 863 1254
rect 867 1250 903 1254
rect 907 1250 927 1254
rect 931 1250 983 1254
rect 987 1250 1047 1254
rect 1051 1250 1095 1254
rect 1099 1250 1119 1254
rect 103 1249 1119 1250
rect 1125 1249 1126 1255
rect 1118 1237 1119 1243
rect 1125 1242 2155 1243
rect 1125 1238 1135 1242
rect 1139 1238 1159 1242
rect 1163 1238 1199 1242
rect 1203 1238 1239 1242
rect 1243 1238 1247 1242
rect 1251 1238 1279 1242
rect 1283 1238 1319 1242
rect 1323 1238 1327 1242
rect 1331 1238 1375 1242
rect 1379 1238 1399 1242
rect 1403 1238 1423 1242
rect 1427 1238 1471 1242
rect 1475 1238 1479 1242
rect 1483 1238 1535 1242
rect 1539 1238 1559 1242
rect 1563 1238 1615 1242
rect 1619 1238 1639 1242
rect 1643 1238 1719 1242
rect 1723 1238 1799 1242
rect 1803 1238 1839 1242
rect 1843 1238 1879 1242
rect 1883 1238 1967 1242
rect 1971 1238 2055 1242
rect 2059 1238 2071 1242
rect 2075 1238 2119 1242
rect 2123 1238 2155 1242
rect 1125 1237 2155 1238
rect 2161 1237 2162 1243
rect 84 1197 85 1203
rect 91 1202 1107 1203
rect 91 1198 111 1202
rect 115 1198 223 1202
rect 227 1198 263 1202
rect 267 1198 279 1202
rect 283 1198 311 1202
rect 315 1198 343 1202
rect 347 1198 359 1202
rect 363 1198 407 1202
rect 411 1198 415 1202
rect 419 1198 479 1202
rect 483 1198 543 1202
rect 547 1198 551 1202
rect 555 1198 607 1202
rect 611 1198 631 1202
rect 635 1198 671 1202
rect 675 1198 711 1202
rect 715 1198 735 1202
rect 739 1198 791 1202
rect 795 1198 799 1202
rect 803 1198 863 1202
rect 867 1198 871 1202
rect 875 1198 927 1202
rect 931 1198 959 1202
rect 963 1198 1095 1202
rect 1099 1198 1107 1202
rect 91 1197 1107 1198
rect 1113 1197 1114 1203
rect 1106 1185 1107 1191
rect 1113 1190 2143 1191
rect 1113 1186 1135 1190
rect 1139 1186 1159 1190
rect 1163 1186 1199 1190
rect 1203 1186 1239 1190
rect 1243 1186 1279 1190
rect 1283 1186 1287 1190
rect 1291 1186 1327 1190
rect 1331 1186 1367 1190
rect 1371 1186 1375 1190
rect 1379 1186 1415 1190
rect 1419 1186 1423 1190
rect 1427 1186 1471 1190
rect 1475 1186 1527 1190
rect 1531 1186 1535 1190
rect 1539 1186 1583 1190
rect 1587 1186 1615 1190
rect 1619 1186 1639 1190
rect 1643 1186 1703 1190
rect 1707 1186 1719 1190
rect 1723 1186 1767 1190
rect 1771 1186 1839 1190
rect 1843 1186 1919 1190
rect 1923 1186 1967 1190
rect 1971 1186 2007 1190
rect 2011 1186 2071 1190
rect 2075 1186 2119 1190
rect 2123 1186 2143 1190
rect 1113 1185 2143 1186
rect 2149 1185 2150 1191
rect 96 1145 97 1151
rect 103 1150 1119 1151
rect 103 1146 111 1150
rect 115 1146 159 1150
rect 163 1146 199 1150
rect 203 1146 223 1150
rect 227 1146 247 1150
rect 251 1146 279 1150
rect 283 1146 303 1150
rect 307 1146 343 1150
rect 347 1146 367 1150
rect 371 1146 407 1150
rect 411 1146 439 1150
rect 443 1146 479 1150
rect 483 1146 511 1150
rect 515 1146 551 1150
rect 555 1146 591 1150
rect 595 1146 631 1150
rect 635 1146 679 1150
rect 683 1146 711 1150
rect 715 1146 775 1150
rect 779 1146 791 1150
rect 795 1146 871 1150
rect 875 1146 879 1150
rect 883 1146 959 1150
rect 963 1146 991 1150
rect 995 1146 1095 1150
rect 1099 1146 1119 1150
rect 103 1145 1119 1146
rect 1125 1145 1126 1151
rect 1118 1125 1119 1131
rect 1125 1130 2155 1131
rect 1125 1126 1135 1130
rect 1139 1126 1287 1130
rect 1291 1126 1327 1130
rect 1331 1126 1367 1130
rect 1371 1126 1383 1130
rect 1387 1126 1415 1130
rect 1419 1126 1423 1130
rect 1427 1126 1471 1130
rect 1475 1126 1527 1130
rect 1531 1126 1583 1130
rect 1587 1126 1591 1130
rect 1595 1126 1639 1130
rect 1643 1126 1655 1130
rect 1659 1126 1703 1130
rect 1707 1126 1711 1130
rect 1715 1126 1767 1130
rect 1771 1126 1823 1130
rect 1827 1126 1839 1130
rect 1843 1126 1871 1130
rect 1875 1126 1919 1130
rect 1923 1126 1927 1130
rect 1931 1126 1983 1130
rect 1987 1126 2007 1130
rect 2011 1126 2031 1130
rect 2035 1126 2071 1130
rect 2075 1126 2119 1130
rect 2123 1126 2155 1130
rect 1125 1125 2155 1126
rect 2161 1125 2162 1131
rect 1398 1100 1404 1101
rect 1550 1100 1556 1101
rect 1398 1096 1399 1100
rect 1403 1096 1551 1100
rect 1555 1096 1556 1100
rect 1398 1095 1404 1096
rect 1550 1095 1556 1096
rect 84 1085 85 1091
rect 91 1090 1107 1091
rect 91 1086 111 1090
rect 115 1086 159 1090
rect 163 1086 199 1090
rect 203 1086 247 1090
rect 251 1086 303 1090
rect 307 1086 367 1090
rect 371 1086 431 1090
rect 435 1086 439 1090
rect 443 1086 503 1090
rect 507 1086 511 1090
rect 515 1086 575 1090
rect 579 1086 591 1090
rect 595 1086 647 1090
rect 651 1086 679 1090
rect 683 1086 719 1090
rect 723 1086 775 1090
rect 779 1086 783 1090
rect 787 1086 839 1090
rect 843 1086 879 1090
rect 883 1086 895 1090
rect 899 1086 951 1090
rect 955 1086 991 1090
rect 995 1086 1007 1090
rect 1011 1086 1047 1090
rect 1051 1086 1095 1090
rect 1099 1086 1107 1090
rect 91 1085 1107 1086
rect 1113 1085 1114 1091
rect 1106 1073 1107 1079
rect 1113 1078 2143 1079
rect 1113 1074 1135 1078
rect 1139 1074 1159 1078
rect 1163 1074 1247 1078
rect 1251 1074 1359 1078
rect 1363 1074 1383 1078
rect 1387 1074 1423 1078
rect 1427 1074 1471 1078
rect 1475 1074 1527 1078
rect 1531 1074 1575 1078
rect 1579 1074 1591 1078
rect 1595 1074 1655 1078
rect 1659 1074 1671 1078
rect 1675 1074 1711 1078
rect 1715 1074 1759 1078
rect 1763 1074 1767 1078
rect 1771 1074 1823 1078
rect 1827 1074 1847 1078
rect 1851 1074 1871 1078
rect 1875 1074 1927 1078
rect 1931 1074 1983 1078
rect 1987 1074 2007 1078
rect 2011 1074 2031 1078
rect 2035 1074 2071 1078
rect 2075 1074 2119 1078
rect 2123 1074 2143 1078
rect 1113 1073 2143 1074
rect 2149 1073 2150 1079
rect 96 1029 97 1035
rect 103 1034 1119 1035
rect 103 1030 111 1034
rect 115 1030 199 1034
rect 203 1030 223 1034
rect 227 1030 247 1034
rect 251 1030 271 1034
rect 275 1030 303 1034
rect 307 1030 335 1034
rect 339 1030 367 1034
rect 371 1030 407 1034
rect 411 1030 431 1034
rect 435 1030 479 1034
rect 483 1030 503 1034
rect 507 1030 559 1034
rect 563 1030 575 1034
rect 579 1030 631 1034
rect 635 1030 647 1034
rect 651 1030 703 1034
rect 707 1030 719 1034
rect 723 1030 775 1034
rect 779 1030 783 1034
rect 787 1030 839 1034
rect 843 1030 895 1034
rect 899 1030 903 1034
rect 907 1030 951 1034
rect 955 1030 967 1034
rect 971 1030 1007 1034
rect 1011 1030 1039 1034
rect 1043 1030 1047 1034
rect 1051 1030 1095 1034
rect 1099 1030 1119 1034
rect 103 1029 1119 1030
rect 1125 1029 1126 1035
rect 1118 1027 1126 1029
rect 1118 1021 1119 1027
rect 1125 1026 2155 1027
rect 1125 1022 1135 1026
rect 1139 1022 1159 1026
rect 1163 1022 1231 1026
rect 1235 1022 1247 1026
rect 1251 1022 1303 1026
rect 1307 1022 1359 1026
rect 1363 1022 1383 1026
rect 1387 1022 1463 1026
rect 1467 1022 1471 1026
rect 1475 1022 1543 1026
rect 1547 1022 1575 1026
rect 1579 1022 1623 1026
rect 1627 1022 1671 1026
rect 1675 1022 1695 1026
rect 1699 1022 1759 1026
rect 1763 1022 1823 1026
rect 1827 1022 1847 1026
rect 1851 1022 1887 1026
rect 1891 1022 1927 1026
rect 1931 1022 1951 1026
rect 1955 1022 2007 1026
rect 2011 1022 2071 1026
rect 2075 1022 2119 1026
rect 2123 1022 2155 1026
rect 1125 1021 2155 1022
rect 2161 1021 2162 1027
rect 84 973 85 979
rect 91 978 1107 979
rect 91 974 111 978
rect 115 974 151 978
rect 155 974 215 978
rect 219 974 223 978
rect 227 974 271 978
rect 275 974 287 978
rect 291 974 335 978
rect 339 974 367 978
rect 371 974 407 978
rect 411 974 447 978
rect 451 974 479 978
rect 483 974 527 978
rect 531 974 559 978
rect 563 974 599 978
rect 603 974 631 978
rect 635 974 671 978
rect 675 974 703 978
rect 707 974 735 978
rect 739 974 775 978
rect 779 974 799 978
rect 803 974 839 978
rect 843 974 863 978
rect 867 974 903 978
rect 907 974 927 978
rect 931 974 967 978
rect 971 974 991 978
rect 995 974 1039 978
rect 1043 974 1047 978
rect 1051 974 1095 978
rect 1099 974 1107 978
rect 91 973 1107 974
rect 1113 975 1114 979
rect 1113 974 2150 975
rect 1113 973 1135 974
rect 1106 970 1135 973
rect 1139 970 1159 974
rect 1163 970 1231 974
rect 1235 970 1239 974
rect 1243 970 1303 974
rect 1307 970 1375 974
rect 1379 970 1383 974
rect 1387 970 1439 974
rect 1443 970 1463 974
rect 1467 970 1511 974
rect 1515 970 1543 974
rect 1547 970 1583 974
rect 1587 970 1623 974
rect 1627 970 1655 974
rect 1659 970 1695 974
rect 1699 970 1727 974
rect 1731 970 1759 974
rect 1763 970 1799 974
rect 1803 970 1823 974
rect 1827 970 1871 974
rect 1875 970 1887 974
rect 1891 970 1943 974
rect 1947 970 1951 974
rect 1955 970 2015 974
rect 2019 970 2071 974
rect 2075 970 2119 974
rect 2123 970 2150 974
rect 1106 969 2150 970
rect 96 921 97 927
rect 103 926 1119 927
rect 103 922 111 926
rect 115 922 135 926
rect 139 922 151 926
rect 155 922 183 926
rect 187 922 215 926
rect 219 922 255 926
rect 259 922 287 926
rect 291 922 327 926
rect 331 922 367 926
rect 371 922 399 926
rect 403 922 447 926
rect 451 922 463 926
rect 467 922 527 926
rect 531 922 599 926
rect 603 922 671 926
rect 675 922 735 926
rect 739 922 743 926
rect 747 922 799 926
rect 803 922 815 926
rect 819 922 863 926
rect 867 922 895 926
rect 899 922 927 926
rect 931 922 983 926
rect 987 922 991 926
rect 995 922 1047 926
rect 1051 922 1095 926
rect 1099 922 1119 926
rect 103 921 1119 922
rect 1125 921 1126 927
rect 1118 919 1126 921
rect 1118 913 1119 919
rect 1125 918 2155 919
rect 1125 914 1135 918
rect 1139 914 1239 918
rect 1243 914 1287 918
rect 1291 914 1303 918
rect 1307 914 1327 918
rect 1331 914 1375 918
rect 1379 914 1423 918
rect 1427 914 1439 918
rect 1443 914 1479 918
rect 1483 914 1511 918
rect 1515 914 1551 918
rect 1555 914 1583 918
rect 1587 914 1623 918
rect 1627 914 1655 918
rect 1659 914 1703 918
rect 1707 914 1727 918
rect 1731 914 1791 918
rect 1795 914 1799 918
rect 1803 914 1871 918
rect 1875 914 1879 918
rect 1883 914 1943 918
rect 1947 914 1967 918
rect 1971 914 2015 918
rect 2019 914 2063 918
rect 2067 914 2071 918
rect 2075 914 2119 918
rect 2123 914 2155 918
rect 1125 913 2155 914
rect 2161 913 2162 919
rect 84 865 85 871
rect 91 870 1107 871
rect 91 866 111 870
rect 115 866 135 870
rect 139 866 175 870
rect 179 866 183 870
rect 187 866 215 870
rect 219 866 255 870
rect 259 866 279 870
rect 283 866 327 870
rect 331 866 343 870
rect 347 866 399 870
rect 403 866 463 870
rect 467 866 527 870
rect 531 866 535 870
rect 539 866 599 870
rect 603 866 615 870
rect 619 866 671 870
rect 675 866 711 870
rect 715 866 743 870
rect 747 866 815 870
rect 819 866 823 870
rect 827 866 895 870
rect 899 866 943 870
rect 947 866 983 870
rect 987 866 1047 870
rect 1051 866 1095 870
rect 1099 866 1107 870
rect 91 865 1107 866
rect 1113 867 1114 871
rect 1113 866 2150 867
rect 1113 865 1135 866
rect 1106 862 1135 865
rect 1139 862 1159 866
rect 1163 862 1199 866
rect 1203 862 1263 866
rect 1267 862 1287 866
rect 1291 862 1327 866
rect 1331 862 1375 866
rect 1379 862 1399 866
rect 1403 862 1423 866
rect 1427 862 1471 866
rect 1475 862 1479 866
rect 1483 862 1543 866
rect 1547 862 1551 866
rect 1555 862 1623 866
rect 1627 862 1703 866
rect 1707 862 1775 866
rect 1779 862 1791 866
rect 1795 862 1855 866
rect 1859 862 1879 866
rect 1883 862 1935 866
rect 1939 862 1967 866
rect 1971 862 2015 866
rect 2019 862 2063 866
rect 2067 862 2071 866
rect 2075 862 2119 866
rect 2123 862 2150 866
rect 1106 861 2150 862
rect 546 852 552 853
rect 846 852 852 853
rect 546 848 547 852
rect 551 848 847 852
rect 851 848 852 852
rect 546 847 552 848
rect 846 847 852 848
rect 478 828 484 829
rect 858 828 864 829
rect 478 824 479 828
rect 483 824 859 828
rect 863 824 864 828
rect 478 823 484 824
rect 858 823 864 824
rect 96 813 97 819
rect 103 818 1119 819
rect 103 814 111 818
rect 115 814 135 818
rect 139 814 175 818
rect 179 814 215 818
rect 219 814 279 818
rect 283 814 335 818
rect 339 814 343 818
rect 347 814 391 818
rect 395 814 399 818
rect 403 814 455 818
rect 459 814 463 818
rect 467 814 519 818
rect 523 814 535 818
rect 539 814 583 818
rect 587 814 615 818
rect 619 814 655 818
rect 659 814 711 818
rect 715 814 735 818
rect 739 814 815 818
rect 819 814 823 818
rect 827 814 895 818
rect 899 814 943 818
rect 947 814 983 818
rect 987 814 1047 818
rect 1051 814 1095 818
rect 1099 814 1119 818
rect 103 813 1119 814
rect 1125 813 1126 819
rect 1118 801 1119 807
rect 1125 806 2155 807
rect 1125 802 1135 806
rect 1139 802 1159 806
rect 1163 802 1199 806
rect 1203 802 1239 806
rect 1243 802 1263 806
rect 1267 802 1327 806
rect 1331 802 1343 806
rect 1347 802 1399 806
rect 1403 802 1447 806
rect 1451 802 1471 806
rect 1475 802 1543 806
rect 1547 802 1551 806
rect 1555 802 1623 806
rect 1627 802 1655 806
rect 1659 802 1703 806
rect 1707 802 1751 806
rect 1755 802 1775 806
rect 1779 802 1839 806
rect 1843 802 1855 806
rect 1859 802 1919 806
rect 1923 802 1935 806
rect 1939 802 2007 806
rect 2011 802 2015 806
rect 2019 802 2071 806
rect 2075 802 2119 806
rect 2123 802 2155 806
rect 1125 801 2155 802
rect 2161 801 2162 807
rect 84 761 85 767
rect 91 766 1107 767
rect 91 762 111 766
rect 115 762 135 766
rect 139 762 175 766
rect 179 762 207 766
rect 211 762 215 766
rect 219 762 279 766
rect 283 762 295 766
rect 299 762 335 766
rect 339 762 375 766
rect 379 762 391 766
rect 395 762 447 766
rect 451 762 455 766
rect 459 762 519 766
rect 523 762 583 766
rect 587 762 639 766
rect 643 762 655 766
rect 659 762 687 766
rect 691 762 735 766
rect 739 762 743 766
rect 747 762 799 766
rect 803 762 815 766
rect 819 762 855 766
rect 859 762 895 766
rect 899 762 983 766
rect 987 762 1047 766
rect 1051 762 1095 766
rect 1099 762 1107 766
rect 91 761 1107 762
rect 1113 761 1114 767
rect 1106 749 1107 755
rect 1113 754 2143 755
rect 1113 750 1135 754
rect 1139 750 1159 754
rect 1163 750 1199 754
rect 1203 750 1239 754
rect 1243 750 1287 754
rect 1291 750 1343 754
rect 1347 750 1359 754
rect 1363 750 1439 754
rect 1443 750 1447 754
rect 1451 750 1527 754
rect 1531 750 1551 754
rect 1555 750 1615 754
rect 1619 750 1655 754
rect 1659 750 1711 754
rect 1715 750 1751 754
rect 1755 750 1807 754
rect 1811 750 1839 754
rect 1843 750 1903 754
rect 1907 750 1919 754
rect 1923 750 1999 754
rect 2003 750 2007 754
rect 2011 750 2071 754
rect 2075 750 2119 754
rect 2123 750 2143 754
rect 1113 749 2143 750
rect 2149 749 2150 755
rect 96 705 97 711
rect 103 710 1119 711
rect 103 706 111 710
rect 115 706 135 710
rect 139 706 183 710
rect 187 706 207 710
rect 211 706 247 710
rect 251 706 295 710
rect 299 706 311 710
rect 315 706 375 710
rect 379 706 383 710
rect 387 706 447 710
rect 451 706 455 710
rect 459 706 519 710
rect 523 706 583 710
rect 587 706 639 710
rect 643 706 647 710
rect 651 706 687 710
rect 691 706 711 710
rect 715 706 743 710
rect 747 706 767 710
rect 771 706 799 710
rect 803 706 823 710
rect 827 706 855 710
rect 859 706 879 710
rect 883 706 943 710
rect 947 706 1095 710
rect 1099 706 1119 710
rect 103 705 1119 706
rect 1125 705 1126 711
rect 1118 693 1119 699
rect 1125 698 2155 699
rect 1125 694 1135 698
rect 1139 694 1159 698
rect 1163 694 1199 698
rect 1203 694 1239 698
rect 1243 694 1287 698
rect 1291 694 1335 698
rect 1339 694 1359 698
rect 1363 694 1391 698
rect 1395 694 1439 698
rect 1443 694 1447 698
rect 1451 694 1511 698
rect 1515 694 1527 698
rect 1531 694 1575 698
rect 1579 694 1615 698
rect 1619 694 1639 698
rect 1643 694 1703 698
rect 1707 694 1711 698
rect 1715 694 1767 698
rect 1771 694 1807 698
rect 1811 694 1831 698
rect 1835 694 1895 698
rect 1899 694 1903 698
rect 1907 694 1959 698
rect 1963 694 1999 698
rect 2003 694 2023 698
rect 2027 694 2071 698
rect 2075 694 2119 698
rect 2123 694 2155 698
rect 1125 693 2155 694
rect 2161 693 2162 699
rect 734 684 740 685
rect 966 684 972 685
rect 734 680 735 684
rect 739 680 967 684
rect 971 680 972 684
rect 734 679 740 680
rect 966 679 972 680
rect 84 645 85 651
rect 91 650 1107 651
rect 91 646 111 650
rect 115 646 135 650
rect 139 646 159 650
rect 163 646 183 650
rect 187 646 215 650
rect 219 646 247 650
rect 251 646 287 650
rect 291 646 311 650
rect 315 646 367 650
rect 371 646 383 650
rect 387 646 455 650
rect 459 646 519 650
rect 523 646 543 650
rect 547 646 583 650
rect 587 646 631 650
rect 635 646 647 650
rect 651 646 711 650
rect 715 646 719 650
rect 723 646 767 650
rect 771 646 799 650
rect 803 646 823 650
rect 827 646 871 650
rect 875 646 879 650
rect 883 646 943 650
rect 947 646 951 650
rect 955 646 1031 650
rect 1035 646 1095 650
rect 1099 646 1107 650
rect 91 645 1107 646
rect 1113 647 1114 651
rect 1113 646 2150 647
rect 1113 645 1135 646
rect 1106 642 1135 645
rect 1139 642 1239 646
rect 1243 642 1279 646
rect 1283 642 1287 646
rect 1291 642 1319 646
rect 1323 642 1335 646
rect 1339 642 1367 646
rect 1371 642 1391 646
rect 1395 642 1423 646
rect 1427 642 1447 646
rect 1451 642 1479 646
rect 1483 642 1511 646
rect 1515 642 1535 646
rect 1539 642 1575 646
rect 1579 642 1591 646
rect 1595 642 1639 646
rect 1643 642 1647 646
rect 1651 642 1703 646
rect 1707 642 1719 646
rect 1723 642 1767 646
rect 1771 642 1799 646
rect 1803 642 1831 646
rect 1835 642 1879 646
rect 1883 642 1895 646
rect 1899 642 1959 646
rect 1963 642 1967 646
rect 1971 642 2023 646
rect 2027 642 2063 646
rect 2067 642 2071 646
rect 2075 642 2119 646
rect 2123 642 2150 646
rect 1106 641 2150 642
rect 726 612 732 613
rect 1038 612 1044 613
rect 726 608 727 612
rect 731 608 1039 612
rect 1043 608 1044 612
rect 726 607 732 608
rect 1038 607 1044 608
rect 96 589 97 595
rect 103 594 1119 595
rect 103 590 111 594
rect 115 590 159 594
rect 163 590 207 594
rect 211 590 215 594
rect 219 590 255 594
rect 259 590 287 594
rect 291 590 311 594
rect 315 590 367 594
rect 371 590 383 594
rect 387 590 455 594
rect 459 590 463 594
rect 467 590 543 594
rect 547 590 623 594
rect 627 590 631 594
rect 635 590 703 594
rect 707 590 719 594
rect 723 590 783 594
rect 787 590 799 594
rect 803 590 855 594
rect 859 590 871 594
rect 875 590 927 594
rect 931 590 951 594
rect 955 590 999 594
rect 1003 590 1031 594
rect 1035 590 1047 594
rect 1051 590 1095 594
rect 1099 590 1119 594
rect 103 589 1119 590
rect 1125 594 2162 595
rect 1125 590 1135 594
rect 1139 590 1279 594
rect 1283 590 1319 594
rect 1323 590 1335 594
rect 1339 590 1367 594
rect 1371 590 1375 594
rect 1379 590 1415 594
rect 1419 590 1423 594
rect 1427 590 1463 594
rect 1467 590 1479 594
rect 1483 590 1519 594
rect 1523 590 1535 594
rect 1539 590 1583 594
rect 1587 590 1591 594
rect 1595 590 1647 594
rect 1651 590 1655 594
rect 1659 590 1719 594
rect 1723 590 1727 594
rect 1731 590 1799 594
rect 1803 590 1807 594
rect 1811 590 1879 594
rect 1883 590 1887 594
rect 1891 590 1967 594
rect 1971 590 1975 594
rect 1979 590 2063 594
rect 2067 590 2119 594
rect 2123 590 2162 594
rect 1125 589 2162 590
rect 1106 538 2150 539
rect 1106 535 1135 538
rect 84 529 85 535
rect 91 534 1107 535
rect 91 530 111 534
rect 115 530 159 534
rect 163 530 167 534
rect 171 530 207 534
rect 211 530 223 534
rect 227 530 255 534
rect 259 530 287 534
rect 291 530 311 534
rect 315 530 359 534
rect 363 530 383 534
rect 387 530 431 534
rect 435 530 463 534
rect 467 530 511 534
rect 515 530 543 534
rect 547 530 591 534
rect 595 530 623 534
rect 627 530 663 534
rect 667 530 703 534
rect 707 530 735 534
rect 739 530 783 534
rect 787 530 807 534
rect 811 530 855 534
rect 859 530 871 534
rect 875 530 927 534
rect 931 530 935 534
rect 939 530 999 534
rect 1003 530 1047 534
rect 1051 530 1095 534
rect 1099 530 1107 534
rect 91 529 1107 530
rect 1113 534 1135 535
rect 1139 534 1191 538
rect 1195 534 1239 538
rect 1243 534 1287 538
rect 1291 534 1335 538
rect 1339 534 1343 538
rect 1347 534 1375 538
rect 1379 534 1407 538
rect 1411 534 1415 538
rect 1419 534 1463 538
rect 1467 534 1479 538
rect 1483 534 1519 538
rect 1523 534 1543 538
rect 1547 534 1583 538
rect 1587 534 1607 538
rect 1611 534 1655 538
rect 1659 534 1671 538
rect 1675 534 1727 538
rect 1731 534 1735 538
rect 1739 534 1799 538
rect 1803 534 1807 538
rect 1811 534 1863 538
rect 1867 534 1887 538
rect 1891 534 1935 538
rect 1939 534 1975 538
rect 1979 534 2007 538
rect 2011 534 2063 538
rect 2067 534 2071 538
rect 2075 534 2119 538
rect 2123 534 2150 538
rect 1113 533 2150 534
rect 1113 529 1114 533
rect 1118 486 2162 487
rect 1118 483 1135 486
rect 96 477 97 483
rect 103 482 1119 483
rect 103 478 111 482
rect 115 478 167 482
rect 171 478 223 482
rect 227 478 231 482
rect 235 478 287 482
rect 291 478 303 482
rect 307 478 359 482
rect 363 478 375 482
rect 379 478 431 482
rect 435 478 455 482
rect 459 478 511 482
rect 515 478 535 482
rect 539 478 591 482
rect 595 478 607 482
rect 611 478 663 482
rect 667 478 679 482
rect 683 478 735 482
rect 739 478 743 482
rect 747 478 799 482
rect 803 478 807 482
rect 811 478 855 482
rect 859 478 871 482
rect 875 478 903 482
rect 907 478 935 482
rect 939 478 959 482
rect 963 478 999 482
rect 1003 478 1007 482
rect 1011 478 1047 482
rect 1051 478 1095 482
rect 1099 478 1119 482
rect 103 477 1119 478
rect 1125 482 1135 483
rect 1139 482 1159 486
rect 1163 482 1191 486
rect 1195 482 1239 486
rect 1243 482 1263 486
rect 1267 482 1287 486
rect 1291 482 1343 486
rect 1347 482 1383 486
rect 1387 482 1407 486
rect 1411 482 1479 486
rect 1483 482 1495 486
rect 1499 482 1543 486
rect 1547 482 1599 486
rect 1603 482 1607 486
rect 1611 482 1671 486
rect 1675 482 1703 486
rect 1707 482 1735 486
rect 1739 482 1799 486
rect 1803 482 1863 486
rect 1867 482 1887 486
rect 1891 482 1935 486
rect 1939 482 1983 486
rect 1987 482 2007 486
rect 2011 482 2071 486
rect 2075 482 2119 486
rect 2123 482 2162 486
rect 1125 481 2162 482
rect 1125 477 1126 481
rect 1106 434 2150 435
rect 1106 431 1135 434
rect 84 425 85 431
rect 91 430 1107 431
rect 91 426 111 430
rect 115 426 151 430
rect 155 426 167 430
rect 171 426 215 430
rect 219 426 231 430
rect 235 426 279 430
rect 283 426 303 430
rect 307 426 351 430
rect 355 426 375 430
rect 379 426 423 430
rect 427 426 455 430
rect 459 426 487 430
rect 491 426 535 430
rect 539 426 551 430
rect 555 426 607 430
rect 611 426 615 430
rect 619 426 671 430
rect 675 426 679 430
rect 683 426 727 430
rect 731 426 743 430
rect 747 426 791 430
rect 795 426 799 430
rect 803 426 855 430
rect 859 426 903 430
rect 907 426 959 430
rect 963 426 1007 430
rect 1011 426 1047 430
rect 1051 426 1095 430
rect 1099 426 1107 430
rect 91 425 1107 426
rect 1113 430 1135 431
rect 1139 430 1159 434
rect 1163 430 1199 434
rect 1203 430 1255 434
rect 1259 430 1263 434
rect 1267 430 1335 434
rect 1339 430 1383 434
rect 1387 430 1415 434
rect 1419 430 1495 434
rect 1499 430 1503 434
rect 1507 430 1591 434
rect 1595 430 1599 434
rect 1603 430 1671 434
rect 1675 430 1703 434
rect 1707 430 1751 434
rect 1755 430 1799 434
rect 1803 430 1823 434
rect 1827 430 1887 434
rect 1891 430 1951 434
rect 1955 430 1983 434
rect 1987 430 2023 434
rect 2027 430 2071 434
rect 2075 430 2119 434
rect 2123 430 2150 434
rect 1113 429 2150 430
rect 1113 425 1114 429
rect 96 373 97 379
rect 103 378 1119 379
rect 103 374 111 378
rect 115 374 135 378
rect 139 374 151 378
rect 155 374 175 378
rect 179 374 215 378
rect 219 374 271 378
rect 275 374 279 378
rect 283 374 335 378
rect 339 374 351 378
rect 355 374 399 378
rect 403 374 423 378
rect 427 374 463 378
rect 467 374 487 378
rect 491 374 519 378
rect 523 374 551 378
rect 555 374 575 378
rect 579 374 615 378
rect 619 374 631 378
rect 635 374 671 378
rect 675 374 687 378
rect 691 374 727 378
rect 731 374 751 378
rect 755 374 791 378
rect 795 374 855 378
rect 859 374 1095 378
rect 1099 374 1119 378
rect 103 373 1119 374
rect 1125 378 2162 379
rect 1125 374 1135 378
rect 1139 374 1159 378
rect 1163 374 1199 378
rect 1203 374 1255 378
rect 1259 374 1303 378
rect 1307 374 1335 378
rect 1339 374 1343 378
rect 1347 374 1383 378
rect 1387 374 1415 378
rect 1419 374 1423 378
rect 1427 374 1463 378
rect 1467 374 1503 378
rect 1507 374 1551 378
rect 1555 374 1591 378
rect 1595 374 1615 378
rect 1619 374 1671 378
rect 1675 374 1679 378
rect 1683 374 1751 378
rect 1755 374 1823 378
rect 1827 374 1831 378
rect 1835 374 1887 378
rect 1891 374 1919 378
rect 1923 374 1951 378
rect 1955 374 2007 378
rect 2011 374 2023 378
rect 2027 374 2071 378
rect 2075 374 2119 378
rect 2123 374 2162 378
rect 1125 373 2162 374
rect 84 317 85 323
rect 91 322 1107 323
rect 91 318 111 322
rect 115 318 135 322
rect 139 318 175 322
rect 179 318 207 322
rect 211 318 215 322
rect 219 318 271 322
rect 275 318 295 322
rect 299 318 335 322
rect 339 318 383 322
rect 387 318 399 322
rect 403 318 463 322
rect 467 318 471 322
rect 475 318 519 322
rect 523 318 551 322
rect 555 318 575 322
rect 579 318 623 322
rect 627 318 631 322
rect 635 318 687 322
rect 691 318 751 322
rect 755 318 807 322
rect 811 318 871 322
rect 875 318 935 322
rect 939 318 1095 322
rect 1099 318 1107 322
rect 91 317 1107 318
rect 1113 322 2150 323
rect 1113 318 1135 322
rect 1139 318 1167 322
rect 1171 318 1207 322
rect 1211 318 1247 322
rect 1251 318 1295 322
rect 1299 318 1303 322
rect 1307 318 1343 322
rect 1347 318 1383 322
rect 1387 318 1391 322
rect 1395 318 1423 322
rect 1427 318 1439 322
rect 1443 318 1463 322
rect 1467 318 1495 322
rect 1499 318 1503 322
rect 1507 318 1551 322
rect 1555 318 1559 322
rect 1563 318 1615 322
rect 1619 318 1623 322
rect 1627 318 1679 322
rect 1683 318 1695 322
rect 1699 318 1751 322
rect 1755 318 1775 322
rect 1779 318 1831 322
rect 1835 318 1855 322
rect 1859 318 1919 322
rect 1923 318 1935 322
rect 1939 318 2007 322
rect 2011 318 2015 322
rect 2019 318 2071 322
rect 2075 318 2119 322
rect 2123 318 2150 322
rect 1113 317 2150 318
rect 96 265 97 271
rect 103 270 1119 271
rect 103 266 111 270
rect 115 266 135 270
rect 139 266 199 270
rect 203 266 207 270
rect 211 266 279 270
rect 283 266 295 270
rect 299 266 359 270
rect 363 266 383 270
rect 387 266 439 270
rect 443 266 471 270
rect 475 266 511 270
rect 515 266 551 270
rect 555 266 583 270
rect 587 266 623 270
rect 627 266 647 270
rect 651 266 687 270
rect 691 266 703 270
rect 707 266 751 270
rect 755 266 759 270
rect 763 266 807 270
rect 811 266 815 270
rect 819 266 871 270
rect 875 266 879 270
rect 883 266 935 270
rect 939 266 1095 270
rect 1099 266 1119 270
rect 103 265 1119 266
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 262 2155 263
rect 1125 258 1135 262
rect 1139 258 1159 262
rect 1163 258 1167 262
rect 1171 258 1207 262
rect 1211 258 1247 262
rect 1251 258 1271 262
rect 1275 258 1295 262
rect 1299 258 1327 262
rect 1331 258 1343 262
rect 1347 258 1391 262
rect 1395 258 1439 262
rect 1443 258 1455 262
rect 1459 258 1495 262
rect 1499 258 1527 262
rect 1531 258 1559 262
rect 1563 258 1607 262
rect 1611 258 1623 262
rect 1627 258 1687 262
rect 1691 258 1695 262
rect 1699 258 1767 262
rect 1771 258 1775 262
rect 1779 258 1839 262
rect 1843 258 1855 262
rect 1859 258 1919 262
rect 1923 258 1935 262
rect 1939 258 1999 262
rect 2003 258 2015 262
rect 2019 258 2071 262
rect 2075 258 2119 262
rect 2123 258 2155 262
rect 1125 257 2155 258
rect 2161 257 2162 263
rect 84 209 85 215
rect 91 214 1107 215
rect 91 210 111 214
rect 115 210 135 214
rect 139 210 183 214
rect 187 210 199 214
rect 203 210 231 214
rect 235 210 279 214
rect 283 210 327 214
rect 331 210 359 214
rect 363 210 375 214
rect 379 210 415 214
rect 419 210 439 214
rect 443 210 455 214
rect 459 210 503 214
rect 507 210 511 214
rect 515 210 551 214
rect 555 210 583 214
rect 587 210 599 214
rect 603 210 647 214
rect 651 210 695 214
rect 699 210 703 214
rect 707 210 743 214
rect 747 210 759 214
rect 763 210 815 214
rect 819 210 879 214
rect 883 210 1095 214
rect 1099 210 1107 214
rect 91 209 1107 210
rect 1113 211 1114 215
rect 1113 210 2150 211
rect 1113 209 1135 210
rect 1106 206 1135 209
rect 1139 206 1159 210
rect 1163 206 1199 210
rect 1203 206 1207 210
rect 1211 206 1263 210
rect 1267 206 1271 210
rect 1275 206 1327 210
rect 1331 206 1391 210
rect 1395 206 1399 210
rect 1403 206 1455 210
rect 1459 206 1471 210
rect 1475 206 1527 210
rect 1531 206 1543 210
rect 1547 206 1607 210
rect 1611 206 1671 210
rect 1675 206 1687 210
rect 1691 206 1735 210
rect 1739 206 1767 210
rect 1771 206 1807 210
rect 1811 206 1839 210
rect 1843 206 1879 210
rect 1883 206 1919 210
rect 1923 206 1951 210
rect 1955 206 1999 210
rect 2003 206 2023 210
rect 2027 206 2071 210
rect 2075 206 2119 210
rect 2123 206 2150 210
rect 1106 205 2150 206
rect 96 133 97 139
rect 103 138 1119 139
rect 103 134 111 138
rect 115 134 135 138
rect 139 134 143 138
rect 147 134 183 138
rect 187 134 223 138
rect 227 134 231 138
rect 235 134 263 138
rect 267 134 279 138
rect 283 134 303 138
rect 307 134 327 138
rect 331 134 343 138
rect 347 134 375 138
rect 379 134 383 138
rect 387 134 415 138
rect 419 134 423 138
rect 427 134 455 138
rect 459 134 463 138
rect 467 134 503 138
rect 507 134 543 138
rect 547 134 551 138
rect 555 134 583 138
rect 587 134 599 138
rect 603 134 623 138
rect 627 134 647 138
rect 651 134 663 138
rect 667 134 695 138
rect 699 134 703 138
rect 707 134 743 138
rect 747 134 783 138
rect 787 134 831 138
rect 835 134 879 138
rect 883 134 927 138
rect 931 134 967 138
rect 971 134 1007 138
rect 1011 134 1047 138
rect 1051 134 1095 138
rect 1099 134 1119 138
rect 103 133 1119 134
rect 1125 138 2162 139
rect 1125 134 1135 138
rect 1139 134 1159 138
rect 1163 134 1199 138
rect 1203 134 1207 138
rect 1211 134 1263 138
rect 1267 134 1271 138
rect 1275 134 1327 138
rect 1331 134 1335 138
rect 1339 134 1399 138
rect 1403 134 1455 138
rect 1459 134 1471 138
rect 1475 134 1511 138
rect 1515 134 1543 138
rect 1547 134 1559 138
rect 1563 134 1607 138
rect 1611 134 1647 138
rect 1651 134 1671 138
rect 1675 134 1687 138
rect 1691 134 1727 138
rect 1731 134 1735 138
rect 1739 134 1767 138
rect 1771 134 1807 138
rect 1811 134 1855 138
rect 1859 134 1879 138
rect 1883 134 1903 138
rect 1907 134 1951 138
rect 1955 134 1991 138
rect 1995 134 2023 138
rect 2027 134 2031 138
rect 2035 134 2071 138
rect 2075 134 2119 138
rect 2123 134 2162 138
rect 1125 133 2162 134
rect 84 81 85 87
rect 91 86 1107 87
rect 91 82 111 86
rect 115 82 143 86
rect 147 82 183 86
rect 187 82 223 86
rect 227 82 263 86
rect 267 82 303 86
rect 307 82 343 86
rect 347 82 383 86
rect 387 82 423 86
rect 427 82 463 86
rect 467 82 503 86
rect 507 82 543 86
rect 547 82 583 86
rect 587 82 623 86
rect 627 82 663 86
rect 667 82 703 86
rect 707 82 743 86
rect 747 82 783 86
rect 787 82 831 86
rect 835 82 879 86
rect 883 82 927 86
rect 931 82 967 86
rect 971 82 1007 86
rect 1011 82 1047 86
rect 1051 82 1095 86
rect 1099 82 1107 86
rect 91 81 1107 82
rect 1113 86 2150 87
rect 1113 82 1135 86
rect 1139 82 1159 86
rect 1163 82 1207 86
rect 1211 82 1271 86
rect 1275 82 1335 86
rect 1339 82 1399 86
rect 1403 82 1455 86
rect 1459 82 1511 86
rect 1515 82 1559 86
rect 1563 82 1607 86
rect 1611 82 1647 86
rect 1651 82 1687 86
rect 1691 82 1727 86
rect 1731 82 1767 86
rect 1771 82 1807 86
rect 1811 82 1855 86
rect 1859 82 1903 86
rect 1907 82 1951 86
rect 1955 82 1991 86
rect 1995 82 2031 86
rect 2035 82 2071 86
rect 2075 82 2119 86
rect 2123 82 2150 86
rect 1113 81 2150 82
<< m5c >>
rect 1119 2225 1125 2231
rect 2155 2225 2161 2231
rect 85 2209 91 2215
rect 1107 2209 1113 2215
rect 1107 2173 1113 2179
rect 2143 2173 2149 2179
rect 97 2149 103 2155
rect 1119 2149 1125 2155
rect 1119 2121 1125 2127
rect 2155 2121 2161 2127
rect 85 2093 91 2099
rect 1107 2093 1113 2099
rect 1107 2069 1113 2075
rect 2143 2069 2149 2075
rect 97 2037 103 2043
rect 1119 2037 1125 2043
rect 1119 2017 1125 2023
rect 2155 2017 2161 2023
rect 85 1985 91 1991
rect 1107 1985 1113 1991
rect 1107 1953 1113 1959
rect 2143 1953 2149 1959
rect 97 1929 103 1935
rect 1119 1929 1125 1935
rect 1119 1901 1125 1907
rect 2155 1901 2161 1907
rect 85 1873 91 1879
rect 1107 1873 1113 1879
rect 1107 1845 1113 1851
rect 2143 1845 2149 1851
rect 97 1817 103 1823
rect 1119 1817 1125 1823
rect 1119 1785 1125 1791
rect 2155 1785 2161 1791
rect 85 1757 91 1763
rect 1107 1757 1113 1763
rect 1107 1729 1113 1735
rect 2143 1729 2149 1735
rect 97 1701 103 1707
rect 1119 1701 1125 1707
rect 1119 1677 1125 1683
rect 2155 1677 2161 1683
rect 85 1645 91 1651
rect 1107 1645 1113 1651
rect 1107 1621 1113 1627
rect 2143 1621 2149 1627
rect 97 1585 103 1591
rect 1119 1585 1125 1591
rect 1119 1569 1125 1575
rect 2155 1569 2161 1575
rect 85 1525 91 1531
rect 1107 1525 1113 1531
rect 1107 1513 1113 1519
rect 2143 1513 2149 1519
rect 97 1465 103 1471
rect 1119 1465 1125 1471
rect 85 1409 91 1415
rect 1107 1409 1113 1415
rect 97 1357 103 1363
rect 1119 1357 1125 1363
rect 1119 1349 1125 1355
rect 2155 1349 2161 1355
rect 85 1305 91 1311
rect 1107 1305 1113 1311
rect 1107 1293 1113 1299
rect 2143 1293 2149 1299
rect 97 1249 103 1255
rect 1119 1249 1125 1255
rect 1119 1237 1125 1243
rect 2155 1237 2161 1243
rect 85 1197 91 1203
rect 1107 1197 1113 1203
rect 1107 1185 1113 1191
rect 2143 1185 2149 1191
rect 97 1145 103 1151
rect 1119 1145 1125 1151
rect 1119 1125 1125 1131
rect 2155 1125 2161 1131
rect 85 1085 91 1091
rect 1107 1085 1113 1091
rect 1107 1073 1113 1079
rect 2143 1073 2149 1079
rect 97 1029 103 1035
rect 1119 1029 1125 1035
rect 1119 1021 1125 1027
rect 2155 1021 2161 1027
rect 85 973 91 979
rect 1107 973 1113 979
rect 97 921 103 927
rect 1119 921 1125 927
rect 1119 913 1125 919
rect 2155 913 2161 919
rect 85 865 91 871
rect 1107 865 1113 871
rect 97 813 103 819
rect 1119 813 1125 819
rect 1119 801 1125 807
rect 2155 801 2161 807
rect 85 761 91 767
rect 1107 761 1113 767
rect 1107 749 1113 755
rect 2143 749 2149 755
rect 97 705 103 711
rect 1119 705 1125 711
rect 1119 693 1125 699
rect 2155 693 2161 699
rect 85 645 91 651
rect 1107 645 1113 651
rect 97 589 103 595
rect 1119 589 1125 595
rect 85 529 91 535
rect 1107 529 1113 535
rect 97 477 103 483
rect 1119 477 1125 483
rect 85 425 91 431
rect 1107 425 1113 431
rect 97 373 103 379
rect 1119 373 1125 379
rect 85 317 91 323
rect 1107 317 1113 323
rect 97 265 103 271
rect 1119 265 1125 271
rect 1119 257 1125 263
rect 2155 257 2161 263
rect 85 209 91 215
rect 1107 209 1113 215
rect 97 133 103 139
rect 1119 133 1125 139
rect 85 81 91 87
rect 1107 81 1113 87
<< m5 >>
rect 84 2215 92 2232
rect 84 2209 85 2215
rect 91 2209 92 2215
rect 84 2099 92 2209
rect 84 2093 85 2099
rect 91 2093 92 2099
rect 84 1991 92 2093
rect 84 1985 85 1991
rect 91 1985 92 1991
rect 84 1879 92 1985
rect 84 1873 85 1879
rect 91 1873 92 1879
rect 84 1763 92 1873
rect 84 1757 85 1763
rect 91 1757 92 1763
rect 84 1651 92 1757
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1531 92 1645
rect 84 1525 85 1531
rect 91 1525 92 1531
rect 84 1415 92 1525
rect 84 1409 85 1415
rect 91 1409 92 1415
rect 84 1311 92 1409
rect 84 1305 85 1311
rect 91 1305 92 1311
rect 84 1203 92 1305
rect 84 1197 85 1203
rect 91 1197 92 1203
rect 84 1091 92 1197
rect 84 1085 85 1091
rect 91 1085 92 1091
rect 84 979 92 1085
rect 84 973 85 979
rect 91 973 92 979
rect 84 871 92 973
rect 84 865 85 871
rect 91 865 92 871
rect 84 767 92 865
rect 84 761 85 767
rect 91 761 92 767
rect 84 651 92 761
rect 84 645 85 651
rect 91 645 92 651
rect 84 535 92 645
rect 84 529 85 535
rect 91 529 92 535
rect 84 431 92 529
rect 84 425 85 431
rect 91 425 92 431
rect 84 323 92 425
rect 84 317 85 323
rect 91 317 92 323
rect 84 215 92 317
rect 84 209 85 215
rect 91 209 92 215
rect 84 87 92 209
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2155 104 2232
rect 96 2149 97 2155
rect 103 2149 104 2155
rect 96 2043 104 2149
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1935 104 2037
rect 96 1929 97 1935
rect 103 1929 104 1935
rect 96 1823 104 1929
rect 96 1817 97 1823
rect 103 1817 104 1823
rect 96 1707 104 1817
rect 96 1701 97 1707
rect 103 1701 104 1707
rect 96 1591 104 1701
rect 96 1585 97 1591
rect 103 1585 104 1591
rect 96 1471 104 1585
rect 96 1465 97 1471
rect 103 1465 104 1471
rect 96 1363 104 1465
rect 96 1357 97 1363
rect 103 1357 104 1363
rect 96 1255 104 1357
rect 96 1249 97 1255
rect 103 1249 104 1255
rect 96 1151 104 1249
rect 96 1145 97 1151
rect 103 1145 104 1151
rect 96 1035 104 1145
rect 96 1029 97 1035
rect 103 1029 104 1035
rect 96 927 104 1029
rect 96 921 97 927
rect 103 921 104 927
rect 96 819 104 921
rect 96 813 97 819
rect 103 813 104 819
rect 96 711 104 813
rect 96 705 97 711
rect 103 705 104 711
rect 96 595 104 705
rect 96 589 97 595
rect 103 589 104 595
rect 96 483 104 589
rect 96 477 97 483
rect 103 477 104 483
rect 96 379 104 477
rect 96 373 97 379
rect 103 373 104 379
rect 96 271 104 373
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1106 2215 1114 2232
rect 1106 2209 1107 2215
rect 1113 2209 1114 2215
rect 1106 2179 1114 2209
rect 1106 2173 1107 2179
rect 1113 2173 1114 2179
rect 1106 2099 1114 2173
rect 1106 2093 1107 2099
rect 1113 2093 1114 2099
rect 1106 2075 1114 2093
rect 1106 2069 1107 2075
rect 1113 2069 1114 2075
rect 1106 1991 1114 2069
rect 1106 1985 1107 1991
rect 1113 1985 1114 1991
rect 1106 1959 1114 1985
rect 1106 1953 1107 1959
rect 1113 1953 1114 1959
rect 1106 1879 1114 1953
rect 1106 1873 1107 1879
rect 1113 1873 1114 1879
rect 1106 1851 1114 1873
rect 1106 1845 1107 1851
rect 1113 1845 1114 1851
rect 1106 1763 1114 1845
rect 1106 1757 1107 1763
rect 1113 1757 1114 1763
rect 1106 1735 1114 1757
rect 1106 1729 1107 1735
rect 1113 1729 1114 1735
rect 1106 1651 1114 1729
rect 1106 1645 1107 1651
rect 1113 1645 1114 1651
rect 1106 1627 1114 1645
rect 1106 1621 1107 1627
rect 1113 1621 1114 1627
rect 1106 1531 1114 1621
rect 1106 1525 1107 1531
rect 1113 1525 1114 1531
rect 1106 1519 1114 1525
rect 1106 1513 1107 1519
rect 1113 1513 1114 1519
rect 1106 1415 1114 1513
rect 1106 1409 1107 1415
rect 1113 1409 1114 1415
rect 1106 1311 1114 1409
rect 1106 1305 1107 1311
rect 1113 1305 1114 1311
rect 1106 1299 1114 1305
rect 1106 1293 1107 1299
rect 1113 1293 1114 1299
rect 1106 1203 1114 1293
rect 1106 1197 1107 1203
rect 1113 1197 1114 1203
rect 1106 1191 1114 1197
rect 1106 1185 1107 1191
rect 1113 1185 1114 1191
rect 1106 1091 1114 1185
rect 1106 1085 1107 1091
rect 1113 1085 1114 1091
rect 1106 1079 1114 1085
rect 1106 1073 1107 1079
rect 1113 1073 1114 1079
rect 1106 979 1114 1073
rect 1106 973 1107 979
rect 1113 973 1114 979
rect 1106 871 1114 973
rect 1106 865 1107 871
rect 1113 865 1114 871
rect 1106 767 1114 865
rect 1106 761 1107 767
rect 1113 761 1114 767
rect 1106 755 1114 761
rect 1106 749 1107 755
rect 1113 749 1114 755
rect 1106 651 1114 749
rect 1106 645 1107 651
rect 1113 645 1114 651
rect 1106 535 1114 645
rect 1106 529 1107 535
rect 1113 529 1114 535
rect 1106 431 1114 529
rect 1106 425 1107 431
rect 1113 425 1114 431
rect 1106 323 1114 425
rect 1106 317 1107 323
rect 1113 317 1114 323
rect 1106 215 1114 317
rect 1106 209 1107 215
rect 1113 209 1114 215
rect 1106 87 1114 209
rect 1106 81 1107 87
rect 1113 81 1114 87
rect 1106 72 1114 81
rect 1118 2231 1126 2232
rect 1118 2225 1119 2231
rect 1125 2225 1126 2231
rect 1118 2155 1126 2225
rect 1118 2149 1119 2155
rect 1125 2149 1126 2155
rect 1118 2127 1126 2149
rect 1118 2121 1119 2127
rect 1125 2121 1126 2127
rect 1118 2043 1126 2121
rect 1118 2037 1119 2043
rect 1125 2037 1126 2043
rect 1118 2023 1126 2037
rect 1118 2017 1119 2023
rect 1125 2017 1126 2023
rect 1118 1935 1126 2017
rect 1118 1929 1119 1935
rect 1125 1929 1126 1935
rect 1118 1907 1126 1929
rect 1118 1901 1119 1907
rect 1125 1901 1126 1907
rect 1118 1823 1126 1901
rect 1118 1817 1119 1823
rect 1125 1817 1126 1823
rect 1118 1791 1126 1817
rect 1118 1785 1119 1791
rect 1125 1785 1126 1791
rect 1118 1707 1126 1785
rect 1118 1701 1119 1707
rect 1125 1701 1126 1707
rect 1118 1683 1126 1701
rect 1118 1677 1119 1683
rect 1125 1677 1126 1683
rect 1118 1591 1126 1677
rect 1118 1585 1119 1591
rect 1125 1585 1126 1591
rect 1118 1575 1126 1585
rect 1118 1569 1119 1575
rect 1125 1569 1126 1575
rect 1118 1471 1126 1569
rect 1118 1465 1119 1471
rect 1125 1465 1126 1471
rect 1118 1363 1126 1465
rect 1118 1357 1119 1363
rect 1125 1357 1126 1363
rect 1118 1355 1126 1357
rect 1118 1349 1119 1355
rect 1125 1349 1126 1355
rect 1118 1255 1126 1349
rect 1118 1249 1119 1255
rect 1125 1249 1126 1255
rect 1118 1243 1126 1249
rect 1118 1237 1119 1243
rect 1125 1237 1126 1243
rect 1118 1151 1126 1237
rect 1118 1145 1119 1151
rect 1125 1145 1126 1151
rect 1118 1131 1126 1145
rect 1118 1125 1119 1131
rect 1125 1125 1126 1131
rect 1118 1035 1126 1125
rect 1118 1029 1119 1035
rect 1125 1029 1126 1035
rect 1118 1027 1126 1029
rect 1118 1021 1119 1027
rect 1125 1021 1126 1027
rect 1118 927 1126 1021
rect 1118 921 1119 927
rect 1125 921 1126 927
rect 1118 919 1126 921
rect 1118 913 1119 919
rect 1125 913 1126 919
rect 1118 819 1126 913
rect 1118 813 1119 819
rect 1125 813 1126 819
rect 1118 807 1126 813
rect 1118 801 1119 807
rect 1125 801 1126 807
rect 1118 711 1126 801
rect 1118 705 1119 711
rect 1125 705 1126 711
rect 1118 699 1126 705
rect 1118 693 1119 699
rect 1125 693 1126 699
rect 1118 595 1126 693
rect 1118 589 1119 595
rect 1125 589 1126 595
rect 1118 483 1126 589
rect 1118 477 1119 483
rect 1125 477 1126 483
rect 1118 379 1126 477
rect 1118 373 1119 379
rect 1125 373 1126 379
rect 1118 271 1126 373
rect 1118 265 1119 271
rect 1125 265 1126 271
rect 1118 263 1126 265
rect 1118 257 1119 263
rect 1125 257 1126 263
rect 1118 139 1126 257
rect 1118 133 1119 139
rect 1125 133 1126 139
rect 1118 72 1126 133
rect 2142 2179 2150 2232
rect 2142 2173 2143 2179
rect 2149 2173 2150 2179
rect 2142 2075 2150 2173
rect 2142 2069 2143 2075
rect 2149 2069 2150 2075
rect 2142 1959 2150 2069
rect 2142 1953 2143 1959
rect 2149 1953 2150 1959
rect 2142 1851 2150 1953
rect 2142 1845 2143 1851
rect 2149 1845 2150 1851
rect 2142 1735 2150 1845
rect 2142 1729 2143 1735
rect 2149 1729 2150 1735
rect 2142 1627 2150 1729
rect 2142 1621 2143 1627
rect 2149 1621 2150 1627
rect 2142 1519 2150 1621
rect 2142 1513 2143 1519
rect 2149 1513 2150 1519
rect 2142 1299 2150 1513
rect 2142 1293 2143 1299
rect 2149 1293 2150 1299
rect 2142 1191 2150 1293
rect 2142 1185 2143 1191
rect 2149 1185 2150 1191
rect 2142 1079 2150 1185
rect 2142 1073 2143 1079
rect 2149 1073 2150 1079
rect 2142 755 2150 1073
rect 2142 749 2143 755
rect 2149 749 2150 755
rect 2142 72 2150 749
rect 2154 2231 2162 2232
rect 2154 2225 2155 2231
rect 2161 2225 2162 2231
rect 2154 2127 2162 2225
rect 2154 2121 2155 2127
rect 2161 2121 2162 2127
rect 2154 2023 2162 2121
rect 2154 2017 2155 2023
rect 2161 2017 2162 2023
rect 2154 1907 2162 2017
rect 2154 1901 2155 1907
rect 2161 1901 2162 1907
rect 2154 1791 2162 1901
rect 2154 1785 2155 1791
rect 2161 1785 2162 1791
rect 2154 1683 2162 1785
rect 2154 1677 2155 1683
rect 2161 1677 2162 1683
rect 2154 1575 2162 1677
rect 2154 1569 2155 1575
rect 2161 1569 2162 1575
rect 2154 1355 2162 1569
rect 2154 1349 2155 1355
rect 2161 1349 2162 1355
rect 2154 1243 2162 1349
rect 2154 1237 2155 1243
rect 2161 1237 2162 1243
rect 2154 1131 2162 1237
rect 2154 1125 2155 1131
rect 2161 1125 2162 1131
rect 2154 1027 2162 1125
rect 2154 1021 2155 1027
rect 2161 1021 2162 1027
rect 2154 919 2162 1021
rect 2154 913 2155 919
rect 2161 913 2162 919
rect 2154 807 2162 913
rect 2154 801 2155 807
rect 2161 801 2162 807
rect 2154 699 2162 801
rect 2154 693 2155 699
rect 2161 693 2162 699
rect 2154 263 2162 693
rect 2154 257 2155 263
rect 2161 257 2162 263
rect 2154 72 2162 257
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__153
timestamp 1731220628
transform 1 0 2112 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220628
transform 1 0 1128 0 1 2180
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220628
transform 1 0 2112 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220628
transform 1 0 1128 0 -1 2172
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220628
transform 1 0 2112 0 1 2076
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220628
transform 1 0 1128 0 1 2076
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220628
transform 1 0 2112 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220628
transform 1 0 1128 0 -1 2068
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220628
transform 1 0 2112 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220628
transform 1 0 1128 0 1 1972
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220628
transform 1 0 2112 0 -1 1952
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220628
transform 1 0 1128 0 -1 1952
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220628
transform 1 0 2112 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220628
transform 1 0 1128 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220628
transform 1 0 2112 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220628
transform 1 0 1128 0 -1 1844
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220628
transform 1 0 2112 0 1 1740
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220628
transform 1 0 1128 0 1 1740
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220628
transform 1 0 2112 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220628
transform 1 0 1128 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220628
transform 1 0 2112 0 1 1632
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220628
transform 1 0 1128 0 1 1632
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220628
transform 1 0 2112 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220628
transform 1 0 1128 0 -1 1620
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220628
transform 1 0 2112 0 1 1524
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220628
transform 1 0 1128 0 1 1524
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220628
transform 1 0 2112 0 -1 1512
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220628
transform 1 0 1128 0 -1 1512
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220628
transform 1 0 2112 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220628
transform 1 0 1128 0 1 1416
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220628
transform 1 0 2112 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220628
transform 1 0 1128 0 -1 1404
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220628
transform 1 0 2112 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220628
transform 1 0 1128 0 1 1304
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220628
transform 1 0 2112 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220628
transform 1 0 1128 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220628
transform 1 0 2112 0 1 1192
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220628
transform 1 0 1128 0 1 1192
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220628
transform 1 0 2112 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220628
transform 1 0 1128 0 -1 1184
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220628
transform 1 0 2112 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220628
transform 1 0 1128 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220628
transform 1 0 2112 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220628
transform 1 0 1128 0 -1 1072
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220628
transform 1 0 2112 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220628
transform 1 0 1128 0 1 976
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220628
transform 1 0 2112 0 -1 968
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220628
transform 1 0 1128 0 -1 968
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220628
transform 1 0 2112 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220628
transform 1 0 1128 0 1 868
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220628
transform 1 0 2112 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220628
transform 1 0 1128 0 -1 860
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220628
transform 1 0 2112 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220628
transform 1 0 1128 0 1 756
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220628
transform 1 0 2112 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220628
transform 1 0 1128 0 -1 748
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220628
transform 1 0 2112 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220628
transform 1 0 1128 0 1 648
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220628
transform 1 0 2112 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220628
transform 1 0 1128 0 -1 640
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220628
transform 1 0 2112 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220628
transform 1 0 1128 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220628
transform 1 0 2112 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220628
transform 1 0 1128 0 -1 532
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220628
transform 1 0 2112 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220628
transform 1 0 1128 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220628
transform 1 0 2112 0 -1 428
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220628
transform 1 0 1128 0 -1 428
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220628
transform 1 0 2112 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220628
transform 1 0 1128 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220628
transform 1 0 2112 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220628
transform 1 0 1128 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220628
transform 1 0 2112 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220628
transform 1 0 1128 0 1 212
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220628
transform 1 0 2112 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220628
transform 1 0 1128 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220628
transform 1 0 2112 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220628
transform 1 0 1128 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220628
transform 1 0 1088 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220628
transform 1 0 104 0 -1 2208
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220628
transform 1 0 1088 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220628
transform 1 0 104 0 1 2104
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220628
transform 1 0 1088 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220628
transform 1 0 104 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220628
transform 1 0 1088 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220628
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220628
transform 1 0 1088 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220628
transform 1 0 104 0 -1 1984
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220628
transform 1 0 1088 0 1 1884
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220628
transform 1 0 104 0 1 1884
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220628
transform 1 0 1088 0 -1 1872
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220628
transform 1 0 104 0 -1 1872
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220628
transform 1 0 1088 0 1 1772
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220628
transform 1 0 104 0 1 1772
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220628
transform 1 0 1088 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220628
transform 1 0 104 0 -1 1756
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220628
transform 1 0 1088 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220628
transform 1 0 104 0 1 1656
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220628
transform 1 0 1088 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220628
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220628
transform 1 0 1088 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220628
transform 1 0 104 0 1 1540
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220628
transform 1 0 1088 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220628
transform 1 0 104 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220628
transform 1 0 1088 0 1 1420
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220628
transform 1 0 104 0 1 1420
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220628
transform 1 0 1088 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220628
transform 1 0 104 0 -1 1408
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220628
transform 1 0 1088 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220628
transform 1 0 104 0 1 1312
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220628
transform 1 0 1088 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220628
transform 1 0 104 0 -1 1304
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220628
transform 1 0 1088 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220628
transform 1 0 104 0 1 1204
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220628
transform 1 0 1088 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220628
transform 1 0 104 0 -1 1196
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220628
transform 1 0 1088 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220628
transform 1 0 104 0 1 1100
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220628
transform 1 0 1088 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220628
transform 1 0 104 0 -1 1084
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220628
transform 1 0 1088 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220628
transform 1 0 104 0 1 984
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220628
transform 1 0 1088 0 -1 972
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220628
transform 1 0 104 0 -1 972
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220628
transform 1 0 1088 0 1 876
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220628
transform 1 0 104 0 1 876
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220628
transform 1 0 1088 0 -1 864
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220628
transform 1 0 104 0 -1 864
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220628
transform 1 0 1088 0 1 768
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220628
transform 1 0 104 0 1 768
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220628
transform 1 0 1088 0 -1 760
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220628
transform 1 0 104 0 -1 760
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220628
transform 1 0 1088 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220628
transform 1 0 104 0 1 660
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220628
transform 1 0 1088 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220628
transform 1 0 104 0 -1 644
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220628
transform 1 0 1088 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220628
transform 1 0 104 0 1 544
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220628
transform 1 0 1088 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220628
transform 1 0 104 0 -1 528
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220628
transform 1 0 1088 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220628
transform 1 0 104 0 1 432
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220628
transform 1 0 1088 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220628
transform 1 0 104 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220628
transform 1 0 1088 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220628
transform 1 0 104 0 1 328
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220628
transform 1 0 1088 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220628
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220628
transform 1 0 1088 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220628
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220628
transform 1 0 1088 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220628
transform 1 0 104 0 -1 208
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220628
transform 1 0 1088 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220628
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0NOR2X1  tst_5999_6
timestamp 1731220628
transform 1 0 1984 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5998_6
timestamp 1731220628
transform 1 0 2024 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5997_6
timestamp 1731220628
transform 1 0 2064 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5996_6
timestamp 1731220628
transform 1 0 2064 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5995_6
timestamp 1731220628
transform 1 0 2064 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5994_6
timestamp 1731220628
transform 1 0 1992 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5993_6
timestamp 1731220628
transform 1 0 2008 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5992_6
timestamp 1731220628
transform 1 0 2064 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5991_6
timestamp 1731220628
transform 1 0 2064 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5990_6
timestamp 1731220628
transform 1 0 2064 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5989_6
timestamp 1731220628
transform 1 0 2016 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5988_6
timestamp 1731220628
transform 1 0 2064 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5987_6
timestamp 1731220628
transform 1 0 2064 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5986_6
timestamp 1731220628
transform 1 0 2000 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5985_6
timestamp 1731220628
transform 1 0 1968 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5984_6
timestamp 1731220628
transform 1 0 2056 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5983_6
timestamp 1731220628
transform 1 0 2056 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5982_6
timestamp 1731220628
transform 1 0 2016 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5981_6
timestamp 1731220628
transform 1 0 2064 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5980_6
timestamp 1731220628
transform 1 0 2064 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5979_6
timestamp 1731220628
transform 1 0 2064 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5978_6
timestamp 1731220628
transform 1 0 2064 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5977_6
timestamp 1731220628
transform 1 0 2008 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5976_6
timestamp 1731220628
transform 1 0 1936 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5975_6
timestamp 1731220628
transform 1 0 2008 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5974_6
timestamp 1731220628
transform 1 0 2064 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5973_6
timestamp 1731220628
transform 1 0 2056 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5972_6
timestamp 1731220628
transform 1 0 1960 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5971_6
timestamp 1731220628
transform 1 0 1872 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5970_6
timestamp 1731220628
transform 1 0 1848 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5969_6
timestamp 1731220628
transform 1 0 1928 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5968_6
timestamp 1731220628
transform 1 0 2000 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5967_6
timestamp 1731220628
transform 1 0 1912 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5966_6
timestamp 1731220628
transform 1 0 1832 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5965_6
timestamp 1731220628
transform 1 0 1800 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5964_6
timestamp 1731220628
transform 1 0 1896 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5963_6
timestamp 1731220628
transform 1 0 1992 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5962_6
timestamp 1731220628
transform 1 0 1952 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5961_6
timestamp 1731220628
transform 1 0 1888 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5960_6
timestamp 1731220628
transform 1 0 1824 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5959_6
timestamp 1731220628
transform 1 0 1760 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5958_6
timestamp 1731220628
transform 1 0 1696 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5957_6
timestamp 1731220628
transform 1 0 1960 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5956_6
timestamp 1731220628
transform 1 0 1872 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5955_6
timestamp 1731220628
transform 1 0 1792 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5954_6
timestamp 1731220628
transform 1 0 1712 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5953_6
timestamp 1731220628
transform 1 0 1640 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5952_6
timestamp 1731220628
transform 1 0 1584 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5951_6
timestamp 1731220628
transform 1 0 1720 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5950_6
timestamp 1731220628
transform 1 0 1800 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5949_6
timestamp 1731220628
transform 1 0 1880 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5948_6
timestamp 1731220628
transform 1 0 1856 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5947_6
timestamp 1731220628
transform 1 0 1792 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5946_6
timestamp 1731220628
transform 1 0 1728 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5945_6
timestamp 1731220628
transform 1 0 1928 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5944_6
timestamp 1731220628
transform 1 0 1976 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5943_6
timestamp 1731220628
transform 1 0 1880 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5942_6
timestamp 1731220628
transform 1 0 1792 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5941_6
timestamp 1731220628
transform 1 0 1816 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5940_6
timestamp 1731220628
transform 1 0 1880 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5939_6
timestamp 1731220628
transform 1 0 1944 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5938_6
timestamp 1731220628
transform 1 0 2000 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5937_6
timestamp 1731220628
transform 1 0 1912 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5936_6
timestamp 1731220628
transform 1 0 1928 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5935_6
timestamp 1731220628
transform 1 0 1848 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5934_6
timestamp 1731220628
transform 1 0 1832 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5933_6
timestamp 1731220628
transform 1 0 1912 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5932_6
timestamp 1731220628
transform 1 0 2016 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5931_6
timestamp 1731220628
transform 1 0 1944 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5930_6
timestamp 1731220628
transform 1 0 1872 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5929_6
timestamp 1731220628
transform 1 0 1800 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5928_6
timestamp 1731220628
transform 1 0 1944 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5927_6
timestamp 1731220628
transform 1 0 1896 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5926_6
timestamp 1731220628
transform 1 0 1848 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5925_6
timestamp 1731220628
transform 1 0 1800 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5924_6
timestamp 1731220628
transform 1 0 1760 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5923_6
timestamp 1731220628
transform 1 0 1720 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5922_6
timestamp 1731220628
transform 1 0 1680 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5921_6
timestamp 1731220628
transform 1 0 1640 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5920_6
timestamp 1731220628
transform 1 0 1600 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5919_6
timestamp 1731220628
transform 1 0 1552 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5918_6
timestamp 1731220628
transform 1 0 1600 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5917_6
timestamp 1731220628
transform 1 0 1664 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5916_6
timestamp 1731220628
transform 1 0 1728 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5915_6
timestamp 1731220628
transform 1 0 1760 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5914_6
timestamp 1731220628
transform 1 0 1680 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5913_6
timestamp 1731220628
transform 1 0 1600 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5912_6
timestamp 1731220628
transform 1 0 1688 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5911_6
timestamp 1731220628
transform 1 0 1768 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5910_6
timestamp 1731220628
transform 1 0 1824 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5909_6
timestamp 1731220628
transform 1 0 1744 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5908_6
timestamp 1731220628
transform 1 0 1664 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5907_6
timestamp 1731220628
transform 1 0 1584 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5906_6
timestamp 1731220628
transform 1 0 1488 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5905_6
timestamp 1731220628
transform 1 0 1592 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5904_6
timestamp 1731220628
transform 1 0 1696 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5903_6
timestamp 1731220628
transform 1 0 1664 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5902_6
timestamp 1731220628
transform 1 0 1600 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5901_6
timestamp 1731220628
transform 1 0 1536 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5900_6
timestamp 1731220628
transform 1 0 1648 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5899_6
timestamp 1731220628
transform 1 0 1576 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5898_6
timestamp 1731220628
transform 1 0 1528 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5897_6
timestamp 1731220628
transform 1 0 1472 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5896_6
timestamp 1731220628
transform 1 0 1440 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5895_6
timestamp 1731220628
transform 1 0 1384 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5894_6
timestamp 1731220628
transform 1 0 1504 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5893_6
timestamp 1731220628
transform 1 0 1568 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5892_6
timestamp 1731220628
transform 1 0 1632 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5891_6
timestamp 1731220628
transform 1 0 1704 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5890_6
timestamp 1731220628
transform 1 0 1608 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5889_6
timestamp 1731220628
transform 1 0 1520 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5888_6
timestamp 1731220628
transform 1 0 1440 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5887_6
timestamp 1731220628
transform 1 0 1544 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5886_6
timestamp 1731220628
transform 1 0 1648 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5885_6
timestamp 1731220628
transform 1 0 1744 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5884_6
timestamp 1731220628
transform 1 0 1768 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5883_6
timestamp 1731220628
transform 1 0 1696 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5882_6
timestamp 1731220628
transform 1 0 1616 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5881_6
timestamp 1731220628
transform 1 0 1536 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5880_6
timestamp 1731220628
transform 1 0 1544 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5879_6
timestamp 1731220628
transform 1 0 1616 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5878_6
timestamp 1731220628
transform 1 0 1696 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5877_6
timestamp 1731220628
transform 1 0 1784 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5876_6
timestamp 1731220628
transform 1 0 1720 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5875_6
timestamp 1731220628
transform 1 0 1648 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5874_6
timestamp 1731220628
transform 1 0 1576 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5873_6
timestamp 1731220628
transform 1 0 1864 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5872_6
timestamp 1731220628
transform 1 0 1792 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5871_6
timestamp 1731220628
transform 1 0 1752 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5870_6
timestamp 1731220628
transform 1 0 1688 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5869_6
timestamp 1731220628
transform 1 0 1616 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5868_6
timestamp 1731220628
transform 1 0 1944 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5867_6
timestamp 1731220628
transform 1 0 1880 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5866_6
timestamp 1731220628
transform 1 0 1816 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5865_6
timestamp 1731220628
transform 1 0 1752 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5864_6
timestamp 1731220628
transform 1 0 1664 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5863_6
timestamp 1731220628
transform 1 0 1840 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5862_6
timestamp 1731220628
transform 1 0 1920 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5861_6
timestamp 1731220628
transform 1 0 2000 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5860_6
timestamp 1731220628
transform 1 0 1976 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5859_6
timestamp 1731220628
transform 1 0 1920 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5858_6
timestamp 1731220628
transform 1 0 1864 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5857_6
timestamp 1731220628
transform 1 0 1816 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5856_6
timestamp 1731220628
transform 1 0 1760 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5855_6
timestamp 1731220628
transform 1 0 1704 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5854_6
timestamp 1731220628
transform 1 0 1912 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5853_6
timestamp 1731220628
transform 1 0 1832 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5852_6
timestamp 1731220628
transform 1 0 1760 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5851_6
timestamp 1731220628
transform 1 0 1696 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5850_6
timestamp 1731220628
transform 1 0 1632 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5849_6
timestamp 1731220628
transform 1 0 1576 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5848_6
timestamp 1731220628
transform 1 0 1712 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5847_6
timestamp 1731220628
transform 1 0 1608 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5846_6
timestamp 1731220628
transform 1 0 1528 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5845_6
timestamp 1731220628
transform 1 0 1464 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5844_6
timestamp 1731220628
transform 1 0 1960 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5843_6
timestamp 1731220628
transform 1 0 1832 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5842_6
timestamp 1731220628
transform 1 0 1712 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5841_6
timestamp 1731220628
transform 1 0 1632 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5840_6
timestamp 1731220628
transform 1 0 1552 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5839_6
timestamp 1731220628
transform 1 0 1792 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5838_6
timestamp 1731220628
transform 1 0 1872 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5837_6
timestamp 1731220628
transform 1 0 1960 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5836_6
timestamp 1731220628
transform 1 0 1896 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5835_6
timestamp 1731220628
transform 1 0 1960 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5834_6
timestamp 1731220628
transform 1 0 2024 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5833_6
timestamp 1731220628
transform 1 0 2048 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5832_6
timestamp 1731220628
transform 1 0 2000 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5831_6
timestamp 1731220628
transform 1 0 2024 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5830_6
timestamp 1731220628
transform 1 0 2064 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5829_6
timestamp 1731220628
transform 1 0 2064 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5828_6
timestamp 1731220628
transform 1 0 2064 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5827_6
timestamp 1731220628
transform 1 0 2064 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5826_6
timestamp 1731220628
transform 1 0 2064 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5825_6
timestamp 1731220628
transform 1 0 2064 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5824_6
timestamp 1731220628
transform 1 0 2064 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5823_6
timestamp 1731220628
transform 1 0 2064 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5822_6
timestamp 1731220628
transform 1 0 1984 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5821_6
timestamp 1731220628
transform 1 0 2008 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5820_6
timestamp 1731220628
transform 1 0 1936 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5819_6
timestamp 1731220628
transform 1 0 1824 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5818_6
timestamp 1731220628
transform 1 0 1752 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5817_6
timestamp 1731220628
transform 1 0 1672 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5816_6
timestamp 1731220628
transform 1 0 1584 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5815_6
timestamp 1731220628
transform 1 0 1864 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5814_6
timestamp 1731220628
transform 1 0 1792 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5813_6
timestamp 1731220628
transform 1 0 1712 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5812_6
timestamp 1731220628
transform 1 0 1624 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5811_6
timestamp 1731220628
transform 1 0 1984 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5810_6
timestamp 1731220628
transform 1 0 1888 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5809_6
timestamp 1731220628
transform 1 0 1800 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5808_6
timestamp 1731220628
transform 1 0 1712 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5807_6
timestamp 1731220628
transform 1 0 1640 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5806_6
timestamp 1731220628
transform 1 0 1576 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5805_6
timestamp 1731220628
transform 1 0 1896 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5804_6
timestamp 1731220628
transform 1 0 1808 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5803_6
timestamp 1731220628
transform 1 0 1728 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5802_6
timestamp 1731220628
transform 1 0 1656 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5801_6
timestamp 1731220628
transform 1 0 1600 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5800_6
timestamp 1731220628
transform 1 0 1552 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5799_6
timestamp 1731220628
transform 1 0 1512 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5798_6
timestamp 1731220628
transform 1 0 1464 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5797_6
timestamp 1731220628
transform 1 0 1560 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5796_6
timestamp 1731220628
transform 1 0 1728 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5795_6
timestamp 1731220628
transform 1 0 1672 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5794_6
timestamp 1731220628
transform 1 0 1616 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5793_6
timestamp 1731220628
transform 1 0 1600 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5792_6
timestamp 1731220628
transform 1 0 1528 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5791_6
timestamp 1731220628
transform 1 0 1672 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5790_6
timestamp 1731220628
transform 1 0 1824 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5789_6
timestamp 1731220628
transform 1 0 1744 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5788_6
timestamp 1731220628
transform 1 0 1672 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5787_6
timestamp 1731220628
transform 1 0 1592 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5786_6
timestamp 1731220628
transform 1 0 1744 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5785_6
timestamp 1731220628
transform 1 0 1808 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5784_6
timestamp 1731220628
transform 1 0 1752 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5783_6
timestamp 1731220628
transform 1 0 1680 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5782_6
timestamp 1731220628
transform 1 0 1824 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5781_6
timestamp 1731220628
transform 1 0 1888 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5780_6
timestamp 1731220628
transform 1 0 1952 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5779_6
timestamp 1731220628
transform 1 0 2016 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5778_6
timestamp 1731220628
transform 1 0 1976 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5777_6
timestamp 1731220628
transform 1 0 1920 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5776_6
timestamp 1731220628
transform 1 0 1864 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5775_6
timestamp 1731220628
transform 1 0 2024 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5774_6
timestamp 1731220628
transform 1 0 2064 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5773_6
timestamp 1731220628
transform 1 0 2064 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5772_6
timestamp 1731220628
transform 1 0 2064 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5771_6
timestamp 1731220628
transform 1 0 2064 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5770_6
timestamp 1731220628
transform 1 0 1976 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5769_6
timestamp 1731220628
transform 1 0 2064 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5768_6
timestamp 1731220628
transform 1 0 2064 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5767_6
timestamp 1731220628
transform 1 0 2000 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5766_6
timestamp 1731220628
transform 1 0 2064 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5765_6
timestamp 1731220628
transform 1 0 2064 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5764_6
timestamp 1731220628
transform 1 0 2016 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5763_6
timestamp 1731220628
transform 1 0 2064 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5762_6
timestamp 1731220628
transform 1 0 2016 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5761_6
timestamp 1731220628
transform 1 0 1944 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5760_6
timestamp 1731220628
transform 1 0 1952 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5759_6
timestamp 1731220628
transform 1 0 2016 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5758_6
timestamp 1731220628
transform 1 0 1952 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5757_6
timestamp 1731220628
transform 1 0 1888 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5756_6
timestamp 1731220628
transform 1 0 1816 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5755_6
timestamp 1731220628
transform 1 0 1736 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5754_6
timestamp 1731220628
transform 1 0 1752 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5753_6
timestamp 1731220628
transform 1 0 1824 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5752_6
timestamp 1731220628
transform 1 0 1888 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5751_6
timestamp 1731220628
transform 1 0 1880 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5750_6
timestamp 1731220628
transform 1 0 1816 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5749_6
timestamp 1731220628
transform 1 0 1744 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5748_6
timestamp 1731220628
transform 1 0 1728 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5747_6
timestamp 1731220628
transform 1 0 1872 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5746_6
timestamp 1731220628
transform 1 0 1800 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5745_6
timestamp 1731220628
transform 1 0 1800 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5744_6
timestamp 1731220628
transform 1 0 1760 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5743_6
timestamp 1731220628
transform 1 0 1720 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5742_6
timestamp 1731220628
transform 1 0 1680 0 1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5741_6
timestamp 1731220628
transform 1 0 1656 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5740_6
timestamp 1731220628
transform 1 0 1584 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5739_6
timestamp 1731220628
transform 1 0 1672 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5738_6
timestamp 1731220628
transform 1 0 1592 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5737_6
timestamp 1731220628
transform 1 0 1584 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5736_6
timestamp 1731220628
transform 1 0 1672 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5735_6
timestamp 1731220628
transform 1 0 1648 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5734_6
timestamp 1731220628
transform 1 0 1624 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5733_6
timestamp 1731220628
transform 1 0 1696 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5732_6
timestamp 1731220628
transform 1 0 1768 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5731_6
timestamp 1731220628
transform 1 0 1840 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5730_6
timestamp 1731220628
transform 1 0 1920 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5729_6
timestamp 1731220628
transform 1 0 1968 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5728_6
timestamp 1731220628
transform 1 0 1856 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5727_6
timestamp 1731220628
transform 1 0 1744 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5726_6
timestamp 1731220628
transform 1 0 1648 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5725_6
timestamp 1731220628
transform 1 0 1568 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5724_6
timestamp 1731220628
transform 1 0 1864 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5723_6
timestamp 1731220628
transform 1 0 1760 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5722_6
timestamp 1731220628
transform 1 0 1664 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5721_6
timestamp 1731220628
transform 1 0 1576 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5720_6
timestamp 1731220628
transform 1 0 1496 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5719_6
timestamp 1731220628
transform 1 0 1424 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5718_6
timestamp 1731220628
transform 1 0 1976 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5717_6
timestamp 1731220628
transform 1 0 1864 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5716_6
timestamp 1731220628
transform 1 0 1760 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5715_6
timestamp 1731220628
transform 1 0 1672 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5714_6
timestamp 1731220628
transform 1 0 1600 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5713_6
timestamp 1731220628
transform 1 0 1544 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5712_6
timestamp 1731220628
transform 1 0 1504 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5711_6
timestamp 1731220628
transform 1 0 1464 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5710_6
timestamp 1731220628
transform 1 0 1424 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5709_6
timestamp 1731220628
transform 1 0 1384 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5708_6
timestamp 1731220628
transform 1 0 1344 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5707_6
timestamp 1731220628
transform 1 0 1304 0 1 1736
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5706_6
timestamp 1731220628
transform 1 0 1608 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5705_6
timestamp 1731220628
transform 1 0 1528 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5704_6
timestamp 1731220628
transform 1 0 1448 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5703_6
timestamp 1731220628
transform 1 0 1376 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5702_6
timestamp 1731220628
transform 1 0 1312 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5701_6
timestamp 1731220628
transform 1 0 1256 0 -1 1732
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5700_6
timestamp 1731220628
transform 1 0 1504 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5699_6
timestamp 1731220628
transform 1 0 1416 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5698_6
timestamp 1731220628
transform 1 0 1328 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5697_6
timestamp 1731220628
transform 1 0 1240 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5696_6
timestamp 1731220628
transform 1 0 1160 0 1 1628
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5695_6
timestamp 1731220628
transform 1 0 1312 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5694_6
timestamp 1731220628
transform 1 0 1240 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5693_6
timestamp 1731220628
transform 1 0 1192 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5692_6
timestamp 1731220628
transform 1 0 1152 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5691_6
timestamp 1731220628
transform 1 0 1456 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5690_6
timestamp 1731220628
transform 1 0 1384 0 -1 1624
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5689_6
timestamp 1731220628
transform 1 0 1320 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5688_6
timestamp 1731220628
transform 1 0 1272 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5687_6
timestamp 1731220628
transform 1 0 1232 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5686_6
timestamp 1731220628
transform 1 0 1368 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5685_6
timestamp 1731220628
transform 1 0 1416 0 1 1520
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5684_6
timestamp 1731220628
transform 1 0 1512 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5683_6
timestamp 1731220628
transform 1 0 1472 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5682_6
timestamp 1731220628
transform 1 0 1432 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5681_6
timestamp 1731220628
transform 1 0 1392 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5680_6
timestamp 1731220628
transform 1 0 1352 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5679_6
timestamp 1731220628
transform 1 0 1312 0 -1 1516
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5678_6
timestamp 1731220628
transform 1 0 1512 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5677_6
timestamp 1731220628
transform 1 0 1448 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5676_6
timestamp 1731220628
transform 1 0 1384 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5675_6
timestamp 1731220628
transform 1 0 1328 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5674_6
timestamp 1731220628
transform 1 0 1272 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5673_6
timestamp 1731220628
transform 1 0 1224 0 1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5672_6
timestamp 1731220628
transform 1 0 1536 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5671_6
timestamp 1731220628
transform 1 0 1440 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5670_6
timestamp 1731220628
transform 1 0 1344 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5669_6
timestamp 1731220628
transform 1 0 1256 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5668_6
timestamp 1731220628
transform 1 0 1192 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5667_6
timestamp 1731220628
transform 1 0 1152 0 -1 1408
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5666_6
timestamp 1731220628
transform 1 0 1480 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5665_6
timestamp 1731220628
transform 1 0 1368 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5664_6
timestamp 1731220628
transform 1 0 1248 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5663_6
timestamp 1731220628
transform 1 0 1152 0 1 1300
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5662_6
timestamp 1731220628
transform 1 0 1040 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5661_6
timestamp 1731220628
transform 1 0 1040 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5660_6
timestamp 1731220628
transform 1 0 1152 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5659_6
timestamp 1731220628
transform 1 0 1192 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5658_6
timestamp 1731220628
transform 1 0 1240 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5657_6
timestamp 1731220628
transform 1 0 1472 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5656_6
timestamp 1731220628
transform 1 0 1392 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5655_6
timestamp 1731220628
transform 1 0 1312 0 -1 1296
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5654_6
timestamp 1731220628
transform 1 0 1232 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5653_6
timestamp 1731220628
transform 1 0 1192 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5652_6
timestamp 1731220628
transform 1 0 1152 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5651_6
timestamp 1731220628
transform 1 0 1272 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5650_6
timestamp 1731220628
transform 1 0 1320 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5649_6
timestamp 1731220628
transform 1 0 1416 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5648_6
timestamp 1731220628
transform 1 0 1368 0 1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5647_6
timestamp 1731220628
transform 1 0 1360 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5646_6
timestamp 1731220628
transform 1 0 1320 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5645_6
timestamp 1731220628
transform 1 0 1280 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5644_6
timestamp 1731220628
transform 1 0 1408 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5643_6
timestamp 1731220628
transform 1 0 1520 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5642_6
timestamp 1731220628
transform 1 0 1464 0 -1 1188
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5641_6
timestamp 1731220628
transform 1 0 1464 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5640_6
timestamp 1731220628
transform 1 0 1416 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5639_6
timestamp 1731220628
transform 1 0 1376 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5638_6
timestamp 1731220628
transform 1 0 1520 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5637_6
timestamp 1731220628
transform 1 0 1648 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5636_6
timestamp 1731220628
transform 1 0 1584 0 1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5635_6
timestamp 1731220628
transform 1 0 1568 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5634_6
timestamp 1731220628
transform 1 0 1464 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5633_6
timestamp 1731220628
transform 1 0 1456 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5632_6
timestamp 1731220628
transform 1 0 1536 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5631_6
timestamp 1731220628
transform 1 0 1504 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5630_6
timestamp 1731220628
transform 1 0 1432 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5629_6
timestamp 1731220628
transform 1 0 1416 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5628_6
timestamp 1731220628
transform 1 0 1472 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5627_6
timestamp 1731220628
transform 1 0 1464 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5626_6
timestamp 1731220628
transform 1 0 1392 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5625_6
timestamp 1731220628
transform 1 0 1320 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5624_6
timestamp 1731220628
transform 1 0 1256 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5623_6
timestamp 1731220628
transform 1 0 1192 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5622_6
timestamp 1731220628
transform 1 0 1280 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5621_6
timestamp 1731220628
transform 1 0 1320 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5620_6
timestamp 1731220628
transform 1 0 1368 0 1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5619_6
timestamp 1731220628
transform 1 0 1368 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5618_6
timestamp 1731220628
transform 1 0 1296 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5617_6
timestamp 1731220628
transform 1 0 1232 0 -1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5616_6
timestamp 1731220628
transform 1 0 1376 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5615_6
timestamp 1731220628
transform 1 0 1296 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5614_6
timestamp 1731220628
transform 1 0 1224 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5613_6
timestamp 1731220628
transform 1 0 1152 0 1 972
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5612_6
timestamp 1731220628
transform 1 0 1352 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5611_6
timestamp 1731220628
transform 1 0 1240 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5610_6
timestamp 1731220628
transform 1 0 1152 0 -1 1076
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5609_6
timestamp 1731220628
transform 1 0 1040 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5608_6
timestamp 1731220628
transform 1 0 1000 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5607_6
timestamp 1731220628
transform 1 0 944 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5606_6
timestamp 1731220628
transform 1 0 888 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5605_6
timestamp 1731220628
transform 1 0 896 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5604_6
timestamp 1731220628
transform 1 0 832 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5603_6
timestamp 1731220628
transform 1 0 768 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5602_6
timestamp 1731220628
transform 1 0 696 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5601_6
timestamp 1731220628
transform 1 0 920 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5600_6
timestamp 1731220628
transform 1 0 856 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5599_6
timestamp 1731220628
transform 1 0 792 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5598_6
timestamp 1731220628
transform 1 0 728 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5597_6
timestamp 1731220628
transform 1 0 664 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5596_6
timestamp 1731220628
transform 1 0 592 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5595_6
timestamp 1731220628
transform 1 0 888 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5594_6
timestamp 1731220628
transform 1 0 808 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5593_6
timestamp 1731220628
transform 1 0 736 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5592_6
timestamp 1731220628
transform 1 0 664 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5591_6
timestamp 1731220628
transform 1 0 592 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5590_6
timestamp 1731220628
transform 1 0 520 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5589_6
timestamp 1731220628
transform 1 0 816 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5588_6
timestamp 1731220628
transform 1 0 704 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5587_6
timestamp 1731220628
transform 1 0 608 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5586_6
timestamp 1731220628
transform 1 0 528 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5585_6
timestamp 1731220628
transform 1 0 648 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5584_6
timestamp 1731220628
transform 1 0 576 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5583_6
timestamp 1731220628
transform 1 0 576 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5582_6
timestamp 1731220628
transform 1 0 640 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5581_6
timestamp 1731220628
transform 1 0 624 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5580_6
timestamp 1731220628
transform 1 0 616 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5579_6
timestamp 1731220628
transform 1 0 696 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5578_6
timestamp 1731220628
transform 1 0 656 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5577_6
timestamp 1731220628
transform 1 0 600 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5576_6
timestamp 1731220628
transform 1 0 544 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5575_6
timestamp 1731220628
transform 1 0 512 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5574_6
timestamp 1731220628
transform 1 0 456 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5573_6
timestamp 1731220628
transform 1 0 376 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5572_6
timestamp 1731220628
transform 1 0 464 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5571_6
timestamp 1731220628
transform 1 0 544 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5570_6
timestamp 1731220628
transform 1 0 504 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5569_6
timestamp 1731220628
transform 1 0 432 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5568_6
timestamp 1731220628
transform 1 0 352 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5567_6
timestamp 1731220628
transform 1 0 320 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5566_6
timestamp 1731220628
transform 1 0 368 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5565_6
timestamp 1731220628
transform 1 0 408 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5564_6
timestamp 1731220628
transform 1 0 496 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5563_6
timestamp 1731220628
transform 1 0 456 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5562_6
timestamp 1731220628
transform 1 0 416 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5561_6
timestamp 1731220628
transform 1 0 376 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5560_6
timestamp 1731220628
transform 1 0 336 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5559_6
timestamp 1731220628
transform 1 0 296 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5558_6
timestamp 1731220628
transform 1 0 256 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5557_6
timestamp 1731220628
transform 1 0 216 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5556_6
timestamp 1731220628
transform 1 0 176 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5555_6
timestamp 1731220628
transform 1 0 136 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5554_6
timestamp 1731220628
transform 1 0 272 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5553_6
timestamp 1731220628
transform 1 0 224 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5552_6
timestamp 1731220628
transform 1 0 176 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5551_6
timestamp 1731220628
transform 1 0 128 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5550_6
timestamp 1731220628
transform 1 0 128 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5549_6
timestamp 1731220628
transform 1 0 192 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5548_6
timestamp 1731220628
transform 1 0 272 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5547_6
timestamp 1731220628
transform 1 0 288 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5546_6
timestamp 1731220628
transform 1 0 200 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5545_6
timestamp 1731220628
transform 1 0 128 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5544_6
timestamp 1731220628
transform 1 0 128 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5543_6
timestamp 1731220628
transform 1 0 168 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5542_6
timestamp 1731220628
transform 1 0 328 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5541_6
timestamp 1731220628
transform 1 0 264 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5540_6
timestamp 1731220628
transform 1 0 208 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5539_6
timestamp 1731220628
transform 1 0 144 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5538_6
timestamp 1731220628
transform 1 0 160 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5537_6
timestamp 1731220628
transform 1 0 160 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5536_6
timestamp 1731220628
transform 1 0 216 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5535_6
timestamp 1731220628
transform 1 0 200 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5534_6
timestamp 1731220628
transform 1 0 248 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5533_6
timestamp 1731220628
transform 1 0 280 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5532_6
timestamp 1731220628
transform 1 0 240 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5531_6
timestamp 1731220628
transform 1 0 304 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5530_6
timestamp 1731220628
transform 1 0 288 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5529_6
timestamp 1731220628
transform 1 0 200 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5528_6
timestamp 1731220628
transform 1 0 272 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5527_6
timestamp 1731220628
transform 1 0 328 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5526_6
timestamp 1731220628
transform 1 0 384 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5525_6
timestamp 1731220628
transform 1 0 392 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5524_6
timestamp 1731220628
transform 1 0 336 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5523_6
timestamp 1731220628
transform 1 0 320 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5522_6
timestamp 1731220628
transform 1 0 392 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5521_6
timestamp 1731220628
transform 1 0 456 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5520_6
timestamp 1731220628
transform 1 0 440 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5519_6
timestamp 1731220628
transform 1 0 520 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5518_6
timestamp 1731220628
transform 1 0 472 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5517_6
timestamp 1731220628
transform 1 0 552 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5516_6
timestamp 1731220628
transform 1 0 624 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5515_6
timestamp 1731220628
transform 1 0 640 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5514_6
timestamp 1731220628
transform 1 0 568 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5513_6
timestamp 1731220628
transform 1 0 496 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5512_6
timestamp 1731220628
transform 1 0 504 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5511_6
timestamp 1731220628
transform 1 0 584 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5510_6
timestamp 1731220628
transform 1 0 672 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5509_6
timestamp 1731220628
transform 1 0 768 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5508_6
timestamp 1731220628
transform 1 0 784 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5507_6
timestamp 1731220628
transform 1 0 704 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5506_6
timestamp 1731220628
transform 1 0 624 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5505_6
timestamp 1731220628
transform 1 0 544 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5504_6
timestamp 1731220628
transform 1 0 600 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5503_6
timestamp 1731220628
transform 1 0 664 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5502_6
timestamp 1731220628
transform 1 0 728 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5501_6
timestamp 1731220628
transform 1 0 792 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5500_6
timestamp 1731220628
transform 1 0 736 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5499_6
timestamp 1731220628
transform 1 0 664 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5498_6
timestamp 1731220628
transform 1 0 816 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5497_6
timestamp 1731220628
transform 1 0 856 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5496_6
timestamp 1731220628
transform 1 0 792 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5495_6
timestamp 1731220628
transform 1 0 728 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5494_6
timestamp 1731220628
transform 1 0 664 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5493_6
timestamp 1731220628
transform 1 0 688 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5492_6
timestamp 1731220628
transform 1 0 752 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5491_6
timestamp 1731220628
transform 1 0 816 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5490_6
timestamp 1731220628
transform 1 0 800 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5489_6
timestamp 1731220628
transform 1 0 744 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5488_6
timestamp 1731220628
transform 1 0 688 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5487_6
timestamp 1731220628
transform 1 0 640 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5486_6
timestamp 1731220628
transform 1 0 768 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5485_6
timestamp 1731220628
transform 1 0 728 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5484_6
timestamp 1731220628
transform 1 0 688 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5483_6
timestamp 1731220628
transform 1 0 648 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5482_6
timestamp 1731220628
transform 1 0 608 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5481_6
timestamp 1731220628
transform 1 0 568 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5480_6
timestamp 1731220628
transform 1 0 512 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5479_6
timestamp 1731220628
transform 1 0 552 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5478_6
timestamp 1731220628
transform 1 0 592 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5477_6
timestamp 1731220628
transform 1 0 624 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5476_6
timestamp 1731220628
transform 1 0 568 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5475_6
timestamp 1731220628
transform 1 0 512 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5474_6
timestamp 1731220628
transform 1 0 464 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5473_6
timestamp 1731220628
transform 1 0 424 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5472_6
timestamp 1731220628
transform 1 0 600 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5471_6
timestamp 1731220628
transform 1 0 536 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5470_6
timestamp 1731220628
transform 1 0 472 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5469_6
timestamp 1731220628
transform 1 0 416 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5468_6
timestamp 1731220628
transform 1 0 368 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5467_6
timestamp 1731220628
transform 1 0 592 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5466_6
timestamp 1731220628
transform 1 0 520 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5465_6
timestamp 1731220628
transform 1 0 448 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5464_6
timestamp 1731220628
transform 1 0 384 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5463_6
timestamp 1731220628
transform 1 0 328 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5462_6
timestamp 1731220628
transform 1 0 536 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5461_6
timestamp 1731220628
transform 1 0 472 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5460_6
timestamp 1731220628
transform 1 0 408 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5459_6
timestamp 1731220628
transform 1 0 352 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5458_6
timestamp 1731220628
transform 1 0 304 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5457_6
timestamp 1731220628
transform 1 0 256 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5456_6
timestamp 1731220628
transform 1 0 472 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5455_6
timestamp 1731220628
transform 1 0 400 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5454_6
timestamp 1731220628
transform 1 0 336 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5453_6
timestamp 1731220628
transform 1 0 272 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5452_6
timestamp 1731220628
transform 1 0 216 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5451_6
timestamp 1731220628
transform 1 0 432 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5450_6
timestamp 1731220628
transform 1 0 360 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5449_6
timestamp 1731220628
transform 1 0 296 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5448_6
timestamp 1731220628
transform 1 0 240 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5447_6
timestamp 1731220628
transform 1 0 192 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5446_6
timestamp 1731220628
transform 1 0 152 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5445_6
timestamp 1731220628
transform 1 0 192 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5444_6
timestamp 1731220628
transform 1 0 240 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5443_6
timestamp 1731220628
transform 1 0 296 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5442_6
timestamp 1731220628
transform 1 0 360 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5441_6
timestamp 1731220628
transform 1 0 424 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5440_6
timestamp 1731220628
transform 1 0 400 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5439_6
timestamp 1731220628
transform 1 0 328 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5438_6
timestamp 1731220628
transform 1 0 264 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5437_6
timestamp 1731220628
transform 1 0 216 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5436_6
timestamp 1731220628
transform 1 0 360 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5435_6
timestamp 1731220628
transform 1 0 280 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5434_6
timestamp 1731220628
transform 1 0 208 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5433_6
timestamp 1731220628
transform 1 0 144 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5432_6
timestamp 1731220628
transform 1 0 128 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5431_6
timestamp 1731220628
transform 1 0 176 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5430_6
timestamp 1731220628
transform 1 0 248 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5429_6
timestamp 1731220628
transform 1 0 272 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5428_6
timestamp 1731220628
transform 1 0 208 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5427_6
timestamp 1731220628
transform 1 0 168 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5426_6
timestamp 1731220628
transform 1 0 128 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5425_6
timestamp 1731220628
transform 1 0 128 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5424_6
timestamp 1731220628
transform 1 0 208 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5423_6
timestamp 1731220628
transform 1 0 168 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5422_6
timestamp 1731220628
transform 1 0 128 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5421_6
timestamp 1731220628
transform 1 0 128 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5420_6
timestamp 1731220628
transform 1 0 176 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5419_6
timestamp 1731220628
transform 1 0 208 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5418_6
timestamp 1731220628
transform 1 0 152 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5417_6
timestamp 1731220628
transform 1 0 152 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5416_6
timestamp 1731220628
transform 1 0 304 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5415_6
timestamp 1731220628
transform 1 0 352 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5414_6
timestamp 1731220628
transform 1 0 280 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5413_6
timestamp 1731220628
transform 1 0 224 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5412_6
timestamp 1731220628
transform 1 0 296 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5411_6
timestamp 1731220628
transform 1 0 272 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5410_6
timestamp 1731220628
transform 1 0 208 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5409_6
timestamp 1731220628
transform 1 0 392 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5408_6
timestamp 1731220628
transform 1 0 344 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5407_6
timestamp 1731220628
transform 1 0 416 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5406_6
timestamp 1731220628
transform 1 0 480 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5405_6
timestamp 1731220628
transform 1 0 528 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5404_6
timestamp 1731220628
transform 1 0 448 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5403_6
timestamp 1731220628
transform 1 0 368 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5402_6
timestamp 1731220628
transform 1 0 424 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5401_6
timestamp 1731220628
transform 1 0 504 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5400_6
timestamp 1731220628
transform 1 0 584 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5399_6
timestamp 1731220628
transform 1 0 536 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5398_6
timestamp 1731220628
transform 1 0 456 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5397_6
timestamp 1731220628
transform 1 0 376 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5396_6
timestamp 1731220628
transform 1 0 360 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5395_6
timestamp 1731220628
transform 1 0 448 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5394_6
timestamp 1731220628
transform 1 0 536 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5393_6
timestamp 1731220628
transform 1 0 512 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5392_6
timestamp 1731220628
transform 1 0 448 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5391_6
timestamp 1731220628
transform 1 0 376 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5390_6
timestamp 1731220628
transform 1 0 368 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5389_6
timestamp 1731220628
transform 1 0 440 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5388_6
timestamp 1731220628
transform 1 0 512 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5387_6
timestamp 1731220628
transform 1 0 576 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5386_6
timestamp 1731220628
transform 1 0 512 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5385_6
timestamp 1731220628
transform 1 0 448 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5384_6
timestamp 1731220628
transform 1 0 456 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5383_6
timestamp 1731220628
transform 1 0 936 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5382_6
timestamp 1731220628
transform 1 0 808 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5381_6
timestamp 1731220628
transform 1 0 728 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5380_6
timestamp 1731220628
transform 1 0 680 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5379_6
timestamp 1731220628
transform 1 0 632 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5378_6
timestamp 1731220628
transform 1 0 736 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5377_6
timestamp 1731220628
transform 1 0 848 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5376_6
timestamp 1731220628
transform 1 0 792 0 -1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5375_6
timestamp 1731220628
transform 1 0 760 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5374_6
timestamp 1731220628
transform 1 0 704 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5373_6
timestamp 1731220628
transform 1 0 936 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5372_6
timestamp 1731220628
transform 1 0 872 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5371_6
timestamp 1731220628
transform 1 0 816 0 1 656
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5370_6
timestamp 1731220628
transform 1 0 792 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5369_6
timestamp 1731220628
transform 1 0 712 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5368_6
timestamp 1731220628
transform 1 0 1024 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5367_6
timestamp 1731220628
transform 1 0 944 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5366_6
timestamp 1731220628
transform 1 0 864 0 -1 648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5365_6
timestamp 1731220628
transform 1 0 848 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5364_6
timestamp 1731220628
transform 1 0 776 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5363_6
timestamp 1731220628
transform 1 0 920 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5362_6
timestamp 1731220628
transform 1 0 992 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5361_6
timestamp 1731220628
transform 1 0 1040 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5360_6
timestamp 1731220628
transform 1 0 1040 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5359_6
timestamp 1731220628
transform 1 0 992 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5358_6
timestamp 1731220628
transform 1 0 928 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5357_6
timestamp 1731220628
transform 1 0 864 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5356_6
timestamp 1731220628
transform 1 0 800 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5355_6
timestamp 1731220628
transform 1 0 728 0 -1 532
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5354_6
timestamp 1731220628
transform 1 0 896 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5353_6
timestamp 1731220628
transform 1 0 848 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5352_6
timestamp 1731220628
transform 1 0 792 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5351_6
timestamp 1731220628
transform 1 0 736 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5350_6
timestamp 1731220628
transform 1 0 672 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5349_6
timestamp 1731220628
transform 1 0 848 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5348_6
timestamp 1731220628
transform 1 0 784 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5347_6
timestamp 1731220628
transform 1 0 720 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5346_6
timestamp 1731220628
transform 1 0 664 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5345_6
timestamp 1731220628
transform 1 0 608 0 -1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5344_6
timestamp 1731220628
transform 1 0 568 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5343_6
timestamp 1731220628
transform 1 0 744 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5342_6
timestamp 1731220628
transform 1 0 680 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5341_6
timestamp 1731220628
transform 1 0 624 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5340_6
timestamp 1731220628
transform 1 0 616 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5339_6
timestamp 1731220628
transform 1 0 680 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5338_6
timestamp 1731220628
transform 1 0 744 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5337_6
timestamp 1731220628
transform 1 0 800 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5336_6
timestamp 1731220628
transform 1 0 864 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5335_6
timestamp 1731220628
transform 1 0 928 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5334_6
timestamp 1731220628
transform 1 0 872 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5333_6
timestamp 1731220628
transform 1 0 808 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5332_6
timestamp 1731220628
transform 1 0 752 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5331_6
timestamp 1731220628
transform 1 0 696 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5330_6
timestamp 1731220628
transform 1 0 640 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5329_6
timestamp 1731220628
transform 1 0 576 0 1 216
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5328_6
timestamp 1731220628
transform 1 0 736 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5327_6
timestamp 1731220628
transform 1 0 688 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5326_6
timestamp 1731220628
transform 1 0 640 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5325_6
timestamp 1731220628
transform 1 0 592 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5324_6
timestamp 1731220628
transform 1 0 544 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5323_6
timestamp 1731220628
transform 1 0 496 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5322_6
timestamp 1731220628
transform 1 0 448 0 -1 212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5321_6
timestamp 1731220628
transform 1 0 536 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5320_6
timestamp 1731220628
transform 1 0 576 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5319_6
timestamp 1731220628
transform 1 0 616 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5318_6
timestamp 1731220628
transform 1 0 656 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5317_6
timestamp 1731220628
transform 1 0 696 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5316_6
timestamp 1731220628
transform 1 0 736 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5315_6
timestamp 1731220628
transform 1 0 776 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5314_6
timestamp 1731220628
transform 1 0 824 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5313_6
timestamp 1731220628
transform 1 0 872 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5312_6
timestamp 1731220628
transform 1 0 920 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5311_6
timestamp 1731220628
transform 1 0 960 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5310_6
timestamp 1731220628
transform 1 0 1000 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5309_6
timestamp 1731220628
transform 1 0 1040 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5308_6
timestamp 1731220628
transform 1 0 1152 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5307_6
timestamp 1731220628
transform 1 0 1152 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5306_6
timestamp 1731220628
transform 1 0 1192 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5305_6
timestamp 1731220628
transform 1 0 1256 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5304_6
timestamp 1731220628
transform 1 0 1264 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5303_6
timestamp 1731220628
transform 1 0 1200 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5302_6
timestamp 1731220628
transform 1 0 1152 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5301_6
timestamp 1731220628
transform 1 0 1160 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5300_6
timestamp 1731220628
transform 1 0 1200 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5299_6
timestamp 1731220628
transform 1 0 1240 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5298_6
timestamp 1731220628
transform 1 0 1288 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5297_6
timestamp 1731220628
transform 1 0 1384 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5296_6
timestamp 1731220628
transform 1 0 1336 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5295_6
timestamp 1731220628
transform 1 0 1320 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5294_6
timestamp 1731220628
transform 1 0 1384 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5293_6
timestamp 1731220628
transform 1 0 1392 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5292_6
timestamp 1731220628
transform 1 0 1320 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5291_6
timestamp 1731220628
transform 1 0 1264 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5290_6
timestamp 1731220628
transform 1 0 1200 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5289_6
timestamp 1731220628
transform 1 0 1328 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5288_6
timestamp 1731220628
transform 1 0 1392 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5287_6
timestamp 1731220628
transform 1 0 1448 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5286_6
timestamp 1731220628
transform 1 0 1504 0 1 84
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5285_6
timestamp 1731220628
transform 1 0 1536 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5284_6
timestamp 1731220628
transform 1 0 1464 0 -1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5283_6
timestamp 1731220628
transform 1 0 1448 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5282_6
timestamp 1731220628
transform 1 0 1520 0 1 208
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5281_6
timestamp 1731220628
transform 1 0 1488 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5280_6
timestamp 1731220628
transform 1 0 1432 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5279_6
timestamp 1731220628
transform 1 0 1616 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5278_6
timestamp 1731220628
transform 1 0 1744 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5277_6
timestamp 1731220628
transform 1 0 1672 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5276_6
timestamp 1731220628
transform 1 0 1608 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5275_6
timestamp 1731220628
transform 1 0 1544 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5274_6
timestamp 1731220628
transform 1 0 1552 0 -1 320
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5273_6
timestamp 1731220628
transform 1 0 1496 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5272_6
timestamp 1731220628
transform 1 0 1456 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5271_6
timestamp 1731220628
transform 1 0 1416 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5270_6
timestamp 1731220628
transform 1 0 1376 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5269_6
timestamp 1731220628
transform 1 0 1336 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5268_6
timestamp 1731220628
transform 1 0 1296 0 1 324
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5267_6
timestamp 1731220628
transform 1 0 1496 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5266_6
timestamp 1731220628
transform 1 0 1408 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5265_6
timestamp 1731220628
transform 1 0 1328 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5264_6
timestamp 1731220628
transform 1 0 1248 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5263_6
timestamp 1731220628
transform 1 0 1192 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5262_6
timestamp 1731220628
transform 1 0 1152 0 -1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5261_6
timestamp 1731220628
transform 1 0 1152 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5260_6
timestamp 1731220628
transform 1 0 1040 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5259_6
timestamp 1731220628
transform 1 0 1000 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5258_6
timestamp 1731220628
transform 1 0 952 0 1 428
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5257_6
timestamp 1731220628
transform 1 0 1256 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5256_6
timestamp 1731220628
transform 1 0 1376 0 1 432
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5255_6
timestamp 1731220628
transform 1 0 1280 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5254_6
timestamp 1731220628
transform 1 0 1232 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5253_6
timestamp 1731220628
transform 1 0 1184 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5252_6
timestamp 1731220628
transform 1 0 1336 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5251_6
timestamp 1731220628
transform 1 0 1400 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5250_6
timestamp 1731220628
transform 1 0 1472 0 -1 536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5249_6
timestamp 1731220628
transform 1 0 1512 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5248_6
timestamp 1731220628
transform 1 0 1456 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5247_6
timestamp 1731220628
transform 1 0 1408 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5246_6
timestamp 1731220628
transform 1 0 1368 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5245_6
timestamp 1731220628
transform 1 0 1328 0 1 540
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5244_6
timestamp 1731220628
transform 1 0 1416 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5243_6
timestamp 1731220628
transform 1 0 1360 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5242_6
timestamp 1731220628
transform 1 0 1312 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5241_6
timestamp 1731220628
transform 1 0 1272 0 -1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5240_6
timestamp 1731220628
transform 1 0 1232 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5239_6
timestamp 1731220628
transform 1 0 1280 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5238_6
timestamp 1731220628
transform 1 0 1328 0 1 644
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5237_6
timestamp 1731220628
transform 1 0 1432 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5236_6
timestamp 1731220628
transform 1 0 1352 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5235_6
timestamp 1731220628
transform 1 0 1280 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5234_6
timestamp 1731220628
transform 1 0 1232 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5233_6
timestamp 1731220628
transform 1 0 1192 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5232_6
timestamp 1731220628
transform 1 0 1152 0 -1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5231_6
timestamp 1731220628
transform 1 0 1336 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5230_6
timestamp 1731220628
transform 1 0 1232 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5229_6
timestamp 1731220628
transform 1 0 1152 0 1 752
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5228_6
timestamp 1731220628
transform 1 0 1040 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5227_6
timestamp 1731220628
transform 1 0 976 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5226_6
timestamp 1731220628
transform 1 0 888 0 1 764
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5225_6
timestamp 1731220628
transform 1 0 1040 0 -1 868
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5224_6
timestamp 1731220628
transform 1 0 1152 0 -1 864
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5223_6
timestamp 1731220628
transform 1 0 1040 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5222_6
timestamp 1731220628
transform 1 0 976 0 1 872
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5221_6
timestamp 1731220628
transform 1 0 984 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5220_6
timestamp 1731220628
transform 1 0 1040 0 -1 976
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5219_6
timestamp 1731220628
transform 1 0 1032 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5218_6
timestamp 1731220628
transform 1 0 960 0 1 980
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5217_6
timestamp 1731220628
transform 1 0 832 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5216_6
timestamp 1731220628
transform 1 0 776 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5215_6
timestamp 1731220628
transform 1 0 712 0 -1 1088
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5214_6
timestamp 1731220628
transform 1 0 872 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5213_6
timestamp 1731220628
transform 1 0 984 0 1 1096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5212_6
timestamp 1731220628
transform 1 0 952 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5211_6
timestamp 1731220628
transform 1 0 864 0 -1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5210_6
timestamp 1731220628
transform 1 0 856 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5209_6
timestamp 1731220628
transform 1 0 920 0 1 1200
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5208_6
timestamp 1731220628
transform 1 0 896 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5207_6
timestamp 1731220628
transform 1 0 976 0 -1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5206_6
timestamp 1731220628
transform 1 0 920 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5205_6
timestamp 1731220628
transform 1 0 992 0 1 1308
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5204_6
timestamp 1731220628
transform 1 0 960 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5203_6
timestamp 1731220628
transform 1 0 888 0 -1 1412
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5202_6
timestamp 1731220628
transform 1 0 864 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5201_6
timestamp 1731220628
transform 1 0 928 0 1 1416
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5200_6
timestamp 1731220628
transform 1 0 880 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5199_6
timestamp 1731220628
transform 1 0 824 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5198_6
timestamp 1731220628
transform 1 0 848 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5197_6
timestamp 1731220628
transform 1 0 784 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5196_6
timestamp 1731220628
transform 1 0 720 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5195_6
timestamp 1731220628
transform 1 0 656 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5194_6
timestamp 1731220628
transform 1 0 600 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5193_6
timestamp 1731220628
transform 1 0 536 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5192_6
timestamp 1731220628
transform 1 0 600 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5191_6
timestamp 1731220628
transform 1 0 544 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5190_6
timestamp 1731220628
transform 1 0 496 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5189_6
timestamp 1731220628
transform 1 0 448 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5188_6
timestamp 1731220628
transform 1 0 712 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5187_6
timestamp 1731220628
transform 1 0 656 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5186_6
timestamp 1731220628
transform 1 0 600 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5185_6
timestamp 1731220628
transform 1 0 664 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5184_6
timestamp 1731220628
transform 1 0 728 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5183_6
timestamp 1731220628
transform 1 0 872 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5182_6
timestamp 1731220628
transform 1 0 800 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5181_6
timestamp 1731220628
transform 1 0 744 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5180_6
timestamp 1731220628
transform 1 0 664 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5179_6
timestamp 1731220628
transform 1 0 816 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5178_6
timestamp 1731220628
transform 1 0 880 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5177_6
timestamp 1731220628
transform 1 0 1024 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5176_6
timestamp 1731220628
transform 1 0 952 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5175_6
timestamp 1731220628
transform 1 0 904 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5174_6
timestamp 1731220628
transform 1 0 832 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5173_6
timestamp 1731220628
transform 1 0 984 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5172_6
timestamp 1731220628
transform 1 0 1040 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5171_6
timestamp 1731220628
transform 1 0 1152 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5170_6
timestamp 1731220628
transform 1 0 1192 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5169_6
timestamp 1731220628
transform 1 0 1232 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5168_6
timestamp 1731220628
transform 1 0 1360 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5167_6
timestamp 1731220628
transform 1 0 1296 0 -1 1848
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5166_6
timestamp 1731220628
transform 1 0 1264 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5165_6
timestamp 1731220628
transform 1 0 1224 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5164_6
timestamp 1731220628
transform 1 0 1312 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5163_6
timestamp 1731220628
transform 1 0 1368 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5162_6
timestamp 1731220628
transform 1 0 1496 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5161_6
timestamp 1731220628
transform 1 0 1432 0 1 1852
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5160_6
timestamp 1731220628
transform 1 0 1416 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5159_6
timestamp 1731220628
transform 1 0 1352 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5158_6
timestamp 1731220628
transform 1 0 1480 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5157_6
timestamp 1731220628
transform 1 0 1552 0 -1 1956
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5156_6
timestamp 1731220628
transform 1 0 1552 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5155_6
timestamp 1731220628
transform 1 0 1448 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5154_6
timestamp 1731220628
transform 1 0 1344 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5153_6
timestamp 1731220628
transform 1 0 1392 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5152_6
timestamp 1731220628
transform 1 0 1488 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5151_6
timestamp 1731220628
transform 1 0 1432 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5150_6
timestamp 1731220628
transform 1 0 1360 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5149_6
timestamp 1731220628
transform 1 0 1512 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5148_6
timestamp 1731220628
transform 1 0 1520 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5147_6
timestamp 1731220628
transform 1 0 1448 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5146_6
timestamp 1731220628
transform 1 0 1384 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5145_6
timestamp 1731220628
transform 1 0 1328 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5144_6
timestamp 1731220628
transform 1 0 1272 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5143_6
timestamp 1731220628
transform 1 0 1232 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5142_6
timestamp 1731220628
transform 1 0 1192 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5141_6
timestamp 1731220628
transform 1 0 1152 0 -1 2176
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5140_6
timestamp 1731220628
transform 1 0 1288 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5139_6
timestamp 1731220628
transform 1 0 1232 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5138_6
timestamp 1731220628
transform 1 0 1192 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5137_6
timestamp 1731220628
transform 1 0 1152 0 1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5136_6
timestamp 1731220628
transform 1 0 1152 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5135_6
timestamp 1731220628
transform 1 0 1208 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5134_6
timestamp 1731220628
transform 1 0 1296 0 -1 2072
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5133_6
timestamp 1731220628
transform 1 0 1232 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5132_6
timestamp 1731220628
transform 1 0 1152 0 1 1968
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5131_6
timestamp 1731220628
transform 1 0 1040 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5130_6
timestamp 1731220628
transform 1 0 1000 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5129_6
timestamp 1731220628
transform 1 0 952 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5128_6
timestamp 1731220628
transform 1 0 904 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5127_6
timestamp 1731220628
transform 1 0 856 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5126_6
timestamp 1731220628
transform 1 0 808 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5125_6
timestamp 1731220628
transform 1 0 856 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5124_6
timestamp 1731220628
transform 1 0 944 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5123_6
timestamp 1731220628
transform 1 0 1032 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5122_6
timestamp 1731220628
transform 1 0 960 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5121_6
timestamp 1731220628
transform 1 0 872 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5120_6
timestamp 1731220628
transform 1 0 792 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5119_6
timestamp 1731220628
transform 1 0 896 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5118_6
timestamp 1731220628
transform 1 0 840 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5117_6
timestamp 1731220628
transform 1 0 784 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5116_6
timestamp 1731220628
transform 1 0 728 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5115_6
timestamp 1731220628
transform 1 0 680 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5114_6
timestamp 1731220628
transform 1 0 624 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5113_6
timestamp 1731220628
transform 1 0 568 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5112_6
timestamp 1731220628
transform 1 0 504 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5111_6
timestamp 1731220628
transform 1 0 552 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5110_6
timestamp 1731220628
transform 1 0 632 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5109_6
timestamp 1731220628
transform 1 0 712 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5108_6
timestamp 1731220628
transform 1 0 696 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5107_6
timestamp 1731220628
transform 1 0 776 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5106_6
timestamp 1731220628
transform 1 0 752 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5105_6
timestamp 1731220628
transform 1 0 688 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5104_6
timestamp 1731220628
transform 1 0 616 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5103_6
timestamp 1731220628
transform 1 0 752 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5102_6
timestamp 1731220628
transform 1 0 824 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5101_6
timestamp 1731220628
transform 1 0 984 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_5100_6
timestamp 1731220628
transform 1 0 904 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_599_6
timestamp 1731220628
transform 1 0 872 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_598_6
timestamp 1731220628
transform 1 0 784 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_597_6
timestamp 1731220628
transform 1 0 824 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_596_6
timestamp 1731220628
transform 1 0 752 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_595_6
timestamp 1731220628
transform 1 0 688 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_594_6
timestamp 1731220628
transform 1 0 760 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_593_6
timestamp 1731220628
transform 1 0 680 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_592_6
timestamp 1731220628
transform 1 0 600 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_591_6
timestamp 1731220628
transform 1 0 560 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_590_6
timestamp 1731220628
transform 1 0 496 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_589_6
timestamp 1731220628
transform 1 0 624 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_588_6
timestamp 1731220628
transform 1 0 608 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_587_6
timestamp 1731220628
transform 1 0 520 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_586_6
timestamp 1731220628
transform 1 0 696 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_585_6
timestamp 1731220628
transform 1 0 680 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_584_6
timestamp 1731220628
transform 1 0 600 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_583_6
timestamp 1731220628
transform 1 0 520 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_582_6
timestamp 1731220628
transform 1 0 440 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_581_6
timestamp 1731220628
transform 1 0 456 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_580_6
timestamp 1731220628
transform 1 0 536 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_579_6
timestamp 1731220628
transform 1 0 616 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_578_6
timestamp 1731220628
transform 1 0 536 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_577_6
timestamp 1731220628
transform 1 0 464 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_576_6
timestamp 1731220628
transform 1 0 400 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_575_6
timestamp 1731220628
transform 1 0 344 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_574_6
timestamp 1731220628
transform 1 0 368 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_573_6
timestamp 1731220628
transform 1 0 368 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_572_6
timestamp 1731220628
transform 1 0 296 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_571_6
timestamp 1731220628
transform 1 0 224 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_570_6
timestamp 1731220628
transform 1 0 440 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_569_6
timestamp 1731220628
transform 1 0 360 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_568_6
timestamp 1731220628
transform 1 0 288 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_567_6
timestamp 1731220628
transform 1 0 224 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_566_6
timestamp 1731220628
transform 1 0 280 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_565_6
timestamp 1731220628
transform 1 0 424 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_564_6
timestamp 1731220628
transform 1 0 352 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_563_6
timestamp 1731220628
transform 1 0 344 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_562_6
timestamp 1731220628
transform 1 0 256 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_561_6
timestamp 1731220628
transform 1 0 432 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_560_6
timestamp 1731220628
transform 1 0 520 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_559_6
timestamp 1731220628
transform 1 0 488 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_558_6
timestamp 1731220628
transform 1 0 392 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_557_6
timestamp 1731220628
transform 1 0 584 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_556_6
timestamp 1731220628
transform 1 0 528 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_555_6
timestamp 1731220628
transform 1 0 456 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_554_6
timestamp 1731220628
transform 1 0 376 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_553_6
timestamp 1731220628
transform 1 0 296 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_552_6
timestamp 1731220628
transform 1 0 296 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_551_6
timestamp 1731220628
transform 1 0 400 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_550_6
timestamp 1731220628
transform 1 0 352 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_549_6
timestamp 1731220628
transform 1 0 344 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_548_6
timestamp 1731220628
transform 1 0 408 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_547_6
timestamp 1731220628
transform 1 0 472 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_546_6
timestamp 1731220628
transform 1 0 528 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_545_6
timestamp 1731220628
transform 1 0 488 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_544_6
timestamp 1731220628
transform 1 0 448 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_543_6
timestamp 1731220628
transform 1 0 408 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_542_6
timestamp 1731220628
transform 1 0 368 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_541_6
timestamp 1731220628
transform 1 0 328 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_540_6
timestamp 1731220628
transform 1 0 288 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_539_6
timestamp 1731220628
transform 1 0 248 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_538_6
timestamp 1731220628
transform 1 0 208 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_537_6
timestamp 1731220628
transform 1 0 168 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_536_6
timestamp 1731220628
transform 1 0 128 0 -1 1528
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_535_6
timestamp 1731220628
transform 1 0 136 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_534_6
timestamp 1731220628
transform 1 0 176 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_533_6
timestamp 1731220628
transform 1 0 224 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_532_6
timestamp 1731220628
transform 1 0 280 0 1 1536
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_531_6
timestamp 1731220628
transform 1 0 248 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_530_6
timestamp 1731220628
transform 1 0 208 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_529_6
timestamp 1731220628
transform 1 0 168 0 -1 1648
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_528_6
timestamp 1731220628
transform 1 0 144 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_527_6
timestamp 1731220628
transform 1 0 216 0 1 1652
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_526_6
timestamp 1731220628
transform 1 0 288 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_525_6
timestamp 1731220628
transform 1 0 192 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_524_6
timestamp 1731220628
transform 1 0 128 0 -1 1760
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_523_6
timestamp 1731220628
transform 1 0 176 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_522_6
timestamp 1731220628
transform 1 0 128 0 1 1768
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_521_6
timestamp 1731220628
transform 1 0 128 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_520_6
timestamp 1731220628
transform 1 0 216 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_519_6
timestamp 1731220628
transform 1 0 168 0 -1 1876
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_518_6
timestamp 1731220628
transform 1 0 128 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_517_6
timestamp 1731220628
transform 1 0 168 0 1 1880
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_516_6
timestamp 1731220628
transform 1 0 152 0 -1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_515_6
timestamp 1731220628
transform 1 0 176 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_514_6
timestamp 1731220628
transform 1 0 272 0 1 1988
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_513_6
timestamp 1731220628
transform 1 0 296 0 -1 2096
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_512_6
timestamp 1731220628
transform 1 0 480 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_511_6
timestamp 1731220628
transform 1 0 416 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_510_6
timestamp 1731220628
transform 1 0 352 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_59_6
timestamp 1731220628
transform 1 0 304 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_58_6
timestamp 1731220628
transform 1 0 264 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_57_6
timestamp 1731220628
transform 1 0 224 0 1 2100
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_56_6
timestamp 1731220628
transform 1 0 440 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_55_6
timestamp 1731220628
transform 1 0 376 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_54_6
timestamp 1731220628
transform 1 0 312 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_53_6
timestamp 1731220628
transform 1 0 248 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_52_6
timestamp 1731220628
transform 1 0 208 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_51_6
timestamp 1731220628
transform 1 0 168 0 -1 2212
box 4 6 36 48
use _0_0std_0_0cells_0_0NOR2X1  tst_50_6
timestamp 1731220628
transform 1 0 128 0 -1 2212
box 4 6 36 48
<< end >>
