magic
tech TSMC180
timestamp 1734144001
<< ndiffusion >>
rect 6 11 12 12
rect 6 9 7 11
rect 9 9 12 11
rect 14 11 20 12
rect 14 9 17 11
rect 19 9 20 11
rect 6 8 10 9
rect 16 8 20 9
<< ndcontact >>
rect 7 9 9 11
rect 17 9 19 11
<< ntransistor >>
rect 12 9 14 12
<< pdiffusion >>
rect 6 31 10 32
rect 16 31 20 32
rect 6 29 7 31
rect 9 29 12 31
rect 6 28 12 29
rect 14 29 17 31
rect 19 29 20 31
rect 14 28 20 29
<< pdcontact >>
rect 7 29 9 31
rect 17 29 19 31
<< ptransistor >>
rect 12 28 14 31
<< polysilicon >>
rect 12 31 14 34
rect 12 12 14 28
rect 12 6 14 9
rect 12 5 20 6
rect 12 3 17 5
rect 19 3 20 5
rect 12 2 20 3
<< polycontact >>
rect 17 3 19 5
<< m1 >>
rect 6 32 9 40
rect 6 31 10 32
rect 6 29 7 31
rect 9 29 10 31
rect 6 28 10 29
rect 16 31 20 32
rect 24 31 27 40
rect 16 29 17 31
rect 19 29 27 31
rect 16 28 27 29
rect 6 12 9 13
rect 6 11 10 12
rect 6 9 7 11
rect 9 9 10 11
rect 6 8 10 9
rect 16 11 20 12
rect 16 9 17 11
rect 19 9 20 11
rect 16 5 20 9
rect 16 3 17 5
rect 19 3 20 5
rect 16 2 20 3
<< labels >>
rlabel m1 s 19 29 27 31 6 Y
port 1 nsew signal output
rlabel m1 s 17 29 19 31 6 Y
port 1 nsew signal output
rlabel m1 s 16 29 17 31 6 Y
port 1 nsew signal output
rlabel m1 s 24 31 27 40 6 Y
port 1 nsew signal output
rlabel m1 s 16 28 27 29 6 Y
port 1 nsew signal output
rlabel m1 s 16 31 20 32 6 Y
port 1 nsew signal output
rlabel m1 s 9 29 10 31 6 Vdd
port 2 nsew power input
rlabel m1 s 7 29 9 31 6 Vdd
port 2 nsew power input
rlabel m1 s 6 28 10 29 6 Vdd
port 2 nsew power input
rlabel m1 s 6 29 7 31 6 Vdd
port 2 nsew power input
rlabel m1 s 6 31 10 32 6 Vdd
port 2 nsew power input
rlabel m1 s 6 32 9 40 6 Vdd
port 2 nsew power input
rlabel m1 s 9 9 10 11 6 GND
port 3 nsew ground input
rlabel m1 s 7 9 9 11 6 GND
port 3 nsew ground input
rlabel m1 s 6 8 10 9 6 GND
port 3 nsew ground input
rlabel m1 s 6 9 7 11 6 GND
port 3 nsew ground input
rlabel m1 s 6 11 10 12 6 GND
port 3 nsew ground input
rlabel m1 s 6 12 9 13 6 GND
port 3 nsew ground input
rlabel space 0 0 30 50 1 prboundary
rlabel ndiffusion 15 10 15 10 3 x
rlabel ndiffusion 15 12 15 12 3 x
rlabel ndiffusion 17 9 17 9 3 x
rlabel ntransistor 13 10 13 10 3 x
rlabel pdiffusion 15 29 15 29 3 Y
rlabel pdiffusion 15 30 15 30 3 Y
rlabel polysilicon 13 32 13 32 3 x
rlabel polysilicon 13 3 13 3 3 x
rlabel polysilicon 13 4 13 4 3 x
rlabel polysilicon 13 6 13 6 3 x
rlabel polysilicon 13 7 13 7 3 x
rlabel polysilicon 13 13 13 13 3 x
rlabel ptransistor 13 29 13 29 3 x
rlabel m1 20 10 20 10 3 x
rlabel m1 20 30 20 30 3 Y
port 1 e default output
rlabel ndcontact 18 10 18 10 3 x
rlabel pdcontact 18 30 18 30 3 Y
port 1 e default output
rlabel m1 20 4 20 4 3 x
rlabel m1 17 10 17 10 3 x
rlabel m1 17 30 17 30 3 Y
port 1 e default output
rlabel m1 25 32 25 32 3 Y
port 1 e
rlabel polycontact 18 4 18 4 3 x
rlabel m1 17 3 17 3 3 x
rlabel m1 17 4 17 4 3 x
rlabel m1 17 6 17 6 3 x
rlabel m1 10 10 10 10 3 GND
rlabel m1 17 12 17 12 3 x
rlabel m1 17 29 17 29 3 Y
port 1 e
rlabel m1 10 30 10 30 3 Vdd
rlabel m1 17 32 17 32 3 Y
port 1 e
rlabel ndcontact 8 10 8 10 3 GND
rlabel pdcontact 8 30 8 30 3 Vdd
rlabel m1 7 9 7 9 3 GND
rlabel m1 7 10 7 10 3 GND
rlabel m1 7 12 7 12 3 GND
rlabel m1 7 13 7 13 3 GND
rlabel m1 7 29 7 29 3 Vdd
rlabel m1 7 30 7 30 3 Vdd
rlabel m1 7 32 7 32 3 Vdd
rlabel m1 7 33 7 33 3 Vdd
<< properties >>
string FIXED_BBOX 0 0 30 50
string LEFclass CORE
string LEFsite CoreSite
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
