magic
tech sky130l
timestamp 1731220403
<< m1 >>
rect 424 2535 428 2571
rect 480 2535 484 2571
rect 816 2535 820 2571
rect 872 2535 876 2571
rect 928 2535 932 2571
rect 2152 2531 2156 2567
rect 2272 2531 2276 2567
rect 512 2483 516 2515
rect 576 2487 580 2515
rect 904 2451 908 2515
rect 984 2475 988 2531
rect 512 2415 516 2451
rect 592 2415 596 2451
rect 968 2335 972 2395
rect 1040 2363 1044 2395
rect 1784 2359 1788 2391
rect 2096 2239 2100 2271
rect 2464 2163 2468 2199
rect 480 2123 484 2155
rect 1000 2123 1004 2155
rect 1216 2123 1220 2155
rect 2384 2115 2388 2147
rect 1800 2051 1804 2087
rect 440 1995 444 2027
rect 496 1995 500 2027
rect 776 1995 780 2027
rect 832 1995 836 2027
rect 888 1995 892 2027
rect 944 1995 948 2027
rect 1000 1995 1004 2027
rect 2032 2003 2036 2035
rect 2472 2003 2476 2035
rect 544 1927 548 1963
rect 2080 1887 2084 1919
rect 1440 1819 1444 1855
rect 1504 1819 1508 1855
rect 1600 1819 1604 1855
rect 680 1723 684 1787
rect 1056 1755 1060 1787
rect 1760 1771 1764 1803
rect 688 1687 692 1723
rect 768 1687 772 1723
rect 1064 1687 1068 1747
rect 1480 1707 1484 1743
rect 1560 1707 1564 1743
rect 1656 1707 1660 1743
rect 1864 1707 1868 1743
rect 424 1635 428 1667
rect 912 1635 916 1667
rect 968 1555 972 1587
rect 1104 1555 1108 1591
rect 1616 1571 1620 1607
rect 1672 1571 1676 1607
rect 1728 1571 1732 1607
rect 1792 1571 1796 1607
rect 1704 1519 1708 1551
rect 2192 1519 2196 1567
rect 528 1439 532 1475
rect 1744 1391 1748 1423
rect 2328 1391 2332 1423
rect 2416 1395 2420 1423
rect 552 1323 556 1359
rect 1848 1319 1852 1355
rect 1736 1263 1740 1303
rect 1864 1203 1868 1239
rect 184 1147 188 1179
rect 536 1147 540 1179
rect 952 1111 956 1179
rect 1728 1079 1732 1115
rect 1936 1079 1940 1139
rect 2384 1079 2388 1115
rect 336 1023 340 1055
rect 1384 1023 1388 1059
rect 1440 1023 1444 1063
rect 1016 955 1020 991
rect 1080 955 1084 991
rect 1144 955 1148 991
rect 1200 955 1204 991
rect 1256 955 1260 991
rect 1864 947 1868 1019
rect 616 903 620 935
rect 1680 863 1684 923
rect 1736 891 1740 923
rect 864 783 868 815
rect 944 787 948 815
rect 1656 771 1660 803
rect 1960 739 1964 803
rect 2360 771 2364 803
rect 304 663 308 691
rect 1536 651 1540 683
rect 1640 651 1644 683
rect 1440 587 1444 623
rect 1952 587 1956 623
rect 224 539 228 567
rect 296 535 300 567
rect 472 499 476 567
rect 1984 531 1988 563
rect 2512 467 2516 503
rect 808 343 812 379
rect 1128 343 1132 379
rect 1216 343 1220 379
rect 792 295 796 323
rect 1992 227 1996 283
rect 2456 227 2460 259
rect 384 175 388 207
rect 2488 179 2492 211
<< m2c >>
rect 528 2631 532 2635
rect 584 2631 588 2635
rect 640 2631 644 2635
rect 696 2631 700 2635
rect 752 2631 756 2635
rect 1528 2627 1532 2631
rect 1584 2627 1588 2631
rect 1640 2627 1644 2631
rect 1696 2627 1700 2631
rect 1752 2627 1756 2631
rect 1808 2627 1812 2631
rect 1864 2627 1868 2631
rect 1920 2627 1924 2631
rect 1976 2627 1980 2631
rect 2032 2627 2036 2631
rect 2088 2627 2092 2631
rect 2144 2627 2148 2631
rect 568 2595 572 2599
rect 624 2595 628 2599
rect 680 2595 684 2599
rect 736 2595 740 2599
rect 792 2595 796 2599
rect 1568 2591 1572 2595
rect 1624 2591 1628 2595
rect 1680 2591 1684 2595
rect 1736 2591 1740 2595
rect 1792 2591 1796 2595
rect 1848 2591 1852 2595
rect 1904 2591 1908 2595
rect 1960 2591 1964 2595
rect 2016 2591 2020 2595
rect 2072 2591 2076 2595
rect 2128 2591 2132 2595
rect 2184 2591 2188 2595
rect 424 2571 428 2575
rect 480 2571 484 2575
rect 816 2571 820 2575
rect 872 2571 876 2575
rect 928 2571 932 2575
rect 248 2567 252 2571
rect 304 2567 308 2571
rect 360 2567 364 2571
rect 416 2567 420 2571
rect 472 2567 476 2571
rect 528 2567 532 2571
rect 584 2567 588 2571
rect 640 2567 644 2571
rect 696 2567 700 2571
rect 752 2567 756 2571
rect 808 2567 812 2571
rect 864 2567 868 2571
rect 920 2567 924 2571
rect 976 2567 980 2571
rect 1032 2567 1036 2571
rect 1088 2567 1092 2571
rect 1144 2567 1148 2571
rect 2152 2567 2156 2571
rect 2272 2567 2276 2571
rect 1472 2563 1476 2567
rect 1576 2563 1580 2567
rect 1688 2563 1692 2567
rect 1800 2563 1804 2567
rect 1912 2563 1916 2567
rect 2024 2563 2028 2567
rect 2144 2563 2148 2567
rect 208 2531 212 2535
rect 264 2531 268 2535
rect 320 2531 324 2535
rect 376 2531 380 2535
rect 424 2531 428 2535
rect 432 2531 436 2535
rect 480 2531 484 2535
rect 488 2531 492 2535
rect 544 2531 548 2535
rect 600 2531 604 2535
rect 656 2531 660 2535
rect 712 2531 716 2535
rect 768 2531 772 2535
rect 816 2531 820 2535
rect 824 2531 828 2535
rect 872 2531 876 2535
rect 880 2531 884 2535
rect 928 2531 932 2535
rect 936 2531 940 2535
rect 984 2531 988 2535
rect 992 2531 996 2535
rect 1048 2531 1052 2535
rect 1104 2531 1108 2535
rect 2264 2563 2268 2567
rect 2384 2563 2388 2567
rect 344 2517 348 2521
rect 400 2515 404 2519
rect 464 2515 468 2519
rect 512 2515 516 2519
rect 528 2515 532 2519
rect 576 2515 580 2519
rect 592 2515 596 2519
rect 656 2515 660 2519
rect 720 2515 724 2519
rect 784 2515 788 2519
rect 848 2515 852 2519
rect 904 2515 908 2519
rect 920 2515 924 2519
rect 384 2479 388 2483
rect 440 2479 444 2483
rect 504 2479 508 2483
rect 512 2479 516 2483
rect 568 2481 572 2485
rect 576 2483 580 2487
rect 632 2479 636 2483
rect 696 2479 700 2483
rect 760 2479 764 2483
rect 824 2479 828 2483
rect 888 2479 892 2483
rect 512 2451 516 2455
rect 592 2451 596 2455
rect 960 2481 964 2485
rect 1432 2527 1436 2531
rect 1536 2527 1540 2531
rect 1648 2527 1652 2531
rect 1760 2527 1764 2531
rect 1872 2527 1876 2531
rect 1984 2527 1988 2531
rect 2104 2527 2108 2531
rect 2152 2527 2156 2531
rect 2224 2527 2228 2531
rect 2272 2527 2276 2531
rect 2344 2527 2348 2531
rect 992 2515 996 2519
rect 1528 2507 1532 2511
rect 1608 2507 1612 2511
rect 1696 2507 1700 2511
rect 1784 2507 1788 2511
rect 1880 2507 1884 2511
rect 1976 2507 1980 2511
rect 2072 2507 2076 2511
rect 2168 2507 2172 2511
rect 2272 2507 2276 2511
rect 2376 2507 2380 2511
rect 1032 2479 1036 2483
rect 984 2471 988 2475
rect 1568 2471 1572 2475
rect 1648 2471 1652 2475
rect 1736 2471 1740 2475
rect 1824 2471 1828 2475
rect 1920 2471 1924 2475
rect 2016 2471 2020 2475
rect 2112 2471 2116 2475
rect 2208 2471 2212 2475
rect 2312 2471 2316 2475
rect 2416 2471 2420 2475
rect 304 2447 308 2451
rect 368 2447 372 2451
rect 432 2447 436 2451
rect 504 2447 508 2451
rect 584 2447 588 2451
rect 664 2447 668 2451
rect 744 2447 748 2451
rect 816 2447 820 2451
rect 896 2447 900 2451
rect 904 2447 908 2451
rect 976 2447 980 2451
rect 1056 2447 1060 2451
rect 1680 2443 1684 2447
rect 1736 2443 1740 2447
rect 1800 2443 1804 2447
rect 1872 2443 1876 2447
rect 1944 2443 1948 2447
rect 2024 2443 2028 2447
rect 2112 2443 2116 2447
rect 2200 2443 2204 2447
rect 2296 2443 2300 2447
rect 2392 2443 2396 2447
rect 2560 2443 2564 2447
rect 264 2411 268 2415
rect 328 2411 332 2415
rect 392 2411 396 2415
rect 464 2411 468 2415
rect 512 2411 516 2415
rect 544 2411 548 2415
rect 592 2411 596 2415
rect 624 2411 628 2415
rect 704 2411 708 2415
rect 776 2411 780 2415
rect 856 2411 860 2415
rect 936 2411 940 2415
rect 1016 2411 1020 2415
rect 1640 2407 1644 2411
rect 1696 2407 1700 2411
rect 1760 2407 1764 2411
rect 1832 2407 1836 2411
rect 1904 2407 1908 2411
rect 1984 2407 1988 2411
rect 2072 2407 2076 2411
rect 2160 2407 2164 2411
rect 2256 2407 2260 2411
rect 2352 2407 2356 2411
rect 2448 2407 2452 2411
rect 2520 2407 2524 2411
rect 224 2395 228 2399
rect 312 2395 316 2399
rect 408 2395 412 2399
rect 504 2395 508 2399
rect 608 2395 612 2399
rect 704 2395 708 2399
rect 800 2395 804 2399
rect 896 2395 900 2399
rect 968 2395 972 2399
rect 992 2395 996 2399
rect 1040 2395 1044 2399
rect 1088 2395 1092 2399
rect 264 2359 268 2363
rect 352 2359 356 2363
rect 448 2359 452 2363
rect 544 2359 548 2363
rect 648 2359 652 2363
rect 744 2359 748 2363
rect 840 2359 844 2363
rect 936 2359 940 2363
rect 1432 2391 1436 2395
rect 1536 2391 1540 2395
rect 1640 2391 1644 2395
rect 1736 2391 1740 2395
rect 1784 2391 1788 2395
rect 1832 2391 1836 2395
rect 1920 2391 1924 2395
rect 2016 2391 2020 2395
rect 2112 2391 2116 2395
rect 2208 2391 2212 2395
rect 2312 2391 2316 2395
rect 2424 2391 2428 2395
rect 2520 2391 2524 2395
rect 1032 2359 1036 2363
rect 1040 2359 1044 2363
rect 1128 2359 1132 2363
rect 1472 2355 1476 2359
rect 1576 2355 1580 2359
rect 1680 2355 1684 2359
rect 1776 2355 1780 2359
rect 1784 2355 1788 2359
rect 1872 2355 1876 2359
rect 1960 2355 1964 2359
rect 2056 2355 2060 2359
rect 2152 2355 2156 2359
rect 2248 2355 2252 2359
rect 2352 2355 2356 2359
rect 2464 2355 2468 2359
rect 2560 2355 2564 2359
rect 192 2331 196 2335
rect 296 2331 300 2335
rect 408 2331 412 2335
rect 520 2331 524 2335
rect 632 2331 636 2335
rect 744 2331 748 2335
rect 848 2331 852 2335
rect 944 2331 948 2335
rect 968 2331 972 2335
rect 1040 2331 1044 2335
rect 1136 2331 1140 2335
rect 1232 2331 1236 2335
rect 1432 2327 1436 2331
rect 1488 2327 1492 2331
rect 1544 2327 1548 2331
rect 1600 2327 1604 2331
rect 1672 2327 1676 2331
rect 1760 2327 1764 2331
rect 1856 2327 1860 2331
rect 1976 2327 1980 2331
rect 2112 2327 2116 2331
rect 2256 2327 2260 2331
rect 2416 2327 2420 2331
rect 2560 2327 2564 2331
rect 152 2295 156 2299
rect 256 2295 260 2299
rect 368 2295 372 2299
rect 480 2295 484 2299
rect 592 2295 596 2299
rect 704 2295 708 2299
rect 808 2295 812 2299
rect 904 2295 908 2299
rect 1000 2295 1004 2299
rect 1096 2295 1100 2299
rect 1192 2295 1196 2299
rect 1392 2291 1396 2295
rect 1448 2291 1452 2295
rect 1504 2291 1508 2295
rect 1560 2291 1564 2295
rect 1632 2291 1636 2295
rect 1720 2291 1724 2295
rect 1816 2291 1820 2295
rect 1936 2291 1940 2295
rect 2072 2291 2076 2295
rect 2216 2291 2220 2295
rect 2376 2291 2380 2295
rect 2520 2291 2524 2295
rect 136 2279 140 2283
rect 224 2279 228 2283
rect 352 2279 356 2283
rect 488 2279 492 2283
rect 616 2279 620 2283
rect 744 2279 748 2283
rect 864 2279 868 2283
rect 976 2279 980 2283
rect 1080 2279 1084 2283
rect 1184 2279 1188 2283
rect 1264 2279 1268 2283
rect 1392 2271 1396 2275
rect 1472 2271 1476 2275
rect 1592 2271 1596 2275
rect 1712 2271 1716 2275
rect 1832 2271 1836 2275
rect 1944 2271 1948 2275
rect 2048 2271 2052 2275
rect 2096 2271 2100 2275
rect 2144 2271 2148 2275
rect 2232 2271 2236 2275
rect 2312 2271 2316 2275
rect 2384 2271 2388 2275
rect 2464 2271 2468 2275
rect 2520 2271 2524 2275
rect 176 2243 180 2247
rect 264 2243 268 2247
rect 392 2245 396 2249
rect 528 2243 532 2247
rect 656 2243 660 2247
rect 784 2243 788 2247
rect 904 2243 908 2247
rect 1016 2243 1020 2247
rect 1120 2243 1124 2247
rect 1224 2243 1228 2247
rect 1304 2243 1308 2247
rect 1432 2235 1436 2239
rect 1512 2235 1516 2239
rect 1632 2235 1636 2239
rect 1752 2235 1756 2239
rect 1872 2235 1876 2239
rect 1984 2235 1988 2239
rect 2088 2235 2092 2239
rect 2096 2235 2100 2239
rect 2184 2235 2188 2239
rect 2272 2235 2276 2239
rect 2352 2235 2356 2239
rect 2424 2235 2428 2239
rect 2504 2235 2508 2239
rect 2560 2235 2564 2239
rect 176 2207 180 2211
rect 264 2207 268 2211
rect 392 2207 396 2211
rect 528 2207 532 2211
rect 656 2207 660 2211
rect 784 2207 788 2211
rect 904 2207 908 2211
rect 1016 2207 1020 2211
rect 1120 2207 1124 2211
rect 1224 2207 1228 2211
rect 1304 2207 1308 2211
rect 2464 2199 2468 2203
rect 1488 2195 1492 2199
rect 1568 2195 1572 2199
rect 1664 2195 1668 2199
rect 1776 2195 1780 2199
rect 1896 2195 1900 2199
rect 2016 2195 2020 2199
rect 2128 2195 2132 2199
rect 2240 2195 2244 2199
rect 2344 2195 2348 2199
rect 2456 2195 2460 2199
rect 136 2171 140 2175
rect 224 2171 228 2175
rect 352 2171 356 2175
rect 488 2171 492 2175
rect 616 2171 620 2175
rect 744 2171 748 2175
rect 864 2171 868 2175
rect 976 2171 980 2175
rect 1080 2171 1084 2175
rect 1184 2171 1188 2175
rect 1264 2171 1268 2175
rect 2560 2195 2564 2199
rect 1448 2159 1452 2163
rect 1528 2159 1532 2163
rect 1624 2159 1628 2163
rect 1736 2159 1740 2163
rect 1856 2159 1860 2163
rect 1976 2159 1980 2163
rect 2088 2159 2092 2163
rect 2200 2159 2204 2163
rect 2304 2159 2308 2163
rect 2416 2159 2420 2163
rect 2464 2159 2468 2163
rect 2520 2159 2524 2163
rect 136 2155 140 2159
rect 192 2155 196 2159
rect 288 2155 292 2159
rect 400 2155 404 2159
rect 480 2155 484 2159
rect 520 2155 524 2159
rect 640 2155 644 2159
rect 752 2155 756 2159
rect 856 2155 860 2159
rect 952 2155 956 2159
rect 1000 2155 1004 2159
rect 1048 2155 1052 2159
rect 1144 2155 1148 2159
rect 1216 2155 1220 2159
rect 1248 2155 1252 2159
rect 1512 2147 1516 2151
rect 1608 2147 1612 2151
rect 1712 2147 1716 2151
rect 1816 2147 1820 2151
rect 1928 2147 1932 2151
rect 2032 2147 2036 2151
rect 2136 2147 2140 2151
rect 2240 2147 2244 2151
rect 2336 2147 2340 2151
rect 2384 2147 2388 2151
rect 2440 2147 2444 2151
rect 2520 2147 2524 2151
rect 176 2119 180 2123
rect 232 2119 236 2123
rect 328 2119 332 2123
rect 440 2119 444 2123
rect 480 2119 484 2123
rect 560 2119 564 2123
rect 680 2119 684 2123
rect 792 2119 796 2123
rect 896 2119 900 2123
rect 992 2119 996 2123
rect 1000 2119 1004 2123
rect 1088 2119 1092 2123
rect 1184 2119 1188 2123
rect 1216 2119 1220 2123
rect 1288 2119 1292 2123
rect 1552 2111 1556 2115
rect 1648 2111 1652 2115
rect 1752 2111 1756 2115
rect 1856 2111 1860 2115
rect 1968 2111 1972 2115
rect 2072 2111 2076 2115
rect 2176 2111 2180 2115
rect 2280 2111 2284 2115
rect 2376 2111 2380 2115
rect 2384 2111 2388 2115
rect 2480 2111 2484 2115
rect 2560 2111 2564 2115
rect 1800 2087 1804 2091
rect 296 2083 300 2087
rect 360 2083 364 2087
rect 432 2083 436 2087
rect 512 2083 516 2087
rect 600 2083 604 2087
rect 688 2083 692 2087
rect 768 2083 772 2087
rect 848 2083 852 2087
rect 920 2083 924 2087
rect 1000 2083 1004 2087
rect 1080 2083 1084 2087
rect 1160 2083 1164 2087
rect 1464 2083 1468 2087
rect 1568 2083 1572 2087
rect 1680 2083 1684 2087
rect 1792 2083 1796 2087
rect 1896 2083 1900 2087
rect 2000 2083 2004 2087
rect 2104 2083 2108 2087
rect 2208 2083 2212 2087
rect 2304 2083 2308 2087
rect 2392 2083 2396 2087
rect 2488 2083 2492 2087
rect 2560 2083 2564 2087
rect 256 2047 260 2051
rect 320 2047 324 2051
rect 392 2047 396 2051
rect 472 2047 476 2051
rect 560 2047 564 2051
rect 648 2047 652 2051
rect 728 2047 732 2051
rect 808 2047 812 2051
rect 880 2047 884 2051
rect 960 2047 964 2051
rect 1040 2047 1044 2051
rect 1120 2047 1124 2051
rect 1424 2047 1428 2051
rect 1528 2047 1532 2051
rect 1640 2047 1644 2051
rect 1752 2047 1756 2051
rect 1800 2047 1804 2051
rect 1856 2047 1860 2051
rect 1960 2047 1964 2051
rect 2064 2047 2068 2051
rect 2168 2047 2172 2051
rect 2264 2047 2268 2051
rect 2352 2047 2356 2051
rect 2448 2047 2452 2051
rect 2520 2047 2524 2051
rect 1392 2035 1396 2039
rect 1480 2035 1484 2039
rect 1584 2035 1588 2039
rect 1688 2035 1692 2039
rect 1784 2035 1788 2039
rect 1880 2035 1884 2039
rect 1984 2035 1988 2039
rect 2032 2035 2036 2039
rect 2088 2035 2092 2039
rect 2192 2035 2196 2039
rect 2304 2035 2308 2039
rect 2424 2035 2428 2039
rect 2472 2035 2476 2039
rect 2520 2035 2524 2039
rect 392 2027 396 2031
rect 440 2027 444 2031
rect 448 2027 452 2031
rect 496 2027 500 2031
rect 504 2027 508 2031
rect 560 2027 564 2031
rect 616 2027 620 2031
rect 672 2027 676 2031
rect 728 2027 732 2031
rect 776 2027 780 2031
rect 784 2027 788 2031
rect 832 2027 836 2031
rect 840 2027 844 2031
rect 888 2027 892 2031
rect 896 2027 900 2031
rect 944 2027 948 2031
rect 952 2027 956 2031
rect 1000 2027 1004 2031
rect 1008 2027 1012 2031
rect 1432 1999 1436 2003
rect 1520 1999 1524 2003
rect 1624 1999 1628 2003
rect 1728 1999 1732 2003
rect 1824 1999 1828 2003
rect 1920 1999 1924 2003
rect 2024 1999 2028 2003
rect 2032 1999 2036 2003
rect 2128 1999 2132 2003
rect 2232 1999 2236 2003
rect 2344 1999 2348 2003
rect 2464 1999 2468 2003
rect 2472 1999 2476 2003
rect 2560 1999 2564 2003
rect 432 1991 436 1995
rect 440 1991 444 1995
rect 488 1991 492 1995
rect 496 1991 500 1995
rect 544 1991 548 1995
rect 600 1991 604 1995
rect 656 1991 660 1995
rect 712 1991 716 1995
rect 768 1991 772 1995
rect 776 1991 780 1995
rect 824 1991 828 1995
rect 832 1991 836 1995
rect 880 1991 884 1995
rect 888 1991 892 1995
rect 936 1991 940 1995
rect 944 1991 948 1995
rect 992 1991 996 1995
rect 1000 1991 1004 1995
rect 1048 1991 1052 1995
rect 1432 1971 1436 1975
rect 1512 1971 1516 1975
rect 1616 1971 1620 1975
rect 1712 1971 1716 1975
rect 1800 1971 1804 1975
rect 1880 1971 1884 1975
rect 1960 1971 1964 1975
rect 2040 1971 2044 1975
rect 2120 1971 2124 1975
rect 544 1963 548 1967
rect 368 1959 372 1963
rect 424 1959 428 1963
rect 480 1959 484 1963
rect 536 1959 540 1963
rect 600 1959 604 1963
rect 680 1959 684 1963
rect 776 1959 780 1963
rect 896 1959 900 1963
rect 1032 1959 1036 1963
rect 1176 1959 1180 1963
rect 1304 1959 1308 1963
rect 1392 1935 1396 1939
rect 1472 1935 1476 1939
rect 1576 1935 1580 1939
rect 1672 1935 1676 1939
rect 1760 1935 1764 1939
rect 1840 1935 1844 1939
rect 1920 1935 1924 1939
rect 2000 1935 2004 1939
rect 2080 1935 2084 1939
rect 328 1923 332 1927
rect 384 1923 388 1927
rect 440 1923 444 1927
rect 496 1923 500 1927
rect 544 1923 548 1927
rect 560 1923 564 1927
rect 640 1923 644 1927
rect 736 1923 740 1927
rect 856 1923 860 1927
rect 992 1923 996 1927
rect 1136 1923 1140 1927
rect 1264 1923 1268 1927
rect 1696 1921 1700 1925
rect 1752 1919 1756 1923
rect 1808 1919 1812 1923
rect 1864 1919 1868 1923
rect 1920 1919 1924 1923
rect 1976 1919 1980 1923
rect 2032 1919 2036 1923
rect 2080 1919 2084 1923
rect 2096 1919 2100 1923
rect 136 1911 140 1915
rect 208 1911 212 1915
rect 304 1911 308 1915
rect 408 1911 412 1915
rect 520 1911 524 1915
rect 632 1911 636 1915
rect 744 1911 748 1915
rect 856 1911 860 1915
rect 960 1911 964 1915
rect 1064 1911 1068 1915
rect 1176 1911 1180 1915
rect 1264 1911 1268 1915
rect 1736 1883 1740 1887
rect 1792 1883 1796 1887
rect 1848 1883 1852 1887
rect 1904 1883 1908 1887
rect 1960 1883 1964 1887
rect 2016 1883 2020 1887
rect 2072 1883 2076 1887
rect 2080 1883 2084 1887
rect 2136 1883 2140 1887
rect 176 1875 180 1879
rect 248 1875 252 1879
rect 344 1875 348 1879
rect 448 1875 452 1879
rect 560 1875 564 1879
rect 672 1875 676 1879
rect 784 1875 788 1879
rect 896 1875 900 1879
rect 1000 1875 1004 1879
rect 1104 1875 1108 1879
rect 1216 1875 1220 1879
rect 1304 1875 1308 1879
rect 1440 1855 1444 1859
rect 1504 1855 1508 1859
rect 1600 1855 1604 1859
rect 1432 1851 1436 1855
rect 176 1839 180 1843
rect 232 1839 236 1843
rect 296 1839 300 1843
rect 384 1839 388 1843
rect 472 1839 476 1843
rect 568 1839 572 1843
rect 656 1839 660 1843
rect 744 1839 748 1843
rect 824 1839 828 1843
rect 904 1839 908 1843
rect 984 1839 988 1843
rect 1072 1839 1076 1843
rect 1496 1851 1500 1855
rect 1592 1851 1596 1855
rect 1688 1851 1692 1855
rect 1776 1851 1780 1855
rect 1864 1851 1868 1855
rect 1952 1851 1956 1855
rect 2040 1851 2044 1855
rect 2128 1851 2132 1855
rect 2216 1851 2220 1855
rect 1392 1815 1396 1819
rect 1440 1815 1444 1819
rect 1456 1815 1460 1819
rect 1504 1815 1508 1819
rect 1552 1815 1556 1819
rect 1600 1815 1604 1819
rect 1648 1815 1652 1819
rect 1736 1815 1740 1819
rect 1824 1815 1828 1819
rect 1912 1815 1916 1819
rect 2000 1815 2004 1819
rect 2088 1815 2092 1819
rect 2176 1815 2180 1819
rect 136 1803 140 1807
rect 192 1803 196 1807
rect 256 1803 260 1807
rect 344 1803 348 1807
rect 432 1803 436 1807
rect 528 1803 532 1807
rect 616 1803 620 1807
rect 704 1803 708 1807
rect 784 1803 788 1807
rect 864 1803 868 1807
rect 944 1803 948 1807
rect 1032 1803 1036 1807
rect 1392 1803 1396 1807
rect 1488 1803 1492 1807
rect 1600 1803 1604 1807
rect 1712 1803 1716 1807
rect 1760 1803 1764 1807
rect 1816 1803 1820 1807
rect 1928 1803 1932 1807
rect 2040 1803 2044 1807
rect 2160 1803 2164 1807
rect 2280 1803 2284 1807
rect 2408 1803 2412 1807
rect 2520 1803 2524 1807
rect 208 1787 212 1791
rect 272 1787 276 1791
rect 344 1787 348 1791
rect 424 1787 428 1791
rect 512 1787 516 1791
rect 600 1787 604 1791
rect 680 1787 684 1791
rect 688 1787 692 1791
rect 768 1787 772 1791
rect 848 1787 852 1791
rect 928 1787 932 1791
rect 1008 1787 1012 1791
rect 1056 1787 1060 1791
rect 1096 1787 1100 1791
rect 248 1751 252 1755
rect 312 1751 316 1755
rect 384 1751 388 1755
rect 464 1751 468 1755
rect 552 1751 556 1755
rect 640 1751 644 1755
rect 728 1751 732 1755
rect 808 1751 812 1755
rect 888 1753 892 1757
rect 1432 1767 1436 1771
rect 1528 1767 1532 1771
rect 1640 1767 1644 1771
rect 1752 1767 1756 1771
rect 1760 1767 1764 1771
rect 1856 1767 1860 1771
rect 1968 1767 1972 1771
rect 2080 1767 2084 1771
rect 2200 1767 2204 1771
rect 2320 1767 2324 1771
rect 2448 1767 2452 1771
rect 2560 1767 2564 1771
rect 968 1751 972 1755
rect 1048 1751 1052 1755
rect 1056 1751 1060 1755
rect 1136 1751 1140 1755
rect 1064 1747 1068 1751
rect 384 1719 388 1723
rect 440 1719 444 1723
rect 504 1719 508 1723
rect 584 1719 588 1723
rect 672 1719 676 1723
rect 680 1719 684 1723
rect 688 1723 692 1727
rect 768 1723 772 1727
rect 760 1719 764 1723
rect 856 1719 860 1723
rect 952 1719 956 1723
rect 1048 1719 1052 1723
rect 1480 1743 1484 1747
rect 1560 1743 1564 1747
rect 1656 1743 1660 1747
rect 1864 1743 1868 1747
rect 1472 1739 1476 1743
rect 1144 1719 1148 1723
rect 1240 1719 1244 1723
rect 1552 1739 1556 1743
rect 1648 1739 1652 1743
rect 1752 1739 1756 1743
rect 1856 1739 1860 1743
rect 1960 1739 1964 1743
rect 2056 1739 2060 1743
rect 2152 1739 2156 1743
rect 2240 1739 2244 1743
rect 2320 1739 2324 1743
rect 2408 1739 2412 1743
rect 2496 1739 2500 1743
rect 2560 1739 2564 1743
rect 1432 1703 1436 1707
rect 1480 1703 1484 1707
rect 1512 1703 1516 1707
rect 1560 1703 1564 1707
rect 1608 1703 1612 1707
rect 1656 1703 1660 1707
rect 1712 1703 1716 1707
rect 1816 1703 1820 1707
rect 1864 1703 1868 1707
rect 1920 1703 1924 1707
rect 2016 1703 2020 1707
rect 2112 1703 2116 1707
rect 2200 1703 2204 1707
rect 2280 1703 2284 1707
rect 2368 1703 2372 1707
rect 2456 1703 2460 1707
rect 2520 1703 2524 1707
rect 344 1683 348 1687
rect 400 1683 404 1687
rect 464 1683 468 1687
rect 544 1683 548 1687
rect 632 1683 636 1687
rect 688 1683 692 1687
rect 720 1683 724 1687
rect 768 1683 772 1687
rect 816 1683 820 1687
rect 912 1683 916 1687
rect 1008 1683 1012 1687
rect 1064 1683 1068 1687
rect 1104 1683 1108 1687
rect 1200 1683 1204 1687
rect 1536 1679 1540 1683
rect 1608 1679 1612 1683
rect 1688 1679 1692 1683
rect 1776 1679 1780 1683
rect 1864 1679 1868 1683
rect 1952 1679 1956 1683
rect 2040 1679 2044 1683
rect 2120 1679 2124 1683
rect 2192 1679 2196 1683
rect 2264 1679 2268 1683
rect 2328 1679 2332 1683
rect 2400 1679 2404 1683
rect 2464 1679 2468 1683
rect 2520 1679 2524 1683
rect 376 1667 380 1671
rect 424 1667 428 1671
rect 432 1667 436 1671
rect 488 1667 492 1671
rect 552 1667 556 1671
rect 624 1667 628 1671
rect 704 1667 708 1671
rect 784 1667 788 1671
rect 864 1667 868 1671
rect 912 1667 916 1671
rect 944 1667 948 1671
rect 1024 1667 1028 1671
rect 1112 1667 1116 1671
rect 1200 1667 1204 1671
rect 1264 1667 1268 1671
rect 416 1631 420 1635
rect 424 1631 428 1635
rect 472 1631 476 1635
rect 528 1631 532 1635
rect 592 1631 596 1635
rect 664 1631 668 1635
rect 744 1633 748 1637
rect 1576 1643 1580 1647
rect 1648 1643 1652 1647
rect 1728 1643 1732 1647
rect 1816 1643 1820 1647
rect 1904 1643 1908 1647
rect 1992 1643 1996 1647
rect 2080 1643 2084 1647
rect 2160 1643 2164 1647
rect 2232 1643 2236 1647
rect 2304 1643 2308 1647
rect 2368 1643 2372 1647
rect 2440 1643 2444 1647
rect 2504 1643 2508 1647
rect 2560 1643 2564 1647
rect 824 1631 828 1635
rect 904 1631 908 1635
rect 912 1631 916 1635
rect 984 1631 988 1635
rect 1064 1631 1068 1635
rect 1152 1631 1156 1635
rect 1240 1631 1244 1635
rect 1304 1631 1308 1635
rect 1616 1607 1620 1611
rect 1672 1607 1676 1611
rect 1728 1607 1732 1611
rect 1792 1607 1796 1611
rect 1608 1603 1612 1607
rect 1104 1591 1108 1595
rect 320 1587 324 1591
rect 400 1587 404 1591
rect 488 1587 492 1591
rect 584 1587 588 1591
rect 680 1587 684 1591
rect 768 1587 772 1591
rect 856 1587 860 1591
rect 936 1587 940 1591
rect 968 1587 972 1591
rect 1016 1587 1020 1591
rect 1096 1587 1100 1591
rect 1184 1587 1188 1591
rect 1664 1603 1668 1607
rect 1720 1603 1724 1607
rect 1784 1603 1788 1607
rect 1864 1603 1868 1607
rect 1952 1603 1956 1607
rect 2040 1603 2044 1607
rect 2136 1603 2140 1607
rect 2240 1603 2244 1607
rect 2352 1603 2356 1607
rect 2464 1603 2468 1607
rect 2560 1603 2564 1607
rect 1568 1567 1572 1571
rect 1616 1567 1620 1571
rect 1624 1567 1628 1571
rect 1672 1567 1676 1571
rect 1680 1567 1684 1571
rect 1728 1567 1732 1571
rect 1744 1567 1748 1571
rect 1792 1567 1796 1571
rect 1824 1567 1828 1571
rect 1912 1567 1916 1571
rect 2000 1567 2004 1571
rect 2096 1567 2100 1571
rect 2192 1567 2196 1571
rect 2200 1567 2204 1571
rect 2312 1567 2316 1571
rect 2424 1567 2428 1571
rect 2520 1567 2524 1571
rect 280 1551 284 1555
rect 360 1551 364 1555
rect 448 1551 452 1555
rect 544 1551 548 1555
rect 640 1551 644 1555
rect 728 1551 732 1555
rect 816 1551 820 1555
rect 896 1551 900 1555
rect 968 1551 972 1555
rect 976 1551 980 1555
rect 1056 1551 1060 1555
rect 1104 1551 1108 1555
rect 1144 1551 1148 1555
rect 1656 1551 1660 1555
rect 1704 1551 1708 1555
rect 1712 1551 1716 1555
rect 1768 1551 1772 1555
rect 1832 1551 1836 1555
rect 1904 1551 1908 1555
rect 1984 1551 1988 1555
rect 2064 1551 2068 1555
rect 2144 1551 2148 1555
rect 256 1539 260 1543
rect 312 1539 316 1543
rect 376 1539 380 1543
rect 448 1539 452 1543
rect 520 1539 524 1543
rect 592 1539 596 1543
rect 664 1539 668 1543
rect 736 1539 740 1543
rect 808 1539 812 1543
rect 880 1539 884 1543
rect 952 1539 956 1543
rect 1032 1539 1036 1543
rect 2224 1551 2228 1555
rect 2304 1551 2308 1555
rect 2384 1551 2388 1555
rect 2464 1551 2468 1555
rect 2520 1551 2524 1555
rect 1696 1515 1700 1519
rect 1704 1515 1708 1519
rect 1752 1515 1756 1519
rect 1808 1515 1812 1519
rect 1872 1515 1876 1519
rect 1944 1515 1948 1519
rect 2024 1515 2028 1519
rect 2104 1515 2108 1519
rect 2184 1515 2188 1519
rect 2192 1515 2196 1519
rect 2264 1515 2268 1519
rect 2344 1515 2348 1519
rect 2424 1515 2428 1519
rect 2504 1515 2508 1519
rect 2560 1515 2564 1519
rect 296 1503 300 1507
rect 352 1503 356 1507
rect 416 1503 420 1507
rect 488 1503 492 1507
rect 560 1503 564 1507
rect 632 1503 636 1507
rect 704 1503 708 1507
rect 776 1503 780 1507
rect 848 1503 852 1507
rect 920 1503 924 1507
rect 992 1503 996 1507
rect 1072 1503 1076 1507
rect 1552 1479 1556 1483
rect 1608 1479 1612 1483
rect 1680 1479 1684 1483
rect 1760 1479 1764 1483
rect 1840 1479 1844 1483
rect 1928 1479 1932 1483
rect 2016 1479 2020 1483
rect 2104 1479 2108 1483
rect 2184 1479 2188 1483
rect 2264 1479 2268 1483
rect 2344 1479 2348 1483
rect 2424 1479 2428 1483
rect 2504 1479 2508 1483
rect 2560 1479 2564 1483
rect 528 1475 532 1479
rect 232 1471 236 1475
rect 320 1471 324 1475
rect 416 1471 420 1475
rect 520 1471 524 1475
rect 616 1471 620 1475
rect 712 1471 716 1475
rect 808 1471 812 1475
rect 896 1471 900 1475
rect 984 1471 988 1475
rect 1072 1471 1076 1475
rect 1168 1471 1172 1475
rect 1512 1443 1516 1447
rect 1568 1443 1572 1447
rect 1640 1443 1644 1447
rect 1720 1443 1724 1447
rect 1800 1443 1804 1447
rect 1888 1443 1892 1447
rect 1976 1443 1980 1447
rect 2064 1443 2068 1447
rect 2144 1443 2148 1447
rect 2224 1443 2228 1447
rect 2304 1443 2308 1447
rect 2384 1443 2388 1447
rect 2464 1443 2468 1447
rect 2520 1443 2524 1447
rect 192 1435 196 1439
rect 280 1435 284 1439
rect 376 1435 380 1439
rect 480 1435 484 1439
rect 528 1435 532 1439
rect 576 1435 580 1439
rect 672 1435 676 1439
rect 768 1435 772 1439
rect 856 1435 860 1439
rect 944 1435 948 1439
rect 1032 1435 1036 1439
rect 1128 1435 1132 1439
rect 1392 1423 1396 1427
rect 1448 1423 1452 1427
rect 1512 1423 1516 1427
rect 1600 1423 1604 1427
rect 1696 1423 1700 1427
rect 1744 1423 1748 1427
rect 1800 1423 1804 1427
rect 1904 1423 1908 1427
rect 2000 1423 2004 1427
rect 2096 1423 2100 1427
rect 2192 1423 2196 1427
rect 2280 1423 2284 1427
rect 2328 1423 2332 1427
rect 2368 1423 2372 1427
rect 2416 1423 2420 1427
rect 2456 1423 2460 1427
rect 2520 1423 2524 1427
rect 136 1419 140 1423
rect 224 1419 228 1423
rect 320 1419 324 1423
rect 424 1419 428 1423
rect 528 1419 532 1423
rect 640 1419 644 1423
rect 744 1419 748 1423
rect 856 1419 860 1423
rect 968 1419 972 1423
rect 1080 1419 1084 1423
rect 1192 1419 1196 1423
rect 1432 1387 1436 1391
rect 1488 1387 1492 1391
rect 1552 1387 1556 1391
rect 1640 1387 1644 1391
rect 1736 1387 1740 1391
rect 1744 1387 1748 1391
rect 1840 1387 1844 1391
rect 1944 1387 1948 1391
rect 2040 1387 2044 1391
rect 2136 1387 2140 1391
rect 2232 1387 2236 1391
rect 2320 1387 2324 1391
rect 2328 1387 2332 1391
rect 2408 1389 2412 1393
rect 2416 1391 2420 1395
rect 2496 1387 2500 1391
rect 2560 1387 2564 1391
rect 176 1383 180 1387
rect 264 1383 268 1387
rect 360 1383 364 1387
rect 464 1383 468 1387
rect 568 1383 572 1387
rect 680 1383 684 1387
rect 784 1383 788 1387
rect 896 1383 900 1387
rect 1008 1383 1012 1387
rect 1120 1383 1124 1387
rect 1232 1383 1236 1387
rect 552 1359 556 1363
rect 176 1355 180 1359
rect 240 1355 244 1359
rect 328 1355 332 1359
rect 432 1355 436 1359
rect 544 1355 548 1359
rect 656 1355 660 1359
rect 768 1355 772 1359
rect 880 1355 884 1359
rect 992 1355 996 1359
rect 1104 1355 1108 1359
rect 1216 1355 1220 1359
rect 1304 1355 1308 1359
rect 1848 1355 1852 1359
rect 1432 1351 1436 1355
rect 1488 1351 1492 1355
rect 1576 1351 1580 1355
rect 1664 1351 1668 1355
rect 1752 1351 1756 1355
rect 1840 1351 1844 1355
rect 136 1319 140 1323
rect 200 1319 204 1323
rect 288 1319 292 1323
rect 392 1319 396 1323
rect 504 1319 508 1323
rect 552 1319 556 1323
rect 616 1319 620 1323
rect 728 1319 732 1323
rect 840 1319 844 1323
rect 952 1319 956 1323
rect 1064 1319 1068 1323
rect 1176 1319 1180 1323
rect 1264 1319 1268 1323
rect 1920 1351 1924 1355
rect 2000 1351 2004 1355
rect 2080 1351 2084 1355
rect 2160 1351 2164 1355
rect 2240 1351 2244 1355
rect 1392 1315 1396 1319
rect 1448 1315 1452 1319
rect 1536 1315 1540 1319
rect 1624 1315 1628 1319
rect 1712 1315 1716 1319
rect 1800 1315 1804 1319
rect 1848 1315 1852 1319
rect 1880 1315 1884 1319
rect 1960 1315 1964 1319
rect 2040 1315 2044 1319
rect 2120 1315 2124 1319
rect 2200 1315 2204 1319
rect 136 1307 140 1311
rect 208 1307 212 1311
rect 304 1307 308 1311
rect 408 1307 412 1311
rect 512 1307 516 1311
rect 608 1307 612 1311
rect 704 1307 708 1311
rect 800 1307 804 1311
rect 888 1307 892 1311
rect 968 1307 972 1311
rect 1048 1307 1052 1311
rect 1128 1307 1132 1311
rect 1208 1307 1212 1311
rect 1264 1307 1268 1311
rect 1736 1303 1740 1307
rect 1648 1299 1652 1303
rect 176 1271 180 1275
rect 248 1271 252 1275
rect 344 1271 348 1275
rect 448 1271 452 1275
rect 552 1271 556 1275
rect 648 1271 652 1275
rect 744 1271 748 1275
rect 840 1271 844 1275
rect 928 1271 932 1275
rect 1008 1271 1012 1275
rect 1088 1273 1092 1277
rect 1168 1271 1172 1275
rect 1248 1271 1252 1275
rect 1304 1271 1308 1275
rect 1688 1263 1692 1267
rect 1744 1299 1748 1303
rect 1840 1299 1844 1303
rect 1936 1299 1940 1303
rect 2024 1299 2028 1303
rect 2112 1299 2116 1303
rect 2208 1299 2212 1303
rect 1784 1263 1788 1267
rect 1880 1263 1884 1267
rect 1976 1263 1980 1267
rect 2064 1263 2068 1267
rect 2152 1263 2156 1267
rect 2248 1263 2252 1267
rect 1736 1259 1740 1263
rect 1864 1239 1868 1243
rect 1528 1235 1532 1239
rect 1592 1235 1596 1239
rect 1656 1235 1660 1239
rect 1720 1235 1724 1239
rect 1792 1235 1796 1239
rect 1856 1235 1860 1239
rect 176 1231 180 1235
rect 232 1231 236 1235
rect 312 1231 316 1235
rect 392 1231 396 1235
rect 472 1231 476 1235
rect 552 1231 556 1235
rect 632 1231 636 1235
rect 704 1231 708 1235
rect 776 1231 780 1235
rect 848 1231 852 1235
rect 928 1231 932 1235
rect 1920 1235 1924 1239
rect 1984 1235 1988 1239
rect 2048 1235 2052 1239
rect 2112 1235 2116 1239
rect 2184 1235 2188 1239
rect 2256 1235 2260 1239
rect 2328 1235 2332 1239
rect 1488 1199 1492 1203
rect 1552 1199 1556 1203
rect 1616 1199 1620 1203
rect 1680 1199 1684 1203
rect 1752 1199 1756 1203
rect 1816 1199 1820 1203
rect 1864 1199 1868 1203
rect 1880 1199 1884 1203
rect 1944 1199 1948 1203
rect 2008 1199 2012 1203
rect 2072 1199 2076 1203
rect 2144 1199 2148 1203
rect 2216 1199 2220 1203
rect 2288 1199 2292 1203
rect 136 1195 140 1199
rect 192 1195 196 1199
rect 272 1195 276 1199
rect 352 1195 356 1199
rect 432 1195 436 1199
rect 512 1195 516 1199
rect 592 1195 596 1199
rect 664 1195 668 1199
rect 736 1195 740 1199
rect 808 1195 812 1199
rect 888 1195 892 1199
rect 136 1179 140 1183
rect 184 1179 188 1183
rect 216 1179 220 1183
rect 304 1179 308 1183
rect 400 1179 404 1183
rect 488 1179 492 1183
rect 536 1179 540 1183
rect 576 1179 580 1183
rect 664 1179 668 1183
rect 744 1179 748 1183
rect 816 1179 820 1183
rect 888 1179 892 1183
rect 952 1179 956 1183
rect 960 1179 964 1183
rect 1040 1179 1044 1183
rect 1392 1179 1396 1183
rect 1480 1179 1484 1183
rect 1576 1181 1580 1185
rect 1680 1179 1684 1183
rect 1784 1179 1788 1183
rect 1888 1179 1892 1183
rect 1992 1179 1996 1183
rect 2088 1179 2092 1183
rect 2184 1179 2188 1183
rect 2280 1179 2284 1183
rect 2376 1179 2380 1183
rect 176 1143 180 1147
rect 184 1143 188 1147
rect 256 1143 260 1147
rect 344 1143 348 1147
rect 440 1143 444 1147
rect 528 1143 532 1147
rect 536 1143 540 1147
rect 616 1143 620 1147
rect 704 1143 708 1147
rect 784 1143 788 1147
rect 856 1143 860 1147
rect 928 1143 932 1147
rect 1000 1143 1004 1147
rect 1080 1143 1084 1147
rect 1432 1143 1436 1147
rect 1520 1143 1524 1147
rect 1616 1143 1620 1147
rect 1720 1143 1724 1147
rect 1824 1143 1828 1147
rect 1928 1143 1932 1147
rect 2032 1143 2036 1147
rect 2128 1143 2132 1147
rect 2224 1143 2228 1147
rect 2320 1143 2324 1147
rect 2416 1143 2420 1147
rect 1936 1139 1940 1143
rect 1728 1115 1732 1119
rect 256 1107 260 1111
rect 352 1107 356 1111
rect 456 1107 460 1111
rect 560 1107 564 1111
rect 664 1107 668 1111
rect 760 1107 764 1111
rect 856 1107 860 1111
rect 944 1107 948 1111
rect 952 1107 956 1111
rect 1024 1107 1028 1111
rect 1112 1107 1116 1111
rect 1200 1109 1204 1113
rect 1432 1111 1436 1115
rect 1512 1111 1516 1115
rect 1616 1111 1620 1115
rect 1720 1111 1724 1115
rect 1824 1111 1828 1115
rect 1920 1111 1924 1115
rect 2384 1115 2388 1119
rect 2008 1111 2012 1115
rect 2096 1111 2100 1115
rect 2176 1111 2180 1115
rect 2248 1111 2252 1115
rect 2312 1111 2316 1115
rect 2376 1111 2380 1115
rect 2440 1111 2444 1115
rect 2504 1111 2508 1115
rect 2560 1111 2564 1115
rect 1392 1075 1396 1079
rect 1472 1075 1476 1079
rect 1576 1075 1580 1079
rect 1680 1075 1684 1079
rect 1728 1075 1732 1079
rect 1784 1075 1788 1079
rect 1880 1075 1884 1079
rect 1936 1075 1940 1079
rect 1968 1075 1972 1079
rect 2056 1075 2060 1079
rect 2136 1075 2140 1079
rect 2208 1075 2212 1079
rect 2272 1075 2276 1079
rect 2336 1075 2340 1079
rect 2384 1075 2388 1079
rect 2400 1075 2404 1079
rect 2464 1075 2468 1079
rect 2520 1075 2524 1079
rect 216 1071 220 1075
rect 312 1071 316 1075
rect 416 1071 420 1075
rect 520 1071 524 1075
rect 624 1071 628 1075
rect 720 1071 724 1075
rect 816 1071 820 1075
rect 904 1071 908 1075
rect 984 1071 988 1075
rect 1072 1071 1076 1075
rect 1160 1071 1164 1075
rect 1440 1063 1444 1067
rect 1384 1059 1388 1063
rect 1392 1059 1396 1063
rect 288 1055 292 1059
rect 336 1055 340 1059
rect 344 1055 348 1059
rect 416 1055 420 1059
rect 496 1055 500 1059
rect 584 1055 588 1059
rect 680 1055 684 1059
rect 776 1055 780 1059
rect 864 1055 868 1059
rect 952 1055 956 1059
rect 1032 1055 1036 1059
rect 1112 1055 1116 1059
rect 1200 1055 1204 1059
rect 1264 1055 1268 1059
rect 1432 1023 1436 1027
rect 1448 1059 1452 1063
rect 1512 1059 1516 1063
rect 1600 1059 1604 1063
rect 1704 1059 1708 1063
rect 1816 1059 1820 1063
rect 1928 1059 1932 1063
rect 2040 1059 2044 1063
rect 2144 1059 2148 1063
rect 2248 1059 2252 1063
rect 2344 1059 2348 1063
rect 2440 1059 2444 1063
rect 2520 1059 2524 1063
rect 1488 1023 1492 1027
rect 1552 1023 1556 1027
rect 1640 1023 1644 1027
rect 1744 1023 1748 1027
rect 1856 1023 1860 1027
rect 1968 1023 1972 1027
rect 2080 1023 2084 1027
rect 2184 1023 2188 1027
rect 2288 1023 2292 1027
rect 2384 1023 2388 1027
rect 2480 1023 2484 1027
rect 2560 1023 2564 1027
rect 328 1019 332 1023
rect 336 1019 340 1023
rect 384 1019 388 1023
rect 456 1019 460 1023
rect 536 1019 540 1023
rect 624 1019 628 1023
rect 720 1019 724 1023
rect 816 1019 820 1023
rect 904 1019 908 1023
rect 992 1019 996 1023
rect 1072 1019 1076 1023
rect 1152 1019 1156 1023
rect 1240 1019 1244 1023
rect 1304 1019 1308 1023
rect 1384 1019 1388 1023
rect 1440 1019 1444 1023
rect 1864 1019 1868 1023
rect 1016 991 1020 995
rect 1080 991 1084 995
rect 1144 991 1148 995
rect 1200 991 1204 995
rect 1256 991 1260 995
rect 448 987 452 991
rect 504 987 508 991
rect 560 987 564 991
rect 624 987 628 991
rect 688 987 692 991
rect 752 987 756 991
rect 816 987 820 991
rect 880 987 884 991
rect 944 987 948 991
rect 1008 987 1012 991
rect 1072 987 1076 991
rect 1136 987 1140 991
rect 1192 987 1196 991
rect 1248 987 1252 991
rect 1304 987 1308 991
rect 1432 979 1436 983
rect 1488 979 1492 983
rect 1544 979 1548 983
rect 1600 979 1604 983
rect 1672 979 1676 983
rect 1752 979 1756 983
rect 1840 979 1844 983
rect 408 951 412 955
rect 464 951 468 955
rect 520 951 524 955
rect 584 951 588 955
rect 648 951 652 955
rect 712 951 716 955
rect 776 951 780 955
rect 840 951 844 955
rect 904 951 908 955
rect 968 951 972 955
rect 1016 951 1020 955
rect 1032 951 1036 955
rect 1080 951 1084 955
rect 1096 951 1100 955
rect 1144 951 1148 955
rect 1152 951 1156 955
rect 1200 951 1204 955
rect 1208 951 1212 955
rect 1256 951 1260 955
rect 1264 951 1268 955
rect 1936 979 1940 983
rect 2048 979 2052 983
rect 2176 979 2180 983
rect 2304 979 2308 983
rect 2440 979 2444 983
rect 2560 979 2564 983
rect 1392 943 1396 947
rect 1448 943 1452 947
rect 1504 943 1508 947
rect 1560 943 1564 947
rect 1632 943 1636 947
rect 1712 943 1716 947
rect 1800 943 1804 947
rect 1864 943 1868 947
rect 1896 943 1900 947
rect 2008 943 2012 947
rect 2136 943 2140 947
rect 2264 943 2268 947
rect 2400 943 2404 947
rect 2520 943 2524 947
rect 400 935 404 939
rect 456 935 460 939
rect 512 935 516 939
rect 568 935 572 939
rect 616 935 620 939
rect 624 935 628 939
rect 680 935 684 939
rect 736 937 740 941
rect 792 935 796 939
rect 1392 923 1396 927
rect 1448 923 1452 927
rect 1504 923 1508 927
rect 1592 923 1596 927
rect 1680 923 1684 927
rect 1688 923 1692 927
rect 1736 923 1740 927
rect 1800 923 1804 927
rect 1920 923 1924 927
rect 2040 923 2044 927
rect 2160 923 2164 927
rect 2288 923 2292 927
rect 2416 923 2420 927
rect 2520 923 2524 927
rect 440 899 444 903
rect 496 899 500 903
rect 552 899 556 903
rect 608 899 612 903
rect 616 899 620 903
rect 664 899 668 903
rect 720 899 724 903
rect 776 899 780 903
rect 832 899 836 903
rect 1432 887 1436 891
rect 1488 887 1492 891
rect 1544 887 1548 891
rect 1632 887 1636 891
rect 312 871 316 875
rect 368 871 372 875
rect 424 871 428 875
rect 488 871 492 875
rect 552 871 556 875
rect 616 871 620 875
rect 680 871 684 875
rect 744 871 748 875
rect 808 871 812 875
rect 880 871 884 875
rect 952 871 956 875
rect 1728 887 1732 891
rect 1736 887 1740 891
rect 1840 887 1844 891
rect 1960 887 1964 891
rect 2080 887 2084 891
rect 2200 887 2204 891
rect 2328 887 2332 891
rect 2456 887 2460 891
rect 2560 887 2564 891
rect 1504 859 1508 863
rect 1584 859 1588 863
rect 1672 859 1676 863
rect 1680 859 1684 863
rect 1760 859 1764 863
rect 1848 859 1852 863
rect 1936 859 1940 863
rect 2024 859 2028 863
rect 2104 859 2108 863
rect 2176 859 2180 863
rect 2248 859 2252 863
rect 2312 859 2316 863
rect 2376 859 2380 863
rect 2440 859 2444 863
rect 2504 859 2508 863
rect 2560 859 2564 863
rect 272 835 276 839
rect 328 835 332 839
rect 384 835 388 839
rect 448 835 452 839
rect 512 835 516 839
rect 576 835 580 839
rect 640 835 644 839
rect 704 835 708 839
rect 768 835 772 839
rect 840 835 844 839
rect 912 835 916 839
rect 1464 823 1468 827
rect 1544 823 1548 827
rect 1632 823 1636 827
rect 1720 823 1724 827
rect 1808 823 1812 827
rect 1896 823 1900 827
rect 1984 823 1988 827
rect 2064 823 2068 827
rect 2136 823 2140 827
rect 2208 823 2212 827
rect 2272 823 2276 827
rect 2336 823 2340 827
rect 2400 823 2404 827
rect 2464 823 2468 827
rect 2520 823 2524 827
rect 144 815 148 819
rect 208 815 212 819
rect 288 815 292 819
rect 376 815 380 819
rect 464 815 468 819
rect 560 815 564 819
rect 648 815 652 819
rect 736 815 740 819
rect 816 815 820 819
rect 864 815 868 819
rect 896 815 900 819
rect 944 815 948 819
rect 984 815 988 819
rect 1072 815 1076 819
rect 1608 803 1612 807
rect 1656 803 1660 807
rect 1664 803 1668 807
rect 1728 803 1732 807
rect 1800 803 1804 807
rect 1880 803 1884 807
rect 1960 803 1964 807
rect 1968 803 1972 807
rect 2048 803 2052 807
rect 2136 803 2140 807
rect 2224 803 2228 807
rect 2312 803 2316 807
rect 2360 803 2364 807
rect 2400 803 2404 807
rect 184 779 188 783
rect 248 779 252 783
rect 328 779 332 783
rect 416 779 420 783
rect 504 779 508 783
rect 600 779 604 783
rect 688 779 692 783
rect 776 779 780 783
rect 856 779 860 783
rect 864 779 868 783
rect 936 781 940 785
rect 944 783 948 787
rect 1024 779 1028 783
rect 1112 779 1116 783
rect 1648 767 1652 771
rect 1656 767 1660 771
rect 1704 767 1708 771
rect 1768 767 1772 771
rect 1840 767 1844 771
rect 1920 767 1924 771
rect 176 743 180 747
rect 232 743 236 747
rect 312 743 316 747
rect 416 743 420 747
rect 520 743 524 747
rect 632 743 636 747
rect 736 743 740 747
rect 840 743 844 747
rect 936 743 940 747
rect 1024 743 1028 747
rect 1112 743 1116 747
rect 1208 743 1212 747
rect 2008 767 2012 771
rect 2088 767 2092 771
rect 2176 767 2180 771
rect 2264 767 2268 771
rect 2352 767 2356 771
rect 2360 767 2364 771
rect 2440 767 2444 771
rect 1600 735 1604 739
rect 1656 735 1660 739
rect 1720 735 1724 739
rect 1792 735 1796 739
rect 1872 735 1876 739
rect 1952 735 1956 739
rect 1960 735 1964 739
rect 2032 735 2036 739
rect 2112 735 2116 739
rect 2192 735 2196 739
rect 2280 735 2284 739
rect 2368 735 2372 739
rect 136 707 140 711
rect 192 707 196 711
rect 272 707 276 711
rect 376 707 380 711
rect 480 707 484 711
rect 592 707 596 711
rect 696 707 700 711
rect 800 707 804 711
rect 896 707 900 711
rect 984 707 988 711
rect 1072 707 1076 711
rect 1168 707 1172 711
rect 1560 699 1564 703
rect 1616 699 1620 703
rect 1680 699 1684 703
rect 1752 699 1756 703
rect 1832 699 1836 703
rect 1912 699 1916 703
rect 1992 699 1996 703
rect 2072 699 2076 703
rect 2152 699 2156 703
rect 2240 699 2244 703
rect 2328 699 2332 703
rect 136 691 140 695
rect 192 691 196 695
rect 256 691 260 695
rect 304 691 308 695
rect 336 691 340 695
rect 424 691 428 695
rect 512 691 516 695
rect 600 691 604 695
rect 688 691 692 695
rect 768 691 772 695
rect 848 691 852 695
rect 928 691 932 695
rect 1016 691 1020 695
rect 1392 683 1396 687
rect 1488 683 1492 687
rect 1536 683 1540 687
rect 1592 683 1596 687
rect 1640 683 1644 687
rect 1696 683 1700 687
rect 1800 683 1804 687
rect 1904 683 1908 687
rect 2000 683 2004 687
rect 2096 683 2100 687
rect 2184 683 2188 687
rect 2272 683 2276 687
rect 2368 683 2372 687
rect 176 655 180 659
rect 232 655 236 659
rect 296 657 300 661
rect 304 659 308 663
rect 376 655 380 659
rect 464 655 468 659
rect 552 655 556 659
rect 640 655 644 659
rect 728 655 732 659
rect 808 655 812 659
rect 888 655 892 659
rect 968 655 972 659
rect 1056 655 1060 659
rect 1432 647 1436 651
rect 1528 647 1532 651
rect 1536 647 1540 651
rect 1632 647 1636 651
rect 1640 647 1644 651
rect 1736 647 1740 651
rect 1840 647 1844 651
rect 1944 647 1948 651
rect 2040 647 2044 651
rect 2136 647 2140 651
rect 2224 647 2228 651
rect 2312 647 2316 651
rect 2408 647 2412 651
rect 1440 623 1444 627
rect 1952 623 1956 627
rect 176 619 180 623
rect 232 619 236 623
rect 288 619 292 623
rect 344 619 348 623
rect 424 619 428 623
rect 512 619 516 623
rect 608 619 612 623
rect 712 619 716 623
rect 816 619 820 623
rect 920 619 924 623
rect 1024 619 1028 623
rect 1120 619 1124 623
rect 1224 619 1228 623
rect 1304 619 1308 623
rect 1432 619 1436 623
rect 1544 619 1548 623
rect 1680 619 1684 623
rect 1816 619 1820 623
rect 1944 619 1948 623
rect 2072 619 2076 623
rect 2192 619 2196 623
rect 2312 619 2316 623
rect 2440 619 2444 623
rect 136 583 140 587
rect 192 583 196 587
rect 248 583 252 587
rect 304 583 308 587
rect 384 583 388 587
rect 472 583 476 587
rect 568 583 572 587
rect 672 583 676 587
rect 776 583 780 587
rect 880 583 884 587
rect 984 583 988 587
rect 1080 583 1084 587
rect 1184 583 1188 587
rect 1264 583 1268 587
rect 1392 583 1396 587
rect 1440 583 1444 587
rect 1504 583 1508 587
rect 1640 583 1644 587
rect 1776 583 1780 587
rect 1904 583 1908 587
rect 1952 583 1956 587
rect 2032 583 2036 587
rect 2152 583 2156 587
rect 2272 583 2276 587
rect 2400 583 2404 587
rect 176 567 180 571
rect 224 567 228 571
rect 240 567 244 571
rect 296 567 300 571
rect 312 567 316 571
rect 392 567 396 571
rect 472 567 476 571
rect 488 567 492 571
rect 592 567 596 571
rect 696 567 700 571
rect 808 567 812 571
rect 920 567 924 571
rect 1040 567 1044 571
rect 1160 567 1164 571
rect 1264 567 1268 571
rect 216 533 220 537
rect 224 535 228 539
rect 280 531 284 535
rect 296 531 300 535
rect 352 531 356 535
rect 432 531 436 535
rect 1392 563 1396 567
rect 1448 563 1452 567
rect 1528 563 1532 567
rect 1624 563 1628 567
rect 1728 563 1732 567
rect 1832 563 1836 567
rect 1936 563 1940 567
rect 1984 563 1988 567
rect 2032 563 2036 567
rect 2128 563 2132 567
rect 2216 563 2220 567
rect 2296 563 2300 567
rect 2376 563 2380 567
rect 2456 563 2460 567
rect 2520 563 2524 567
rect 528 531 532 535
rect 632 531 636 535
rect 736 531 740 535
rect 848 531 852 535
rect 960 531 964 535
rect 1080 531 1084 535
rect 1200 531 1204 535
rect 1304 531 1308 535
rect 1432 527 1436 531
rect 1488 527 1492 531
rect 1568 527 1572 531
rect 1664 527 1668 531
rect 1768 527 1772 531
rect 1872 527 1876 531
rect 1976 527 1980 531
rect 1984 527 1988 531
rect 2072 527 2076 531
rect 2168 527 2172 531
rect 2256 527 2260 531
rect 2336 527 2340 531
rect 2416 527 2420 531
rect 2496 527 2500 531
rect 2560 527 2564 531
rect 2512 503 2516 507
rect 1568 499 1572 503
rect 1632 499 1636 503
rect 1704 499 1708 503
rect 1784 499 1788 503
rect 1872 499 1876 503
rect 1960 499 1964 503
rect 2048 499 2052 503
rect 2128 499 2132 503
rect 2208 499 2212 503
rect 2288 499 2292 503
rect 2360 499 2364 503
rect 2432 499 2436 503
rect 2504 499 2508 503
rect 336 495 340 499
rect 392 495 396 499
rect 456 495 460 499
rect 472 495 476 499
rect 528 495 532 499
rect 608 495 612 499
rect 680 495 684 499
rect 752 495 756 499
rect 824 495 828 499
rect 896 495 900 499
rect 968 495 972 499
rect 1040 495 1044 499
rect 1120 495 1124 499
rect 2560 499 2564 503
rect 1528 463 1532 467
rect 1592 463 1596 467
rect 1664 463 1668 467
rect 1744 463 1748 467
rect 1832 463 1836 467
rect 1920 463 1924 467
rect 2008 463 2012 467
rect 2088 463 2092 467
rect 2168 463 2172 467
rect 2248 463 2252 467
rect 2320 463 2324 467
rect 2392 463 2396 467
rect 2464 463 2468 467
rect 2512 463 2516 467
rect 2520 463 2524 467
rect 296 459 300 463
rect 352 459 356 463
rect 416 459 420 463
rect 488 459 492 463
rect 568 459 572 463
rect 640 459 644 463
rect 712 459 716 463
rect 784 459 788 463
rect 856 459 860 463
rect 928 459 932 463
rect 1000 459 1004 463
rect 1080 459 1084 463
rect 432 443 436 447
rect 488 443 492 447
rect 552 443 556 447
rect 624 443 628 447
rect 704 443 708 447
rect 776 443 780 447
rect 848 443 852 447
rect 920 443 924 447
rect 992 443 996 447
rect 1064 443 1068 447
rect 1136 443 1140 447
rect 1216 443 1220 447
rect 1624 443 1628 447
rect 1680 443 1684 447
rect 1736 443 1740 447
rect 1792 443 1796 447
rect 1848 443 1852 447
rect 1904 443 1908 447
rect 1976 443 1980 447
rect 2064 443 2068 447
rect 2168 443 2172 447
rect 2288 443 2292 447
rect 2416 443 2420 447
rect 2520 443 2524 447
rect 472 407 476 411
rect 528 407 532 411
rect 592 407 596 411
rect 664 407 668 411
rect 744 407 748 411
rect 816 407 820 411
rect 888 407 892 411
rect 960 407 964 411
rect 1032 407 1036 411
rect 1104 409 1108 413
rect 1176 407 1180 411
rect 1256 407 1260 411
rect 1664 407 1668 411
rect 1720 407 1724 411
rect 1776 407 1780 411
rect 1832 407 1836 411
rect 1888 407 1892 411
rect 1944 407 1948 411
rect 2016 407 2020 411
rect 2104 407 2108 411
rect 2208 407 2212 411
rect 2328 407 2332 411
rect 2456 407 2460 411
rect 2560 407 2564 411
rect 808 379 812 383
rect 1128 379 1132 383
rect 1216 379 1220 383
rect 1688 379 1692 383
rect 1744 379 1748 383
rect 1800 379 1804 383
rect 1856 379 1860 383
rect 1912 379 1916 383
rect 1984 379 1988 383
rect 2072 379 2076 383
rect 2184 379 2188 383
rect 2312 379 2316 383
rect 2448 379 2452 383
rect 2560 379 2564 383
rect 448 375 452 379
rect 504 375 508 379
rect 568 375 572 379
rect 640 375 644 379
rect 720 375 724 379
rect 800 375 804 379
rect 880 375 884 379
rect 960 375 964 379
rect 1040 375 1044 379
rect 1120 375 1124 379
rect 1208 375 1212 379
rect 1296 375 1300 379
rect 1648 343 1652 347
rect 1704 343 1708 347
rect 1760 343 1764 347
rect 1816 343 1820 347
rect 1872 343 1876 347
rect 1944 343 1948 347
rect 2032 343 2036 347
rect 2144 343 2148 347
rect 2272 343 2276 347
rect 2408 343 2412 347
rect 2520 343 2524 347
rect 408 339 412 343
rect 464 339 468 343
rect 528 339 532 343
rect 600 339 604 343
rect 680 339 684 343
rect 760 339 764 343
rect 808 339 812 343
rect 840 339 844 343
rect 920 339 924 343
rect 1000 339 1004 343
rect 1080 339 1084 343
rect 1128 339 1132 343
rect 1168 339 1172 343
rect 1216 339 1220 343
rect 1256 339 1260 343
rect 440 323 444 327
rect 496 323 500 327
rect 552 323 556 327
rect 608 323 612 327
rect 672 323 676 327
rect 744 323 748 327
rect 792 323 796 327
rect 824 323 828 327
rect 904 323 908 327
rect 992 323 996 327
rect 1088 323 1092 327
rect 1192 323 1196 327
rect 1608 323 1612 327
rect 1664 323 1668 327
rect 1720 323 1724 327
rect 1784 323 1788 327
rect 1864 323 1868 327
rect 1944 323 1948 327
rect 2032 323 2036 327
rect 2120 323 2124 327
rect 2208 323 2212 327
rect 2288 323 2292 327
rect 2368 323 2372 327
rect 2456 323 2460 327
rect 2520 323 2524 327
rect 480 287 484 291
rect 536 287 540 291
rect 592 287 596 291
rect 648 287 652 291
rect 712 287 716 291
rect 784 289 788 293
rect 792 291 796 295
rect 864 287 868 291
rect 944 287 948 291
rect 1032 287 1036 291
rect 1128 287 1132 291
rect 1232 287 1236 291
rect 1648 287 1652 291
rect 1704 287 1708 291
rect 1760 287 1764 291
rect 1824 287 1828 291
rect 1904 287 1908 291
rect 1984 287 1988 291
rect 2072 287 2076 291
rect 2160 287 2164 291
rect 2248 287 2252 291
rect 2328 287 2332 291
rect 2408 287 2412 291
rect 2496 287 2500 291
rect 2560 287 2564 291
rect 1992 283 1996 287
rect 1568 259 1572 263
rect 1640 259 1644 263
rect 1720 259 1724 263
rect 1808 259 1812 263
rect 1896 259 1900 263
rect 1984 259 1988 263
rect 320 255 324 259
rect 392 255 396 259
rect 472 255 476 259
rect 560 255 564 259
rect 656 255 660 259
rect 752 255 756 259
rect 856 255 860 259
rect 960 255 964 259
rect 1064 255 1068 259
rect 1176 255 1180 259
rect 1288 255 1292 259
rect 2072 259 2076 263
rect 2152 259 2156 263
rect 2232 259 2236 263
rect 2304 259 2308 263
rect 2368 259 2372 263
rect 2440 259 2444 263
rect 2456 259 2460 263
rect 2504 259 2508 263
rect 2560 259 2564 263
rect 1528 223 1532 227
rect 1600 223 1604 227
rect 1680 223 1684 227
rect 1768 223 1772 227
rect 1856 223 1860 227
rect 1944 223 1948 227
rect 1992 223 1996 227
rect 2032 223 2036 227
rect 2112 223 2116 227
rect 2192 223 2196 227
rect 2264 223 2268 227
rect 2328 223 2332 227
rect 2400 223 2404 227
rect 2456 223 2460 227
rect 2464 223 2468 227
rect 2520 223 2524 227
rect 280 219 284 223
rect 352 219 356 223
rect 432 219 436 223
rect 520 219 524 223
rect 616 219 620 223
rect 712 219 716 223
rect 816 219 820 223
rect 920 219 924 223
rect 1024 219 1028 223
rect 1136 219 1140 223
rect 1248 219 1252 223
rect 1392 211 1396 215
rect 1456 211 1460 215
rect 1536 211 1540 215
rect 1632 211 1636 215
rect 1728 211 1732 215
rect 1832 211 1836 215
rect 1936 211 1940 215
rect 2040 211 2044 215
rect 2144 211 2148 215
rect 2240 211 2244 215
rect 2336 211 2340 215
rect 2440 211 2444 215
rect 2488 211 2492 215
rect 2520 211 2524 215
rect 176 207 180 211
rect 248 207 252 211
rect 336 207 340 211
rect 384 207 388 211
rect 440 207 444 211
rect 544 207 548 211
rect 656 207 660 211
rect 768 207 772 211
rect 888 207 892 211
rect 1008 207 1012 211
rect 1128 207 1132 211
rect 1248 207 1252 211
rect 1432 175 1436 179
rect 1496 175 1500 179
rect 1576 175 1580 179
rect 1672 175 1676 179
rect 1768 175 1772 179
rect 1872 175 1876 179
rect 1976 175 1980 179
rect 2080 175 2084 179
rect 2184 175 2188 179
rect 2280 175 2284 179
rect 2376 175 2380 179
rect 2480 175 2484 179
rect 2488 175 2492 179
rect 2560 175 2564 179
rect 216 171 220 175
rect 288 171 292 175
rect 376 171 380 175
rect 384 171 388 175
rect 480 171 484 175
rect 584 171 588 175
rect 696 171 700 175
rect 808 171 812 175
rect 928 171 932 175
rect 1048 171 1052 175
rect 1168 171 1172 175
rect 1288 171 1292 175
rect 1432 131 1436 135
rect 1488 131 1492 135
rect 1544 131 1548 135
rect 1600 131 1604 135
rect 1664 131 1668 135
rect 1744 131 1748 135
rect 1824 131 1828 135
rect 1904 131 1908 135
rect 1976 131 1980 135
rect 2048 131 2052 135
rect 2112 131 2116 135
rect 2176 131 2180 135
rect 2240 131 2244 135
rect 2304 131 2308 135
rect 2376 131 2380 135
rect 2448 131 2452 135
rect 176 119 180 123
rect 232 119 236 123
rect 288 119 292 123
rect 344 119 348 123
rect 400 119 404 123
rect 456 119 460 123
rect 512 119 516 123
rect 568 119 572 123
rect 624 119 628 123
rect 680 119 684 123
rect 736 119 740 123
rect 792 119 796 123
rect 856 119 860 123
rect 920 119 924 123
rect 984 119 988 123
rect 1048 119 1052 123
rect 1112 119 1116 123
rect 1184 119 1188 123
rect 1248 119 1252 123
rect 1304 119 1308 123
rect 1392 95 1396 99
rect 1448 95 1452 99
rect 1504 95 1508 99
rect 1560 95 1564 99
rect 1624 95 1628 99
rect 1704 95 1708 99
rect 1784 95 1788 99
rect 1864 95 1868 99
rect 1936 95 1940 99
rect 2008 95 2012 99
rect 2072 95 2076 99
rect 2136 95 2140 99
rect 2200 95 2204 99
rect 2264 95 2268 99
rect 2336 95 2340 99
rect 2408 95 2412 99
rect 192 83 196 87
rect 248 83 252 87
rect 304 83 308 87
rect 360 83 364 87
rect 416 83 420 87
rect 472 83 476 87
rect 528 83 532 87
rect 584 83 588 87
rect 640 83 644 87
rect 696 83 700 87
rect 752 83 756 87
rect 816 83 820 87
rect 880 83 884 87
rect 944 83 948 87
rect 1008 83 1012 87
rect 1072 83 1076 87
rect 1144 83 1148 87
rect 1208 83 1212 87
rect 1264 83 1268 87
<< m2 >>
rect 622 2643 628 2644
rect 622 2642 623 2643
rect 545 2640 623 2642
rect 527 2635 533 2636
rect 527 2631 528 2635
rect 532 2634 533 2635
rect 545 2634 547 2640
rect 622 2639 623 2640
rect 627 2639 628 2643
rect 734 2643 740 2644
rect 734 2642 735 2643
rect 622 2638 628 2639
rect 656 2640 735 2642
rect 532 2632 547 2634
rect 582 2635 589 2636
rect 532 2631 533 2632
rect 582 2631 583 2635
rect 588 2631 589 2635
rect 639 2635 645 2636
rect 639 2631 640 2635
rect 644 2634 645 2635
rect 656 2634 658 2640
rect 734 2639 735 2640
rect 739 2639 740 2643
rect 734 2638 740 2639
rect 1622 2639 1628 2640
rect 1622 2638 1623 2639
rect 1544 2636 1623 2638
rect 644 2632 658 2634
rect 694 2635 701 2636
rect 644 2631 645 2632
rect 694 2631 695 2635
rect 700 2631 701 2635
rect 750 2635 757 2636
rect 750 2631 751 2635
rect 756 2631 757 2635
rect 1527 2631 1533 2632
rect 527 2630 533 2631
rect 550 2630 556 2631
rect 582 2630 589 2631
rect 606 2630 612 2631
rect 639 2630 645 2631
rect 662 2630 668 2631
rect 694 2630 701 2631
rect 718 2630 724 2631
rect 750 2630 757 2631
rect 774 2630 780 2631
rect 550 2626 551 2630
rect 555 2626 556 2630
rect 550 2625 556 2626
rect 606 2626 607 2630
rect 611 2626 612 2630
rect 606 2625 612 2626
rect 662 2626 663 2630
rect 667 2626 668 2630
rect 662 2625 668 2626
rect 718 2626 719 2630
rect 723 2626 724 2630
rect 718 2625 724 2626
rect 774 2626 775 2630
rect 779 2626 780 2630
rect 1527 2627 1528 2631
rect 1532 2630 1533 2631
rect 1544 2630 1546 2636
rect 1622 2635 1623 2636
rect 1627 2635 1628 2639
rect 1734 2639 1740 2640
rect 1734 2638 1735 2639
rect 1622 2634 1628 2635
rect 1656 2636 1735 2638
rect 1532 2628 1546 2630
rect 1582 2631 1589 2632
rect 1532 2627 1533 2628
rect 1582 2627 1583 2631
rect 1588 2627 1589 2631
rect 1639 2631 1645 2632
rect 1639 2627 1640 2631
rect 1644 2630 1645 2631
rect 1656 2630 1658 2636
rect 1734 2635 1735 2636
rect 1739 2635 1740 2639
rect 1838 2639 1844 2640
rect 1838 2638 1839 2639
rect 1734 2634 1740 2635
rect 1768 2636 1839 2638
rect 1644 2628 1658 2630
rect 1694 2631 1701 2632
rect 1644 2627 1645 2628
rect 1694 2627 1695 2631
rect 1700 2627 1701 2631
rect 1751 2631 1757 2632
rect 1751 2627 1752 2631
rect 1756 2630 1757 2631
rect 1768 2630 1770 2636
rect 1838 2635 1839 2636
rect 1843 2635 1844 2639
rect 1958 2639 1964 2640
rect 1958 2638 1959 2639
rect 1838 2634 1844 2635
rect 1881 2636 1959 2638
rect 1756 2628 1770 2630
rect 1806 2631 1813 2632
rect 1756 2627 1757 2628
rect 1806 2627 1807 2631
rect 1812 2627 1813 2631
rect 1863 2631 1869 2632
rect 1863 2627 1864 2631
rect 1868 2630 1869 2631
rect 1881 2630 1883 2636
rect 1958 2635 1959 2636
rect 1963 2635 1964 2639
rect 2182 2639 2188 2640
rect 2182 2638 2183 2639
rect 1958 2634 1964 2635
rect 1999 2636 2183 2638
rect 1999 2634 2001 2636
rect 2182 2635 2183 2636
rect 2187 2635 2188 2639
rect 2182 2634 2188 2635
rect 1988 2632 2001 2634
rect 1868 2628 1883 2630
rect 1918 2631 1925 2632
rect 1868 2627 1869 2628
rect 1918 2627 1919 2631
rect 1924 2627 1925 2631
rect 1975 2631 1981 2632
rect 1975 2627 1976 2631
rect 1980 2630 1981 2631
rect 1988 2630 1990 2632
rect 1980 2628 1990 2630
rect 2026 2631 2037 2632
rect 1980 2627 1981 2628
rect 2026 2627 2027 2631
rect 2031 2627 2032 2631
rect 2036 2627 2037 2631
rect 2074 2631 2080 2632
rect 2074 2627 2075 2631
rect 2079 2630 2080 2631
rect 2087 2631 2093 2632
rect 2087 2630 2088 2631
rect 2079 2628 2088 2630
rect 2079 2627 2080 2628
rect 1527 2626 1533 2627
rect 1550 2626 1556 2627
rect 1582 2626 1589 2627
rect 1606 2626 1612 2627
rect 1639 2626 1645 2627
rect 1662 2626 1668 2627
rect 1694 2626 1701 2627
rect 1718 2626 1724 2627
rect 1751 2626 1757 2627
rect 1774 2626 1780 2627
rect 1806 2626 1813 2627
rect 1830 2626 1836 2627
rect 1863 2626 1869 2627
rect 1886 2626 1892 2627
rect 1918 2626 1925 2627
rect 1942 2626 1948 2627
rect 1975 2626 1981 2627
rect 1998 2626 2004 2627
rect 2026 2626 2037 2627
rect 2054 2626 2060 2627
rect 2074 2626 2080 2627
rect 2087 2627 2088 2628
rect 2092 2627 2093 2631
rect 2130 2631 2136 2632
rect 2130 2627 2131 2631
rect 2135 2630 2136 2631
rect 2143 2631 2149 2632
rect 2143 2630 2144 2631
rect 2135 2628 2144 2630
rect 2135 2627 2136 2628
rect 2087 2626 2093 2627
rect 2110 2626 2116 2627
rect 2130 2626 2136 2627
rect 2143 2627 2144 2628
rect 2148 2627 2149 2631
rect 2143 2626 2149 2627
rect 2166 2626 2172 2627
rect 774 2625 780 2626
rect 1550 2622 1551 2626
rect 1555 2622 1556 2626
rect 110 2621 116 2622
rect 110 2617 111 2621
rect 115 2617 116 2621
rect 110 2616 116 2617
rect 1326 2621 1332 2622
rect 1550 2621 1556 2622
rect 1606 2622 1607 2626
rect 1611 2622 1612 2626
rect 1606 2621 1612 2622
rect 1662 2622 1663 2626
rect 1667 2622 1668 2626
rect 1662 2621 1668 2622
rect 1718 2622 1719 2626
rect 1723 2622 1724 2626
rect 1718 2621 1724 2622
rect 1774 2622 1775 2626
rect 1779 2622 1780 2626
rect 1774 2621 1780 2622
rect 1830 2622 1831 2626
rect 1835 2622 1836 2626
rect 1830 2621 1836 2622
rect 1886 2622 1887 2626
rect 1891 2622 1892 2626
rect 1886 2621 1892 2622
rect 1942 2622 1943 2626
rect 1947 2622 1948 2626
rect 1942 2621 1948 2622
rect 1998 2622 1999 2626
rect 2003 2622 2004 2626
rect 1998 2621 2004 2622
rect 2054 2622 2055 2626
rect 2059 2622 2060 2626
rect 2054 2621 2060 2622
rect 2110 2622 2111 2626
rect 2115 2622 2116 2626
rect 2110 2621 2116 2622
rect 2166 2622 2167 2626
rect 2171 2622 2172 2626
rect 2166 2621 2172 2622
rect 1326 2617 1327 2621
rect 1331 2617 1332 2621
rect 1326 2616 1332 2617
rect 1366 2617 1372 2618
rect 1366 2613 1367 2617
rect 1371 2613 1372 2617
rect 1366 2612 1372 2613
rect 2582 2617 2588 2618
rect 2582 2613 2583 2617
rect 2587 2613 2588 2617
rect 2582 2612 2588 2613
rect 582 2611 588 2612
rect 582 2607 583 2611
rect 587 2610 588 2611
rect 694 2611 700 2612
rect 587 2608 674 2610
rect 587 2607 588 2608
rect 582 2606 588 2607
rect 110 2604 116 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 534 2603 540 2604
rect 534 2599 535 2603
rect 539 2599 540 2603
rect 590 2603 596 2604
rect 534 2598 540 2599
rect 558 2599 564 2600
rect 558 2595 559 2599
rect 563 2598 564 2599
rect 567 2599 573 2600
rect 567 2598 568 2599
rect 563 2596 568 2598
rect 563 2595 564 2596
rect 558 2594 564 2595
rect 567 2595 568 2596
rect 572 2595 573 2599
rect 590 2599 591 2603
rect 595 2599 596 2603
rect 646 2603 652 2604
rect 590 2598 596 2599
rect 622 2599 629 2600
rect 567 2594 573 2595
rect 622 2595 623 2599
rect 628 2595 629 2599
rect 646 2599 647 2603
rect 651 2599 652 2603
rect 646 2598 652 2599
rect 672 2598 674 2608
rect 694 2607 695 2611
rect 699 2610 700 2611
rect 699 2608 786 2610
rect 699 2607 700 2608
rect 694 2606 700 2607
rect 702 2603 708 2604
rect 679 2599 685 2600
rect 679 2598 680 2599
rect 672 2596 680 2598
rect 622 2594 629 2595
rect 679 2595 680 2596
rect 684 2595 685 2599
rect 702 2599 703 2603
rect 707 2599 708 2603
rect 758 2603 764 2604
rect 702 2598 708 2599
rect 734 2599 741 2600
rect 679 2594 685 2595
rect 734 2595 735 2599
rect 740 2595 741 2599
rect 758 2599 759 2603
rect 763 2599 764 2603
rect 758 2598 764 2599
rect 784 2598 786 2608
rect 1582 2607 1588 2608
rect 1326 2604 1332 2605
rect 1326 2600 1327 2604
rect 1331 2600 1332 2604
rect 1582 2603 1583 2607
rect 1587 2606 1588 2607
rect 1694 2607 1700 2608
rect 1587 2604 1674 2606
rect 1587 2603 1588 2604
rect 1582 2602 1588 2603
rect 791 2599 797 2600
rect 1326 2599 1332 2600
rect 1366 2600 1372 2601
rect 791 2598 792 2599
rect 784 2596 792 2598
rect 734 2594 741 2595
rect 791 2595 792 2596
rect 796 2595 797 2599
rect 1366 2596 1367 2600
rect 1371 2596 1372 2600
rect 1366 2595 1372 2596
rect 1534 2599 1540 2600
rect 1534 2595 1535 2599
rect 1539 2595 1540 2599
rect 1590 2599 1596 2600
rect 791 2594 797 2595
rect 1534 2594 1540 2595
rect 1567 2595 1573 2596
rect 1567 2594 1568 2595
rect 1544 2592 1568 2594
rect 1446 2591 1452 2592
rect 1446 2587 1447 2591
rect 1451 2590 1452 2591
rect 1544 2590 1546 2592
rect 1567 2591 1568 2592
rect 1572 2591 1573 2595
rect 1590 2595 1591 2599
rect 1595 2595 1596 2599
rect 1646 2599 1652 2600
rect 1590 2594 1596 2595
rect 1622 2595 1629 2596
rect 1567 2590 1573 2591
rect 1622 2591 1623 2595
rect 1628 2591 1629 2595
rect 1646 2595 1647 2599
rect 1651 2595 1652 2599
rect 1646 2594 1652 2595
rect 1672 2594 1674 2604
rect 1694 2603 1695 2607
rect 1699 2606 1700 2607
rect 1806 2607 1812 2608
rect 1699 2604 1786 2606
rect 1699 2603 1700 2604
rect 1694 2602 1700 2603
rect 1702 2599 1708 2600
rect 1679 2595 1685 2596
rect 1679 2594 1680 2595
rect 1672 2592 1680 2594
rect 1622 2590 1629 2591
rect 1679 2591 1680 2592
rect 1684 2591 1685 2595
rect 1702 2595 1703 2599
rect 1707 2595 1708 2599
rect 1758 2599 1764 2600
rect 1702 2594 1708 2595
rect 1734 2595 1741 2596
rect 1679 2590 1685 2591
rect 1734 2591 1735 2595
rect 1740 2591 1741 2595
rect 1758 2595 1759 2599
rect 1763 2595 1764 2599
rect 1758 2594 1764 2595
rect 1784 2594 1786 2604
rect 1806 2603 1807 2607
rect 1811 2606 1812 2607
rect 1918 2607 1924 2608
rect 1811 2604 1898 2606
rect 1811 2603 1812 2604
rect 1806 2602 1812 2603
rect 1814 2599 1820 2600
rect 1791 2595 1797 2596
rect 1791 2594 1792 2595
rect 1784 2592 1792 2594
rect 1734 2590 1741 2591
rect 1791 2591 1792 2592
rect 1796 2591 1797 2595
rect 1814 2595 1815 2599
rect 1819 2595 1820 2599
rect 1870 2599 1876 2600
rect 1814 2594 1820 2595
rect 1838 2595 1844 2596
rect 1791 2590 1797 2591
rect 1838 2591 1839 2595
rect 1843 2594 1844 2595
rect 1847 2595 1853 2596
rect 1847 2594 1848 2595
rect 1843 2592 1848 2594
rect 1843 2591 1844 2592
rect 1838 2590 1844 2591
rect 1847 2591 1848 2592
rect 1852 2591 1853 2595
rect 1870 2595 1871 2599
rect 1875 2595 1876 2599
rect 1870 2594 1876 2595
rect 1896 2594 1898 2604
rect 1918 2603 1919 2607
rect 1923 2606 1924 2607
rect 1923 2604 2010 2606
rect 1923 2603 1924 2604
rect 1918 2602 1924 2603
rect 1926 2599 1932 2600
rect 1903 2595 1909 2596
rect 1903 2594 1904 2595
rect 1896 2592 1904 2594
rect 1847 2590 1853 2591
rect 1903 2591 1904 2592
rect 1908 2591 1909 2595
rect 1926 2595 1927 2599
rect 1931 2595 1932 2599
rect 1982 2599 1988 2600
rect 1926 2594 1932 2595
rect 1958 2595 1965 2596
rect 1903 2590 1909 2591
rect 1958 2591 1959 2595
rect 1964 2591 1965 2595
rect 1982 2595 1983 2599
rect 1987 2595 1988 2599
rect 1982 2594 1988 2595
rect 2008 2594 2010 2604
rect 2582 2600 2588 2601
rect 2038 2599 2044 2600
rect 2015 2595 2021 2596
rect 2015 2594 2016 2595
rect 2008 2592 2016 2594
rect 1958 2590 1965 2591
rect 2015 2591 2016 2592
rect 2020 2591 2021 2595
rect 2038 2595 2039 2599
rect 2043 2595 2044 2599
rect 2094 2599 2100 2600
rect 2038 2594 2044 2595
rect 2071 2595 2080 2596
rect 2015 2590 2021 2591
rect 2071 2591 2072 2595
rect 2079 2591 2080 2595
rect 2094 2595 2095 2599
rect 2099 2595 2100 2599
rect 2150 2599 2156 2600
rect 2094 2594 2100 2595
rect 2127 2595 2136 2596
rect 2071 2590 2080 2591
rect 2127 2591 2128 2595
rect 2135 2591 2136 2595
rect 2150 2595 2151 2599
rect 2155 2595 2156 2599
rect 2582 2596 2583 2600
rect 2587 2596 2588 2600
rect 2150 2594 2156 2595
rect 2182 2595 2189 2596
rect 2582 2595 2588 2596
rect 2127 2590 2136 2591
rect 2182 2591 2183 2595
rect 2188 2591 2189 2595
rect 2182 2590 2189 2591
rect 1451 2588 1546 2590
rect 1451 2587 1452 2588
rect 1446 2586 1452 2587
rect 238 2579 244 2580
rect 238 2575 239 2579
rect 243 2578 244 2579
rect 526 2579 532 2580
rect 243 2576 410 2578
rect 243 2575 244 2576
rect 238 2574 244 2575
rect 247 2571 253 2572
rect 214 2569 220 2570
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 247 2567 248 2571
rect 252 2570 253 2571
rect 262 2571 268 2572
rect 262 2570 263 2571
rect 252 2568 263 2570
rect 252 2567 253 2568
rect 247 2566 253 2567
rect 262 2567 263 2568
rect 267 2567 268 2571
rect 303 2571 309 2572
rect 262 2566 268 2567
rect 270 2569 276 2570
rect 214 2564 220 2565
rect 270 2565 271 2569
rect 275 2565 276 2569
rect 303 2567 304 2571
rect 308 2570 309 2571
rect 318 2571 324 2572
rect 318 2570 319 2571
rect 308 2568 319 2570
rect 308 2567 309 2568
rect 303 2566 309 2567
rect 318 2567 319 2568
rect 323 2567 324 2571
rect 354 2571 365 2572
rect 318 2566 324 2567
rect 326 2569 332 2570
rect 270 2564 276 2565
rect 326 2565 327 2569
rect 331 2565 332 2569
rect 354 2567 355 2571
rect 359 2567 360 2571
rect 364 2567 365 2571
rect 408 2570 410 2576
rect 423 2575 429 2576
rect 415 2571 421 2572
rect 415 2570 416 2571
rect 354 2566 365 2567
rect 382 2569 388 2570
rect 326 2564 332 2565
rect 382 2565 383 2569
rect 387 2565 388 2569
rect 408 2568 416 2570
rect 415 2567 416 2568
rect 420 2567 421 2571
rect 423 2571 424 2575
rect 428 2574 429 2575
rect 479 2575 485 2576
rect 428 2572 466 2574
rect 428 2571 429 2572
rect 423 2570 429 2571
rect 464 2570 466 2572
rect 471 2571 477 2572
rect 471 2570 472 2571
rect 415 2566 421 2567
rect 438 2569 444 2570
rect 382 2564 388 2565
rect 438 2565 439 2569
rect 443 2565 444 2569
rect 464 2568 472 2570
rect 471 2567 472 2568
rect 476 2567 477 2571
rect 479 2571 480 2575
rect 484 2574 485 2575
rect 526 2575 527 2579
rect 531 2578 532 2579
rect 686 2579 692 2580
rect 531 2576 634 2578
rect 531 2575 532 2576
rect 526 2574 532 2575
rect 484 2572 522 2574
rect 484 2571 485 2572
rect 479 2570 485 2571
rect 520 2570 522 2572
rect 527 2571 533 2572
rect 527 2570 528 2571
rect 471 2566 477 2567
rect 494 2569 500 2570
rect 438 2564 444 2565
rect 494 2565 495 2569
rect 499 2565 500 2569
rect 520 2568 528 2570
rect 527 2567 528 2568
rect 532 2567 533 2571
rect 583 2571 589 2572
rect 527 2566 533 2567
rect 550 2569 556 2570
rect 494 2564 500 2565
rect 550 2565 551 2569
rect 555 2565 556 2569
rect 583 2567 584 2571
rect 588 2570 589 2571
rect 598 2571 604 2572
rect 598 2570 599 2571
rect 588 2568 599 2570
rect 588 2567 589 2568
rect 583 2566 589 2567
rect 598 2567 599 2568
rect 603 2567 604 2571
rect 632 2570 634 2576
rect 686 2575 687 2579
rect 691 2578 692 2579
rect 974 2579 980 2580
rect 691 2576 802 2578
rect 691 2575 692 2576
rect 686 2574 692 2575
rect 639 2571 645 2572
rect 639 2570 640 2571
rect 598 2566 604 2567
rect 606 2569 612 2570
rect 550 2564 556 2565
rect 606 2565 607 2569
rect 611 2565 612 2569
rect 632 2568 640 2570
rect 639 2567 640 2568
rect 644 2567 645 2571
rect 695 2571 701 2572
rect 639 2566 645 2567
rect 662 2569 668 2570
rect 606 2564 612 2565
rect 662 2565 663 2569
rect 667 2565 668 2569
rect 695 2567 696 2571
rect 700 2570 701 2571
rect 710 2571 716 2572
rect 710 2570 711 2571
rect 700 2568 711 2570
rect 700 2567 701 2568
rect 695 2566 701 2567
rect 710 2567 711 2568
rect 715 2567 716 2571
rect 750 2571 757 2572
rect 710 2566 716 2567
rect 718 2569 724 2570
rect 662 2564 668 2565
rect 718 2565 719 2569
rect 723 2565 724 2569
rect 750 2567 751 2571
rect 756 2567 757 2571
rect 800 2570 802 2576
rect 815 2575 821 2576
rect 807 2571 813 2572
rect 807 2570 808 2571
rect 750 2566 757 2567
rect 774 2569 780 2570
rect 718 2564 724 2565
rect 774 2565 775 2569
rect 779 2565 780 2569
rect 800 2568 808 2570
rect 807 2567 808 2568
rect 812 2567 813 2571
rect 815 2571 816 2575
rect 820 2574 821 2575
rect 871 2575 877 2576
rect 820 2572 858 2574
rect 820 2571 821 2572
rect 815 2570 821 2571
rect 856 2570 858 2572
rect 863 2571 869 2572
rect 863 2570 864 2571
rect 807 2566 813 2567
rect 830 2569 836 2570
rect 774 2564 780 2565
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 856 2568 864 2570
rect 863 2567 864 2568
rect 868 2567 869 2571
rect 871 2571 872 2575
rect 876 2574 877 2575
rect 927 2575 933 2576
rect 876 2572 914 2574
rect 876 2571 877 2572
rect 871 2570 877 2571
rect 912 2570 914 2572
rect 919 2571 925 2572
rect 919 2570 920 2571
rect 863 2566 869 2567
rect 886 2569 892 2570
rect 830 2564 836 2565
rect 886 2565 887 2569
rect 891 2565 892 2569
rect 912 2568 920 2570
rect 919 2567 920 2568
rect 924 2567 925 2571
rect 927 2571 928 2575
rect 932 2574 933 2575
rect 974 2575 975 2579
rect 979 2578 980 2579
rect 979 2576 1138 2578
rect 979 2575 980 2576
rect 974 2574 980 2575
rect 932 2572 970 2574
rect 932 2571 933 2572
rect 927 2570 933 2571
rect 968 2570 970 2572
rect 975 2571 981 2572
rect 975 2570 976 2571
rect 919 2566 925 2567
rect 942 2569 948 2570
rect 886 2564 892 2565
rect 942 2565 943 2569
rect 947 2565 948 2569
rect 968 2568 976 2570
rect 975 2567 976 2568
rect 980 2567 981 2571
rect 1031 2571 1037 2572
rect 975 2566 981 2567
rect 998 2569 1004 2570
rect 942 2564 948 2565
rect 998 2565 999 2569
rect 1003 2565 1004 2569
rect 1031 2567 1032 2571
rect 1036 2570 1037 2571
rect 1046 2571 1052 2572
rect 1046 2570 1047 2571
rect 1036 2568 1047 2570
rect 1036 2567 1037 2568
rect 1031 2566 1037 2567
rect 1046 2567 1047 2568
rect 1051 2567 1052 2571
rect 1087 2571 1093 2572
rect 1046 2566 1052 2567
rect 1054 2569 1060 2570
rect 998 2564 1004 2565
rect 1054 2565 1055 2569
rect 1059 2565 1060 2569
rect 1087 2567 1088 2571
rect 1092 2570 1093 2571
rect 1102 2571 1108 2572
rect 1102 2570 1103 2571
rect 1092 2568 1103 2570
rect 1092 2567 1093 2568
rect 1087 2566 1093 2567
rect 1102 2567 1103 2568
rect 1107 2567 1108 2571
rect 1136 2570 1138 2576
rect 1143 2571 1149 2572
rect 1143 2570 1144 2571
rect 1102 2566 1108 2567
rect 1110 2569 1116 2570
rect 1054 2564 1060 2565
rect 1110 2565 1111 2569
rect 1115 2565 1116 2569
rect 1136 2568 1144 2570
rect 1143 2567 1144 2568
rect 1148 2567 1149 2571
rect 2070 2571 2076 2572
rect 1143 2566 1149 2567
rect 1326 2568 1332 2569
rect 1110 2564 1116 2565
rect 1326 2564 1327 2568
rect 1331 2564 1332 2568
rect 1471 2567 1477 2568
rect 1438 2565 1444 2566
rect 110 2563 116 2564
rect 1326 2563 1332 2564
rect 1366 2564 1372 2565
rect 1366 2560 1367 2564
rect 1371 2560 1372 2564
rect 1438 2561 1439 2565
rect 1443 2561 1444 2565
rect 1471 2563 1472 2567
rect 1476 2566 1477 2567
rect 1534 2567 1540 2568
rect 1534 2566 1535 2567
rect 1476 2564 1535 2566
rect 1476 2563 1477 2564
rect 1471 2562 1477 2563
rect 1534 2563 1535 2564
rect 1539 2563 1540 2567
rect 1575 2567 1581 2568
rect 1534 2562 1540 2563
rect 1542 2565 1548 2566
rect 1438 2560 1444 2561
rect 1542 2561 1543 2565
rect 1547 2561 1548 2565
rect 1575 2563 1576 2567
rect 1580 2566 1581 2567
rect 1646 2567 1652 2568
rect 1646 2566 1647 2567
rect 1580 2564 1647 2566
rect 1580 2563 1581 2564
rect 1575 2562 1581 2563
rect 1646 2563 1647 2564
rect 1651 2563 1652 2567
rect 1687 2567 1693 2568
rect 1646 2562 1652 2563
rect 1654 2565 1660 2566
rect 1542 2560 1548 2561
rect 1654 2561 1655 2565
rect 1659 2561 1660 2565
rect 1687 2563 1688 2567
rect 1692 2566 1693 2567
rect 1758 2567 1764 2568
rect 1758 2566 1759 2567
rect 1692 2564 1759 2566
rect 1692 2563 1693 2564
rect 1687 2562 1693 2563
rect 1758 2563 1759 2564
rect 1763 2563 1764 2567
rect 1799 2567 1805 2568
rect 1758 2562 1764 2563
rect 1766 2565 1772 2566
rect 1654 2560 1660 2561
rect 1766 2561 1767 2565
rect 1771 2561 1772 2565
rect 1799 2563 1800 2567
rect 1804 2566 1805 2567
rect 1870 2567 1876 2568
rect 1870 2566 1871 2567
rect 1804 2564 1871 2566
rect 1804 2563 1805 2564
rect 1799 2562 1805 2563
rect 1870 2563 1871 2564
rect 1875 2563 1876 2567
rect 1902 2567 1908 2568
rect 1870 2562 1876 2563
rect 1878 2565 1884 2566
rect 1766 2560 1772 2561
rect 1878 2561 1879 2565
rect 1883 2561 1884 2565
rect 1902 2563 1903 2567
rect 1907 2566 1908 2567
rect 1911 2567 1917 2568
rect 1911 2566 1912 2567
rect 1907 2564 1912 2566
rect 1907 2563 1908 2564
rect 1902 2562 1908 2563
rect 1911 2563 1912 2564
rect 1916 2563 1917 2567
rect 2023 2567 2032 2568
rect 1911 2562 1917 2563
rect 1990 2565 1996 2566
rect 1878 2560 1884 2561
rect 1990 2561 1991 2565
rect 1995 2561 1996 2565
rect 2023 2563 2024 2567
rect 2031 2563 2032 2567
rect 2070 2567 2071 2571
rect 2075 2570 2076 2571
rect 2151 2571 2157 2572
rect 2075 2568 2138 2570
rect 2075 2567 2076 2568
rect 2070 2566 2076 2567
rect 2136 2566 2138 2568
rect 2143 2567 2149 2568
rect 2143 2566 2144 2567
rect 2023 2562 2032 2563
rect 2110 2565 2116 2566
rect 1990 2560 1996 2561
rect 2110 2561 2111 2565
rect 2115 2561 2116 2565
rect 2136 2564 2144 2566
rect 2143 2563 2144 2564
rect 2148 2563 2149 2567
rect 2151 2567 2152 2571
rect 2156 2570 2157 2571
rect 2271 2571 2277 2572
rect 2156 2568 2258 2570
rect 2156 2567 2157 2568
rect 2151 2566 2157 2567
rect 2256 2566 2258 2568
rect 2263 2567 2269 2568
rect 2263 2566 2264 2567
rect 2143 2562 2149 2563
rect 2230 2565 2236 2566
rect 2110 2560 2116 2561
rect 2230 2561 2231 2565
rect 2235 2561 2236 2565
rect 2256 2564 2264 2566
rect 2263 2563 2264 2564
rect 2268 2563 2269 2567
rect 2271 2567 2272 2571
rect 2276 2570 2277 2571
rect 2276 2568 2378 2570
rect 2276 2567 2277 2568
rect 2271 2566 2277 2567
rect 2376 2566 2378 2568
rect 2383 2567 2389 2568
rect 2383 2566 2384 2567
rect 2263 2562 2269 2563
rect 2350 2565 2356 2566
rect 2230 2560 2236 2561
rect 2350 2561 2351 2565
rect 2355 2561 2356 2565
rect 2376 2564 2384 2566
rect 2383 2563 2384 2564
rect 2388 2563 2389 2567
rect 2383 2562 2389 2563
rect 2582 2564 2588 2565
rect 2350 2560 2356 2561
rect 2582 2560 2583 2564
rect 2587 2560 2588 2564
rect 1366 2559 1372 2560
rect 2582 2559 2588 2560
rect 110 2551 116 2552
rect 110 2547 111 2551
rect 115 2547 116 2551
rect 110 2546 116 2547
rect 1326 2551 1332 2552
rect 1326 2547 1327 2551
rect 1331 2547 1332 2551
rect 1326 2546 1332 2547
rect 1366 2547 1372 2548
rect 1366 2543 1367 2547
rect 1371 2543 1372 2547
rect 230 2542 236 2543
rect 230 2538 231 2542
rect 235 2538 236 2542
rect 230 2537 236 2538
rect 286 2542 292 2543
rect 286 2538 287 2542
rect 291 2538 292 2542
rect 286 2537 292 2538
rect 342 2542 348 2543
rect 342 2538 343 2542
rect 347 2538 348 2542
rect 342 2537 348 2538
rect 398 2542 404 2543
rect 398 2538 399 2542
rect 403 2538 404 2542
rect 398 2537 404 2538
rect 454 2542 460 2543
rect 454 2538 455 2542
rect 459 2538 460 2542
rect 454 2537 460 2538
rect 510 2542 516 2543
rect 510 2538 511 2542
rect 515 2538 516 2542
rect 510 2537 516 2538
rect 566 2542 572 2543
rect 566 2538 567 2542
rect 571 2538 572 2542
rect 566 2537 572 2538
rect 622 2542 628 2543
rect 622 2538 623 2542
rect 627 2538 628 2542
rect 622 2537 628 2538
rect 678 2542 684 2543
rect 678 2538 679 2542
rect 683 2538 684 2542
rect 678 2537 684 2538
rect 734 2542 740 2543
rect 734 2538 735 2542
rect 739 2538 740 2542
rect 734 2537 740 2538
rect 790 2542 796 2543
rect 790 2538 791 2542
rect 795 2538 796 2542
rect 790 2537 796 2538
rect 846 2542 852 2543
rect 846 2538 847 2542
rect 851 2538 852 2542
rect 846 2537 852 2538
rect 902 2542 908 2543
rect 902 2538 903 2542
rect 907 2538 908 2542
rect 902 2537 908 2538
rect 958 2542 964 2543
rect 958 2538 959 2542
rect 963 2538 964 2542
rect 958 2537 964 2538
rect 1014 2542 1020 2543
rect 1014 2538 1015 2542
rect 1019 2538 1020 2542
rect 1014 2537 1020 2538
rect 1070 2542 1076 2543
rect 1070 2538 1071 2542
rect 1075 2538 1076 2542
rect 1070 2537 1076 2538
rect 1126 2542 1132 2543
rect 1366 2542 1372 2543
rect 2582 2547 2588 2548
rect 2582 2543 2583 2547
rect 2587 2543 2588 2547
rect 2582 2542 2588 2543
rect 1126 2538 1127 2542
rect 1131 2538 1132 2542
rect 1126 2537 1132 2538
rect 1454 2538 1460 2539
rect 207 2535 213 2536
rect 207 2531 208 2535
rect 212 2534 213 2535
rect 238 2535 244 2536
rect 238 2534 239 2535
rect 212 2532 239 2534
rect 212 2531 213 2532
rect 207 2530 213 2531
rect 238 2531 239 2532
rect 243 2531 244 2535
rect 238 2530 244 2531
rect 262 2535 269 2536
rect 262 2531 263 2535
rect 268 2531 269 2535
rect 262 2530 269 2531
rect 318 2535 325 2536
rect 318 2531 319 2535
rect 324 2531 325 2535
rect 318 2530 325 2531
rect 375 2535 381 2536
rect 375 2531 376 2535
rect 380 2534 381 2535
rect 423 2535 429 2536
rect 423 2534 424 2535
rect 380 2532 424 2534
rect 380 2531 381 2532
rect 375 2530 381 2531
rect 423 2531 424 2532
rect 428 2531 429 2535
rect 423 2530 429 2531
rect 431 2535 437 2536
rect 431 2531 432 2535
rect 436 2534 437 2535
rect 479 2535 485 2536
rect 479 2534 480 2535
rect 436 2532 480 2534
rect 436 2531 437 2532
rect 431 2530 437 2531
rect 479 2531 480 2532
rect 484 2531 485 2535
rect 479 2530 485 2531
rect 487 2535 493 2536
rect 487 2531 488 2535
rect 492 2534 493 2535
rect 526 2535 532 2536
rect 526 2534 527 2535
rect 492 2532 527 2534
rect 492 2531 493 2532
rect 487 2530 493 2531
rect 526 2531 527 2532
rect 531 2531 532 2535
rect 526 2530 532 2531
rect 543 2535 549 2536
rect 543 2531 544 2535
rect 548 2534 549 2535
rect 558 2535 564 2536
rect 558 2534 559 2535
rect 548 2532 559 2534
rect 548 2531 549 2532
rect 543 2530 549 2531
rect 558 2531 559 2532
rect 563 2531 564 2535
rect 558 2530 564 2531
rect 598 2535 605 2536
rect 598 2531 599 2535
rect 604 2531 605 2535
rect 598 2530 605 2531
rect 655 2535 661 2536
rect 655 2531 656 2535
rect 660 2534 661 2535
rect 686 2535 692 2536
rect 686 2534 687 2535
rect 660 2532 687 2534
rect 660 2531 661 2532
rect 655 2530 661 2531
rect 686 2531 687 2532
rect 691 2531 692 2535
rect 686 2530 692 2531
rect 710 2535 717 2536
rect 710 2531 711 2535
rect 716 2531 717 2535
rect 710 2530 717 2531
rect 767 2535 773 2536
rect 767 2531 768 2535
rect 772 2534 773 2535
rect 815 2535 821 2536
rect 815 2534 816 2535
rect 772 2532 816 2534
rect 772 2531 773 2532
rect 767 2530 773 2531
rect 815 2531 816 2532
rect 820 2531 821 2535
rect 815 2530 821 2531
rect 823 2535 829 2536
rect 823 2531 824 2535
rect 828 2534 829 2535
rect 871 2535 877 2536
rect 871 2534 872 2535
rect 828 2532 872 2534
rect 828 2531 829 2532
rect 823 2530 829 2531
rect 871 2531 872 2532
rect 876 2531 877 2535
rect 871 2530 877 2531
rect 879 2535 885 2536
rect 879 2531 880 2535
rect 884 2534 885 2535
rect 927 2535 933 2536
rect 927 2534 928 2535
rect 884 2532 928 2534
rect 884 2531 885 2532
rect 879 2530 885 2531
rect 927 2531 928 2532
rect 932 2531 933 2535
rect 927 2530 933 2531
rect 935 2535 941 2536
rect 935 2531 936 2535
rect 940 2534 941 2535
rect 974 2535 980 2536
rect 974 2534 975 2535
rect 940 2532 975 2534
rect 940 2531 941 2532
rect 935 2530 941 2531
rect 974 2531 975 2532
rect 979 2531 980 2535
rect 974 2530 980 2531
rect 983 2535 989 2536
rect 983 2531 984 2535
rect 988 2534 989 2535
rect 991 2535 997 2536
rect 991 2534 992 2535
rect 988 2532 992 2534
rect 988 2531 989 2532
rect 983 2530 989 2531
rect 991 2531 992 2532
rect 996 2531 997 2535
rect 991 2530 997 2531
rect 1046 2535 1053 2536
rect 1046 2531 1047 2535
rect 1052 2531 1053 2535
rect 1046 2530 1053 2531
rect 1102 2535 1109 2536
rect 1102 2531 1103 2535
rect 1108 2531 1109 2535
rect 1454 2534 1455 2538
rect 1459 2534 1460 2538
rect 1454 2533 1460 2534
rect 1558 2538 1564 2539
rect 1558 2534 1559 2538
rect 1563 2534 1564 2538
rect 1558 2533 1564 2534
rect 1670 2538 1676 2539
rect 1670 2534 1671 2538
rect 1675 2534 1676 2538
rect 1670 2533 1676 2534
rect 1782 2538 1788 2539
rect 1782 2534 1783 2538
rect 1787 2534 1788 2538
rect 1782 2533 1788 2534
rect 1894 2538 1900 2539
rect 1894 2534 1895 2538
rect 1899 2534 1900 2538
rect 1894 2533 1900 2534
rect 2006 2538 2012 2539
rect 2006 2534 2007 2538
rect 2011 2534 2012 2538
rect 2006 2533 2012 2534
rect 2126 2538 2132 2539
rect 2126 2534 2127 2538
rect 2131 2534 2132 2538
rect 2126 2533 2132 2534
rect 2246 2538 2252 2539
rect 2246 2534 2247 2538
rect 2251 2534 2252 2538
rect 2246 2533 2252 2534
rect 2366 2538 2372 2539
rect 2366 2534 2367 2538
rect 2371 2534 2372 2538
rect 2366 2533 2372 2534
rect 1102 2530 1109 2531
rect 1431 2531 1437 2532
rect 1022 2527 1028 2528
rect 1022 2526 1023 2527
rect 864 2524 1023 2526
rect 354 2523 360 2524
rect 354 2522 355 2523
rect 343 2521 355 2522
rect 343 2517 344 2521
rect 348 2520 355 2521
rect 348 2517 349 2520
rect 354 2519 355 2520
rect 359 2519 360 2523
rect 354 2518 360 2519
rect 386 2519 392 2520
rect 343 2516 349 2517
rect 386 2515 387 2519
rect 391 2518 392 2519
rect 399 2519 405 2520
rect 399 2518 400 2519
rect 391 2516 400 2518
rect 391 2515 392 2516
rect 366 2514 372 2515
rect 386 2514 392 2515
rect 399 2515 400 2516
rect 404 2515 405 2519
rect 442 2519 448 2520
rect 442 2515 443 2519
rect 447 2518 448 2519
rect 463 2519 469 2520
rect 463 2518 464 2519
rect 447 2516 464 2518
rect 447 2515 448 2516
rect 399 2514 405 2515
rect 422 2514 428 2515
rect 442 2514 448 2515
rect 463 2515 464 2516
rect 468 2515 469 2519
rect 511 2519 517 2520
rect 511 2515 512 2519
rect 516 2518 517 2519
rect 527 2519 533 2520
rect 527 2518 528 2519
rect 516 2516 528 2518
rect 516 2515 517 2516
rect 463 2514 469 2515
rect 486 2514 492 2515
rect 511 2514 517 2515
rect 527 2515 528 2516
rect 532 2515 533 2519
rect 575 2519 581 2520
rect 575 2515 576 2519
rect 580 2518 581 2519
rect 591 2519 597 2520
rect 591 2518 592 2519
rect 580 2516 592 2518
rect 580 2515 581 2516
rect 527 2514 533 2515
rect 550 2514 556 2515
rect 575 2514 581 2515
rect 591 2515 592 2516
rect 596 2515 597 2519
rect 654 2519 661 2520
rect 654 2515 655 2519
rect 660 2515 661 2519
rect 706 2519 712 2520
rect 706 2515 707 2519
rect 711 2518 712 2519
rect 719 2519 725 2520
rect 719 2518 720 2519
rect 711 2516 720 2518
rect 711 2515 712 2516
rect 591 2514 597 2515
rect 614 2514 620 2515
rect 654 2514 661 2515
rect 678 2514 684 2515
rect 706 2514 712 2515
rect 719 2515 720 2516
rect 724 2515 725 2519
rect 758 2519 764 2520
rect 758 2515 759 2519
rect 763 2518 764 2519
rect 783 2519 789 2520
rect 783 2518 784 2519
rect 763 2516 784 2518
rect 763 2515 764 2516
rect 719 2514 725 2515
rect 742 2514 748 2515
rect 758 2514 764 2515
rect 783 2515 784 2516
rect 788 2515 789 2519
rect 847 2519 853 2520
rect 847 2515 848 2519
rect 852 2518 853 2519
rect 864 2518 866 2524
rect 1022 2523 1023 2524
rect 1027 2523 1028 2527
rect 1431 2527 1432 2531
rect 1436 2530 1437 2531
rect 1446 2531 1452 2532
rect 1446 2530 1447 2531
rect 1436 2528 1447 2530
rect 1436 2527 1437 2528
rect 1431 2526 1437 2527
rect 1446 2527 1447 2528
rect 1451 2527 1452 2531
rect 1446 2526 1452 2527
rect 1534 2531 1541 2532
rect 1534 2527 1535 2531
rect 1540 2527 1541 2531
rect 1534 2526 1541 2527
rect 1646 2531 1653 2532
rect 1646 2527 1647 2531
rect 1652 2527 1653 2531
rect 1646 2526 1653 2527
rect 1758 2531 1765 2532
rect 1758 2527 1759 2531
rect 1764 2527 1765 2531
rect 1758 2526 1765 2527
rect 1870 2531 1877 2532
rect 1870 2527 1871 2531
rect 1876 2527 1877 2531
rect 1870 2526 1877 2527
rect 1983 2531 1989 2532
rect 1983 2527 1984 2531
rect 1988 2530 1989 2531
rect 2070 2531 2076 2532
rect 2070 2530 2071 2531
rect 1988 2528 2071 2530
rect 1988 2527 1989 2528
rect 1983 2526 1989 2527
rect 2070 2527 2071 2528
rect 2075 2527 2076 2531
rect 2070 2526 2076 2527
rect 2103 2531 2109 2532
rect 2103 2527 2104 2531
rect 2108 2530 2109 2531
rect 2151 2531 2157 2532
rect 2151 2530 2152 2531
rect 2108 2528 2152 2530
rect 2108 2527 2109 2528
rect 2103 2526 2109 2527
rect 2151 2527 2152 2528
rect 2156 2527 2157 2531
rect 2151 2526 2157 2527
rect 2223 2531 2229 2532
rect 2223 2527 2224 2531
rect 2228 2530 2229 2531
rect 2271 2531 2277 2532
rect 2271 2530 2272 2531
rect 2228 2528 2272 2530
rect 2228 2527 2229 2528
rect 2223 2526 2229 2527
rect 2271 2527 2272 2528
rect 2276 2527 2277 2531
rect 2271 2526 2277 2527
rect 2314 2531 2320 2532
rect 2314 2527 2315 2531
rect 2319 2530 2320 2531
rect 2343 2531 2349 2532
rect 2343 2530 2344 2531
rect 2319 2528 2344 2530
rect 2319 2527 2320 2528
rect 2314 2526 2320 2527
rect 2343 2527 2344 2528
rect 2348 2527 2349 2531
rect 2343 2526 2349 2527
rect 1022 2522 1028 2523
rect 852 2516 866 2518
rect 903 2519 909 2520
rect 852 2515 853 2516
rect 903 2515 904 2519
rect 908 2518 909 2519
rect 919 2519 925 2520
rect 919 2518 920 2519
rect 908 2516 920 2518
rect 908 2515 909 2516
rect 783 2514 789 2515
rect 806 2514 812 2515
rect 847 2514 853 2515
rect 870 2514 876 2515
rect 903 2514 909 2515
rect 919 2515 920 2516
rect 924 2515 925 2519
rect 978 2519 984 2520
rect 978 2515 979 2519
rect 983 2518 984 2519
rect 991 2519 997 2520
rect 991 2518 992 2519
rect 983 2516 992 2518
rect 983 2515 984 2516
rect 919 2514 925 2515
rect 942 2514 948 2515
rect 978 2514 984 2515
rect 991 2515 992 2516
rect 996 2515 997 2519
rect 991 2514 997 2515
rect 1014 2514 1020 2515
rect 366 2510 367 2514
rect 371 2510 372 2514
rect 366 2509 372 2510
rect 422 2510 423 2514
rect 427 2510 428 2514
rect 422 2509 428 2510
rect 486 2510 487 2514
rect 491 2510 492 2514
rect 486 2509 492 2510
rect 550 2510 551 2514
rect 555 2510 556 2514
rect 550 2509 556 2510
rect 614 2510 615 2514
rect 619 2510 620 2514
rect 614 2509 620 2510
rect 678 2510 679 2514
rect 683 2510 684 2514
rect 678 2509 684 2510
rect 742 2510 743 2514
rect 747 2510 748 2514
rect 742 2509 748 2510
rect 806 2510 807 2514
rect 811 2510 812 2514
rect 806 2509 812 2510
rect 870 2510 871 2514
rect 875 2510 876 2514
rect 870 2509 876 2510
rect 942 2510 943 2514
rect 947 2510 948 2514
rect 942 2509 948 2510
rect 1014 2510 1015 2514
rect 1019 2510 1020 2514
rect 1014 2509 1020 2510
rect 1527 2511 1533 2512
rect 1527 2507 1528 2511
rect 1532 2510 1533 2511
rect 1542 2511 1548 2512
rect 1542 2510 1543 2511
rect 1532 2508 1543 2510
rect 1532 2507 1533 2508
rect 1527 2506 1533 2507
rect 1542 2507 1543 2508
rect 1547 2507 1548 2511
rect 1570 2511 1576 2512
rect 1570 2507 1571 2511
rect 1575 2510 1576 2511
rect 1607 2511 1613 2512
rect 1607 2510 1608 2511
rect 1575 2508 1608 2510
rect 1575 2507 1576 2508
rect 1542 2506 1548 2507
rect 1550 2506 1556 2507
rect 1570 2506 1576 2507
rect 1607 2507 1608 2508
rect 1612 2507 1613 2511
rect 1650 2511 1656 2512
rect 1650 2507 1651 2511
rect 1655 2510 1656 2511
rect 1695 2511 1701 2512
rect 1695 2510 1696 2511
rect 1655 2508 1696 2510
rect 1655 2507 1656 2508
rect 1607 2506 1613 2507
rect 1630 2506 1636 2507
rect 1650 2506 1656 2507
rect 1695 2507 1696 2508
rect 1700 2507 1701 2511
rect 1738 2511 1744 2512
rect 1738 2507 1739 2511
rect 1743 2510 1744 2511
rect 1783 2511 1789 2512
rect 1783 2510 1784 2511
rect 1743 2508 1784 2510
rect 1743 2507 1744 2508
rect 1695 2506 1701 2507
rect 1718 2506 1724 2507
rect 1738 2506 1744 2507
rect 1783 2507 1784 2508
rect 1788 2507 1789 2511
rect 1826 2511 1832 2512
rect 1826 2507 1827 2511
rect 1831 2510 1832 2511
rect 1879 2511 1885 2512
rect 1879 2510 1880 2511
rect 1831 2508 1880 2510
rect 1831 2507 1832 2508
rect 1783 2506 1789 2507
rect 1806 2506 1812 2507
rect 1826 2506 1832 2507
rect 1879 2507 1880 2508
rect 1884 2507 1885 2511
rect 1974 2511 1981 2512
rect 1974 2507 1975 2511
rect 1980 2507 1981 2511
rect 2018 2511 2024 2512
rect 2018 2507 2019 2511
rect 2023 2510 2024 2511
rect 2071 2511 2077 2512
rect 2071 2510 2072 2511
rect 2023 2508 2072 2510
rect 2023 2507 2024 2508
rect 1879 2506 1885 2507
rect 1902 2506 1908 2507
rect 1974 2506 1981 2507
rect 1998 2506 2004 2507
rect 2018 2506 2024 2507
rect 2071 2507 2072 2508
rect 2076 2507 2077 2511
rect 2114 2511 2120 2512
rect 2114 2507 2115 2511
rect 2119 2510 2120 2511
rect 2167 2511 2173 2512
rect 2167 2510 2168 2511
rect 2119 2508 2168 2510
rect 2119 2507 2120 2508
rect 2071 2506 2077 2507
rect 2094 2506 2100 2507
rect 2114 2506 2120 2507
rect 2167 2507 2168 2508
rect 2172 2507 2173 2511
rect 2270 2511 2277 2512
rect 2270 2507 2271 2511
rect 2276 2507 2277 2511
rect 2375 2511 2381 2512
rect 2375 2507 2376 2511
rect 2380 2510 2381 2511
rect 2390 2511 2396 2512
rect 2390 2510 2391 2511
rect 2380 2508 2391 2510
rect 2380 2507 2381 2508
rect 2167 2506 2173 2507
rect 2190 2506 2196 2507
rect 2270 2506 2277 2507
rect 2294 2506 2300 2507
rect 2375 2506 2381 2507
rect 2390 2507 2391 2508
rect 2395 2507 2396 2511
rect 2390 2506 2396 2507
rect 2398 2506 2404 2507
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 1326 2505 1332 2506
rect 1326 2501 1327 2505
rect 1331 2501 1332 2505
rect 1550 2502 1551 2506
rect 1555 2502 1556 2506
rect 1550 2501 1556 2502
rect 1630 2502 1631 2506
rect 1635 2502 1636 2506
rect 1630 2501 1636 2502
rect 1718 2502 1719 2506
rect 1723 2502 1724 2506
rect 1718 2501 1724 2502
rect 1806 2502 1807 2506
rect 1811 2502 1812 2506
rect 1806 2501 1812 2502
rect 1902 2502 1903 2506
rect 1907 2502 1908 2506
rect 1902 2501 1908 2502
rect 1998 2502 1999 2506
rect 2003 2502 2004 2506
rect 1998 2501 2004 2502
rect 2094 2502 2095 2506
rect 2099 2502 2100 2506
rect 2094 2501 2100 2502
rect 2190 2502 2191 2506
rect 2195 2502 2196 2506
rect 2190 2501 2196 2502
rect 2294 2502 2295 2506
rect 2299 2502 2300 2506
rect 2294 2501 2300 2502
rect 2398 2502 2399 2506
rect 2403 2502 2404 2506
rect 2398 2501 2404 2502
rect 1326 2500 1332 2501
rect 1366 2497 1372 2498
rect 654 2495 660 2496
rect 654 2491 655 2495
rect 659 2494 660 2495
rect 659 2492 882 2494
rect 1366 2493 1367 2497
rect 1371 2493 1372 2497
rect 1366 2492 1372 2493
rect 2582 2497 2588 2498
rect 2582 2493 2583 2497
rect 2587 2493 2588 2497
rect 2582 2492 2588 2493
rect 659 2491 660 2492
rect 654 2490 660 2491
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 350 2487 356 2488
rect 350 2483 351 2487
rect 355 2483 356 2487
rect 406 2487 412 2488
rect 350 2482 356 2483
rect 383 2483 392 2484
rect 383 2479 384 2483
rect 391 2479 392 2483
rect 406 2483 407 2487
rect 411 2483 412 2487
rect 470 2487 476 2488
rect 406 2482 412 2483
rect 439 2483 448 2484
rect 383 2478 392 2479
rect 439 2479 440 2483
rect 447 2479 448 2483
rect 470 2483 471 2487
rect 475 2483 476 2487
rect 534 2487 540 2488
rect 470 2482 476 2483
rect 503 2483 509 2484
rect 439 2478 448 2479
rect 503 2479 504 2483
rect 508 2482 509 2483
rect 511 2483 517 2484
rect 511 2482 512 2483
rect 508 2480 512 2482
rect 508 2479 509 2480
rect 503 2478 509 2479
rect 511 2479 512 2480
rect 516 2479 517 2483
rect 534 2483 535 2487
rect 539 2483 540 2487
rect 575 2487 581 2488
rect 575 2486 576 2487
rect 534 2482 540 2483
rect 567 2485 576 2486
rect 567 2481 568 2485
rect 572 2484 576 2485
rect 572 2481 573 2484
rect 575 2483 576 2484
rect 580 2483 581 2487
rect 575 2482 581 2483
rect 598 2487 604 2488
rect 598 2483 599 2487
rect 603 2483 604 2487
rect 662 2487 668 2488
rect 598 2482 604 2483
rect 622 2483 628 2484
rect 567 2480 573 2481
rect 511 2478 517 2479
rect 622 2479 623 2483
rect 627 2482 628 2483
rect 631 2483 637 2484
rect 631 2482 632 2483
rect 627 2480 632 2482
rect 627 2479 628 2480
rect 622 2478 628 2479
rect 631 2479 632 2480
rect 636 2479 637 2483
rect 662 2483 663 2487
rect 667 2483 668 2487
rect 726 2487 732 2488
rect 662 2482 668 2483
rect 695 2483 701 2484
rect 631 2478 637 2479
rect 695 2479 696 2483
rect 700 2482 701 2483
rect 706 2483 712 2484
rect 706 2482 707 2483
rect 700 2480 707 2482
rect 700 2479 701 2480
rect 695 2478 701 2479
rect 706 2479 707 2480
rect 711 2479 712 2483
rect 726 2483 727 2487
rect 731 2483 732 2487
rect 790 2487 796 2488
rect 726 2482 732 2483
rect 758 2483 765 2484
rect 706 2478 712 2479
rect 758 2479 759 2483
rect 764 2479 765 2483
rect 790 2483 791 2487
rect 795 2483 796 2487
rect 854 2487 860 2488
rect 790 2482 796 2483
rect 823 2483 829 2484
rect 758 2478 765 2479
rect 823 2479 824 2483
rect 828 2482 829 2483
rect 854 2483 855 2487
rect 859 2483 860 2487
rect 854 2482 860 2483
rect 880 2482 882 2492
rect 1326 2488 1332 2489
rect 926 2487 932 2488
rect 887 2483 893 2484
rect 887 2482 888 2483
rect 828 2480 846 2482
rect 880 2480 888 2482
rect 828 2479 829 2480
rect 823 2478 829 2479
rect 844 2474 846 2480
rect 887 2479 888 2480
rect 892 2479 893 2483
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 978 2487 984 2488
rect 978 2486 979 2487
rect 926 2482 932 2483
rect 959 2485 979 2486
rect 959 2481 960 2485
rect 964 2484 979 2485
rect 964 2481 965 2484
rect 978 2483 979 2484
rect 983 2483 984 2487
rect 978 2482 984 2483
rect 998 2487 1004 2488
rect 998 2483 999 2487
rect 1003 2483 1004 2487
rect 1326 2484 1327 2488
rect 1331 2484 1332 2488
rect 998 2482 1004 2483
rect 1022 2483 1028 2484
rect 959 2480 965 2481
rect 887 2478 893 2479
rect 1022 2479 1023 2483
rect 1027 2482 1028 2483
rect 1031 2483 1037 2484
rect 1326 2483 1332 2484
rect 2270 2487 2276 2488
rect 2270 2483 2271 2487
rect 2275 2486 2276 2487
rect 2275 2484 2410 2486
rect 2275 2483 2276 2484
rect 1031 2482 1032 2483
rect 1027 2480 1032 2482
rect 1027 2479 1028 2480
rect 1022 2478 1028 2479
rect 1031 2479 1032 2480
rect 1036 2479 1037 2483
rect 2270 2482 2276 2483
rect 1031 2478 1037 2479
rect 1366 2480 1372 2481
rect 1366 2476 1367 2480
rect 1371 2476 1372 2480
rect 983 2475 989 2476
rect 1366 2475 1372 2476
rect 1534 2479 1540 2480
rect 1534 2475 1535 2479
rect 1539 2475 1540 2479
rect 1614 2479 1620 2480
rect 983 2474 984 2475
rect 844 2472 984 2474
rect 983 2471 984 2472
rect 988 2471 989 2475
rect 1534 2474 1540 2475
rect 1567 2475 1576 2476
rect 983 2470 989 2471
rect 1567 2471 1568 2475
rect 1575 2471 1576 2475
rect 1614 2475 1615 2479
rect 1619 2475 1620 2479
rect 1702 2479 1708 2480
rect 1614 2474 1620 2475
rect 1647 2475 1656 2476
rect 1567 2470 1576 2471
rect 1647 2471 1648 2475
rect 1655 2471 1656 2475
rect 1702 2475 1703 2479
rect 1707 2475 1708 2479
rect 1790 2479 1796 2480
rect 1702 2474 1708 2475
rect 1735 2475 1744 2476
rect 1647 2470 1656 2471
rect 1735 2471 1736 2475
rect 1743 2471 1744 2475
rect 1790 2475 1791 2479
rect 1795 2475 1796 2479
rect 1886 2479 1892 2480
rect 1790 2474 1796 2475
rect 1823 2475 1832 2476
rect 1735 2470 1744 2471
rect 1823 2471 1824 2475
rect 1831 2471 1832 2475
rect 1886 2475 1887 2479
rect 1891 2475 1892 2479
rect 1982 2479 1988 2480
rect 1886 2474 1892 2475
rect 1919 2475 1925 2476
rect 1919 2474 1920 2475
rect 1823 2470 1832 2471
rect 1896 2472 1920 2474
rect 1654 2467 1660 2468
rect 1654 2463 1655 2467
rect 1659 2466 1660 2467
rect 1896 2466 1898 2472
rect 1919 2471 1920 2472
rect 1924 2471 1925 2475
rect 1982 2475 1983 2479
rect 1987 2475 1988 2479
rect 2078 2479 2084 2480
rect 1982 2474 1988 2475
rect 2015 2475 2024 2476
rect 1919 2470 1925 2471
rect 2015 2471 2016 2475
rect 2023 2471 2024 2475
rect 2078 2475 2079 2479
rect 2083 2475 2084 2479
rect 2174 2479 2180 2480
rect 2078 2474 2084 2475
rect 2111 2475 2120 2476
rect 2015 2470 2024 2471
rect 2111 2471 2112 2475
rect 2119 2471 2120 2475
rect 2174 2475 2175 2479
rect 2179 2475 2180 2479
rect 2278 2479 2284 2480
rect 2174 2474 2180 2475
rect 2207 2475 2213 2476
rect 2111 2470 2120 2471
rect 2207 2471 2208 2475
rect 2212 2474 2213 2475
rect 2254 2475 2260 2476
rect 2254 2474 2255 2475
rect 2212 2472 2255 2474
rect 2212 2471 2213 2472
rect 2207 2470 2213 2471
rect 2254 2471 2255 2472
rect 2259 2471 2260 2475
rect 2278 2475 2279 2479
rect 2283 2475 2284 2479
rect 2382 2479 2388 2480
rect 2278 2474 2284 2475
rect 2311 2475 2320 2476
rect 2254 2470 2260 2471
rect 2311 2471 2312 2475
rect 2319 2471 2320 2475
rect 2382 2475 2383 2479
rect 2387 2475 2388 2479
rect 2382 2474 2388 2475
rect 2408 2474 2410 2484
rect 2582 2480 2588 2481
rect 2582 2476 2583 2480
rect 2587 2476 2588 2480
rect 2415 2475 2421 2476
rect 2582 2475 2588 2476
rect 2415 2474 2416 2475
rect 2408 2472 2416 2474
rect 2311 2470 2320 2471
rect 2415 2471 2416 2472
rect 2420 2471 2421 2475
rect 2415 2470 2421 2471
rect 1659 2464 1898 2466
rect 1659 2463 1660 2464
rect 1654 2462 1660 2463
rect 278 2459 284 2460
rect 278 2455 279 2459
rect 283 2458 284 2459
rect 718 2459 724 2460
rect 283 2456 498 2458
rect 283 2455 284 2456
rect 278 2454 284 2455
rect 303 2451 309 2452
rect 270 2449 276 2450
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 270 2445 271 2449
rect 275 2445 276 2449
rect 303 2447 304 2451
rect 308 2450 309 2451
rect 326 2451 332 2452
rect 326 2450 327 2451
rect 308 2448 327 2450
rect 308 2447 309 2448
rect 303 2446 309 2447
rect 326 2447 327 2448
rect 331 2447 332 2451
rect 367 2451 373 2452
rect 326 2446 332 2447
rect 334 2449 340 2450
rect 270 2444 276 2445
rect 334 2445 335 2449
rect 339 2445 340 2449
rect 367 2447 368 2451
rect 372 2450 373 2451
rect 390 2451 396 2452
rect 390 2450 391 2451
rect 372 2448 391 2450
rect 372 2447 373 2448
rect 367 2446 373 2447
rect 390 2447 391 2448
rect 395 2447 396 2451
rect 422 2451 428 2452
rect 390 2446 396 2447
rect 398 2449 404 2450
rect 334 2444 340 2445
rect 398 2445 399 2449
rect 403 2445 404 2449
rect 422 2447 423 2451
rect 427 2450 428 2451
rect 431 2451 437 2452
rect 431 2450 432 2451
rect 427 2448 432 2450
rect 427 2447 428 2448
rect 422 2446 428 2447
rect 431 2447 432 2448
rect 436 2447 437 2451
rect 496 2450 498 2456
rect 511 2455 517 2456
rect 503 2451 509 2452
rect 503 2450 504 2451
rect 431 2446 437 2447
rect 470 2449 476 2450
rect 398 2444 404 2445
rect 470 2445 471 2449
rect 475 2445 476 2449
rect 496 2448 504 2450
rect 503 2447 504 2448
rect 508 2447 509 2451
rect 511 2451 512 2455
rect 516 2454 517 2455
rect 591 2455 597 2456
rect 516 2452 578 2454
rect 516 2451 517 2452
rect 511 2450 517 2451
rect 576 2450 578 2452
rect 583 2451 589 2452
rect 583 2450 584 2451
rect 503 2446 509 2447
rect 550 2449 556 2450
rect 470 2444 476 2445
rect 550 2445 551 2449
rect 555 2445 556 2449
rect 576 2448 584 2450
rect 583 2447 584 2448
rect 588 2447 589 2451
rect 591 2451 592 2455
rect 596 2454 597 2455
rect 718 2455 719 2459
rect 723 2458 724 2459
rect 723 2456 1050 2458
rect 723 2455 724 2456
rect 718 2454 724 2455
rect 596 2452 658 2454
rect 596 2451 597 2452
rect 591 2450 597 2451
rect 656 2450 658 2452
rect 663 2451 669 2452
rect 663 2450 664 2451
rect 583 2446 589 2447
rect 630 2449 636 2450
rect 550 2444 556 2445
rect 630 2445 631 2449
rect 635 2445 636 2449
rect 656 2448 664 2450
rect 663 2447 664 2448
rect 668 2447 669 2451
rect 743 2451 749 2452
rect 663 2446 669 2447
rect 710 2449 716 2450
rect 630 2444 636 2445
rect 710 2445 711 2449
rect 715 2445 716 2449
rect 743 2447 744 2451
rect 748 2450 749 2451
rect 774 2451 780 2452
rect 774 2450 775 2451
rect 748 2448 775 2450
rect 748 2447 749 2448
rect 743 2446 749 2447
rect 774 2447 775 2448
rect 779 2447 780 2451
rect 815 2451 821 2452
rect 774 2446 780 2447
rect 782 2449 788 2450
rect 710 2444 716 2445
rect 782 2445 783 2449
rect 787 2445 788 2449
rect 815 2447 816 2451
rect 820 2450 821 2451
rect 854 2451 860 2452
rect 854 2450 855 2451
rect 820 2448 855 2450
rect 820 2447 821 2448
rect 815 2446 821 2447
rect 854 2447 855 2448
rect 859 2447 860 2451
rect 895 2451 901 2452
rect 854 2446 860 2447
rect 862 2449 868 2450
rect 782 2444 788 2445
rect 862 2445 863 2449
rect 867 2445 868 2449
rect 895 2447 896 2451
rect 900 2450 901 2451
rect 903 2451 909 2452
rect 903 2450 904 2451
rect 900 2448 904 2450
rect 900 2447 901 2448
rect 895 2446 901 2447
rect 903 2447 904 2448
rect 908 2447 909 2451
rect 975 2451 981 2452
rect 903 2446 909 2447
rect 942 2449 948 2450
rect 862 2444 868 2445
rect 942 2445 943 2449
rect 947 2445 948 2449
rect 975 2447 976 2451
rect 980 2450 981 2451
rect 1014 2451 1020 2452
rect 1014 2450 1015 2451
rect 980 2448 1015 2450
rect 980 2447 981 2448
rect 975 2446 981 2447
rect 1014 2447 1015 2448
rect 1019 2447 1020 2451
rect 1048 2450 1050 2456
rect 1974 2455 1980 2456
rect 1055 2451 1061 2452
rect 1055 2450 1056 2451
rect 1014 2446 1020 2447
rect 1022 2449 1028 2450
rect 942 2444 948 2445
rect 1022 2445 1023 2449
rect 1027 2445 1028 2449
rect 1048 2448 1056 2450
rect 1055 2447 1056 2448
rect 1060 2447 1061 2451
rect 1974 2451 1975 2455
rect 1979 2454 1980 2455
rect 1979 2452 2194 2454
rect 1979 2451 1980 2452
rect 1974 2450 1980 2451
rect 1055 2446 1061 2447
rect 1326 2448 1332 2449
rect 1022 2444 1028 2445
rect 1326 2444 1327 2448
rect 1331 2444 1332 2448
rect 1679 2447 1685 2448
rect 1646 2445 1652 2446
rect 110 2443 116 2444
rect 1326 2443 1332 2444
rect 1366 2444 1372 2445
rect 1366 2440 1367 2444
rect 1371 2440 1372 2444
rect 1646 2441 1647 2445
rect 1651 2441 1652 2445
rect 1679 2443 1680 2447
rect 1684 2446 1685 2447
rect 1694 2447 1700 2448
rect 1694 2446 1695 2447
rect 1684 2444 1695 2446
rect 1684 2443 1685 2444
rect 1679 2442 1685 2443
rect 1694 2443 1695 2444
rect 1699 2443 1700 2447
rect 1735 2447 1741 2448
rect 1694 2442 1700 2443
rect 1702 2445 1708 2446
rect 1646 2440 1652 2441
rect 1702 2441 1703 2445
rect 1707 2441 1708 2445
rect 1735 2443 1736 2447
rect 1740 2446 1741 2447
rect 1758 2447 1764 2448
rect 1758 2446 1759 2447
rect 1740 2444 1759 2446
rect 1740 2443 1741 2444
rect 1735 2442 1741 2443
rect 1758 2443 1759 2444
rect 1763 2443 1764 2447
rect 1799 2447 1805 2448
rect 1758 2442 1764 2443
rect 1766 2445 1772 2446
rect 1702 2440 1708 2441
rect 1766 2441 1767 2445
rect 1771 2441 1772 2445
rect 1799 2443 1800 2447
rect 1804 2446 1805 2447
rect 1830 2447 1836 2448
rect 1830 2446 1831 2447
rect 1804 2444 1831 2446
rect 1804 2443 1805 2444
rect 1799 2442 1805 2443
rect 1830 2443 1831 2444
rect 1835 2443 1836 2447
rect 1871 2447 1877 2448
rect 1830 2442 1836 2443
rect 1838 2445 1844 2446
rect 1766 2440 1772 2441
rect 1838 2441 1839 2445
rect 1843 2441 1844 2445
rect 1871 2443 1872 2447
rect 1876 2446 1877 2447
rect 1902 2447 1908 2448
rect 1902 2446 1903 2447
rect 1876 2444 1903 2446
rect 1876 2443 1877 2444
rect 1871 2442 1877 2443
rect 1902 2443 1903 2444
rect 1907 2443 1908 2447
rect 1934 2447 1940 2448
rect 1902 2442 1908 2443
rect 1910 2445 1916 2446
rect 1838 2440 1844 2441
rect 1910 2441 1911 2445
rect 1915 2441 1916 2445
rect 1934 2443 1935 2447
rect 1939 2446 1940 2447
rect 1943 2447 1949 2448
rect 1943 2446 1944 2447
rect 1939 2444 1944 2446
rect 1939 2443 1940 2444
rect 1934 2442 1940 2443
rect 1943 2443 1944 2444
rect 1948 2443 1949 2447
rect 2023 2447 2029 2448
rect 1943 2442 1949 2443
rect 1990 2445 1996 2446
rect 1910 2440 1916 2441
rect 1990 2441 1991 2445
rect 1995 2441 1996 2445
rect 2023 2443 2024 2447
rect 2028 2446 2029 2447
rect 2070 2447 2076 2448
rect 2070 2446 2071 2447
rect 2028 2444 2071 2446
rect 2028 2443 2029 2444
rect 2023 2442 2029 2443
rect 2070 2443 2071 2444
rect 2075 2443 2076 2447
rect 2111 2447 2117 2448
rect 2070 2442 2076 2443
rect 2078 2445 2084 2446
rect 1990 2440 1996 2441
rect 2078 2441 2079 2445
rect 2083 2441 2084 2445
rect 2111 2443 2112 2447
rect 2116 2446 2117 2447
rect 2158 2447 2164 2448
rect 2158 2446 2159 2447
rect 2116 2444 2159 2446
rect 2116 2443 2117 2444
rect 2111 2442 2117 2443
rect 2158 2443 2159 2444
rect 2163 2443 2164 2447
rect 2192 2446 2194 2452
rect 2210 2451 2216 2452
rect 2199 2447 2205 2448
rect 2199 2446 2200 2447
rect 2158 2442 2164 2443
rect 2166 2445 2172 2446
rect 2078 2440 2084 2441
rect 2166 2441 2167 2445
rect 2171 2441 2172 2445
rect 2192 2444 2200 2446
rect 2199 2443 2200 2444
rect 2204 2443 2205 2447
rect 2210 2447 2211 2451
rect 2215 2450 2216 2451
rect 2462 2451 2468 2452
rect 2215 2448 2290 2450
rect 2215 2447 2216 2448
rect 2210 2446 2216 2447
rect 2288 2446 2290 2448
rect 2295 2447 2301 2448
rect 2295 2446 2296 2447
rect 2199 2442 2205 2443
rect 2262 2445 2268 2446
rect 2166 2440 2172 2441
rect 2262 2441 2263 2445
rect 2267 2441 2268 2445
rect 2288 2444 2296 2446
rect 2295 2443 2296 2444
rect 2300 2443 2301 2447
rect 2390 2447 2397 2448
rect 2295 2442 2301 2443
rect 2358 2445 2364 2446
rect 2262 2440 2268 2441
rect 2358 2441 2359 2445
rect 2363 2441 2364 2445
rect 2390 2443 2391 2447
rect 2396 2443 2397 2447
rect 2462 2447 2463 2451
rect 2467 2450 2468 2451
rect 2467 2448 2554 2450
rect 2467 2447 2468 2448
rect 2462 2446 2468 2447
rect 2552 2446 2554 2448
rect 2559 2447 2565 2448
rect 2559 2446 2560 2447
rect 2390 2442 2397 2443
rect 2454 2445 2460 2446
rect 2358 2440 2364 2441
rect 2454 2441 2455 2445
rect 2459 2441 2460 2445
rect 2454 2440 2460 2441
rect 2526 2445 2532 2446
rect 2526 2441 2527 2445
rect 2531 2441 2532 2445
rect 2552 2444 2560 2446
rect 2559 2443 2560 2444
rect 2564 2443 2565 2447
rect 2559 2442 2565 2443
rect 2582 2444 2588 2445
rect 2526 2440 2532 2441
rect 2582 2440 2583 2444
rect 2587 2440 2588 2444
rect 1366 2439 1372 2440
rect 2582 2439 2588 2440
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 1326 2431 1332 2432
rect 1326 2427 1327 2431
rect 1331 2427 1332 2431
rect 1326 2426 1332 2427
rect 1366 2427 1372 2428
rect 1366 2423 1367 2427
rect 1371 2423 1372 2427
rect 286 2422 292 2423
rect 286 2418 287 2422
rect 291 2418 292 2422
rect 286 2417 292 2418
rect 350 2422 356 2423
rect 350 2418 351 2422
rect 355 2418 356 2422
rect 350 2417 356 2418
rect 414 2422 420 2423
rect 414 2418 415 2422
rect 419 2418 420 2422
rect 414 2417 420 2418
rect 486 2422 492 2423
rect 486 2418 487 2422
rect 491 2418 492 2422
rect 486 2417 492 2418
rect 566 2422 572 2423
rect 566 2418 567 2422
rect 571 2418 572 2422
rect 566 2417 572 2418
rect 646 2422 652 2423
rect 646 2418 647 2422
rect 651 2418 652 2422
rect 646 2417 652 2418
rect 726 2422 732 2423
rect 726 2418 727 2422
rect 731 2418 732 2422
rect 726 2417 732 2418
rect 798 2422 804 2423
rect 798 2418 799 2422
rect 803 2418 804 2422
rect 798 2417 804 2418
rect 878 2422 884 2423
rect 878 2418 879 2422
rect 883 2418 884 2422
rect 878 2417 884 2418
rect 958 2422 964 2423
rect 958 2418 959 2422
rect 963 2418 964 2422
rect 958 2417 964 2418
rect 1038 2422 1044 2423
rect 1366 2422 1372 2423
rect 2582 2427 2588 2428
rect 2582 2423 2583 2427
rect 2587 2423 2588 2427
rect 2582 2422 2588 2423
rect 1038 2418 1039 2422
rect 1043 2418 1044 2422
rect 1038 2417 1044 2418
rect 1662 2418 1668 2419
rect 263 2415 269 2416
rect 263 2411 264 2415
rect 268 2414 269 2415
rect 278 2415 284 2416
rect 278 2414 279 2415
rect 268 2412 279 2414
rect 268 2411 269 2412
rect 263 2410 269 2411
rect 278 2411 279 2412
rect 283 2411 284 2415
rect 278 2410 284 2411
rect 326 2415 333 2416
rect 326 2411 327 2415
rect 332 2411 333 2415
rect 326 2410 333 2411
rect 390 2415 397 2416
rect 390 2411 391 2415
rect 396 2411 397 2415
rect 390 2410 397 2411
rect 463 2415 469 2416
rect 463 2411 464 2415
rect 468 2414 469 2415
rect 511 2415 517 2416
rect 511 2414 512 2415
rect 468 2412 512 2414
rect 468 2411 469 2412
rect 463 2410 469 2411
rect 511 2411 512 2412
rect 516 2411 517 2415
rect 511 2410 517 2411
rect 543 2415 549 2416
rect 543 2411 544 2415
rect 548 2414 549 2415
rect 591 2415 597 2416
rect 591 2414 592 2415
rect 548 2412 592 2414
rect 548 2411 549 2412
rect 543 2410 549 2411
rect 591 2411 592 2412
rect 596 2411 597 2415
rect 591 2410 597 2411
rect 622 2415 629 2416
rect 622 2411 623 2415
rect 628 2411 629 2415
rect 622 2410 629 2411
rect 703 2415 709 2416
rect 703 2411 704 2415
rect 708 2414 709 2415
rect 718 2415 724 2416
rect 718 2414 719 2415
rect 708 2412 719 2414
rect 708 2411 709 2412
rect 703 2410 709 2411
rect 718 2411 719 2412
rect 723 2411 724 2415
rect 718 2410 724 2411
rect 774 2415 781 2416
rect 774 2411 775 2415
rect 780 2411 781 2415
rect 774 2410 781 2411
rect 854 2415 861 2416
rect 854 2411 855 2415
rect 860 2411 861 2415
rect 854 2410 861 2411
rect 934 2415 941 2416
rect 934 2411 935 2415
rect 940 2411 941 2415
rect 934 2410 941 2411
rect 1014 2415 1021 2416
rect 1014 2411 1015 2415
rect 1020 2411 1021 2415
rect 1662 2414 1663 2418
rect 1667 2414 1668 2418
rect 1662 2413 1668 2414
rect 1718 2418 1724 2419
rect 1718 2414 1719 2418
rect 1723 2414 1724 2418
rect 1718 2413 1724 2414
rect 1782 2418 1788 2419
rect 1782 2414 1783 2418
rect 1787 2414 1788 2418
rect 1782 2413 1788 2414
rect 1854 2418 1860 2419
rect 1854 2414 1855 2418
rect 1859 2414 1860 2418
rect 1854 2413 1860 2414
rect 1926 2418 1932 2419
rect 1926 2414 1927 2418
rect 1931 2414 1932 2418
rect 1926 2413 1932 2414
rect 2006 2418 2012 2419
rect 2006 2414 2007 2418
rect 2011 2414 2012 2418
rect 2006 2413 2012 2414
rect 2094 2418 2100 2419
rect 2094 2414 2095 2418
rect 2099 2414 2100 2418
rect 2094 2413 2100 2414
rect 2182 2418 2188 2419
rect 2182 2414 2183 2418
rect 2187 2414 2188 2418
rect 2182 2413 2188 2414
rect 2278 2418 2284 2419
rect 2278 2414 2279 2418
rect 2283 2414 2284 2418
rect 2278 2413 2284 2414
rect 2374 2418 2380 2419
rect 2374 2414 2375 2418
rect 2379 2414 2380 2418
rect 2374 2413 2380 2414
rect 2470 2418 2476 2419
rect 2470 2414 2471 2418
rect 2475 2414 2476 2418
rect 2470 2413 2476 2414
rect 2542 2418 2548 2419
rect 2542 2414 2543 2418
rect 2547 2414 2548 2418
rect 2542 2413 2548 2414
rect 1014 2410 1021 2411
rect 1639 2411 1645 2412
rect 1639 2407 1640 2411
rect 1644 2410 1645 2411
rect 1654 2411 1660 2412
rect 1654 2410 1655 2411
rect 1644 2408 1655 2410
rect 1644 2407 1645 2408
rect 1639 2406 1645 2407
rect 1654 2407 1655 2408
rect 1659 2407 1660 2411
rect 1654 2406 1660 2407
rect 1694 2411 1701 2412
rect 1694 2407 1695 2411
rect 1700 2407 1701 2411
rect 1694 2406 1701 2407
rect 1758 2411 1765 2412
rect 1758 2407 1759 2411
rect 1764 2407 1765 2411
rect 1758 2406 1765 2407
rect 1830 2411 1837 2412
rect 1830 2407 1831 2411
rect 1836 2407 1837 2411
rect 1830 2406 1837 2407
rect 1902 2411 1909 2412
rect 1902 2407 1903 2411
rect 1908 2407 1909 2411
rect 1962 2411 1968 2412
rect 1902 2406 1909 2407
rect 1934 2407 1940 2408
rect 1934 2403 1935 2407
rect 1939 2403 1940 2407
rect 1962 2407 1963 2411
rect 1967 2410 1968 2411
rect 1983 2411 1989 2412
rect 1983 2410 1984 2411
rect 1967 2408 1984 2410
rect 1967 2407 1968 2408
rect 1962 2406 1968 2407
rect 1983 2407 1984 2408
rect 1988 2407 1989 2411
rect 1983 2406 1989 2407
rect 2070 2411 2077 2412
rect 2070 2407 2071 2411
rect 2076 2407 2077 2411
rect 2070 2406 2077 2407
rect 2158 2411 2165 2412
rect 2158 2407 2159 2411
rect 2164 2407 2165 2411
rect 2158 2406 2165 2407
rect 2254 2411 2261 2412
rect 2254 2407 2255 2411
rect 2260 2407 2261 2411
rect 2254 2406 2261 2407
rect 2351 2411 2357 2412
rect 2351 2407 2352 2411
rect 2356 2410 2357 2411
rect 2438 2411 2444 2412
rect 2438 2410 2439 2411
rect 2356 2408 2439 2410
rect 2356 2407 2357 2408
rect 2351 2406 2357 2407
rect 2438 2407 2439 2408
rect 2443 2407 2444 2411
rect 2438 2406 2444 2407
rect 2447 2411 2453 2412
rect 2447 2407 2448 2411
rect 2452 2410 2453 2411
rect 2462 2411 2468 2412
rect 2462 2410 2463 2411
rect 2452 2408 2463 2410
rect 2452 2407 2453 2408
rect 2447 2406 2453 2407
rect 2462 2407 2463 2408
rect 2467 2407 2468 2411
rect 2462 2406 2468 2407
rect 2519 2411 2525 2412
rect 2519 2407 2520 2411
rect 2524 2410 2525 2411
rect 2558 2411 2564 2412
rect 2558 2410 2559 2411
rect 2524 2408 2559 2410
rect 2524 2407 2525 2408
rect 2519 2406 2525 2407
rect 2558 2407 2559 2408
rect 2563 2407 2564 2411
rect 2558 2406 2564 2407
rect 1934 2402 1940 2403
rect 2054 2403 2060 2404
rect 2054 2402 2055 2403
rect 1552 2400 1938 2402
rect 1999 2400 2055 2402
rect 223 2399 229 2400
rect 223 2395 224 2399
rect 228 2398 229 2399
rect 238 2399 244 2400
rect 238 2398 239 2399
rect 228 2396 239 2398
rect 228 2395 229 2396
rect 223 2394 229 2395
rect 238 2395 239 2396
rect 243 2395 244 2399
rect 266 2399 272 2400
rect 266 2395 267 2399
rect 271 2398 272 2399
rect 311 2399 317 2400
rect 311 2398 312 2399
rect 271 2396 312 2398
rect 271 2395 272 2396
rect 238 2394 244 2395
rect 246 2394 252 2395
rect 266 2394 272 2395
rect 311 2395 312 2396
rect 316 2395 317 2399
rect 407 2399 413 2400
rect 407 2395 408 2399
rect 412 2398 413 2399
rect 422 2399 428 2400
rect 422 2398 423 2399
rect 412 2396 423 2398
rect 412 2395 413 2396
rect 311 2394 317 2395
rect 334 2394 340 2395
rect 407 2394 413 2395
rect 422 2395 423 2396
rect 427 2395 428 2399
rect 450 2399 456 2400
rect 450 2395 451 2399
rect 455 2398 456 2399
rect 503 2399 509 2400
rect 503 2398 504 2399
rect 455 2396 504 2398
rect 455 2395 456 2396
rect 422 2394 428 2395
rect 430 2394 436 2395
rect 450 2394 456 2395
rect 503 2395 504 2396
rect 508 2395 509 2399
rect 546 2399 552 2400
rect 546 2395 547 2399
rect 551 2398 552 2399
rect 607 2399 613 2400
rect 607 2398 608 2399
rect 551 2396 608 2398
rect 551 2395 552 2396
rect 503 2394 509 2395
rect 526 2394 532 2395
rect 546 2394 552 2395
rect 607 2395 608 2396
rect 612 2395 613 2399
rect 702 2399 709 2400
rect 702 2395 703 2399
rect 708 2395 709 2399
rect 746 2399 752 2400
rect 746 2395 747 2399
rect 751 2398 752 2399
rect 799 2399 805 2400
rect 799 2398 800 2399
rect 751 2396 800 2398
rect 751 2395 752 2396
rect 607 2394 613 2395
rect 630 2394 636 2395
rect 702 2394 709 2395
rect 726 2394 732 2395
rect 746 2394 752 2395
rect 799 2395 800 2396
rect 804 2395 805 2399
rect 842 2399 848 2400
rect 842 2395 843 2399
rect 847 2398 848 2399
rect 895 2399 901 2400
rect 895 2398 896 2399
rect 847 2396 896 2398
rect 847 2395 848 2396
rect 799 2394 805 2395
rect 822 2394 828 2395
rect 842 2394 848 2395
rect 895 2395 896 2396
rect 900 2395 901 2399
rect 967 2399 973 2400
rect 967 2395 968 2399
rect 972 2398 973 2399
rect 991 2399 997 2400
rect 991 2398 992 2399
rect 972 2396 992 2398
rect 972 2395 973 2396
rect 895 2394 901 2395
rect 918 2394 924 2395
rect 967 2394 973 2395
rect 991 2395 992 2396
rect 996 2395 997 2399
rect 1039 2399 1045 2400
rect 1039 2395 1040 2399
rect 1044 2398 1045 2399
rect 1087 2399 1093 2400
rect 1087 2398 1088 2399
rect 1044 2396 1088 2398
rect 1044 2395 1045 2396
rect 991 2394 997 2395
rect 1014 2394 1020 2395
rect 1039 2394 1045 2395
rect 1087 2395 1088 2396
rect 1092 2395 1093 2399
rect 1431 2395 1437 2396
rect 1087 2394 1093 2395
rect 1110 2394 1116 2395
rect 246 2390 247 2394
rect 251 2390 252 2394
rect 246 2389 252 2390
rect 334 2390 335 2394
rect 339 2390 340 2394
rect 334 2389 340 2390
rect 430 2390 431 2394
rect 435 2390 436 2394
rect 430 2389 436 2390
rect 526 2390 527 2394
rect 531 2390 532 2394
rect 526 2389 532 2390
rect 630 2390 631 2394
rect 635 2390 636 2394
rect 630 2389 636 2390
rect 726 2390 727 2394
rect 731 2390 732 2394
rect 726 2389 732 2390
rect 822 2390 823 2394
rect 827 2390 828 2394
rect 822 2389 828 2390
rect 918 2390 919 2394
rect 923 2390 924 2394
rect 918 2389 924 2390
rect 1014 2390 1015 2394
rect 1019 2390 1020 2394
rect 1014 2389 1020 2390
rect 1110 2390 1111 2394
rect 1115 2390 1116 2394
rect 1431 2391 1432 2395
rect 1436 2394 1437 2395
rect 1446 2395 1452 2396
rect 1446 2394 1447 2395
rect 1436 2392 1447 2394
rect 1436 2391 1437 2392
rect 1431 2390 1437 2391
rect 1446 2391 1447 2392
rect 1451 2391 1452 2395
rect 1535 2395 1541 2396
rect 1535 2391 1536 2395
rect 1540 2394 1541 2395
rect 1552 2394 1554 2400
rect 1999 2398 2001 2400
rect 2054 2399 2055 2400
rect 2059 2399 2060 2403
rect 2054 2398 2060 2399
rect 1936 2396 2001 2398
rect 1540 2392 1554 2394
rect 1578 2395 1584 2396
rect 1540 2391 1541 2392
rect 1578 2391 1579 2395
rect 1583 2394 1584 2395
rect 1639 2395 1645 2396
rect 1639 2394 1640 2395
rect 1583 2392 1640 2394
rect 1583 2391 1584 2392
rect 1446 2390 1452 2391
rect 1454 2390 1460 2391
rect 1535 2390 1541 2391
rect 1558 2390 1564 2391
rect 1578 2390 1584 2391
rect 1639 2391 1640 2392
rect 1644 2391 1645 2395
rect 1682 2395 1688 2396
rect 1682 2391 1683 2395
rect 1687 2394 1688 2395
rect 1735 2395 1741 2396
rect 1735 2394 1736 2395
rect 1687 2392 1736 2394
rect 1687 2391 1688 2392
rect 1639 2390 1645 2391
rect 1662 2390 1668 2391
rect 1682 2390 1688 2391
rect 1735 2391 1736 2392
rect 1740 2391 1741 2395
rect 1783 2395 1789 2396
rect 1783 2391 1784 2395
rect 1788 2394 1789 2395
rect 1831 2395 1837 2396
rect 1831 2394 1832 2395
rect 1788 2392 1832 2394
rect 1788 2391 1789 2392
rect 1735 2390 1741 2391
rect 1758 2390 1764 2391
rect 1783 2390 1789 2391
rect 1831 2391 1832 2392
rect 1836 2391 1837 2395
rect 1919 2395 1925 2396
rect 1919 2391 1920 2395
rect 1924 2394 1925 2395
rect 1936 2394 1938 2396
rect 1924 2392 1938 2394
rect 2014 2395 2021 2396
rect 1924 2391 1925 2392
rect 2014 2391 2015 2395
rect 2020 2391 2021 2395
rect 2111 2395 2117 2396
rect 2111 2391 2112 2395
rect 2116 2394 2117 2395
rect 2126 2395 2132 2396
rect 2126 2394 2127 2395
rect 2116 2392 2127 2394
rect 2116 2391 2117 2392
rect 1831 2390 1837 2391
rect 1854 2390 1860 2391
rect 1919 2390 1925 2391
rect 1942 2390 1948 2391
rect 2014 2390 2021 2391
rect 2038 2390 2044 2391
rect 2111 2390 2117 2391
rect 2126 2391 2127 2392
rect 2131 2391 2132 2395
rect 2207 2395 2216 2396
rect 2207 2391 2208 2395
rect 2215 2391 2216 2395
rect 2246 2395 2252 2396
rect 2246 2391 2247 2395
rect 2251 2394 2252 2395
rect 2311 2395 2317 2396
rect 2311 2394 2312 2395
rect 2251 2392 2312 2394
rect 2251 2391 2252 2392
rect 2126 2390 2132 2391
rect 2134 2390 2140 2391
rect 2207 2390 2216 2391
rect 2230 2390 2236 2391
rect 2246 2390 2252 2391
rect 2311 2391 2312 2392
rect 2316 2391 2317 2395
rect 2422 2395 2429 2396
rect 2422 2391 2423 2395
rect 2428 2391 2429 2395
rect 2519 2395 2525 2396
rect 2519 2391 2520 2395
rect 2524 2394 2525 2395
rect 2534 2395 2540 2396
rect 2534 2394 2535 2395
rect 2524 2392 2535 2394
rect 2524 2391 2525 2392
rect 2311 2390 2317 2391
rect 2334 2390 2340 2391
rect 2422 2390 2429 2391
rect 2446 2390 2452 2391
rect 2519 2390 2525 2391
rect 2534 2391 2535 2392
rect 2539 2391 2540 2395
rect 2534 2390 2540 2391
rect 2542 2390 2548 2391
rect 1110 2389 1116 2390
rect 1454 2386 1455 2390
rect 1459 2386 1460 2390
rect 110 2385 116 2386
rect 110 2381 111 2385
rect 115 2381 116 2385
rect 110 2380 116 2381
rect 1326 2385 1332 2386
rect 1454 2385 1460 2386
rect 1558 2386 1559 2390
rect 1563 2386 1564 2390
rect 1558 2385 1564 2386
rect 1662 2386 1663 2390
rect 1667 2386 1668 2390
rect 1662 2385 1668 2386
rect 1758 2386 1759 2390
rect 1763 2386 1764 2390
rect 1758 2385 1764 2386
rect 1854 2386 1855 2390
rect 1859 2386 1860 2390
rect 1854 2385 1860 2386
rect 1942 2386 1943 2390
rect 1947 2386 1948 2390
rect 1942 2385 1948 2386
rect 2038 2386 2039 2390
rect 2043 2386 2044 2390
rect 2038 2385 2044 2386
rect 2134 2386 2135 2390
rect 2139 2386 2140 2390
rect 2134 2385 2140 2386
rect 2230 2386 2231 2390
rect 2235 2386 2236 2390
rect 2230 2385 2236 2386
rect 2334 2386 2335 2390
rect 2339 2386 2340 2390
rect 2334 2385 2340 2386
rect 2446 2386 2447 2390
rect 2451 2386 2452 2390
rect 2446 2385 2452 2386
rect 2542 2386 2543 2390
rect 2547 2386 2548 2390
rect 2542 2385 2548 2386
rect 1326 2381 1327 2385
rect 1331 2381 1332 2385
rect 1326 2380 1332 2381
rect 1366 2381 1372 2382
rect 1366 2377 1367 2381
rect 1371 2377 1372 2381
rect 1366 2376 1372 2377
rect 2582 2381 2588 2382
rect 2582 2377 2583 2381
rect 2587 2377 2588 2381
rect 2582 2376 2588 2377
rect 702 2375 708 2376
rect 702 2371 703 2375
rect 707 2374 708 2375
rect 707 2372 1122 2374
rect 707 2371 708 2372
rect 702 2370 708 2371
rect 110 2368 116 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 230 2367 236 2368
rect 230 2363 231 2367
rect 235 2363 236 2367
rect 318 2367 324 2368
rect 230 2362 236 2363
rect 263 2363 272 2364
rect 263 2359 264 2363
rect 271 2359 272 2363
rect 318 2363 319 2367
rect 323 2363 324 2367
rect 414 2367 420 2368
rect 318 2362 324 2363
rect 351 2363 360 2364
rect 263 2358 272 2359
rect 351 2359 352 2363
rect 359 2359 360 2363
rect 414 2363 415 2367
rect 419 2363 420 2367
rect 510 2367 516 2368
rect 414 2362 420 2363
rect 447 2363 456 2364
rect 351 2358 360 2359
rect 447 2359 448 2363
rect 455 2359 456 2363
rect 510 2363 511 2367
rect 515 2363 516 2367
rect 614 2367 620 2368
rect 510 2362 516 2363
rect 543 2363 552 2364
rect 447 2358 456 2359
rect 543 2359 544 2363
rect 551 2359 552 2363
rect 614 2363 615 2367
rect 619 2363 620 2367
rect 710 2367 716 2368
rect 614 2362 620 2363
rect 646 2363 653 2364
rect 543 2358 552 2359
rect 646 2359 647 2363
rect 652 2359 653 2363
rect 710 2363 711 2367
rect 715 2363 716 2367
rect 806 2367 812 2368
rect 710 2362 716 2363
rect 743 2363 752 2364
rect 646 2358 653 2359
rect 743 2359 744 2363
rect 751 2359 752 2363
rect 806 2363 807 2367
rect 811 2363 812 2367
rect 902 2367 908 2368
rect 806 2362 812 2363
rect 839 2363 848 2364
rect 743 2358 752 2359
rect 839 2359 840 2363
rect 847 2359 848 2363
rect 902 2363 903 2367
rect 907 2363 908 2367
rect 998 2367 1004 2368
rect 902 2362 908 2363
rect 934 2363 941 2364
rect 839 2358 848 2359
rect 934 2359 935 2363
rect 940 2359 941 2363
rect 998 2363 999 2367
rect 1003 2363 1004 2367
rect 1094 2367 1100 2368
rect 998 2362 1004 2363
rect 1031 2363 1037 2364
rect 934 2358 941 2359
rect 1031 2359 1032 2363
rect 1036 2362 1037 2363
rect 1039 2363 1045 2364
rect 1039 2362 1040 2363
rect 1036 2360 1040 2362
rect 1036 2359 1037 2360
rect 1031 2358 1037 2359
rect 1039 2359 1040 2360
rect 1044 2359 1045 2363
rect 1094 2363 1095 2367
rect 1099 2363 1100 2367
rect 1094 2362 1100 2363
rect 1120 2362 1122 2372
rect 2014 2371 2020 2372
rect 1326 2368 1332 2369
rect 1326 2364 1327 2368
rect 1331 2364 1332 2368
rect 2014 2367 2015 2371
rect 2019 2370 2020 2371
rect 2019 2368 2146 2370
rect 2019 2367 2020 2368
rect 2014 2366 2020 2367
rect 1127 2363 1133 2364
rect 1326 2363 1332 2364
rect 1366 2364 1372 2365
rect 1127 2362 1128 2363
rect 1120 2360 1128 2362
rect 1039 2358 1045 2359
rect 1127 2359 1128 2360
rect 1132 2359 1133 2363
rect 1366 2360 1367 2364
rect 1371 2360 1372 2364
rect 1366 2359 1372 2360
rect 1438 2363 1444 2364
rect 1438 2359 1439 2363
rect 1443 2359 1444 2363
rect 1542 2363 1548 2364
rect 1127 2358 1133 2359
rect 1438 2358 1444 2359
rect 1471 2359 1477 2360
rect 1471 2355 1472 2359
rect 1476 2358 1477 2359
rect 1534 2359 1540 2360
rect 1534 2358 1535 2359
rect 1476 2356 1535 2358
rect 1476 2355 1477 2356
rect 1471 2354 1477 2355
rect 1534 2355 1535 2356
rect 1539 2355 1540 2359
rect 1542 2359 1543 2363
rect 1547 2359 1548 2363
rect 1646 2363 1652 2364
rect 1542 2358 1548 2359
rect 1575 2359 1584 2360
rect 1534 2354 1540 2355
rect 1575 2355 1576 2359
rect 1583 2355 1584 2359
rect 1646 2359 1647 2363
rect 1651 2359 1652 2363
rect 1742 2363 1748 2364
rect 1646 2358 1652 2359
rect 1679 2359 1688 2360
rect 1575 2354 1584 2355
rect 1679 2355 1680 2359
rect 1687 2355 1688 2359
rect 1742 2359 1743 2363
rect 1747 2359 1748 2363
rect 1838 2363 1844 2364
rect 1742 2358 1748 2359
rect 1775 2359 1781 2360
rect 1679 2354 1688 2355
rect 1775 2355 1776 2359
rect 1780 2358 1781 2359
rect 1783 2359 1789 2360
rect 1783 2358 1784 2359
rect 1780 2356 1784 2358
rect 1780 2355 1781 2356
rect 1775 2354 1781 2355
rect 1783 2355 1784 2356
rect 1788 2355 1789 2359
rect 1838 2359 1839 2363
rect 1843 2359 1844 2363
rect 1926 2363 1932 2364
rect 1838 2358 1844 2359
rect 1862 2359 1868 2360
rect 1783 2354 1789 2355
rect 1862 2355 1863 2359
rect 1867 2358 1868 2359
rect 1871 2359 1877 2360
rect 1871 2358 1872 2359
rect 1867 2356 1872 2358
rect 1867 2355 1868 2356
rect 1862 2354 1868 2355
rect 1871 2355 1872 2356
rect 1876 2355 1877 2359
rect 1926 2359 1927 2363
rect 1931 2359 1932 2363
rect 2022 2363 2028 2364
rect 1926 2358 1932 2359
rect 1959 2359 1968 2360
rect 1871 2354 1877 2355
rect 1959 2355 1960 2359
rect 1967 2355 1968 2359
rect 2022 2359 2023 2363
rect 2027 2359 2028 2363
rect 2118 2363 2124 2364
rect 2022 2358 2028 2359
rect 2054 2359 2061 2360
rect 1959 2354 1968 2355
rect 2054 2355 2055 2359
rect 2060 2355 2061 2359
rect 2118 2359 2119 2363
rect 2123 2359 2124 2363
rect 2118 2358 2124 2359
rect 2144 2358 2146 2368
rect 2582 2364 2588 2365
rect 2214 2363 2220 2364
rect 2151 2359 2157 2360
rect 2151 2358 2152 2359
rect 2144 2356 2152 2358
rect 2054 2354 2061 2355
rect 2151 2355 2152 2356
rect 2156 2355 2157 2359
rect 2214 2359 2215 2363
rect 2219 2359 2220 2363
rect 2318 2363 2324 2364
rect 2214 2358 2220 2359
rect 2246 2359 2253 2360
rect 2151 2354 2157 2355
rect 2246 2355 2247 2359
rect 2252 2355 2253 2359
rect 2318 2359 2319 2363
rect 2323 2359 2324 2363
rect 2430 2363 2436 2364
rect 2318 2358 2324 2359
rect 2351 2359 2357 2360
rect 2246 2354 2253 2355
rect 2351 2355 2352 2359
rect 2356 2358 2357 2359
rect 2374 2359 2380 2360
rect 2374 2358 2375 2359
rect 2356 2356 2375 2358
rect 2356 2355 2357 2356
rect 2351 2354 2357 2355
rect 2374 2355 2375 2356
rect 2379 2355 2380 2359
rect 2430 2359 2431 2363
rect 2435 2359 2436 2363
rect 2526 2363 2532 2364
rect 2430 2358 2436 2359
rect 2463 2359 2469 2360
rect 2463 2358 2464 2359
rect 2440 2356 2464 2358
rect 2374 2354 2380 2355
rect 2438 2355 2444 2356
rect 2438 2351 2439 2355
rect 2443 2351 2444 2355
rect 2463 2355 2464 2356
rect 2468 2355 2469 2359
rect 2526 2359 2527 2363
rect 2531 2359 2532 2363
rect 2582 2360 2583 2364
rect 2587 2360 2588 2364
rect 2526 2358 2532 2359
rect 2558 2359 2565 2360
rect 2582 2359 2588 2360
rect 2463 2354 2469 2355
rect 2558 2355 2559 2359
rect 2564 2355 2565 2359
rect 2558 2354 2565 2355
rect 2438 2350 2444 2351
rect 166 2343 172 2344
rect 166 2339 167 2343
rect 171 2342 172 2343
rect 734 2343 740 2344
rect 171 2340 626 2342
rect 171 2339 172 2340
rect 166 2338 172 2339
rect 191 2335 197 2336
rect 158 2333 164 2334
rect 110 2332 116 2333
rect 110 2328 111 2332
rect 115 2328 116 2332
rect 158 2329 159 2333
rect 163 2329 164 2333
rect 191 2331 192 2335
rect 196 2334 197 2335
rect 254 2335 260 2336
rect 254 2334 255 2335
rect 196 2332 255 2334
rect 196 2331 197 2332
rect 191 2330 197 2331
rect 254 2331 255 2332
rect 259 2331 260 2335
rect 295 2335 301 2336
rect 254 2330 260 2331
rect 262 2333 268 2334
rect 158 2328 164 2329
rect 262 2329 263 2333
rect 267 2329 268 2333
rect 295 2331 296 2335
rect 300 2334 301 2335
rect 346 2335 352 2336
rect 346 2334 347 2335
rect 300 2332 347 2334
rect 300 2331 301 2332
rect 295 2330 301 2331
rect 346 2331 347 2332
rect 351 2331 352 2335
rect 407 2335 413 2336
rect 346 2330 352 2331
rect 374 2333 380 2334
rect 262 2328 268 2329
rect 374 2329 375 2333
rect 379 2329 380 2333
rect 407 2331 408 2335
rect 412 2334 413 2335
rect 478 2335 484 2336
rect 478 2334 479 2335
rect 412 2332 479 2334
rect 412 2331 413 2332
rect 407 2330 413 2331
rect 478 2331 479 2332
rect 483 2331 484 2335
rect 519 2335 525 2336
rect 478 2330 484 2331
rect 486 2333 492 2334
rect 374 2328 380 2329
rect 486 2329 487 2333
rect 491 2329 492 2333
rect 519 2331 520 2335
rect 524 2334 525 2335
rect 590 2335 596 2336
rect 590 2334 591 2335
rect 524 2332 591 2334
rect 524 2331 525 2332
rect 519 2330 525 2331
rect 590 2331 591 2332
rect 595 2331 596 2335
rect 624 2334 626 2340
rect 734 2339 735 2343
rect 739 2342 740 2343
rect 739 2340 1226 2342
rect 739 2339 740 2340
rect 734 2338 740 2339
rect 631 2335 637 2336
rect 631 2334 632 2335
rect 590 2330 596 2331
rect 598 2333 604 2334
rect 486 2328 492 2329
rect 598 2329 599 2333
rect 603 2329 604 2333
rect 624 2332 632 2334
rect 631 2331 632 2332
rect 636 2331 637 2335
rect 743 2335 749 2336
rect 631 2330 637 2331
rect 710 2333 716 2334
rect 598 2328 604 2329
rect 710 2329 711 2333
rect 715 2329 716 2333
rect 743 2331 744 2335
rect 748 2334 749 2335
rect 806 2335 812 2336
rect 806 2334 807 2335
rect 748 2332 807 2334
rect 748 2331 749 2332
rect 743 2330 749 2331
rect 806 2331 807 2332
rect 811 2331 812 2335
rect 847 2335 853 2336
rect 806 2330 812 2331
rect 814 2333 820 2334
rect 710 2328 716 2329
rect 814 2329 815 2333
rect 819 2329 820 2333
rect 847 2331 848 2335
rect 852 2334 853 2335
rect 902 2335 908 2336
rect 902 2334 903 2335
rect 852 2332 903 2334
rect 852 2331 853 2332
rect 847 2330 853 2331
rect 902 2331 903 2332
rect 907 2331 908 2335
rect 943 2335 949 2336
rect 902 2330 908 2331
rect 910 2333 916 2334
rect 814 2328 820 2329
rect 910 2329 911 2333
rect 915 2329 916 2333
rect 943 2331 944 2335
rect 948 2334 949 2335
rect 967 2335 973 2336
rect 967 2334 968 2335
rect 948 2332 968 2334
rect 948 2331 949 2332
rect 943 2330 949 2331
rect 967 2331 968 2332
rect 972 2331 973 2335
rect 1039 2335 1045 2336
rect 967 2330 973 2331
rect 1006 2333 1012 2334
rect 910 2328 916 2329
rect 1006 2329 1007 2333
rect 1011 2329 1012 2333
rect 1039 2331 1040 2335
rect 1044 2334 1045 2335
rect 1094 2335 1100 2336
rect 1094 2334 1095 2335
rect 1044 2332 1095 2334
rect 1044 2331 1045 2332
rect 1039 2330 1045 2331
rect 1094 2331 1095 2332
rect 1099 2331 1100 2335
rect 1135 2335 1141 2336
rect 1094 2330 1100 2331
rect 1102 2333 1108 2334
rect 1006 2328 1012 2329
rect 1102 2329 1103 2333
rect 1107 2329 1108 2333
rect 1135 2331 1136 2335
rect 1140 2334 1141 2335
rect 1190 2335 1196 2336
rect 1190 2334 1191 2335
rect 1140 2332 1191 2334
rect 1140 2331 1141 2332
rect 1135 2330 1141 2331
rect 1190 2331 1191 2332
rect 1195 2331 1196 2335
rect 1224 2334 1226 2340
rect 1446 2339 1452 2340
rect 1231 2335 1237 2336
rect 1231 2334 1232 2335
rect 1190 2330 1196 2331
rect 1198 2333 1204 2334
rect 1102 2328 1108 2329
rect 1198 2329 1199 2333
rect 1203 2329 1204 2333
rect 1224 2332 1232 2334
rect 1231 2331 1232 2332
rect 1236 2331 1237 2335
rect 1446 2335 1447 2339
rect 1451 2338 1452 2339
rect 2126 2339 2132 2340
rect 1451 2336 1538 2338
rect 1451 2335 1452 2336
rect 1446 2334 1452 2335
rect 1231 2330 1237 2331
rect 1326 2332 1332 2333
rect 1198 2328 1204 2329
rect 1326 2328 1327 2332
rect 1331 2328 1332 2332
rect 1431 2331 1437 2332
rect 1398 2329 1404 2330
rect 110 2327 116 2328
rect 1326 2327 1332 2328
rect 1366 2328 1372 2329
rect 1366 2324 1367 2328
rect 1371 2324 1372 2328
rect 1398 2325 1399 2329
rect 1403 2325 1404 2329
rect 1431 2327 1432 2331
rect 1436 2330 1437 2331
rect 1446 2331 1452 2332
rect 1446 2330 1447 2331
rect 1436 2328 1447 2330
rect 1436 2327 1437 2328
rect 1431 2326 1437 2327
rect 1446 2327 1447 2328
rect 1451 2327 1452 2331
rect 1487 2331 1493 2332
rect 1446 2326 1452 2327
rect 1454 2329 1460 2330
rect 1398 2324 1404 2325
rect 1454 2325 1455 2329
rect 1459 2325 1460 2329
rect 1487 2327 1488 2331
rect 1492 2330 1493 2331
rect 1502 2331 1508 2332
rect 1502 2330 1503 2331
rect 1492 2328 1503 2330
rect 1492 2327 1493 2328
rect 1487 2326 1493 2327
rect 1502 2327 1503 2328
rect 1507 2327 1508 2331
rect 1536 2330 1538 2336
rect 2126 2335 2127 2339
rect 2131 2338 2132 2339
rect 2131 2336 2250 2338
rect 2131 2335 2132 2336
rect 2126 2334 2132 2335
rect 1543 2331 1549 2332
rect 1543 2330 1544 2331
rect 1502 2326 1508 2327
rect 1510 2329 1516 2330
rect 1454 2324 1460 2325
rect 1510 2325 1511 2329
rect 1515 2325 1516 2329
rect 1536 2328 1544 2330
rect 1543 2327 1544 2328
rect 1548 2327 1549 2331
rect 1599 2331 1605 2332
rect 1543 2326 1549 2327
rect 1566 2329 1572 2330
rect 1510 2324 1516 2325
rect 1566 2325 1567 2329
rect 1571 2325 1572 2329
rect 1599 2327 1600 2331
rect 1604 2330 1605 2331
rect 1630 2331 1636 2332
rect 1630 2330 1631 2331
rect 1604 2328 1631 2330
rect 1604 2327 1605 2328
rect 1599 2326 1605 2327
rect 1630 2327 1631 2328
rect 1635 2327 1636 2331
rect 1671 2331 1677 2332
rect 1630 2326 1636 2327
rect 1638 2329 1644 2330
rect 1566 2324 1572 2325
rect 1638 2325 1639 2329
rect 1643 2325 1644 2329
rect 1671 2327 1672 2331
rect 1676 2330 1677 2331
rect 1718 2331 1724 2332
rect 1718 2330 1719 2331
rect 1676 2328 1719 2330
rect 1676 2327 1677 2328
rect 1671 2326 1677 2327
rect 1718 2327 1719 2328
rect 1723 2327 1724 2331
rect 1759 2331 1765 2332
rect 1718 2326 1724 2327
rect 1726 2329 1732 2330
rect 1638 2324 1644 2325
rect 1726 2325 1727 2329
rect 1731 2325 1732 2329
rect 1759 2327 1760 2331
rect 1764 2330 1765 2331
rect 1814 2331 1820 2332
rect 1814 2330 1815 2331
rect 1764 2328 1815 2330
rect 1764 2327 1765 2328
rect 1759 2326 1765 2327
rect 1814 2327 1815 2328
rect 1819 2327 1820 2331
rect 1855 2331 1861 2332
rect 1814 2326 1820 2327
rect 1822 2329 1828 2330
rect 1726 2324 1732 2325
rect 1822 2325 1823 2329
rect 1827 2325 1828 2329
rect 1855 2327 1856 2331
rect 1860 2330 1861 2331
rect 1934 2331 1940 2332
rect 1934 2330 1935 2331
rect 1860 2328 1935 2330
rect 1860 2327 1861 2328
rect 1855 2326 1861 2327
rect 1934 2327 1935 2328
rect 1939 2327 1940 2331
rect 1975 2331 1981 2332
rect 1934 2326 1940 2327
rect 1942 2329 1948 2330
rect 1822 2324 1828 2325
rect 1942 2325 1943 2329
rect 1947 2325 1948 2329
rect 1975 2327 1976 2331
rect 1980 2330 1981 2331
rect 2070 2331 2076 2332
rect 2070 2330 2071 2331
rect 1980 2328 2071 2330
rect 1980 2327 1981 2328
rect 1975 2326 1981 2327
rect 2070 2327 2071 2328
rect 2075 2327 2076 2331
rect 2111 2331 2117 2332
rect 2070 2326 2076 2327
rect 2078 2329 2084 2330
rect 1942 2324 1948 2325
rect 2078 2325 2079 2329
rect 2083 2325 2084 2329
rect 2111 2327 2112 2331
rect 2116 2330 2117 2331
rect 2214 2331 2220 2332
rect 2214 2330 2215 2331
rect 2116 2328 2215 2330
rect 2116 2327 2117 2328
rect 2111 2326 2117 2327
rect 2214 2327 2215 2328
rect 2219 2327 2220 2331
rect 2248 2330 2250 2336
rect 2534 2335 2540 2336
rect 2255 2331 2261 2332
rect 2255 2330 2256 2331
rect 2214 2326 2220 2327
rect 2222 2329 2228 2330
rect 2078 2324 2084 2325
rect 2222 2325 2223 2329
rect 2227 2325 2228 2329
rect 2248 2328 2256 2330
rect 2255 2327 2256 2328
rect 2260 2327 2261 2331
rect 2414 2331 2421 2332
rect 2255 2326 2261 2327
rect 2382 2329 2388 2330
rect 2222 2324 2228 2325
rect 2382 2325 2383 2329
rect 2387 2325 2388 2329
rect 2414 2327 2415 2331
rect 2420 2327 2421 2331
rect 2534 2331 2535 2335
rect 2539 2334 2540 2335
rect 2539 2332 2554 2334
rect 2539 2331 2540 2332
rect 2534 2330 2540 2331
rect 2552 2330 2554 2332
rect 2559 2331 2565 2332
rect 2559 2330 2560 2331
rect 2414 2326 2421 2327
rect 2526 2329 2532 2330
rect 2382 2324 2388 2325
rect 2526 2325 2527 2329
rect 2531 2325 2532 2329
rect 2552 2328 2560 2330
rect 2559 2327 2560 2328
rect 2564 2327 2565 2331
rect 2559 2326 2565 2327
rect 2582 2328 2588 2329
rect 2526 2324 2532 2325
rect 2582 2324 2583 2328
rect 2587 2324 2588 2328
rect 1366 2323 1372 2324
rect 2582 2323 2588 2324
rect 110 2315 116 2316
rect 110 2311 111 2315
rect 115 2311 116 2315
rect 110 2310 116 2311
rect 1326 2315 1332 2316
rect 1326 2311 1327 2315
rect 1331 2311 1332 2315
rect 1326 2310 1332 2311
rect 1366 2311 1372 2312
rect 1366 2307 1367 2311
rect 1371 2307 1372 2311
rect 174 2306 180 2307
rect 174 2302 175 2306
rect 179 2302 180 2306
rect 174 2301 180 2302
rect 278 2306 284 2307
rect 278 2302 279 2306
rect 283 2302 284 2306
rect 278 2301 284 2302
rect 390 2306 396 2307
rect 390 2302 391 2306
rect 395 2302 396 2306
rect 390 2301 396 2302
rect 502 2306 508 2307
rect 502 2302 503 2306
rect 507 2302 508 2306
rect 502 2301 508 2302
rect 614 2306 620 2307
rect 614 2302 615 2306
rect 619 2302 620 2306
rect 614 2301 620 2302
rect 726 2306 732 2307
rect 726 2302 727 2306
rect 731 2302 732 2306
rect 726 2301 732 2302
rect 830 2306 836 2307
rect 830 2302 831 2306
rect 835 2302 836 2306
rect 830 2301 836 2302
rect 926 2306 932 2307
rect 926 2302 927 2306
rect 931 2302 932 2306
rect 926 2301 932 2302
rect 1022 2306 1028 2307
rect 1022 2302 1023 2306
rect 1027 2302 1028 2306
rect 1022 2301 1028 2302
rect 1118 2306 1124 2307
rect 1118 2302 1119 2306
rect 1123 2302 1124 2306
rect 1118 2301 1124 2302
rect 1214 2306 1220 2307
rect 1366 2306 1372 2307
rect 2582 2311 2588 2312
rect 2582 2307 2583 2311
rect 2587 2307 2588 2311
rect 2582 2306 2588 2307
rect 1214 2302 1215 2306
rect 1219 2302 1220 2306
rect 1214 2301 1220 2302
rect 1414 2302 1420 2303
rect 151 2299 157 2300
rect 151 2295 152 2299
rect 156 2298 157 2299
rect 166 2299 172 2300
rect 166 2298 167 2299
rect 156 2296 167 2298
rect 156 2295 157 2296
rect 151 2294 157 2295
rect 166 2295 167 2296
rect 171 2295 172 2299
rect 166 2294 172 2295
rect 254 2299 261 2300
rect 254 2295 255 2299
rect 260 2295 261 2299
rect 254 2294 261 2295
rect 354 2299 360 2300
rect 354 2295 355 2299
rect 359 2298 360 2299
rect 367 2299 373 2300
rect 367 2298 368 2299
rect 359 2296 368 2298
rect 359 2295 360 2296
rect 354 2294 360 2295
rect 367 2295 368 2296
rect 372 2295 373 2299
rect 367 2294 373 2295
rect 478 2299 485 2300
rect 478 2295 479 2299
rect 484 2295 485 2299
rect 478 2294 485 2295
rect 590 2299 597 2300
rect 590 2295 591 2299
rect 596 2295 597 2299
rect 590 2294 597 2295
rect 703 2299 709 2300
rect 703 2295 704 2299
rect 708 2298 709 2299
rect 734 2299 740 2300
rect 734 2298 735 2299
rect 708 2296 735 2298
rect 708 2295 709 2296
rect 703 2294 709 2295
rect 734 2295 735 2296
rect 739 2295 740 2299
rect 734 2294 740 2295
rect 806 2299 813 2300
rect 806 2295 807 2299
rect 812 2295 813 2299
rect 806 2294 813 2295
rect 902 2299 909 2300
rect 902 2295 903 2299
rect 908 2295 909 2299
rect 902 2294 909 2295
rect 999 2299 1005 2300
rect 999 2295 1000 2299
rect 1004 2298 1005 2299
rect 1014 2299 1020 2300
rect 1014 2298 1015 2299
rect 1004 2296 1015 2298
rect 1004 2295 1005 2296
rect 999 2294 1005 2295
rect 1014 2295 1015 2296
rect 1019 2295 1020 2299
rect 1014 2294 1020 2295
rect 1094 2299 1101 2300
rect 1094 2295 1095 2299
rect 1100 2295 1101 2299
rect 1094 2294 1101 2295
rect 1190 2299 1197 2300
rect 1190 2295 1191 2299
rect 1196 2295 1197 2299
rect 1414 2298 1415 2302
rect 1419 2298 1420 2302
rect 1414 2297 1420 2298
rect 1470 2302 1476 2303
rect 1470 2298 1471 2302
rect 1475 2298 1476 2302
rect 1470 2297 1476 2298
rect 1526 2302 1532 2303
rect 1526 2298 1527 2302
rect 1531 2298 1532 2302
rect 1526 2297 1532 2298
rect 1582 2302 1588 2303
rect 1582 2298 1583 2302
rect 1587 2298 1588 2302
rect 1582 2297 1588 2298
rect 1654 2302 1660 2303
rect 1654 2298 1655 2302
rect 1659 2298 1660 2302
rect 1654 2297 1660 2298
rect 1742 2302 1748 2303
rect 1742 2298 1743 2302
rect 1747 2298 1748 2302
rect 1742 2297 1748 2298
rect 1838 2302 1844 2303
rect 1838 2298 1839 2302
rect 1843 2298 1844 2302
rect 1838 2297 1844 2298
rect 1958 2302 1964 2303
rect 1958 2298 1959 2302
rect 1963 2298 1964 2302
rect 1958 2297 1964 2298
rect 2094 2302 2100 2303
rect 2094 2298 2095 2302
rect 2099 2298 2100 2302
rect 2094 2297 2100 2298
rect 2238 2302 2244 2303
rect 2238 2298 2239 2302
rect 2243 2298 2244 2302
rect 2238 2297 2244 2298
rect 2398 2302 2404 2303
rect 2398 2298 2399 2302
rect 2403 2298 2404 2302
rect 2398 2297 2404 2298
rect 2542 2302 2548 2303
rect 2542 2298 2543 2302
rect 2547 2298 2548 2302
rect 2542 2297 2548 2298
rect 1190 2294 1197 2295
rect 1306 2295 1312 2296
rect 646 2291 652 2292
rect 646 2290 647 2291
rect 319 2288 647 2290
rect 319 2286 321 2288
rect 646 2287 647 2288
rect 651 2287 652 2291
rect 1110 2291 1116 2292
rect 1110 2290 1111 2291
rect 646 2286 652 2287
rect 760 2288 1111 2290
rect 240 2284 321 2286
rect 134 2283 141 2284
rect 134 2279 135 2283
rect 140 2279 141 2283
rect 223 2283 229 2284
rect 223 2279 224 2283
rect 228 2282 229 2283
rect 240 2282 242 2284
rect 228 2280 242 2282
rect 346 2283 357 2284
rect 228 2279 229 2280
rect 346 2279 347 2283
rect 351 2279 352 2283
rect 356 2279 357 2283
rect 442 2283 448 2284
rect 442 2279 443 2283
rect 447 2282 448 2283
rect 487 2283 493 2284
rect 487 2282 488 2283
rect 447 2280 488 2282
rect 447 2279 448 2280
rect 134 2278 141 2279
rect 158 2278 164 2279
rect 223 2278 229 2279
rect 246 2278 252 2279
rect 346 2278 357 2279
rect 374 2278 380 2279
rect 442 2278 448 2279
rect 487 2279 488 2280
rect 492 2279 493 2283
rect 530 2283 536 2284
rect 530 2279 531 2283
rect 535 2282 536 2283
rect 615 2283 621 2284
rect 615 2282 616 2283
rect 535 2280 616 2282
rect 535 2279 536 2280
rect 487 2278 493 2279
rect 510 2278 516 2279
rect 530 2278 536 2279
rect 615 2279 616 2280
rect 620 2279 621 2283
rect 743 2283 749 2284
rect 743 2279 744 2283
rect 748 2282 749 2283
rect 760 2282 762 2288
rect 1110 2287 1111 2288
rect 1115 2287 1116 2291
rect 1306 2291 1307 2295
rect 1311 2294 1312 2295
rect 1391 2295 1397 2296
rect 1391 2294 1392 2295
rect 1311 2292 1392 2294
rect 1311 2291 1312 2292
rect 1306 2290 1312 2291
rect 1391 2291 1392 2292
rect 1396 2291 1397 2295
rect 1391 2290 1397 2291
rect 1446 2295 1453 2296
rect 1446 2291 1447 2295
rect 1452 2291 1453 2295
rect 1446 2290 1453 2291
rect 1502 2295 1509 2296
rect 1502 2291 1503 2295
rect 1508 2291 1509 2295
rect 1502 2290 1509 2291
rect 1534 2295 1540 2296
rect 1534 2291 1535 2295
rect 1539 2294 1540 2295
rect 1559 2295 1565 2296
rect 1559 2294 1560 2295
rect 1539 2292 1560 2294
rect 1539 2291 1540 2292
rect 1534 2290 1540 2291
rect 1559 2291 1560 2292
rect 1564 2291 1565 2295
rect 1559 2290 1565 2291
rect 1630 2295 1637 2296
rect 1630 2291 1631 2295
rect 1636 2291 1637 2295
rect 1630 2290 1637 2291
rect 1718 2295 1725 2296
rect 1718 2291 1719 2295
rect 1724 2291 1725 2295
rect 1718 2290 1725 2291
rect 1815 2295 1821 2296
rect 1815 2291 1816 2295
rect 1820 2294 1821 2295
rect 1862 2295 1868 2296
rect 1862 2294 1863 2295
rect 1820 2292 1863 2294
rect 1820 2291 1821 2292
rect 1815 2290 1821 2291
rect 1862 2291 1863 2292
rect 1867 2291 1868 2295
rect 1862 2290 1868 2291
rect 1934 2295 1941 2296
rect 1934 2291 1935 2295
rect 1940 2291 1941 2295
rect 1934 2290 1941 2291
rect 2070 2295 2077 2296
rect 2070 2291 2071 2295
rect 2076 2291 2077 2295
rect 2070 2290 2077 2291
rect 2214 2295 2221 2296
rect 2214 2291 2215 2295
rect 2220 2291 2221 2295
rect 2214 2290 2221 2291
rect 2374 2295 2381 2296
rect 2374 2291 2375 2295
rect 2380 2291 2381 2295
rect 2374 2290 2381 2291
rect 2519 2295 2525 2296
rect 2519 2291 2520 2295
rect 2524 2294 2525 2295
rect 2558 2295 2564 2296
rect 2558 2294 2559 2295
rect 2524 2292 2559 2294
rect 2524 2291 2525 2292
rect 2519 2290 2525 2291
rect 2558 2291 2559 2292
rect 2563 2291 2564 2295
rect 2558 2290 2564 2291
rect 1110 2286 1116 2287
rect 748 2280 762 2282
rect 822 2283 828 2284
rect 748 2279 749 2280
rect 822 2279 823 2283
rect 827 2282 828 2283
rect 863 2283 869 2284
rect 863 2282 864 2283
rect 827 2280 864 2282
rect 827 2279 828 2280
rect 615 2278 621 2279
rect 638 2278 644 2279
rect 743 2278 749 2279
rect 766 2278 772 2279
rect 822 2278 828 2279
rect 863 2279 864 2280
rect 868 2279 869 2283
rect 906 2283 912 2284
rect 906 2279 907 2283
rect 911 2282 912 2283
rect 975 2283 981 2284
rect 975 2282 976 2283
rect 911 2280 976 2282
rect 911 2279 912 2280
rect 863 2278 869 2279
rect 886 2278 892 2279
rect 906 2278 912 2279
rect 975 2279 976 2280
rect 980 2279 981 2283
rect 1078 2283 1085 2284
rect 1078 2279 1079 2283
rect 1084 2279 1085 2283
rect 1183 2283 1189 2284
rect 1183 2279 1184 2283
rect 1188 2282 1189 2283
rect 1198 2283 1204 2284
rect 1198 2282 1199 2283
rect 1188 2280 1199 2282
rect 1188 2279 1189 2280
rect 975 2278 981 2279
rect 998 2278 1004 2279
rect 1078 2278 1085 2279
rect 1102 2278 1108 2279
rect 1183 2278 1189 2279
rect 1198 2279 1199 2280
rect 1203 2279 1204 2283
rect 1263 2283 1269 2284
rect 1263 2279 1264 2283
rect 1268 2282 1269 2283
rect 1278 2283 1284 2284
rect 1278 2282 1279 2283
rect 1268 2280 1279 2282
rect 1268 2279 1269 2280
rect 1198 2278 1204 2279
rect 1206 2278 1212 2279
rect 1263 2278 1269 2279
rect 1278 2279 1279 2280
rect 1283 2279 1284 2283
rect 2414 2283 2420 2284
rect 2414 2282 2415 2283
rect 1961 2280 2415 2282
rect 1662 2279 1668 2280
rect 1278 2278 1284 2279
rect 1286 2278 1292 2279
rect 1662 2278 1663 2279
rect 158 2274 159 2278
rect 163 2274 164 2278
rect 158 2273 164 2274
rect 246 2274 247 2278
rect 251 2274 252 2278
rect 246 2273 252 2274
rect 374 2274 375 2278
rect 379 2274 380 2278
rect 374 2273 380 2274
rect 510 2274 511 2278
rect 515 2274 516 2278
rect 510 2273 516 2274
rect 638 2274 639 2278
rect 643 2274 644 2278
rect 638 2273 644 2274
rect 766 2274 767 2278
rect 771 2274 772 2278
rect 766 2273 772 2274
rect 886 2274 887 2278
rect 891 2274 892 2278
rect 886 2273 892 2274
rect 998 2274 999 2278
rect 1003 2274 1004 2278
rect 998 2273 1004 2274
rect 1102 2274 1103 2278
rect 1107 2274 1108 2278
rect 1102 2273 1108 2274
rect 1206 2274 1207 2278
rect 1211 2274 1212 2278
rect 1206 2273 1212 2274
rect 1286 2274 1287 2278
rect 1291 2274 1292 2278
rect 1608 2276 1663 2278
rect 1286 2273 1292 2274
rect 1390 2275 1397 2276
rect 1390 2271 1391 2275
rect 1396 2271 1397 2275
rect 1471 2275 1477 2276
rect 1471 2271 1472 2275
rect 1476 2274 1477 2275
rect 1486 2275 1492 2276
rect 1486 2274 1487 2275
rect 1476 2272 1487 2274
rect 1476 2271 1477 2272
rect 1390 2270 1397 2271
rect 1414 2270 1420 2271
rect 1471 2270 1477 2271
rect 1486 2271 1487 2272
rect 1491 2271 1492 2275
rect 1591 2275 1597 2276
rect 1591 2271 1592 2275
rect 1596 2274 1597 2275
rect 1608 2274 1610 2276
rect 1662 2275 1663 2276
rect 1667 2275 1668 2279
rect 1662 2274 1668 2275
rect 1710 2275 1717 2276
rect 1596 2272 1610 2274
rect 1596 2271 1597 2272
rect 1710 2271 1711 2275
rect 1716 2271 1717 2275
rect 1814 2275 1820 2276
rect 1814 2271 1815 2275
rect 1819 2274 1820 2275
rect 1831 2275 1837 2276
rect 1831 2274 1832 2275
rect 1819 2272 1832 2274
rect 1819 2271 1820 2272
rect 1486 2270 1492 2271
rect 1494 2270 1500 2271
rect 1591 2270 1597 2271
rect 1614 2270 1620 2271
rect 1710 2270 1717 2271
rect 1734 2270 1740 2271
rect 1814 2270 1820 2271
rect 1831 2271 1832 2272
rect 1836 2271 1837 2275
rect 1943 2275 1949 2276
rect 1943 2271 1944 2275
rect 1948 2274 1949 2275
rect 1961 2274 1963 2280
rect 2414 2279 2415 2280
rect 2419 2279 2420 2283
rect 2414 2278 2420 2279
rect 1948 2272 1963 2274
rect 1986 2275 1992 2276
rect 1948 2271 1949 2272
rect 1986 2271 1987 2275
rect 1991 2274 1992 2275
rect 2047 2275 2053 2276
rect 2047 2274 2048 2275
rect 1991 2272 2048 2274
rect 1991 2271 1992 2272
rect 1831 2270 1837 2271
rect 1854 2270 1860 2271
rect 1943 2270 1949 2271
rect 1966 2270 1972 2271
rect 1986 2270 1992 2271
rect 2047 2271 2048 2272
rect 2052 2271 2053 2275
rect 2095 2275 2101 2276
rect 2095 2271 2096 2275
rect 2100 2274 2101 2275
rect 2143 2275 2149 2276
rect 2143 2274 2144 2275
rect 2100 2272 2144 2274
rect 2100 2271 2101 2272
rect 2047 2270 2053 2271
rect 2070 2270 2076 2271
rect 2095 2270 2101 2271
rect 2143 2271 2144 2272
rect 2148 2271 2149 2275
rect 2186 2275 2192 2276
rect 2186 2271 2187 2275
rect 2191 2274 2192 2275
rect 2231 2275 2237 2276
rect 2231 2274 2232 2275
rect 2191 2272 2232 2274
rect 2191 2271 2192 2272
rect 2143 2270 2149 2271
rect 2166 2270 2172 2271
rect 2186 2270 2192 2271
rect 2231 2271 2232 2272
rect 2236 2271 2237 2275
rect 2274 2275 2280 2276
rect 2274 2271 2275 2275
rect 2279 2274 2280 2275
rect 2311 2275 2317 2276
rect 2311 2274 2312 2275
rect 2279 2272 2312 2274
rect 2279 2271 2280 2272
rect 2231 2270 2237 2271
rect 2254 2270 2260 2271
rect 2274 2270 2280 2271
rect 2311 2271 2312 2272
rect 2316 2271 2317 2275
rect 2382 2275 2389 2276
rect 2382 2271 2383 2275
rect 2388 2271 2389 2275
rect 2414 2275 2420 2276
rect 2414 2271 2415 2275
rect 2419 2274 2420 2275
rect 2463 2275 2469 2276
rect 2463 2274 2464 2275
rect 2419 2272 2464 2274
rect 2419 2271 2420 2272
rect 2311 2270 2317 2271
rect 2334 2270 2340 2271
rect 2382 2270 2389 2271
rect 2406 2270 2412 2271
rect 2414 2270 2420 2271
rect 2463 2271 2464 2272
rect 2468 2271 2469 2275
rect 2506 2275 2512 2276
rect 2506 2271 2507 2275
rect 2511 2274 2512 2275
rect 2519 2275 2525 2276
rect 2519 2274 2520 2275
rect 2511 2272 2520 2274
rect 2511 2271 2512 2272
rect 2463 2270 2469 2271
rect 2486 2270 2492 2271
rect 2506 2270 2512 2271
rect 2519 2271 2520 2272
rect 2524 2271 2525 2275
rect 2519 2270 2525 2271
rect 2542 2270 2548 2271
rect 110 2269 116 2270
rect 110 2265 111 2269
rect 115 2265 116 2269
rect 110 2264 116 2265
rect 1326 2269 1332 2270
rect 1326 2265 1327 2269
rect 1331 2265 1332 2269
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1494 2266 1495 2270
rect 1499 2266 1500 2270
rect 1494 2265 1500 2266
rect 1614 2266 1615 2270
rect 1619 2266 1620 2270
rect 1614 2265 1620 2266
rect 1734 2266 1735 2270
rect 1739 2266 1740 2270
rect 1734 2265 1740 2266
rect 1854 2266 1855 2270
rect 1859 2266 1860 2270
rect 1854 2265 1860 2266
rect 1966 2266 1967 2270
rect 1971 2266 1972 2270
rect 1966 2265 1972 2266
rect 2070 2266 2071 2270
rect 2075 2266 2076 2270
rect 2070 2265 2076 2266
rect 2166 2266 2167 2270
rect 2171 2266 2172 2270
rect 2166 2265 2172 2266
rect 2254 2266 2255 2270
rect 2259 2266 2260 2270
rect 2254 2265 2260 2266
rect 2334 2266 2335 2270
rect 2339 2266 2340 2270
rect 2334 2265 2340 2266
rect 2406 2266 2407 2270
rect 2411 2266 2412 2270
rect 2406 2265 2412 2266
rect 2486 2266 2487 2270
rect 2491 2266 2492 2270
rect 2486 2265 2492 2266
rect 2542 2266 2543 2270
rect 2547 2266 2548 2270
rect 2542 2265 2548 2266
rect 1326 2264 1332 2265
rect 1366 2261 1372 2262
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2258 140 2259
rect 1078 2259 1084 2260
rect 139 2256 258 2258
rect 139 2255 140 2256
rect 134 2254 140 2255
rect 110 2252 116 2253
rect 110 2248 111 2252
rect 115 2248 116 2252
rect 110 2247 116 2248
rect 142 2251 148 2252
rect 142 2247 143 2251
rect 147 2247 148 2251
rect 230 2251 236 2252
rect 142 2246 148 2247
rect 166 2247 172 2248
rect 166 2243 167 2247
rect 171 2246 172 2247
rect 175 2247 181 2248
rect 175 2246 176 2247
rect 171 2244 176 2246
rect 171 2243 172 2244
rect 166 2242 172 2243
rect 175 2243 176 2244
rect 180 2243 181 2247
rect 230 2247 231 2251
rect 235 2247 236 2251
rect 230 2246 236 2247
rect 256 2246 258 2256
rect 1078 2255 1079 2259
rect 1083 2258 1084 2259
rect 1083 2256 1218 2258
rect 1366 2257 1367 2261
rect 1371 2257 1372 2261
rect 1366 2256 1372 2257
rect 2582 2261 2588 2262
rect 2582 2257 2583 2261
rect 2587 2257 2588 2261
rect 2582 2256 2588 2257
rect 1083 2255 1084 2256
rect 1078 2254 1084 2255
rect 358 2251 364 2252
rect 263 2247 269 2248
rect 263 2246 264 2247
rect 256 2244 264 2246
rect 175 2242 181 2243
rect 263 2243 264 2244
rect 268 2243 269 2247
rect 358 2247 359 2251
rect 363 2247 364 2251
rect 442 2251 448 2252
rect 442 2250 443 2251
rect 358 2246 364 2247
rect 391 2249 443 2250
rect 391 2245 392 2249
rect 396 2248 443 2249
rect 396 2245 397 2248
rect 442 2247 443 2248
rect 447 2247 448 2251
rect 442 2246 448 2247
rect 494 2251 500 2252
rect 494 2247 495 2251
rect 499 2247 500 2251
rect 622 2251 628 2252
rect 494 2246 500 2247
rect 527 2247 536 2248
rect 391 2244 397 2245
rect 263 2242 269 2243
rect 527 2243 528 2247
rect 535 2243 536 2247
rect 622 2247 623 2251
rect 627 2247 628 2251
rect 750 2251 756 2252
rect 622 2246 628 2247
rect 646 2247 652 2248
rect 527 2242 536 2243
rect 646 2243 647 2247
rect 651 2246 652 2247
rect 655 2247 661 2248
rect 655 2246 656 2247
rect 651 2244 656 2246
rect 651 2243 652 2244
rect 646 2242 652 2243
rect 655 2243 656 2244
rect 660 2243 661 2247
rect 750 2247 751 2251
rect 755 2247 756 2251
rect 870 2251 876 2252
rect 750 2246 756 2247
rect 783 2247 789 2248
rect 655 2242 661 2243
rect 783 2243 784 2247
rect 788 2246 789 2247
rect 822 2247 828 2248
rect 822 2246 823 2247
rect 788 2244 823 2246
rect 788 2243 789 2244
rect 783 2242 789 2243
rect 822 2243 823 2244
rect 827 2243 828 2247
rect 870 2247 871 2251
rect 875 2247 876 2251
rect 982 2251 988 2252
rect 870 2246 876 2247
rect 903 2247 912 2248
rect 822 2242 828 2243
rect 903 2243 904 2247
rect 911 2243 912 2247
rect 982 2247 983 2251
rect 987 2247 988 2251
rect 1086 2251 1092 2252
rect 982 2246 988 2247
rect 1014 2247 1021 2248
rect 903 2242 912 2243
rect 1014 2243 1015 2247
rect 1020 2243 1021 2247
rect 1086 2247 1087 2251
rect 1091 2247 1092 2251
rect 1190 2251 1196 2252
rect 1086 2246 1092 2247
rect 1110 2247 1116 2248
rect 1014 2242 1021 2243
rect 1110 2243 1111 2247
rect 1115 2246 1116 2247
rect 1119 2247 1125 2248
rect 1119 2246 1120 2247
rect 1115 2244 1120 2246
rect 1115 2243 1116 2244
rect 1110 2242 1116 2243
rect 1119 2243 1120 2244
rect 1124 2243 1125 2247
rect 1190 2247 1191 2251
rect 1195 2247 1196 2251
rect 1190 2246 1196 2247
rect 1216 2246 1218 2256
rect 1326 2252 1332 2253
rect 1270 2251 1276 2252
rect 1223 2247 1229 2248
rect 1223 2246 1224 2247
rect 1216 2244 1224 2246
rect 1119 2242 1125 2243
rect 1223 2243 1224 2244
rect 1228 2243 1229 2247
rect 1270 2247 1271 2251
rect 1275 2247 1276 2251
rect 1326 2248 1327 2252
rect 1331 2248 1332 2252
rect 1270 2246 1276 2247
rect 1303 2247 1312 2248
rect 1326 2247 1332 2248
rect 1390 2251 1396 2252
rect 1390 2247 1391 2251
rect 1395 2250 1396 2251
rect 1710 2251 1716 2252
rect 1395 2248 1515 2250
rect 1395 2247 1396 2248
rect 1223 2242 1229 2243
rect 1303 2243 1304 2247
rect 1311 2243 1312 2247
rect 1390 2246 1396 2247
rect 1303 2242 1312 2243
rect 1366 2244 1372 2245
rect 1366 2240 1367 2244
rect 1371 2240 1372 2244
rect 1366 2239 1372 2240
rect 1398 2243 1404 2244
rect 1398 2239 1399 2243
rect 1403 2239 1404 2243
rect 1478 2243 1484 2244
rect 1398 2238 1404 2239
rect 1431 2239 1437 2240
rect 1278 2235 1284 2236
rect 1278 2231 1279 2235
rect 1283 2234 1284 2235
rect 1431 2235 1432 2239
rect 1436 2235 1437 2239
rect 1478 2239 1479 2243
rect 1483 2239 1484 2243
rect 1513 2240 1515 2248
rect 1710 2247 1711 2251
rect 1715 2250 1716 2251
rect 1715 2248 1866 2250
rect 1715 2247 1716 2248
rect 1710 2246 1716 2247
rect 1598 2243 1604 2244
rect 1478 2238 1484 2239
rect 1511 2239 1517 2240
rect 1431 2234 1437 2235
rect 1511 2235 1512 2239
rect 1516 2235 1517 2239
rect 1598 2239 1599 2243
rect 1603 2239 1604 2243
rect 1718 2243 1724 2244
rect 1598 2238 1604 2239
rect 1631 2239 1637 2240
rect 1631 2238 1632 2239
rect 1511 2234 1517 2235
rect 1608 2236 1632 2238
rect 1283 2232 1435 2234
rect 1283 2231 1284 2232
rect 1278 2230 1284 2231
rect 1486 2231 1492 2232
rect 1486 2227 1487 2231
rect 1491 2230 1492 2231
rect 1608 2230 1610 2236
rect 1631 2235 1632 2236
rect 1636 2235 1637 2239
rect 1718 2239 1719 2243
rect 1723 2239 1724 2243
rect 1838 2243 1844 2244
rect 1718 2238 1724 2239
rect 1750 2239 1757 2240
rect 1631 2234 1637 2235
rect 1750 2235 1751 2239
rect 1756 2235 1757 2239
rect 1838 2239 1839 2243
rect 1843 2239 1844 2243
rect 1838 2238 1844 2239
rect 1864 2238 1866 2248
rect 2582 2244 2588 2245
rect 1950 2243 1956 2244
rect 1871 2239 1877 2240
rect 1871 2238 1872 2239
rect 1864 2236 1872 2238
rect 1750 2234 1757 2235
rect 1871 2235 1872 2236
rect 1876 2235 1877 2239
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 2054 2243 2060 2244
rect 1950 2238 1956 2239
rect 1983 2239 1992 2240
rect 1871 2234 1877 2235
rect 1983 2235 1984 2239
rect 1991 2235 1992 2239
rect 2054 2239 2055 2243
rect 2059 2239 2060 2243
rect 2150 2243 2156 2244
rect 2054 2238 2060 2239
rect 2087 2239 2093 2240
rect 1983 2234 1992 2235
rect 2087 2235 2088 2239
rect 2092 2238 2093 2239
rect 2095 2239 2101 2240
rect 2095 2238 2096 2239
rect 2092 2236 2096 2238
rect 2092 2235 2093 2236
rect 2087 2234 2093 2235
rect 2095 2235 2096 2236
rect 2100 2235 2101 2239
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2238 2243 2244 2244
rect 2150 2238 2156 2239
rect 2183 2239 2192 2240
rect 2095 2234 2101 2235
rect 2183 2235 2184 2239
rect 2191 2235 2192 2239
rect 2238 2239 2239 2243
rect 2243 2239 2244 2243
rect 2318 2243 2324 2244
rect 2238 2238 2244 2239
rect 2271 2239 2280 2240
rect 2183 2234 2192 2235
rect 2271 2235 2272 2239
rect 2279 2235 2280 2239
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2390 2243 2396 2244
rect 2318 2238 2324 2239
rect 2351 2239 2357 2240
rect 2271 2234 2280 2235
rect 2351 2235 2352 2239
rect 2356 2238 2357 2239
rect 2390 2239 2391 2243
rect 2395 2239 2396 2243
rect 2470 2243 2476 2244
rect 2390 2238 2396 2239
rect 2422 2239 2429 2240
rect 2356 2236 2386 2238
rect 2356 2235 2357 2236
rect 2351 2234 2357 2235
rect 2384 2234 2386 2236
rect 2414 2235 2420 2236
rect 2414 2234 2415 2235
rect 2384 2232 2415 2234
rect 2414 2231 2415 2232
rect 2419 2231 2420 2235
rect 2422 2235 2423 2239
rect 2428 2235 2429 2239
rect 2470 2239 2471 2243
rect 2475 2239 2476 2243
rect 2526 2243 2532 2244
rect 2470 2238 2476 2239
rect 2503 2239 2512 2240
rect 2422 2234 2429 2235
rect 2503 2235 2504 2239
rect 2511 2235 2512 2239
rect 2526 2239 2527 2243
rect 2531 2239 2532 2243
rect 2582 2240 2583 2244
rect 2587 2240 2588 2244
rect 2526 2238 2532 2239
rect 2558 2239 2565 2240
rect 2582 2239 2588 2240
rect 2503 2234 2512 2235
rect 2558 2235 2559 2239
rect 2564 2235 2565 2239
rect 2558 2234 2565 2235
rect 2414 2230 2420 2231
rect 1491 2228 1610 2230
rect 1491 2227 1492 2228
rect 1486 2226 1492 2227
rect 1198 2219 1204 2220
rect 1198 2215 1199 2219
rect 1203 2218 1204 2219
rect 1203 2216 1298 2218
rect 1203 2215 1204 2216
rect 1198 2214 1204 2215
rect 175 2211 181 2212
rect 142 2209 148 2210
rect 110 2208 116 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 142 2205 143 2209
rect 147 2205 148 2209
rect 175 2207 176 2211
rect 180 2210 181 2211
rect 222 2211 228 2212
rect 222 2210 223 2211
rect 180 2208 223 2210
rect 180 2207 181 2208
rect 175 2206 181 2207
rect 222 2207 223 2208
rect 227 2207 228 2211
rect 263 2211 269 2212
rect 222 2206 228 2207
rect 230 2209 236 2210
rect 142 2204 148 2205
rect 230 2205 231 2209
rect 235 2205 236 2209
rect 263 2207 264 2211
rect 268 2210 269 2211
rect 350 2211 356 2212
rect 350 2210 351 2211
rect 268 2208 351 2210
rect 268 2207 269 2208
rect 263 2206 269 2207
rect 350 2207 351 2208
rect 355 2207 356 2211
rect 391 2211 397 2212
rect 350 2206 356 2207
rect 358 2209 364 2210
rect 230 2204 236 2205
rect 358 2205 359 2209
rect 363 2205 364 2209
rect 391 2207 392 2211
rect 396 2210 397 2211
rect 486 2211 492 2212
rect 486 2210 487 2211
rect 396 2208 487 2210
rect 396 2207 397 2208
rect 391 2206 397 2207
rect 486 2207 487 2208
rect 491 2207 492 2211
rect 527 2211 533 2212
rect 486 2206 492 2207
rect 494 2209 500 2210
rect 358 2204 364 2205
rect 494 2205 495 2209
rect 499 2205 500 2209
rect 527 2207 528 2211
rect 532 2210 533 2211
rect 614 2211 620 2212
rect 614 2210 615 2211
rect 532 2208 615 2210
rect 532 2207 533 2208
rect 527 2206 533 2207
rect 614 2207 615 2208
rect 619 2207 620 2211
rect 646 2211 652 2212
rect 614 2206 620 2207
rect 622 2209 628 2210
rect 494 2204 500 2205
rect 622 2205 623 2209
rect 627 2205 628 2209
rect 646 2207 647 2211
rect 651 2210 652 2211
rect 655 2211 661 2212
rect 655 2210 656 2211
rect 651 2208 656 2210
rect 651 2207 652 2208
rect 646 2206 652 2207
rect 655 2207 656 2208
rect 660 2207 661 2211
rect 783 2211 789 2212
rect 655 2206 661 2207
rect 750 2209 756 2210
rect 622 2204 628 2205
rect 750 2205 751 2209
rect 755 2205 756 2209
rect 783 2207 784 2211
rect 788 2210 789 2211
rect 862 2211 868 2212
rect 862 2210 863 2211
rect 788 2208 863 2210
rect 788 2207 789 2208
rect 783 2206 789 2207
rect 862 2207 863 2208
rect 867 2207 868 2211
rect 903 2211 909 2212
rect 862 2206 868 2207
rect 870 2209 876 2210
rect 750 2204 756 2205
rect 870 2205 871 2209
rect 875 2205 876 2209
rect 903 2207 904 2211
rect 908 2210 909 2211
rect 974 2211 980 2212
rect 974 2210 975 2211
rect 908 2208 975 2210
rect 908 2207 909 2208
rect 903 2206 909 2207
rect 974 2207 975 2208
rect 979 2207 980 2211
rect 1015 2211 1021 2212
rect 974 2206 980 2207
rect 982 2209 988 2210
rect 870 2204 876 2205
rect 982 2205 983 2209
rect 987 2205 988 2209
rect 1015 2207 1016 2211
rect 1020 2210 1021 2211
rect 1078 2211 1084 2212
rect 1078 2210 1079 2211
rect 1020 2208 1079 2210
rect 1020 2207 1021 2208
rect 1015 2206 1021 2207
rect 1078 2207 1079 2208
rect 1083 2207 1084 2211
rect 1119 2211 1125 2212
rect 1078 2206 1084 2207
rect 1086 2209 1092 2210
rect 982 2204 988 2205
rect 1086 2205 1087 2209
rect 1091 2205 1092 2209
rect 1119 2207 1120 2211
rect 1124 2210 1125 2211
rect 1182 2211 1188 2212
rect 1182 2210 1183 2211
rect 1124 2208 1183 2210
rect 1124 2207 1125 2208
rect 1119 2206 1125 2207
rect 1182 2207 1183 2208
rect 1187 2207 1188 2211
rect 1223 2211 1229 2212
rect 1182 2206 1188 2207
rect 1190 2209 1196 2210
rect 1086 2204 1092 2205
rect 1190 2205 1191 2209
rect 1195 2205 1196 2209
rect 1223 2207 1224 2211
rect 1228 2210 1229 2211
rect 1262 2211 1268 2212
rect 1262 2210 1263 2211
rect 1228 2208 1263 2210
rect 1228 2207 1229 2208
rect 1223 2206 1229 2207
rect 1262 2207 1263 2208
rect 1267 2207 1268 2211
rect 1296 2210 1298 2216
rect 1303 2211 1309 2212
rect 1303 2210 1304 2211
rect 1262 2206 1268 2207
rect 1270 2209 1276 2210
rect 1190 2204 1196 2205
rect 1270 2205 1271 2209
rect 1275 2205 1276 2209
rect 1296 2208 1304 2210
rect 1303 2207 1304 2208
rect 1308 2207 1309 2211
rect 1303 2206 1309 2207
rect 1326 2208 1332 2209
rect 1270 2204 1276 2205
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 110 2203 116 2204
rect 1326 2203 1332 2204
rect 2382 2203 2388 2204
rect 1487 2199 1493 2200
rect 1454 2197 1460 2198
rect 1366 2196 1372 2197
rect 1366 2192 1367 2196
rect 1371 2192 1372 2196
rect 1454 2193 1455 2197
rect 1459 2193 1460 2197
rect 1487 2195 1488 2199
rect 1492 2198 1493 2199
rect 1526 2199 1532 2200
rect 1526 2198 1527 2199
rect 1492 2196 1527 2198
rect 1492 2195 1493 2196
rect 1487 2194 1493 2195
rect 1526 2195 1527 2196
rect 1531 2195 1532 2199
rect 1567 2199 1573 2200
rect 1526 2194 1532 2195
rect 1534 2197 1540 2198
rect 1454 2192 1460 2193
rect 1534 2193 1535 2197
rect 1539 2193 1540 2197
rect 1567 2195 1568 2199
rect 1572 2198 1573 2199
rect 1622 2199 1628 2200
rect 1622 2198 1623 2199
rect 1572 2196 1623 2198
rect 1572 2195 1573 2196
rect 1567 2194 1573 2195
rect 1622 2195 1623 2196
rect 1627 2195 1628 2199
rect 1662 2199 1669 2200
rect 1622 2194 1628 2195
rect 1630 2197 1636 2198
rect 1534 2192 1540 2193
rect 1630 2193 1631 2197
rect 1635 2193 1636 2197
rect 1662 2195 1663 2199
rect 1668 2195 1669 2199
rect 1775 2199 1781 2200
rect 1662 2194 1669 2195
rect 1742 2197 1748 2198
rect 1630 2192 1636 2193
rect 1742 2193 1743 2197
rect 1747 2193 1748 2197
rect 1775 2195 1776 2199
rect 1780 2198 1781 2199
rect 1854 2199 1860 2200
rect 1854 2198 1855 2199
rect 1780 2196 1855 2198
rect 1780 2195 1781 2196
rect 1775 2194 1781 2195
rect 1854 2195 1855 2196
rect 1859 2195 1860 2199
rect 1895 2199 1901 2200
rect 1854 2194 1860 2195
rect 1862 2197 1868 2198
rect 1742 2192 1748 2193
rect 1862 2193 1863 2197
rect 1867 2193 1868 2197
rect 1895 2195 1896 2199
rect 1900 2198 1901 2199
rect 1974 2199 1980 2200
rect 1974 2198 1975 2199
rect 1900 2196 1975 2198
rect 1900 2195 1901 2196
rect 1895 2194 1901 2195
rect 1974 2195 1975 2196
rect 1979 2195 1980 2199
rect 2006 2199 2012 2200
rect 1974 2194 1980 2195
rect 1982 2197 1988 2198
rect 1862 2192 1868 2193
rect 1982 2193 1983 2197
rect 1987 2193 1988 2197
rect 2006 2195 2007 2199
rect 2011 2198 2012 2199
rect 2015 2199 2021 2200
rect 2015 2198 2016 2199
rect 2011 2196 2016 2198
rect 2011 2195 2012 2196
rect 2006 2194 2012 2195
rect 2015 2195 2016 2196
rect 2020 2195 2021 2199
rect 2127 2199 2133 2200
rect 2015 2194 2021 2195
rect 2094 2197 2100 2198
rect 1982 2192 1988 2193
rect 2094 2193 2095 2197
rect 2099 2193 2100 2197
rect 2127 2195 2128 2199
rect 2132 2198 2133 2199
rect 2198 2199 2204 2200
rect 2198 2198 2199 2199
rect 2132 2196 2199 2198
rect 2132 2195 2133 2196
rect 2127 2194 2133 2195
rect 2198 2195 2199 2196
rect 2203 2195 2204 2199
rect 2239 2199 2245 2200
rect 2198 2194 2204 2195
rect 2206 2197 2212 2198
rect 2094 2192 2100 2193
rect 2206 2193 2207 2197
rect 2211 2193 2212 2197
rect 2239 2195 2240 2199
rect 2244 2198 2245 2199
rect 2302 2199 2308 2200
rect 2302 2198 2303 2199
rect 2244 2196 2303 2198
rect 2244 2195 2245 2196
rect 2239 2194 2245 2195
rect 2302 2195 2303 2196
rect 2307 2195 2308 2199
rect 2338 2199 2349 2200
rect 2302 2194 2308 2195
rect 2310 2197 2316 2198
rect 2206 2192 2212 2193
rect 2310 2193 2311 2197
rect 2315 2193 2316 2197
rect 2338 2195 2339 2199
rect 2343 2195 2344 2199
rect 2348 2195 2349 2199
rect 2382 2199 2383 2203
rect 2387 2202 2388 2203
rect 2463 2203 2469 2204
rect 2387 2200 2450 2202
rect 2387 2199 2388 2200
rect 2382 2198 2388 2199
rect 2448 2198 2450 2200
rect 2455 2199 2461 2200
rect 2455 2198 2456 2199
rect 2338 2194 2349 2195
rect 2422 2197 2428 2198
rect 2310 2192 2316 2193
rect 2422 2193 2423 2197
rect 2427 2193 2428 2197
rect 2448 2196 2456 2198
rect 2455 2195 2456 2196
rect 2460 2195 2461 2199
rect 2463 2199 2464 2203
rect 2468 2202 2469 2203
rect 2468 2200 2554 2202
rect 2468 2199 2469 2200
rect 2463 2198 2469 2199
rect 2552 2198 2554 2200
rect 2559 2199 2565 2200
rect 2559 2198 2560 2199
rect 2455 2194 2461 2195
rect 2526 2197 2532 2198
rect 2422 2192 2428 2193
rect 2526 2193 2527 2197
rect 2531 2193 2532 2197
rect 2552 2196 2560 2198
rect 2559 2195 2560 2196
rect 2564 2195 2565 2199
rect 2559 2194 2565 2195
rect 2582 2196 2588 2197
rect 2526 2192 2532 2193
rect 2582 2192 2583 2196
rect 2587 2192 2588 2196
rect 110 2191 116 2192
rect 110 2187 111 2191
rect 115 2187 116 2191
rect 110 2186 116 2187
rect 1326 2191 1332 2192
rect 1366 2191 1372 2192
rect 2582 2191 2588 2192
rect 1326 2187 1327 2191
rect 1331 2187 1332 2191
rect 1326 2186 1332 2187
rect 158 2182 164 2183
rect 158 2178 159 2182
rect 163 2178 164 2182
rect 158 2177 164 2178
rect 246 2182 252 2183
rect 246 2178 247 2182
rect 251 2178 252 2182
rect 246 2177 252 2178
rect 374 2182 380 2183
rect 374 2178 375 2182
rect 379 2178 380 2182
rect 374 2177 380 2178
rect 510 2182 516 2183
rect 510 2178 511 2182
rect 515 2178 516 2182
rect 510 2177 516 2178
rect 638 2182 644 2183
rect 638 2178 639 2182
rect 643 2178 644 2182
rect 638 2177 644 2178
rect 766 2182 772 2183
rect 766 2178 767 2182
rect 771 2178 772 2182
rect 766 2177 772 2178
rect 886 2182 892 2183
rect 886 2178 887 2182
rect 891 2178 892 2182
rect 886 2177 892 2178
rect 998 2182 1004 2183
rect 998 2178 999 2182
rect 1003 2178 1004 2182
rect 998 2177 1004 2178
rect 1102 2182 1108 2183
rect 1102 2178 1103 2182
rect 1107 2178 1108 2182
rect 1102 2177 1108 2178
rect 1206 2182 1212 2183
rect 1206 2178 1207 2182
rect 1211 2178 1212 2182
rect 1206 2177 1212 2178
rect 1286 2182 1292 2183
rect 1286 2178 1287 2182
rect 1291 2178 1292 2182
rect 1286 2177 1292 2178
rect 1366 2179 1372 2180
rect 135 2175 141 2176
rect 135 2171 136 2175
rect 140 2174 141 2175
rect 166 2175 172 2176
rect 166 2174 167 2175
rect 140 2172 167 2174
rect 140 2171 141 2172
rect 135 2170 141 2171
rect 166 2171 167 2172
rect 171 2171 172 2175
rect 166 2170 172 2171
rect 222 2175 229 2176
rect 222 2171 223 2175
rect 228 2171 229 2175
rect 222 2170 229 2171
rect 350 2175 357 2176
rect 350 2171 351 2175
rect 356 2171 357 2175
rect 350 2170 357 2171
rect 486 2175 493 2176
rect 486 2171 487 2175
rect 492 2171 493 2175
rect 486 2170 493 2171
rect 614 2175 621 2176
rect 614 2171 615 2175
rect 620 2171 621 2175
rect 614 2170 621 2171
rect 743 2175 749 2176
rect 743 2171 744 2175
rect 748 2174 749 2175
rect 854 2175 860 2176
rect 854 2174 855 2175
rect 748 2172 855 2174
rect 748 2171 749 2172
rect 743 2170 749 2171
rect 854 2171 855 2172
rect 859 2171 860 2175
rect 854 2170 860 2171
rect 862 2175 869 2176
rect 862 2171 863 2175
rect 868 2171 869 2175
rect 862 2170 869 2171
rect 974 2175 981 2176
rect 974 2171 975 2175
rect 980 2171 981 2175
rect 974 2170 981 2171
rect 1078 2175 1085 2176
rect 1078 2171 1079 2175
rect 1084 2171 1085 2175
rect 1078 2170 1085 2171
rect 1182 2175 1189 2176
rect 1182 2171 1183 2175
rect 1188 2171 1189 2175
rect 1182 2170 1189 2171
rect 1262 2175 1269 2176
rect 1262 2171 1263 2175
rect 1268 2171 1269 2175
rect 1366 2175 1367 2179
rect 1371 2175 1372 2179
rect 1366 2174 1372 2175
rect 2582 2179 2588 2180
rect 2582 2175 2583 2179
rect 2587 2175 2588 2179
rect 2582 2174 2588 2175
rect 1262 2170 1269 2171
rect 1470 2170 1476 2171
rect 1470 2166 1471 2170
rect 1475 2166 1476 2170
rect 1470 2165 1476 2166
rect 1550 2170 1556 2171
rect 1550 2166 1551 2170
rect 1555 2166 1556 2170
rect 1550 2165 1556 2166
rect 1646 2170 1652 2171
rect 1646 2166 1647 2170
rect 1651 2166 1652 2170
rect 1646 2165 1652 2166
rect 1758 2170 1764 2171
rect 1758 2166 1759 2170
rect 1763 2166 1764 2170
rect 1758 2165 1764 2166
rect 1878 2170 1884 2171
rect 1878 2166 1879 2170
rect 1883 2166 1884 2170
rect 1878 2165 1884 2166
rect 1998 2170 2004 2171
rect 1998 2166 1999 2170
rect 2003 2166 2004 2170
rect 1998 2165 2004 2166
rect 2110 2170 2116 2171
rect 2110 2166 2111 2170
rect 2115 2166 2116 2170
rect 2110 2165 2116 2166
rect 2222 2170 2228 2171
rect 2222 2166 2223 2170
rect 2227 2166 2228 2170
rect 2222 2165 2228 2166
rect 2326 2170 2332 2171
rect 2326 2166 2327 2170
rect 2331 2166 2332 2170
rect 2326 2165 2332 2166
rect 2438 2170 2444 2171
rect 2438 2166 2439 2170
rect 2443 2166 2444 2170
rect 2438 2165 2444 2166
rect 2542 2170 2548 2171
rect 2542 2166 2543 2170
rect 2547 2166 2548 2170
rect 2542 2165 2548 2166
rect 1447 2163 1453 2164
rect 135 2159 144 2160
rect 135 2155 136 2159
rect 143 2155 144 2159
rect 178 2159 184 2160
rect 178 2155 179 2159
rect 183 2158 184 2159
rect 191 2159 197 2160
rect 191 2158 192 2159
rect 183 2156 192 2158
rect 183 2155 184 2156
rect 135 2154 144 2155
rect 158 2154 164 2155
rect 178 2154 184 2155
rect 191 2155 192 2156
rect 196 2155 197 2159
rect 234 2159 240 2160
rect 234 2155 235 2159
rect 239 2158 240 2159
rect 287 2159 293 2160
rect 287 2158 288 2159
rect 239 2156 288 2158
rect 239 2155 240 2156
rect 191 2154 197 2155
rect 214 2154 220 2155
rect 234 2154 240 2155
rect 287 2155 288 2156
rect 292 2155 293 2159
rect 330 2159 336 2160
rect 330 2155 331 2159
rect 335 2158 336 2159
rect 399 2159 405 2160
rect 399 2158 400 2159
rect 335 2156 400 2158
rect 335 2155 336 2156
rect 287 2154 293 2155
rect 310 2154 316 2155
rect 330 2154 336 2155
rect 399 2155 400 2156
rect 404 2155 405 2159
rect 479 2159 485 2160
rect 479 2155 480 2159
rect 484 2158 485 2159
rect 519 2159 525 2160
rect 519 2158 520 2159
rect 484 2156 520 2158
rect 484 2155 485 2156
rect 399 2154 405 2155
rect 422 2154 428 2155
rect 479 2154 485 2155
rect 519 2155 520 2156
rect 524 2155 525 2159
rect 562 2159 568 2160
rect 562 2155 563 2159
rect 567 2158 568 2159
rect 639 2159 645 2160
rect 639 2158 640 2159
rect 567 2156 640 2158
rect 567 2155 568 2156
rect 519 2154 525 2155
rect 542 2154 548 2155
rect 562 2154 568 2155
rect 639 2155 640 2156
rect 644 2155 645 2159
rect 750 2159 757 2160
rect 750 2155 751 2159
rect 756 2155 757 2159
rect 794 2159 800 2160
rect 794 2155 795 2159
rect 799 2158 800 2159
rect 855 2159 861 2160
rect 855 2158 856 2159
rect 799 2156 856 2158
rect 799 2155 800 2156
rect 639 2154 645 2155
rect 662 2154 668 2155
rect 750 2154 757 2155
rect 774 2154 780 2155
rect 794 2154 800 2155
rect 855 2155 856 2156
rect 860 2155 861 2159
rect 898 2159 904 2160
rect 898 2155 899 2159
rect 903 2158 904 2159
rect 951 2159 957 2160
rect 951 2158 952 2159
rect 903 2156 952 2158
rect 903 2155 904 2156
rect 855 2154 861 2155
rect 878 2154 884 2155
rect 898 2154 904 2155
rect 951 2155 952 2156
rect 956 2155 957 2159
rect 999 2159 1005 2160
rect 999 2155 1000 2159
rect 1004 2158 1005 2159
rect 1047 2159 1053 2160
rect 1047 2158 1048 2159
rect 1004 2156 1048 2158
rect 1004 2155 1005 2156
rect 951 2154 957 2155
rect 974 2154 980 2155
rect 999 2154 1005 2155
rect 1047 2155 1048 2156
rect 1052 2155 1053 2159
rect 1090 2159 1096 2160
rect 1090 2155 1091 2159
rect 1095 2158 1096 2159
rect 1143 2159 1149 2160
rect 1143 2158 1144 2159
rect 1095 2156 1144 2158
rect 1095 2155 1096 2156
rect 1047 2154 1053 2155
rect 1070 2154 1076 2155
rect 1090 2154 1096 2155
rect 1143 2155 1144 2156
rect 1148 2155 1149 2159
rect 1215 2159 1221 2160
rect 1215 2155 1216 2159
rect 1220 2158 1221 2159
rect 1247 2159 1253 2160
rect 1247 2158 1248 2159
rect 1220 2156 1248 2158
rect 1220 2155 1221 2156
rect 1143 2154 1149 2155
rect 1166 2154 1172 2155
rect 1215 2154 1221 2155
rect 1247 2155 1248 2156
rect 1252 2155 1253 2159
rect 1447 2159 1448 2163
rect 1452 2162 1453 2163
rect 1526 2163 1533 2164
rect 1452 2160 1522 2162
rect 1452 2159 1453 2160
rect 1447 2158 1453 2159
rect 1247 2154 1253 2155
rect 1270 2154 1276 2155
rect 158 2150 159 2154
rect 163 2150 164 2154
rect 158 2149 164 2150
rect 214 2150 215 2154
rect 219 2150 220 2154
rect 214 2149 220 2150
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 422 2150 423 2154
rect 427 2150 428 2154
rect 422 2149 428 2150
rect 542 2150 543 2154
rect 547 2150 548 2154
rect 542 2149 548 2150
rect 662 2150 663 2154
rect 667 2150 668 2154
rect 662 2149 668 2150
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 878 2150 879 2154
rect 883 2150 884 2154
rect 878 2149 884 2150
rect 974 2150 975 2154
rect 979 2150 980 2154
rect 974 2149 980 2150
rect 1070 2150 1071 2154
rect 1075 2150 1076 2154
rect 1070 2149 1076 2150
rect 1166 2150 1167 2154
rect 1171 2150 1172 2154
rect 1166 2149 1172 2150
rect 1270 2150 1271 2154
rect 1275 2150 1276 2154
rect 1520 2154 1522 2160
rect 1526 2159 1527 2163
rect 1532 2159 1533 2163
rect 1526 2158 1533 2159
rect 1622 2163 1629 2164
rect 1622 2159 1623 2163
rect 1628 2159 1629 2163
rect 1622 2158 1629 2159
rect 1735 2163 1741 2164
rect 1735 2159 1736 2163
rect 1740 2162 1741 2163
rect 1750 2163 1756 2164
rect 1750 2162 1751 2163
rect 1740 2160 1751 2162
rect 1740 2159 1741 2160
rect 1735 2158 1741 2159
rect 1750 2159 1751 2160
rect 1755 2159 1756 2163
rect 1750 2158 1756 2159
rect 1854 2163 1861 2164
rect 1854 2159 1855 2163
rect 1860 2159 1861 2163
rect 1854 2158 1861 2159
rect 1974 2163 1981 2164
rect 1974 2159 1975 2163
rect 1980 2159 1981 2163
rect 1974 2158 1981 2159
rect 2074 2163 2080 2164
rect 2074 2159 2075 2163
rect 2079 2162 2080 2163
rect 2087 2163 2093 2164
rect 2087 2162 2088 2163
rect 2079 2160 2088 2162
rect 2079 2159 2080 2160
rect 2074 2158 2080 2159
rect 2087 2159 2088 2160
rect 2092 2159 2093 2163
rect 2087 2158 2093 2159
rect 2198 2163 2205 2164
rect 2198 2159 2199 2163
rect 2204 2159 2205 2163
rect 2198 2158 2205 2159
rect 2302 2163 2309 2164
rect 2302 2159 2303 2163
rect 2308 2159 2309 2163
rect 2302 2158 2309 2159
rect 2415 2163 2421 2164
rect 2415 2159 2416 2163
rect 2420 2162 2421 2163
rect 2463 2163 2469 2164
rect 2463 2162 2464 2163
rect 2420 2160 2464 2162
rect 2420 2159 2421 2160
rect 2415 2158 2421 2159
rect 2463 2159 2464 2160
rect 2468 2159 2469 2163
rect 2463 2158 2469 2159
rect 2519 2163 2525 2164
rect 2519 2159 2520 2163
rect 2524 2162 2525 2163
rect 2558 2163 2564 2164
rect 2558 2162 2559 2163
rect 2524 2160 2559 2162
rect 2524 2159 2525 2160
rect 2519 2158 2525 2159
rect 2558 2159 2559 2160
rect 2563 2159 2564 2163
rect 2558 2158 2564 2159
rect 1542 2155 1548 2156
rect 1542 2154 1543 2155
rect 1520 2152 1543 2154
rect 1270 2149 1276 2150
rect 1510 2151 1517 2152
rect 1510 2147 1511 2151
rect 1516 2147 1517 2151
rect 1542 2151 1543 2152
rect 1547 2151 1548 2155
rect 2006 2155 2012 2156
rect 2006 2154 2007 2155
rect 1944 2152 2007 2154
rect 1542 2150 1548 2151
rect 1607 2151 1613 2152
rect 1607 2147 1608 2151
rect 1612 2150 1613 2151
rect 1622 2151 1628 2152
rect 1622 2150 1623 2151
rect 1612 2148 1623 2150
rect 1612 2147 1613 2148
rect 1510 2146 1517 2147
rect 1534 2146 1540 2147
rect 1607 2146 1613 2147
rect 1622 2147 1623 2148
rect 1627 2147 1628 2151
rect 1682 2151 1688 2152
rect 1682 2147 1683 2151
rect 1687 2150 1688 2151
rect 1711 2151 1717 2152
rect 1711 2150 1712 2151
rect 1687 2148 1712 2150
rect 1687 2147 1688 2148
rect 1622 2146 1628 2147
rect 1630 2146 1636 2147
rect 1682 2146 1688 2147
rect 1711 2147 1712 2148
rect 1716 2147 1717 2151
rect 1814 2151 1821 2152
rect 1814 2147 1815 2151
rect 1820 2147 1821 2151
rect 1927 2151 1933 2152
rect 1927 2147 1928 2151
rect 1932 2150 1933 2151
rect 1944 2150 1946 2152
rect 2006 2151 2007 2152
rect 2011 2151 2012 2155
rect 2294 2155 2300 2156
rect 2294 2154 2295 2155
rect 2256 2152 2295 2154
rect 2006 2150 2012 2151
rect 2031 2151 2037 2152
rect 1932 2148 1946 2150
rect 1932 2147 1933 2148
rect 2031 2147 2032 2151
rect 2036 2150 2037 2151
rect 2046 2151 2052 2152
rect 2046 2150 2047 2151
rect 2036 2148 2047 2150
rect 2036 2147 2037 2148
rect 1711 2146 1717 2147
rect 1734 2146 1740 2147
rect 1814 2146 1821 2147
rect 1838 2146 1844 2147
rect 1927 2146 1933 2147
rect 1950 2146 1956 2147
rect 2031 2146 2037 2147
rect 2046 2147 2047 2148
rect 2051 2147 2052 2151
rect 2134 2151 2141 2152
rect 2134 2147 2135 2151
rect 2140 2147 2141 2151
rect 2239 2151 2245 2152
rect 2239 2147 2240 2151
rect 2244 2150 2245 2151
rect 2256 2150 2258 2152
rect 2294 2151 2295 2152
rect 2299 2151 2300 2155
rect 2294 2150 2300 2151
rect 2335 2151 2344 2152
rect 2244 2148 2258 2150
rect 2244 2147 2245 2148
rect 2335 2147 2336 2151
rect 2343 2147 2344 2151
rect 2383 2151 2389 2152
rect 2383 2147 2384 2151
rect 2388 2150 2389 2151
rect 2439 2151 2445 2152
rect 2439 2150 2440 2151
rect 2388 2148 2440 2150
rect 2388 2147 2389 2148
rect 2046 2146 2052 2147
rect 2054 2146 2060 2147
rect 2134 2146 2141 2147
rect 2158 2146 2164 2147
rect 2239 2146 2245 2147
rect 2262 2146 2268 2147
rect 2335 2146 2344 2147
rect 2358 2146 2364 2147
rect 2383 2146 2389 2147
rect 2439 2147 2440 2148
rect 2444 2147 2445 2151
rect 2519 2151 2525 2152
rect 2519 2147 2520 2151
rect 2524 2150 2525 2151
rect 2534 2151 2540 2152
rect 2534 2150 2535 2151
rect 2524 2148 2535 2150
rect 2524 2147 2525 2148
rect 2439 2146 2445 2147
rect 2462 2146 2468 2147
rect 2519 2146 2525 2147
rect 2534 2147 2535 2148
rect 2539 2147 2540 2151
rect 2534 2146 2540 2147
rect 2542 2146 2548 2147
rect 110 2145 116 2146
rect 110 2141 111 2145
rect 115 2141 116 2145
rect 110 2140 116 2141
rect 1326 2145 1332 2146
rect 1326 2141 1327 2145
rect 1331 2141 1332 2145
rect 1534 2142 1535 2146
rect 1539 2142 1540 2146
rect 1534 2141 1540 2142
rect 1630 2142 1631 2146
rect 1635 2142 1636 2146
rect 1630 2141 1636 2142
rect 1734 2142 1735 2146
rect 1739 2142 1740 2146
rect 1734 2141 1740 2142
rect 1838 2142 1839 2146
rect 1843 2142 1844 2146
rect 1838 2141 1844 2142
rect 1950 2142 1951 2146
rect 1955 2142 1956 2146
rect 1950 2141 1956 2142
rect 2054 2142 2055 2146
rect 2059 2142 2060 2146
rect 2054 2141 2060 2142
rect 2158 2142 2159 2146
rect 2163 2142 2164 2146
rect 2158 2141 2164 2142
rect 2262 2142 2263 2146
rect 2267 2142 2268 2146
rect 2262 2141 2268 2142
rect 2358 2142 2359 2146
rect 2363 2142 2364 2146
rect 2358 2141 2364 2142
rect 2462 2142 2463 2146
rect 2467 2142 2468 2146
rect 2462 2141 2468 2142
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 1326 2140 1332 2141
rect 1366 2137 1372 2138
rect 1366 2133 1367 2137
rect 1371 2133 1372 2137
rect 1366 2132 1372 2133
rect 2582 2137 2588 2138
rect 2582 2133 2583 2137
rect 2587 2133 2588 2137
rect 2582 2132 2588 2133
rect 110 2128 116 2129
rect 1326 2128 1332 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 142 2127 148 2128
rect 142 2123 143 2127
rect 147 2123 148 2127
rect 198 2127 204 2128
rect 142 2122 148 2123
rect 175 2123 184 2124
rect 175 2119 176 2123
rect 183 2119 184 2123
rect 198 2123 199 2127
rect 203 2123 204 2127
rect 294 2127 300 2128
rect 198 2122 204 2123
rect 231 2123 240 2124
rect 175 2118 184 2119
rect 231 2119 232 2123
rect 239 2119 240 2123
rect 294 2123 295 2127
rect 299 2123 300 2127
rect 406 2127 412 2128
rect 294 2122 300 2123
rect 327 2123 336 2124
rect 231 2118 240 2119
rect 327 2119 328 2123
rect 335 2119 336 2123
rect 406 2123 407 2127
rect 411 2123 412 2127
rect 526 2127 532 2128
rect 406 2122 412 2123
rect 439 2123 445 2124
rect 327 2118 336 2119
rect 439 2119 440 2123
rect 444 2122 445 2123
rect 479 2123 485 2124
rect 479 2122 480 2123
rect 444 2120 480 2122
rect 444 2119 445 2120
rect 439 2118 445 2119
rect 479 2119 480 2120
rect 484 2119 485 2123
rect 526 2123 527 2127
rect 531 2123 532 2127
rect 646 2127 652 2128
rect 526 2122 532 2123
rect 559 2123 568 2124
rect 479 2118 485 2119
rect 559 2119 560 2123
rect 567 2119 568 2123
rect 646 2123 647 2127
rect 651 2123 652 2127
rect 758 2127 764 2128
rect 646 2122 652 2123
rect 670 2123 676 2124
rect 559 2118 568 2119
rect 670 2119 671 2123
rect 675 2122 676 2123
rect 679 2123 685 2124
rect 679 2122 680 2123
rect 675 2120 680 2122
rect 675 2119 676 2120
rect 670 2118 676 2119
rect 679 2119 680 2120
rect 684 2119 685 2123
rect 758 2123 759 2127
rect 763 2123 764 2127
rect 862 2127 868 2128
rect 758 2122 764 2123
rect 791 2123 800 2124
rect 679 2118 685 2119
rect 791 2119 792 2123
rect 799 2119 800 2123
rect 862 2123 863 2127
rect 867 2123 868 2127
rect 958 2127 964 2128
rect 862 2122 868 2123
rect 895 2123 904 2124
rect 791 2118 800 2119
rect 895 2119 896 2123
rect 903 2119 904 2123
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 1054 2127 1060 2128
rect 958 2122 964 2123
rect 991 2123 997 2124
rect 895 2118 904 2119
rect 991 2119 992 2123
rect 996 2122 997 2123
rect 999 2123 1005 2124
rect 999 2122 1000 2123
rect 996 2120 1000 2122
rect 996 2119 997 2120
rect 991 2118 997 2119
rect 999 2119 1000 2120
rect 1004 2119 1005 2123
rect 1054 2123 1055 2127
rect 1059 2123 1060 2127
rect 1150 2127 1156 2128
rect 1054 2122 1060 2123
rect 1087 2123 1096 2124
rect 999 2118 1005 2119
rect 1087 2119 1088 2123
rect 1095 2119 1096 2123
rect 1150 2123 1151 2127
rect 1155 2123 1156 2127
rect 1254 2127 1260 2128
rect 1150 2122 1156 2123
rect 1183 2123 1189 2124
rect 1087 2118 1096 2119
rect 1183 2119 1184 2123
rect 1188 2122 1189 2123
rect 1215 2123 1221 2124
rect 1215 2122 1216 2123
rect 1188 2120 1216 2122
rect 1188 2119 1189 2120
rect 1183 2118 1189 2119
rect 1215 2119 1216 2120
rect 1220 2119 1221 2123
rect 1254 2123 1255 2127
rect 1259 2123 1260 2127
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1254 2122 1260 2123
rect 1286 2123 1293 2124
rect 1326 2123 1332 2124
rect 1510 2127 1516 2128
rect 1510 2123 1511 2127
rect 1515 2126 1516 2127
rect 1814 2127 1820 2128
rect 1515 2124 1642 2126
rect 1515 2123 1516 2124
rect 1215 2118 1221 2119
rect 1286 2119 1287 2123
rect 1292 2119 1293 2123
rect 1510 2122 1516 2123
rect 1286 2118 1293 2119
rect 1366 2120 1372 2121
rect 1366 2116 1367 2120
rect 1371 2116 1372 2120
rect 1366 2115 1372 2116
rect 1518 2119 1524 2120
rect 1518 2115 1519 2119
rect 1523 2115 1524 2119
rect 1614 2119 1620 2120
rect 1518 2114 1524 2115
rect 1542 2115 1548 2116
rect 1542 2111 1543 2115
rect 1547 2114 1548 2115
rect 1551 2115 1557 2116
rect 1551 2114 1552 2115
rect 1547 2112 1552 2114
rect 1547 2111 1548 2112
rect 1542 2110 1548 2111
rect 1551 2111 1552 2112
rect 1556 2111 1557 2115
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1640 2114 1642 2124
rect 1814 2123 1815 2127
rect 1819 2126 1820 2127
rect 2134 2127 2140 2128
rect 1819 2124 1962 2126
rect 1819 2123 1820 2124
rect 1814 2122 1820 2123
rect 1718 2119 1724 2120
rect 1647 2115 1653 2116
rect 1647 2114 1648 2115
rect 1640 2112 1648 2114
rect 1551 2110 1557 2111
rect 1647 2111 1648 2112
rect 1652 2111 1653 2115
rect 1718 2115 1719 2119
rect 1723 2115 1724 2119
rect 1822 2119 1828 2120
rect 1718 2114 1724 2115
rect 1751 2115 1757 2116
rect 1751 2114 1752 2115
rect 1647 2110 1653 2111
rect 1728 2112 1752 2114
rect 1622 2107 1628 2108
rect 1622 2103 1623 2107
rect 1627 2106 1628 2107
rect 1728 2106 1730 2112
rect 1751 2111 1752 2112
rect 1756 2111 1757 2115
rect 1822 2115 1823 2119
rect 1827 2115 1828 2119
rect 1934 2119 1940 2120
rect 1822 2114 1828 2115
rect 1854 2115 1861 2116
rect 1751 2110 1757 2111
rect 1854 2111 1855 2115
rect 1860 2111 1861 2115
rect 1934 2115 1935 2119
rect 1939 2115 1940 2119
rect 1934 2114 1940 2115
rect 1960 2114 1962 2124
rect 2134 2123 2135 2127
rect 2139 2126 2140 2127
rect 2139 2124 2274 2126
rect 2139 2123 2140 2124
rect 2134 2122 2140 2123
rect 2038 2119 2044 2120
rect 1967 2115 1973 2116
rect 1967 2114 1968 2115
rect 1960 2112 1968 2114
rect 1854 2110 1861 2111
rect 1967 2111 1968 2112
rect 1972 2111 1973 2115
rect 2038 2115 2039 2119
rect 2043 2115 2044 2119
rect 2142 2119 2148 2120
rect 2038 2114 2044 2115
rect 2071 2115 2080 2116
rect 1967 2110 1973 2111
rect 2071 2111 2072 2115
rect 2079 2111 2080 2115
rect 2142 2115 2143 2119
rect 2147 2115 2148 2119
rect 2246 2119 2252 2120
rect 2142 2114 2148 2115
rect 2175 2115 2181 2116
rect 2175 2114 2176 2115
rect 2071 2110 2080 2111
rect 2152 2112 2176 2114
rect 1627 2104 1730 2106
rect 2046 2107 2052 2108
rect 1627 2103 1628 2104
rect 1622 2102 1628 2103
rect 2046 2103 2047 2107
rect 2051 2106 2052 2107
rect 2152 2106 2154 2112
rect 2175 2111 2176 2112
rect 2180 2111 2181 2115
rect 2246 2115 2247 2119
rect 2251 2115 2252 2119
rect 2246 2114 2252 2115
rect 2272 2114 2274 2124
rect 2582 2120 2588 2121
rect 2342 2119 2348 2120
rect 2279 2115 2285 2116
rect 2279 2114 2280 2115
rect 2272 2112 2280 2114
rect 2175 2110 2181 2111
rect 2279 2111 2280 2112
rect 2284 2111 2285 2115
rect 2342 2115 2343 2119
rect 2347 2115 2348 2119
rect 2446 2119 2452 2120
rect 2342 2114 2348 2115
rect 2375 2115 2381 2116
rect 2279 2110 2285 2111
rect 2375 2111 2376 2115
rect 2380 2114 2381 2115
rect 2383 2115 2389 2116
rect 2383 2114 2384 2115
rect 2380 2112 2384 2114
rect 2380 2111 2381 2112
rect 2375 2110 2381 2111
rect 2383 2111 2384 2112
rect 2388 2111 2389 2115
rect 2446 2115 2447 2119
rect 2451 2115 2452 2119
rect 2526 2119 2532 2120
rect 2446 2114 2452 2115
rect 2478 2115 2485 2116
rect 2383 2110 2389 2111
rect 2478 2111 2479 2115
rect 2484 2111 2485 2115
rect 2526 2115 2527 2119
rect 2531 2115 2532 2119
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2526 2114 2532 2115
rect 2558 2115 2565 2116
rect 2582 2115 2588 2116
rect 2478 2110 2485 2111
rect 2558 2111 2559 2115
rect 2564 2111 2565 2115
rect 2558 2110 2565 2111
rect 2051 2104 2154 2106
rect 2051 2103 2052 2104
rect 2046 2102 2052 2103
rect 750 2095 756 2096
rect 750 2091 751 2095
rect 755 2094 756 2095
rect 755 2092 1161 2094
rect 755 2091 756 2092
rect 750 2090 756 2091
rect 1159 2088 1161 2092
rect 1799 2091 1805 2092
rect 295 2087 301 2088
rect 262 2085 268 2086
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 262 2081 263 2085
rect 267 2081 268 2085
rect 295 2083 296 2087
rect 300 2086 301 2087
rect 318 2087 324 2088
rect 318 2086 319 2087
rect 300 2084 319 2086
rect 300 2083 301 2084
rect 295 2082 301 2083
rect 318 2083 319 2084
rect 323 2083 324 2087
rect 359 2087 365 2088
rect 318 2082 324 2083
rect 326 2085 332 2086
rect 262 2080 268 2081
rect 326 2081 327 2085
rect 331 2081 332 2085
rect 359 2083 360 2087
rect 364 2086 365 2087
rect 390 2087 396 2088
rect 390 2086 391 2087
rect 364 2084 391 2086
rect 364 2083 365 2084
rect 359 2082 365 2083
rect 390 2083 391 2084
rect 395 2083 396 2087
rect 431 2087 437 2088
rect 390 2082 396 2083
rect 398 2085 404 2086
rect 326 2080 332 2081
rect 398 2081 399 2085
rect 403 2081 404 2085
rect 431 2083 432 2087
rect 436 2086 437 2087
rect 470 2087 476 2088
rect 470 2086 471 2087
rect 436 2084 471 2086
rect 436 2083 437 2084
rect 431 2082 437 2083
rect 470 2083 471 2084
rect 475 2083 476 2087
rect 511 2087 517 2088
rect 470 2082 476 2083
rect 478 2085 484 2086
rect 398 2080 404 2081
rect 478 2081 479 2085
rect 483 2081 484 2085
rect 511 2083 512 2087
rect 516 2086 517 2087
rect 558 2087 564 2088
rect 558 2086 559 2087
rect 516 2084 559 2086
rect 516 2083 517 2084
rect 511 2082 517 2083
rect 558 2083 559 2084
rect 563 2083 564 2087
rect 599 2087 605 2088
rect 558 2082 564 2083
rect 566 2085 572 2086
rect 478 2080 484 2081
rect 566 2081 567 2085
rect 571 2081 572 2085
rect 599 2083 600 2087
rect 604 2086 605 2087
rect 646 2087 652 2088
rect 646 2086 647 2087
rect 604 2084 647 2086
rect 604 2083 605 2084
rect 599 2082 605 2083
rect 646 2083 647 2084
rect 651 2083 652 2087
rect 678 2087 684 2088
rect 646 2082 652 2083
rect 654 2085 660 2086
rect 566 2080 572 2081
rect 654 2081 655 2085
rect 659 2081 660 2085
rect 678 2083 679 2087
rect 683 2086 684 2087
rect 687 2087 693 2088
rect 687 2086 688 2087
rect 683 2084 688 2086
rect 683 2083 684 2084
rect 678 2082 684 2083
rect 687 2083 688 2084
rect 692 2083 693 2087
rect 767 2087 773 2088
rect 687 2082 693 2083
rect 734 2085 740 2086
rect 654 2080 660 2081
rect 734 2081 735 2085
rect 739 2081 740 2085
rect 767 2083 768 2087
rect 772 2086 773 2087
rect 806 2087 812 2088
rect 806 2086 807 2087
rect 772 2084 807 2086
rect 772 2083 773 2084
rect 767 2082 773 2083
rect 806 2083 807 2084
rect 811 2083 812 2087
rect 847 2087 853 2088
rect 806 2082 812 2083
rect 814 2085 820 2086
rect 734 2080 740 2081
rect 814 2081 815 2085
rect 819 2081 820 2085
rect 847 2083 848 2087
rect 852 2086 853 2087
rect 878 2087 884 2088
rect 878 2086 879 2087
rect 852 2084 879 2086
rect 852 2083 853 2084
rect 847 2082 853 2083
rect 878 2083 879 2084
rect 883 2083 884 2087
rect 919 2087 925 2088
rect 878 2082 884 2083
rect 886 2085 892 2086
rect 814 2080 820 2081
rect 886 2081 887 2085
rect 891 2081 892 2085
rect 919 2083 920 2087
rect 924 2086 925 2087
rect 958 2087 964 2088
rect 958 2086 959 2087
rect 924 2084 959 2086
rect 924 2083 925 2084
rect 919 2082 925 2083
rect 958 2083 959 2084
rect 963 2083 964 2087
rect 999 2087 1005 2088
rect 958 2082 964 2083
rect 966 2085 972 2086
rect 886 2080 892 2081
rect 966 2081 967 2085
rect 971 2081 972 2085
rect 999 2083 1000 2087
rect 1004 2086 1005 2087
rect 1038 2087 1044 2088
rect 1038 2086 1039 2087
rect 1004 2084 1039 2086
rect 1004 2083 1005 2084
rect 999 2082 1005 2083
rect 1038 2083 1039 2084
rect 1043 2083 1044 2087
rect 1079 2087 1085 2088
rect 1038 2082 1044 2083
rect 1046 2085 1052 2086
rect 966 2080 972 2081
rect 1046 2081 1047 2085
rect 1051 2081 1052 2085
rect 1079 2083 1080 2087
rect 1084 2086 1085 2087
rect 1118 2087 1124 2088
rect 1118 2086 1119 2087
rect 1084 2084 1119 2086
rect 1084 2083 1085 2084
rect 1079 2082 1085 2083
rect 1118 2083 1119 2084
rect 1123 2083 1124 2087
rect 1159 2087 1165 2088
rect 1118 2082 1124 2083
rect 1126 2085 1132 2086
rect 1046 2080 1052 2081
rect 1126 2081 1127 2085
rect 1131 2081 1132 2085
rect 1159 2083 1160 2087
rect 1164 2083 1165 2087
rect 1463 2087 1469 2088
rect 1430 2085 1436 2086
rect 1159 2082 1165 2083
rect 1326 2084 1332 2085
rect 1126 2080 1132 2081
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 110 2079 116 2080
rect 1326 2079 1332 2080
rect 1366 2084 1372 2085
rect 1366 2080 1367 2084
rect 1371 2080 1372 2084
rect 1430 2081 1431 2085
rect 1435 2081 1436 2085
rect 1463 2083 1464 2087
rect 1468 2086 1469 2087
rect 1526 2087 1532 2088
rect 1526 2086 1527 2087
rect 1468 2084 1527 2086
rect 1468 2083 1469 2084
rect 1463 2082 1469 2083
rect 1526 2083 1527 2084
rect 1531 2083 1532 2087
rect 1567 2087 1573 2088
rect 1526 2082 1532 2083
rect 1534 2085 1540 2086
rect 1430 2080 1436 2081
rect 1534 2081 1535 2085
rect 1539 2081 1540 2085
rect 1567 2083 1568 2087
rect 1572 2086 1573 2087
rect 1638 2087 1644 2088
rect 1638 2086 1639 2087
rect 1572 2084 1639 2086
rect 1572 2083 1573 2084
rect 1567 2082 1573 2083
rect 1638 2083 1639 2084
rect 1643 2083 1644 2087
rect 1679 2087 1688 2088
rect 1638 2082 1644 2083
rect 1646 2085 1652 2086
rect 1534 2080 1540 2081
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1679 2083 1680 2087
rect 1687 2083 1688 2087
rect 1786 2087 1797 2088
rect 1679 2082 1688 2083
rect 1758 2085 1764 2086
rect 1646 2080 1652 2081
rect 1758 2081 1759 2085
rect 1763 2081 1764 2085
rect 1786 2083 1787 2087
rect 1791 2083 1792 2087
rect 1796 2083 1797 2087
rect 1799 2087 1800 2091
rect 1804 2090 1805 2091
rect 2430 2091 2436 2092
rect 1804 2088 1890 2090
rect 1804 2087 1805 2088
rect 1799 2086 1805 2087
rect 1888 2086 1890 2088
rect 1895 2087 1901 2088
rect 1895 2086 1896 2087
rect 1786 2082 1797 2083
rect 1862 2085 1868 2086
rect 1758 2080 1764 2081
rect 1862 2081 1863 2085
rect 1867 2081 1868 2085
rect 1888 2084 1896 2086
rect 1895 2083 1896 2084
rect 1900 2083 1901 2087
rect 1999 2087 2005 2088
rect 1895 2082 1901 2083
rect 1966 2085 1972 2086
rect 1862 2080 1868 2081
rect 1966 2081 1967 2085
rect 1971 2081 1972 2085
rect 1999 2083 2000 2087
rect 2004 2086 2005 2087
rect 2062 2087 2068 2088
rect 2062 2086 2063 2087
rect 2004 2084 2063 2086
rect 2004 2083 2005 2084
rect 1999 2082 2005 2083
rect 2062 2083 2063 2084
rect 2067 2083 2068 2087
rect 2103 2087 2109 2088
rect 2062 2082 2068 2083
rect 2070 2085 2076 2086
rect 1966 2080 1972 2081
rect 2070 2081 2071 2085
rect 2075 2081 2076 2085
rect 2103 2083 2104 2087
rect 2108 2086 2109 2087
rect 2166 2087 2172 2088
rect 2166 2086 2167 2087
rect 2108 2084 2167 2086
rect 2108 2083 2109 2084
rect 2103 2082 2109 2083
rect 2166 2083 2167 2084
rect 2171 2083 2172 2087
rect 2207 2087 2213 2088
rect 2166 2082 2172 2083
rect 2174 2085 2180 2086
rect 2070 2080 2076 2081
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2207 2083 2208 2087
rect 2212 2086 2213 2087
rect 2262 2087 2268 2088
rect 2262 2086 2263 2087
rect 2212 2084 2263 2086
rect 2212 2083 2213 2084
rect 2207 2082 2213 2083
rect 2262 2083 2263 2084
rect 2267 2083 2268 2087
rect 2294 2087 2300 2088
rect 2262 2082 2268 2083
rect 2270 2085 2276 2086
rect 2174 2080 2180 2081
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2294 2083 2295 2087
rect 2299 2086 2300 2087
rect 2303 2087 2309 2088
rect 2303 2086 2304 2087
rect 2299 2084 2304 2086
rect 2299 2083 2300 2084
rect 2294 2082 2300 2083
rect 2303 2083 2304 2084
rect 2308 2083 2309 2087
rect 2391 2087 2397 2088
rect 2303 2082 2309 2083
rect 2358 2085 2364 2086
rect 2270 2080 2276 2081
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2391 2083 2392 2087
rect 2396 2086 2397 2087
rect 2422 2087 2428 2088
rect 2422 2086 2423 2087
rect 2396 2084 2423 2086
rect 2396 2083 2397 2084
rect 2391 2082 2397 2083
rect 2422 2083 2423 2084
rect 2427 2083 2428 2087
rect 2430 2087 2431 2091
rect 2435 2090 2436 2091
rect 2534 2091 2540 2092
rect 2435 2088 2482 2090
rect 2435 2087 2436 2088
rect 2430 2086 2436 2087
rect 2480 2086 2482 2088
rect 2487 2087 2493 2088
rect 2487 2086 2488 2087
rect 2422 2082 2428 2083
rect 2454 2085 2460 2086
rect 2358 2080 2364 2081
rect 2454 2081 2455 2085
rect 2459 2081 2460 2085
rect 2480 2084 2488 2086
rect 2487 2083 2488 2084
rect 2492 2083 2493 2087
rect 2534 2087 2535 2091
rect 2539 2090 2540 2091
rect 2539 2088 2554 2090
rect 2539 2087 2540 2088
rect 2534 2086 2540 2087
rect 2552 2086 2554 2088
rect 2559 2087 2565 2088
rect 2559 2086 2560 2087
rect 2487 2082 2493 2083
rect 2526 2085 2532 2086
rect 2454 2080 2460 2081
rect 2526 2081 2527 2085
rect 2531 2081 2532 2085
rect 2552 2084 2560 2086
rect 2559 2083 2560 2084
rect 2564 2083 2565 2087
rect 2559 2082 2565 2083
rect 2582 2084 2588 2085
rect 2526 2080 2532 2081
rect 2582 2080 2583 2084
rect 2587 2080 2588 2084
rect 1366 2079 1372 2080
rect 2582 2079 2588 2080
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 110 2062 116 2063
rect 1326 2067 1332 2068
rect 1326 2063 1327 2067
rect 1331 2063 1332 2067
rect 1326 2062 1332 2063
rect 1366 2067 1372 2068
rect 1366 2063 1367 2067
rect 1371 2063 1372 2067
rect 1366 2062 1372 2063
rect 2582 2067 2588 2068
rect 2582 2063 2583 2067
rect 2587 2063 2588 2067
rect 2582 2062 2588 2063
rect 278 2058 284 2059
rect 278 2054 279 2058
rect 283 2054 284 2058
rect 278 2053 284 2054
rect 342 2058 348 2059
rect 342 2054 343 2058
rect 347 2054 348 2058
rect 342 2053 348 2054
rect 414 2058 420 2059
rect 414 2054 415 2058
rect 419 2054 420 2058
rect 414 2053 420 2054
rect 494 2058 500 2059
rect 494 2054 495 2058
rect 499 2054 500 2058
rect 494 2053 500 2054
rect 582 2058 588 2059
rect 582 2054 583 2058
rect 587 2054 588 2058
rect 582 2053 588 2054
rect 670 2058 676 2059
rect 670 2054 671 2058
rect 675 2054 676 2058
rect 670 2053 676 2054
rect 750 2058 756 2059
rect 750 2054 751 2058
rect 755 2054 756 2058
rect 750 2053 756 2054
rect 830 2058 836 2059
rect 830 2054 831 2058
rect 835 2054 836 2058
rect 830 2053 836 2054
rect 902 2058 908 2059
rect 902 2054 903 2058
rect 907 2054 908 2058
rect 902 2053 908 2054
rect 982 2058 988 2059
rect 982 2054 983 2058
rect 987 2054 988 2058
rect 982 2053 988 2054
rect 1062 2058 1068 2059
rect 1062 2054 1063 2058
rect 1067 2054 1068 2058
rect 1062 2053 1068 2054
rect 1142 2058 1148 2059
rect 1142 2054 1143 2058
rect 1147 2054 1148 2058
rect 1142 2053 1148 2054
rect 1446 2058 1452 2059
rect 1446 2054 1447 2058
rect 1451 2054 1452 2058
rect 1446 2053 1452 2054
rect 1550 2058 1556 2059
rect 1550 2054 1551 2058
rect 1555 2054 1556 2058
rect 1550 2053 1556 2054
rect 1662 2058 1668 2059
rect 1662 2054 1663 2058
rect 1667 2054 1668 2058
rect 1662 2053 1668 2054
rect 1774 2058 1780 2059
rect 1774 2054 1775 2058
rect 1779 2054 1780 2058
rect 1774 2053 1780 2054
rect 1878 2058 1884 2059
rect 1878 2054 1879 2058
rect 1883 2054 1884 2058
rect 1878 2053 1884 2054
rect 1982 2058 1988 2059
rect 1982 2054 1983 2058
rect 1987 2054 1988 2058
rect 1982 2053 1988 2054
rect 2086 2058 2092 2059
rect 2086 2054 2087 2058
rect 2091 2054 2092 2058
rect 2086 2053 2092 2054
rect 2190 2058 2196 2059
rect 2190 2054 2191 2058
rect 2195 2054 2196 2058
rect 2190 2053 2196 2054
rect 2286 2058 2292 2059
rect 2286 2054 2287 2058
rect 2291 2054 2292 2058
rect 2286 2053 2292 2054
rect 2374 2058 2380 2059
rect 2374 2054 2375 2058
rect 2379 2054 2380 2058
rect 2374 2053 2380 2054
rect 2470 2058 2476 2059
rect 2470 2054 2471 2058
rect 2475 2054 2476 2058
rect 2470 2053 2476 2054
rect 2542 2058 2548 2059
rect 2542 2054 2543 2058
rect 2547 2054 2548 2058
rect 2542 2053 2548 2054
rect 255 2051 264 2052
rect 255 2047 256 2051
rect 263 2047 264 2051
rect 255 2046 264 2047
rect 318 2051 325 2052
rect 318 2047 319 2051
rect 324 2047 325 2051
rect 318 2046 325 2047
rect 390 2051 397 2052
rect 390 2047 391 2051
rect 396 2047 397 2051
rect 390 2046 397 2047
rect 470 2051 477 2052
rect 470 2047 471 2051
rect 476 2047 477 2051
rect 470 2046 477 2047
rect 558 2051 565 2052
rect 558 2047 559 2051
rect 564 2047 565 2051
rect 558 2046 565 2047
rect 646 2051 653 2052
rect 646 2047 647 2051
rect 652 2047 653 2051
rect 646 2046 653 2047
rect 727 2051 733 2052
rect 727 2047 728 2051
rect 732 2050 733 2051
rect 806 2051 813 2052
rect 732 2048 802 2050
rect 732 2047 733 2048
rect 727 2046 733 2047
rect 800 2042 802 2048
rect 806 2047 807 2051
rect 812 2047 813 2051
rect 806 2046 813 2047
rect 878 2051 885 2052
rect 878 2047 879 2051
rect 884 2047 885 2051
rect 878 2046 885 2047
rect 958 2051 965 2052
rect 958 2047 959 2051
rect 964 2047 965 2051
rect 958 2046 965 2047
rect 1038 2051 1045 2052
rect 1038 2047 1039 2051
rect 1044 2047 1045 2051
rect 1038 2046 1045 2047
rect 1118 2051 1125 2052
rect 1118 2047 1119 2051
rect 1124 2047 1125 2051
rect 1118 2046 1125 2047
rect 1423 2051 1432 2052
rect 1423 2047 1424 2051
rect 1431 2047 1432 2051
rect 1423 2046 1432 2047
rect 1526 2051 1533 2052
rect 1526 2047 1527 2051
rect 1532 2047 1533 2051
rect 1526 2046 1533 2047
rect 1638 2051 1645 2052
rect 1638 2047 1639 2051
rect 1644 2047 1645 2051
rect 1638 2046 1645 2047
rect 1751 2051 1757 2052
rect 1751 2047 1752 2051
rect 1756 2050 1757 2051
rect 1799 2051 1805 2052
rect 1799 2050 1800 2051
rect 1756 2048 1800 2050
rect 1756 2047 1757 2048
rect 1751 2046 1757 2047
rect 1799 2047 1800 2048
rect 1804 2047 1805 2051
rect 1799 2046 1805 2047
rect 1854 2051 1861 2052
rect 1854 2047 1855 2051
rect 1860 2047 1861 2051
rect 1854 2046 1861 2047
rect 1959 2051 1965 2052
rect 1959 2047 1960 2051
rect 1964 2050 1965 2051
rect 2054 2051 2060 2052
rect 2054 2050 2055 2051
rect 1964 2048 2055 2050
rect 1964 2047 1965 2048
rect 1959 2046 1965 2047
rect 2054 2047 2055 2048
rect 2059 2047 2060 2051
rect 2054 2046 2060 2047
rect 2062 2051 2069 2052
rect 2062 2047 2063 2051
rect 2068 2047 2069 2051
rect 2062 2046 2069 2047
rect 2166 2051 2173 2052
rect 2166 2047 2167 2051
rect 2172 2047 2173 2051
rect 2166 2046 2173 2047
rect 2262 2051 2269 2052
rect 2262 2047 2263 2051
rect 2268 2047 2269 2051
rect 2262 2046 2269 2047
rect 2351 2051 2357 2052
rect 2351 2047 2352 2051
rect 2356 2050 2357 2051
rect 2430 2051 2436 2052
rect 2430 2050 2431 2051
rect 2356 2048 2431 2050
rect 2356 2047 2357 2048
rect 2351 2046 2357 2047
rect 2430 2047 2431 2048
rect 2435 2047 2436 2051
rect 2430 2046 2436 2047
rect 2447 2051 2453 2052
rect 2447 2047 2448 2051
rect 2452 2050 2453 2051
rect 2478 2051 2484 2052
rect 2478 2050 2479 2051
rect 2452 2048 2479 2050
rect 2452 2047 2453 2048
rect 2447 2046 2453 2047
rect 2478 2047 2479 2048
rect 2483 2047 2484 2051
rect 2478 2046 2484 2047
rect 2519 2051 2525 2052
rect 2519 2047 2520 2051
rect 2524 2050 2525 2051
rect 2558 2051 2564 2052
rect 2558 2050 2559 2051
rect 2524 2048 2559 2050
rect 2524 2047 2525 2048
rect 2519 2046 2525 2047
rect 2558 2047 2559 2048
rect 2563 2047 2564 2051
rect 2558 2046 2564 2047
rect 1046 2043 1052 2044
rect 1046 2042 1047 2043
rect 800 2040 1047 2042
rect 678 2039 684 2040
rect 678 2038 679 2039
rect 408 2036 679 2038
rect 391 2031 397 2032
rect 391 2027 392 2031
rect 396 2030 397 2031
rect 408 2030 410 2036
rect 678 2035 679 2036
rect 683 2035 684 2039
rect 1046 2039 1047 2040
rect 1051 2039 1052 2043
rect 1046 2038 1052 2039
rect 1390 2039 1397 2040
rect 678 2034 684 2035
rect 1390 2035 1391 2039
rect 1396 2035 1397 2039
rect 1479 2039 1485 2040
rect 1479 2035 1480 2039
rect 1484 2038 1485 2039
rect 1494 2039 1500 2040
rect 1494 2038 1495 2039
rect 1484 2036 1495 2038
rect 1484 2035 1485 2036
rect 1390 2034 1397 2035
rect 1414 2034 1420 2035
rect 1479 2034 1485 2035
rect 1494 2035 1495 2036
rect 1499 2035 1500 2039
rect 1522 2039 1528 2040
rect 1522 2035 1523 2039
rect 1527 2038 1528 2039
rect 1583 2039 1589 2040
rect 1583 2038 1584 2039
rect 1527 2036 1584 2038
rect 1527 2035 1528 2036
rect 1494 2034 1500 2035
rect 1502 2034 1508 2035
rect 1522 2034 1528 2035
rect 1583 2035 1584 2036
rect 1588 2035 1589 2039
rect 1686 2039 1693 2040
rect 1686 2035 1687 2039
rect 1692 2035 1693 2039
rect 1783 2039 1792 2040
rect 1783 2035 1784 2039
rect 1791 2035 1792 2039
rect 1879 2039 1885 2040
rect 1879 2035 1880 2039
rect 1884 2038 1885 2039
rect 1894 2039 1900 2040
rect 1894 2038 1895 2039
rect 1884 2036 1895 2038
rect 1884 2035 1885 2036
rect 1583 2034 1589 2035
rect 1606 2034 1612 2035
rect 1686 2034 1693 2035
rect 1710 2034 1716 2035
rect 1783 2034 1792 2035
rect 1806 2034 1812 2035
rect 1879 2034 1885 2035
rect 1894 2035 1895 2036
rect 1899 2035 1900 2039
rect 1918 2039 1924 2040
rect 1918 2035 1919 2039
rect 1923 2038 1924 2039
rect 1983 2039 1989 2040
rect 1983 2038 1984 2039
rect 1923 2036 1984 2038
rect 1923 2035 1924 2036
rect 1894 2034 1900 2035
rect 1902 2034 1908 2035
rect 1918 2034 1924 2035
rect 1983 2035 1984 2036
rect 1988 2035 1989 2039
rect 2031 2039 2037 2040
rect 2031 2035 2032 2039
rect 2036 2038 2037 2039
rect 2087 2039 2093 2040
rect 2087 2038 2088 2039
rect 2036 2036 2088 2038
rect 2036 2035 2037 2036
rect 1983 2034 1989 2035
rect 2006 2034 2012 2035
rect 2031 2034 2037 2035
rect 2087 2035 2088 2036
rect 2092 2035 2093 2039
rect 2130 2039 2136 2040
rect 2130 2035 2131 2039
rect 2135 2038 2136 2039
rect 2191 2039 2197 2040
rect 2191 2038 2192 2039
rect 2135 2036 2192 2038
rect 2135 2035 2136 2036
rect 2087 2034 2093 2035
rect 2110 2034 2116 2035
rect 2130 2034 2136 2035
rect 2191 2035 2192 2036
rect 2196 2035 2197 2039
rect 2234 2039 2240 2040
rect 2234 2035 2235 2039
rect 2239 2038 2240 2039
rect 2303 2039 2309 2040
rect 2303 2038 2304 2039
rect 2239 2036 2304 2038
rect 2239 2035 2240 2036
rect 2191 2034 2197 2035
rect 2214 2034 2220 2035
rect 2234 2034 2240 2035
rect 2303 2035 2304 2036
rect 2308 2035 2309 2039
rect 2422 2039 2429 2040
rect 2422 2035 2423 2039
rect 2428 2035 2429 2039
rect 2471 2039 2477 2040
rect 2471 2035 2472 2039
rect 2476 2038 2477 2039
rect 2519 2039 2525 2040
rect 2519 2038 2520 2039
rect 2476 2036 2520 2038
rect 2476 2035 2477 2036
rect 2303 2034 2309 2035
rect 2326 2034 2332 2035
rect 2422 2034 2429 2035
rect 2446 2034 2452 2035
rect 2471 2034 2477 2035
rect 2519 2035 2520 2036
rect 2524 2035 2525 2039
rect 2519 2034 2525 2035
rect 2542 2034 2548 2035
rect 396 2028 410 2030
rect 439 2031 445 2032
rect 396 2027 397 2028
rect 439 2027 440 2031
rect 444 2030 445 2031
rect 447 2031 453 2032
rect 447 2030 448 2031
rect 444 2028 448 2030
rect 444 2027 445 2028
rect 391 2026 397 2027
rect 414 2026 420 2027
rect 439 2026 445 2027
rect 447 2027 448 2028
rect 452 2027 453 2031
rect 495 2031 501 2032
rect 495 2027 496 2031
rect 500 2030 501 2031
rect 503 2031 509 2032
rect 503 2030 504 2031
rect 500 2028 504 2030
rect 500 2027 501 2028
rect 447 2026 453 2027
rect 470 2026 476 2027
rect 495 2026 501 2027
rect 503 2027 504 2028
rect 508 2027 509 2031
rect 546 2031 552 2032
rect 546 2027 547 2031
rect 551 2030 552 2031
rect 559 2031 565 2032
rect 559 2030 560 2031
rect 551 2028 560 2030
rect 551 2027 552 2028
rect 503 2026 509 2027
rect 526 2026 532 2027
rect 546 2026 552 2027
rect 559 2027 560 2028
rect 564 2027 565 2031
rect 602 2031 608 2032
rect 602 2027 603 2031
rect 607 2030 608 2031
rect 615 2031 621 2032
rect 615 2030 616 2031
rect 607 2028 616 2030
rect 607 2027 608 2028
rect 559 2026 565 2027
rect 582 2026 588 2027
rect 602 2026 608 2027
rect 615 2027 616 2028
rect 620 2027 621 2031
rect 658 2031 664 2032
rect 658 2027 659 2031
rect 663 2030 664 2031
rect 671 2031 677 2032
rect 671 2030 672 2031
rect 663 2028 672 2030
rect 663 2027 664 2028
rect 615 2026 621 2027
rect 638 2026 644 2027
rect 658 2026 664 2027
rect 671 2027 672 2028
rect 676 2027 677 2031
rect 727 2031 733 2032
rect 727 2027 728 2031
rect 732 2030 733 2031
rect 742 2031 748 2032
rect 742 2030 743 2031
rect 732 2028 743 2030
rect 732 2027 733 2028
rect 671 2026 677 2027
rect 694 2026 700 2027
rect 727 2026 733 2027
rect 742 2027 743 2028
rect 747 2027 748 2031
rect 775 2031 781 2032
rect 775 2027 776 2031
rect 780 2030 781 2031
rect 783 2031 789 2032
rect 783 2030 784 2031
rect 780 2028 784 2030
rect 780 2027 781 2028
rect 742 2026 748 2027
rect 750 2026 756 2027
rect 775 2026 781 2027
rect 783 2027 784 2028
rect 788 2027 789 2031
rect 831 2031 837 2032
rect 831 2027 832 2031
rect 836 2030 837 2031
rect 839 2031 845 2032
rect 839 2030 840 2031
rect 836 2028 840 2030
rect 836 2027 837 2028
rect 783 2026 789 2027
rect 806 2026 812 2027
rect 831 2026 837 2027
rect 839 2027 840 2028
rect 844 2027 845 2031
rect 887 2031 893 2032
rect 887 2027 888 2031
rect 892 2030 893 2031
rect 895 2031 901 2032
rect 895 2030 896 2031
rect 892 2028 896 2030
rect 892 2027 893 2028
rect 839 2026 845 2027
rect 862 2026 868 2027
rect 887 2026 893 2027
rect 895 2027 896 2028
rect 900 2027 901 2031
rect 943 2031 949 2032
rect 943 2027 944 2031
rect 948 2030 949 2031
rect 951 2031 957 2032
rect 951 2030 952 2031
rect 948 2028 952 2030
rect 948 2027 949 2028
rect 895 2026 901 2027
rect 918 2026 924 2027
rect 943 2026 949 2027
rect 951 2027 952 2028
rect 956 2027 957 2031
rect 999 2031 1005 2032
rect 999 2027 1000 2031
rect 1004 2030 1005 2031
rect 1007 2031 1013 2032
rect 1007 2030 1008 2031
rect 1004 2028 1008 2030
rect 1004 2027 1005 2028
rect 951 2026 957 2027
rect 974 2026 980 2027
rect 999 2026 1005 2027
rect 1007 2027 1008 2028
rect 1012 2027 1013 2031
rect 1414 2030 1415 2034
rect 1419 2030 1420 2034
rect 1414 2029 1420 2030
rect 1502 2030 1503 2034
rect 1507 2030 1508 2034
rect 1502 2029 1508 2030
rect 1606 2030 1607 2034
rect 1611 2030 1612 2034
rect 1606 2029 1612 2030
rect 1710 2030 1711 2034
rect 1715 2030 1716 2034
rect 1710 2029 1716 2030
rect 1806 2030 1807 2034
rect 1811 2030 1812 2034
rect 1806 2029 1812 2030
rect 1902 2030 1903 2034
rect 1907 2030 1908 2034
rect 1902 2029 1908 2030
rect 2006 2030 2007 2034
rect 2011 2030 2012 2034
rect 2006 2029 2012 2030
rect 2110 2030 2111 2034
rect 2115 2030 2116 2034
rect 2110 2029 2116 2030
rect 2214 2030 2215 2034
rect 2219 2030 2220 2034
rect 2214 2029 2220 2030
rect 2326 2030 2327 2034
rect 2331 2030 2332 2034
rect 2326 2029 2332 2030
rect 2446 2030 2447 2034
rect 2451 2030 2452 2034
rect 2446 2029 2452 2030
rect 2542 2030 2543 2034
rect 2547 2030 2548 2034
rect 2542 2029 2548 2030
rect 1007 2026 1013 2027
rect 1030 2026 1036 2027
rect 414 2022 415 2026
rect 419 2022 420 2026
rect 414 2021 420 2022
rect 470 2022 471 2026
rect 475 2022 476 2026
rect 470 2021 476 2022
rect 526 2022 527 2026
rect 531 2022 532 2026
rect 526 2021 532 2022
rect 582 2022 583 2026
rect 587 2022 588 2026
rect 582 2021 588 2022
rect 638 2022 639 2026
rect 643 2022 644 2026
rect 638 2021 644 2022
rect 694 2022 695 2026
rect 699 2022 700 2026
rect 694 2021 700 2022
rect 750 2022 751 2026
rect 755 2022 756 2026
rect 750 2021 756 2022
rect 806 2022 807 2026
rect 811 2022 812 2026
rect 806 2021 812 2022
rect 862 2022 863 2026
rect 867 2022 868 2026
rect 862 2021 868 2022
rect 918 2022 919 2026
rect 923 2022 924 2026
rect 918 2021 924 2022
rect 974 2022 975 2026
rect 979 2022 980 2026
rect 974 2021 980 2022
rect 1030 2022 1031 2026
rect 1035 2022 1036 2026
rect 1030 2021 1036 2022
rect 1366 2025 1372 2026
rect 1366 2021 1367 2025
rect 1371 2021 1372 2025
rect 1366 2020 1372 2021
rect 2582 2025 2588 2026
rect 2582 2021 2583 2025
rect 2587 2021 2588 2025
rect 2582 2020 2588 2021
rect 110 2017 116 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 1326 2017 1332 2018
rect 1326 2013 1327 2017
rect 1331 2013 1332 2017
rect 1326 2012 1332 2013
rect 1390 2015 1396 2016
rect 1390 2011 1391 2015
rect 1395 2014 1396 2015
rect 1686 2015 1692 2016
rect 1395 2012 1618 2014
rect 1395 2011 1396 2012
rect 1390 2010 1396 2011
rect 1366 2008 1372 2009
rect 1366 2004 1367 2008
rect 1371 2004 1372 2008
rect 1366 2003 1372 2004
rect 1398 2007 1404 2008
rect 1398 2003 1399 2007
rect 1403 2003 1404 2007
rect 1486 2007 1492 2008
rect 1398 2002 1404 2003
rect 1426 2003 1437 2004
rect 110 2000 116 2001
rect 1326 2000 1332 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 398 1999 404 2000
rect 398 1995 399 1999
rect 403 1995 404 1999
rect 454 1999 460 2000
rect 398 1994 404 1995
rect 431 1995 437 1996
rect 431 1991 432 1995
rect 436 1994 437 1995
rect 439 1995 445 1996
rect 439 1994 440 1995
rect 436 1992 440 1994
rect 436 1991 437 1992
rect 431 1990 437 1991
rect 439 1991 440 1992
rect 444 1991 445 1995
rect 454 1995 455 1999
rect 459 1995 460 1999
rect 510 1999 516 2000
rect 454 1994 460 1995
rect 487 1995 493 1996
rect 439 1990 445 1991
rect 487 1991 488 1995
rect 492 1994 493 1995
rect 495 1995 501 1996
rect 495 1994 496 1995
rect 492 1992 496 1994
rect 492 1991 493 1992
rect 487 1990 493 1991
rect 495 1991 496 1992
rect 500 1991 501 1995
rect 510 1995 511 1999
rect 515 1995 516 1999
rect 566 1999 572 2000
rect 510 1994 516 1995
rect 543 1995 552 1996
rect 495 1990 501 1991
rect 543 1991 544 1995
rect 551 1991 552 1995
rect 566 1995 567 1999
rect 571 1995 572 1999
rect 622 1999 628 2000
rect 566 1994 572 1995
rect 599 1995 608 1996
rect 543 1990 552 1991
rect 599 1991 600 1995
rect 607 1991 608 1995
rect 622 1995 623 1999
rect 627 1995 628 1999
rect 678 1999 684 2000
rect 622 1994 628 1995
rect 655 1995 664 1996
rect 599 1990 608 1991
rect 655 1991 656 1995
rect 663 1991 664 1995
rect 678 1995 679 1999
rect 683 1995 684 1999
rect 734 1999 740 2000
rect 678 1994 684 1995
rect 711 1995 717 1996
rect 711 1994 712 1995
rect 655 1990 664 1991
rect 696 1992 712 1994
rect 590 1987 596 1988
rect 590 1983 591 1987
rect 595 1986 596 1987
rect 696 1986 698 1992
rect 711 1991 712 1992
rect 716 1991 717 1995
rect 734 1995 735 1999
rect 739 1995 740 1999
rect 790 1999 796 2000
rect 734 1994 740 1995
rect 767 1995 773 1996
rect 711 1990 717 1991
rect 767 1991 768 1995
rect 772 1994 773 1995
rect 775 1995 781 1996
rect 775 1994 776 1995
rect 772 1992 776 1994
rect 772 1991 773 1992
rect 767 1990 773 1991
rect 775 1991 776 1992
rect 780 1991 781 1995
rect 790 1995 791 1999
rect 795 1995 796 1999
rect 846 1999 852 2000
rect 790 1994 796 1995
rect 823 1995 829 1996
rect 775 1990 781 1991
rect 823 1991 824 1995
rect 828 1994 829 1995
rect 831 1995 837 1996
rect 831 1994 832 1995
rect 828 1992 832 1994
rect 828 1991 829 1992
rect 823 1990 829 1991
rect 831 1991 832 1992
rect 836 1991 837 1995
rect 846 1995 847 1999
rect 851 1995 852 1999
rect 902 1999 908 2000
rect 846 1994 852 1995
rect 879 1995 885 1996
rect 831 1990 837 1991
rect 879 1991 880 1995
rect 884 1994 885 1995
rect 887 1995 893 1996
rect 887 1994 888 1995
rect 884 1992 888 1994
rect 884 1991 885 1992
rect 879 1990 885 1991
rect 887 1991 888 1992
rect 892 1991 893 1995
rect 902 1995 903 1999
rect 907 1995 908 1999
rect 958 1999 964 2000
rect 902 1994 908 1995
rect 935 1995 941 1996
rect 887 1990 893 1991
rect 935 1991 936 1995
rect 940 1994 941 1995
rect 943 1995 949 1996
rect 943 1994 944 1995
rect 940 1992 944 1994
rect 940 1991 941 1992
rect 935 1990 941 1991
rect 943 1991 944 1992
rect 948 1991 949 1995
rect 958 1995 959 1999
rect 963 1995 964 1999
rect 1014 1999 1020 2000
rect 958 1994 964 1995
rect 991 1995 997 1996
rect 943 1990 949 1991
rect 991 1991 992 1995
rect 996 1994 997 1995
rect 999 1995 1005 1996
rect 999 1994 1000 1995
rect 996 1992 1000 1994
rect 996 1991 997 1992
rect 991 1990 997 1991
rect 999 1991 1000 1992
rect 1004 1991 1005 1995
rect 1014 1995 1015 1999
rect 1019 1995 1020 1999
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1426 1999 1427 2003
rect 1431 1999 1432 2003
rect 1436 1999 1437 2003
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1590 2007 1596 2008
rect 1486 2002 1492 2003
rect 1519 2003 1528 2004
rect 1426 1998 1437 1999
rect 1519 1999 1520 2003
rect 1527 1999 1528 2003
rect 1590 2003 1591 2007
rect 1595 2003 1596 2007
rect 1590 2002 1596 2003
rect 1616 2002 1618 2012
rect 1686 2011 1687 2015
rect 1691 2014 1692 2015
rect 2054 2015 2060 2016
rect 1691 2012 1818 2014
rect 1691 2011 1692 2012
rect 1686 2010 1692 2011
rect 1694 2007 1700 2008
rect 1623 2003 1629 2004
rect 1623 2002 1624 2003
rect 1616 2000 1624 2002
rect 1519 1998 1528 1999
rect 1623 1999 1624 2000
rect 1628 1999 1629 2003
rect 1694 2003 1695 2007
rect 1699 2003 1700 2007
rect 1790 2007 1796 2008
rect 1694 2002 1700 2003
rect 1727 2003 1733 2004
rect 1623 1998 1629 1999
rect 1727 1999 1728 2003
rect 1732 2002 1733 2003
rect 1758 2003 1764 2004
rect 1758 2002 1759 2003
rect 1732 2000 1759 2002
rect 1732 1999 1733 2000
rect 1727 1998 1733 1999
rect 1758 1999 1759 2000
rect 1763 1999 1764 2003
rect 1790 2003 1791 2007
rect 1795 2003 1796 2007
rect 1790 2002 1796 2003
rect 1816 2002 1818 2012
rect 2054 2011 2055 2015
rect 2059 2014 2060 2015
rect 2059 2012 2338 2014
rect 2059 2011 2060 2012
rect 2054 2010 2060 2011
rect 1886 2007 1892 2008
rect 1823 2003 1829 2004
rect 1823 2002 1824 2003
rect 1816 2000 1824 2002
rect 1758 1998 1764 1999
rect 1823 1999 1824 2000
rect 1828 1999 1829 2003
rect 1886 2003 1887 2007
rect 1891 2003 1892 2007
rect 1990 2007 1996 2008
rect 1886 2002 1892 2003
rect 1918 2003 1925 2004
rect 1823 1998 1829 1999
rect 1918 1999 1919 2003
rect 1924 1999 1925 2003
rect 1990 2003 1991 2007
rect 1995 2003 1996 2007
rect 2094 2007 2100 2008
rect 1990 2002 1996 2003
rect 2023 2003 2029 2004
rect 1918 1998 1925 1999
rect 2023 1999 2024 2003
rect 2028 2002 2029 2003
rect 2031 2003 2037 2004
rect 2031 2002 2032 2003
rect 2028 2000 2032 2002
rect 2028 1999 2029 2000
rect 2023 1998 2029 1999
rect 2031 1999 2032 2000
rect 2036 1999 2037 2003
rect 2094 2003 2095 2007
rect 2099 2003 2100 2007
rect 2198 2007 2204 2008
rect 2094 2002 2100 2003
rect 2127 2003 2136 2004
rect 2031 1998 2037 1999
rect 2127 1999 2128 2003
rect 2135 1999 2136 2003
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2310 2007 2316 2008
rect 2198 2002 2204 2003
rect 2231 2003 2240 2004
rect 2127 1998 2136 1999
rect 2231 1999 2232 2003
rect 2239 1999 2240 2003
rect 2310 2003 2311 2007
rect 2315 2003 2316 2007
rect 2310 2002 2316 2003
rect 2336 2002 2338 2012
rect 2582 2008 2588 2009
rect 2430 2007 2436 2008
rect 2343 2003 2349 2004
rect 2343 2002 2344 2003
rect 2336 2000 2344 2002
rect 2231 1998 2240 1999
rect 2343 1999 2344 2000
rect 2348 1999 2349 2003
rect 2430 2003 2431 2007
rect 2435 2003 2436 2007
rect 2526 2007 2532 2008
rect 2430 2002 2436 2003
rect 2463 2003 2469 2004
rect 2343 1998 2349 1999
rect 2463 1999 2464 2003
rect 2468 2002 2469 2003
rect 2471 2003 2477 2004
rect 2471 2002 2472 2003
rect 2468 2000 2472 2002
rect 2468 1999 2469 2000
rect 2463 1998 2469 1999
rect 2471 1999 2472 2000
rect 2476 1999 2477 2003
rect 2526 2003 2527 2007
rect 2531 2003 2532 2007
rect 2582 2004 2583 2008
rect 2587 2004 2588 2008
rect 2526 2002 2532 2003
rect 2558 2003 2565 2004
rect 2582 2003 2588 2004
rect 2471 1998 2477 1999
rect 2558 1999 2559 2003
rect 2564 1999 2565 2003
rect 2558 1998 2565 1999
rect 1014 1994 1020 1995
rect 1046 1995 1053 1996
rect 1326 1995 1332 1996
rect 999 1990 1005 1991
rect 1046 1991 1047 1995
rect 1052 1991 1053 1995
rect 1046 1990 1053 1991
rect 595 1984 698 1986
rect 595 1983 596 1984
rect 590 1982 596 1983
rect 1606 1983 1612 1984
rect 1494 1979 1500 1980
rect 1431 1975 1437 1976
rect 1398 1973 1404 1974
rect 1366 1972 1372 1973
rect 358 1971 364 1972
rect 358 1967 359 1971
rect 363 1970 364 1971
rect 363 1968 539 1970
rect 1366 1968 1367 1972
rect 1371 1968 1372 1972
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1431 1971 1432 1975
rect 1436 1974 1437 1975
rect 1470 1975 1476 1976
rect 1470 1974 1471 1975
rect 1436 1972 1471 1974
rect 1436 1971 1437 1972
rect 1431 1970 1437 1971
rect 1470 1971 1471 1972
rect 1475 1971 1476 1975
rect 1494 1975 1495 1979
rect 1499 1978 1500 1979
rect 1606 1979 1607 1983
rect 1611 1982 1612 1983
rect 1894 1983 1900 1984
rect 1611 1980 1794 1982
rect 1611 1979 1612 1980
rect 1606 1978 1612 1979
rect 1499 1976 1506 1978
rect 1499 1975 1500 1976
rect 1494 1974 1500 1975
rect 1504 1974 1506 1976
rect 1511 1975 1517 1976
rect 1511 1974 1512 1975
rect 1470 1970 1476 1971
rect 1478 1973 1484 1974
rect 1398 1968 1404 1969
rect 1478 1969 1479 1973
rect 1483 1969 1484 1973
rect 1504 1972 1512 1974
rect 1511 1971 1512 1972
rect 1516 1971 1517 1975
rect 1615 1975 1621 1976
rect 1511 1970 1517 1971
rect 1582 1973 1588 1974
rect 1478 1968 1484 1969
rect 1582 1969 1583 1973
rect 1587 1969 1588 1973
rect 1615 1971 1616 1975
rect 1620 1974 1621 1975
rect 1670 1975 1676 1976
rect 1670 1974 1671 1975
rect 1620 1972 1671 1974
rect 1620 1971 1621 1972
rect 1615 1970 1621 1971
rect 1670 1971 1671 1972
rect 1675 1971 1676 1975
rect 1706 1975 1717 1976
rect 1670 1970 1676 1971
rect 1678 1973 1684 1974
rect 1582 1968 1588 1969
rect 1678 1969 1679 1973
rect 1683 1969 1684 1973
rect 1706 1971 1707 1975
rect 1711 1971 1712 1975
rect 1716 1971 1717 1975
rect 1792 1974 1794 1980
rect 1894 1979 1895 1983
rect 1899 1982 1900 1983
rect 1899 1980 2114 1982
rect 1899 1979 1900 1980
rect 1894 1978 1900 1979
rect 1799 1975 1805 1976
rect 1799 1974 1800 1975
rect 1706 1970 1717 1971
rect 1766 1973 1772 1974
rect 1678 1968 1684 1969
rect 1766 1969 1767 1973
rect 1771 1969 1772 1973
rect 1792 1972 1800 1974
rect 1799 1971 1800 1972
rect 1804 1971 1805 1975
rect 1879 1975 1885 1976
rect 1799 1970 1805 1971
rect 1846 1973 1852 1974
rect 1766 1968 1772 1969
rect 1846 1969 1847 1973
rect 1851 1969 1852 1973
rect 1879 1971 1880 1975
rect 1884 1974 1885 1975
rect 1918 1975 1924 1976
rect 1918 1974 1919 1975
rect 1884 1972 1919 1974
rect 1884 1971 1885 1972
rect 1879 1970 1885 1971
rect 1918 1971 1919 1972
rect 1923 1971 1924 1975
rect 1959 1975 1965 1976
rect 1918 1970 1924 1971
rect 1926 1973 1932 1974
rect 1846 1968 1852 1969
rect 1926 1969 1927 1973
rect 1931 1969 1932 1973
rect 1959 1971 1960 1975
rect 1964 1974 1965 1975
rect 1998 1975 2004 1976
rect 1998 1974 1999 1975
rect 1964 1972 1999 1974
rect 1964 1971 1965 1972
rect 1959 1970 1965 1971
rect 1998 1971 1999 1972
rect 2003 1971 2004 1975
rect 2039 1975 2045 1976
rect 1998 1970 2004 1971
rect 2006 1973 2012 1974
rect 1926 1968 1932 1969
rect 2006 1969 2007 1973
rect 2011 1969 2012 1973
rect 2039 1971 2040 1975
rect 2044 1974 2045 1975
rect 2078 1975 2084 1976
rect 2078 1974 2079 1975
rect 2044 1972 2079 1974
rect 2044 1971 2045 1972
rect 2039 1970 2045 1971
rect 2078 1971 2079 1972
rect 2083 1971 2084 1975
rect 2112 1974 2114 1980
rect 2119 1975 2125 1976
rect 2119 1974 2120 1975
rect 2078 1970 2084 1971
rect 2086 1973 2092 1974
rect 2006 1968 2012 1969
rect 2086 1969 2087 1973
rect 2091 1969 2092 1973
rect 2112 1972 2120 1974
rect 2119 1971 2120 1972
rect 2124 1971 2125 1975
rect 2119 1970 2125 1971
rect 2582 1972 2588 1973
rect 2086 1968 2092 1969
rect 2582 1968 2583 1972
rect 2587 1968 2588 1972
rect 363 1967 364 1968
rect 358 1966 364 1967
rect 537 1964 539 1968
rect 543 1967 549 1968
rect 1366 1967 1372 1968
rect 2582 1967 2588 1968
rect 367 1963 373 1964
rect 334 1961 340 1962
rect 110 1960 116 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 334 1957 335 1961
rect 339 1957 340 1961
rect 367 1959 368 1963
rect 372 1962 373 1963
rect 382 1963 388 1964
rect 382 1962 383 1963
rect 372 1960 383 1962
rect 372 1959 373 1960
rect 367 1958 373 1959
rect 382 1959 383 1960
rect 387 1959 388 1963
rect 423 1963 429 1964
rect 382 1958 388 1959
rect 390 1961 396 1962
rect 334 1956 340 1957
rect 390 1957 391 1961
rect 395 1957 396 1961
rect 423 1959 424 1963
rect 428 1962 429 1963
rect 438 1963 444 1964
rect 438 1962 439 1963
rect 428 1960 439 1962
rect 428 1959 429 1960
rect 423 1958 429 1959
rect 438 1959 439 1960
rect 443 1959 444 1963
rect 479 1963 485 1964
rect 438 1958 444 1959
rect 446 1961 452 1962
rect 390 1956 396 1957
rect 446 1957 447 1961
rect 451 1957 452 1961
rect 479 1959 480 1963
rect 484 1962 485 1963
rect 494 1963 500 1964
rect 494 1962 495 1963
rect 484 1960 495 1962
rect 484 1959 485 1960
rect 479 1958 485 1959
rect 494 1959 495 1960
rect 499 1959 500 1963
rect 535 1963 541 1964
rect 494 1958 500 1959
rect 502 1961 508 1962
rect 446 1956 452 1957
rect 502 1957 503 1961
rect 507 1957 508 1961
rect 535 1959 536 1963
rect 540 1959 541 1963
rect 543 1963 544 1967
rect 548 1966 549 1967
rect 548 1964 603 1966
rect 548 1963 549 1964
rect 543 1962 549 1963
rect 599 1963 605 1964
rect 535 1958 541 1959
rect 566 1961 572 1962
rect 502 1956 508 1957
rect 566 1957 567 1961
rect 571 1957 572 1961
rect 599 1959 600 1963
rect 604 1959 605 1963
rect 679 1963 685 1964
rect 599 1958 605 1959
rect 646 1961 652 1962
rect 566 1956 572 1957
rect 646 1957 647 1961
rect 651 1957 652 1961
rect 679 1959 680 1963
rect 684 1962 685 1963
rect 734 1963 740 1964
rect 734 1962 735 1963
rect 684 1960 735 1962
rect 684 1959 685 1960
rect 679 1958 685 1959
rect 734 1959 735 1960
rect 739 1959 740 1963
rect 775 1963 781 1964
rect 734 1958 740 1959
rect 742 1961 748 1962
rect 646 1956 652 1957
rect 742 1957 743 1961
rect 747 1957 748 1961
rect 775 1959 776 1963
rect 780 1962 781 1963
rect 854 1963 860 1964
rect 854 1962 855 1963
rect 780 1960 855 1962
rect 780 1959 781 1960
rect 775 1958 781 1959
rect 854 1959 855 1960
rect 859 1959 860 1963
rect 895 1963 901 1964
rect 854 1958 860 1959
rect 862 1961 868 1962
rect 742 1956 748 1957
rect 862 1957 863 1961
rect 867 1957 868 1961
rect 895 1959 896 1963
rect 900 1962 901 1963
rect 990 1963 996 1964
rect 990 1962 991 1963
rect 900 1960 991 1962
rect 900 1959 901 1960
rect 895 1958 901 1959
rect 990 1959 991 1960
rect 995 1959 996 1963
rect 1031 1963 1037 1964
rect 990 1958 996 1959
rect 998 1961 1004 1962
rect 862 1956 868 1957
rect 998 1957 999 1961
rect 1003 1957 1004 1961
rect 1031 1959 1032 1963
rect 1036 1962 1037 1963
rect 1134 1963 1140 1964
rect 1134 1962 1135 1963
rect 1036 1960 1135 1962
rect 1036 1959 1037 1960
rect 1031 1958 1037 1959
rect 1134 1959 1135 1960
rect 1139 1959 1140 1963
rect 1174 1963 1181 1964
rect 1134 1958 1140 1959
rect 1142 1961 1148 1962
rect 998 1956 1004 1957
rect 1142 1957 1143 1961
rect 1147 1957 1148 1961
rect 1174 1959 1175 1963
rect 1180 1959 1181 1963
rect 1303 1963 1309 1964
rect 1174 1958 1181 1959
rect 1270 1961 1276 1962
rect 1142 1956 1148 1957
rect 1270 1957 1271 1961
rect 1275 1957 1276 1961
rect 1303 1959 1304 1963
rect 1308 1962 1309 1963
rect 1308 1960 1322 1962
rect 1308 1959 1309 1960
rect 1303 1958 1309 1959
rect 1270 1956 1276 1957
rect 110 1955 116 1956
rect 1320 1950 1322 1960
rect 1326 1960 1332 1961
rect 1326 1956 1327 1960
rect 1331 1956 1332 1960
rect 1326 1955 1332 1956
rect 1366 1955 1372 1956
rect 1366 1951 1367 1955
rect 1371 1951 1372 1955
rect 1366 1950 1372 1951
rect 2582 1955 2588 1956
rect 2582 1951 2583 1955
rect 2587 1951 2588 1955
rect 2582 1950 2588 1951
rect 1320 1948 1350 1950
rect 110 1943 116 1944
rect 110 1939 111 1943
rect 115 1939 116 1943
rect 110 1938 116 1939
rect 1326 1943 1332 1944
rect 1326 1939 1327 1943
rect 1331 1939 1332 1943
rect 1326 1938 1332 1939
rect 1348 1938 1350 1948
rect 1414 1946 1420 1947
rect 1414 1942 1415 1946
rect 1419 1942 1420 1946
rect 1414 1941 1420 1942
rect 1494 1946 1500 1947
rect 1494 1942 1495 1946
rect 1499 1942 1500 1946
rect 1494 1941 1500 1942
rect 1598 1946 1604 1947
rect 1598 1942 1599 1946
rect 1603 1942 1604 1946
rect 1598 1941 1604 1942
rect 1694 1946 1700 1947
rect 1694 1942 1695 1946
rect 1699 1942 1700 1946
rect 1694 1941 1700 1942
rect 1782 1946 1788 1947
rect 1782 1942 1783 1946
rect 1787 1942 1788 1946
rect 1782 1941 1788 1942
rect 1862 1946 1868 1947
rect 1862 1942 1863 1946
rect 1867 1942 1868 1946
rect 1862 1941 1868 1942
rect 1942 1946 1948 1947
rect 1942 1942 1943 1946
rect 1947 1942 1948 1946
rect 1942 1941 1948 1942
rect 2022 1946 2028 1947
rect 2022 1942 2023 1946
rect 2027 1942 2028 1946
rect 2022 1941 2028 1942
rect 2102 1946 2108 1947
rect 2102 1942 2103 1946
rect 2107 1942 2108 1946
rect 2102 1941 2108 1942
rect 1391 1939 1397 1940
rect 1391 1938 1392 1939
rect 1348 1936 1392 1938
rect 1391 1935 1392 1936
rect 1396 1935 1397 1939
rect 350 1934 356 1935
rect 350 1930 351 1934
rect 355 1930 356 1934
rect 350 1929 356 1930
rect 406 1934 412 1935
rect 406 1930 407 1934
rect 411 1930 412 1934
rect 406 1929 412 1930
rect 462 1934 468 1935
rect 462 1930 463 1934
rect 467 1930 468 1934
rect 462 1929 468 1930
rect 518 1934 524 1935
rect 518 1930 519 1934
rect 523 1930 524 1934
rect 518 1929 524 1930
rect 582 1934 588 1935
rect 582 1930 583 1934
rect 587 1930 588 1934
rect 582 1929 588 1930
rect 662 1934 668 1935
rect 662 1930 663 1934
rect 667 1930 668 1934
rect 662 1929 668 1930
rect 758 1934 764 1935
rect 758 1930 759 1934
rect 763 1930 764 1934
rect 758 1929 764 1930
rect 878 1934 884 1935
rect 878 1930 879 1934
rect 883 1930 884 1934
rect 878 1929 884 1930
rect 1014 1934 1020 1935
rect 1014 1930 1015 1934
rect 1019 1930 1020 1934
rect 1014 1929 1020 1930
rect 1158 1934 1164 1935
rect 1158 1930 1159 1934
rect 1163 1930 1164 1934
rect 1158 1929 1164 1930
rect 1286 1934 1292 1935
rect 1391 1934 1397 1935
rect 1470 1939 1477 1940
rect 1470 1935 1471 1939
rect 1476 1935 1477 1939
rect 1470 1934 1477 1935
rect 1575 1939 1581 1940
rect 1575 1935 1576 1939
rect 1580 1938 1581 1939
rect 1606 1939 1612 1940
rect 1606 1938 1607 1939
rect 1580 1936 1607 1938
rect 1580 1935 1581 1936
rect 1575 1934 1581 1935
rect 1606 1935 1607 1936
rect 1611 1935 1612 1939
rect 1606 1934 1612 1935
rect 1670 1939 1677 1940
rect 1670 1935 1671 1939
rect 1676 1935 1677 1939
rect 1670 1934 1677 1935
rect 1758 1939 1765 1940
rect 1758 1935 1759 1939
rect 1764 1935 1765 1939
rect 1758 1934 1765 1935
rect 1839 1939 1848 1940
rect 1839 1935 1840 1939
rect 1847 1935 1848 1939
rect 1839 1934 1848 1935
rect 1918 1939 1925 1940
rect 1918 1935 1919 1939
rect 1924 1935 1925 1939
rect 1918 1934 1925 1935
rect 1998 1939 2005 1940
rect 1998 1935 1999 1939
rect 2004 1935 2005 1939
rect 1998 1934 2005 1935
rect 2078 1939 2085 1940
rect 2078 1935 2079 1939
rect 2084 1935 2085 1939
rect 2078 1934 2085 1935
rect 1286 1930 1287 1934
rect 1291 1930 1292 1934
rect 1958 1931 1964 1932
rect 1958 1930 1959 1931
rect 1286 1929 1292 1930
rect 1880 1928 1959 1930
rect 327 1927 333 1928
rect 327 1923 328 1927
rect 332 1926 333 1927
rect 358 1927 364 1928
rect 358 1926 359 1927
rect 332 1924 359 1926
rect 332 1923 333 1924
rect 327 1922 333 1923
rect 358 1923 359 1924
rect 363 1923 364 1927
rect 358 1922 364 1923
rect 382 1927 389 1928
rect 382 1923 383 1927
rect 388 1923 389 1927
rect 382 1922 389 1923
rect 438 1927 445 1928
rect 438 1923 439 1927
rect 444 1923 445 1927
rect 438 1922 445 1923
rect 495 1927 501 1928
rect 495 1923 496 1927
rect 500 1926 501 1927
rect 543 1927 549 1928
rect 543 1926 544 1927
rect 500 1924 544 1926
rect 500 1923 501 1924
rect 495 1922 501 1923
rect 543 1923 544 1924
rect 548 1923 549 1927
rect 543 1922 549 1923
rect 559 1927 565 1928
rect 559 1923 560 1927
rect 564 1926 565 1927
rect 590 1927 596 1928
rect 590 1926 591 1927
rect 564 1924 591 1926
rect 564 1923 565 1924
rect 559 1922 565 1923
rect 590 1923 591 1924
rect 595 1923 596 1927
rect 590 1922 596 1923
rect 639 1927 645 1928
rect 639 1923 640 1927
rect 644 1926 645 1927
rect 670 1927 676 1928
rect 670 1926 671 1927
rect 644 1924 671 1926
rect 644 1923 645 1924
rect 639 1922 645 1923
rect 670 1923 671 1924
rect 675 1923 676 1927
rect 670 1922 676 1923
rect 734 1927 741 1928
rect 734 1923 735 1927
rect 740 1923 741 1927
rect 734 1922 741 1923
rect 854 1927 861 1928
rect 854 1923 855 1927
rect 860 1923 861 1927
rect 854 1922 861 1923
rect 990 1927 997 1928
rect 990 1923 991 1927
rect 996 1923 997 1927
rect 990 1922 997 1923
rect 1134 1927 1141 1928
rect 1134 1923 1135 1927
rect 1140 1923 1141 1927
rect 1134 1922 1141 1923
rect 1218 1927 1224 1928
rect 1218 1923 1219 1927
rect 1223 1926 1224 1927
rect 1263 1927 1269 1928
rect 1263 1926 1264 1927
rect 1223 1924 1264 1926
rect 1223 1923 1224 1924
rect 1218 1922 1224 1923
rect 1263 1923 1264 1924
rect 1268 1923 1269 1927
rect 1706 1927 1712 1928
rect 1706 1926 1707 1927
rect 1263 1922 1269 1923
rect 1695 1925 1707 1926
rect 1695 1921 1696 1925
rect 1700 1924 1707 1925
rect 1700 1921 1701 1924
rect 1706 1923 1707 1924
rect 1711 1923 1712 1927
rect 1706 1922 1712 1923
rect 1738 1923 1744 1924
rect 1695 1920 1701 1921
rect 846 1919 852 1920
rect 1738 1919 1739 1923
rect 1743 1922 1744 1923
rect 1751 1923 1757 1924
rect 1751 1922 1752 1923
rect 1743 1920 1752 1922
rect 1743 1919 1744 1920
rect 846 1918 847 1919
rect 760 1916 847 1918
rect 134 1915 141 1916
rect 134 1911 135 1915
rect 140 1911 141 1915
rect 207 1915 213 1916
rect 207 1911 208 1915
rect 212 1914 213 1915
rect 222 1915 228 1916
rect 222 1914 223 1915
rect 212 1912 223 1914
rect 212 1911 213 1912
rect 134 1910 141 1911
rect 158 1910 164 1911
rect 207 1910 213 1911
rect 222 1911 223 1912
rect 227 1911 228 1915
rect 302 1915 309 1916
rect 302 1911 303 1915
rect 308 1911 309 1915
rect 407 1915 413 1916
rect 407 1911 408 1915
rect 412 1914 413 1915
rect 422 1915 428 1916
rect 422 1914 423 1915
rect 412 1912 423 1914
rect 412 1911 413 1912
rect 222 1910 228 1911
rect 230 1910 236 1911
rect 302 1910 309 1911
rect 326 1910 332 1911
rect 407 1910 413 1911
rect 422 1911 423 1912
rect 427 1911 428 1915
rect 494 1915 500 1916
rect 494 1911 495 1915
rect 499 1914 500 1915
rect 519 1915 525 1916
rect 519 1914 520 1915
rect 499 1912 520 1914
rect 499 1911 500 1912
rect 422 1910 428 1911
rect 430 1910 436 1911
rect 494 1910 500 1911
rect 519 1911 520 1912
rect 524 1911 525 1915
rect 630 1915 637 1916
rect 630 1911 631 1915
rect 636 1911 637 1915
rect 743 1915 749 1916
rect 743 1911 744 1915
rect 748 1914 749 1915
rect 760 1914 762 1916
rect 846 1915 847 1916
rect 851 1915 852 1919
rect 1718 1918 1724 1919
rect 1738 1918 1744 1919
rect 1751 1919 1752 1920
rect 1756 1919 1757 1923
rect 1806 1923 1813 1924
rect 1806 1919 1807 1923
rect 1812 1919 1813 1923
rect 1863 1923 1869 1924
rect 1863 1919 1864 1923
rect 1868 1922 1869 1923
rect 1880 1922 1882 1928
rect 1958 1927 1959 1928
rect 1963 1927 1964 1931
rect 2134 1931 2140 1932
rect 2134 1930 2135 1931
rect 1958 1926 1964 1927
rect 1999 1928 2135 1930
rect 1999 1926 2001 1928
rect 2134 1927 2135 1928
rect 2139 1927 2140 1931
rect 2134 1926 2140 1927
rect 1988 1924 2001 1926
rect 1868 1920 1882 1922
rect 1918 1923 1925 1924
rect 1868 1919 1869 1920
rect 1918 1919 1919 1923
rect 1924 1919 1925 1923
rect 1975 1923 1981 1924
rect 1975 1919 1976 1923
rect 1980 1922 1981 1923
rect 1988 1922 1990 1924
rect 1980 1920 1990 1922
rect 2030 1923 2037 1924
rect 1980 1919 1981 1920
rect 2030 1919 2031 1923
rect 2036 1919 2037 1923
rect 2079 1923 2085 1924
rect 2079 1919 2080 1923
rect 2084 1922 2085 1923
rect 2095 1923 2101 1924
rect 2095 1922 2096 1923
rect 2084 1920 2096 1922
rect 2084 1919 2085 1920
rect 1751 1918 1757 1919
rect 1774 1918 1780 1919
rect 1806 1918 1813 1919
rect 1830 1918 1836 1919
rect 1863 1918 1869 1919
rect 1886 1918 1892 1919
rect 1918 1918 1925 1919
rect 1942 1918 1948 1919
rect 1975 1918 1981 1919
rect 1998 1918 2004 1919
rect 2030 1918 2037 1919
rect 2054 1918 2060 1919
rect 2079 1918 2085 1919
rect 2095 1919 2096 1920
rect 2100 1919 2101 1923
rect 2095 1918 2101 1919
rect 2118 1918 2124 1919
rect 846 1914 852 1915
rect 854 1915 861 1916
rect 748 1912 762 1914
rect 748 1911 749 1912
rect 854 1911 855 1915
rect 860 1911 861 1915
rect 959 1915 965 1916
rect 959 1911 960 1915
rect 964 1914 965 1915
rect 974 1915 980 1916
rect 974 1914 975 1915
rect 964 1912 975 1914
rect 964 1911 965 1912
rect 519 1910 525 1911
rect 542 1910 548 1911
rect 630 1910 637 1911
rect 654 1910 660 1911
rect 743 1910 749 1911
rect 766 1910 772 1911
rect 854 1910 861 1911
rect 878 1910 884 1911
rect 959 1910 965 1911
rect 974 1911 975 1912
rect 979 1911 980 1915
rect 1062 1915 1069 1916
rect 1062 1911 1063 1915
rect 1068 1911 1069 1915
rect 1106 1915 1112 1916
rect 1106 1911 1107 1915
rect 1111 1914 1112 1915
rect 1175 1915 1181 1916
rect 1175 1914 1176 1915
rect 1111 1912 1176 1914
rect 1111 1911 1112 1912
rect 974 1910 980 1911
rect 982 1910 988 1911
rect 1062 1910 1069 1911
rect 1086 1910 1092 1911
rect 1106 1910 1112 1911
rect 1175 1911 1176 1912
rect 1180 1911 1181 1915
rect 1263 1915 1269 1916
rect 1263 1911 1264 1915
rect 1268 1914 1269 1915
rect 1278 1915 1284 1916
rect 1278 1914 1279 1915
rect 1268 1912 1279 1914
rect 1268 1911 1269 1912
rect 1175 1910 1181 1911
rect 1198 1910 1204 1911
rect 1263 1910 1269 1911
rect 1278 1911 1279 1912
rect 1283 1911 1284 1915
rect 1718 1914 1719 1918
rect 1723 1914 1724 1918
rect 1718 1913 1724 1914
rect 1774 1914 1775 1918
rect 1779 1914 1780 1918
rect 1774 1913 1780 1914
rect 1830 1914 1831 1918
rect 1835 1914 1836 1918
rect 1830 1913 1836 1914
rect 1886 1914 1887 1918
rect 1891 1914 1892 1918
rect 1886 1913 1892 1914
rect 1942 1914 1943 1918
rect 1947 1914 1948 1918
rect 1942 1913 1948 1914
rect 1998 1914 1999 1918
rect 2003 1914 2004 1918
rect 1998 1913 2004 1914
rect 2054 1914 2055 1918
rect 2059 1914 2060 1918
rect 2054 1913 2060 1914
rect 2118 1914 2119 1918
rect 2123 1914 2124 1918
rect 2118 1913 2124 1914
rect 1278 1910 1284 1911
rect 1286 1910 1292 1911
rect 158 1906 159 1910
rect 163 1906 164 1910
rect 158 1905 164 1906
rect 230 1906 231 1910
rect 235 1906 236 1910
rect 230 1905 236 1906
rect 326 1906 327 1910
rect 331 1906 332 1910
rect 326 1905 332 1906
rect 430 1906 431 1910
rect 435 1906 436 1910
rect 430 1905 436 1906
rect 542 1906 543 1910
rect 547 1906 548 1910
rect 542 1905 548 1906
rect 654 1906 655 1910
rect 659 1906 660 1910
rect 654 1905 660 1906
rect 766 1906 767 1910
rect 771 1906 772 1910
rect 766 1905 772 1906
rect 878 1906 879 1910
rect 883 1906 884 1910
rect 878 1905 884 1906
rect 982 1906 983 1910
rect 987 1906 988 1910
rect 982 1905 988 1906
rect 1086 1906 1087 1910
rect 1091 1906 1092 1910
rect 1086 1905 1092 1906
rect 1198 1906 1199 1910
rect 1203 1906 1204 1910
rect 1198 1905 1204 1906
rect 1286 1906 1287 1910
rect 1291 1906 1292 1910
rect 1286 1905 1292 1906
rect 1366 1909 1372 1910
rect 1366 1905 1367 1909
rect 1371 1905 1372 1909
rect 1366 1904 1372 1905
rect 2582 1909 2588 1910
rect 2582 1905 2583 1909
rect 2587 1905 2588 1909
rect 2582 1904 2588 1905
rect 110 1901 116 1902
rect 110 1897 111 1901
rect 115 1897 116 1901
rect 110 1896 116 1897
rect 1326 1901 1332 1902
rect 1326 1897 1327 1901
rect 1331 1897 1332 1901
rect 1326 1896 1332 1897
rect 1806 1899 1812 1900
rect 1806 1895 1807 1899
rect 1811 1898 1812 1899
rect 1918 1899 1924 1900
rect 1811 1896 1898 1898
rect 1811 1895 1812 1896
rect 1806 1894 1812 1895
rect 1366 1892 1372 1893
rect 134 1891 140 1892
rect 134 1887 135 1891
rect 139 1890 140 1891
rect 302 1891 308 1892
rect 139 1888 242 1890
rect 139 1887 140 1888
rect 134 1886 140 1887
rect 110 1884 116 1885
rect 110 1880 111 1884
rect 115 1880 116 1884
rect 110 1879 116 1880
rect 142 1883 148 1884
rect 142 1879 143 1883
rect 147 1879 148 1883
rect 214 1883 220 1884
rect 142 1878 148 1879
rect 166 1879 172 1880
rect 166 1875 167 1879
rect 171 1878 172 1879
rect 175 1879 181 1880
rect 175 1878 176 1879
rect 171 1876 176 1878
rect 171 1875 172 1876
rect 166 1874 172 1875
rect 175 1875 176 1876
rect 180 1875 181 1879
rect 214 1879 215 1883
rect 219 1879 220 1883
rect 214 1878 220 1879
rect 240 1878 242 1888
rect 302 1887 303 1891
rect 307 1890 308 1891
rect 630 1891 636 1892
rect 307 1888 442 1890
rect 307 1887 308 1888
rect 302 1886 308 1887
rect 310 1883 316 1884
rect 247 1879 253 1880
rect 247 1878 248 1879
rect 240 1876 248 1878
rect 175 1874 181 1875
rect 247 1875 248 1876
rect 252 1875 253 1879
rect 310 1879 311 1883
rect 315 1879 316 1883
rect 414 1883 420 1884
rect 310 1878 316 1879
rect 343 1879 349 1880
rect 343 1878 344 1879
rect 247 1874 253 1875
rect 319 1876 344 1878
rect 222 1871 228 1872
rect 222 1867 223 1871
rect 227 1870 228 1871
rect 319 1870 321 1876
rect 343 1875 344 1876
rect 348 1875 349 1879
rect 414 1879 415 1883
rect 419 1879 420 1883
rect 414 1878 420 1879
rect 440 1878 442 1888
rect 630 1887 631 1891
rect 635 1890 636 1891
rect 854 1891 860 1892
rect 635 1888 787 1890
rect 635 1887 636 1888
rect 630 1886 636 1887
rect 526 1883 532 1884
rect 447 1879 453 1880
rect 447 1878 448 1879
rect 440 1876 448 1878
rect 343 1874 349 1875
rect 447 1875 448 1876
rect 452 1875 453 1879
rect 526 1879 527 1883
rect 531 1879 532 1883
rect 638 1883 644 1884
rect 526 1878 532 1879
rect 559 1879 565 1880
rect 559 1878 560 1879
rect 447 1874 453 1875
rect 536 1876 560 1878
rect 227 1868 321 1870
rect 422 1871 428 1872
rect 227 1867 228 1868
rect 222 1866 228 1867
rect 422 1867 423 1871
rect 427 1870 428 1871
rect 536 1870 538 1876
rect 559 1875 560 1876
rect 564 1875 565 1879
rect 638 1879 639 1883
rect 643 1879 644 1883
rect 750 1883 756 1884
rect 638 1878 644 1879
rect 670 1879 677 1880
rect 559 1874 565 1875
rect 670 1875 671 1879
rect 676 1875 677 1879
rect 750 1879 751 1883
rect 755 1879 756 1883
rect 785 1880 787 1888
rect 854 1887 855 1891
rect 859 1890 860 1891
rect 1062 1891 1068 1892
rect 859 1888 1003 1890
rect 859 1887 860 1888
rect 854 1886 860 1887
rect 862 1883 868 1884
rect 750 1878 756 1879
rect 783 1879 789 1880
rect 670 1874 677 1875
rect 783 1875 784 1879
rect 788 1875 789 1879
rect 862 1879 863 1883
rect 867 1879 868 1883
rect 966 1883 972 1884
rect 862 1878 868 1879
rect 895 1879 901 1880
rect 895 1878 896 1879
rect 872 1876 896 1878
rect 783 1874 789 1875
rect 846 1875 852 1876
rect 846 1871 847 1875
rect 851 1874 852 1875
rect 872 1874 874 1876
rect 895 1875 896 1876
rect 900 1875 901 1879
rect 966 1879 967 1883
rect 971 1879 972 1883
rect 1001 1880 1003 1888
rect 1062 1887 1063 1891
rect 1067 1890 1068 1891
rect 1067 1888 1298 1890
rect 1067 1887 1068 1888
rect 1062 1886 1068 1887
rect 1070 1883 1076 1884
rect 966 1878 972 1879
rect 999 1879 1005 1880
rect 895 1874 901 1875
rect 999 1875 1000 1879
rect 1004 1875 1005 1879
rect 1070 1879 1071 1883
rect 1075 1879 1076 1883
rect 1182 1883 1188 1884
rect 1070 1878 1076 1879
rect 1103 1879 1112 1880
rect 999 1874 1005 1875
rect 1103 1875 1104 1879
rect 1111 1875 1112 1879
rect 1182 1879 1183 1883
rect 1187 1879 1188 1883
rect 1270 1883 1276 1884
rect 1182 1878 1188 1879
rect 1215 1879 1224 1880
rect 1103 1874 1112 1875
rect 1215 1875 1216 1879
rect 1223 1875 1224 1879
rect 1270 1879 1271 1883
rect 1275 1879 1276 1883
rect 1270 1878 1276 1879
rect 1296 1878 1298 1888
rect 1366 1888 1367 1892
rect 1371 1888 1372 1892
rect 1366 1887 1372 1888
rect 1702 1891 1708 1892
rect 1702 1887 1703 1891
rect 1707 1887 1708 1891
rect 1758 1891 1764 1892
rect 1702 1886 1708 1887
rect 1735 1887 1744 1888
rect 1326 1884 1332 1885
rect 1326 1880 1327 1884
rect 1331 1880 1332 1884
rect 1735 1883 1736 1887
rect 1743 1883 1744 1887
rect 1758 1887 1759 1891
rect 1763 1887 1764 1891
rect 1814 1891 1820 1892
rect 1758 1886 1764 1887
rect 1782 1887 1788 1888
rect 1735 1882 1744 1883
rect 1782 1883 1783 1887
rect 1787 1886 1788 1887
rect 1791 1887 1797 1888
rect 1791 1886 1792 1887
rect 1787 1884 1792 1886
rect 1787 1883 1788 1884
rect 1782 1882 1788 1883
rect 1791 1883 1792 1884
rect 1796 1883 1797 1887
rect 1814 1887 1815 1891
rect 1819 1887 1820 1891
rect 1870 1891 1876 1892
rect 1814 1886 1820 1887
rect 1842 1887 1853 1888
rect 1791 1882 1797 1883
rect 1842 1883 1843 1887
rect 1847 1883 1848 1887
rect 1852 1883 1853 1887
rect 1870 1887 1871 1891
rect 1875 1887 1876 1891
rect 1870 1886 1876 1887
rect 1896 1886 1898 1896
rect 1918 1895 1919 1899
rect 1923 1898 1924 1899
rect 1923 1896 2010 1898
rect 1923 1895 1924 1896
rect 1918 1894 1924 1895
rect 1926 1891 1932 1892
rect 1903 1887 1909 1888
rect 1903 1886 1904 1887
rect 1896 1884 1904 1886
rect 1842 1882 1853 1883
rect 1903 1883 1904 1884
rect 1908 1883 1909 1887
rect 1926 1887 1927 1891
rect 1931 1887 1932 1891
rect 1982 1891 1988 1892
rect 1926 1886 1932 1887
rect 1958 1887 1965 1888
rect 1903 1882 1909 1883
rect 1958 1883 1959 1887
rect 1964 1883 1965 1887
rect 1982 1887 1983 1891
rect 1987 1887 1988 1891
rect 1982 1886 1988 1887
rect 2008 1886 2010 1896
rect 2582 1892 2588 1893
rect 2038 1891 2044 1892
rect 2015 1887 2021 1888
rect 2015 1886 2016 1887
rect 2008 1884 2016 1886
rect 1958 1882 1965 1883
rect 2015 1883 2016 1884
rect 2020 1883 2021 1887
rect 2038 1887 2039 1891
rect 2043 1887 2044 1891
rect 2102 1891 2108 1892
rect 2038 1886 2044 1887
rect 2071 1887 2077 1888
rect 2015 1882 2021 1883
rect 2071 1883 2072 1887
rect 2076 1886 2077 1887
rect 2079 1887 2085 1888
rect 2079 1886 2080 1887
rect 2076 1884 2080 1886
rect 2076 1883 2077 1884
rect 2071 1882 2077 1883
rect 2079 1883 2080 1884
rect 2084 1883 2085 1887
rect 2102 1887 2103 1891
rect 2107 1887 2108 1891
rect 2582 1888 2583 1892
rect 2587 1888 2588 1892
rect 2102 1886 2108 1887
rect 2134 1887 2141 1888
rect 2582 1887 2588 1888
rect 2079 1882 2085 1883
rect 2134 1883 2135 1887
rect 2140 1883 2141 1887
rect 2134 1882 2141 1883
rect 1303 1879 1309 1880
rect 1326 1879 1332 1880
rect 1303 1878 1304 1879
rect 1296 1876 1304 1878
rect 1215 1874 1224 1875
rect 1303 1875 1304 1876
rect 1308 1875 1309 1879
rect 1303 1874 1309 1875
rect 851 1872 874 1874
rect 851 1871 852 1872
rect 846 1870 852 1871
rect 427 1868 538 1870
rect 427 1867 428 1868
rect 422 1866 428 1867
rect 1278 1859 1284 1860
rect 1278 1855 1279 1859
rect 1283 1858 1284 1859
rect 1439 1859 1445 1860
rect 1283 1856 1435 1858
rect 1283 1855 1284 1856
rect 1278 1854 1284 1855
rect 1431 1855 1437 1856
rect 1398 1853 1404 1854
rect 1366 1852 1372 1853
rect 974 1851 980 1852
rect 974 1847 975 1851
rect 979 1850 980 1851
rect 979 1848 1066 1850
rect 979 1847 980 1848
rect 974 1846 980 1847
rect 175 1843 181 1844
rect 142 1841 148 1842
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 142 1837 143 1841
rect 147 1837 148 1841
rect 175 1839 176 1843
rect 180 1842 181 1843
rect 190 1843 196 1844
rect 190 1842 191 1843
rect 180 1840 191 1842
rect 180 1839 181 1840
rect 175 1838 181 1839
rect 190 1839 191 1840
rect 195 1839 196 1843
rect 231 1843 237 1844
rect 190 1838 196 1839
rect 198 1841 204 1842
rect 142 1836 148 1837
rect 198 1837 199 1841
rect 203 1837 204 1841
rect 231 1839 232 1843
rect 236 1842 237 1843
rect 254 1843 260 1844
rect 254 1842 255 1843
rect 236 1840 255 1842
rect 236 1839 237 1840
rect 231 1838 237 1839
rect 254 1839 255 1840
rect 259 1839 260 1843
rect 295 1843 301 1844
rect 254 1838 260 1839
rect 262 1841 268 1842
rect 198 1836 204 1837
rect 262 1837 263 1841
rect 267 1837 268 1841
rect 295 1839 296 1843
rect 300 1842 301 1843
rect 342 1843 348 1844
rect 342 1842 343 1843
rect 300 1840 343 1842
rect 300 1839 301 1840
rect 295 1838 301 1839
rect 342 1839 343 1840
rect 347 1839 348 1843
rect 383 1843 389 1844
rect 342 1838 348 1839
rect 350 1841 356 1842
rect 262 1836 268 1837
rect 350 1837 351 1841
rect 355 1837 356 1841
rect 383 1839 384 1843
rect 388 1842 389 1843
rect 430 1843 436 1844
rect 430 1842 431 1843
rect 388 1840 431 1842
rect 388 1839 389 1840
rect 383 1838 389 1839
rect 430 1839 431 1840
rect 435 1839 436 1843
rect 471 1843 477 1844
rect 430 1838 436 1839
rect 438 1841 444 1842
rect 350 1836 356 1837
rect 438 1837 439 1841
rect 443 1837 444 1841
rect 471 1839 472 1843
rect 476 1842 477 1843
rect 526 1843 532 1844
rect 526 1842 527 1843
rect 476 1840 527 1842
rect 476 1839 477 1840
rect 471 1838 477 1839
rect 526 1839 527 1840
rect 531 1839 532 1843
rect 558 1843 564 1844
rect 526 1838 532 1839
rect 534 1841 540 1842
rect 438 1836 444 1837
rect 534 1837 535 1841
rect 539 1837 540 1841
rect 558 1839 559 1843
rect 563 1842 564 1843
rect 567 1843 573 1844
rect 567 1842 568 1843
rect 563 1840 568 1842
rect 563 1839 564 1840
rect 558 1838 564 1839
rect 567 1839 568 1840
rect 572 1839 573 1843
rect 655 1843 661 1844
rect 567 1838 573 1839
rect 622 1841 628 1842
rect 534 1836 540 1837
rect 622 1837 623 1841
rect 627 1837 628 1841
rect 655 1839 656 1843
rect 660 1842 661 1843
rect 702 1843 708 1844
rect 702 1842 703 1843
rect 660 1840 703 1842
rect 660 1839 661 1840
rect 655 1838 661 1839
rect 702 1839 703 1840
rect 707 1839 708 1843
rect 743 1843 749 1844
rect 702 1838 708 1839
rect 710 1841 716 1842
rect 622 1836 628 1837
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 743 1839 744 1843
rect 748 1842 749 1843
rect 782 1843 788 1844
rect 782 1842 783 1843
rect 748 1840 783 1842
rect 748 1839 749 1840
rect 743 1838 749 1839
rect 782 1839 783 1840
rect 787 1839 788 1843
rect 823 1843 829 1844
rect 782 1838 788 1839
rect 790 1841 796 1842
rect 710 1836 716 1837
rect 790 1837 791 1841
rect 795 1837 796 1841
rect 823 1839 824 1843
rect 828 1842 829 1843
rect 862 1843 868 1844
rect 862 1842 863 1843
rect 828 1840 863 1842
rect 828 1839 829 1840
rect 823 1838 829 1839
rect 862 1839 863 1840
rect 867 1839 868 1843
rect 903 1843 909 1844
rect 862 1838 868 1839
rect 870 1841 876 1842
rect 790 1836 796 1837
rect 870 1837 871 1841
rect 875 1837 876 1841
rect 903 1839 904 1843
rect 908 1842 909 1843
rect 942 1843 948 1844
rect 942 1842 943 1843
rect 908 1840 943 1842
rect 908 1839 909 1840
rect 903 1838 909 1839
rect 942 1839 943 1840
rect 947 1839 948 1843
rect 983 1843 989 1844
rect 942 1838 948 1839
rect 950 1841 956 1842
rect 870 1836 876 1837
rect 950 1837 951 1841
rect 955 1837 956 1841
rect 983 1839 984 1843
rect 988 1842 989 1843
rect 1030 1843 1036 1844
rect 1030 1842 1031 1843
rect 988 1840 1031 1842
rect 988 1839 989 1840
rect 983 1838 989 1839
rect 1030 1839 1031 1840
rect 1035 1839 1036 1843
rect 1064 1842 1066 1848
rect 1366 1848 1367 1852
rect 1371 1848 1372 1852
rect 1398 1849 1399 1853
rect 1403 1849 1404 1853
rect 1431 1851 1432 1855
rect 1436 1851 1437 1855
rect 1439 1855 1440 1859
rect 1444 1858 1445 1859
rect 1503 1859 1509 1860
rect 1444 1856 1490 1858
rect 1444 1855 1445 1856
rect 1439 1854 1445 1855
rect 1488 1854 1490 1856
rect 1495 1855 1501 1856
rect 1495 1854 1496 1855
rect 1431 1850 1437 1851
rect 1462 1853 1468 1854
rect 1398 1848 1404 1849
rect 1462 1849 1463 1853
rect 1467 1849 1468 1853
rect 1488 1852 1496 1854
rect 1495 1851 1496 1852
rect 1500 1851 1501 1855
rect 1503 1855 1504 1859
rect 1508 1858 1509 1859
rect 1599 1859 1605 1860
rect 1508 1856 1586 1858
rect 1508 1855 1509 1856
rect 1503 1854 1509 1855
rect 1584 1854 1586 1856
rect 1591 1855 1597 1856
rect 1591 1854 1592 1855
rect 1495 1850 1501 1851
rect 1558 1853 1564 1854
rect 1462 1848 1468 1849
rect 1558 1849 1559 1853
rect 1563 1849 1564 1853
rect 1584 1852 1592 1854
rect 1591 1851 1592 1852
rect 1596 1851 1597 1855
rect 1599 1855 1600 1859
rect 1604 1858 1605 1859
rect 1714 1859 1720 1860
rect 1604 1856 1682 1858
rect 1604 1855 1605 1856
rect 1599 1854 1605 1855
rect 1680 1854 1682 1856
rect 1687 1855 1693 1856
rect 1687 1854 1688 1855
rect 1591 1850 1597 1851
rect 1654 1853 1660 1854
rect 1558 1848 1564 1849
rect 1654 1849 1655 1853
rect 1659 1849 1660 1853
rect 1680 1852 1688 1854
rect 1687 1851 1688 1852
rect 1692 1851 1693 1855
rect 1714 1855 1715 1859
rect 1719 1858 1720 1859
rect 1719 1856 1770 1858
rect 1719 1855 1720 1856
rect 1714 1854 1720 1855
rect 1768 1854 1770 1856
rect 1775 1855 1781 1856
rect 1775 1854 1776 1855
rect 1687 1850 1693 1851
rect 1742 1853 1748 1854
rect 1654 1848 1660 1849
rect 1742 1849 1743 1853
rect 1747 1849 1748 1853
rect 1768 1852 1776 1854
rect 1775 1851 1776 1852
rect 1780 1851 1781 1855
rect 1863 1855 1869 1856
rect 1775 1850 1781 1851
rect 1830 1853 1836 1854
rect 1742 1848 1748 1849
rect 1830 1849 1831 1853
rect 1835 1849 1836 1853
rect 1863 1851 1864 1855
rect 1868 1854 1869 1855
rect 1910 1855 1916 1856
rect 1910 1854 1911 1855
rect 1868 1852 1911 1854
rect 1868 1851 1869 1852
rect 1863 1850 1869 1851
rect 1910 1851 1911 1852
rect 1915 1851 1916 1855
rect 1951 1855 1957 1856
rect 1910 1850 1916 1851
rect 1918 1853 1924 1854
rect 1830 1848 1836 1849
rect 1918 1849 1919 1853
rect 1923 1849 1924 1853
rect 1951 1851 1952 1855
rect 1956 1854 1957 1855
rect 1998 1855 2004 1856
rect 1998 1854 1999 1855
rect 1956 1852 1999 1854
rect 1956 1851 1957 1852
rect 1951 1850 1957 1851
rect 1998 1851 1999 1852
rect 2003 1851 2004 1855
rect 2030 1855 2036 1856
rect 1998 1850 2004 1851
rect 2006 1853 2012 1854
rect 1918 1848 1924 1849
rect 2006 1849 2007 1853
rect 2011 1849 2012 1853
rect 2030 1851 2031 1855
rect 2035 1854 2036 1855
rect 2039 1855 2045 1856
rect 2039 1854 2040 1855
rect 2035 1852 2040 1854
rect 2035 1851 2036 1852
rect 2030 1850 2036 1851
rect 2039 1851 2040 1852
rect 2044 1851 2045 1855
rect 2127 1855 2133 1856
rect 2039 1850 2045 1851
rect 2094 1853 2100 1854
rect 2006 1848 2012 1849
rect 2094 1849 2095 1853
rect 2099 1849 2100 1853
rect 2127 1851 2128 1855
rect 2132 1854 2133 1855
rect 2174 1855 2180 1856
rect 2174 1854 2175 1855
rect 2132 1852 2175 1854
rect 2132 1851 2133 1852
rect 2127 1850 2133 1851
rect 2174 1851 2175 1852
rect 2179 1851 2180 1855
rect 2206 1855 2212 1856
rect 2174 1850 2180 1851
rect 2182 1853 2188 1854
rect 2094 1848 2100 1849
rect 2182 1849 2183 1853
rect 2187 1849 2188 1853
rect 2206 1851 2207 1855
rect 2211 1854 2212 1855
rect 2215 1855 2221 1856
rect 2215 1854 2216 1855
rect 2211 1852 2216 1854
rect 2211 1851 2212 1852
rect 2206 1850 2212 1851
rect 2215 1851 2216 1852
rect 2220 1851 2221 1855
rect 2215 1850 2221 1851
rect 2582 1852 2588 1853
rect 2182 1848 2188 1849
rect 2582 1848 2583 1852
rect 2587 1848 2588 1852
rect 1366 1847 1372 1848
rect 2582 1847 2588 1848
rect 1071 1843 1077 1844
rect 1071 1842 1072 1843
rect 1030 1838 1036 1839
rect 1038 1841 1044 1842
rect 950 1836 956 1837
rect 1038 1837 1039 1841
rect 1043 1837 1044 1841
rect 1064 1840 1072 1842
rect 1071 1839 1072 1840
rect 1076 1839 1077 1843
rect 1071 1838 1077 1839
rect 1326 1840 1332 1841
rect 1038 1836 1044 1837
rect 1326 1836 1327 1840
rect 1331 1836 1332 1840
rect 110 1835 116 1836
rect 1326 1835 1332 1836
rect 1366 1835 1372 1836
rect 1366 1831 1367 1835
rect 1371 1831 1372 1835
rect 1366 1830 1372 1831
rect 2582 1835 2588 1836
rect 2582 1831 2583 1835
rect 2587 1831 2588 1835
rect 2582 1830 2588 1831
rect 1414 1826 1420 1827
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 110 1818 116 1819
rect 1326 1823 1332 1824
rect 1326 1819 1327 1823
rect 1331 1819 1332 1823
rect 1414 1822 1415 1826
rect 1419 1822 1420 1826
rect 1414 1821 1420 1822
rect 1478 1826 1484 1827
rect 1478 1822 1479 1826
rect 1483 1822 1484 1826
rect 1478 1821 1484 1822
rect 1574 1826 1580 1827
rect 1574 1822 1575 1826
rect 1579 1822 1580 1826
rect 1574 1821 1580 1822
rect 1670 1826 1676 1827
rect 1670 1822 1671 1826
rect 1675 1822 1676 1826
rect 1670 1821 1676 1822
rect 1758 1826 1764 1827
rect 1758 1822 1759 1826
rect 1763 1822 1764 1826
rect 1758 1821 1764 1822
rect 1846 1826 1852 1827
rect 1846 1822 1847 1826
rect 1851 1822 1852 1826
rect 1846 1821 1852 1822
rect 1934 1826 1940 1827
rect 1934 1822 1935 1826
rect 1939 1822 1940 1826
rect 1934 1821 1940 1822
rect 2022 1826 2028 1827
rect 2022 1822 2023 1826
rect 2027 1822 2028 1826
rect 2022 1821 2028 1822
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2110 1821 2116 1822
rect 2198 1826 2204 1827
rect 2198 1822 2199 1826
rect 2203 1822 2204 1826
rect 2198 1821 2204 1822
rect 1326 1818 1332 1819
rect 1391 1819 1397 1820
rect 1391 1815 1392 1819
rect 1396 1818 1397 1819
rect 1439 1819 1445 1820
rect 1439 1818 1440 1819
rect 1396 1816 1440 1818
rect 1396 1815 1397 1816
rect 158 1814 164 1815
rect 158 1810 159 1814
rect 163 1810 164 1814
rect 158 1809 164 1810
rect 214 1814 220 1815
rect 214 1810 215 1814
rect 219 1810 220 1814
rect 214 1809 220 1810
rect 278 1814 284 1815
rect 278 1810 279 1814
rect 283 1810 284 1814
rect 278 1809 284 1810
rect 366 1814 372 1815
rect 366 1810 367 1814
rect 371 1810 372 1814
rect 366 1809 372 1810
rect 454 1814 460 1815
rect 454 1810 455 1814
rect 459 1810 460 1814
rect 454 1809 460 1810
rect 550 1814 556 1815
rect 550 1810 551 1814
rect 555 1810 556 1814
rect 550 1809 556 1810
rect 638 1814 644 1815
rect 638 1810 639 1814
rect 643 1810 644 1814
rect 638 1809 644 1810
rect 726 1814 732 1815
rect 726 1810 727 1814
rect 731 1810 732 1814
rect 726 1809 732 1810
rect 806 1814 812 1815
rect 806 1810 807 1814
rect 811 1810 812 1814
rect 806 1809 812 1810
rect 886 1814 892 1815
rect 886 1810 887 1814
rect 891 1810 892 1814
rect 886 1809 892 1810
rect 966 1814 972 1815
rect 966 1810 967 1814
rect 971 1810 972 1814
rect 966 1809 972 1810
rect 1054 1814 1060 1815
rect 1391 1814 1397 1815
rect 1439 1815 1440 1816
rect 1444 1815 1445 1819
rect 1439 1814 1445 1815
rect 1455 1819 1461 1820
rect 1455 1815 1456 1819
rect 1460 1818 1461 1819
rect 1503 1819 1509 1820
rect 1503 1818 1504 1819
rect 1460 1816 1504 1818
rect 1460 1815 1461 1816
rect 1455 1814 1461 1815
rect 1503 1815 1504 1816
rect 1508 1815 1509 1819
rect 1503 1814 1509 1815
rect 1551 1819 1557 1820
rect 1551 1815 1552 1819
rect 1556 1818 1557 1819
rect 1599 1819 1605 1820
rect 1599 1818 1600 1819
rect 1556 1816 1600 1818
rect 1556 1815 1557 1816
rect 1551 1814 1557 1815
rect 1599 1815 1600 1816
rect 1604 1815 1605 1819
rect 1599 1814 1605 1815
rect 1642 1819 1653 1820
rect 1642 1815 1643 1819
rect 1647 1815 1648 1819
rect 1652 1815 1653 1819
rect 1642 1814 1653 1815
rect 1735 1819 1741 1820
rect 1735 1815 1736 1819
rect 1740 1818 1741 1819
rect 1782 1819 1788 1820
rect 1782 1818 1783 1819
rect 1740 1816 1783 1818
rect 1740 1815 1741 1816
rect 1735 1814 1741 1815
rect 1782 1815 1783 1816
rect 1787 1815 1788 1819
rect 1782 1814 1788 1815
rect 1823 1819 1832 1820
rect 1823 1815 1824 1819
rect 1831 1815 1832 1819
rect 1823 1814 1832 1815
rect 1910 1819 1917 1820
rect 1910 1815 1911 1819
rect 1916 1815 1917 1819
rect 1910 1814 1917 1815
rect 1998 1819 2005 1820
rect 1998 1815 1999 1819
rect 2004 1815 2005 1819
rect 1998 1814 2005 1815
rect 2082 1819 2093 1820
rect 2082 1815 2083 1819
rect 2087 1815 2088 1819
rect 2092 1815 2093 1819
rect 2082 1814 2093 1815
rect 2174 1819 2181 1820
rect 2174 1815 2175 1819
rect 2180 1815 2181 1819
rect 2174 1814 2181 1815
rect 1054 1810 1055 1814
rect 1059 1810 1060 1814
rect 1054 1809 1060 1810
rect 135 1807 141 1808
rect 135 1803 136 1807
rect 140 1806 141 1807
rect 166 1807 172 1808
rect 166 1806 167 1807
rect 140 1804 167 1806
rect 140 1803 141 1804
rect 135 1802 141 1803
rect 166 1803 167 1804
rect 171 1803 172 1807
rect 166 1802 172 1803
rect 190 1807 197 1808
rect 190 1803 191 1807
rect 196 1803 197 1807
rect 190 1802 197 1803
rect 254 1807 261 1808
rect 254 1803 255 1807
rect 260 1803 261 1807
rect 254 1802 261 1803
rect 342 1807 349 1808
rect 342 1803 343 1807
rect 348 1803 349 1807
rect 342 1802 349 1803
rect 430 1807 437 1808
rect 430 1803 431 1807
rect 436 1803 437 1807
rect 430 1802 437 1803
rect 526 1807 533 1808
rect 526 1803 527 1807
rect 532 1803 533 1807
rect 526 1802 533 1803
rect 615 1807 621 1808
rect 615 1803 616 1807
rect 620 1806 621 1807
rect 630 1807 636 1808
rect 630 1806 631 1807
rect 620 1804 631 1806
rect 620 1803 621 1804
rect 615 1802 621 1803
rect 630 1803 631 1804
rect 635 1803 636 1807
rect 630 1802 636 1803
rect 702 1807 709 1808
rect 702 1803 703 1807
rect 708 1803 709 1807
rect 702 1802 709 1803
rect 782 1807 789 1808
rect 782 1803 783 1807
rect 788 1803 789 1807
rect 782 1802 789 1803
rect 862 1807 869 1808
rect 862 1803 863 1807
rect 868 1803 869 1807
rect 862 1802 869 1803
rect 943 1807 949 1808
rect 943 1803 944 1807
rect 948 1806 949 1807
rect 958 1807 964 1808
rect 958 1806 959 1807
rect 948 1804 959 1806
rect 948 1803 949 1804
rect 943 1802 949 1803
rect 958 1803 959 1804
rect 963 1803 964 1807
rect 958 1802 964 1803
rect 1030 1807 1037 1808
rect 1030 1803 1031 1807
rect 1036 1803 1037 1807
rect 1030 1802 1037 1803
rect 1391 1807 1397 1808
rect 1391 1803 1392 1807
rect 1396 1806 1397 1807
rect 1406 1807 1412 1808
rect 1406 1806 1407 1807
rect 1396 1804 1407 1806
rect 1396 1803 1397 1804
rect 1391 1802 1397 1803
rect 1406 1803 1407 1804
rect 1411 1803 1412 1807
rect 1434 1807 1440 1808
rect 1434 1803 1435 1807
rect 1439 1806 1440 1807
rect 1487 1807 1493 1808
rect 1487 1806 1488 1807
rect 1439 1804 1488 1806
rect 1439 1803 1440 1804
rect 1406 1802 1412 1803
rect 1414 1802 1420 1803
rect 1434 1802 1440 1803
rect 1487 1803 1488 1804
rect 1492 1803 1493 1807
rect 1530 1807 1536 1808
rect 1530 1803 1531 1807
rect 1535 1806 1536 1807
rect 1599 1807 1605 1808
rect 1599 1806 1600 1807
rect 1535 1804 1600 1806
rect 1535 1803 1536 1804
rect 1487 1802 1493 1803
rect 1510 1802 1516 1803
rect 1530 1802 1536 1803
rect 1599 1803 1600 1804
rect 1604 1803 1605 1807
rect 1711 1807 1720 1808
rect 1711 1803 1712 1807
rect 1719 1803 1720 1807
rect 1759 1807 1765 1808
rect 1759 1803 1760 1807
rect 1764 1806 1765 1807
rect 1815 1807 1821 1808
rect 1815 1806 1816 1807
rect 1764 1804 1816 1806
rect 1764 1803 1765 1804
rect 1599 1802 1605 1803
rect 1622 1802 1628 1803
rect 1711 1802 1720 1803
rect 1734 1802 1740 1803
rect 1759 1802 1765 1803
rect 1815 1803 1816 1804
rect 1820 1803 1821 1807
rect 1926 1807 1933 1808
rect 1926 1803 1927 1807
rect 1932 1803 1933 1807
rect 1970 1807 1976 1808
rect 1970 1803 1971 1807
rect 1975 1806 1976 1807
rect 2039 1807 2045 1808
rect 2039 1806 2040 1807
rect 1975 1804 2040 1806
rect 1975 1803 1976 1804
rect 1815 1802 1821 1803
rect 1838 1802 1844 1803
rect 1926 1802 1933 1803
rect 1950 1802 1956 1803
rect 1970 1802 1976 1803
rect 2039 1803 2040 1804
rect 2044 1803 2045 1807
rect 2154 1807 2165 1808
rect 2154 1803 2155 1807
rect 2159 1803 2160 1807
rect 2164 1803 2165 1807
rect 2234 1807 2240 1808
rect 2234 1803 2235 1807
rect 2239 1806 2240 1807
rect 2279 1807 2285 1808
rect 2279 1806 2280 1807
rect 2239 1804 2280 1806
rect 2239 1803 2240 1804
rect 2039 1802 2045 1803
rect 2062 1802 2068 1803
rect 2154 1802 2165 1803
rect 2182 1802 2188 1803
rect 2234 1802 2240 1803
rect 2279 1803 2280 1804
rect 2284 1803 2285 1807
rect 2322 1807 2328 1808
rect 2322 1803 2323 1807
rect 2327 1806 2328 1807
rect 2407 1807 2413 1808
rect 2407 1806 2408 1807
rect 2327 1804 2408 1806
rect 2327 1803 2328 1804
rect 2279 1802 2285 1803
rect 2302 1802 2308 1803
rect 2322 1802 2328 1803
rect 2407 1803 2408 1804
rect 2412 1803 2413 1807
rect 2519 1807 2525 1808
rect 2519 1803 2520 1807
rect 2524 1806 2525 1807
rect 2534 1807 2540 1808
rect 2534 1806 2535 1807
rect 2524 1804 2535 1806
rect 2524 1803 2525 1804
rect 2407 1802 2413 1803
rect 2430 1802 2436 1803
rect 2519 1802 2525 1803
rect 2534 1803 2535 1804
rect 2539 1803 2540 1807
rect 2534 1802 2540 1803
rect 2542 1802 2548 1803
rect 558 1799 564 1800
rect 558 1798 559 1799
rect 224 1796 559 1798
rect 207 1791 213 1792
rect 207 1787 208 1791
rect 212 1790 213 1791
rect 224 1790 226 1796
rect 558 1795 559 1796
rect 563 1795 564 1799
rect 1414 1798 1415 1802
rect 1419 1798 1420 1802
rect 1414 1797 1420 1798
rect 1510 1798 1511 1802
rect 1515 1798 1516 1802
rect 1510 1797 1516 1798
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1734 1798 1735 1802
rect 1739 1798 1740 1802
rect 1734 1797 1740 1798
rect 1838 1798 1839 1802
rect 1843 1798 1844 1802
rect 1838 1797 1844 1798
rect 1950 1798 1951 1802
rect 1955 1798 1956 1802
rect 1950 1797 1956 1798
rect 2062 1798 2063 1802
rect 2067 1798 2068 1802
rect 2062 1797 2068 1798
rect 2182 1798 2183 1802
rect 2187 1798 2188 1802
rect 2182 1797 2188 1798
rect 2302 1798 2303 1802
rect 2307 1798 2308 1802
rect 2302 1797 2308 1798
rect 2430 1798 2431 1802
rect 2435 1798 2436 1802
rect 2430 1797 2436 1798
rect 2542 1798 2543 1802
rect 2547 1798 2548 1802
rect 2542 1797 2548 1798
rect 558 1794 564 1795
rect 942 1795 948 1796
rect 212 1788 226 1790
rect 250 1791 256 1792
rect 212 1787 213 1788
rect 250 1787 251 1791
rect 255 1790 256 1791
rect 271 1791 277 1792
rect 271 1790 272 1791
rect 255 1788 272 1790
rect 255 1787 256 1788
rect 207 1786 213 1787
rect 230 1786 236 1787
rect 250 1786 256 1787
rect 271 1787 272 1788
rect 276 1787 277 1791
rect 314 1791 320 1792
rect 314 1787 315 1791
rect 319 1790 320 1791
rect 343 1791 349 1792
rect 343 1790 344 1791
rect 319 1788 344 1790
rect 319 1787 320 1788
rect 271 1786 277 1787
rect 294 1786 300 1787
rect 314 1786 320 1787
rect 343 1787 344 1788
rect 348 1787 349 1791
rect 386 1791 392 1792
rect 386 1787 387 1791
rect 391 1790 392 1791
rect 423 1791 429 1792
rect 423 1790 424 1791
rect 391 1788 424 1790
rect 391 1787 392 1788
rect 343 1786 349 1787
rect 366 1786 372 1787
rect 386 1786 392 1787
rect 423 1787 424 1788
rect 428 1787 429 1791
rect 466 1791 472 1792
rect 466 1787 467 1791
rect 471 1790 472 1791
rect 511 1791 517 1792
rect 511 1790 512 1791
rect 471 1788 512 1790
rect 471 1787 472 1788
rect 423 1786 429 1787
rect 446 1786 452 1787
rect 466 1786 472 1787
rect 511 1787 512 1788
rect 516 1787 517 1791
rect 598 1791 605 1792
rect 598 1787 599 1791
rect 604 1787 605 1791
rect 679 1791 685 1792
rect 679 1787 680 1791
rect 684 1790 685 1791
rect 687 1791 693 1792
rect 687 1790 688 1791
rect 684 1788 688 1790
rect 684 1787 685 1788
rect 511 1786 517 1787
rect 534 1786 540 1787
rect 598 1786 605 1787
rect 622 1786 628 1787
rect 679 1786 685 1787
rect 687 1787 688 1788
rect 692 1787 693 1791
rect 767 1791 773 1792
rect 767 1790 768 1791
rect 728 1788 768 1790
rect 726 1787 732 1788
rect 687 1786 693 1787
rect 710 1786 716 1787
rect 230 1782 231 1786
rect 235 1782 236 1786
rect 230 1781 236 1782
rect 294 1782 295 1786
rect 299 1782 300 1786
rect 294 1781 300 1782
rect 366 1782 367 1786
rect 371 1782 372 1786
rect 366 1781 372 1782
rect 446 1782 447 1786
rect 451 1782 452 1786
rect 446 1781 452 1782
rect 534 1782 535 1786
rect 539 1782 540 1786
rect 534 1781 540 1782
rect 622 1782 623 1786
rect 627 1782 628 1786
rect 622 1781 628 1782
rect 710 1782 711 1786
rect 715 1782 716 1786
rect 726 1783 727 1787
rect 731 1783 732 1787
rect 767 1787 768 1788
rect 772 1787 773 1791
rect 847 1791 853 1792
rect 847 1787 848 1791
rect 852 1790 853 1791
rect 862 1791 868 1792
rect 862 1790 863 1791
rect 852 1788 863 1790
rect 852 1787 853 1788
rect 767 1786 773 1787
rect 790 1786 796 1787
rect 847 1786 853 1787
rect 862 1787 863 1788
rect 867 1787 868 1791
rect 910 1791 916 1792
rect 910 1787 911 1791
rect 915 1790 916 1791
rect 927 1791 933 1792
rect 927 1790 928 1791
rect 915 1788 928 1790
rect 915 1787 916 1788
rect 862 1786 868 1787
rect 870 1786 876 1787
rect 910 1786 916 1787
rect 927 1787 928 1788
rect 932 1787 933 1791
rect 942 1791 943 1795
rect 947 1794 948 1795
rect 947 1792 962 1794
rect 1366 1793 1372 1794
rect 947 1791 948 1792
rect 942 1790 948 1791
rect 960 1790 962 1792
rect 1007 1791 1013 1792
rect 1007 1790 1008 1791
rect 960 1788 1008 1790
rect 1007 1787 1008 1788
rect 1012 1787 1013 1791
rect 1055 1791 1061 1792
rect 1055 1787 1056 1791
rect 1060 1790 1061 1791
rect 1095 1791 1101 1792
rect 1095 1790 1096 1791
rect 1060 1788 1096 1790
rect 1060 1787 1061 1788
rect 927 1786 933 1787
rect 950 1786 956 1787
rect 1007 1786 1013 1787
rect 1030 1786 1036 1787
rect 1055 1786 1061 1787
rect 1095 1787 1096 1788
rect 1100 1787 1101 1791
rect 1366 1789 1367 1793
rect 1371 1789 1372 1793
rect 1366 1788 1372 1789
rect 2582 1793 2588 1794
rect 2582 1789 2583 1793
rect 2587 1789 2588 1793
rect 2582 1788 2588 1789
rect 1095 1786 1101 1787
rect 1118 1786 1124 1787
rect 726 1782 732 1783
rect 790 1782 791 1786
rect 795 1782 796 1786
rect 710 1781 716 1782
rect 790 1781 796 1782
rect 870 1782 871 1786
rect 875 1782 876 1786
rect 870 1781 876 1782
rect 950 1782 951 1786
rect 955 1782 956 1786
rect 950 1781 956 1782
rect 1030 1782 1031 1786
rect 1035 1782 1036 1786
rect 1030 1781 1036 1782
rect 1118 1782 1119 1786
rect 1123 1782 1124 1786
rect 1118 1781 1124 1782
rect 1926 1783 1932 1784
rect 1926 1779 1927 1783
rect 1931 1782 1932 1783
rect 1931 1780 2442 1782
rect 1931 1779 1932 1780
rect 1926 1778 1932 1779
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 1326 1777 1332 1778
rect 1326 1773 1327 1777
rect 1331 1773 1332 1777
rect 1326 1772 1332 1773
rect 1366 1776 1372 1777
rect 1366 1772 1367 1776
rect 1371 1772 1372 1776
rect 1366 1771 1372 1772
rect 1398 1775 1404 1776
rect 1398 1771 1399 1775
rect 1403 1771 1404 1775
rect 1494 1775 1500 1776
rect 1398 1770 1404 1771
rect 1431 1771 1440 1772
rect 598 1767 604 1768
rect 598 1763 599 1767
rect 603 1766 604 1767
rect 1431 1767 1432 1771
rect 1439 1767 1440 1771
rect 1494 1771 1495 1775
rect 1499 1771 1500 1775
rect 1606 1775 1612 1776
rect 1494 1770 1500 1771
rect 1527 1771 1536 1772
rect 1431 1766 1440 1767
rect 1527 1767 1528 1771
rect 1535 1767 1536 1771
rect 1606 1771 1607 1775
rect 1611 1771 1612 1775
rect 1718 1775 1724 1776
rect 1606 1770 1612 1771
rect 1639 1771 1648 1772
rect 1527 1766 1536 1767
rect 1639 1767 1640 1771
rect 1647 1767 1648 1771
rect 1718 1771 1719 1775
rect 1723 1771 1724 1775
rect 1822 1775 1828 1776
rect 1718 1770 1724 1771
rect 1751 1771 1757 1772
rect 1639 1766 1648 1767
rect 1751 1767 1752 1771
rect 1756 1770 1757 1771
rect 1759 1771 1765 1772
rect 1759 1770 1760 1771
rect 1756 1768 1760 1770
rect 1756 1767 1757 1768
rect 1751 1766 1757 1767
rect 1759 1767 1760 1768
rect 1764 1767 1765 1771
rect 1822 1771 1823 1775
rect 1827 1771 1828 1775
rect 1934 1775 1940 1776
rect 1822 1770 1828 1771
rect 1855 1771 1861 1772
rect 1759 1766 1765 1767
rect 1855 1767 1856 1771
rect 1860 1770 1861 1771
rect 1918 1771 1924 1772
rect 1918 1770 1919 1771
rect 1860 1768 1919 1770
rect 1860 1767 1861 1768
rect 1855 1766 1861 1767
rect 1918 1767 1919 1768
rect 1923 1767 1924 1771
rect 1934 1771 1935 1775
rect 1939 1771 1940 1775
rect 2046 1775 2052 1776
rect 1934 1770 1940 1771
rect 1967 1771 1976 1772
rect 1918 1766 1924 1767
rect 1967 1767 1968 1771
rect 1975 1767 1976 1771
rect 2046 1771 2047 1775
rect 2051 1771 2052 1775
rect 2166 1775 2172 1776
rect 2046 1770 2052 1771
rect 2079 1771 2088 1772
rect 1967 1766 1976 1767
rect 2079 1767 2080 1771
rect 2087 1767 2088 1771
rect 2166 1771 2167 1775
rect 2171 1771 2172 1775
rect 2286 1775 2292 1776
rect 2166 1770 2172 1771
rect 2199 1771 2205 1772
rect 2079 1766 2088 1767
rect 2199 1767 2200 1771
rect 2204 1770 2205 1771
rect 2234 1771 2240 1772
rect 2234 1770 2235 1771
rect 2204 1768 2235 1770
rect 2204 1767 2205 1768
rect 2199 1766 2205 1767
rect 2234 1767 2235 1768
rect 2239 1767 2240 1771
rect 2286 1771 2287 1775
rect 2291 1771 2292 1775
rect 2414 1775 2420 1776
rect 2286 1770 2292 1771
rect 2319 1771 2328 1772
rect 2234 1766 2240 1767
rect 2319 1767 2320 1771
rect 2327 1767 2328 1771
rect 2414 1771 2415 1775
rect 2419 1771 2420 1775
rect 2414 1770 2420 1771
rect 2440 1770 2442 1780
rect 2582 1776 2588 1777
rect 2526 1775 2532 1776
rect 2447 1771 2453 1772
rect 2447 1770 2448 1771
rect 2440 1768 2448 1770
rect 2319 1766 2328 1767
rect 2447 1767 2448 1768
rect 2452 1767 2453 1771
rect 2526 1771 2527 1775
rect 2531 1771 2532 1775
rect 2582 1772 2583 1776
rect 2587 1772 2588 1776
rect 2526 1770 2532 1771
rect 2559 1771 2565 1772
rect 2582 1771 2588 1772
rect 2447 1766 2453 1767
rect 2470 1767 2476 1768
rect 603 1764 802 1766
rect 603 1763 604 1764
rect 598 1762 604 1763
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 278 1759 284 1760
rect 214 1754 220 1755
rect 247 1755 256 1756
rect 247 1751 248 1755
rect 255 1751 256 1755
rect 278 1755 279 1759
rect 283 1755 284 1759
rect 350 1759 356 1760
rect 278 1754 284 1755
rect 311 1755 320 1756
rect 247 1750 256 1751
rect 311 1751 312 1755
rect 319 1751 320 1755
rect 350 1755 351 1759
rect 355 1755 356 1759
rect 430 1759 436 1760
rect 350 1754 356 1755
rect 383 1755 392 1756
rect 311 1750 320 1751
rect 383 1751 384 1755
rect 391 1751 392 1755
rect 430 1755 431 1759
rect 435 1755 436 1759
rect 518 1759 524 1760
rect 430 1754 436 1755
rect 463 1755 472 1756
rect 383 1750 392 1751
rect 463 1751 464 1755
rect 471 1751 472 1755
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 606 1759 612 1760
rect 518 1754 524 1755
rect 551 1755 557 1756
rect 551 1754 552 1755
rect 463 1750 472 1751
rect 528 1752 552 1754
rect 358 1747 364 1748
rect 358 1743 359 1747
rect 363 1746 364 1747
rect 528 1746 530 1752
rect 551 1751 552 1752
rect 556 1751 557 1755
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 694 1759 700 1760
rect 606 1754 612 1755
rect 630 1755 636 1756
rect 551 1750 557 1751
rect 630 1751 631 1755
rect 635 1754 636 1755
rect 639 1755 645 1756
rect 639 1754 640 1755
rect 635 1752 640 1754
rect 635 1751 636 1752
rect 630 1750 636 1751
rect 639 1751 640 1752
rect 644 1751 645 1755
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 774 1759 780 1760
rect 694 1754 700 1755
rect 726 1755 733 1756
rect 639 1750 645 1751
rect 726 1751 727 1755
rect 732 1751 733 1755
rect 774 1755 775 1759
rect 779 1755 780 1759
rect 774 1754 780 1755
rect 800 1754 802 1764
rect 2470 1763 2471 1767
rect 2475 1766 2476 1767
rect 2559 1767 2560 1771
rect 2564 1767 2565 1771
rect 2559 1766 2565 1767
rect 2475 1764 2563 1766
rect 2475 1763 2476 1764
rect 2470 1762 2476 1763
rect 1326 1760 1332 1761
rect 854 1759 860 1760
rect 807 1755 813 1756
rect 807 1754 808 1755
rect 800 1752 808 1754
rect 726 1750 733 1751
rect 807 1751 808 1752
rect 812 1751 813 1755
rect 854 1755 855 1759
rect 859 1755 860 1759
rect 910 1759 916 1760
rect 910 1758 911 1759
rect 854 1754 860 1755
rect 887 1757 911 1758
rect 887 1753 888 1757
rect 892 1756 911 1757
rect 892 1753 893 1756
rect 910 1755 911 1756
rect 915 1755 916 1759
rect 910 1754 916 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 1014 1759 1020 1760
rect 934 1754 940 1755
rect 958 1755 964 1756
rect 887 1752 893 1753
rect 807 1750 813 1751
rect 958 1751 959 1755
rect 963 1754 964 1755
rect 967 1755 973 1756
rect 967 1754 968 1755
rect 963 1752 968 1754
rect 963 1751 964 1752
rect 958 1750 964 1751
rect 967 1751 968 1752
rect 972 1751 973 1755
rect 1014 1755 1015 1759
rect 1019 1755 1020 1759
rect 1102 1759 1108 1760
rect 1014 1754 1020 1755
rect 1047 1755 1053 1756
rect 967 1750 973 1751
rect 1047 1751 1048 1755
rect 1052 1754 1053 1755
rect 1055 1755 1061 1756
rect 1055 1754 1056 1755
rect 1052 1752 1056 1754
rect 1052 1751 1053 1752
rect 1047 1750 1053 1751
rect 1055 1751 1056 1752
rect 1060 1751 1061 1755
rect 1102 1755 1103 1759
rect 1107 1755 1108 1759
rect 1326 1756 1327 1760
rect 1331 1756 1332 1760
rect 1102 1754 1108 1755
rect 1135 1755 1141 1756
rect 1326 1755 1332 1756
rect 1135 1754 1136 1755
rect 1112 1752 1136 1754
rect 1055 1750 1061 1751
rect 1063 1751 1069 1752
rect 1063 1747 1064 1751
rect 1068 1750 1069 1751
rect 1112 1750 1114 1752
rect 1135 1751 1136 1752
rect 1140 1751 1141 1755
rect 1135 1750 1141 1751
rect 1068 1748 1114 1750
rect 1068 1747 1069 1748
rect 1063 1746 1069 1747
rect 1406 1747 1412 1748
rect 363 1744 530 1746
rect 363 1743 364 1744
rect 358 1742 364 1743
rect 1406 1743 1407 1747
rect 1411 1746 1412 1747
rect 1479 1747 1485 1748
rect 1411 1744 1466 1746
rect 1411 1743 1412 1744
rect 1406 1742 1412 1743
rect 1464 1742 1466 1744
rect 1471 1743 1477 1744
rect 1471 1742 1472 1743
rect 1438 1741 1444 1742
rect 1366 1740 1372 1741
rect 1366 1736 1367 1740
rect 1371 1736 1372 1740
rect 1438 1737 1439 1741
rect 1443 1737 1444 1741
rect 1464 1740 1472 1742
rect 1471 1739 1472 1740
rect 1476 1739 1477 1743
rect 1479 1743 1480 1747
rect 1484 1746 1485 1747
rect 1559 1747 1565 1748
rect 1484 1744 1546 1746
rect 1484 1743 1485 1744
rect 1479 1742 1485 1743
rect 1544 1742 1546 1744
rect 1551 1743 1557 1744
rect 1551 1742 1552 1743
rect 1471 1738 1477 1739
rect 1518 1741 1524 1742
rect 1438 1736 1444 1737
rect 1518 1737 1519 1741
rect 1523 1737 1524 1741
rect 1544 1740 1552 1742
rect 1551 1739 1552 1740
rect 1556 1739 1557 1743
rect 1559 1743 1560 1747
rect 1564 1746 1565 1747
rect 1655 1747 1661 1748
rect 1564 1744 1642 1746
rect 1564 1743 1565 1744
rect 1559 1742 1565 1743
rect 1640 1742 1642 1744
rect 1647 1743 1653 1744
rect 1647 1742 1648 1743
rect 1551 1738 1557 1739
rect 1614 1741 1620 1742
rect 1518 1736 1524 1737
rect 1614 1737 1615 1741
rect 1619 1737 1620 1741
rect 1640 1740 1648 1742
rect 1647 1739 1648 1740
rect 1652 1739 1653 1743
rect 1655 1743 1656 1747
rect 1660 1746 1661 1747
rect 1774 1747 1780 1748
rect 1660 1744 1746 1746
rect 1660 1743 1661 1744
rect 1655 1742 1661 1743
rect 1744 1742 1746 1744
rect 1751 1743 1757 1744
rect 1751 1742 1752 1743
rect 1647 1738 1653 1739
rect 1718 1741 1724 1742
rect 1614 1736 1620 1737
rect 1718 1737 1719 1741
rect 1723 1737 1724 1741
rect 1744 1740 1752 1742
rect 1751 1739 1752 1740
rect 1756 1739 1757 1743
rect 1774 1743 1775 1747
rect 1779 1746 1780 1747
rect 1863 1747 1869 1748
rect 1779 1744 1850 1746
rect 1779 1743 1780 1744
rect 1774 1742 1780 1743
rect 1848 1742 1850 1744
rect 1855 1743 1861 1744
rect 1855 1742 1856 1743
rect 1751 1738 1757 1739
rect 1822 1741 1828 1742
rect 1718 1736 1724 1737
rect 1822 1737 1823 1741
rect 1827 1737 1828 1741
rect 1848 1740 1856 1742
rect 1855 1739 1856 1740
rect 1860 1739 1861 1743
rect 1863 1743 1864 1747
rect 1868 1746 1869 1747
rect 2534 1747 2540 1748
rect 1868 1744 1954 1746
rect 1868 1743 1869 1744
rect 1863 1742 1869 1743
rect 1952 1742 1954 1744
rect 1959 1743 1965 1744
rect 1959 1742 1960 1743
rect 1855 1738 1861 1739
rect 1926 1741 1932 1742
rect 1822 1736 1828 1737
rect 1926 1737 1927 1741
rect 1931 1737 1932 1741
rect 1952 1740 1960 1742
rect 1959 1739 1960 1740
rect 1964 1739 1965 1743
rect 2055 1743 2061 1744
rect 1959 1738 1965 1739
rect 2022 1741 2028 1742
rect 1926 1736 1932 1737
rect 2022 1737 2023 1741
rect 2027 1737 2028 1741
rect 2055 1739 2056 1743
rect 2060 1742 2061 1743
rect 2110 1743 2116 1744
rect 2110 1742 2111 1743
rect 2060 1740 2111 1742
rect 2060 1739 2061 1740
rect 2055 1738 2061 1739
rect 2110 1739 2111 1740
rect 2115 1739 2116 1743
rect 2151 1743 2160 1744
rect 2110 1738 2116 1739
rect 2118 1741 2124 1742
rect 2022 1736 2028 1737
rect 2118 1737 2119 1741
rect 2123 1737 2124 1741
rect 2151 1739 2152 1743
rect 2159 1739 2160 1743
rect 2239 1743 2245 1744
rect 2151 1738 2160 1739
rect 2206 1741 2212 1742
rect 2118 1736 2124 1737
rect 2206 1737 2207 1741
rect 2211 1737 2212 1741
rect 2239 1739 2240 1743
rect 2244 1742 2245 1743
rect 2278 1743 2284 1744
rect 2278 1742 2279 1743
rect 2244 1740 2279 1742
rect 2244 1739 2245 1740
rect 2239 1738 2245 1739
rect 2278 1739 2279 1740
rect 2283 1739 2284 1743
rect 2319 1743 2325 1744
rect 2278 1738 2284 1739
rect 2286 1741 2292 1742
rect 2206 1736 2212 1737
rect 2286 1737 2287 1741
rect 2291 1737 2292 1741
rect 2319 1739 2320 1743
rect 2324 1742 2325 1743
rect 2366 1743 2372 1744
rect 2366 1742 2367 1743
rect 2324 1740 2367 1742
rect 2324 1739 2325 1740
rect 2319 1738 2325 1739
rect 2366 1739 2367 1740
rect 2371 1739 2372 1743
rect 2398 1743 2404 1744
rect 2366 1738 2372 1739
rect 2374 1741 2380 1742
rect 2286 1736 2292 1737
rect 2374 1737 2375 1741
rect 2379 1737 2380 1741
rect 2398 1739 2399 1743
rect 2403 1742 2404 1743
rect 2407 1743 2413 1744
rect 2407 1742 2408 1743
rect 2403 1740 2408 1742
rect 2403 1739 2404 1740
rect 2398 1738 2404 1739
rect 2407 1739 2408 1740
rect 2412 1739 2413 1743
rect 2494 1743 2501 1744
rect 2407 1738 2413 1739
rect 2462 1741 2468 1742
rect 2374 1736 2380 1737
rect 2462 1737 2463 1741
rect 2467 1737 2468 1741
rect 2494 1739 2495 1743
rect 2500 1739 2501 1743
rect 2534 1743 2535 1747
rect 2539 1746 2540 1747
rect 2539 1744 2563 1746
rect 2539 1743 2540 1744
rect 2534 1742 2540 1743
rect 2559 1743 2565 1744
rect 2494 1738 2501 1739
rect 2526 1741 2532 1742
rect 2462 1736 2468 1737
rect 2526 1737 2527 1741
rect 2531 1737 2532 1741
rect 2559 1739 2560 1743
rect 2564 1739 2565 1743
rect 2559 1738 2565 1739
rect 2582 1740 2588 1741
rect 2526 1736 2532 1737
rect 2582 1736 2583 1740
rect 2587 1736 2588 1740
rect 1366 1735 1372 1736
rect 2582 1735 2588 1736
rect 862 1731 868 1732
rect 687 1727 693 1728
rect 383 1723 389 1724
rect 350 1721 356 1722
rect 110 1720 116 1721
rect 110 1716 111 1720
rect 115 1716 116 1720
rect 350 1717 351 1721
rect 355 1717 356 1721
rect 383 1719 384 1723
rect 388 1722 389 1723
rect 398 1723 404 1724
rect 398 1722 399 1723
rect 388 1720 399 1722
rect 388 1719 389 1720
rect 383 1718 389 1719
rect 398 1719 399 1720
rect 403 1719 404 1723
rect 439 1723 445 1724
rect 398 1718 404 1719
rect 406 1721 412 1722
rect 350 1716 356 1717
rect 406 1717 407 1721
rect 411 1717 412 1721
rect 439 1719 440 1723
rect 444 1722 445 1723
rect 462 1723 468 1724
rect 462 1722 463 1723
rect 444 1720 463 1722
rect 444 1719 445 1720
rect 439 1718 445 1719
rect 462 1719 463 1720
rect 467 1719 468 1723
rect 503 1723 509 1724
rect 462 1718 468 1719
rect 470 1721 476 1722
rect 406 1716 412 1717
rect 470 1717 471 1721
rect 475 1717 476 1721
rect 503 1719 504 1723
rect 508 1722 509 1723
rect 542 1723 548 1724
rect 542 1722 543 1723
rect 508 1720 543 1722
rect 508 1719 509 1720
rect 503 1718 509 1719
rect 542 1719 543 1720
rect 547 1719 548 1723
rect 582 1723 589 1724
rect 542 1718 548 1719
rect 550 1721 556 1722
rect 470 1716 476 1717
rect 550 1717 551 1721
rect 555 1717 556 1721
rect 582 1719 583 1723
rect 588 1719 589 1723
rect 671 1723 677 1724
rect 582 1718 589 1719
rect 638 1721 644 1722
rect 550 1716 556 1717
rect 638 1717 639 1721
rect 643 1717 644 1721
rect 671 1719 672 1723
rect 676 1722 677 1723
rect 679 1723 685 1724
rect 679 1722 680 1723
rect 676 1720 680 1722
rect 676 1719 677 1720
rect 671 1718 677 1719
rect 679 1719 680 1720
rect 684 1719 685 1723
rect 687 1723 688 1727
rect 692 1726 693 1727
rect 767 1727 773 1728
rect 692 1724 754 1726
rect 692 1723 693 1724
rect 687 1722 693 1723
rect 752 1722 754 1724
rect 759 1723 765 1724
rect 759 1722 760 1723
rect 679 1718 685 1719
rect 726 1721 732 1722
rect 638 1716 644 1717
rect 726 1717 727 1721
rect 731 1717 732 1721
rect 752 1720 760 1722
rect 759 1719 760 1720
rect 764 1719 765 1723
rect 767 1723 768 1727
rect 772 1726 773 1727
rect 862 1727 863 1731
rect 867 1727 868 1731
rect 862 1726 868 1727
rect 772 1724 859 1726
rect 864 1724 946 1726
rect 772 1723 773 1724
rect 767 1722 773 1723
rect 855 1723 861 1724
rect 759 1718 765 1719
rect 822 1721 828 1722
rect 726 1716 732 1717
rect 822 1717 823 1721
rect 827 1717 828 1721
rect 855 1719 856 1723
rect 860 1719 861 1723
rect 944 1722 946 1724
rect 951 1723 957 1724
rect 951 1722 952 1723
rect 855 1718 861 1719
rect 918 1721 924 1722
rect 822 1716 828 1717
rect 918 1717 919 1721
rect 923 1717 924 1721
rect 944 1720 952 1722
rect 951 1719 952 1720
rect 956 1719 957 1723
rect 1047 1723 1053 1724
rect 951 1718 957 1719
rect 1014 1721 1020 1722
rect 918 1716 924 1717
rect 1014 1717 1015 1721
rect 1019 1717 1020 1721
rect 1047 1719 1048 1723
rect 1052 1722 1053 1723
rect 1102 1723 1108 1724
rect 1102 1722 1103 1723
rect 1052 1720 1103 1722
rect 1052 1719 1053 1720
rect 1047 1718 1053 1719
rect 1102 1719 1103 1720
rect 1107 1719 1108 1723
rect 1143 1723 1149 1724
rect 1102 1718 1108 1719
rect 1110 1721 1116 1722
rect 1014 1716 1020 1717
rect 1110 1717 1111 1721
rect 1115 1717 1116 1721
rect 1143 1719 1144 1723
rect 1148 1722 1149 1723
rect 1198 1723 1204 1724
rect 1198 1722 1199 1723
rect 1148 1720 1199 1722
rect 1148 1719 1149 1720
rect 1143 1718 1149 1719
rect 1198 1719 1199 1720
rect 1203 1719 1204 1723
rect 1230 1723 1236 1724
rect 1198 1718 1204 1719
rect 1206 1721 1212 1722
rect 1110 1716 1116 1717
rect 1206 1717 1207 1721
rect 1211 1717 1212 1721
rect 1230 1719 1231 1723
rect 1235 1722 1236 1723
rect 1239 1723 1245 1724
rect 1239 1722 1240 1723
rect 1235 1720 1240 1722
rect 1235 1719 1236 1720
rect 1230 1718 1236 1719
rect 1239 1719 1240 1720
rect 1244 1719 1245 1723
rect 1366 1723 1372 1724
rect 1239 1718 1245 1719
rect 1326 1720 1332 1721
rect 1206 1716 1212 1717
rect 1326 1716 1327 1720
rect 1331 1716 1332 1720
rect 1366 1719 1367 1723
rect 1371 1719 1372 1723
rect 1366 1718 1372 1719
rect 2582 1723 2588 1724
rect 2582 1719 2583 1723
rect 2587 1719 2588 1723
rect 2582 1718 2588 1719
rect 110 1715 116 1716
rect 1326 1715 1332 1716
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1534 1714 1540 1715
rect 1534 1710 1535 1714
rect 1539 1710 1540 1714
rect 1534 1709 1540 1710
rect 1630 1714 1636 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 1734 1714 1740 1715
rect 1734 1710 1735 1714
rect 1739 1710 1740 1714
rect 1734 1709 1740 1710
rect 1838 1714 1844 1715
rect 1838 1710 1839 1714
rect 1843 1710 1844 1714
rect 1838 1709 1844 1710
rect 1942 1714 1948 1715
rect 1942 1710 1943 1714
rect 1947 1710 1948 1714
rect 1942 1709 1948 1710
rect 2038 1714 2044 1715
rect 2038 1710 2039 1714
rect 2043 1710 2044 1714
rect 2038 1709 2044 1710
rect 2134 1714 2140 1715
rect 2134 1710 2135 1714
rect 2139 1710 2140 1714
rect 2134 1709 2140 1710
rect 2222 1714 2228 1715
rect 2222 1710 2223 1714
rect 2227 1710 2228 1714
rect 2222 1709 2228 1710
rect 2302 1714 2308 1715
rect 2302 1710 2303 1714
rect 2307 1710 2308 1714
rect 2302 1709 2308 1710
rect 2390 1714 2396 1715
rect 2390 1710 2391 1714
rect 2395 1710 2396 1714
rect 2390 1709 2396 1710
rect 2478 1714 2484 1715
rect 2478 1710 2479 1714
rect 2483 1710 2484 1714
rect 2478 1709 2484 1710
rect 2542 1714 2548 1715
rect 2542 1710 2543 1714
rect 2547 1710 2548 1714
rect 2542 1709 2548 1710
rect 1431 1707 1437 1708
rect 110 1703 116 1704
rect 110 1699 111 1703
rect 115 1699 116 1703
rect 110 1698 116 1699
rect 1326 1703 1332 1704
rect 1326 1699 1327 1703
rect 1331 1699 1332 1703
rect 1431 1703 1432 1707
rect 1436 1706 1437 1707
rect 1479 1707 1485 1708
rect 1479 1706 1480 1707
rect 1436 1704 1480 1706
rect 1436 1703 1437 1704
rect 1431 1702 1437 1703
rect 1479 1703 1480 1704
rect 1484 1703 1485 1707
rect 1479 1702 1485 1703
rect 1511 1707 1517 1708
rect 1511 1703 1512 1707
rect 1516 1706 1517 1707
rect 1559 1707 1565 1708
rect 1559 1706 1560 1707
rect 1516 1704 1560 1706
rect 1516 1703 1517 1704
rect 1511 1702 1517 1703
rect 1559 1703 1560 1704
rect 1564 1703 1565 1707
rect 1559 1702 1565 1703
rect 1607 1707 1613 1708
rect 1607 1703 1608 1707
rect 1612 1706 1613 1707
rect 1655 1707 1661 1708
rect 1655 1706 1656 1707
rect 1612 1704 1656 1706
rect 1612 1703 1613 1704
rect 1607 1702 1613 1703
rect 1655 1703 1656 1704
rect 1660 1703 1661 1707
rect 1655 1702 1661 1703
rect 1711 1707 1717 1708
rect 1711 1703 1712 1707
rect 1716 1706 1717 1707
rect 1722 1707 1728 1708
rect 1722 1706 1723 1707
rect 1716 1704 1723 1706
rect 1716 1703 1717 1704
rect 1711 1702 1717 1703
rect 1722 1703 1723 1704
rect 1727 1703 1728 1707
rect 1722 1702 1728 1703
rect 1815 1707 1821 1708
rect 1815 1703 1816 1707
rect 1820 1706 1821 1707
rect 1863 1707 1869 1708
rect 1863 1706 1864 1707
rect 1820 1704 1864 1706
rect 1820 1703 1821 1704
rect 1815 1702 1821 1703
rect 1863 1703 1864 1704
rect 1868 1703 1869 1707
rect 1863 1702 1869 1703
rect 1918 1707 1925 1708
rect 1918 1703 1919 1707
rect 1924 1703 1925 1707
rect 1918 1702 1925 1703
rect 2015 1707 2024 1708
rect 2015 1703 2016 1707
rect 2023 1703 2024 1707
rect 2015 1702 2024 1703
rect 2110 1707 2117 1708
rect 2110 1703 2111 1707
rect 2116 1703 2117 1707
rect 2110 1702 2117 1703
rect 2199 1707 2205 1708
rect 2199 1703 2200 1707
rect 2204 1706 2205 1707
rect 2230 1707 2236 1708
rect 2230 1706 2231 1707
rect 2204 1704 2231 1706
rect 2204 1703 2205 1704
rect 2199 1702 2205 1703
rect 2230 1703 2231 1704
rect 2235 1703 2236 1707
rect 2230 1702 2236 1703
rect 2278 1707 2285 1708
rect 2278 1703 2279 1707
rect 2284 1703 2285 1707
rect 2278 1702 2285 1703
rect 2366 1707 2373 1708
rect 2366 1703 2367 1707
rect 2372 1703 2373 1707
rect 2366 1702 2373 1703
rect 2455 1707 2461 1708
rect 2455 1703 2456 1707
rect 2460 1706 2461 1707
rect 2470 1707 2476 1708
rect 2470 1706 2471 1707
rect 2460 1704 2471 1706
rect 2460 1703 2461 1704
rect 2455 1702 2461 1703
rect 2470 1703 2471 1704
rect 2475 1703 2476 1707
rect 2470 1702 2476 1703
rect 2519 1707 2525 1708
rect 2519 1703 2520 1707
rect 2524 1706 2525 1707
rect 2558 1707 2564 1708
rect 2558 1706 2559 1707
rect 2524 1704 2559 1706
rect 2524 1703 2525 1704
rect 2519 1702 2525 1703
rect 2558 1703 2559 1704
rect 2563 1703 2564 1707
rect 2558 1702 2564 1703
rect 1326 1698 1332 1699
rect 366 1694 372 1695
rect 366 1690 367 1694
rect 371 1690 372 1694
rect 366 1689 372 1690
rect 422 1694 428 1695
rect 422 1690 423 1694
rect 427 1690 428 1694
rect 422 1689 428 1690
rect 486 1694 492 1695
rect 486 1690 487 1694
rect 491 1690 492 1694
rect 486 1689 492 1690
rect 566 1694 572 1695
rect 566 1690 567 1694
rect 571 1690 572 1694
rect 566 1689 572 1690
rect 654 1694 660 1695
rect 654 1690 655 1694
rect 659 1690 660 1694
rect 654 1689 660 1690
rect 742 1694 748 1695
rect 742 1690 743 1694
rect 747 1690 748 1694
rect 742 1689 748 1690
rect 838 1694 844 1695
rect 838 1690 839 1694
rect 843 1690 844 1694
rect 838 1689 844 1690
rect 934 1694 940 1695
rect 934 1690 935 1694
rect 939 1690 940 1694
rect 934 1689 940 1690
rect 1030 1694 1036 1695
rect 1030 1690 1031 1694
rect 1035 1690 1036 1694
rect 1030 1689 1036 1690
rect 1126 1694 1132 1695
rect 1126 1690 1127 1694
rect 1131 1690 1132 1694
rect 1126 1689 1132 1690
rect 1222 1694 1228 1695
rect 1222 1690 1223 1694
rect 1227 1690 1228 1694
rect 2294 1691 2300 1692
rect 2294 1690 2295 1691
rect 1222 1689 1228 1690
rect 2056 1688 2295 1690
rect 343 1687 349 1688
rect 343 1683 344 1687
rect 348 1686 349 1687
rect 358 1687 364 1688
rect 358 1686 359 1687
rect 348 1684 359 1686
rect 348 1683 349 1684
rect 343 1682 349 1683
rect 358 1683 359 1684
rect 363 1683 364 1687
rect 358 1682 364 1683
rect 398 1687 405 1688
rect 398 1683 399 1687
rect 404 1683 405 1687
rect 398 1682 405 1683
rect 462 1687 469 1688
rect 462 1683 463 1687
rect 468 1683 469 1687
rect 462 1682 469 1683
rect 542 1687 549 1688
rect 542 1683 543 1687
rect 548 1683 549 1687
rect 542 1682 549 1683
rect 631 1687 637 1688
rect 631 1683 632 1687
rect 636 1686 637 1687
rect 687 1687 693 1688
rect 687 1686 688 1687
rect 636 1684 688 1686
rect 636 1683 637 1684
rect 631 1682 637 1683
rect 687 1683 688 1684
rect 692 1683 693 1687
rect 687 1682 693 1683
rect 719 1687 725 1688
rect 719 1683 720 1687
rect 724 1686 725 1687
rect 767 1687 773 1688
rect 767 1686 768 1687
rect 724 1684 768 1686
rect 724 1683 725 1684
rect 719 1682 725 1683
rect 767 1683 768 1684
rect 772 1683 773 1687
rect 767 1682 773 1683
rect 815 1687 824 1688
rect 815 1683 816 1687
rect 823 1683 824 1687
rect 815 1682 824 1683
rect 911 1687 917 1688
rect 911 1683 912 1687
rect 916 1686 917 1687
rect 982 1687 988 1688
rect 982 1686 983 1687
rect 916 1684 983 1686
rect 916 1683 917 1684
rect 911 1682 917 1683
rect 982 1683 983 1684
rect 987 1683 988 1687
rect 982 1682 988 1683
rect 1007 1687 1013 1688
rect 1007 1683 1008 1687
rect 1012 1686 1013 1687
rect 1063 1687 1069 1688
rect 1063 1686 1064 1687
rect 1012 1684 1064 1686
rect 1012 1683 1013 1684
rect 1007 1682 1013 1683
rect 1063 1683 1064 1684
rect 1068 1683 1069 1687
rect 1063 1682 1069 1683
rect 1102 1687 1109 1688
rect 1102 1683 1103 1687
rect 1108 1683 1109 1687
rect 1102 1682 1109 1683
rect 1198 1687 1205 1688
rect 1198 1683 1199 1687
rect 1204 1683 1205 1687
rect 1198 1682 1205 1683
rect 1535 1683 1541 1684
rect 582 1679 588 1680
rect 582 1678 583 1679
rect 392 1676 583 1678
rect 375 1671 381 1672
rect 375 1667 376 1671
rect 380 1670 381 1671
rect 392 1670 394 1676
rect 582 1675 583 1676
rect 587 1675 588 1679
rect 1535 1679 1536 1683
rect 1540 1682 1541 1683
rect 1550 1683 1556 1684
rect 1550 1682 1551 1683
rect 1540 1680 1551 1682
rect 1540 1679 1541 1680
rect 1535 1678 1541 1679
rect 1550 1679 1551 1680
rect 1555 1679 1556 1683
rect 1578 1683 1584 1684
rect 1578 1679 1579 1683
rect 1583 1682 1584 1683
rect 1607 1683 1613 1684
rect 1607 1682 1608 1683
rect 1583 1680 1608 1682
rect 1583 1679 1584 1680
rect 1550 1678 1556 1679
rect 1558 1678 1564 1679
rect 1578 1678 1584 1679
rect 1607 1679 1608 1680
rect 1612 1679 1613 1683
rect 1650 1683 1656 1684
rect 1650 1679 1651 1683
rect 1655 1682 1656 1683
rect 1687 1683 1693 1684
rect 1687 1682 1688 1683
rect 1655 1680 1688 1682
rect 1655 1679 1656 1680
rect 1607 1678 1613 1679
rect 1630 1678 1636 1679
rect 1650 1678 1656 1679
rect 1687 1679 1688 1680
rect 1692 1679 1693 1683
rect 1774 1683 1781 1684
rect 1774 1679 1775 1683
rect 1780 1679 1781 1683
rect 1818 1683 1824 1684
rect 1818 1679 1819 1683
rect 1823 1682 1824 1683
rect 1863 1683 1869 1684
rect 1863 1682 1864 1683
rect 1823 1680 1864 1682
rect 1823 1679 1824 1680
rect 1687 1678 1693 1679
rect 1710 1678 1716 1679
rect 1774 1678 1781 1679
rect 1798 1678 1804 1679
rect 1818 1678 1824 1679
rect 1863 1679 1864 1680
rect 1868 1679 1869 1683
rect 1902 1683 1908 1684
rect 1902 1679 1903 1683
rect 1907 1682 1908 1683
rect 1951 1683 1957 1684
rect 1951 1682 1952 1683
rect 1907 1680 1952 1682
rect 1907 1679 1908 1680
rect 1863 1678 1869 1679
rect 1886 1678 1892 1679
rect 1902 1678 1908 1679
rect 1951 1679 1952 1680
rect 1956 1679 1957 1683
rect 2039 1683 2045 1684
rect 2039 1679 2040 1683
rect 2044 1682 2045 1683
rect 2056 1682 2058 1688
rect 2294 1687 2295 1688
rect 2299 1687 2300 1691
rect 2434 1691 2440 1692
rect 2434 1690 2435 1691
rect 2294 1686 2300 1687
rect 2345 1688 2435 1690
rect 2044 1680 2058 1682
rect 2082 1683 2088 1684
rect 2044 1679 2045 1680
rect 2082 1679 2083 1683
rect 2087 1682 2088 1683
rect 2119 1683 2125 1684
rect 2119 1682 2120 1683
rect 2087 1680 2120 1682
rect 2087 1679 2088 1680
rect 1951 1678 1957 1679
rect 1974 1678 1980 1679
rect 2039 1678 2045 1679
rect 2062 1678 2068 1679
rect 2082 1678 2088 1679
rect 2119 1679 2120 1680
rect 2124 1679 2125 1683
rect 2162 1683 2168 1684
rect 2162 1679 2163 1683
rect 2167 1682 2168 1683
rect 2191 1683 2197 1684
rect 2191 1682 2192 1683
rect 2167 1680 2192 1682
rect 2167 1679 2168 1680
rect 2119 1678 2125 1679
rect 2142 1678 2148 1679
rect 2162 1678 2168 1679
rect 2191 1679 2192 1680
rect 2196 1679 2197 1683
rect 2262 1683 2269 1684
rect 2262 1679 2263 1683
rect 2268 1679 2269 1683
rect 2327 1683 2333 1684
rect 2327 1679 2328 1683
rect 2332 1682 2333 1683
rect 2345 1682 2347 1688
rect 2434 1687 2435 1688
rect 2439 1687 2440 1691
rect 2434 1686 2440 1687
rect 2494 1687 2500 1688
rect 2494 1686 2495 1687
rect 2465 1684 2495 1686
rect 2332 1680 2347 1682
rect 2398 1683 2405 1684
rect 2332 1679 2333 1680
rect 2398 1679 2399 1683
rect 2404 1679 2405 1683
rect 2463 1683 2469 1684
rect 2463 1679 2464 1683
rect 2468 1679 2469 1683
rect 2494 1683 2495 1684
rect 2499 1683 2500 1687
rect 2494 1682 2500 1683
rect 2519 1683 2525 1684
rect 2519 1679 2520 1683
rect 2524 1682 2525 1683
rect 2534 1683 2540 1684
rect 2534 1682 2535 1683
rect 2524 1680 2535 1682
rect 2524 1679 2525 1680
rect 2191 1678 2197 1679
rect 2214 1678 2220 1679
rect 2262 1678 2269 1679
rect 2286 1678 2292 1679
rect 2327 1678 2333 1679
rect 2350 1678 2356 1679
rect 2398 1678 2405 1679
rect 2422 1678 2428 1679
rect 2463 1678 2469 1679
rect 2486 1678 2492 1679
rect 2519 1678 2525 1679
rect 2534 1679 2535 1680
rect 2539 1679 2540 1683
rect 2534 1678 2540 1679
rect 2542 1678 2548 1679
rect 582 1674 588 1675
rect 1230 1675 1236 1676
rect 1230 1674 1231 1675
rect 1216 1672 1231 1674
rect 380 1668 394 1670
rect 423 1671 429 1672
rect 380 1667 381 1668
rect 423 1667 424 1671
rect 428 1670 429 1671
rect 431 1671 437 1672
rect 431 1670 432 1671
rect 428 1668 432 1670
rect 428 1667 429 1668
rect 375 1666 381 1667
rect 398 1666 404 1667
rect 423 1666 429 1667
rect 431 1667 432 1668
rect 436 1667 437 1671
rect 470 1671 476 1672
rect 470 1667 471 1671
rect 475 1670 476 1671
rect 487 1671 493 1672
rect 487 1670 488 1671
rect 475 1668 488 1670
rect 475 1667 476 1668
rect 431 1666 437 1667
rect 454 1666 460 1667
rect 470 1666 476 1667
rect 487 1667 488 1668
rect 492 1667 493 1671
rect 530 1671 536 1672
rect 530 1667 531 1671
rect 535 1670 536 1671
rect 551 1671 557 1672
rect 551 1670 552 1671
rect 535 1668 552 1670
rect 535 1667 536 1668
rect 487 1666 493 1667
rect 510 1666 516 1667
rect 530 1666 536 1667
rect 551 1667 552 1668
rect 556 1667 557 1671
rect 594 1671 600 1672
rect 594 1667 595 1671
rect 599 1670 600 1671
rect 623 1671 629 1672
rect 623 1670 624 1671
rect 599 1668 624 1670
rect 599 1667 600 1668
rect 551 1666 557 1667
rect 574 1666 580 1667
rect 594 1666 600 1667
rect 623 1667 624 1668
rect 628 1667 629 1671
rect 666 1671 672 1672
rect 666 1667 667 1671
rect 671 1670 672 1671
rect 703 1671 709 1672
rect 703 1670 704 1671
rect 671 1668 704 1670
rect 671 1667 672 1668
rect 623 1666 629 1667
rect 646 1666 652 1667
rect 666 1666 672 1667
rect 703 1667 704 1668
rect 708 1667 709 1671
rect 766 1671 772 1672
rect 766 1667 767 1671
rect 771 1670 772 1671
rect 783 1671 789 1672
rect 783 1670 784 1671
rect 771 1668 784 1670
rect 771 1667 772 1668
rect 703 1666 709 1667
rect 726 1666 732 1667
rect 766 1666 772 1667
rect 783 1667 784 1668
rect 788 1667 789 1671
rect 854 1671 860 1672
rect 854 1667 855 1671
rect 859 1670 860 1671
rect 863 1671 869 1672
rect 863 1670 864 1671
rect 859 1668 864 1670
rect 859 1667 860 1668
rect 783 1666 789 1667
rect 806 1666 812 1667
rect 854 1666 860 1667
rect 863 1667 864 1668
rect 868 1667 869 1671
rect 911 1671 917 1672
rect 911 1667 912 1671
rect 916 1670 917 1671
rect 943 1671 949 1672
rect 943 1670 944 1671
rect 916 1668 944 1670
rect 916 1667 917 1668
rect 863 1666 869 1667
rect 886 1666 892 1667
rect 911 1666 917 1667
rect 943 1667 944 1668
rect 948 1667 949 1671
rect 1022 1671 1029 1672
rect 1022 1667 1023 1671
rect 1028 1667 1029 1671
rect 1066 1671 1072 1672
rect 1066 1667 1067 1671
rect 1071 1670 1072 1671
rect 1111 1671 1117 1672
rect 1111 1670 1112 1671
rect 1071 1668 1112 1670
rect 1071 1667 1072 1668
rect 943 1666 949 1667
rect 966 1666 972 1667
rect 1022 1666 1029 1667
rect 1046 1666 1052 1667
rect 1066 1666 1072 1667
rect 1111 1667 1112 1668
rect 1116 1667 1117 1671
rect 1199 1671 1205 1672
rect 1199 1667 1200 1671
rect 1204 1670 1205 1671
rect 1216 1670 1218 1672
rect 1230 1671 1231 1672
rect 1235 1671 1236 1675
rect 1558 1674 1559 1678
rect 1563 1674 1564 1678
rect 1558 1673 1564 1674
rect 1630 1674 1631 1678
rect 1635 1674 1636 1678
rect 1630 1673 1636 1674
rect 1710 1674 1711 1678
rect 1715 1674 1716 1678
rect 1710 1673 1716 1674
rect 1798 1674 1799 1678
rect 1803 1674 1804 1678
rect 1798 1673 1804 1674
rect 1886 1674 1887 1678
rect 1891 1674 1892 1678
rect 1886 1673 1892 1674
rect 1974 1674 1975 1678
rect 1979 1674 1980 1678
rect 1974 1673 1980 1674
rect 2062 1674 2063 1678
rect 2067 1674 2068 1678
rect 2062 1673 2068 1674
rect 2142 1674 2143 1678
rect 2147 1674 2148 1678
rect 2142 1673 2148 1674
rect 2214 1674 2215 1678
rect 2219 1674 2220 1678
rect 2214 1673 2220 1674
rect 2286 1674 2287 1678
rect 2291 1674 2292 1678
rect 2286 1673 2292 1674
rect 2350 1674 2351 1678
rect 2355 1674 2356 1678
rect 2350 1673 2356 1674
rect 2422 1674 2423 1678
rect 2427 1674 2428 1678
rect 2422 1673 2428 1674
rect 2486 1674 2487 1678
rect 2491 1674 2492 1678
rect 2486 1673 2492 1674
rect 2542 1674 2543 1678
rect 2547 1674 2548 1678
rect 2542 1673 2548 1674
rect 1230 1670 1236 1671
rect 1242 1671 1248 1672
rect 1204 1668 1218 1670
rect 1204 1667 1205 1668
rect 1242 1667 1243 1671
rect 1247 1670 1248 1671
rect 1263 1671 1269 1672
rect 1263 1670 1264 1671
rect 1247 1668 1264 1670
rect 1247 1667 1248 1668
rect 1111 1666 1117 1667
rect 1134 1666 1140 1667
rect 1199 1666 1205 1667
rect 1222 1666 1228 1667
rect 1242 1666 1248 1667
rect 1263 1667 1264 1668
rect 1268 1667 1269 1671
rect 1366 1669 1372 1670
rect 1263 1666 1269 1667
rect 1286 1666 1292 1667
rect 398 1662 399 1666
rect 403 1662 404 1666
rect 398 1661 404 1662
rect 454 1662 455 1666
rect 459 1662 460 1666
rect 454 1661 460 1662
rect 510 1662 511 1666
rect 515 1662 516 1666
rect 510 1661 516 1662
rect 574 1662 575 1666
rect 579 1662 580 1666
rect 574 1661 580 1662
rect 646 1662 647 1666
rect 651 1662 652 1666
rect 646 1661 652 1662
rect 726 1662 727 1666
rect 731 1662 732 1666
rect 726 1661 732 1662
rect 806 1662 807 1666
rect 811 1662 812 1666
rect 806 1661 812 1662
rect 886 1662 887 1666
rect 891 1662 892 1666
rect 886 1661 892 1662
rect 966 1662 967 1666
rect 971 1662 972 1666
rect 966 1661 972 1662
rect 1046 1662 1047 1666
rect 1051 1662 1052 1666
rect 1046 1661 1052 1662
rect 1134 1662 1135 1666
rect 1139 1662 1140 1666
rect 1134 1661 1140 1662
rect 1222 1662 1223 1666
rect 1227 1662 1228 1666
rect 1222 1661 1228 1662
rect 1286 1662 1287 1666
rect 1291 1662 1292 1666
rect 1366 1665 1367 1669
rect 1371 1665 1372 1669
rect 1366 1664 1372 1665
rect 2582 1669 2588 1670
rect 2582 1665 2583 1669
rect 2587 1665 2588 1669
rect 2582 1664 2588 1665
rect 1286 1661 1292 1662
rect 2262 1659 2268 1660
rect 110 1657 116 1658
rect 110 1653 111 1657
rect 115 1653 116 1657
rect 110 1652 116 1653
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 2262 1655 2263 1659
rect 2267 1658 2268 1659
rect 2398 1659 2404 1660
rect 2267 1656 2362 1658
rect 2267 1655 2268 1656
rect 2262 1654 2268 1655
rect 1326 1652 1332 1653
rect 1366 1652 1372 1653
rect 1366 1648 1367 1652
rect 1371 1648 1372 1652
rect 1022 1647 1028 1648
rect 1366 1647 1372 1648
rect 1542 1651 1548 1652
rect 1542 1647 1543 1651
rect 1547 1647 1548 1651
rect 1614 1651 1620 1652
rect 1022 1643 1023 1647
rect 1027 1646 1028 1647
rect 1542 1646 1548 1647
rect 1575 1647 1584 1648
rect 1027 1644 1298 1646
rect 1027 1643 1028 1644
rect 1022 1642 1028 1643
rect 110 1640 116 1641
rect 110 1636 111 1640
rect 115 1636 116 1640
rect 110 1635 116 1636
rect 382 1639 388 1640
rect 382 1635 383 1639
rect 387 1635 388 1639
rect 438 1639 444 1640
rect 382 1634 388 1635
rect 415 1635 421 1636
rect 415 1631 416 1635
rect 420 1634 421 1635
rect 423 1635 429 1636
rect 423 1634 424 1635
rect 420 1632 424 1634
rect 420 1631 421 1632
rect 415 1630 421 1631
rect 423 1631 424 1632
rect 428 1631 429 1635
rect 438 1635 439 1639
rect 443 1635 444 1639
rect 494 1639 500 1640
rect 438 1634 444 1635
rect 470 1635 477 1636
rect 423 1630 429 1631
rect 470 1631 471 1635
rect 476 1631 477 1635
rect 494 1635 495 1639
rect 499 1635 500 1639
rect 558 1639 564 1640
rect 494 1634 500 1635
rect 527 1635 536 1636
rect 470 1630 477 1631
rect 527 1631 528 1635
rect 535 1631 536 1635
rect 558 1635 559 1639
rect 563 1635 564 1639
rect 630 1639 636 1640
rect 558 1634 564 1635
rect 591 1635 600 1636
rect 527 1630 536 1631
rect 591 1631 592 1635
rect 599 1631 600 1635
rect 630 1635 631 1639
rect 635 1635 636 1639
rect 710 1639 716 1640
rect 630 1634 636 1635
rect 663 1635 672 1636
rect 591 1630 600 1631
rect 663 1631 664 1635
rect 671 1631 672 1635
rect 710 1635 711 1639
rect 715 1635 716 1639
rect 766 1639 772 1640
rect 766 1638 767 1639
rect 710 1634 716 1635
rect 743 1637 767 1638
rect 743 1633 744 1637
rect 748 1636 767 1637
rect 748 1633 749 1636
rect 766 1635 767 1636
rect 771 1635 772 1639
rect 766 1634 772 1635
rect 790 1639 796 1640
rect 790 1635 791 1639
rect 795 1635 796 1639
rect 870 1639 876 1640
rect 790 1634 796 1635
rect 818 1635 829 1636
rect 743 1632 749 1633
rect 663 1630 672 1631
rect 818 1631 819 1635
rect 823 1631 824 1635
rect 828 1631 829 1635
rect 870 1635 871 1639
rect 875 1635 876 1639
rect 950 1639 956 1640
rect 870 1634 876 1635
rect 903 1635 909 1636
rect 818 1630 829 1631
rect 903 1631 904 1635
rect 908 1634 909 1635
rect 911 1635 917 1636
rect 911 1634 912 1635
rect 908 1632 912 1634
rect 908 1631 909 1632
rect 903 1630 909 1631
rect 911 1631 912 1632
rect 916 1631 917 1635
rect 950 1635 951 1639
rect 955 1635 956 1639
rect 1030 1639 1036 1640
rect 950 1634 956 1635
rect 982 1635 989 1636
rect 911 1630 917 1631
rect 982 1631 983 1635
rect 988 1631 989 1635
rect 1030 1635 1031 1639
rect 1035 1635 1036 1639
rect 1118 1639 1124 1640
rect 1030 1634 1036 1635
rect 1063 1635 1072 1636
rect 982 1630 989 1631
rect 1063 1631 1064 1635
rect 1071 1631 1072 1635
rect 1118 1635 1119 1639
rect 1123 1635 1124 1639
rect 1206 1639 1212 1640
rect 1118 1634 1124 1635
rect 1142 1635 1148 1636
rect 1063 1630 1072 1631
rect 1142 1631 1143 1635
rect 1147 1634 1148 1635
rect 1151 1635 1157 1636
rect 1151 1634 1152 1635
rect 1147 1632 1152 1634
rect 1147 1631 1148 1632
rect 1142 1630 1148 1631
rect 1151 1631 1152 1632
rect 1156 1631 1157 1635
rect 1206 1635 1207 1639
rect 1211 1635 1212 1639
rect 1270 1639 1276 1640
rect 1206 1634 1212 1635
rect 1239 1635 1248 1636
rect 1151 1630 1157 1631
rect 1239 1631 1240 1635
rect 1247 1631 1248 1635
rect 1270 1635 1271 1639
rect 1275 1635 1276 1639
rect 1270 1634 1276 1635
rect 1296 1634 1298 1644
rect 1575 1643 1576 1647
rect 1583 1643 1584 1647
rect 1614 1647 1615 1651
rect 1619 1647 1620 1651
rect 1694 1651 1700 1652
rect 1614 1646 1620 1647
rect 1647 1647 1656 1648
rect 1575 1642 1584 1643
rect 1647 1643 1648 1647
rect 1655 1643 1656 1647
rect 1694 1647 1695 1651
rect 1699 1647 1700 1651
rect 1782 1651 1788 1652
rect 1694 1646 1700 1647
rect 1722 1647 1733 1648
rect 1647 1642 1656 1643
rect 1722 1643 1723 1647
rect 1727 1643 1728 1647
rect 1732 1643 1733 1647
rect 1782 1647 1783 1651
rect 1787 1647 1788 1651
rect 1870 1651 1876 1652
rect 1782 1646 1788 1647
rect 1815 1647 1824 1648
rect 1722 1642 1733 1643
rect 1815 1643 1816 1647
rect 1823 1643 1824 1647
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 1958 1651 1964 1652
rect 1870 1646 1876 1647
rect 1902 1647 1909 1648
rect 1815 1642 1824 1643
rect 1902 1643 1903 1647
rect 1908 1643 1909 1647
rect 1958 1647 1959 1651
rect 1963 1647 1964 1651
rect 2046 1651 2052 1652
rect 1958 1646 1964 1647
rect 1982 1647 1988 1648
rect 1902 1642 1909 1643
rect 1982 1643 1983 1647
rect 1987 1646 1988 1647
rect 1991 1647 1997 1648
rect 1991 1646 1992 1647
rect 1987 1644 1992 1646
rect 1987 1643 1988 1644
rect 1982 1642 1988 1643
rect 1991 1643 1992 1644
rect 1996 1643 1997 1647
rect 2046 1647 2047 1651
rect 2051 1647 2052 1651
rect 2126 1651 2132 1652
rect 2046 1646 2052 1647
rect 2079 1647 2088 1648
rect 1991 1642 1997 1643
rect 2079 1643 2080 1647
rect 2087 1643 2088 1647
rect 2126 1647 2127 1651
rect 2131 1647 2132 1651
rect 2198 1651 2204 1652
rect 2126 1646 2132 1647
rect 2159 1647 2168 1648
rect 2079 1642 2088 1643
rect 2159 1643 2160 1647
rect 2167 1643 2168 1647
rect 2198 1647 2199 1651
rect 2203 1647 2204 1651
rect 2270 1651 2276 1652
rect 2198 1646 2204 1647
rect 2230 1647 2237 1648
rect 2159 1642 2168 1643
rect 2230 1643 2231 1647
rect 2236 1643 2237 1647
rect 2270 1647 2271 1651
rect 2275 1647 2276 1651
rect 2334 1651 2340 1652
rect 2270 1646 2276 1647
rect 2294 1647 2300 1648
rect 2230 1642 2237 1643
rect 2294 1643 2295 1647
rect 2299 1646 2300 1647
rect 2303 1647 2309 1648
rect 2303 1646 2304 1647
rect 2299 1644 2304 1646
rect 2299 1643 2300 1644
rect 2294 1642 2300 1643
rect 2303 1643 2304 1644
rect 2308 1643 2309 1647
rect 2334 1647 2335 1651
rect 2339 1647 2340 1651
rect 2334 1646 2340 1647
rect 2360 1646 2362 1656
rect 2398 1655 2399 1659
rect 2403 1658 2404 1659
rect 2403 1656 2498 1658
rect 2403 1655 2404 1656
rect 2398 1654 2404 1655
rect 2406 1651 2412 1652
rect 2367 1647 2373 1648
rect 2367 1646 2368 1647
rect 2360 1644 2368 1646
rect 2303 1642 2309 1643
rect 2367 1643 2368 1644
rect 2372 1643 2373 1647
rect 2406 1647 2407 1651
rect 2411 1647 2412 1651
rect 2470 1651 2476 1652
rect 2406 1646 2412 1647
rect 2434 1647 2445 1648
rect 2367 1642 2373 1643
rect 2434 1643 2435 1647
rect 2439 1643 2440 1647
rect 2444 1643 2445 1647
rect 2470 1647 2471 1651
rect 2475 1647 2476 1651
rect 2470 1646 2476 1647
rect 2496 1646 2498 1656
rect 2582 1652 2588 1653
rect 2526 1651 2532 1652
rect 2503 1647 2509 1648
rect 2503 1646 2504 1647
rect 2496 1644 2504 1646
rect 2434 1642 2445 1643
rect 2503 1643 2504 1644
rect 2508 1643 2509 1647
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2582 1648 2583 1652
rect 2587 1648 2588 1652
rect 2526 1646 2532 1647
rect 2558 1647 2565 1648
rect 2582 1647 2588 1648
rect 2503 1642 2509 1643
rect 2558 1643 2559 1647
rect 2564 1643 2565 1647
rect 2558 1642 2565 1643
rect 1326 1640 1332 1641
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1303 1635 1309 1636
rect 1326 1635 1332 1636
rect 1303 1634 1304 1635
rect 1296 1632 1304 1634
rect 1239 1630 1248 1631
rect 1303 1631 1304 1632
rect 1308 1631 1309 1635
rect 1303 1630 1309 1631
rect 1550 1611 1556 1612
rect 1550 1607 1551 1611
rect 1555 1610 1556 1611
rect 1615 1611 1621 1612
rect 1555 1608 1602 1610
rect 1555 1607 1556 1608
rect 1550 1606 1556 1607
rect 1600 1606 1602 1608
rect 1607 1607 1613 1608
rect 1607 1606 1608 1607
rect 1574 1605 1580 1606
rect 1366 1604 1372 1605
rect 1366 1600 1367 1604
rect 1371 1600 1372 1604
rect 1574 1601 1575 1605
rect 1579 1601 1580 1605
rect 1600 1604 1608 1606
rect 1607 1603 1608 1604
rect 1612 1603 1613 1607
rect 1615 1607 1616 1611
rect 1620 1610 1621 1611
rect 1671 1611 1677 1612
rect 1620 1608 1658 1610
rect 1620 1607 1621 1608
rect 1615 1606 1621 1607
rect 1656 1606 1658 1608
rect 1663 1607 1669 1608
rect 1663 1606 1664 1607
rect 1607 1602 1613 1603
rect 1630 1605 1636 1606
rect 1574 1600 1580 1601
rect 1630 1601 1631 1605
rect 1635 1601 1636 1605
rect 1656 1604 1664 1606
rect 1663 1603 1664 1604
rect 1668 1603 1669 1607
rect 1671 1607 1672 1611
rect 1676 1610 1677 1611
rect 1727 1611 1733 1612
rect 1676 1608 1723 1610
rect 1676 1607 1677 1608
rect 1671 1606 1677 1607
rect 1719 1607 1725 1608
rect 1663 1602 1669 1603
rect 1686 1605 1692 1606
rect 1630 1600 1636 1601
rect 1686 1601 1687 1605
rect 1691 1601 1692 1605
rect 1719 1603 1720 1607
rect 1724 1603 1725 1607
rect 1727 1607 1728 1611
rect 1732 1610 1733 1611
rect 1791 1611 1797 1612
rect 1732 1608 1778 1610
rect 1732 1607 1733 1608
rect 1727 1606 1733 1607
rect 1776 1606 1778 1608
rect 1783 1607 1789 1608
rect 1783 1606 1784 1607
rect 1719 1602 1725 1603
rect 1750 1605 1756 1606
rect 1686 1600 1692 1601
rect 1750 1601 1751 1605
rect 1755 1601 1756 1605
rect 1776 1604 1784 1606
rect 1783 1603 1784 1604
rect 1788 1603 1789 1607
rect 1791 1607 1792 1611
rect 1796 1610 1797 1611
rect 2534 1611 2540 1612
rect 1796 1608 1858 1610
rect 1796 1607 1797 1608
rect 1791 1606 1797 1607
rect 1856 1606 1858 1608
rect 1863 1607 1869 1608
rect 1863 1606 1864 1607
rect 1783 1602 1789 1603
rect 1830 1605 1836 1606
rect 1750 1600 1756 1601
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1856 1604 1864 1606
rect 1863 1603 1864 1604
rect 1868 1603 1869 1607
rect 1951 1607 1957 1608
rect 1863 1602 1869 1603
rect 1918 1605 1924 1606
rect 1830 1600 1836 1601
rect 1918 1601 1919 1605
rect 1923 1601 1924 1605
rect 1951 1603 1952 1607
rect 1956 1606 1957 1607
rect 1998 1607 2004 1608
rect 1998 1606 1999 1607
rect 1956 1604 1999 1606
rect 1956 1603 1957 1604
rect 1951 1602 1957 1603
rect 1998 1603 1999 1604
rect 2003 1603 2004 1607
rect 2039 1607 2045 1608
rect 1998 1602 2004 1603
rect 2006 1605 2012 1606
rect 1918 1600 1924 1601
rect 2006 1601 2007 1605
rect 2011 1601 2012 1605
rect 2039 1603 2040 1607
rect 2044 1606 2045 1607
rect 2094 1607 2100 1608
rect 2094 1606 2095 1607
rect 2044 1604 2095 1606
rect 2044 1603 2045 1604
rect 2039 1602 2045 1603
rect 2094 1603 2095 1604
rect 2099 1603 2100 1607
rect 2126 1607 2132 1608
rect 2094 1602 2100 1603
rect 2102 1605 2108 1606
rect 2006 1600 2012 1601
rect 2102 1601 2103 1605
rect 2107 1601 2108 1605
rect 2126 1603 2127 1607
rect 2131 1606 2132 1607
rect 2135 1607 2141 1608
rect 2135 1606 2136 1607
rect 2131 1604 2136 1606
rect 2131 1603 2132 1604
rect 2126 1602 2132 1603
rect 2135 1603 2136 1604
rect 2140 1603 2141 1607
rect 2239 1607 2245 1608
rect 2135 1602 2141 1603
rect 2206 1605 2212 1606
rect 2102 1600 2108 1601
rect 2206 1601 2207 1605
rect 2211 1601 2212 1605
rect 2239 1603 2240 1607
rect 2244 1606 2245 1607
rect 2310 1607 2316 1608
rect 2310 1606 2311 1607
rect 2244 1604 2311 1606
rect 2244 1603 2245 1604
rect 2239 1602 2245 1603
rect 2310 1603 2311 1604
rect 2315 1603 2316 1607
rect 2351 1607 2357 1608
rect 2310 1602 2316 1603
rect 2318 1605 2324 1606
rect 2206 1600 2212 1601
rect 2318 1601 2319 1605
rect 2323 1601 2324 1605
rect 2351 1603 2352 1607
rect 2356 1606 2357 1607
rect 2422 1607 2428 1608
rect 2422 1606 2423 1607
rect 2356 1604 2423 1606
rect 2356 1603 2357 1604
rect 2351 1602 2357 1603
rect 2422 1603 2423 1604
rect 2427 1603 2428 1607
rect 2462 1607 2469 1608
rect 2422 1602 2428 1603
rect 2430 1605 2436 1606
rect 2318 1600 2324 1601
rect 2430 1601 2431 1605
rect 2435 1601 2436 1605
rect 2462 1603 2463 1607
rect 2468 1603 2469 1607
rect 2534 1607 2535 1611
rect 2539 1610 2540 1611
rect 2539 1608 2563 1610
rect 2539 1607 2540 1608
rect 2534 1606 2540 1607
rect 2559 1607 2565 1608
rect 2462 1602 2469 1603
rect 2526 1605 2532 1606
rect 2430 1600 2436 1601
rect 2526 1601 2527 1605
rect 2531 1601 2532 1605
rect 2559 1603 2560 1607
rect 2564 1603 2565 1607
rect 2559 1602 2565 1603
rect 2582 1604 2588 1605
rect 2526 1600 2532 1601
rect 2582 1600 2583 1604
rect 2587 1600 2588 1604
rect 910 1599 916 1600
rect 1366 1599 1372 1600
rect 2582 1599 2588 1600
rect 910 1595 911 1599
rect 915 1598 916 1599
rect 915 1596 1090 1598
rect 915 1595 916 1596
rect 910 1594 916 1595
rect 319 1591 325 1592
rect 286 1589 292 1590
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 286 1585 287 1589
rect 291 1585 292 1589
rect 319 1587 320 1591
rect 324 1590 325 1591
rect 358 1591 364 1592
rect 358 1590 359 1591
rect 324 1588 359 1590
rect 324 1587 325 1588
rect 319 1586 325 1587
rect 358 1587 359 1588
rect 363 1587 364 1591
rect 399 1591 405 1592
rect 358 1586 364 1587
rect 366 1589 372 1590
rect 286 1584 292 1585
rect 366 1585 367 1589
rect 371 1585 372 1589
rect 399 1587 400 1591
rect 404 1590 405 1591
rect 446 1591 452 1592
rect 446 1590 447 1591
rect 404 1588 447 1590
rect 404 1587 405 1588
rect 399 1586 405 1587
rect 446 1587 447 1588
rect 451 1587 452 1591
rect 487 1591 493 1592
rect 446 1586 452 1587
rect 454 1589 460 1590
rect 366 1584 372 1585
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 487 1587 488 1591
rect 492 1590 493 1591
rect 534 1591 540 1592
rect 534 1590 535 1591
rect 492 1588 535 1590
rect 492 1587 493 1588
rect 487 1586 493 1587
rect 534 1587 535 1588
rect 539 1587 540 1591
rect 583 1591 589 1592
rect 534 1586 540 1587
rect 550 1589 556 1590
rect 454 1584 460 1585
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 583 1587 584 1591
rect 588 1590 589 1591
rect 638 1591 644 1592
rect 638 1590 639 1591
rect 588 1588 639 1590
rect 588 1587 589 1588
rect 583 1586 589 1587
rect 638 1587 639 1588
rect 643 1587 644 1591
rect 670 1591 676 1592
rect 638 1586 644 1587
rect 646 1589 652 1590
rect 550 1584 556 1585
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 670 1587 671 1591
rect 675 1590 676 1591
rect 679 1591 685 1592
rect 679 1590 680 1591
rect 675 1588 680 1590
rect 675 1587 676 1588
rect 670 1586 676 1587
rect 679 1587 680 1588
rect 684 1587 685 1591
rect 767 1591 773 1592
rect 679 1586 685 1587
rect 734 1589 740 1590
rect 646 1584 652 1585
rect 734 1585 735 1589
rect 739 1585 740 1589
rect 767 1587 768 1591
rect 772 1590 773 1591
rect 814 1591 820 1592
rect 814 1590 815 1591
rect 772 1588 815 1590
rect 772 1587 773 1588
rect 767 1586 773 1587
rect 814 1587 815 1588
rect 819 1587 820 1591
rect 854 1591 861 1592
rect 814 1586 820 1587
rect 822 1589 828 1590
rect 734 1584 740 1585
rect 822 1585 823 1589
rect 827 1585 828 1589
rect 854 1587 855 1591
rect 860 1587 861 1591
rect 935 1591 941 1592
rect 854 1586 861 1587
rect 902 1589 908 1590
rect 822 1584 828 1585
rect 902 1585 903 1589
rect 907 1585 908 1589
rect 935 1587 936 1591
rect 940 1590 941 1591
rect 967 1591 973 1592
rect 967 1590 968 1591
rect 940 1588 968 1590
rect 940 1587 941 1588
rect 935 1586 941 1587
rect 967 1587 968 1588
rect 972 1587 973 1591
rect 1015 1591 1021 1592
rect 967 1586 973 1587
rect 982 1589 988 1590
rect 902 1584 908 1585
rect 982 1585 983 1589
rect 987 1585 988 1589
rect 1015 1587 1016 1591
rect 1020 1590 1021 1591
rect 1030 1591 1036 1592
rect 1030 1590 1031 1591
rect 1020 1588 1031 1590
rect 1020 1587 1021 1588
rect 1015 1586 1021 1587
rect 1030 1587 1031 1588
rect 1035 1587 1036 1591
rect 1088 1590 1090 1596
rect 1103 1595 1109 1596
rect 1095 1591 1101 1592
rect 1095 1590 1096 1591
rect 1030 1586 1036 1587
rect 1062 1589 1068 1590
rect 982 1584 988 1585
rect 1062 1585 1063 1589
rect 1067 1585 1068 1589
rect 1088 1588 1096 1590
rect 1095 1587 1096 1588
rect 1100 1587 1101 1591
rect 1103 1591 1104 1595
rect 1108 1594 1109 1595
rect 1108 1592 1178 1594
rect 1108 1591 1109 1592
rect 1103 1590 1109 1591
rect 1176 1590 1178 1592
rect 1183 1591 1189 1592
rect 1183 1590 1184 1591
rect 1095 1586 1101 1587
rect 1150 1589 1156 1590
rect 1062 1584 1068 1585
rect 1150 1585 1151 1589
rect 1155 1585 1156 1589
rect 1176 1588 1184 1590
rect 1183 1587 1184 1588
rect 1188 1587 1189 1591
rect 1183 1586 1189 1587
rect 1326 1588 1332 1589
rect 1150 1584 1156 1585
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 110 1583 116 1584
rect 1326 1583 1332 1584
rect 1366 1587 1372 1588
rect 1366 1583 1367 1587
rect 1371 1583 1372 1587
rect 1366 1582 1372 1583
rect 2582 1587 2588 1588
rect 2582 1583 2583 1587
rect 2587 1583 2588 1587
rect 2582 1582 2588 1583
rect 1590 1578 1596 1579
rect 1590 1574 1591 1578
rect 1595 1574 1596 1578
rect 1590 1573 1596 1574
rect 1646 1578 1652 1579
rect 1646 1574 1647 1578
rect 1651 1574 1652 1578
rect 1646 1573 1652 1574
rect 1702 1578 1708 1579
rect 1702 1574 1703 1578
rect 1707 1574 1708 1578
rect 1702 1573 1708 1574
rect 1766 1578 1772 1579
rect 1766 1574 1767 1578
rect 1771 1574 1772 1578
rect 1766 1573 1772 1574
rect 1846 1578 1852 1579
rect 1846 1574 1847 1578
rect 1851 1574 1852 1578
rect 1846 1573 1852 1574
rect 1934 1578 1940 1579
rect 1934 1574 1935 1578
rect 1939 1574 1940 1578
rect 1934 1573 1940 1574
rect 2022 1578 2028 1579
rect 2022 1574 2023 1578
rect 2027 1574 2028 1578
rect 2022 1573 2028 1574
rect 2118 1578 2124 1579
rect 2118 1574 2119 1578
rect 2123 1574 2124 1578
rect 2118 1573 2124 1574
rect 2222 1578 2228 1579
rect 2222 1574 2223 1578
rect 2227 1574 2228 1578
rect 2222 1573 2228 1574
rect 2334 1578 2340 1579
rect 2334 1574 2335 1578
rect 2339 1574 2340 1578
rect 2334 1573 2340 1574
rect 2446 1578 2452 1579
rect 2446 1574 2447 1578
rect 2451 1574 2452 1578
rect 2446 1573 2452 1574
rect 2542 1578 2548 1579
rect 2542 1574 2543 1578
rect 2547 1574 2548 1578
rect 2542 1573 2548 1574
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 110 1566 116 1567
rect 1326 1571 1332 1572
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 1326 1566 1332 1567
rect 1567 1571 1573 1572
rect 1567 1567 1568 1571
rect 1572 1570 1573 1571
rect 1615 1571 1621 1572
rect 1615 1570 1616 1571
rect 1572 1568 1616 1570
rect 1572 1567 1573 1568
rect 1567 1566 1573 1567
rect 1615 1567 1616 1568
rect 1620 1567 1621 1571
rect 1615 1566 1621 1567
rect 1623 1571 1629 1572
rect 1623 1567 1624 1571
rect 1628 1570 1629 1571
rect 1671 1571 1677 1572
rect 1671 1570 1672 1571
rect 1628 1568 1672 1570
rect 1628 1567 1629 1568
rect 1623 1566 1629 1567
rect 1671 1567 1672 1568
rect 1676 1567 1677 1571
rect 1671 1566 1677 1567
rect 1679 1571 1685 1572
rect 1679 1567 1680 1571
rect 1684 1570 1685 1571
rect 1727 1571 1733 1572
rect 1727 1570 1728 1571
rect 1684 1568 1728 1570
rect 1684 1567 1685 1568
rect 1679 1566 1685 1567
rect 1727 1567 1728 1568
rect 1732 1567 1733 1571
rect 1727 1566 1733 1567
rect 1743 1571 1749 1572
rect 1743 1567 1744 1571
rect 1748 1570 1749 1571
rect 1791 1571 1797 1572
rect 1791 1570 1792 1571
rect 1748 1568 1792 1570
rect 1748 1567 1749 1568
rect 1743 1566 1749 1567
rect 1791 1567 1792 1568
rect 1796 1567 1797 1571
rect 1791 1566 1797 1567
rect 1823 1571 1829 1572
rect 1823 1567 1824 1571
rect 1828 1570 1829 1571
rect 1902 1571 1908 1572
rect 1902 1570 1903 1571
rect 1828 1568 1903 1570
rect 1828 1567 1829 1568
rect 1823 1566 1829 1567
rect 1902 1567 1903 1568
rect 1907 1567 1908 1571
rect 1902 1566 1908 1567
rect 1911 1571 1917 1572
rect 1911 1567 1912 1571
rect 1916 1570 1917 1571
rect 1982 1571 1988 1572
rect 1982 1570 1983 1571
rect 1916 1568 1983 1570
rect 1916 1567 1917 1568
rect 1911 1566 1917 1567
rect 1982 1567 1983 1568
rect 1987 1567 1988 1571
rect 1982 1566 1988 1567
rect 1998 1571 2005 1572
rect 1998 1567 1999 1571
rect 2004 1567 2005 1571
rect 1998 1566 2005 1567
rect 2094 1571 2101 1572
rect 2094 1567 2095 1571
rect 2100 1567 2101 1571
rect 2094 1566 2101 1567
rect 2191 1571 2197 1572
rect 2191 1567 2192 1571
rect 2196 1570 2197 1571
rect 2199 1571 2205 1572
rect 2199 1570 2200 1571
rect 2196 1568 2200 1570
rect 2196 1567 2197 1568
rect 2191 1566 2197 1567
rect 2199 1567 2200 1568
rect 2204 1567 2205 1571
rect 2199 1566 2205 1567
rect 2310 1571 2317 1572
rect 2310 1567 2311 1571
rect 2316 1567 2317 1571
rect 2310 1566 2317 1567
rect 2422 1571 2429 1572
rect 2422 1567 2423 1571
rect 2428 1567 2429 1571
rect 2422 1566 2429 1567
rect 2519 1571 2525 1572
rect 2519 1567 2520 1571
rect 2524 1570 2525 1571
rect 2558 1571 2564 1572
rect 2558 1570 2559 1571
rect 2524 1568 2559 1570
rect 2524 1567 2525 1568
rect 2519 1566 2525 1567
rect 2558 1567 2559 1568
rect 2563 1567 2564 1571
rect 2558 1566 2564 1567
rect 2342 1563 2348 1564
rect 302 1562 308 1563
rect 302 1558 303 1562
rect 307 1558 308 1562
rect 302 1557 308 1558
rect 382 1562 388 1563
rect 382 1558 383 1562
rect 387 1558 388 1562
rect 382 1557 388 1558
rect 470 1562 476 1563
rect 470 1558 471 1562
rect 475 1558 476 1562
rect 470 1557 476 1558
rect 566 1562 572 1563
rect 566 1558 567 1562
rect 571 1558 572 1562
rect 566 1557 572 1558
rect 662 1562 668 1563
rect 662 1558 663 1562
rect 667 1558 668 1562
rect 662 1557 668 1558
rect 750 1562 756 1563
rect 750 1558 751 1562
rect 755 1558 756 1562
rect 750 1557 756 1558
rect 838 1562 844 1563
rect 838 1558 839 1562
rect 843 1558 844 1562
rect 838 1557 844 1558
rect 918 1562 924 1563
rect 918 1558 919 1562
rect 923 1558 924 1562
rect 918 1557 924 1558
rect 998 1562 1004 1563
rect 998 1558 999 1562
rect 1003 1558 1004 1562
rect 998 1557 1004 1558
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1166 1562 1172 1563
rect 2342 1562 2343 1563
rect 1166 1558 1167 1562
rect 1171 1558 1172 1562
rect 2225 1560 2343 1562
rect 2126 1559 2132 1560
rect 2126 1558 2127 1559
rect 1166 1557 1172 1558
rect 2080 1556 2127 1558
rect 279 1555 285 1556
rect 279 1551 280 1555
rect 284 1554 285 1555
rect 294 1555 300 1556
rect 294 1554 295 1555
rect 284 1552 295 1554
rect 284 1551 285 1552
rect 279 1550 285 1551
rect 294 1551 295 1552
rect 299 1551 300 1555
rect 294 1550 300 1551
rect 358 1555 365 1556
rect 358 1551 359 1555
rect 364 1551 365 1555
rect 446 1555 453 1556
rect 358 1550 365 1551
rect 414 1551 420 1552
rect 414 1550 415 1551
rect 368 1548 415 1550
rect 368 1546 370 1548
rect 414 1547 415 1548
rect 419 1547 420 1551
rect 446 1551 447 1555
rect 452 1551 453 1555
rect 446 1550 453 1551
rect 534 1555 540 1556
rect 534 1551 535 1555
rect 539 1554 540 1555
rect 543 1555 549 1556
rect 543 1554 544 1555
rect 539 1552 544 1554
rect 539 1551 540 1552
rect 534 1550 540 1551
rect 543 1551 544 1552
rect 548 1551 549 1555
rect 543 1550 549 1551
rect 638 1555 645 1556
rect 638 1551 639 1555
rect 644 1551 645 1555
rect 706 1555 712 1556
rect 638 1550 645 1551
rect 670 1551 676 1552
rect 670 1550 671 1551
rect 414 1546 420 1547
rect 648 1548 671 1550
rect 648 1546 650 1548
rect 670 1547 671 1548
rect 675 1547 676 1551
rect 706 1551 707 1555
rect 711 1554 712 1555
rect 727 1555 733 1556
rect 727 1554 728 1555
rect 711 1552 728 1554
rect 711 1551 712 1552
rect 706 1550 712 1551
rect 727 1551 728 1552
rect 732 1551 733 1555
rect 727 1550 733 1551
rect 814 1555 821 1556
rect 814 1551 815 1555
rect 820 1551 821 1555
rect 814 1550 821 1551
rect 895 1555 901 1556
rect 895 1551 896 1555
rect 900 1554 901 1555
rect 910 1555 916 1556
rect 910 1554 911 1555
rect 900 1552 911 1554
rect 900 1551 901 1552
rect 895 1550 901 1551
rect 910 1551 911 1552
rect 915 1551 916 1555
rect 910 1550 916 1551
rect 967 1555 973 1556
rect 967 1551 968 1555
rect 972 1554 973 1555
rect 975 1555 981 1556
rect 975 1554 976 1555
rect 972 1552 976 1554
rect 972 1551 973 1552
rect 967 1550 973 1551
rect 975 1551 976 1552
rect 980 1551 981 1555
rect 975 1550 981 1551
rect 1055 1555 1061 1556
rect 1055 1551 1056 1555
rect 1060 1554 1061 1555
rect 1103 1555 1109 1556
rect 1103 1554 1104 1555
rect 1060 1552 1104 1554
rect 1060 1551 1061 1552
rect 1055 1550 1061 1551
rect 1103 1551 1104 1552
rect 1108 1551 1109 1555
rect 1103 1550 1109 1551
rect 1142 1555 1149 1556
rect 1142 1551 1143 1555
rect 1148 1551 1149 1555
rect 1142 1550 1149 1551
rect 1655 1555 1661 1556
rect 1655 1551 1656 1555
rect 1660 1554 1661 1555
rect 1670 1555 1676 1556
rect 1670 1554 1671 1555
rect 1660 1552 1671 1554
rect 1660 1551 1661 1552
rect 1655 1550 1661 1551
rect 1670 1551 1671 1552
rect 1675 1551 1676 1555
rect 1703 1555 1709 1556
rect 1703 1551 1704 1555
rect 1708 1554 1709 1555
rect 1711 1555 1717 1556
rect 1711 1554 1712 1555
rect 1708 1552 1712 1554
rect 1708 1551 1709 1552
rect 1670 1550 1676 1551
rect 1678 1550 1684 1551
rect 1703 1550 1709 1551
rect 1711 1551 1712 1552
rect 1716 1551 1717 1555
rect 1754 1555 1760 1556
rect 1754 1551 1755 1555
rect 1759 1554 1760 1555
rect 1767 1555 1773 1556
rect 1767 1554 1768 1555
rect 1759 1552 1768 1554
rect 1759 1551 1760 1552
rect 1711 1550 1717 1551
rect 1734 1550 1740 1551
rect 1754 1550 1760 1551
rect 1767 1551 1768 1552
rect 1772 1551 1773 1555
rect 1810 1555 1816 1556
rect 1810 1551 1811 1555
rect 1815 1554 1816 1555
rect 1831 1555 1837 1556
rect 1831 1554 1832 1555
rect 1815 1552 1832 1554
rect 1815 1551 1816 1552
rect 1767 1550 1773 1551
rect 1790 1550 1796 1551
rect 1810 1550 1816 1551
rect 1831 1551 1832 1552
rect 1836 1551 1837 1555
rect 1874 1555 1880 1556
rect 1874 1551 1875 1555
rect 1879 1554 1880 1555
rect 1903 1555 1909 1556
rect 1903 1554 1904 1555
rect 1879 1552 1904 1554
rect 1879 1551 1880 1552
rect 1831 1550 1837 1551
rect 1854 1550 1860 1551
rect 1874 1550 1880 1551
rect 1903 1551 1904 1552
rect 1908 1551 1909 1555
rect 1946 1555 1952 1556
rect 1946 1551 1947 1555
rect 1951 1554 1952 1555
rect 1983 1555 1989 1556
rect 1983 1554 1984 1555
rect 1951 1552 1984 1554
rect 1951 1551 1952 1552
rect 1903 1550 1909 1551
rect 1926 1550 1932 1551
rect 1946 1550 1952 1551
rect 1983 1551 1984 1552
rect 1988 1551 1989 1555
rect 2063 1555 2069 1556
rect 2063 1551 2064 1555
rect 2068 1554 2069 1555
rect 2080 1554 2082 1556
rect 2126 1555 2127 1556
rect 2131 1555 2132 1559
rect 2225 1556 2227 1560
rect 2342 1559 2343 1560
rect 2347 1559 2348 1563
rect 2342 1558 2348 1559
rect 2126 1554 2132 1555
rect 2142 1555 2149 1556
rect 2068 1552 2082 1554
rect 2068 1551 2069 1552
rect 2142 1551 2143 1555
rect 2148 1551 2149 1555
rect 2223 1555 2229 1556
rect 2223 1551 2224 1555
rect 2228 1551 2229 1555
rect 2266 1555 2272 1556
rect 2266 1551 2267 1555
rect 2271 1554 2272 1555
rect 2303 1555 2309 1556
rect 2303 1554 2304 1555
rect 2271 1552 2304 1554
rect 2271 1551 2272 1552
rect 1983 1550 1989 1551
rect 2006 1550 2012 1551
rect 2063 1550 2069 1551
rect 2086 1550 2092 1551
rect 2142 1550 2149 1551
rect 2166 1550 2172 1551
rect 2223 1550 2229 1551
rect 2246 1550 2252 1551
rect 2266 1550 2272 1551
rect 2303 1551 2304 1552
rect 2308 1551 2309 1555
rect 2382 1555 2389 1556
rect 2382 1551 2383 1555
rect 2388 1551 2389 1555
rect 2462 1555 2469 1556
rect 2462 1551 2463 1555
rect 2468 1551 2469 1555
rect 2519 1555 2525 1556
rect 2519 1551 2520 1555
rect 2524 1554 2525 1555
rect 2534 1555 2540 1556
rect 2534 1554 2535 1555
rect 2524 1552 2535 1554
rect 2524 1551 2525 1552
rect 2303 1550 2309 1551
rect 2326 1550 2332 1551
rect 2382 1550 2389 1551
rect 2406 1550 2412 1551
rect 2462 1550 2469 1551
rect 2486 1550 2492 1551
rect 2519 1550 2525 1551
rect 2534 1551 2535 1552
rect 2539 1551 2540 1555
rect 2534 1550 2540 1551
rect 2542 1550 2548 1551
rect 670 1546 676 1547
rect 1678 1546 1679 1550
rect 1683 1546 1684 1550
rect 319 1544 370 1546
rect 608 1544 650 1546
rect 1678 1545 1684 1546
rect 1734 1546 1735 1550
rect 1739 1546 1740 1550
rect 1734 1545 1740 1546
rect 1790 1546 1791 1550
rect 1795 1546 1796 1550
rect 1790 1545 1796 1546
rect 1854 1546 1855 1550
rect 1859 1546 1860 1550
rect 1854 1545 1860 1546
rect 1926 1546 1927 1550
rect 1931 1546 1932 1550
rect 1926 1545 1932 1546
rect 2006 1546 2007 1550
rect 2011 1546 2012 1550
rect 2006 1545 2012 1546
rect 2086 1546 2087 1550
rect 2091 1546 2092 1550
rect 2086 1545 2092 1546
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2246 1546 2247 1550
rect 2251 1546 2252 1550
rect 2246 1545 2252 1546
rect 2326 1546 2327 1550
rect 2331 1546 2332 1550
rect 2326 1545 2332 1546
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2486 1546 2487 1550
rect 2491 1546 2492 1550
rect 2486 1545 2492 1546
rect 2542 1546 2543 1550
rect 2547 1546 2548 1550
rect 2542 1545 2548 1546
rect 254 1543 261 1544
rect 254 1539 255 1543
rect 260 1539 261 1543
rect 311 1543 317 1544
rect 311 1539 312 1543
rect 316 1542 317 1543
rect 319 1542 321 1544
rect 316 1540 321 1542
rect 375 1543 381 1544
rect 316 1539 317 1540
rect 375 1539 376 1543
rect 380 1542 381 1543
rect 390 1543 396 1544
rect 390 1542 391 1543
rect 380 1540 391 1542
rect 380 1539 381 1540
rect 254 1538 261 1539
rect 278 1538 284 1539
rect 311 1538 317 1539
rect 334 1538 340 1539
rect 375 1538 381 1539
rect 390 1539 391 1540
rect 395 1539 396 1543
rect 446 1543 453 1544
rect 446 1539 447 1543
rect 452 1539 453 1543
rect 490 1543 496 1544
rect 490 1539 491 1543
rect 495 1542 496 1543
rect 519 1543 525 1544
rect 519 1542 520 1543
rect 495 1540 520 1542
rect 495 1539 496 1540
rect 390 1538 396 1539
rect 398 1538 404 1539
rect 446 1538 453 1539
rect 470 1538 476 1539
rect 490 1538 496 1539
rect 519 1539 520 1540
rect 524 1539 525 1543
rect 591 1543 597 1544
rect 591 1539 592 1543
rect 596 1542 597 1543
rect 608 1542 610 1544
rect 596 1540 610 1542
rect 663 1543 669 1544
rect 596 1539 597 1540
rect 663 1539 664 1543
rect 668 1542 669 1543
rect 678 1543 684 1544
rect 678 1542 679 1543
rect 668 1540 679 1542
rect 668 1539 669 1540
rect 519 1538 525 1539
rect 542 1538 548 1539
rect 591 1538 597 1539
rect 614 1538 620 1539
rect 663 1538 669 1539
rect 678 1539 679 1540
rect 683 1539 684 1543
rect 734 1543 741 1544
rect 734 1539 735 1543
rect 740 1539 741 1543
rect 806 1543 813 1544
rect 806 1539 807 1543
rect 812 1539 813 1543
rect 878 1543 885 1544
rect 878 1539 879 1543
rect 884 1539 885 1543
rect 951 1543 957 1544
rect 951 1539 952 1543
rect 956 1542 957 1543
rect 966 1543 972 1544
rect 966 1542 967 1543
rect 956 1540 967 1542
rect 956 1539 957 1540
rect 678 1538 684 1539
rect 686 1538 692 1539
rect 734 1538 741 1539
rect 758 1538 764 1539
rect 806 1538 813 1539
rect 830 1538 836 1539
rect 878 1538 885 1539
rect 902 1538 908 1539
rect 951 1538 957 1539
rect 966 1539 967 1540
rect 971 1539 972 1543
rect 1030 1543 1037 1544
rect 1030 1539 1031 1543
rect 1036 1539 1037 1543
rect 1366 1541 1372 1542
rect 966 1538 972 1539
rect 974 1538 980 1539
rect 1030 1538 1037 1539
rect 1054 1538 1060 1539
rect 278 1534 279 1538
rect 283 1534 284 1538
rect 278 1533 284 1534
rect 334 1534 335 1538
rect 339 1534 340 1538
rect 334 1533 340 1534
rect 398 1534 399 1538
rect 403 1534 404 1538
rect 398 1533 404 1534
rect 470 1534 471 1538
rect 475 1534 476 1538
rect 470 1533 476 1534
rect 542 1534 543 1538
rect 547 1534 548 1538
rect 542 1533 548 1534
rect 614 1534 615 1538
rect 619 1534 620 1538
rect 614 1533 620 1534
rect 686 1534 687 1538
rect 691 1534 692 1538
rect 686 1533 692 1534
rect 758 1534 759 1538
rect 763 1534 764 1538
rect 758 1533 764 1534
rect 830 1534 831 1538
rect 835 1534 836 1538
rect 830 1533 836 1534
rect 902 1534 903 1538
rect 907 1534 908 1538
rect 902 1533 908 1534
rect 974 1534 975 1538
rect 979 1534 980 1538
rect 974 1533 980 1534
rect 1054 1534 1055 1538
rect 1059 1534 1060 1538
rect 1366 1537 1367 1541
rect 1371 1537 1372 1541
rect 1366 1536 1372 1537
rect 2582 1541 2588 1542
rect 2582 1537 2583 1541
rect 2587 1537 2588 1541
rect 2582 1536 2588 1537
rect 1054 1533 1060 1534
rect 1902 1531 1908 1532
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 1326 1529 1332 1530
rect 1326 1525 1327 1529
rect 1331 1525 1332 1529
rect 1902 1527 1903 1531
rect 1907 1530 1908 1531
rect 2142 1531 2148 1532
rect 1907 1528 2027 1530
rect 1907 1527 1908 1528
rect 1902 1526 1908 1527
rect 1326 1524 1332 1525
rect 1366 1524 1372 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 254 1519 260 1520
rect 254 1515 255 1519
rect 259 1518 260 1519
rect 446 1519 452 1520
rect 259 1516 346 1518
rect 259 1515 260 1516
rect 254 1514 260 1515
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 262 1511 268 1512
rect 262 1507 263 1511
rect 267 1507 268 1511
rect 318 1511 324 1512
rect 262 1506 268 1507
rect 294 1507 301 1508
rect 294 1503 295 1507
rect 300 1503 301 1507
rect 318 1507 319 1511
rect 323 1507 324 1511
rect 318 1506 324 1507
rect 344 1506 346 1516
rect 446 1515 447 1519
rect 451 1518 452 1519
rect 734 1519 740 1520
rect 451 1516 626 1518
rect 451 1515 452 1516
rect 446 1514 452 1515
rect 382 1511 388 1512
rect 351 1507 357 1508
rect 351 1506 352 1507
rect 344 1504 352 1506
rect 294 1502 301 1503
rect 351 1503 352 1504
rect 356 1503 357 1507
rect 382 1507 383 1511
rect 387 1507 388 1511
rect 454 1511 460 1512
rect 382 1506 388 1507
rect 414 1507 421 1508
rect 351 1502 357 1503
rect 414 1503 415 1507
rect 420 1503 421 1507
rect 454 1507 455 1511
rect 459 1507 460 1511
rect 526 1511 532 1512
rect 454 1506 460 1507
rect 487 1507 496 1508
rect 414 1502 421 1503
rect 487 1503 488 1507
rect 495 1503 496 1507
rect 526 1507 527 1511
rect 531 1507 532 1511
rect 598 1511 604 1512
rect 526 1506 532 1507
rect 559 1507 565 1508
rect 487 1502 496 1503
rect 559 1503 560 1507
rect 564 1506 565 1507
rect 574 1507 580 1508
rect 574 1506 575 1507
rect 564 1504 575 1506
rect 564 1503 565 1504
rect 559 1502 565 1503
rect 574 1503 575 1504
rect 579 1503 580 1507
rect 598 1507 599 1511
rect 603 1507 604 1511
rect 598 1506 604 1507
rect 624 1506 626 1516
rect 734 1515 735 1519
rect 739 1518 740 1519
rect 878 1519 884 1520
rect 1366 1519 1372 1520
rect 1662 1523 1668 1524
rect 1662 1519 1663 1523
rect 1667 1519 1668 1523
rect 1718 1523 1724 1524
rect 739 1516 842 1518
rect 739 1515 740 1516
rect 734 1514 740 1515
rect 670 1511 676 1512
rect 631 1507 637 1508
rect 631 1506 632 1507
rect 624 1504 632 1506
rect 574 1502 580 1503
rect 631 1503 632 1504
rect 636 1503 637 1507
rect 670 1507 671 1511
rect 675 1507 676 1511
rect 742 1511 748 1512
rect 670 1506 676 1507
rect 703 1507 712 1508
rect 631 1502 637 1503
rect 703 1503 704 1507
rect 711 1503 712 1507
rect 742 1507 743 1511
rect 747 1507 748 1511
rect 814 1511 820 1512
rect 742 1506 748 1507
rect 775 1507 781 1508
rect 775 1506 776 1507
rect 703 1502 712 1503
rect 752 1504 776 1506
rect 678 1499 684 1500
rect 678 1495 679 1499
rect 683 1498 684 1499
rect 752 1498 754 1504
rect 775 1503 776 1504
rect 780 1503 781 1507
rect 814 1507 815 1511
rect 819 1507 820 1511
rect 814 1506 820 1507
rect 840 1506 842 1516
rect 878 1515 879 1519
rect 883 1518 884 1519
rect 1662 1518 1668 1519
rect 1695 1519 1701 1520
rect 883 1516 995 1518
rect 883 1515 884 1516
rect 878 1514 884 1515
rect 886 1511 892 1512
rect 847 1507 853 1508
rect 847 1506 848 1507
rect 840 1504 848 1506
rect 775 1502 781 1503
rect 847 1503 848 1504
rect 852 1503 853 1507
rect 886 1507 887 1511
rect 891 1507 892 1511
rect 958 1511 964 1512
rect 886 1506 892 1507
rect 910 1507 916 1508
rect 847 1502 853 1503
rect 910 1503 911 1507
rect 915 1506 916 1507
rect 919 1507 925 1508
rect 919 1506 920 1507
rect 915 1504 920 1506
rect 915 1503 916 1504
rect 910 1502 916 1503
rect 919 1503 920 1504
rect 924 1503 925 1507
rect 958 1507 959 1511
rect 963 1507 964 1511
rect 993 1508 995 1516
rect 1695 1515 1696 1519
rect 1700 1518 1701 1519
rect 1703 1519 1709 1520
rect 1703 1518 1704 1519
rect 1700 1516 1704 1518
rect 1700 1515 1701 1516
rect 1695 1514 1701 1515
rect 1703 1515 1704 1516
rect 1708 1515 1709 1519
rect 1718 1519 1719 1523
rect 1723 1519 1724 1523
rect 1774 1523 1780 1524
rect 1718 1518 1724 1519
rect 1751 1519 1760 1520
rect 1703 1514 1709 1515
rect 1751 1515 1752 1519
rect 1759 1515 1760 1519
rect 1774 1519 1775 1523
rect 1779 1519 1780 1523
rect 1838 1523 1844 1524
rect 1774 1518 1780 1519
rect 1807 1519 1816 1520
rect 1751 1514 1760 1515
rect 1807 1515 1808 1519
rect 1815 1515 1816 1519
rect 1838 1519 1839 1523
rect 1843 1519 1844 1523
rect 1910 1523 1916 1524
rect 1838 1518 1844 1519
rect 1871 1519 1880 1520
rect 1807 1514 1816 1515
rect 1871 1515 1872 1519
rect 1879 1515 1880 1519
rect 1910 1519 1911 1523
rect 1915 1519 1916 1523
rect 1990 1523 1996 1524
rect 1910 1518 1916 1519
rect 1943 1519 1952 1520
rect 1871 1514 1880 1515
rect 1943 1515 1944 1519
rect 1951 1515 1952 1519
rect 1990 1519 1991 1523
rect 1995 1519 1996 1523
rect 2025 1520 2027 1528
rect 2142 1527 2143 1531
rect 2147 1530 2148 1531
rect 2382 1531 2388 1532
rect 2147 1528 2258 1530
rect 2147 1527 2148 1528
rect 2142 1526 2148 1527
rect 2070 1523 2076 1524
rect 1990 1518 1996 1519
rect 2023 1519 2029 1520
rect 1943 1514 1952 1515
rect 2023 1515 2024 1519
rect 2028 1515 2029 1519
rect 2070 1519 2071 1523
rect 2075 1519 2076 1523
rect 2150 1523 2156 1524
rect 2070 1518 2076 1519
rect 2103 1519 2109 1520
rect 2103 1518 2104 1519
rect 2080 1516 2104 1518
rect 2023 1514 2029 1515
rect 2034 1515 2040 1516
rect 1326 1512 1332 1513
rect 1038 1511 1044 1512
rect 958 1506 964 1507
rect 991 1507 997 1508
rect 919 1502 925 1503
rect 991 1503 992 1507
rect 996 1503 997 1507
rect 1038 1507 1039 1511
rect 1043 1507 1044 1511
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 2034 1511 2035 1515
rect 2039 1514 2040 1515
rect 2080 1514 2082 1516
rect 2103 1515 2104 1516
rect 2108 1515 2109 1519
rect 2150 1519 2151 1523
rect 2155 1519 2156 1523
rect 2230 1523 2236 1524
rect 2150 1518 2156 1519
rect 2183 1519 2189 1520
rect 2103 1514 2109 1515
rect 2183 1515 2184 1519
rect 2188 1518 2189 1519
rect 2191 1519 2197 1520
rect 2191 1518 2192 1519
rect 2188 1516 2192 1518
rect 2188 1515 2189 1516
rect 2183 1514 2189 1515
rect 2191 1515 2192 1516
rect 2196 1515 2197 1519
rect 2230 1519 2231 1523
rect 2235 1519 2236 1523
rect 2230 1518 2236 1519
rect 2256 1518 2258 1528
rect 2382 1527 2383 1531
rect 2387 1530 2388 1531
rect 2387 1528 2498 1530
rect 2387 1527 2388 1528
rect 2382 1526 2388 1527
rect 2310 1523 2316 1524
rect 2263 1519 2269 1520
rect 2263 1518 2264 1519
rect 2256 1516 2264 1518
rect 2191 1514 2197 1515
rect 2263 1515 2264 1516
rect 2268 1515 2269 1519
rect 2310 1519 2311 1523
rect 2315 1519 2316 1523
rect 2390 1523 2396 1524
rect 2310 1518 2316 1519
rect 2342 1519 2349 1520
rect 2263 1514 2269 1515
rect 2342 1515 2343 1519
rect 2348 1515 2349 1519
rect 2390 1519 2391 1523
rect 2395 1519 2396 1523
rect 2470 1523 2476 1524
rect 2390 1518 2396 1519
rect 2414 1519 2420 1520
rect 2342 1514 2349 1515
rect 2414 1515 2415 1519
rect 2419 1518 2420 1519
rect 2423 1519 2429 1520
rect 2423 1518 2424 1519
rect 2419 1516 2424 1518
rect 2419 1515 2420 1516
rect 2414 1514 2420 1515
rect 2423 1515 2424 1516
rect 2428 1515 2429 1519
rect 2470 1519 2471 1523
rect 2475 1519 2476 1523
rect 2470 1518 2476 1519
rect 2496 1518 2498 1528
rect 2582 1524 2588 1525
rect 2526 1523 2532 1524
rect 2503 1519 2509 1520
rect 2503 1518 2504 1519
rect 2496 1516 2504 1518
rect 2423 1514 2429 1515
rect 2503 1515 2504 1516
rect 2508 1515 2509 1519
rect 2526 1519 2527 1523
rect 2531 1519 2532 1523
rect 2582 1520 2583 1524
rect 2587 1520 2588 1524
rect 2526 1518 2532 1519
rect 2558 1519 2565 1520
rect 2582 1519 2588 1520
rect 2503 1514 2509 1515
rect 2558 1515 2559 1519
rect 2564 1515 2565 1519
rect 2558 1514 2565 1515
rect 2039 1512 2082 1514
rect 2039 1511 2040 1512
rect 2034 1510 2040 1511
rect 1038 1506 1044 1507
rect 1071 1507 1077 1508
rect 1326 1507 1332 1508
rect 1071 1506 1072 1507
rect 991 1502 997 1503
rect 1048 1504 1072 1506
rect 683 1496 754 1498
rect 966 1499 972 1500
rect 683 1495 684 1496
rect 678 1494 684 1495
rect 966 1495 967 1499
rect 971 1498 972 1499
rect 1048 1498 1050 1504
rect 1071 1503 1072 1504
rect 1076 1503 1077 1507
rect 1071 1502 1077 1503
rect 971 1496 1050 1498
rect 971 1495 972 1496
rect 966 1494 972 1495
rect 1670 1491 1676 1492
rect 1670 1487 1671 1491
rect 1675 1490 1676 1491
rect 1675 1488 1931 1490
rect 1675 1487 1676 1488
rect 1670 1486 1676 1487
rect 1929 1484 1931 1488
rect 2282 1487 2288 1488
rect 1551 1483 1557 1484
rect 1518 1481 1524 1482
rect 1366 1480 1372 1481
rect 390 1479 396 1480
rect 231 1475 237 1476
rect 198 1473 204 1474
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 198 1469 199 1473
rect 203 1469 204 1473
rect 231 1471 232 1475
rect 236 1474 237 1475
rect 278 1475 284 1476
rect 278 1474 279 1475
rect 236 1472 279 1474
rect 236 1471 237 1472
rect 231 1470 237 1471
rect 278 1471 279 1472
rect 283 1471 284 1475
rect 319 1475 325 1476
rect 278 1470 284 1471
rect 286 1473 292 1474
rect 198 1468 204 1469
rect 286 1469 287 1473
rect 291 1469 292 1473
rect 319 1471 320 1475
rect 324 1474 325 1475
rect 374 1475 380 1476
rect 374 1474 375 1475
rect 324 1472 375 1474
rect 324 1471 325 1472
rect 319 1470 325 1471
rect 374 1471 375 1472
rect 379 1471 380 1475
rect 390 1475 391 1479
rect 395 1478 396 1479
rect 527 1479 533 1480
rect 395 1476 410 1478
rect 395 1475 396 1476
rect 390 1474 396 1475
rect 408 1474 410 1476
rect 415 1475 421 1476
rect 415 1474 416 1475
rect 374 1470 380 1471
rect 382 1473 388 1474
rect 286 1468 292 1469
rect 382 1469 383 1473
rect 387 1469 388 1473
rect 408 1472 416 1474
rect 415 1471 416 1472
rect 420 1471 421 1475
rect 510 1475 516 1476
rect 415 1470 421 1471
rect 486 1473 492 1474
rect 382 1468 388 1469
rect 486 1469 487 1473
rect 491 1469 492 1473
rect 510 1471 511 1475
rect 515 1474 516 1475
rect 519 1475 525 1476
rect 519 1474 520 1475
rect 515 1472 520 1474
rect 515 1471 516 1472
rect 510 1470 516 1471
rect 519 1471 520 1472
rect 524 1471 525 1475
rect 527 1475 528 1479
rect 532 1478 533 1479
rect 532 1476 619 1478
rect 1366 1476 1367 1480
rect 1371 1476 1372 1480
rect 1518 1477 1519 1481
rect 1523 1477 1524 1481
rect 1551 1479 1552 1483
rect 1556 1482 1557 1483
rect 1566 1483 1572 1484
rect 1566 1482 1567 1483
rect 1556 1480 1567 1482
rect 1556 1479 1557 1480
rect 1551 1478 1557 1479
rect 1566 1479 1567 1480
rect 1571 1479 1572 1483
rect 1607 1483 1613 1484
rect 1566 1478 1572 1479
rect 1574 1481 1580 1482
rect 1518 1476 1524 1477
rect 1574 1477 1575 1481
rect 1579 1477 1580 1481
rect 1607 1479 1608 1483
rect 1612 1482 1613 1483
rect 1638 1483 1644 1484
rect 1638 1482 1639 1483
rect 1612 1480 1639 1482
rect 1612 1479 1613 1480
rect 1607 1478 1613 1479
rect 1638 1479 1639 1480
rect 1643 1479 1644 1483
rect 1679 1483 1685 1484
rect 1638 1478 1644 1479
rect 1646 1481 1652 1482
rect 1574 1476 1580 1477
rect 1646 1477 1647 1481
rect 1651 1477 1652 1481
rect 1679 1479 1680 1483
rect 1684 1482 1685 1483
rect 1718 1483 1724 1484
rect 1718 1482 1719 1483
rect 1684 1480 1719 1482
rect 1684 1479 1685 1480
rect 1679 1478 1685 1479
rect 1718 1479 1719 1480
rect 1723 1479 1724 1483
rect 1759 1483 1765 1484
rect 1718 1478 1724 1479
rect 1726 1481 1732 1482
rect 1646 1476 1652 1477
rect 1726 1477 1727 1481
rect 1731 1477 1732 1481
rect 1759 1479 1760 1483
rect 1764 1482 1765 1483
rect 1798 1483 1804 1484
rect 1798 1482 1799 1483
rect 1764 1480 1799 1482
rect 1764 1479 1765 1480
rect 1759 1478 1765 1479
rect 1798 1479 1799 1480
rect 1803 1479 1804 1483
rect 1839 1483 1845 1484
rect 1798 1478 1804 1479
rect 1806 1481 1812 1482
rect 1726 1476 1732 1477
rect 1806 1477 1807 1481
rect 1811 1477 1812 1481
rect 1839 1479 1840 1483
rect 1844 1482 1845 1483
rect 1886 1483 1892 1484
rect 1886 1482 1887 1483
rect 1844 1480 1887 1482
rect 1844 1479 1845 1480
rect 1839 1478 1845 1479
rect 1886 1479 1887 1480
rect 1891 1479 1892 1483
rect 1927 1483 1933 1484
rect 1886 1478 1892 1479
rect 1894 1481 1900 1482
rect 1806 1476 1812 1477
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1927 1479 1928 1483
rect 1932 1479 1933 1483
rect 2006 1483 2012 1484
rect 1927 1478 1933 1479
rect 1982 1481 1988 1482
rect 1894 1476 1900 1477
rect 1982 1477 1983 1481
rect 1987 1477 1988 1481
rect 2006 1479 2007 1483
rect 2011 1482 2012 1483
rect 2015 1483 2021 1484
rect 2015 1482 2016 1483
rect 2011 1480 2016 1482
rect 2011 1479 2012 1480
rect 2006 1478 2012 1479
rect 2015 1479 2016 1480
rect 2020 1479 2021 1483
rect 2103 1483 2109 1484
rect 2015 1478 2021 1479
rect 2070 1481 2076 1482
rect 1982 1476 1988 1477
rect 2070 1477 2071 1481
rect 2075 1477 2076 1481
rect 2103 1479 2104 1483
rect 2108 1482 2109 1483
rect 2142 1483 2148 1484
rect 2142 1482 2143 1483
rect 2108 1480 2143 1482
rect 2108 1479 2109 1480
rect 2103 1478 2109 1479
rect 2142 1479 2143 1480
rect 2147 1479 2148 1483
rect 2183 1483 2189 1484
rect 2142 1478 2148 1479
rect 2150 1481 2156 1482
rect 2070 1476 2076 1477
rect 2150 1477 2151 1481
rect 2155 1477 2156 1481
rect 2183 1479 2184 1483
rect 2188 1482 2189 1483
rect 2222 1483 2228 1484
rect 2222 1482 2223 1483
rect 2188 1480 2223 1482
rect 2188 1479 2189 1480
rect 2183 1478 2189 1479
rect 2222 1479 2223 1480
rect 2227 1479 2228 1483
rect 2263 1483 2272 1484
rect 2222 1478 2228 1479
rect 2230 1481 2236 1482
rect 2150 1476 2156 1477
rect 2230 1477 2231 1481
rect 2235 1477 2236 1481
rect 2263 1479 2264 1483
rect 2271 1479 2272 1483
rect 2282 1483 2283 1487
rect 2287 1486 2288 1487
rect 2354 1487 2360 1488
rect 2287 1484 2347 1486
rect 2287 1483 2288 1484
rect 2282 1482 2288 1483
rect 2343 1483 2349 1484
rect 2263 1478 2272 1479
rect 2310 1481 2316 1482
rect 2230 1476 2236 1477
rect 2310 1477 2311 1481
rect 2315 1477 2316 1481
rect 2343 1479 2344 1483
rect 2348 1479 2349 1483
rect 2354 1483 2355 1487
rect 2359 1486 2360 1487
rect 2534 1487 2540 1488
rect 2359 1484 2418 1486
rect 2359 1483 2360 1484
rect 2354 1482 2360 1483
rect 2416 1482 2418 1484
rect 2423 1483 2429 1484
rect 2423 1482 2424 1483
rect 2343 1478 2349 1479
rect 2390 1481 2396 1482
rect 2310 1476 2316 1477
rect 2390 1477 2391 1481
rect 2395 1477 2396 1481
rect 2416 1480 2424 1482
rect 2423 1479 2424 1480
rect 2428 1479 2429 1483
rect 2503 1483 2509 1484
rect 2423 1478 2429 1479
rect 2470 1481 2476 1482
rect 2390 1476 2396 1477
rect 2470 1477 2471 1481
rect 2475 1477 2476 1481
rect 2503 1479 2504 1483
rect 2508 1482 2509 1483
rect 2518 1483 2524 1484
rect 2518 1482 2519 1483
rect 2508 1480 2519 1482
rect 2508 1479 2509 1480
rect 2503 1478 2509 1479
rect 2518 1479 2519 1480
rect 2523 1479 2524 1483
rect 2534 1483 2535 1487
rect 2539 1486 2540 1487
rect 2539 1484 2563 1486
rect 2539 1483 2540 1484
rect 2534 1482 2540 1483
rect 2559 1483 2565 1484
rect 2518 1478 2524 1479
rect 2526 1481 2532 1482
rect 2470 1476 2476 1477
rect 2526 1477 2527 1481
rect 2531 1477 2532 1481
rect 2559 1479 2560 1483
rect 2564 1479 2565 1483
rect 2559 1478 2565 1479
rect 2582 1480 2588 1481
rect 2526 1476 2532 1477
rect 2582 1476 2583 1480
rect 2587 1476 2588 1480
rect 532 1475 533 1476
rect 527 1474 533 1475
rect 615 1475 621 1476
rect 519 1470 525 1471
rect 582 1473 588 1474
rect 486 1468 492 1469
rect 582 1469 583 1473
rect 587 1469 588 1473
rect 615 1471 616 1475
rect 620 1471 621 1475
rect 711 1475 717 1476
rect 615 1470 621 1471
rect 678 1473 684 1474
rect 582 1468 588 1469
rect 678 1469 679 1473
rect 683 1469 684 1473
rect 711 1471 712 1475
rect 716 1474 717 1475
rect 766 1475 772 1476
rect 766 1474 767 1475
rect 716 1472 767 1474
rect 716 1471 717 1472
rect 711 1470 717 1471
rect 766 1471 767 1472
rect 771 1471 772 1475
rect 806 1475 813 1476
rect 766 1470 772 1471
rect 774 1473 780 1474
rect 678 1468 684 1469
rect 774 1469 775 1473
rect 779 1469 780 1473
rect 806 1471 807 1475
rect 812 1471 813 1475
rect 895 1475 901 1476
rect 806 1470 813 1471
rect 862 1473 868 1474
rect 774 1468 780 1469
rect 862 1469 863 1473
rect 867 1469 868 1473
rect 895 1471 896 1475
rect 900 1474 901 1475
rect 942 1475 948 1476
rect 942 1474 943 1475
rect 900 1472 943 1474
rect 900 1471 901 1472
rect 895 1470 901 1471
rect 942 1471 943 1472
rect 947 1471 948 1475
rect 983 1475 989 1476
rect 942 1470 948 1471
rect 950 1473 956 1474
rect 862 1468 868 1469
rect 950 1469 951 1473
rect 955 1469 956 1473
rect 983 1471 984 1475
rect 988 1474 989 1475
rect 1030 1475 1036 1476
rect 1030 1474 1031 1475
rect 988 1472 1031 1474
rect 988 1471 989 1472
rect 983 1470 989 1471
rect 1030 1471 1031 1472
rect 1035 1471 1036 1475
rect 1071 1475 1077 1476
rect 1030 1470 1036 1471
rect 1038 1473 1044 1474
rect 950 1468 956 1469
rect 1038 1469 1039 1473
rect 1043 1469 1044 1473
rect 1071 1471 1072 1475
rect 1076 1474 1077 1475
rect 1126 1475 1132 1476
rect 1126 1474 1127 1475
rect 1076 1472 1127 1474
rect 1076 1471 1077 1472
rect 1071 1470 1077 1471
rect 1126 1471 1127 1472
rect 1131 1471 1132 1475
rect 1167 1475 1173 1476
rect 1126 1470 1132 1471
rect 1134 1473 1140 1474
rect 1038 1468 1044 1469
rect 1134 1469 1135 1473
rect 1139 1469 1140 1473
rect 1167 1471 1168 1475
rect 1172 1474 1173 1475
rect 1190 1475 1196 1476
rect 1366 1475 1372 1476
rect 2582 1475 2588 1476
rect 1190 1474 1191 1475
rect 1172 1472 1191 1474
rect 1172 1471 1173 1472
rect 1167 1470 1173 1471
rect 1190 1471 1191 1472
rect 1195 1471 1196 1475
rect 1190 1470 1196 1471
rect 1326 1472 1332 1473
rect 1134 1468 1140 1469
rect 1326 1468 1327 1472
rect 1331 1468 1332 1472
rect 110 1467 116 1468
rect 1326 1467 1332 1468
rect 1366 1463 1372 1464
rect 1366 1459 1367 1463
rect 1371 1459 1372 1463
rect 1366 1458 1372 1459
rect 2582 1463 2588 1464
rect 2582 1459 2583 1463
rect 2587 1459 2588 1463
rect 2582 1458 2588 1459
rect 110 1455 116 1456
rect 110 1451 111 1455
rect 115 1451 116 1455
rect 110 1450 116 1451
rect 1326 1455 1332 1456
rect 1326 1451 1327 1455
rect 1331 1451 1332 1455
rect 1326 1450 1332 1451
rect 1534 1454 1540 1455
rect 1534 1450 1535 1454
rect 1539 1450 1540 1454
rect 1534 1449 1540 1450
rect 1590 1454 1596 1455
rect 1590 1450 1591 1454
rect 1595 1450 1596 1454
rect 1590 1449 1596 1450
rect 1662 1454 1668 1455
rect 1662 1450 1663 1454
rect 1667 1450 1668 1454
rect 1662 1449 1668 1450
rect 1742 1454 1748 1455
rect 1742 1450 1743 1454
rect 1747 1450 1748 1454
rect 1742 1449 1748 1450
rect 1822 1454 1828 1455
rect 1822 1450 1823 1454
rect 1827 1450 1828 1454
rect 1822 1449 1828 1450
rect 1910 1454 1916 1455
rect 1910 1450 1911 1454
rect 1915 1450 1916 1454
rect 1910 1449 1916 1450
rect 1998 1454 2004 1455
rect 1998 1450 1999 1454
rect 2003 1450 2004 1454
rect 1998 1449 2004 1450
rect 2086 1454 2092 1455
rect 2086 1450 2087 1454
rect 2091 1450 2092 1454
rect 2086 1449 2092 1450
rect 2166 1454 2172 1455
rect 2166 1450 2167 1454
rect 2171 1450 2172 1454
rect 2166 1449 2172 1450
rect 2246 1454 2252 1455
rect 2246 1450 2247 1454
rect 2251 1450 2252 1454
rect 2246 1449 2252 1450
rect 2326 1454 2332 1455
rect 2326 1450 2327 1454
rect 2331 1450 2332 1454
rect 2326 1449 2332 1450
rect 2406 1454 2412 1455
rect 2406 1450 2407 1454
rect 2411 1450 2412 1454
rect 2406 1449 2412 1450
rect 2486 1454 2492 1455
rect 2486 1450 2487 1454
rect 2491 1450 2492 1454
rect 2486 1449 2492 1450
rect 2542 1454 2548 1455
rect 2542 1450 2543 1454
rect 2547 1450 2548 1454
rect 2542 1449 2548 1450
rect 1511 1447 1517 1448
rect 214 1446 220 1447
rect 214 1442 215 1446
rect 219 1442 220 1446
rect 214 1441 220 1442
rect 302 1446 308 1447
rect 302 1442 303 1446
rect 307 1442 308 1446
rect 302 1441 308 1442
rect 398 1446 404 1447
rect 398 1442 399 1446
rect 403 1442 404 1446
rect 398 1441 404 1442
rect 502 1446 508 1447
rect 502 1442 503 1446
rect 507 1442 508 1446
rect 502 1441 508 1442
rect 598 1446 604 1447
rect 598 1442 599 1446
rect 603 1442 604 1446
rect 598 1441 604 1442
rect 694 1446 700 1447
rect 694 1442 695 1446
rect 699 1442 700 1446
rect 694 1441 700 1442
rect 790 1446 796 1447
rect 790 1442 791 1446
rect 795 1442 796 1446
rect 790 1441 796 1442
rect 878 1446 884 1447
rect 878 1442 879 1446
rect 883 1442 884 1446
rect 878 1441 884 1442
rect 966 1446 972 1447
rect 966 1442 967 1446
rect 971 1442 972 1446
rect 966 1441 972 1442
rect 1054 1446 1060 1447
rect 1054 1442 1055 1446
rect 1059 1442 1060 1446
rect 1054 1441 1060 1442
rect 1150 1446 1156 1447
rect 1150 1442 1151 1446
rect 1155 1442 1156 1446
rect 1511 1443 1512 1447
rect 1516 1446 1517 1447
rect 1566 1447 1573 1448
rect 1516 1444 1562 1446
rect 1516 1443 1517 1444
rect 1511 1442 1517 1443
rect 1150 1441 1156 1442
rect 174 1439 180 1440
rect 174 1435 175 1439
rect 179 1438 180 1439
rect 191 1439 197 1440
rect 191 1438 192 1439
rect 179 1436 192 1438
rect 179 1435 180 1436
rect 174 1434 180 1435
rect 191 1435 192 1436
rect 196 1435 197 1439
rect 191 1434 197 1435
rect 278 1439 285 1440
rect 278 1435 279 1439
rect 284 1435 285 1439
rect 278 1434 285 1435
rect 374 1439 381 1440
rect 374 1435 375 1439
rect 380 1435 381 1439
rect 374 1434 381 1435
rect 479 1439 485 1440
rect 479 1435 480 1439
rect 484 1438 485 1439
rect 527 1439 533 1440
rect 527 1438 528 1439
rect 484 1436 528 1438
rect 484 1435 485 1436
rect 479 1434 485 1435
rect 527 1435 528 1436
rect 532 1435 533 1439
rect 527 1434 533 1435
rect 574 1439 581 1440
rect 574 1435 575 1439
rect 580 1435 581 1439
rect 574 1434 581 1435
rect 671 1439 677 1440
rect 671 1435 672 1439
rect 676 1438 677 1439
rect 758 1439 764 1440
rect 758 1438 759 1439
rect 676 1436 759 1438
rect 676 1435 677 1436
rect 671 1434 677 1435
rect 758 1435 759 1436
rect 763 1435 764 1439
rect 758 1434 764 1435
rect 766 1439 773 1440
rect 766 1435 767 1439
rect 772 1435 773 1439
rect 766 1434 773 1435
rect 855 1439 861 1440
rect 855 1435 856 1439
rect 860 1438 861 1439
rect 910 1439 916 1440
rect 910 1438 911 1439
rect 860 1436 911 1438
rect 860 1435 861 1436
rect 855 1434 861 1435
rect 910 1435 911 1436
rect 915 1435 916 1439
rect 910 1434 916 1435
rect 942 1439 949 1440
rect 942 1435 943 1439
rect 948 1435 949 1439
rect 942 1434 949 1435
rect 1030 1439 1037 1440
rect 1030 1435 1031 1439
rect 1036 1435 1037 1439
rect 1030 1434 1037 1435
rect 1126 1439 1133 1440
rect 1126 1435 1127 1439
rect 1132 1435 1133 1439
rect 1560 1438 1562 1444
rect 1566 1443 1567 1447
rect 1572 1443 1573 1447
rect 1566 1442 1573 1443
rect 1638 1447 1645 1448
rect 1638 1443 1639 1447
rect 1644 1443 1645 1447
rect 1638 1442 1645 1443
rect 1718 1447 1725 1448
rect 1718 1443 1719 1447
rect 1724 1443 1725 1447
rect 1718 1442 1725 1443
rect 1798 1447 1805 1448
rect 1798 1443 1799 1447
rect 1804 1443 1805 1447
rect 1798 1442 1805 1443
rect 1886 1447 1893 1448
rect 1886 1443 1887 1447
rect 1892 1443 1893 1447
rect 1886 1442 1893 1443
rect 1975 1447 1981 1448
rect 1975 1443 1976 1447
rect 1980 1446 1981 1447
rect 2034 1447 2040 1448
rect 2034 1446 2035 1447
rect 1980 1444 2035 1446
rect 1980 1443 1981 1444
rect 1975 1442 1981 1443
rect 2034 1443 2035 1444
rect 2039 1443 2040 1447
rect 2034 1442 2040 1443
rect 2042 1447 2048 1448
rect 2042 1443 2043 1447
rect 2047 1446 2048 1447
rect 2063 1447 2069 1448
rect 2063 1446 2064 1447
rect 2047 1444 2064 1446
rect 2047 1443 2048 1444
rect 2042 1442 2048 1443
rect 2063 1443 2064 1444
rect 2068 1443 2069 1447
rect 2063 1442 2069 1443
rect 2142 1447 2149 1448
rect 2142 1443 2143 1447
rect 2148 1443 2149 1447
rect 2142 1442 2149 1443
rect 2222 1447 2229 1448
rect 2222 1443 2223 1447
rect 2228 1443 2229 1447
rect 2222 1442 2229 1443
rect 2303 1447 2309 1448
rect 2303 1443 2304 1447
rect 2308 1446 2309 1447
rect 2354 1447 2360 1448
rect 2354 1446 2355 1447
rect 2308 1444 2355 1446
rect 2308 1443 2309 1444
rect 2303 1442 2309 1443
rect 2354 1443 2355 1444
rect 2359 1443 2360 1447
rect 2354 1442 2360 1443
rect 2383 1447 2389 1448
rect 2383 1443 2384 1447
rect 2388 1446 2389 1447
rect 2414 1447 2420 1448
rect 2414 1446 2415 1447
rect 2388 1444 2415 1446
rect 2388 1443 2389 1444
rect 2383 1442 2389 1443
rect 2414 1443 2415 1444
rect 2419 1443 2420 1447
rect 2414 1442 2420 1443
rect 2463 1447 2469 1448
rect 2463 1443 2464 1447
rect 2468 1443 2469 1447
rect 2463 1442 2469 1443
rect 2518 1447 2525 1448
rect 2518 1443 2519 1447
rect 2524 1443 2525 1447
rect 2518 1442 2525 1443
rect 1838 1439 1844 1440
rect 1838 1438 1839 1439
rect 1560 1436 1839 1438
rect 1126 1434 1133 1435
rect 1838 1435 1839 1436
rect 1843 1435 1844 1439
rect 2465 1438 2467 1442
rect 2558 1439 2564 1440
rect 2558 1438 2559 1439
rect 2465 1436 2559 1438
rect 1838 1434 1844 1435
rect 2006 1435 2012 1436
rect 2006 1434 2007 1435
rect 1916 1432 2007 1434
rect 358 1431 364 1432
rect 358 1430 359 1431
rect 240 1428 359 1430
rect 134 1423 141 1424
rect 134 1419 135 1423
rect 140 1419 141 1423
rect 223 1423 229 1424
rect 223 1419 224 1423
rect 228 1422 229 1423
rect 240 1422 242 1428
rect 358 1427 359 1428
rect 363 1427 364 1431
rect 510 1431 516 1432
rect 510 1430 511 1431
rect 358 1426 364 1427
rect 441 1428 511 1430
rect 228 1420 242 1422
rect 319 1423 325 1424
rect 228 1419 229 1420
rect 319 1419 320 1423
rect 324 1422 325 1423
rect 334 1423 340 1424
rect 334 1422 335 1423
rect 324 1420 335 1422
rect 324 1419 325 1420
rect 134 1418 141 1419
rect 158 1418 164 1419
rect 223 1418 229 1419
rect 246 1418 252 1419
rect 319 1418 325 1419
rect 334 1419 335 1420
rect 339 1419 340 1423
rect 423 1423 429 1424
rect 423 1419 424 1423
rect 428 1422 429 1423
rect 441 1422 443 1428
rect 510 1427 511 1428
rect 515 1427 516 1431
rect 1118 1431 1124 1432
rect 1118 1430 1119 1431
rect 510 1426 516 1427
rect 984 1428 1119 1430
rect 428 1420 443 1422
rect 466 1423 472 1424
rect 428 1419 429 1420
rect 466 1419 467 1423
rect 471 1422 472 1423
rect 527 1423 533 1424
rect 527 1422 528 1423
rect 471 1420 528 1422
rect 471 1419 472 1420
rect 334 1418 340 1419
rect 342 1418 348 1419
rect 423 1418 429 1419
rect 446 1418 452 1419
rect 466 1418 472 1419
rect 527 1419 528 1420
rect 532 1419 533 1423
rect 570 1423 576 1424
rect 570 1419 571 1423
rect 575 1422 576 1423
rect 639 1423 645 1424
rect 639 1422 640 1423
rect 575 1420 640 1422
rect 575 1419 576 1420
rect 527 1418 533 1419
rect 550 1418 556 1419
rect 570 1418 576 1419
rect 639 1419 640 1420
rect 644 1419 645 1423
rect 742 1423 749 1424
rect 742 1419 743 1423
rect 748 1419 749 1423
rect 855 1423 861 1424
rect 855 1419 856 1423
rect 860 1422 861 1423
rect 870 1423 876 1424
rect 870 1422 871 1423
rect 860 1420 871 1422
rect 860 1419 861 1420
rect 639 1418 645 1419
rect 662 1418 668 1419
rect 742 1418 749 1419
rect 766 1418 772 1419
rect 855 1418 861 1419
rect 870 1419 871 1420
rect 875 1419 876 1423
rect 967 1423 973 1424
rect 967 1419 968 1423
rect 972 1422 973 1423
rect 984 1422 986 1428
rect 1118 1427 1119 1428
rect 1123 1427 1124 1431
rect 1118 1426 1124 1427
rect 1391 1427 1397 1428
rect 972 1420 986 1422
rect 1078 1423 1085 1424
rect 972 1419 973 1420
rect 1078 1419 1079 1423
rect 1084 1419 1085 1423
rect 1190 1423 1197 1424
rect 1190 1419 1191 1423
rect 1196 1419 1197 1423
rect 1391 1423 1392 1427
rect 1396 1426 1397 1427
rect 1406 1427 1412 1428
rect 1406 1426 1407 1427
rect 1396 1424 1407 1426
rect 1396 1423 1397 1424
rect 1391 1422 1397 1423
rect 1406 1423 1407 1424
rect 1411 1423 1412 1427
rect 1434 1427 1440 1428
rect 1434 1423 1435 1427
rect 1439 1426 1440 1427
rect 1447 1427 1453 1428
rect 1447 1426 1448 1427
rect 1439 1424 1448 1426
rect 1439 1423 1440 1424
rect 1406 1422 1412 1423
rect 1414 1422 1420 1423
rect 1434 1422 1440 1423
rect 1447 1423 1448 1424
rect 1452 1423 1453 1427
rect 1502 1427 1508 1428
rect 1502 1423 1503 1427
rect 1507 1426 1508 1427
rect 1511 1427 1517 1428
rect 1511 1426 1512 1427
rect 1507 1424 1512 1426
rect 1507 1423 1508 1424
rect 1447 1422 1453 1423
rect 1470 1422 1476 1423
rect 1502 1422 1508 1423
rect 1511 1423 1512 1424
rect 1516 1423 1517 1427
rect 1554 1427 1560 1428
rect 1554 1423 1555 1427
rect 1559 1426 1560 1427
rect 1599 1427 1605 1428
rect 1599 1426 1600 1427
rect 1559 1424 1600 1426
rect 1559 1423 1560 1424
rect 1511 1422 1517 1423
rect 1534 1422 1540 1423
rect 1554 1422 1560 1423
rect 1599 1423 1600 1424
rect 1604 1423 1605 1427
rect 1642 1427 1648 1428
rect 1642 1423 1643 1427
rect 1647 1426 1648 1427
rect 1695 1427 1701 1428
rect 1695 1426 1696 1427
rect 1647 1424 1696 1426
rect 1647 1423 1648 1424
rect 1599 1422 1605 1423
rect 1622 1422 1628 1423
rect 1642 1422 1648 1423
rect 1695 1423 1696 1424
rect 1700 1423 1701 1427
rect 1743 1427 1749 1428
rect 1743 1423 1744 1427
rect 1748 1426 1749 1427
rect 1799 1427 1805 1428
rect 1799 1426 1800 1427
rect 1748 1424 1800 1426
rect 1748 1423 1749 1424
rect 1695 1422 1701 1423
rect 1718 1422 1724 1423
rect 1743 1422 1749 1423
rect 1799 1423 1800 1424
rect 1804 1423 1805 1427
rect 1903 1427 1909 1428
rect 1903 1423 1904 1427
rect 1908 1426 1909 1427
rect 1916 1426 1918 1432
rect 2006 1431 2007 1432
rect 2011 1431 2012 1435
rect 2134 1435 2140 1436
rect 2134 1434 2135 1435
rect 2006 1430 2012 1431
rect 2016 1432 2135 1434
rect 1908 1424 1918 1426
rect 1999 1427 2005 1428
rect 1908 1423 1909 1424
rect 1999 1423 2000 1427
rect 2004 1426 2005 1427
rect 2016 1426 2018 1432
rect 2134 1431 2135 1432
rect 2139 1431 2140 1435
rect 2558 1435 2559 1436
rect 2563 1435 2564 1439
rect 2558 1434 2564 1435
rect 2134 1430 2140 1431
rect 2238 1431 2244 1432
rect 2238 1430 2239 1431
rect 2208 1428 2239 1430
rect 2004 1424 2018 1426
rect 2094 1427 2101 1428
rect 2004 1423 2005 1424
rect 2094 1423 2095 1427
rect 2100 1423 2101 1427
rect 2191 1427 2197 1428
rect 2191 1423 2192 1427
rect 2196 1426 2197 1427
rect 2208 1426 2210 1428
rect 2238 1427 2239 1428
rect 2243 1427 2244 1431
rect 2238 1426 2244 1427
rect 2279 1427 2288 1428
rect 2196 1424 2210 1426
rect 2196 1423 2197 1424
rect 2279 1423 2280 1427
rect 2287 1423 2288 1427
rect 2327 1427 2333 1428
rect 2327 1423 2328 1427
rect 2332 1426 2333 1427
rect 2367 1427 2373 1428
rect 2367 1426 2368 1427
rect 2332 1424 2368 1426
rect 2332 1423 2333 1424
rect 1799 1422 1805 1423
rect 1822 1422 1828 1423
rect 1903 1422 1909 1423
rect 1926 1422 1932 1423
rect 1999 1422 2005 1423
rect 2022 1422 2028 1423
rect 2094 1422 2101 1423
rect 2118 1422 2124 1423
rect 2191 1422 2197 1423
rect 2214 1422 2220 1423
rect 2279 1422 2288 1423
rect 2302 1422 2308 1423
rect 2327 1422 2333 1423
rect 2367 1423 2368 1424
rect 2372 1423 2373 1427
rect 2415 1427 2421 1428
rect 2415 1423 2416 1427
rect 2420 1426 2421 1427
rect 2455 1427 2461 1428
rect 2455 1426 2456 1427
rect 2420 1424 2456 1426
rect 2420 1423 2421 1424
rect 2367 1422 2373 1423
rect 2390 1422 2396 1423
rect 2415 1422 2421 1423
rect 2455 1423 2456 1424
rect 2460 1423 2461 1427
rect 2506 1427 2512 1428
rect 2506 1423 2507 1427
rect 2511 1426 2512 1427
rect 2519 1427 2525 1428
rect 2519 1426 2520 1427
rect 2511 1424 2520 1426
rect 2511 1423 2512 1424
rect 2455 1422 2461 1423
rect 2478 1422 2484 1423
rect 2506 1422 2512 1423
rect 2519 1423 2520 1424
rect 2524 1423 2525 1427
rect 2519 1422 2525 1423
rect 2542 1422 2548 1423
rect 870 1418 876 1419
rect 878 1418 884 1419
rect 967 1418 973 1419
rect 990 1418 996 1419
rect 1078 1418 1085 1419
rect 1102 1418 1108 1419
rect 1190 1418 1197 1419
rect 1214 1418 1220 1419
rect 158 1414 159 1418
rect 163 1414 164 1418
rect 158 1413 164 1414
rect 246 1414 247 1418
rect 251 1414 252 1418
rect 246 1413 252 1414
rect 342 1414 343 1418
rect 347 1414 348 1418
rect 342 1413 348 1414
rect 446 1414 447 1418
rect 451 1414 452 1418
rect 446 1413 452 1414
rect 550 1414 551 1418
rect 555 1414 556 1418
rect 550 1413 556 1414
rect 662 1414 663 1418
rect 667 1414 668 1418
rect 662 1413 668 1414
rect 766 1414 767 1418
rect 771 1414 772 1418
rect 766 1413 772 1414
rect 878 1414 879 1418
rect 883 1414 884 1418
rect 878 1413 884 1414
rect 990 1414 991 1418
rect 995 1414 996 1418
rect 990 1413 996 1414
rect 1102 1414 1103 1418
rect 1107 1414 1108 1418
rect 1102 1413 1108 1414
rect 1214 1414 1215 1418
rect 1219 1414 1220 1418
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1414 1417 1420 1418
rect 1470 1418 1471 1422
rect 1475 1418 1476 1422
rect 1470 1417 1476 1418
rect 1534 1418 1535 1422
rect 1539 1418 1540 1422
rect 1534 1417 1540 1418
rect 1622 1418 1623 1422
rect 1627 1418 1628 1422
rect 1622 1417 1628 1418
rect 1718 1418 1719 1422
rect 1723 1418 1724 1422
rect 1718 1417 1724 1418
rect 1822 1418 1823 1422
rect 1827 1418 1828 1422
rect 1822 1417 1828 1418
rect 1926 1418 1927 1422
rect 1931 1418 1932 1422
rect 1926 1417 1932 1418
rect 2022 1418 2023 1422
rect 2027 1418 2028 1422
rect 2022 1417 2028 1418
rect 2118 1418 2119 1422
rect 2123 1418 2124 1422
rect 2118 1417 2124 1418
rect 2214 1418 2215 1422
rect 2219 1418 2220 1422
rect 2214 1417 2220 1418
rect 2302 1418 2303 1422
rect 2307 1418 2308 1422
rect 2302 1417 2308 1418
rect 2390 1418 2391 1422
rect 2395 1418 2396 1422
rect 2390 1417 2396 1418
rect 2478 1418 2479 1422
rect 2483 1418 2484 1422
rect 2478 1417 2484 1418
rect 2542 1418 2543 1422
rect 2547 1418 2548 1422
rect 2542 1417 2548 1418
rect 1214 1413 1220 1414
rect 1366 1413 1372 1414
rect 110 1409 116 1410
rect 110 1405 111 1409
rect 115 1405 116 1409
rect 110 1404 116 1405
rect 1326 1409 1332 1410
rect 1326 1405 1327 1409
rect 1331 1405 1332 1409
rect 1366 1409 1367 1413
rect 1371 1409 1372 1413
rect 1366 1408 1372 1409
rect 2582 1413 2588 1414
rect 2582 1409 2583 1413
rect 2587 1409 2588 1413
rect 2582 1408 2588 1409
rect 1326 1404 1332 1405
rect 2094 1403 2100 1404
rect 134 1399 140 1400
rect 134 1395 135 1399
rect 139 1398 140 1399
rect 742 1399 748 1400
rect 139 1396 258 1398
rect 139 1395 140 1396
rect 134 1394 140 1395
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 142 1391 148 1392
rect 142 1387 143 1391
rect 147 1387 148 1391
rect 230 1391 236 1392
rect 142 1386 148 1387
rect 174 1387 181 1388
rect 174 1383 175 1387
rect 180 1383 181 1387
rect 230 1387 231 1391
rect 235 1387 236 1391
rect 230 1386 236 1387
rect 256 1386 258 1396
rect 742 1395 743 1399
rect 747 1398 748 1399
rect 1078 1399 1084 1400
rect 747 1396 890 1398
rect 747 1395 748 1396
rect 742 1394 748 1395
rect 326 1391 332 1392
rect 263 1387 269 1388
rect 263 1386 264 1387
rect 256 1384 264 1386
rect 174 1382 181 1383
rect 263 1383 264 1384
rect 268 1383 269 1387
rect 326 1387 327 1391
rect 331 1387 332 1391
rect 430 1391 436 1392
rect 326 1386 332 1387
rect 358 1387 365 1388
rect 263 1382 269 1383
rect 358 1383 359 1387
rect 364 1383 365 1387
rect 430 1387 431 1391
rect 435 1387 436 1391
rect 534 1391 540 1392
rect 430 1386 436 1387
rect 463 1387 472 1388
rect 358 1382 365 1383
rect 463 1383 464 1387
rect 471 1383 472 1387
rect 534 1387 535 1391
rect 539 1387 540 1391
rect 646 1391 652 1392
rect 534 1386 540 1387
rect 567 1387 576 1388
rect 463 1382 472 1383
rect 567 1383 568 1387
rect 575 1383 576 1387
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 750 1391 756 1392
rect 646 1386 652 1387
rect 670 1387 676 1388
rect 567 1382 576 1383
rect 670 1383 671 1387
rect 675 1386 676 1387
rect 679 1387 685 1388
rect 679 1386 680 1387
rect 675 1384 680 1386
rect 675 1383 676 1384
rect 670 1382 676 1383
rect 679 1383 680 1384
rect 684 1383 685 1387
rect 750 1387 751 1391
rect 755 1387 756 1391
rect 862 1391 868 1392
rect 750 1386 756 1387
rect 783 1387 789 1388
rect 679 1382 685 1383
rect 758 1383 764 1384
rect 758 1379 759 1383
rect 763 1382 764 1383
rect 783 1383 784 1387
rect 788 1383 789 1387
rect 862 1387 863 1391
rect 867 1387 868 1391
rect 862 1386 868 1387
rect 888 1386 890 1396
rect 1078 1395 1079 1399
rect 1083 1398 1084 1399
rect 2094 1399 2095 1403
rect 2099 1402 2100 1403
rect 2099 1400 2235 1402
rect 2099 1399 2100 1400
rect 2094 1398 2100 1399
rect 1083 1396 1226 1398
rect 1083 1395 1084 1396
rect 1078 1394 1084 1395
rect 974 1391 980 1392
rect 895 1387 901 1388
rect 895 1386 896 1387
rect 888 1384 896 1386
rect 783 1382 789 1383
rect 895 1383 896 1384
rect 900 1383 901 1387
rect 974 1387 975 1391
rect 979 1387 980 1391
rect 1086 1391 1092 1392
rect 974 1386 980 1387
rect 998 1387 1004 1388
rect 895 1382 901 1383
rect 998 1383 999 1387
rect 1003 1386 1004 1387
rect 1007 1387 1013 1388
rect 1007 1386 1008 1387
rect 1003 1384 1008 1386
rect 1003 1383 1004 1384
rect 998 1382 1004 1383
rect 1007 1383 1008 1384
rect 1012 1383 1013 1387
rect 1086 1387 1087 1391
rect 1091 1387 1092 1391
rect 1198 1391 1204 1392
rect 1086 1386 1092 1387
rect 1118 1387 1125 1388
rect 1007 1382 1013 1383
rect 1118 1383 1119 1387
rect 1124 1383 1125 1387
rect 1198 1387 1199 1391
rect 1203 1387 1204 1391
rect 1198 1386 1204 1387
rect 1224 1386 1226 1396
rect 1366 1396 1372 1397
rect 1326 1392 1332 1393
rect 1326 1388 1327 1392
rect 1331 1388 1332 1392
rect 1366 1392 1367 1396
rect 1371 1392 1372 1396
rect 1366 1391 1372 1392
rect 1398 1395 1404 1396
rect 1398 1391 1399 1395
rect 1403 1391 1404 1395
rect 1454 1395 1460 1396
rect 1398 1390 1404 1391
rect 1431 1391 1440 1392
rect 1231 1387 1237 1388
rect 1326 1387 1332 1388
rect 1431 1387 1432 1391
rect 1439 1387 1440 1391
rect 1454 1391 1455 1395
rect 1459 1391 1460 1395
rect 1518 1395 1524 1396
rect 1454 1390 1460 1391
rect 1487 1391 1493 1392
rect 1231 1386 1232 1387
rect 1224 1384 1232 1386
rect 1118 1382 1125 1383
rect 1231 1383 1232 1384
rect 1236 1383 1237 1387
rect 1431 1386 1440 1387
rect 1487 1387 1488 1391
rect 1492 1390 1493 1391
rect 1502 1391 1508 1392
rect 1502 1390 1503 1391
rect 1492 1388 1503 1390
rect 1492 1387 1493 1388
rect 1487 1386 1493 1387
rect 1502 1387 1503 1388
rect 1507 1387 1508 1391
rect 1518 1391 1519 1395
rect 1523 1391 1524 1395
rect 1606 1395 1612 1396
rect 1518 1390 1524 1391
rect 1551 1391 1560 1392
rect 1502 1386 1508 1387
rect 1551 1387 1552 1391
rect 1559 1387 1560 1391
rect 1606 1391 1607 1395
rect 1611 1391 1612 1395
rect 1702 1395 1708 1396
rect 1606 1390 1612 1391
rect 1639 1391 1648 1392
rect 1551 1386 1560 1387
rect 1639 1387 1640 1391
rect 1647 1387 1648 1391
rect 1702 1391 1703 1395
rect 1707 1391 1708 1395
rect 1806 1395 1812 1396
rect 1702 1390 1708 1391
rect 1735 1391 1741 1392
rect 1639 1386 1648 1387
rect 1735 1387 1736 1391
rect 1740 1390 1741 1391
rect 1743 1391 1749 1392
rect 1743 1390 1744 1391
rect 1740 1388 1744 1390
rect 1740 1387 1741 1388
rect 1735 1386 1741 1387
rect 1743 1387 1744 1388
rect 1748 1387 1749 1391
rect 1806 1391 1807 1395
rect 1811 1391 1812 1395
rect 1910 1395 1916 1396
rect 1806 1390 1812 1391
rect 1838 1391 1845 1392
rect 1743 1386 1749 1387
rect 1838 1387 1839 1391
rect 1844 1387 1845 1391
rect 1910 1391 1911 1395
rect 1915 1391 1916 1395
rect 2006 1395 2012 1396
rect 1910 1390 1916 1391
rect 1934 1391 1940 1392
rect 1838 1386 1845 1387
rect 1934 1387 1935 1391
rect 1939 1390 1940 1391
rect 1943 1391 1949 1392
rect 1943 1390 1944 1391
rect 1939 1388 1944 1390
rect 1939 1387 1940 1388
rect 1934 1386 1940 1387
rect 1943 1387 1944 1388
rect 1948 1387 1949 1391
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2102 1395 2108 1396
rect 2006 1390 2012 1391
rect 2039 1391 2048 1392
rect 1943 1386 1949 1387
rect 2039 1387 2040 1391
rect 2047 1387 2048 1391
rect 2102 1391 2103 1395
rect 2107 1391 2108 1395
rect 2198 1395 2204 1396
rect 2102 1390 2108 1391
rect 2134 1391 2141 1392
rect 2039 1386 2048 1387
rect 2134 1387 2135 1391
rect 2140 1387 2141 1391
rect 2198 1391 2199 1395
rect 2203 1391 2204 1395
rect 2233 1392 2235 1400
rect 2582 1396 2588 1397
rect 2286 1395 2292 1396
rect 2198 1390 2204 1391
rect 2231 1391 2237 1392
rect 2134 1386 2141 1387
rect 2231 1387 2232 1391
rect 2236 1387 2237 1391
rect 2286 1391 2287 1395
rect 2291 1391 2292 1395
rect 2374 1395 2380 1396
rect 2286 1390 2292 1391
rect 2319 1391 2325 1392
rect 2231 1386 2237 1387
rect 2319 1387 2320 1391
rect 2324 1390 2325 1391
rect 2327 1391 2333 1392
rect 2327 1390 2328 1391
rect 2324 1388 2328 1390
rect 2324 1387 2325 1388
rect 2319 1386 2325 1387
rect 2327 1387 2328 1388
rect 2332 1387 2333 1391
rect 2374 1391 2375 1395
rect 2379 1391 2380 1395
rect 2415 1395 2421 1396
rect 2415 1394 2416 1395
rect 2374 1390 2380 1391
rect 2407 1393 2416 1394
rect 2407 1389 2408 1393
rect 2412 1392 2416 1393
rect 2412 1389 2413 1392
rect 2415 1391 2416 1392
rect 2420 1391 2421 1395
rect 2415 1390 2421 1391
rect 2462 1395 2468 1396
rect 2462 1391 2463 1395
rect 2467 1391 2468 1395
rect 2526 1395 2532 1396
rect 2462 1390 2468 1391
rect 2495 1391 2501 1392
rect 2407 1388 2413 1389
rect 2327 1386 2333 1387
rect 2495 1387 2496 1391
rect 2500 1390 2501 1391
rect 2506 1391 2512 1392
rect 2506 1390 2507 1391
rect 2500 1388 2507 1390
rect 2500 1387 2501 1388
rect 2495 1386 2501 1387
rect 2506 1387 2507 1388
rect 2511 1387 2512 1391
rect 2526 1391 2527 1395
rect 2531 1391 2532 1395
rect 2582 1392 2583 1396
rect 2587 1392 2588 1396
rect 2526 1390 2532 1391
rect 2558 1391 2565 1392
rect 2582 1391 2588 1392
rect 2506 1386 2512 1387
rect 2558 1387 2559 1391
rect 2564 1387 2565 1391
rect 2558 1386 2565 1387
rect 1231 1382 1237 1383
rect 763 1380 787 1382
rect 763 1379 764 1380
rect 758 1378 764 1379
rect 334 1367 340 1368
rect 334 1363 335 1367
rect 339 1366 340 1367
rect 339 1364 435 1366
rect 339 1363 340 1364
rect 334 1362 340 1363
rect 433 1360 435 1364
rect 474 1363 480 1364
rect 175 1359 181 1360
rect 142 1357 148 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 142 1353 143 1357
rect 147 1353 148 1357
rect 175 1355 176 1359
rect 180 1358 181 1359
rect 198 1359 204 1360
rect 198 1358 199 1359
rect 180 1356 199 1358
rect 180 1355 181 1356
rect 175 1354 181 1355
rect 198 1355 199 1356
rect 203 1355 204 1359
rect 239 1359 245 1360
rect 198 1354 204 1355
rect 206 1357 212 1358
rect 142 1352 148 1353
rect 206 1353 207 1357
rect 211 1353 212 1357
rect 239 1355 240 1359
rect 244 1358 245 1359
rect 286 1359 292 1360
rect 286 1358 287 1359
rect 244 1356 287 1358
rect 244 1355 245 1356
rect 239 1354 245 1355
rect 286 1355 287 1356
rect 291 1355 292 1359
rect 327 1359 333 1360
rect 286 1354 292 1355
rect 294 1357 300 1358
rect 206 1352 212 1353
rect 294 1353 295 1357
rect 299 1353 300 1357
rect 327 1355 328 1359
rect 332 1358 333 1359
rect 390 1359 396 1360
rect 390 1358 391 1359
rect 332 1356 391 1358
rect 332 1355 333 1356
rect 327 1354 333 1355
rect 390 1355 391 1356
rect 395 1355 396 1359
rect 431 1359 437 1360
rect 390 1354 396 1355
rect 398 1357 404 1358
rect 294 1352 300 1353
rect 398 1353 399 1357
rect 403 1353 404 1357
rect 431 1355 432 1359
rect 436 1355 437 1359
rect 474 1359 475 1363
rect 479 1362 480 1363
rect 551 1363 557 1364
rect 479 1360 547 1362
rect 479 1359 480 1360
rect 474 1358 480 1359
rect 543 1359 549 1360
rect 431 1354 437 1355
rect 510 1357 516 1358
rect 398 1352 404 1353
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 543 1355 544 1359
rect 548 1355 549 1359
rect 551 1359 552 1363
rect 556 1362 557 1363
rect 556 1360 659 1362
rect 556 1359 557 1360
rect 551 1358 557 1359
rect 655 1359 661 1360
rect 543 1354 549 1355
rect 622 1357 628 1358
rect 510 1352 516 1353
rect 622 1353 623 1357
rect 627 1353 628 1357
rect 655 1355 656 1359
rect 660 1355 661 1359
rect 767 1359 773 1360
rect 655 1354 661 1355
rect 734 1357 740 1358
rect 622 1352 628 1353
rect 734 1353 735 1357
rect 739 1353 740 1357
rect 767 1355 768 1359
rect 772 1358 773 1359
rect 838 1359 844 1360
rect 838 1358 839 1359
rect 772 1356 839 1358
rect 772 1355 773 1356
rect 767 1354 773 1355
rect 838 1355 839 1356
rect 843 1355 844 1359
rect 870 1359 876 1360
rect 838 1354 844 1355
rect 846 1357 852 1358
rect 734 1352 740 1353
rect 846 1353 847 1357
rect 851 1353 852 1357
rect 870 1355 871 1359
rect 875 1358 876 1359
rect 879 1359 885 1360
rect 879 1358 880 1359
rect 875 1356 880 1358
rect 875 1355 876 1356
rect 870 1354 876 1355
rect 879 1355 880 1356
rect 884 1355 885 1359
rect 991 1359 997 1360
rect 879 1354 885 1355
rect 958 1357 964 1358
rect 846 1352 852 1353
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 991 1355 992 1359
rect 996 1358 997 1359
rect 1062 1359 1068 1360
rect 1062 1358 1063 1359
rect 996 1356 1063 1358
rect 996 1355 997 1356
rect 991 1354 997 1355
rect 1062 1355 1063 1356
rect 1067 1355 1068 1359
rect 1103 1359 1109 1360
rect 1062 1354 1068 1355
rect 1070 1357 1076 1358
rect 958 1352 964 1353
rect 1070 1353 1071 1357
rect 1075 1353 1076 1357
rect 1103 1355 1104 1359
rect 1108 1358 1109 1359
rect 1174 1359 1180 1360
rect 1174 1358 1175 1359
rect 1108 1356 1175 1358
rect 1108 1355 1109 1356
rect 1103 1354 1109 1355
rect 1174 1355 1175 1356
rect 1179 1355 1180 1359
rect 1215 1359 1221 1360
rect 1174 1354 1180 1355
rect 1182 1357 1188 1358
rect 1070 1352 1076 1353
rect 1182 1353 1183 1357
rect 1187 1353 1188 1357
rect 1215 1355 1216 1359
rect 1220 1358 1221 1359
rect 1262 1359 1268 1360
rect 1262 1358 1263 1359
rect 1220 1356 1263 1358
rect 1220 1355 1221 1356
rect 1215 1354 1221 1355
rect 1262 1355 1263 1356
rect 1267 1355 1268 1359
rect 1294 1359 1300 1360
rect 1262 1354 1268 1355
rect 1270 1357 1276 1358
rect 1182 1352 1188 1353
rect 1270 1353 1271 1357
rect 1275 1353 1276 1357
rect 1294 1355 1295 1359
rect 1299 1358 1300 1359
rect 1303 1359 1309 1360
rect 1303 1358 1304 1359
rect 1299 1356 1304 1358
rect 1299 1355 1300 1356
rect 1294 1354 1300 1355
rect 1303 1355 1304 1356
rect 1308 1355 1309 1359
rect 1847 1359 1853 1360
rect 1303 1354 1309 1355
rect 1326 1356 1332 1357
rect 1270 1352 1276 1353
rect 1326 1352 1327 1356
rect 1331 1352 1332 1356
rect 1431 1355 1437 1356
rect 1398 1353 1404 1354
rect 110 1351 116 1352
rect 1326 1351 1332 1352
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1431 1351 1432 1355
rect 1436 1354 1437 1355
rect 1446 1355 1452 1356
rect 1446 1354 1447 1355
rect 1436 1352 1447 1354
rect 1436 1351 1437 1352
rect 1431 1350 1437 1351
rect 1446 1351 1447 1352
rect 1451 1351 1452 1355
rect 1487 1355 1493 1356
rect 1446 1350 1452 1351
rect 1454 1353 1460 1354
rect 1398 1348 1404 1349
rect 1454 1349 1455 1353
rect 1459 1349 1460 1353
rect 1487 1351 1488 1355
rect 1492 1354 1493 1355
rect 1534 1355 1540 1356
rect 1534 1354 1535 1355
rect 1492 1352 1535 1354
rect 1492 1351 1493 1352
rect 1487 1350 1493 1351
rect 1534 1351 1535 1352
rect 1539 1351 1540 1355
rect 1575 1355 1581 1356
rect 1534 1350 1540 1351
rect 1542 1353 1548 1354
rect 1454 1348 1460 1349
rect 1542 1349 1543 1353
rect 1547 1349 1548 1353
rect 1575 1351 1576 1355
rect 1580 1354 1581 1355
rect 1622 1355 1628 1356
rect 1622 1354 1623 1355
rect 1580 1352 1623 1354
rect 1580 1351 1581 1352
rect 1575 1350 1581 1351
rect 1622 1351 1623 1352
rect 1627 1351 1628 1355
rect 1663 1355 1669 1356
rect 1622 1350 1628 1351
rect 1630 1353 1636 1354
rect 1542 1348 1548 1349
rect 1630 1349 1631 1353
rect 1635 1349 1636 1353
rect 1663 1351 1664 1355
rect 1668 1354 1669 1355
rect 1710 1355 1716 1356
rect 1710 1354 1711 1355
rect 1668 1352 1711 1354
rect 1668 1351 1669 1352
rect 1663 1350 1669 1351
rect 1710 1351 1711 1352
rect 1715 1351 1716 1355
rect 1750 1355 1757 1356
rect 1710 1350 1716 1351
rect 1718 1353 1724 1354
rect 1630 1348 1636 1349
rect 1718 1349 1719 1353
rect 1723 1349 1724 1353
rect 1750 1351 1751 1355
rect 1756 1351 1757 1355
rect 1838 1355 1845 1356
rect 1750 1350 1757 1351
rect 1806 1353 1812 1354
rect 1718 1348 1724 1349
rect 1806 1349 1807 1353
rect 1811 1349 1812 1353
rect 1838 1351 1839 1355
rect 1844 1351 1845 1355
rect 1847 1355 1848 1359
rect 1852 1358 1853 1359
rect 1852 1356 1923 1358
rect 1852 1355 1853 1356
rect 1847 1354 1853 1355
rect 1919 1355 1925 1356
rect 1838 1350 1845 1351
rect 1886 1353 1892 1354
rect 1806 1348 1812 1349
rect 1886 1349 1887 1353
rect 1891 1349 1892 1353
rect 1919 1351 1920 1355
rect 1924 1351 1925 1355
rect 1999 1355 2005 1356
rect 1919 1350 1925 1351
rect 1966 1353 1972 1354
rect 1886 1348 1892 1349
rect 1966 1349 1967 1353
rect 1971 1349 1972 1353
rect 1999 1351 2000 1355
rect 2004 1354 2005 1355
rect 2038 1355 2044 1356
rect 2038 1354 2039 1355
rect 2004 1352 2039 1354
rect 2004 1351 2005 1352
rect 1999 1350 2005 1351
rect 2038 1351 2039 1352
rect 2043 1351 2044 1355
rect 2079 1355 2085 1356
rect 2038 1350 2044 1351
rect 2046 1353 2052 1354
rect 1966 1348 1972 1349
rect 2046 1349 2047 1353
rect 2051 1349 2052 1353
rect 2079 1351 2080 1355
rect 2084 1354 2085 1355
rect 2118 1355 2124 1356
rect 2118 1354 2119 1355
rect 2084 1352 2119 1354
rect 2084 1351 2085 1352
rect 2079 1350 2085 1351
rect 2118 1351 2119 1352
rect 2123 1351 2124 1355
rect 2159 1355 2165 1356
rect 2118 1350 2124 1351
rect 2126 1353 2132 1354
rect 2046 1348 2052 1349
rect 2126 1349 2127 1353
rect 2131 1349 2132 1353
rect 2159 1351 2160 1355
rect 2164 1354 2165 1355
rect 2198 1355 2204 1356
rect 2198 1354 2199 1355
rect 2164 1352 2199 1354
rect 2164 1351 2165 1352
rect 2159 1350 2165 1351
rect 2198 1351 2199 1352
rect 2203 1351 2204 1355
rect 2238 1355 2245 1356
rect 2198 1350 2204 1351
rect 2206 1353 2212 1354
rect 2126 1348 2132 1349
rect 2206 1349 2207 1353
rect 2211 1349 2212 1353
rect 2238 1351 2239 1355
rect 2244 1351 2245 1355
rect 2238 1350 2245 1351
rect 2582 1352 2588 1353
rect 2206 1348 2212 1349
rect 2582 1348 2583 1352
rect 2587 1348 2588 1352
rect 1366 1347 1372 1348
rect 2582 1347 2588 1348
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 110 1334 116 1335
rect 1326 1339 1332 1340
rect 1326 1335 1327 1339
rect 1331 1335 1332 1339
rect 1326 1334 1332 1335
rect 1366 1335 1372 1336
rect 1366 1331 1367 1335
rect 1371 1331 1372 1335
rect 158 1330 164 1331
rect 158 1326 159 1330
rect 163 1326 164 1330
rect 158 1325 164 1326
rect 222 1330 228 1331
rect 222 1326 223 1330
rect 227 1326 228 1330
rect 222 1325 228 1326
rect 310 1330 316 1331
rect 310 1326 311 1330
rect 315 1326 316 1330
rect 310 1325 316 1326
rect 414 1330 420 1331
rect 414 1326 415 1330
rect 419 1326 420 1330
rect 414 1325 420 1326
rect 526 1330 532 1331
rect 526 1326 527 1330
rect 531 1326 532 1330
rect 526 1325 532 1326
rect 638 1330 644 1331
rect 638 1326 639 1330
rect 643 1326 644 1330
rect 638 1325 644 1326
rect 750 1330 756 1331
rect 750 1326 751 1330
rect 755 1326 756 1330
rect 750 1325 756 1326
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 862 1325 868 1326
rect 974 1330 980 1331
rect 974 1326 975 1330
rect 979 1326 980 1330
rect 974 1325 980 1326
rect 1086 1330 1092 1331
rect 1086 1326 1087 1330
rect 1091 1326 1092 1330
rect 1086 1325 1092 1326
rect 1198 1330 1204 1331
rect 1198 1326 1199 1330
rect 1203 1326 1204 1330
rect 1198 1325 1204 1326
rect 1286 1330 1292 1331
rect 1366 1330 1372 1331
rect 2582 1335 2588 1336
rect 2582 1331 2583 1335
rect 2587 1331 2588 1335
rect 2582 1330 2588 1331
rect 1286 1326 1287 1330
rect 1291 1326 1292 1330
rect 1286 1325 1292 1326
rect 1414 1326 1420 1327
rect 135 1323 141 1324
rect 135 1319 136 1323
rect 140 1322 141 1323
rect 174 1323 180 1324
rect 174 1322 175 1323
rect 140 1320 175 1322
rect 140 1319 141 1320
rect 135 1318 141 1319
rect 174 1319 175 1320
rect 179 1319 180 1323
rect 174 1318 180 1319
rect 198 1323 205 1324
rect 198 1319 199 1323
rect 204 1319 205 1323
rect 198 1318 205 1319
rect 286 1323 293 1324
rect 286 1319 287 1323
rect 292 1319 293 1323
rect 390 1323 397 1324
rect 286 1318 293 1319
rect 342 1319 348 1320
rect 342 1318 343 1319
rect 296 1316 343 1318
rect 296 1314 298 1316
rect 342 1315 343 1316
rect 347 1315 348 1319
rect 390 1319 391 1323
rect 396 1319 397 1323
rect 390 1318 397 1319
rect 503 1323 509 1324
rect 503 1319 504 1323
rect 508 1322 509 1323
rect 551 1323 557 1324
rect 551 1322 552 1323
rect 508 1320 552 1322
rect 508 1319 509 1320
rect 503 1318 509 1319
rect 551 1319 552 1320
rect 556 1319 557 1323
rect 551 1318 557 1319
rect 615 1323 621 1324
rect 615 1319 616 1323
rect 620 1322 621 1323
rect 670 1323 676 1324
rect 670 1322 671 1323
rect 620 1320 671 1322
rect 620 1319 621 1320
rect 615 1318 621 1319
rect 670 1319 671 1320
rect 675 1319 676 1323
rect 670 1318 676 1319
rect 727 1323 733 1324
rect 727 1319 728 1323
rect 732 1322 733 1323
rect 742 1323 748 1324
rect 742 1322 743 1323
rect 732 1320 743 1322
rect 732 1319 733 1320
rect 727 1318 733 1319
rect 742 1319 743 1320
rect 747 1319 748 1323
rect 742 1318 748 1319
rect 838 1323 845 1324
rect 838 1319 839 1323
rect 844 1319 845 1323
rect 838 1318 845 1319
rect 951 1323 957 1324
rect 951 1319 952 1323
rect 956 1322 957 1323
rect 998 1323 1004 1324
rect 998 1322 999 1323
rect 956 1320 999 1322
rect 956 1319 957 1320
rect 951 1318 957 1319
rect 998 1319 999 1320
rect 1003 1319 1004 1323
rect 998 1318 1004 1319
rect 1062 1323 1069 1324
rect 1062 1319 1063 1323
rect 1068 1319 1069 1323
rect 1062 1318 1069 1319
rect 1174 1323 1181 1324
rect 1174 1319 1175 1323
rect 1180 1319 1181 1323
rect 1174 1318 1181 1319
rect 1262 1323 1269 1324
rect 1262 1319 1263 1323
rect 1268 1319 1269 1323
rect 1414 1322 1415 1326
rect 1419 1322 1420 1326
rect 1414 1321 1420 1322
rect 1470 1326 1476 1327
rect 1470 1322 1471 1326
rect 1475 1322 1476 1326
rect 1470 1321 1476 1322
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1646 1326 1652 1327
rect 1646 1322 1647 1326
rect 1651 1322 1652 1326
rect 1646 1321 1652 1322
rect 1734 1326 1740 1327
rect 1734 1322 1735 1326
rect 1739 1322 1740 1326
rect 1734 1321 1740 1322
rect 1822 1326 1828 1327
rect 1822 1322 1823 1326
rect 1827 1322 1828 1326
rect 1822 1321 1828 1322
rect 1902 1326 1908 1327
rect 1902 1322 1903 1326
rect 1907 1322 1908 1326
rect 1902 1321 1908 1322
rect 1982 1326 1988 1327
rect 1982 1322 1983 1326
rect 1987 1322 1988 1326
rect 1982 1321 1988 1322
rect 2062 1326 2068 1327
rect 2062 1322 2063 1326
rect 2067 1322 2068 1326
rect 2062 1321 2068 1322
rect 2142 1326 2148 1327
rect 2142 1322 2143 1326
rect 2147 1322 2148 1326
rect 2142 1321 2148 1322
rect 2222 1326 2228 1327
rect 2222 1322 2223 1326
rect 2227 1322 2228 1326
rect 2222 1321 2228 1322
rect 1262 1318 1269 1319
rect 1306 1319 1312 1320
rect 342 1314 348 1315
rect 474 1315 480 1316
rect 474 1314 475 1315
rect 224 1312 298 1314
rect 424 1312 475 1314
rect 134 1311 141 1312
rect 134 1307 135 1311
rect 140 1307 141 1311
rect 207 1311 213 1312
rect 207 1307 208 1311
rect 212 1310 213 1311
rect 224 1310 226 1312
rect 212 1308 226 1310
rect 302 1311 309 1312
rect 212 1307 213 1308
rect 302 1307 303 1311
rect 308 1307 309 1311
rect 407 1311 413 1312
rect 407 1307 408 1311
rect 412 1310 413 1311
rect 424 1310 426 1312
rect 474 1311 475 1312
rect 479 1311 480 1315
rect 1306 1315 1307 1319
rect 1311 1318 1312 1319
rect 1391 1319 1397 1320
rect 1391 1318 1392 1319
rect 1311 1316 1392 1318
rect 1311 1315 1312 1316
rect 1306 1314 1312 1315
rect 1391 1315 1392 1316
rect 1396 1315 1397 1319
rect 1391 1314 1397 1315
rect 1446 1319 1453 1320
rect 1446 1315 1447 1319
rect 1452 1315 1453 1319
rect 1446 1314 1453 1315
rect 1534 1319 1541 1320
rect 1534 1315 1535 1319
rect 1540 1315 1541 1319
rect 1534 1314 1541 1315
rect 1622 1319 1629 1320
rect 1622 1315 1623 1319
rect 1628 1315 1629 1319
rect 1622 1314 1629 1315
rect 1710 1319 1717 1320
rect 1710 1315 1711 1319
rect 1716 1315 1717 1319
rect 1710 1314 1717 1315
rect 1799 1319 1805 1320
rect 1799 1315 1800 1319
rect 1804 1318 1805 1319
rect 1847 1319 1853 1320
rect 1847 1318 1848 1319
rect 1804 1316 1848 1318
rect 1804 1315 1805 1316
rect 1799 1314 1805 1315
rect 1847 1315 1848 1316
rect 1852 1315 1853 1319
rect 1847 1314 1853 1315
rect 1879 1319 1885 1320
rect 1879 1315 1880 1319
rect 1884 1318 1885 1319
rect 1934 1319 1940 1320
rect 1934 1318 1935 1319
rect 1884 1316 1935 1318
rect 1884 1315 1885 1316
rect 1879 1314 1885 1315
rect 1934 1315 1935 1316
rect 1939 1315 1940 1319
rect 1934 1314 1940 1315
rect 1959 1319 1965 1320
rect 1959 1315 1960 1319
rect 1964 1318 1965 1319
rect 1974 1319 1980 1320
rect 1974 1318 1975 1319
rect 1964 1316 1975 1318
rect 1964 1315 1965 1316
rect 1959 1314 1965 1315
rect 1974 1315 1975 1316
rect 1979 1315 1980 1319
rect 1974 1314 1980 1315
rect 2038 1319 2045 1320
rect 2038 1315 2039 1319
rect 2044 1315 2045 1319
rect 2038 1314 2045 1315
rect 2118 1319 2125 1320
rect 2118 1315 2119 1319
rect 2124 1315 2125 1319
rect 2118 1314 2125 1315
rect 2198 1319 2205 1320
rect 2198 1315 2199 1319
rect 2204 1315 2205 1319
rect 2198 1314 2205 1315
rect 474 1310 480 1311
rect 482 1311 488 1312
rect 412 1308 426 1310
rect 412 1307 413 1308
rect 482 1307 483 1311
rect 487 1310 488 1311
rect 511 1311 517 1312
rect 511 1310 512 1311
rect 487 1308 512 1310
rect 487 1307 488 1308
rect 134 1306 141 1307
rect 158 1306 164 1307
rect 207 1306 213 1307
rect 230 1306 236 1307
rect 302 1306 309 1307
rect 326 1306 332 1307
rect 407 1306 413 1307
rect 430 1306 436 1307
rect 482 1306 488 1307
rect 511 1307 512 1308
rect 516 1307 517 1311
rect 606 1311 613 1312
rect 606 1307 607 1311
rect 612 1307 613 1311
rect 650 1311 656 1312
rect 650 1307 651 1311
rect 655 1310 656 1311
rect 703 1311 709 1312
rect 703 1310 704 1311
rect 655 1308 704 1310
rect 655 1307 656 1308
rect 511 1306 517 1307
rect 534 1306 540 1307
rect 606 1306 613 1307
rect 630 1306 636 1307
rect 650 1306 656 1307
rect 703 1307 704 1308
rect 708 1307 709 1311
rect 778 1311 784 1312
rect 778 1307 779 1311
rect 783 1310 784 1311
rect 799 1311 805 1312
rect 799 1310 800 1311
rect 783 1308 800 1310
rect 783 1307 784 1308
rect 703 1306 709 1307
rect 726 1306 732 1307
rect 778 1306 784 1307
rect 799 1307 800 1308
rect 804 1307 805 1311
rect 887 1311 896 1312
rect 887 1307 888 1311
rect 895 1307 896 1311
rect 930 1311 936 1312
rect 930 1307 931 1311
rect 935 1310 936 1311
rect 967 1311 973 1312
rect 967 1310 968 1311
rect 935 1308 968 1310
rect 935 1307 936 1308
rect 799 1306 805 1307
rect 822 1306 828 1307
rect 887 1306 896 1307
rect 910 1306 916 1307
rect 930 1306 936 1307
rect 967 1307 968 1308
rect 972 1307 973 1311
rect 1010 1311 1016 1312
rect 1010 1307 1011 1311
rect 1015 1310 1016 1311
rect 1047 1311 1053 1312
rect 1047 1310 1048 1311
rect 1015 1308 1048 1310
rect 1015 1307 1016 1308
rect 967 1306 973 1307
rect 990 1306 996 1307
rect 1010 1306 1016 1307
rect 1047 1307 1048 1308
rect 1052 1307 1053 1311
rect 1110 1311 1116 1312
rect 1110 1307 1111 1311
rect 1115 1310 1116 1311
rect 1127 1311 1133 1312
rect 1127 1310 1128 1311
rect 1115 1308 1128 1310
rect 1115 1307 1116 1308
rect 1047 1306 1053 1307
rect 1070 1306 1076 1307
rect 1110 1306 1116 1307
rect 1127 1307 1128 1308
rect 1132 1307 1133 1311
rect 1170 1311 1176 1312
rect 1170 1307 1171 1311
rect 1175 1310 1176 1311
rect 1207 1311 1213 1312
rect 1207 1310 1208 1311
rect 1175 1308 1208 1310
rect 1175 1307 1176 1308
rect 1127 1306 1133 1307
rect 1150 1306 1156 1307
rect 1170 1306 1176 1307
rect 1207 1307 1208 1308
rect 1212 1307 1213 1311
rect 1250 1311 1256 1312
rect 1250 1307 1251 1311
rect 1255 1310 1256 1311
rect 1263 1311 1269 1312
rect 1263 1310 1264 1311
rect 1255 1308 1264 1310
rect 1255 1307 1256 1308
rect 1207 1306 1213 1307
rect 1230 1306 1236 1307
rect 1250 1306 1256 1307
rect 1263 1307 1264 1308
rect 1268 1307 1269 1311
rect 2054 1311 2060 1312
rect 2054 1310 2055 1311
rect 1999 1308 2055 1310
rect 1735 1307 1741 1308
rect 1263 1306 1269 1307
rect 1286 1306 1292 1307
rect 1735 1306 1736 1307
rect 158 1302 159 1306
rect 163 1302 164 1306
rect 158 1301 164 1302
rect 230 1302 231 1306
rect 235 1302 236 1306
rect 230 1301 236 1302
rect 326 1302 327 1306
rect 331 1302 332 1306
rect 326 1301 332 1302
rect 430 1302 431 1306
rect 435 1302 436 1306
rect 430 1301 436 1302
rect 534 1302 535 1306
rect 539 1302 540 1306
rect 534 1301 540 1302
rect 630 1302 631 1306
rect 635 1302 636 1306
rect 630 1301 636 1302
rect 726 1302 727 1306
rect 731 1302 732 1306
rect 726 1301 732 1302
rect 822 1302 823 1306
rect 827 1302 828 1306
rect 822 1301 828 1302
rect 910 1302 911 1306
rect 915 1302 916 1306
rect 910 1301 916 1302
rect 990 1302 991 1306
rect 995 1302 996 1306
rect 990 1301 996 1302
rect 1070 1302 1071 1306
rect 1075 1302 1076 1306
rect 1070 1301 1076 1302
rect 1150 1302 1151 1306
rect 1155 1302 1156 1306
rect 1150 1301 1156 1302
rect 1230 1302 1231 1306
rect 1235 1302 1236 1306
rect 1230 1301 1236 1302
rect 1286 1302 1287 1306
rect 1291 1302 1292 1306
rect 1664 1304 1736 1306
rect 1286 1301 1292 1302
rect 1647 1303 1653 1304
rect 1647 1299 1648 1303
rect 1652 1302 1653 1303
rect 1664 1302 1666 1304
rect 1735 1303 1736 1304
rect 1740 1303 1741 1307
rect 1790 1307 1796 1308
rect 1790 1306 1791 1307
rect 1760 1304 1791 1306
rect 1735 1302 1741 1303
rect 1743 1303 1749 1304
rect 1652 1300 1666 1302
rect 1652 1299 1653 1300
rect 1743 1299 1744 1303
rect 1748 1302 1749 1303
rect 1760 1302 1762 1304
rect 1790 1303 1791 1304
rect 1795 1303 1796 1307
rect 1999 1306 2001 1308
rect 2054 1307 2055 1308
rect 2059 1307 2060 1311
rect 2246 1311 2252 1312
rect 2246 1310 2247 1311
rect 2054 1306 2060 1307
rect 2129 1308 2247 1310
rect 1937 1304 2001 1306
rect 1790 1302 1796 1303
rect 1838 1303 1845 1304
rect 1748 1300 1762 1302
rect 1748 1299 1749 1300
rect 1838 1299 1839 1303
rect 1844 1299 1845 1303
rect 1935 1303 1941 1304
rect 1935 1299 1936 1303
rect 1940 1299 1941 1303
rect 2022 1303 2029 1304
rect 2022 1299 2023 1303
rect 2028 1299 2029 1303
rect 2111 1303 2117 1304
rect 2111 1299 2112 1303
rect 2116 1302 2117 1303
rect 2129 1302 2131 1308
rect 2246 1307 2247 1308
rect 2251 1307 2252 1311
rect 2246 1306 2252 1307
rect 2116 1300 2131 1302
rect 2186 1303 2192 1304
rect 2116 1299 2117 1300
rect 2186 1299 2187 1303
rect 2191 1302 2192 1303
rect 2207 1303 2213 1304
rect 2207 1302 2208 1303
rect 2191 1300 2208 1302
rect 2191 1299 2192 1300
rect 1647 1298 1653 1299
rect 1670 1298 1676 1299
rect 1743 1298 1749 1299
rect 1766 1298 1772 1299
rect 1838 1298 1845 1299
rect 1862 1298 1868 1299
rect 1935 1298 1941 1299
rect 1958 1298 1964 1299
rect 2022 1298 2029 1299
rect 2046 1298 2052 1299
rect 2111 1298 2117 1299
rect 2134 1298 2140 1299
rect 2186 1298 2192 1299
rect 2207 1299 2208 1300
rect 2212 1299 2213 1303
rect 2207 1298 2213 1299
rect 2230 1298 2236 1299
rect 110 1297 116 1298
rect 110 1293 111 1297
rect 115 1293 116 1297
rect 110 1292 116 1293
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1670 1294 1671 1298
rect 1675 1294 1676 1298
rect 1670 1293 1676 1294
rect 1766 1294 1767 1298
rect 1771 1294 1772 1298
rect 1766 1293 1772 1294
rect 1862 1294 1863 1298
rect 1867 1294 1868 1298
rect 1862 1293 1868 1294
rect 1958 1294 1959 1298
rect 1963 1294 1964 1298
rect 1958 1293 1964 1294
rect 2046 1294 2047 1298
rect 2051 1294 2052 1298
rect 2046 1293 2052 1294
rect 2134 1294 2135 1298
rect 2139 1294 2140 1298
rect 2134 1293 2140 1294
rect 2230 1294 2231 1298
rect 2235 1294 2236 1298
rect 2230 1293 2236 1294
rect 1326 1292 1332 1293
rect 1366 1289 1372 1290
rect 134 1287 140 1288
rect 134 1283 135 1287
rect 139 1286 140 1287
rect 606 1287 612 1288
rect 139 1284 242 1286
rect 139 1283 140 1284
rect 134 1282 140 1283
rect 110 1280 116 1281
rect 110 1276 111 1280
rect 115 1276 116 1280
rect 110 1275 116 1276
rect 142 1279 148 1280
rect 142 1275 143 1279
rect 147 1275 148 1279
rect 214 1279 220 1280
rect 142 1274 148 1275
rect 174 1275 181 1276
rect 174 1271 175 1275
rect 180 1271 181 1275
rect 214 1275 215 1279
rect 219 1275 220 1279
rect 214 1274 220 1275
rect 240 1274 242 1284
rect 606 1283 607 1287
rect 611 1286 612 1287
rect 611 1284 834 1286
rect 1366 1285 1367 1289
rect 1371 1285 1372 1289
rect 1366 1284 1372 1285
rect 2582 1289 2588 1290
rect 2582 1285 2583 1289
rect 2587 1285 2588 1289
rect 2582 1284 2588 1285
rect 611 1283 612 1284
rect 606 1282 612 1283
rect 310 1279 316 1280
rect 247 1275 253 1276
rect 247 1274 248 1275
rect 240 1272 248 1274
rect 174 1270 181 1271
rect 247 1271 248 1272
rect 252 1271 253 1275
rect 310 1275 311 1279
rect 315 1275 316 1279
rect 414 1279 420 1280
rect 310 1274 316 1275
rect 342 1275 349 1276
rect 247 1270 253 1271
rect 342 1271 343 1275
rect 348 1271 349 1275
rect 414 1275 415 1279
rect 419 1275 420 1279
rect 518 1279 524 1280
rect 414 1274 420 1275
rect 447 1275 453 1276
rect 342 1270 349 1271
rect 447 1271 448 1275
rect 452 1274 453 1275
rect 482 1275 488 1276
rect 482 1274 483 1275
rect 452 1272 483 1274
rect 452 1271 453 1272
rect 447 1270 453 1271
rect 482 1271 483 1272
rect 487 1271 488 1275
rect 518 1275 519 1279
rect 523 1275 524 1279
rect 614 1279 620 1280
rect 518 1274 524 1275
rect 542 1275 548 1276
rect 482 1270 488 1271
rect 542 1271 543 1275
rect 547 1274 548 1275
rect 551 1275 557 1276
rect 551 1274 552 1275
rect 547 1272 552 1274
rect 547 1271 548 1272
rect 542 1270 548 1271
rect 551 1271 552 1272
rect 556 1271 557 1275
rect 614 1275 615 1279
rect 619 1275 620 1279
rect 710 1279 716 1280
rect 614 1274 620 1275
rect 647 1275 656 1276
rect 551 1270 557 1271
rect 647 1271 648 1275
rect 655 1271 656 1275
rect 710 1275 711 1279
rect 715 1275 716 1279
rect 806 1279 812 1280
rect 710 1274 716 1275
rect 742 1275 749 1276
rect 647 1270 656 1271
rect 742 1271 743 1275
rect 748 1271 749 1275
rect 806 1275 807 1279
rect 811 1275 812 1279
rect 806 1274 812 1275
rect 832 1274 834 1284
rect 1326 1280 1332 1281
rect 894 1279 900 1280
rect 839 1275 845 1276
rect 839 1274 840 1275
rect 832 1272 840 1274
rect 742 1270 749 1271
rect 839 1271 840 1272
rect 844 1271 845 1275
rect 894 1275 895 1279
rect 899 1275 900 1279
rect 974 1279 980 1280
rect 894 1274 900 1275
rect 927 1275 936 1276
rect 839 1270 845 1271
rect 927 1271 928 1275
rect 935 1271 936 1275
rect 974 1275 975 1279
rect 979 1275 980 1279
rect 1054 1279 1060 1280
rect 974 1274 980 1275
rect 1007 1275 1016 1276
rect 927 1270 936 1271
rect 1007 1271 1008 1275
rect 1015 1271 1016 1275
rect 1054 1275 1055 1279
rect 1059 1275 1060 1279
rect 1110 1279 1116 1280
rect 1110 1278 1111 1279
rect 1054 1274 1060 1275
rect 1087 1277 1111 1278
rect 1087 1273 1088 1277
rect 1092 1276 1111 1277
rect 1092 1273 1093 1276
rect 1110 1275 1111 1276
rect 1115 1275 1116 1279
rect 1110 1274 1116 1275
rect 1134 1279 1140 1280
rect 1134 1275 1135 1279
rect 1139 1275 1140 1279
rect 1214 1279 1220 1280
rect 1134 1274 1140 1275
rect 1167 1275 1176 1276
rect 1087 1272 1093 1273
rect 1007 1270 1016 1271
rect 1167 1271 1168 1275
rect 1175 1271 1176 1275
rect 1214 1275 1215 1279
rect 1219 1275 1220 1279
rect 1270 1279 1276 1280
rect 1214 1274 1220 1275
rect 1247 1275 1256 1276
rect 1167 1270 1176 1271
rect 1247 1271 1248 1275
rect 1255 1271 1256 1275
rect 1270 1275 1271 1279
rect 1275 1275 1276 1279
rect 1326 1276 1327 1280
rect 1331 1276 1332 1280
rect 1270 1274 1276 1275
rect 1303 1275 1312 1276
rect 1326 1275 1332 1276
rect 2022 1279 2028 1280
rect 2022 1275 2023 1279
rect 2027 1278 2028 1279
rect 2027 1276 2146 1278
rect 2027 1275 2028 1276
rect 1247 1270 1256 1271
rect 1303 1271 1304 1275
rect 1311 1271 1312 1275
rect 2022 1274 2028 1275
rect 1303 1270 1312 1271
rect 1366 1272 1372 1273
rect 1366 1268 1367 1272
rect 1371 1268 1372 1272
rect 1366 1267 1372 1268
rect 1654 1271 1660 1272
rect 1654 1267 1655 1271
rect 1659 1267 1660 1271
rect 1750 1271 1756 1272
rect 1654 1266 1660 1267
rect 1687 1267 1693 1268
rect 1687 1266 1688 1267
rect 1664 1264 1688 1266
rect 1662 1263 1668 1264
rect 1662 1259 1663 1263
rect 1667 1259 1668 1263
rect 1687 1263 1688 1264
rect 1692 1263 1693 1267
rect 1750 1267 1751 1271
rect 1755 1267 1756 1271
rect 1846 1271 1852 1272
rect 1750 1266 1756 1267
rect 1783 1267 1789 1268
rect 1783 1266 1784 1267
rect 1760 1264 1784 1266
rect 1687 1262 1693 1263
rect 1735 1263 1741 1264
rect 1662 1258 1668 1259
rect 1735 1259 1736 1263
rect 1740 1262 1741 1263
rect 1760 1262 1762 1264
rect 1783 1263 1784 1264
rect 1788 1263 1789 1267
rect 1846 1267 1847 1271
rect 1851 1267 1852 1271
rect 1942 1271 1948 1272
rect 1846 1266 1852 1267
rect 1879 1267 1885 1268
rect 1783 1262 1789 1263
rect 1879 1263 1880 1267
rect 1884 1266 1885 1267
rect 1934 1267 1940 1268
rect 1934 1266 1935 1267
rect 1884 1264 1935 1266
rect 1884 1263 1885 1264
rect 1879 1262 1885 1263
rect 1934 1263 1935 1264
rect 1939 1263 1940 1267
rect 1942 1267 1943 1271
rect 1947 1267 1948 1271
rect 2030 1271 2036 1272
rect 1942 1266 1948 1267
rect 1974 1267 1981 1268
rect 1934 1262 1940 1263
rect 1974 1263 1975 1267
rect 1980 1263 1981 1267
rect 2030 1267 2031 1271
rect 2035 1267 2036 1271
rect 2118 1271 2124 1272
rect 2030 1266 2036 1267
rect 2054 1267 2060 1268
rect 1974 1262 1981 1263
rect 2054 1263 2055 1267
rect 2059 1266 2060 1267
rect 2063 1267 2069 1268
rect 2063 1266 2064 1267
rect 2059 1264 2064 1266
rect 2059 1263 2060 1264
rect 2054 1262 2060 1263
rect 2063 1263 2064 1264
rect 2068 1263 2069 1267
rect 2118 1267 2119 1271
rect 2123 1267 2124 1271
rect 2118 1266 2124 1267
rect 2144 1266 2146 1276
rect 2582 1272 2588 1273
rect 2214 1271 2220 1272
rect 2151 1267 2157 1268
rect 2151 1266 2152 1267
rect 2144 1264 2152 1266
rect 2063 1262 2069 1263
rect 2151 1263 2152 1264
rect 2156 1263 2157 1267
rect 2214 1267 2215 1271
rect 2219 1267 2220 1271
rect 2582 1268 2583 1272
rect 2587 1268 2588 1272
rect 2214 1266 2220 1267
rect 2246 1267 2253 1268
rect 2582 1267 2588 1268
rect 2151 1262 2157 1263
rect 2246 1263 2247 1267
rect 2252 1263 2253 1267
rect 2246 1262 2253 1263
rect 1740 1260 1762 1262
rect 1740 1259 1741 1260
rect 1735 1258 1741 1259
rect 1518 1247 1524 1248
rect 150 1243 156 1244
rect 150 1239 151 1243
rect 155 1242 156 1243
rect 822 1243 828 1244
rect 155 1240 321 1242
rect 155 1239 156 1240
rect 150 1238 156 1239
rect 319 1238 321 1240
rect 494 1239 500 1240
rect 319 1236 386 1238
rect 175 1235 181 1236
rect 142 1233 148 1234
rect 110 1232 116 1233
rect 110 1228 111 1232
rect 115 1228 116 1232
rect 142 1229 143 1233
rect 147 1229 148 1233
rect 175 1231 176 1235
rect 180 1234 181 1235
rect 190 1235 196 1236
rect 190 1234 191 1235
rect 180 1232 191 1234
rect 180 1231 181 1232
rect 175 1230 181 1231
rect 190 1231 191 1232
rect 195 1231 196 1235
rect 231 1235 237 1236
rect 190 1230 196 1231
rect 198 1233 204 1234
rect 142 1228 148 1229
rect 198 1229 199 1233
rect 203 1229 204 1233
rect 231 1231 232 1235
rect 236 1234 237 1235
rect 270 1235 276 1236
rect 270 1234 271 1235
rect 236 1232 271 1234
rect 236 1231 237 1232
rect 231 1230 237 1231
rect 270 1231 271 1232
rect 275 1231 276 1235
rect 302 1235 308 1236
rect 270 1230 276 1231
rect 278 1233 284 1234
rect 198 1228 204 1229
rect 278 1229 279 1233
rect 283 1229 284 1233
rect 302 1231 303 1235
rect 307 1234 308 1235
rect 311 1235 317 1236
rect 311 1234 312 1235
rect 307 1232 312 1234
rect 307 1231 308 1232
rect 302 1230 308 1231
rect 311 1231 312 1232
rect 316 1231 317 1235
rect 384 1234 386 1236
rect 391 1235 397 1236
rect 391 1234 392 1235
rect 311 1230 317 1231
rect 358 1233 364 1234
rect 278 1228 284 1229
rect 358 1229 359 1233
rect 363 1229 364 1233
rect 384 1232 392 1234
rect 391 1231 392 1232
rect 396 1231 397 1235
rect 471 1235 477 1236
rect 391 1230 397 1231
rect 438 1233 444 1234
rect 358 1228 364 1229
rect 438 1229 439 1233
rect 443 1229 444 1233
rect 471 1231 472 1235
rect 476 1234 477 1235
rect 486 1235 492 1236
rect 486 1234 487 1235
rect 476 1232 487 1234
rect 476 1231 477 1232
rect 471 1230 477 1231
rect 486 1231 487 1232
rect 491 1231 492 1235
rect 494 1235 495 1239
rect 499 1238 500 1239
rect 822 1239 823 1243
rect 827 1242 828 1243
rect 1518 1243 1519 1247
rect 1523 1246 1524 1247
rect 1694 1247 1700 1248
rect 1523 1244 1650 1246
rect 1523 1243 1524 1244
rect 1518 1242 1524 1243
rect 827 1240 931 1242
rect 827 1239 828 1240
rect 822 1238 828 1239
rect 499 1236 546 1238
rect 929 1236 931 1240
rect 1527 1239 1533 1240
rect 1494 1237 1500 1238
rect 1366 1236 1372 1237
rect 499 1235 500 1236
rect 494 1234 500 1235
rect 544 1234 546 1236
rect 551 1235 557 1236
rect 551 1234 552 1235
rect 486 1230 492 1231
rect 518 1233 524 1234
rect 438 1228 444 1229
rect 518 1229 519 1233
rect 523 1229 524 1233
rect 544 1232 552 1234
rect 551 1231 552 1232
rect 556 1231 557 1235
rect 631 1235 637 1236
rect 551 1230 557 1231
rect 598 1233 604 1234
rect 518 1228 524 1229
rect 598 1229 599 1233
rect 603 1229 604 1233
rect 631 1231 632 1235
rect 636 1234 637 1235
rect 662 1235 668 1236
rect 662 1234 663 1235
rect 636 1232 663 1234
rect 636 1231 637 1232
rect 631 1230 637 1231
rect 662 1231 663 1232
rect 667 1231 668 1235
rect 703 1235 709 1236
rect 662 1230 668 1231
rect 670 1233 676 1234
rect 598 1228 604 1229
rect 670 1229 671 1233
rect 675 1229 676 1233
rect 703 1231 704 1235
rect 708 1234 709 1235
rect 734 1235 740 1236
rect 734 1234 735 1235
rect 708 1232 735 1234
rect 708 1231 709 1232
rect 703 1230 709 1231
rect 734 1231 735 1232
rect 739 1231 740 1235
rect 775 1235 784 1236
rect 734 1230 740 1231
rect 742 1233 748 1234
rect 670 1228 676 1229
rect 742 1229 743 1233
rect 747 1229 748 1233
rect 775 1231 776 1235
rect 783 1231 784 1235
rect 846 1235 853 1236
rect 775 1230 784 1231
rect 814 1233 820 1234
rect 742 1228 748 1229
rect 814 1229 815 1233
rect 819 1229 820 1233
rect 846 1231 847 1235
rect 852 1231 853 1235
rect 927 1235 933 1236
rect 846 1230 853 1231
rect 894 1233 900 1234
rect 814 1228 820 1229
rect 894 1229 895 1233
rect 899 1229 900 1233
rect 927 1231 928 1235
rect 932 1231 933 1235
rect 927 1230 933 1231
rect 1326 1232 1332 1233
rect 894 1228 900 1229
rect 1326 1228 1327 1232
rect 1331 1228 1332 1232
rect 1366 1232 1367 1236
rect 1371 1232 1372 1236
rect 1494 1233 1495 1237
rect 1499 1233 1500 1237
rect 1527 1235 1528 1239
rect 1532 1238 1533 1239
rect 1550 1239 1556 1240
rect 1550 1238 1551 1239
rect 1532 1236 1551 1238
rect 1532 1235 1533 1236
rect 1527 1234 1533 1235
rect 1550 1235 1551 1236
rect 1555 1235 1556 1239
rect 1586 1239 1597 1240
rect 1550 1234 1556 1235
rect 1558 1237 1564 1238
rect 1494 1232 1500 1233
rect 1558 1233 1559 1237
rect 1563 1233 1564 1237
rect 1586 1235 1587 1239
rect 1591 1235 1592 1239
rect 1596 1235 1597 1239
rect 1648 1238 1650 1244
rect 1694 1243 1695 1247
rect 1699 1246 1700 1247
rect 2086 1247 2092 1248
rect 1699 1244 1850 1246
rect 1699 1243 1700 1244
rect 1694 1242 1700 1243
rect 1655 1239 1661 1240
rect 1655 1238 1656 1239
rect 1586 1234 1597 1235
rect 1622 1237 1628 1238
rect 1558 1232 1564 1233
rect 1622 1233 1623 1237
rect 1627 1233 1628 1237
rect 1648 1236 1656 1238
rect 1655 1235 1656 1236
rect 1660 1235 1661 1239
rect 1719 1239 1725 1240
rect 1655 1234 1661 1235
rect 1686 1237 1692 1238
rect 1622 1232 1628 1233
rect 1686 1233 1687 1237
rect 1691 1233 1692 1237
rect 1719 1235 1720 1239
rect 1724 1238 1725 1239
rect 1750 1239 1756 1240
rect 1750 1238 1751 1239
rect 1724 1236 1751 1238
rect 1724 1235 1725 1236
rect 1719 1234 1725 1235
rect 1750 1235 1751 1236
rect 1755 1235 1756 1239
rect 1790 1239 1797 1240
rect 1750 1234 1756 1235
rect 1758 1237 1764 1238
rect 1686 1232 1692 1233
rect 1758 1233 1759 1237
rect 1763 1233 1764 1237
rect 1790 1235 1791 1239
rect 1796 1235 1797 1239
rect 1848 1238 1850 1244
rect 1863 1243 1869 1244
rect 1855 1239 1861 1240
rect 1855 1238 1856 1239
rect 1790 1234 1797 1235
rect 1822 1237 1828 1238
rect 1758 1232 1764 1233
rect 1822 1233 1823 1237
rect 1827 1233 1828 1237
rect 1848 1236 1856 1238
rect 1855 1235 1856 1236
rect 1860 1235 1861 1239
rect 1863 1239 1864 1243
rect 1868 1242 1869 1243
rect 2086 1243 2087 1247
rect 2091 1246 2092 1247
rect 2091 1244 2322 1246
rect 2091 1243 2092 1244
rect 2086 1242 2092 1243
rect 1868 1240 1923 1242
rect 1868 1239 1869 1240
rect 1863 1238 1869 1239
rect 1919 1239 1925 1240
rect 1855 1234 1861 1235
rect 1886 1237 1892 1238
rect 1822 1232 1828 1233
rect 1886 1233 1887 1237
rect 1891 1233 1892 1237
rect 1919 1235 1920 1239
rect 1924 1235 1925 1239
rect 1983 1239 1989 1240
rect 1919 1234 1925 1235
rect 1950 1237 1956 1238
rect 1886 1232 1892 1233
rect 1950 1233 1951 1237
rect 1955 1233 1956 1237
rect 1983 1235 1984 1239
rect 1988 1238 1989 1239
rect 2006 1239 2012 1240
rect 2006 1238 2007 1239
rect 1988 1236 2007 1238
rect 1988 1235 1989 1236
rect 1983 1234 1989 1235
rect 2006 1235 2007 1236
rect 2011 1235 2012 1239
rect 2038 1239 2044 1240
rect 2006 1234 2012 1235
rect 2014 1237 2020 1238
rect 1950 1232 1956 1233
rect 2014 1233 2015 1237
rect 2019 1233 2020 1237
rect 2038 1235 2039 1239
rect 2043 1238 2044 1239
rect 2047 1239 2053 1240
rect 2047 1238 2048 1239
rect 2043 1236 2048 1238
rect 2043 1235 2044 1236
rect 2038 1234 2044 1235
rect 2047 1235 2048 1236
rect 2052 1235 2053 1239
rect 2111 1239 2117 1240
rect 2047 1234 2053 1235
rect 2078 1237 2084 1238
rect 2014 1232 2020 1233
rect 2078 1233 2079 1237
rect 2083 1233 2084 1237
rect 2111 1235 2112 1239
rect 2116 1238 2117 1239
rect 2138 1239 2144 1240
rect 2138 1238 2139 1239
rect 2116 1236 2139 1238
rect 2116 1235 2117 1236
rect 2111 1234 2117 1235
rect 2138 1235 2139 1236
rect 2143 1235 2144 1239
rect 2183 1239 2192 1240
rect 2138 1234 2144 1235
rect 2150 1237 2156 1238
rect 2078 1232 2084 1233
rect 2150 1233 2151 1237
rect 2155 1233 2156 1237
rect 2183 1235 2184 1239
rect 2191 1235 2192 1239
rect 2255 1239 2261 1240
rect 2183 1234 2192 1235
rect 2222 1237 2228 1238
rect 2150 1232 2156 1233
rect 2222 1233 2223 1237
rect 2227 1233 2228 1237
rect 2255 1235 2256 1239
rect 2260 1238 2261 1239
rect 2286 1239 2292 1240
rect 2286 1238 2287 1239
rect 2260 1236 2287 1238
rect 2260 1235 2261 1236
rect 2255 1234 2261 1235
rect 2286 1235 2287 1236
rect 2291 1235 2292 1239
rect 2320 1238 2322 1244
rect 2327 1239 2333 1240
rect 2327 1238 2328 1239
rect 2286 1234 2292 1235
rect 2294 1237 2300 1238
rect 2222 1232 2228 1233
rect 2294 1233 2295 1237
rect 2299 1233 2300 1237
rect 2320 1236 2328 1238
rect 2327 1235 2328 1236
rect 2332 1235 2333 1239
rect 2327 1234 2333 1235
rect 2582 1236 2588 1237
rect 2294 1232 2300 1233
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 1366 1231 1372 1232
rect 2582 1231 2588 1232
rect 110 1227 116 1228
rect 1326 1227 1332 1228
rect 1366 1219 1372 1220
rect 110 1215 116 1216
rect 110 1211 111 1215
rect 115 1211 116 1215
rect 110 1210 116 1211
rect 1326 1215 1332 1216
rect 1326 1211 1327 1215
rect 1331 1211 1332 1215
rect 1366 1215 1367 1219
rect 1371 1215 1372 1219
rect 1366 1214 1372 1215
rect 2582 1219 2588 1220
rect 2582 1215 2583 1219
rect 2587 1215 2588 1219
rect 2582 1214 2588 1215
rect 1326 1210 1332 1211
rect 1510 1210 1516 1211
rect 158 1206 164 1207
rect 158 1202 159 1206
rect 163 1202 164 1206
rect 158 1201 164 1202
rect 214 1206 220 1207
rect 214 1202 215 1206
rect 219 1202 220 1206
rect 214 1201 220 1202
rect 294 1206 300 1207
rect 294 1202 295 1206
rect 299 1202 300 1206
rect 294 1201 300 1202
rect 374 1206 380 1207
rect 374 1202 375 1206
rect 379 1202 380 1206
rect 374 1201 380 1202
rect 454 1206 460 1207
rect 454 1202 455 1206
rect 459 1202 460 1206
rect 454 1201 460 1202
rect 534 1206 540 1207
rect 534 1202 535 1206
rect 539 1202 540 1206
rect 534 1201 540 1202
rect 614 1206 620 1207
rect 614 1202 615 1206
rect 619 1202 620 1206
rect 614 1201 620 1202
rect 686 1206 692 1207
rect 686 1202 687 1206
rect 691 1202 692 1206
rect 686 1201 692 1202
rect 758 1206 764 1207
rect 758 1202 759 1206
rect 763 1202 764 1206
rect 758 1201 764 1202
rect 830 1206 836 1207
rect 830 1202 831 1206
rect 835 1202 836 1206
rect 830 1201 836 1202
rect 910 1206 916 1207
rect 910 1202 911 1206
rect 915 1202 916 1206
rect 1510 1206 1511 1210
rect 1515 1206 1516 1210
rect 1510 1205 1516 1206
rect 1574 1210 1580 1211
rect 1574 1206 1575 1210
rect 1579 1206 1580 1210
rect 1574 1205 1580 1206
rect 1638 1210 1644 1211
rect 1638 1206 1639 1210
rect 1643 1206 1644 1210
rect 1638 1205 1644 1206
rect 1702 1210 1708 1211
rect 1702 1206 1703 1210
rect 1707 1206 1708 1210
rect 1702 1205 1708 1206
rect 1774 1210 1780 1211
rect 1774 1206 1775 1210
rect 1779 1206 1780 1210
rect 1774 1205 1780 1206
rect 1838 1210 1844 1211
rect 1838 1206 1839 1210
rect 1843 1206 1844 1210
rect 1838 1205 1844 1206
rect 1902 1210 1908 1211
rect 1902 1206 1903 1210
rect 1907 1206 1908 1210
rect 1902 1205 1908 1206
rect 1966 1210 1972 1211
rect 1966 1206 1967 1210
rect 1971 1206 1972 1210
rect 1966 1205 1972 1206
rect 2030 1210 2036 1211
rect 2030 1206 2031 1210
rect 2035 1206 2036 1210
rect 2030 1205 2036 1206
rect 2094 1210 2100 1211
rect 2094 1206 2095 1210
rect 2099 1206 2100 1210
rect 2094 1205 2100 1206
rect 2166 1210 2172 1211
rect 2166 1206 2167 1210
rect 2171 1206 2172 1210
rect 2166 1205 2172 1206
rect 2238 1210 2244 1211
rect 2238 1206 2239 1210
rect 2243 1206 2244 1210
rect 2238 1205 2244 1206
rect 2310 1210 2316 1211
rect 2310 1206 2311 1210
rect 2315 1206 2316 1210
rect 2310 1205 2316 1206
rect 910 1201 916 1202
rect 1487 1203 1493 1204
rect 135 1199 141 1200
rect 135 1195 136 1199
rect 140 1198 141 1199
rect 150 1199 156 1200
rect 150 1198 151 1199
rect 140 1196 151 1198
rect 140 1195 141 1196
rect 135 1194 141 1195
rect 150 1195 151 1196
rect 155 1195 156 1199
rect 150 1194 156 1195
rect 190 1199 197 1200
rect 190 1195 191 1199
rect 196 1195 197 1199
rect 190 1194 197 1195
rect 270 1199 277 1200
rect 270 1195 271 1199
rect 276 1195 277 1199
rect 270 1194 277 1195
rect 346 1199 357 1200
rect 346 1195 347 1199
rect 351 1195 352 1199
rect 356 1195 357 1199
rect 346 1194 357 1195
rect 431 1199 437 1200
rect 431 1195 432 1199
rect 436 1198 437 1199
rect 494 1199 500 1200
rect 494 1198 495 1199
rect 436 1196 495 1198
rect 436 1195 437 1196
rect 431 1194 437 1195
rect 494 1195 495 1196
rect 499 1195 500 1199
rect 494 1194 500 1195
rect 511 1199 517 1200
rect 511 1195 512 1199
rect 516 1198 517 1199
rect 542 1199 548 1200
rect 542 1198 543 1199
rect 516 1196 543 1198
rect 516 1195 517 1196
rect 511 1194 517 1195
rect 542 1195 543 1196
rect 547 1195 548 1199
rect 542 1194 548 1195
rect 591 1199 597 1200
rect 591 1195 592 1199
rect 596 1198 597 1199
rect 662 1199 669 1200
rect 596 1196 659 1198
rect 596 1195 597 1196
rect 591 1194 597 1195
rect 657 1190 659 1196
rect 662 1195 663 1199
rect 668 1195 669 1199
rect 662 1194 669 1195
rect 734 1199 741 1200
rect 734 1195 735 1199
rect 740 1195 741 1199
rect 734 1194 741 1195
rect 807 1199 813 1200
rect 807 1195 808 1199
rect 812 1198 813 1199
rect 822 1199 828 1200
rect 822 1198 823 1199
rect 812 1196 823 1198
rect 812 1195 813 1196
rect 807 1194 813 1195
rect 822 1195 823 1196
rect 827 1195 828 1199
rect 822 1194 828 1195
rect 858 1199 864 1200
rect 858 1195 859 1199
rect 863 1198 864 1199
rect 887 1199 893 1200
rect 887 1198 888 1199
rect 863 1196 888 1198
rect 863 1195 864 1196
rect 858 1194 864 1195
rect 887 1195 888 1196
rect 892 1195 893 1199
rect 1487 1199 1488 1203
rect 1492 1202 1493 1203
rect 1518 1203 1524 1204
rect 1518 1202 1519 1203
rect 1492 1200 1519 1202
rect 1492 1199 1493 1200
rect 1487 1198 1493 1199
rect 1518 1199 1519 1200
rect 1523 1199 1524 1203
rect 1518 1198 1524 1199
rect 1550 1203 1557 1204
rect 1550 1199 1551 1203
rect 1556 1199 1557 1203
rect 1550 1198 1557 1199
rect 1615 1203 1621 1204
rect 1615 1199 1616 1203
rect 1620 1202 1621 1203
rect 1662 1203 1668 1204
rect 1662 1202 1663 1203
rect 1620 1200 1663 1202
rect 1620 1199 1621 1200
rect 1615 1198 1621 1199
rect 1662 1199 1663 1200
rect 1667 1199 1668 1203
rect 1662 1198 1668 1199
rect 1679 1203 1685 1204
rect 1679 1199 1680 1203
rect 1684 1202 1685 1203
rect 1694 1203 1700 1204
rect 1694 1202 1695 1203
rect 1684 1200 1695 1202
rect 1684 1199 1685 1200
rect 1679 1198 1685 1199
rect 1694 1199 1695 1200
rect 1699 1199 1700 1203
rect 1694 1198 1700 1199
rect 1750 1203 1757 1204
rect 1750 1199 1751 1203
rect 1756 1199 1757 1203
rect 1750 1198 1757 1199
rect 1815 1203 1821 1204
rect 1815 1199 1816 1203
rect 1820 1202 1821 1203
rect 1863 1203 1869 1204
rect 1863 1202 1864 1203
rect 1820 1200 1864 1202
rect 1820 1199 1821 1200
rect 1815 1198 1821 1199
rect 1863 1199 1864 1200
rect 1868 1199 1869 1203
rect 1863 1198 1869 1199
rect 1879 1203 1885 1204
rect 1879 1199 1880 1203
rect 1884 1202 1885 1203
rect 1926 1203 1932 1204
rect 1926 1202 1927 1203
rect 1884 1200 1927 1202
rect 1884 1199 1885 1200
rect 1879 1198 1885 1199
rect 1926 1199 1927 1200
rect 1931 1199 1932 1203
rect 1926 1198 1932 1199
rect 1934 1203 1940 1204
rect 1934 1199 1935 1203
rect 1939 1202 1940 1203
rect 1943 1203 1949 1204
rect 1943 1202 1944 1203
rect 1939 1200 1944 1202
rect 1939 1199 1940 1200
rect 1934 1198 1940 1199
rect 1943 1199 1944 1200
rect 1948 1199 1949 1203
rect 1943 1198 1949 1199
rect 2006 1203 2013 1204
rect 2006 1199 2007 1203
rect 2012 1199 2013 1203
rect 2006 1198 2013 1199
rect 2071 1203 2077 1204
rect 2071 1199 2072 1203
rect 2076 1202 2077 1203
rect 2086 1203 2092 1204
rect 2086 1202 2087 1203
rect 2076 1200 2087 1202
rect 2076 1199 2077 1200
rect 2071 1198 2077 1199
rect 2086 1199 2087 1200
rect 2091 1199 2092 1203
rect 2086 1198 2092 1199
rect 2138 1203 2149 1204
rect 2138 1199 2139 1203
rect 2143 1199 2144 1203
rect 2148 1199 2149 1203
rect 2138 1198 2149 1199
rect 2215 1203 2224 1204
rect 2215 1199 2216 1203
rect 2223 1199 2224 1203
rect 2215 1198 2224 1199
rect 2286 1203 2293 1204
rect 2286 1199 2287 1203
rect 2292 1199 2293 1203
rect 2286 1198 2293 1199
rect 887 1194 893 1195
rect 846 1191 852 1192
rect 846 1190 847 1191
rect 657 1188 847 1190
rect 846 1187 847 1188
rect 851 1187 852 1191
rect 846 1186 852 1187
rect 1586 1187 1592 1188
rect 1586 1186 1587 1187
rect 1575 1185 1587 1186
rect 134 1183 141 1184
rect 134 1179 135 1183
rect 140 1179 141 1183
rect 183 1183 189 1184
rect 183 1179 184 1183
rect 188 1182 189 1183
rect 215 1183 221 1184
rect 215 1182 216 1183
rect 188 1180 216 1182
rect 188 1179 189 1180
rect 134 1178 141 1179
rect 158 1178 164 1179
rect 183 1178 189 1179
rect 215 1179 216 1180
rect 220 1179 221 1183
rect 258 1183 264 1184
rect 258 1179 259 1183
rect 263 1182 264 1183
rect 303 1183 309 1184
rect 303 1182 304 1183
rect 263 1180 304 1182
rect 263 1179 264 1180
rect 215 1178 221 1179
rect 238 1178 244 1179
rect 258 1178 264 1179
rect 303 1179 304 1180
rect 308 1179 309 1183
rect 354 1183 360 1184
rect 354 1179 355 1183
rect 359 1182 360 1183
rect 399 1183 405 1184
rect 399 1182 400 1183
rect 359 1180 400 1182
rect 359 1179 360 1180
rect 303 1178 309 1179
rect 326 1178 332 1179
rect 354 1178 360 1179
rect 399 1179 400 1180
rect 404 1179 405 1183
rect 486 1183 493 1184
rect 486 1179 487 1183
rect 492 1179 493 1183
rect 535 1183 541 1184
rect 535 1179 536 1183
rect 540 1182 541 1183
rect 575 1183 581 1184
rect 575 1182 576 1183
rect 540 1180 576 1182
rect 540 1179 541 1180
rect 399 1178 405 1179
rect 422 1178 428 1179
rect 486 1178 493 1179
rect 510 1178 516 1179
rect 535 1178 541 1179
rect 575 1179 576 1180
rect 580 1179 581 1183
rect 663 1183 669 1184
rect 663 1179 664 1183
rect 668 1182 669 1183
rect 678 1183 684 1184
rect 678 1182 679 1183
rect 668 1180 679 1182
rect 668 1179 669 1180
rect 575 1178 581 1179
rect 598 1178 604 1179
rect 663 1178 669 1179
rect 678 1179 679 1180
rect 683 1179 684 1183
rect 706 1183 712 1184
rect 706 1179 707 1183
rect 711 1182 712 1183
rect 743 1183 749 1184
rect 743 1182 744 1183
rect 711 1180 744 1182
rect 711 1179 712 1180
rect 678 1178 684 1179
rect 686 1178 692 1179
rect 706 1178 712 1179
rect 743 1179 744 1180
rect 748 1179 749 1183
rect 786 1183 792 1184
rect 786 1179 787 1183
rect 791 1182 792 1183
rect 815 1183 821 1184
rect 815 1182 816 1183
rect 791 1180 816 1182
rect 791 1179 792 1180
rect 743 1178 749 1179
rect 766 1178 772 1179
rect 786 1178 792 1179
rect 815 1179 816 1180
rect 820 1179 821 1183
rect 886 1183 893 1184
rect 886 1179 887 1183
rect 892 1179 893 1183
rect 951 1183 957 1184
rect 951 1179 952 1183
rect 956 1182 957 1183
rect 959 1183 965 1184
rect 959 1182 960 1183
rect 956 1180 960 1182
rect 956 1179 957 1180
rect 815 1178 821 1179
rect 838 1178 844 1179
rect 886 1178 893 1179
rect 910 1178 916 1179
rect 951 1178 957 1179
rect 959 1179 960 1180
rect 964 1179 965 1183
rect 1002 1183 1008 1184
rect 1002 1179 1003 1183
rect 1007 1182 1008 1183
rect 1039 1183 1045 1184
rect 1039 1182 1040 1183
rect 1007 1180 1040 1182
rect 1007 1179 1008 1180
rect 959 1178 965 1179
rect 982 1178 988 1179
rect 1002 1178 1008 1179
rect 1039 1179 1040 1180
rect 1044 1179 1045 1183
rect 1390 1183 1397 1184
rect 1390 1179 1391 1183
rect 1396 1179 1397 1183
rect 1479 1183 1485 1184
rect 1479 1179 1480 1183
rect 1484 1182 1485 1183
rect 1494 1183 1500 1184
rect 1494 1182 1495 1183
rect 1484 1180 1495 1182
rect 1484 1179 1485 1180
rect 1039 1178 1045 1179
rect 1062 1178 1068 1179
rect 1390 1178 1397 1179
rect 1414 1178 1420 1179
rect 1479 1178 1485 1179
rect 1494 1179 1495 1180
rect 1499 1179 1500 1183
rect 1575 1181 1576 1185
rect 1580 1184 1587 1185
rect 1580 1181 1581 1184
rect 1586 1183 1587 1184
rect 1591 1183 1592 1187
rect 2038 1187 2044 1188
rect 2038 1186 2039 1187
rect 1999 1184 2039 1186
rect 1586 1182 1592 1183
rect 1618 1183 1624 1184
rect 1575 1180 1581 1181
rect 1618 1179 1619 1183
rect 1623 1182 1624 1183
rect 1679 1183 1685 1184
rect 1679 1182 1680 1183
rect 1623 1180 1680 1182
rect 1623 1179 1624 1180
rect 1494 1178 1500 1179
rect 1502 1178 1508 1179
rect 158 1174 159 1178
rect 163 1174 164 1178
rect 158 1173 164 1174
rect 238 1174 239 1178
rect 243 1174 244 1178
rect 238 1173 244 1174
rect 326 1174 327 1178
rect 331 1174 332 1178
rect 326 1173 332 1174
rect 422 1174 423 1178
rect 427 1174 428 1178
rect 422 1173 428 1174
rect 510 1174 511 1178
rect 515 1174 516 1178
rect 510 1173 516 1174
rect 598 1174 599 1178
rect 603 1174 604 1178
rect 598 1173 604 1174
rect 686 1174 687 1178
rect 691 1174 692 1178
rect 686 1173 692 1174
rect 766 1174 767 1178
rect 771 1174 772 1178
rect 766 1173 772 1174
rect 838 1174 839 1178
rect 843 1174 844 1178
rect 838 1173 844 1174
rect 910 1174 911 1178
rect 915 1174 916 1178
rect 910 1173 916 1174
rect 982 1174 983 1178
rect 987 1174 988 1178
rect 982 1173 988 1174
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1414 1174 1415 1178
rect 1419 1174 1420 1178
rect 1414 1173 1420 1174
rect 1502 1174 1503 1178
rect 1507 1174 1508 1178
rect 1502 1173 1508 1174
rect 1598 1178 1604 1179
rect 1618 1178 1624 1179
rect 1679 1179 1680 1180
rect 1684 1179 1685 1183
rect 1722 1183 1728 1184
rect 1722 1179 1723 1183
rect 1727 1182 1728 1183
rect 1783 1183 1789 1184
rect 1783 1182 1784 1183
rect 1727 1180 1784 1182
rect 1727 1179 1728 1180
rect 1679 1178 1685 1179
rect 1702 1178 1708 1179
rect 1722 1178 1728 1179
rect 1783 1179 1784 1180
rect 1788 1179 1789 1183
rect 1826 1183 1832 1184
rect 1826 1179 1827 1183
rect 1831 1182 1832 1183
rect 1887 1183 1893 1184
rect 1887 1182 1888 1183
rect 1831 1180 1888 1182
rect 1831 1179 1832 1180
rect 1783 1178 1789 1179
rect 1806 1178 1812 1179
rect 1826 1178 1832 1179
rect 1887 1179 1888 1180
rect 1892 1179 1893 1183
rect 1991 1183 1997 1184
rect 1991 1179 1992 1183
rect 1996 1182 1997 1183
rect 1999 1182 2001 1184
rect 2038 1183 2039 1184
rect 2043 1183 2044 1187
rect 2038 1182 2044 1183
rect 2086 1183 2093 1184
rect 1996 1180 2001 1182
rect 1996 1179 1997 1180
rect 2086 1179 2087 1183
rect 2092 1179 2093 1183
rect 2130 1183 2136 1184
rect 2130 1179 2131 1183
rect 2135 1182 2136 1183
rect 2183 1183 2189 1184
rect 2183 1182 2184 1183
rect 2135 1180 2184 1182
rect 2135 1179 2136 1180
rect 1887 1178 1893 1179
rect 1910 1178 1916 1179
rect 1991 1178 1997 1179
rect 2014 1178 2020 1179
rect 2086 1178 2093 1179
rect 2110 1178 2116 1179
rect 2130 1178 2136 1179
rect 2183 1179 2184 1180
rect 2188 1179 2189 1183
rect 2279 1183 2285 1184
rect 2279 1179 2280 1183
rect 2284 1182 2285 1183
rect 2294 1183 2300 1184
rect 2294 1182 2295 1183
rect 2284 1180 2295 1182
rect 2284 1179 2285 1180
rect 2183 1178 2189 1179
rect 2206 1178 2212 1179
rect 2279 1178 2285 1179
rect 2294 1179 2295 1180
rect 2299 1179 2300 1183
rect 2322 1183 2328 1184
rect 2322 1179 2323 1183
rect 2327 1182 2328 1183
rect 2375 1183 2381 1184
rect 2375 1182 2376 1183
rect 2327 1180 2376 1182
rect 2327 1179 2328 1180
rect 2294 1178 2300 1179
rect 2302 1178 2308 1179
rect 2322 1178 2328 1179
rect 2375 1179 2376 1180
rect 2380 1179 2381 1183
rect 2375 1178 2381 1179
rect 2398 1178 2404 1179
rect 1598 1174 1599 1178
rect 1603 1174 1604 1178
rect 1598 1173 1604 1174
rect 1702 1174 1703 1178
rect 1707 1174 1708 1178
rect 1702 1173 1708 1174
rect 1806 1174 1807 1178
rect 1811 1174 1812 1178
rect 1806 1173 1812 1174
rect 1910 1174 1911 1178
rect 1915 1174 1916 1178
rect 1910 1173 1916 1174
rect 2014 1174 2015 1178
rect 2019 1174 2020 1178
rect 2014 1173 2020 1174
rect 2110 1174 2111 1178
rect 2115 1174 2116 1178
rect 2110 1173 2116 1174
rect 2206 1174 2207 1178
rect 2211 1174 2212 1178
rect 2206 1173 2212 1174
rect 2302 1174 2303 1178
rect 2307 1174 2308 1178
rect 2302 1173 2308 1174
rect 2398 1174 2399 1178
rect 2403 1174 2404 1178
rect 2398 1173 2404 1174
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 110 1164 116 1165
rect 1326 1169 1332 1170
rect 1326 1165 1327 1169
rect 1331 1165 1332 1169
rect 1326 1164 1332 1165
rect 1366 1169 1372 1170
rect 1366 1165 1367 1169
rect 1371 1165 1372 1169
rect 1366 1164 1372 1165
rect 2582 1169 2588 1170
rect 2582 1165 2583 1169
rect 2587 1165 2588 1169
rect 2582 1164 2588 1165
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1158 140 1159
rect 886 1159 892 1160
rect 139 1156 434 1158
rect 139 1155 140 1156
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 110 1147 116 1148
rect 142 1151 148 1152
rect 142 1147 143 1151
rect 147 1147 148 1151
rect 222 1151 228 1152
rect 142 1146 148 1147
rect 175 1147 181 1148
rect 175 1143 176 1147
rect 180 1146 181 1147
rect 183 1147 189 1148
rect 183 1146 184 1147
rect 180 1144 184 1146
rect 180 1143 181 1144
rect 175 1142 181 1143
rect 183 1143 184 1144
rect 188 1143 189 1147
rect 222 1147 223 1151
rect 227 1147 228 1151
rect 310 1151 316 1152
rect 222 1146 228 1147
rect 255 1147 264 1148
rect 183 1142 189 1143
rect 255 1143 256 1147
rect 263 1143 264 1147
rect 310 1147 311 1151
rect 315 1147 316 1151
rect 406 1151 412 1152
rect 310 1146 316 1147
rect 343 1147 352 1148
rect 255 1142 264 1143
rect 343 1143 344 1147
rect 351 1143 352 1147
rect 406 1147 407 1151
rect 411 1147 412 1151
rect 406 1146 412 1147
rect 432 1146 434 1156
rect 886 1155 887 1159
rect 891 1158 892 1159
rect 1390 1159 1396 1160
rect 891 1156 1074 1158
rect 891 1155 892 1156
rect 886 1154 892 1155
rect 494 1151 500 1152
rect 439 1147 445 1148
rect 439 1146 440 1147
rect 432 1144 440 1146
rect 343 1142 352 1143
rect 439 1143 440 1144
rect 444 1143 445 1147
rect 494 1147 495 1151
rect 499 1147 500 1151
rect 582 1151 588 1152
rect 494 1146 500 1147
rect 527 1147 533 1148
rect 439 1142 445 1143
rect 527 1143 528 1147
rect 532 1146 533 1147
rect 535 1147 541 1148
rect 535 1146 536 1147
rect 532 1144 536 1146
rect 532 1143 533 1144
rect 527 1142 533 1143
rect 535 1143 536 1144
rect 540 1143 541 1147
rect 582 1147 583 1151
rect 587 1147 588 1151
rect 670 1151 676 1152
rect 582 1146 588 1147
rect 615 1147 624 1148
rect 535 1142 541 1143
rect 615 1143 616 1147
rect 623 1143 624 1147
rect 670 1147 671 1151
rect 675 1147 676 1151
rect 750 1151 756 1152
rect 670 1146 676 1147
rect 703 1147 712 1148
rect 615 1142 624 1143
rect 703 1143 704 1147
rect 711 1143 712 1147
rect 750 1147 751 1151
rect 755 1147 756 1151
rect 822 1151 828 1152
rect 750 1146 756 1147
rect 783 1147 792 1148
rect 703 1142 712 1143
rect 783 1143 784 1147
rect 791 1143 792 1147
rect 822 1147 823 1151
rect 827 1147 828 1151
rect 894 1151 900 1152
rect 822 1146 828 1147
rect 855 1147 864 1148
rect 783 1142 792 1143
rect 855 1143 856 1147
rect 863 1143 864 1147
rect 894 1147 895 1151
rect 899 1147 900 1151
rect 966 1151 972 1152
rect 894 1146 900 1147
rect 927 1147 933 1148
rect 927 1146 928 1147
rect 855 1142 864 1143
rect 904 1144 928 1146
rect 678 1139 684 1140
rect 678 1135 679 1139
rect 683 1138 684 1139
rect 904 1138 906 1144
rect 927 1143 928 1144
rect 932 1143 933 1147
rect 966 1147 967 1151
rect 971 1147 972 1151
rect 1046 1151 1052 1152
rect 966 1146 972 1147
rect 999 1147 1008 1148
rect 927 1142 933 1143
rect 999 1143 1000 1147
rect 1007 1143 1008 1147
rect 1046 1147 1047 1151
rect 1051 1147 1052 1151
rect 1046 1146 1052 1147
rect 1072 1146 1074 1156
rect 1390 1155 1391 1159
rect 1395 1158 1396 1159
rect 2086 1159 2092 1160
rect 1395 1156 1521 1158
rect 1395 1155 1396 1156
rect 1390 1154 1396 1155
rect 1326 1152 1332 1153
rect 1326 1148 1327 1152
rect 1331 1148 1332 1152
rect 1079 1147 1085 1148
rect 1326 1147 1332 1148
rect 1366 1152 1372 1153
rect 1366 1148 1367 1152
rect 1371 1148 1372 1152
rect 1366 1147 1372 1148
rect 1398 1151 1404 1152
rect 1398 1147 1399 1151
rect 1403 1147 1404 1151
rect 1486 1151 1492 1152
rect 1079 1146 1080 1147
rect 1072 1144 1080 1146
rect 999 1142 1008 1143
rect 1079 1143 1080 1144
rect 1084 1143 1085 1147
rect 1398 1146 1404 1147
rect 1422 1147 1428 1148
rect 1079 1142 1085 1143
rect 1422 1143 1423 1147
rect 1427 1146 1428 1147
rect 1431 1147 1437 1148
rect 1431 1146 1432 1147
rect 1427 1144 1432 1146
rect 1427 1143 1428 1144
rect 1422 1142 1428 1143
rect 1431 1143 1432 1144
rect 1436 1143 1437 1147
rect 1486 1147 1487 1151
rect 1491 1147 1492 1151
rect 1486 1146 1492 1147
rect 1519 1148 1521 1156
rect 2086 1155 2087 1159
rect 2091 1158 2092 1159
rect 2091 1156 2410 1158
rect 2091 1155 2092 1156
rect 2086 1154 2092 1155
rect 1582 1151 1588 1152
rect 1519 1147 1525 1148
rect 1431 1142 1437 1143
rect 1519 1143 1520 1147
rect 1524 1143 1525 1147
rect 1582 1147 1583 1151
rect 1587 1147 1588 1151
rect 1686 1151 1692 1152
rect 1582 1146 1588 1147
rect 1615 1147 1621 1148
rect 1615 1146 1616 1147
rect 1519 1142 1525 1143
rect 1592 1144 1616 1146
rect 683 1136 906 1138
rect 1494 1139 1500 1140
rect 683 1135 684 1136
rect 678 1134 684 1135
rect 1494 1135 1495 1139
rect 1499 1138 1500 1139
rect 1592 1138 1594 1144
rect 1615 1143 1616 1144
rect 1620 1143 1621 1147
rect 1686 1147 1687 1151
rect 1691 1147 1692 1151
rect 1790 1151 1796 1152
rect 1686 1146 1692 1147
rect 1719 1147 1728 1148
rect 1615 1142 1621 1143
rect 1719 1143 1720 1147
rect 1727 1143 1728 1147
rect 1790 1147 1791 1151
rect 1795 1147 1796 1151
rect 1894 1151 1900 1152
rect 1790 1146 1796 1147
rect 1823 1147 1832 1148
rect 1719 1142 1728 1143
rect 1823 1143 1824 1147
rect 1831 1143 1832 1147
rect 1894 1147 1895 1151
rect 1899 1147 1900 1151
rect 1998 1151 2004 1152
rect 1894 1146 1900 1147
rect 1926 1147 1933 1148
rect 1823 1142 1832 1143
rect 1926 1143 1927 1147
rect 1932 1143 1933 1147
rect 1998 1147 1999 1151
rect 2003 1147 2004 1151
rect 2094 1151 2100 1152
rect 1998 1146 2004 1147
rect 2031 1147 2037 1148
rect 2031 1146 2032 1147
rect 2012 1144 2032 1146
rect 1926 1142 1933 1143
rect 1935 1143 1941 1144
rect 1935 1139 1936 1143
rect 1940 1142 1941 1143
rect 2012 1142 2014 1144
rect 2031 1143 2032 1144
rect 2036 1143 2037 1147
rect 2094 1147 2095 1151
rect 2099 1147 2100 1151
rect 2190 1151 2196 1152
rect 2094 1146 2100 1147
rect 2127 1147 2136 1148
rect 2031 1142 2037 1143
rect 2127 1143 2128 1147
rect 2135 1143 2136 1147
rect 2190 1147 2191 1151
rect 2195 1147 2196 1151
rect 2286 1151 2292 1152
rect 2190 1146 2196 1147
rect 2218 1147 2229 1148
rect 2127 1142 2136 1143
rect 2218 1143 2219 1147
rect 2223 1143 2224 1147
rect 2228 1143 2229 1147
rect 2286 1147 2287 1151
rect 2291 1147 2292 1151
rect 2382 1151 2388 1152
rect 2286 1146 2292 1147
rect 2319 1147 2328 1148
rect 2218 1142 2229 1143
rect 2319 1143 2320 1147
rect 2327 1143 2328 1147
rect 2382 1147 2383 1151
rect 2387 1147 2388 1151
rect 2382 1146 2388 1147
rect 2408 1146 2410 1156
rect 2582 1152 2588 1153
rect 2582 1148 2583 1152
rect 2587 1148 2588 1152
rect 2415 1147 2421 1148
rect 2582 1147 2588 1148
rect 2415 1146 2416 1147
rect 2408 1144 2416 1146
rect 2319 1142 2328 1143
rect 2415 1143 2416 1144
rect 2420 1143 2421 1147
rect 2415 1142 2421 1143
rect 1940 1140 2014 1142
rect 1940 1139 1941 1140
rect 1935 1138 1941 1139
rect 1499 1136 1594 1138
rect 1499 1135 1500 1136
rect 1494 1134 1500 1135
rect 2438 1123 2444 1124
rect 1014 1119 1020 1120
rect 1014 1115 1015 1119
rect 1019 1118 1020 1119
rect 1626 1119 1632 1120
rect 1019 1116 1202 1118
rect 1019 1115 1020 1116
rect 1014 1114 1020 1115
rect 1200 1114 1202 1116
rect 1431 1115 1437 1116
rect 1199 1113 1205 1114
rect 1398 1113 1404 1114
rect 255 1111 261 1112
rect 222 1109 228 1110
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 222 1105 223 1109
rect 227 1105 228 1109
rect 255 1107 256 1111
rect 260 1110 261 1111
rect 310 1111 316 1112
rect 310 1110 311 1111
rect 260 1108 311 1110
rect 260 1107 261 1108
rect 255 1106 261 1107
rect 310 1107 311 1108
rect 315 1107 316 1111
rect 351 1111 360 1112
rect 310 1106 316 1107
rect 318 1109 324 1110
rect 222 1104 228 1105
rect 318 1105 319 1109
rect 323 1105 324 1109
rect 351 1107 352 1111
rect 359 1107 360 1111
rect 455 1111 461 1112
rect 351 1106 360 1107
rect 422 1109 428 1110
rect 318 1104 324 1105
rect 422 1105 423 1109
rect 427 1105 428 1109
rect 455 1107 456 1111
rect 460 1110 461 1111
rect 518 1111 524 1112
rect 518 1110 519 1111
rect 460 1108 519 1110
rect 460 1107 461 1108
rect 455 1106 461 1107
rect 518 1107 519 1108
rect 523 1107 524 1111
rect 550 1111 556 1112
rect 518 1106 524 1107
rect 526 1109 532 1110
rect 422 1104 428 1105
rect 526 1105 527 1109
rect 531 1105 532 1109
rect 550 1107 551 1111
rect 555 1110 556 1111
rect 559 1111 565 1112
rect 559 1110 560 1111
rect 555 1108 560 1110
rect 555 1107 556 1108
rect 550 1106 556 1107
rect 559 1107 560 1108
rect 564 1107 565 1111
rect 663 1111 669 1112
rect 559 1106 565 1107
rect 630 1109 636 1110
rect 526 1104 532 1105
rect 630 1105 631 1109
rect 635 1105 636 1109
rect 663 1107 664 1111
rect 668 1110 669 1111
rect 678 1111 684 1112
rect 678 1110 679 1111
rect 668 1108 679 1110
rect 668 1107 669 1108
rect 663 1106 669 1107
rect 678 1107 679 1108
rect 683 1107 684 1111
rect 759 1111 765 1112
rect 678 1106 684 1107
rect 726 1109 732 1110
rect 630 1104 636 1105
rect 726 1105 727 1109
rect 731 1105 732 1109
rect 759 1107 760 1111
rect 764 1110 765 1111
rect 814 1111 820 1112
rect 814 1110 815 1111
rect 764 1108 815 1110
rect 764 1107 765 1108
rect 759 1106 765 1107
rect 814 1107 815 1108
rect 819 1107 820 1111
rect 855 1111 861 1112
rect 814 1106 820 1107
rect 822 1109 828 1110
rect 726 1104 732 1105
rect 822 1105 823 1109
rect 827 1105 828 1109
rect 855 1107 856 1111
rect 860 1110 861 1111
rect 902 1111 908 1112
rect 902 1110 903 1111
rect 860 1108 903 1110
rect 860 1107 861 1108
rect 855 1106 861 1107
rect 902 1107 903 1108
rect 907 1107 908 1111
rect 943 1111 949 1112
rect 902 1106 908 1107
rect 910 1109 916 1110
rect 822 1104 828 1105
rect 910 1105 911 1109
rect 915 1105 916 1109
rect 943 1107 944 1111
rect 948 1110 949 1111
rect 951 1111 957 1112
rect 951 1110 952 1111
rect 948 1108 952 1110
rect 948 1107 949 1108
rect 943 1106 949 1107
rect 951 1107 952 1108
rect 956 1107 957 1111
rect 1022 1111 1029 1112
rect 951 1106 957 1107
rect 990 1109 996 1110
rect 910 1104 916 1105
rect 990 1105 991 1109
rect 995 1105 996 1109
rect 1022 1107 1023 1111
rect 1028 1107 1029 1111
rect 1111 1111 1117 1112
rect 1022 1106 1029 1107
rect 1078 1109 1084 1110
rect 990 1104 996 1105
rect 1078 1105 1079 1109
rect 1083 1105 1084 1109
rect 1111 1107 1112 1111
rect 1116 1110 1117 1111
rect 1158 1111 1164 1112
rect 1158 1110 1159 1111
rect 1116 1108 1159 1110
rect 1116 1107 1117 1108
rect 1111 1106 1117 1107
rect 1158 1107 1159 1108
rect 1163 1107 1164 1111
rect 1158 1106 1164 1107
rect 1166 1109 1172 1110
rect 1078 1104 1084 1105
rect 1166 1105 1167 1109
rect 1171 1105 1172 1109
rect 1199 1109 1200 1113
rect 1204 1109 1205 1113
rect 1366 1112 1372 1113
rect 1199 1108 1205 1109
rect 1326 1108 1332 1109
rect 1166 1104 1172 1105
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1366 1108 1367 1112
rect 1371 1108 1372 1112
rect 1398 1109 1399 1113
rect 1403 1109 1404 1113
rect 1431 1111 1432 1115
rect 1436 1114 1437 1115
rect 1470 1115 1476 1116
rect 1470 1114 1471 1115
rect 1436 1112 1471 1114
rect 1436 1111 1437 1112
rect 1431 1110 1437 1111
rect 1470 1111 1471 1112
rect 1475 1111 1476 1115
rect 1502 1115 1508 1116
rect 1470 1110 1476 1111
rect 1478 1113 1484 1114
rect 1398 1108 1404 1109
rect 1478 1109 1479 1113
rect 1483 1109 1484 1113
rect 1502 1111 1503 1115
rect 1507 1114 1508 1115
rect 1511 1115 1517 1116
rect 1511 1114 1512 1115
rect 1507 1112 1512 1114
rect 1507 1111 1508 1112
rect 1502 1110 1508 1111
rect 1511 1111 1512 1112
rect 1516 1111 1517 1115
rect 1615 1115 1624 1116
rect 1511 1110 1517 1111
rect 1582 1113 1588 1114
rect 1478 1108 1484 1109
rect 1582 1109 1583 1113
rect 1587 1109 1588 1113
rect 1615 1111 1616 1115
rect 1623 1111 1624 1115
rect 1626 1115 1627 1119
rect 1631 1118 1632 1119
rect 1727 1119 1733 1120
rect 1631 1116 1714 1118
rect 1631 1115 1632 1116
rect 1626 1114 1632 1115
rect 1712 1114 1714 1116
rect 1719 1115 1725 1116
rect 1719 1114 1720 1115
rect 1615 1110 1624 1111
rect 1686 1113 1692 1114
rect 1582 1108 1588 1109
rect 1686 1109 1687 1113
rect 1691 1109 1692 1113
rect 1712 1112 1720 1114
rect 1719 1111 1720 1112
rect 1724 1111 1725 1115
rect 1727 1115 1728 1119
rect 1732 1118 1733 1119
rect 2294 1119 2300 1120
rect 1732 1116 1827 1118
rect 1732 1115 1733 1116
rect 1727 1114 1733 1115
rect 1823 1115 1829 1116
rect 1719 1110 1725 1111
rect 1790 1113 1796 1114
rect 1686 1108 1692 1109
rect 1790 1109 1791 1113
rect 1795 1109 1796 1113
rect 1823 1111 1824 1115
rect 1828 1111 1829 1115
rect 1919 1115 1925 1116
rect 1823 1110 1829 1111
rect 1886 1113 1892 1114
rect 1790 1108 1796 1109
rect 1886 1109 1887 1113
rect 1891 1109 1892 1113
rect 1919 1111 1920 1115
rect 1924 1114 1925 1115
rect 1966 1115 1972 1116
rect 1966 1114 1967 1115
rect 1924 1112 1967 1114
rect 1924 1111 1925 1112
rect 1919 1110 1925 1111
rect 1966 1111 1967 1112
rect 1971 1111 1972 1115
rect 2007 1115 2013 1116
rect 1966 1110 1972 1111
rect 1974 1113 1980 1114
rect 1886 1108 1892 1109
rect 1974 1109 1975 1113
rect 1979 1109 1980 1113
rect 2007 1111 2008 1115
rect 2012 1114 2013 1115
rect 2038 1115 2044 1116
rect 2038 1114 2039 1115
rect 2012 1112 2039 1114
rect 2012 1111 2013 1112
rect 2007 1110 2013 1111
rect 2038 1111 2039 1112
rect 2043 1111 2044 1115
rect 2095 1115 2101 1116
rect 2038 1110 2044 1111
rect 2062 1113 2068 1114
rect 1974 1108 1980 1109
rect 2062 1109 2063 1113
rect 2067 1109 2068 1113
rect 2095 1111 2096 1115
rect 2100 1114 2101 1115
rect 2134 1115 2140 1116
rect 2134 1114 2135 1115
rect 2100 1112 2135 1114
rect 2100 1111 2101 1112
rect 2095 1110 2101 1111
rect 2134 1111 2135 1112
rect 2139 1111 2140 1115
rect 2175 1115 2181 1116
rect 2134 1110 2140 1111
rect 2142 1113 2148 1114
rect 2062 1108 2068 1109
rect 2142 1109 2143 1113
rect 2147 1109 2148 1113
rect 2175 1111 2176 1115
rect 2180 1114 2181 1115
rect 2206 1115 2212 1116
rect 2206 1114 2207 1115
rect 2180 1112 2207 1114
rect 2180 1111 2181 1112
rect 2175 1110 2181 1111
rect 2206 1111 2207 1112
rect 2211 1111 2212 1115
rect 2247 1115 2253 1116
rect 2206 1110 2212 1111
rect 2214 1113 2220 1114
rect 2142 1108 2148 1109
rect 2214 1109 2215 1113
rect 2219 1109 2220 1113
rect 2247 1111 2248 1115
rect 2252 1114 2253 1115
rect 2270 1115 2276 1116
rect 2270 1114 2271 1115
rect 2252 1112 2271 1114
rect 2252 1111 2253 1112
rect 2247 1110 2253 1111
rect 2270 1111 2271 1112
rect 2275 1111 2276 1115
rect 2294 1115 2295 1119
rect 2299 1118 2300 1119
rect 2383 1119 2389 1120
rect 2299 1116 2306 1118
rect 2299 1115 2300 1116
rect 2294 1114 2300 1115
rect 2304 1114 2306 1116
rect 2311 1115 2317 1116
rect 2311 1114 2312 1115
rect 2270 1110 2276 1111
rect 2278 1113 2284 1114
rect 2214 1108 2220 1109
rect 2278 1109 2279 1113
rect 2283 1109 2284 1113
rect 2304 1112 2312 1114
rect 2311 1111 2312 1112
rect 2316 1111 2317 1115
rect 2374 1115 2381 1116
rect 2311 1110 2317 1111
rect 2342 1113 2348 1114
rect 2278 1108 2284 1109
rect 2342 1109 2343 1113
rect 2347 1109 2348 1113
rect 2374 1111 2375 1115
rect 2380 1111 2381 1115
rect 2383 1115 2384 1119
rect 2388 1118 2389 1119
rect 2438 1119 2439 1123
rect 2443 1122 2444 1123
rect 2443 1120 2563 1122
rect 2443 1119 2444 1120
rect 2438 1118 2444 1119
rect 2388 1116 2434 1118
rect 2561 1116 2563 1120
rect 2388 1115 2389 1116
rect 2383 1114 2389 1115
rect 2432 1114 2434 1116
rect 2439 1115 2445 1116
rect 2439 1114 2440 1115
rect 2374 1110 2381 1111
rect 2406 1113 2412 1114
rect 2342 1108 2348 1109
rect 2406 1109 2407 1113
rect 2411 1109 2412 1113
rect 2432 1112 2440 1114
rect 2439 1111 2440 1112
rect 2444 1111 2445 1115
rect 2503 1115 2509 1116
rect 2439 1110 2445 1111
rect 2470 1113 2476 1114
rect 2406 1108 2412 1109
rect 2470 1109 2471 1113
rect 2475 1109 2476 1113
rect 2503 1111 2504 1115
rect 2508 1114 2509 1115
rect 2518 1115 2524 1116
rect 2518 1114 2519 1115
rect 2508 1112 2519 1114
rect 2508 1111 2509 1112
rect 2503 1110 2509 1111
rect 2518 1111 2519 1112
rect 2523 1111 2524 1115
rect 2559 1115 2565 1116
rect 2518 1110 2524 1111
rect 2526 1113 2532 1114
rect 2470 1108 2476 1109
rect 2526 1109 2527 1113
rect 2531 1109 2532 1113
rect 2559 1111 2560 1115
rect 2564 1111 2565 1115
rect 2559 1110 2565 1111
rect 2582 1112 2588 1113
rect 2526 1108 2532 1109
rect 2582 1108 2583 1112
rect 2587 1108 2588 1112
rect 1366 1107 1372 1108
rect 2582 1107 2588 1108
rect 110 1103 116 1104
rect 1326 1103 1332 1104
rect 1366 1095 1372 1096
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 1326 1091 1332 1092
rect 1326 1087 1327 1091
rect 1331 1087 1332 1091
rect 1366 1091 1367 1095
rect 1371 1091 1372 1095
rect 1366 1090 1372 1091
rect 2582 1095 2588 1096
rect 2582 1091 2583 1095
rect 2587 1091 2588 1095
rect 2582 1090 2588 1091
rect 1326 1086 1332 1087
rect 1414 1086 1420 1087
rect 238 1082 244 1083
rect 238 1078 239 1082
rect 243 1078 244 1082
rect 238 1077 244 1078
rect 334 1082 340 1083
rect 334 1078 335 1082
rect 339 1078 340 1082
rect 334 1077 340 1078
rect 438 1082 444 1083
rect 438 1078 439 1082
rect 443 1078 444 1082
rect 438 1077 444 1078
rect 542 1082 548 1083
rect 542 1078 543 1082
rect 547 1078 548 1082
rect 542 1077 548 1078
rect 646 1082 652 1083
rect 646 1078 647 1082
rect 651 1078 652 1082
rect 646 1077 652 1078
rect 742 1082 748 1083
rect 742 1078 743 1082
rect 747 1078 748 1082
rect 742 1077 748 1078
rect 838 1082 844 1083
rect 838 1078 839 1082
rect 843 1078 844 1082
rect 838 1077 844 1078
rect 926 1082 932 1083
rect 926 1078 927 1082
rect 931 1078 932 1082
rect 926 1077 932 1078
rect 1006 1082 1012 1083
rect 1006 1078 1007 1082
rect 1011 1078 1012 1082
rect 1006 1077 1012 1078
rect 1094 1082 1100 1083
rect 1094 1078 1095 1082
rect 1099 1078 1100 1082
rect 1094 1077 1100 1078
rect 1182 1082 1188 1083
rect 1182 1078 1183 1082
rect 1187 1078 1188 1082
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1494 1086 1500 1087
rect 1494 1082 1495 1086
rect 1499 1082 1500 1086
rect 1494 1081 1500 1082
rect 1598 1086 1604 1087
rect 1598 1082 1599 1086
rect 1603 1082 1604 1086
rect 1598 1081 1604 1082
rect 1702 1086 1708 1087
rect 1702 1082 1703 1086
rect 1707 1082 1708 1086
rect 1702 1081 1708 1082
rect 1806 1086 1812 1087
rect 1806 1082 1807 1086
rect 1811 1082 1812 1086
rect 1806 1081 1812 1082
rect 1902 1086 1908 1087
rect 1902 1082 1903 1086
rect 1907 1082 1908 1086
rect 1902 1081 1908 1082
rect 1990 1086 1996 1087
rect 1990 1082 1991 1086
rect 1995 1082 1996 1086
rect 1990 1081 1996 1082
rect 2078 1086 2084 1087
rect 2078 1082 2079 1086
rect 2083 1082 2084 1086
rect 2078 1081 2084 1082
rect 2158 1086 2164 1087
rect 2158 1082 2159 1086
rect 2163 1082 2164 1086
rect 2158 1081 2164 1082
rect 2230 1086 2236 1087
rect 2230 1082 2231 1086
rect 2235 1082 2236 1086
rect 2230 1081 2236 1082
rect 2294 1086 2300 1087
rect 2294 1082 2295 1086
rect 2299 1082 2300 1086
rect 2294 1081 2300 1082
rect 2358 1086 2364 1087
rect 2358 1082 2359 1086
rect 2363 1082 2364 1086
rect 2358 1081 2364 1082
rect 2422 1086 2428 1087
rect 2422 1082 2423 1086
rect 2427 1082 2428 1086
rect 2422 1081 2428 1082
rect 2486 1086 2492 1087
rect 2486 1082 2487 1086
rect 2491 1082 2492 1086
rect 2486 1081 2492 1082
rect 2542 1086 2548 1087
rect 2542 1082 2543 1086
rect 2547 1082 2548 1086
rect 2542 1081 2548 1082
rect 1182 1077 1188 1078
rect 1391 1079 1397 1080
rect 215 1075 224 1076
rect 215 1071 216 1075
rect 223 1071 224 1075
rect 215 1070 224 1071
rect 310 1075 317 1076
rect 310 1071 311 1075
rect 316 1071 317 1075
rect 310 1070 317 1071
rect 415 1075 421 1076
rect 415 1071 416 1075
rect 420 1074 421 1075
rect 454 1075 460 1076
rect 454 1074 455 1075
rect 420 1072 455 1074
rect 420 1071 421 1072
rect 415 1070 421 1071
rect 454 1071 455 1072
rect 459 1071 460 1075
rect 454 1070 460 1071
rect 518 1075 525 1076
rect 518 1071 519 1075
rect 524 1071 525 1075
rect 518 1070 525 1071
rect 618 1075 629 1076
rect 618 1071 619 1075
rect 623 1071 624 1075
rect 628 1071 629 1075
rect 618 1070 629 1071
rect 719 1075 725 1076
rect 719 1071 720 1075
rect 724 1074 725 1075
rect 814 1075 821 1076
rect 724 1072 810 1074
rect 724 1071 725 1072
rect 719 1070 725 1071
rect 534 1067 540 1068
rect 534 1066 535 1067
rect 319 1064 535 1066
rect 319 1062 321 1064
rect 534 1063 535 1064
rect 539 1063 540 1067
rect 808 1066 810 1072
rect 814 1071 815 1075
rect 820 1071 821 1075
rect 814 1070 821 1071
rect 902 1075 909 1076
rect 902 1071 903 1075
rect 908 1071 909 1075
rect 902 1070 909 1071
rect 983 1075 989 1076
rect 983 1071 984 1075
rect 988 1074 989 1075
rect 1014 1075 1020 1076
rect 1014 1074 1015 1075
rect 988 1072 1015 1074
rect 988 1071 989 1072
rect 983 1070 989 1071
rect 1014 1071 1015 1072
rect 1019 1071 1020 1075
rect 1014 1070 1020 1071
rect 1070 1075 1077 1076
rect 1070 1071 1071 1075
rect 1076 1071 1077 1075
rect 1070 1070 1077 1071
rect 1158 1075 1165 1076
rect 1158 1071 1159 1075
rect 1164 1071 1165 1075
rect 1391 1075 1392 1079
rect 1396 1078 1397 1079
rect 1422 1079 1428 1080
rect 1422 1078 1423 1079
rect 1396 1076 1423 1078
rect 1396 1075 1397 1076
rect 1391 1074 1397 1075
rect 1422 1075 1423 1076
rect 1427 1075 1428 1079
rect 1422 1074 1428 1075
rect 1470 1079 1477 1080
rect 1470 1075 1471 1079
rect 1476 1075 1477 1079
rect 1470 1074 1477 1075
rect 1575 1079 1581 1080
rect 1575 1075 1576 1079
rect 1580 1078 1581 1079
rect 1626 1079 1632 1080
rect 1626 1078 1627 1079
rect 1580 1076 1627 1078
rect 1580 1075 1581 1076
rect 1575 1074 1581 1075
rect 1626 1075 1627 1076
rect 1631 1075 1632 1079
rect 1626 1074 1632 1075
rect 1679 1079 1685 1080
rect 1679 1075 1680 1079
rect 1684 1078 1685 1079
rect 1727 1079 1733 1080
rect 1727 1078 1728 1079
rect 1684 1076 1728 1078
rect 1684 1075 1685 1076
rect 1679 1074 1685 1075
rect 1727 1075 1728 1076
rect 1732 1075 1733 1079
rect 1727 1074 1733 1075
rect 1783 1079 1789 1080
rect 1783 1075 1784 1079
rect 1788 1078 1789 1079
rect 1854 1079 1860 1080
rect 1854 1078 1855 1079
rect 1788 1076 1855 1078
rect 1788 1075 1789 1076
rect 1783 1074 1789 1075
rect 1854 1075 1855 1076
rect 1859 1075 1860 1079
rect 1854 1074 1860 1075
rect 1879 1079 1885 1080
rect 1879 1075 1880 1079
rect 1884 1078 1885 1079
rect 1935 1079 1941 1080
rect 1935 1078 1936 1079
rect 1884 1076 1936 1078
rect 1884 1075 1885 1076
rect 1879 1074 1885 1075
rect 1935 1075 1936 1076
rect 1940 1075 1941 1079
rect 1935 1074 1941 1075
rect 1966 1079 1973 1080
rect 1966 1075 1967 1079
rect 1972 1075 1973 1079
rect 1966 1074 1973 1075
rect 2055 1079 2061 1080
rect 2055 1075 2056 1079
rect 2060 1078 2061 1079
rect 2126 1079 2132 1080
rect 2126 1078 2127 1079
rect 2060 1076 2127 1078
rect 2060 1075 2061 1076
rect 2055 1074 2061 1075
rect 2126 1075 2127 1076
rect 2131 1075 2132 1079
rect 2126 1074 2132 1075
rect 2134 1079 2141 1080
rect 2134 1075 2135 1079
rect 2140 1075 2141 1079
rect 2134 1074 2141 1075
rect 2206 1079 2213 1080
rect 2206 1075 2207 1079
rect 2212 1075 2213 1079
rect 2206 1074 2213 1075
rect 2270 1079 2277 1080
rect 2270 1075 2271 1079
rect 2276 1075 2277 1079
rect 2270 1074 2277 1075
rect 2335 1079 2341 1080
rect 2335 1075 2336 1079
rect 2340 1078 2341 1079
rect 2383 1079 2389 1080
rect 2383 1078 2384 1079
rect 2340 1076 2384 1078
rect 2340 1075 2341 1076
rect 2335 1074 2341 1075
rect 2383 1075 2384 1076
rect 2388 1075 2389 1079
rect 2383 1074 2389 1075
rect 2399 1079 2405 1080
rect 2399 1075 2400 1079
rect 2404 1078 2405 1079
rect 2438 1079 2444 1080
rect 2438 1078 2439 1079
rect 2404 1076 2439 1078
rect 2404 1075 2405 1076
rect 2399 1074 2405 1075
rect 2438 1075 2439 1076
rect 2443 1075 2444 1079
rect 2438 1074 2444 1075
rect 2463 1079 2469 1080
rect 2463 1075 2464 1079
rect 2468 1078 2469 1079
rect 2478 1079 2484 1080
rect 2478 1078 2479 1079
rect 2468 1076 2479 1078
rect 2468 1075 2469 1076
rect 2463 1074 2469 1075
rect 2478 1075 2479 1076
rect 2483 1075 2484 1079
rect 2478 1074 2484 1075
rect 2518 1079 2525 1080
rect 2518 1075 2519 1079
rect 2524 1075 2525 1079
rect 2518 1074 2525 1075
rect 1158 1070 1165 1071
rect 2286 1071 2292 1072
rect 2286 1070 2287 1071
rect 2161 1068 2287 1070
rect 1022 1067 1028 1068
rect 1022 1066 1023 1067
rect 808 1064 1023 1066
rect 534 1062 540 1063
rect 1022 1063 1023 1064
rect 1027 1063 1028 1067
rect 1439 1067 1445 1068
rect 1439 1066 1440 1067
rect 1408 1064 1440 1066
rect 1022 1062 1028 1063
rect 1383 1063 1389 1064
rect 1383 1062 1384 1063
rect 304 1060 321 1062
rect 1280 1060 1384 1062
rect 287 1059 293 1060
rect 287 1055 288 1059
rect 292 1058 293 1059
rect 304 1058 306 1060
rect 292 1056 306 1058
rect 335 1059 341 1060
rect 292 1055 293 1056
rect 335 1055 336 1059
rect 340 1058 341 1059
rect 343 1059 349 1060
rect 343 1058 344 1059
rect 340 1056 344 1058
rect 340 1055 341 1056
rect 287 1054 293 1055
rect 310 1054 316 1055
rect 335 1054 341 1055
rect 343 1055 344 1056
rect 348 1055 349 1059
rect 386 1059 392 1060
rect 386 1055 387 1059
rect 391 1058 392 1059
rect 415 1059 421 1060
rect 415 1058 416 1059
rect 391 1056 416 1058
rect 391 1055 392 1056
rect 343 1054 349 1055
rect 366 1054 372 1055
rect 386 1054 392 1055
rect 415 1055 416 1056
rect 420 1055 421 1059
rect 494 1059 501 1060
rect 494 1055 495 1059
rect 500 1055 501 1059
rect 562 1059 568 1060
rect 562 1055 563 1059
rect 567 1058 568 1059
rect 583 1059 589 1060
rect 583 1058 584 1059
rect 567 1056 584 1058
rect 567 1055 568 1056
rect 415 1054 421 1055
rect 438 1054 444 1055
rect 494 1054 501 1055
rect 518 1054 524 1055
rect 562 1054 568 1055
rect 583 1055 584 1056
rect 588 1055 589 1059
rect 678 1059 685 1060
rect 678 1055 679 1059
rect 684 1055 685 1059
rect 722 1059 728 1060
rect 722 1055 723 1059
rect 727 1058 728 1059
rect 775 1059 781 1060
rect 775 1058 776 1059
rect 727 1056 776 1058
rect 727 1055 728 1056
rect 583 1054 589 1055
rect 606 1054 612 1055
rect 678 1054 685 1055
rect 702 1054 708 1055
rect 722 1054 728 1055
rect 775 1055 776 1056
rect 780 1055 781 1059
rect 863 1059 869 1060
rect 863 1055 864 1059
rect 868 1058 869 1059
rect 878 1059 884 1060
rect 878 1058 879 1059
rect 868 1056 879 1058
rect 868 1055 869 1056
rect 775 1054 781 1055
rect 798 1054 804 1055
rect 863 1054 869 1055
rect 878 1055 879 1056
rect 883 1055 884 1059
rect 906 1059 912 1060
rect 906 1055 907 1059
rect 911 1058 912 1059
rect 951 1059 957 1060
rect 951 1058 952 1059
rect 911 1056 952 1058
rect 911 1055 912 1056
rect 878 1054 884 1055
rect 886 1054 892 1055
rect 906 1054 912 1055
rect 951 1055 952 1056
rect 956 1055 957 1059
rect 994 1059 1000 1060
rect 994 1055 995 1059
rect 999 1058 1000 1059
rect 1031 1059 1037 1060
rect 1031 1058 1032 1059
rect 999 1056 1032 1058
rect 999 1055 1000 1056
rect 951 1054 957 1055
rect 974 1054 980 1055
rect 994 1054 1000 1055
rect 1031 1055 1032 1056
rect 1036 1055 1037 1059
rect 1062 1059 1068 1060
rect 1062 1055 1063 1059
rect 1067 1058 1068 1059
rect 1111 1059 1117 1060
rect 1111 1058 1112 1059
rect 1067 1056 1112 1058
rect 1067 1055 1068 1056
rect 1031 1054 1037 1055
rect 1054 1054 1060 1055
rect 1062 1054 1068 1055
rect 1111 1055 1112 1056
rect 1116 1055 1117 1059
rect 1154 1059 1160 1060
rect 1154 1055 1155 1059
rect 1159 1058 1160 1059
rect 1199 1059 1205 1060
rect 1199 1058 1200 1059
rect 1159 1056 1200 1058
rect 1159 1055 1160 1056
rect 1111 1054 1117 1055
rect 1134 1054 1140 1055
rect 1154 1054 1160 1055
rect 1199 1055 1200 1056
rect 1204 1055 1205 1059
rect 1263 1059 1269 1060
rect 1263 1055 1264 1059
rect 1268 1058 1269 1059
rect 1280 1058 1282 1060
rect 1383 1059 1384 1060
rect 1388 1059 1389 1063
rect 1383 1058 1389 1059
rect 1391 1063 1397 1064
rect 1391 1059 1392 1063
rect 1396 1062 1397 1063
rect 1408 1062 1410 1064
rect 1439 1063 1440 1064
rect 1444 1063 1445 1067
rect 1502 1067 1508 1068
rect 1502 1066 1503 1067
rect 1464 1064 1503 1066
rect 1439 1062 1445 1063
rect 1447 1063 1453 1064
rect 1396 1060 1410 1062
rect 1396 1059 1397 1060
rect 1447 1059 1448 1063
rect 1452 1062 1453 1063
rect 1464 1062 1466 1064
rect 1502 1063 1503 1064
rect 1507 1063 1508 1067
rect 1502 1062 1508 1063
rect 1511 1063 1517 1064
rect 1452 1060 1466 1062
rect 1452 1059 1453 1060
rect 1511 1059 1512 1063
rect 1516 1062 1517 1063
rect 1526 1063 1532 1064
rect 1526 1062 1527 1063
rect 1516 1060 1527 1062
rect 1516 1059 1517 1060
rect 1391 1058 1397 1059
rect 1414 1058 1420 1059
rect 1447 1058 1453 1059
rect 1470 1058 1476 1059
rect 1511 1058 1517 1059
rect 1526 1059 1527 1060
rect 1531 1059 1532 1063
rect 1554 1063 1560 1064
rect 1554 1059 1555 1063
rect 1559 1062 1560 1063
rect 1599 1063 1605 1064
rect 1599 1062 1600 1063
rect 1559 1060 1600 1062
rect 1559 1059 1560 1060
rect 1526 1058 1532 1059
rect 1534 1058 1540 1059
rect 1554 1058 1560 1059
rect 1599 1059 1600 1060
rect 1604 1059 1605 1063
rect 1642 1063 1648 1064
rect 1642 1059 1643 1063
rect 1647 1062 1648 1063
rect 1703 1063 1709 1064
rect 1703 1062 1704 1063
rect 1647 1060 1704 1062
rect 1647 1059 1648 1060
rect 1599 1058 1605 1059
rect 1622 1058 1628 1059
rect 1642 1058 1648 1059
rect 1703 1059 1704 1060
rect 1708 1059 1709 1063
rect 1746 1063 1752 1064
rect 1746 1059 1747 1063
rect 1751 1062 1752 1063
rect 1815 1063 1821 1064
rect 1815 1062 1816 1063
rect 1751 1060 1816 1062
rect 1751 1059 1752 1060
rect 1703 1058 1709 1059
rect 1726 1058 1732 1059
rect 1746 1058 1752 1059
rect 1815 1059 1816 1060
rect 1820 1059 1821 1063
rect 1926 1063 1933 1064
rect 1926 1059 1927 1063
rect 1932 1059 1933 1063
rect 2038 1063 2045 1064
rect 2038 1059 2039 1063
rect 2044 1059 2045 1063
rect 2143 1063 2149 1064
rect 2143 1059 2144 1063
rect 2148 1062 2149 1063
rect 2161 1062 2163 1068
rect 2286 1067 2287 1068
rect 2291 1067 2292 1071
rect 2286 1066 2292 1067
rect 2374 1067 2380 1068
rect 2374 1066 2375 1067
rect 2360 1064 2375 1066
rect 2148 1060 2163 1062
rect 2246 1063 2253 1064
rect 2148 1059 2149 1060
rect 2246 1059 2247 1063
rect 2252 1059 2253 1063
rect 2343 1063 2349 1064
rect 2343 1059 2344 1063
rect 2348 1062 2349 1063
rect 2360 1062 2362 1064
rect 2374 1063 2375 1064
rect 2379 1063 2380 1067
rect 2374 1062 2380 1063
rect 2438 1063 2445 1064
rect 2348 1060 2362 1062
rect 2348 1059 2349 1060
rect 2438 1059 2439 1063
rect 2444 1059 2445 1063
rect 2519 1063 2525 1064
rect 2519 1059 2520 1063
rect 2524 1062 2525 1063
rect 2534 1063 2540 1064
rect 2534 1062 2535 1063
rect 2524 1060 2535 1062
rect 2524 1059 2525 1060
rect 1815 1058 1821 1059
rect 1838 1058 1844 1059
rect 1926 1058 1933 1059
rect 1950 1058 1956 1059
rect 2038 1058 2045 1059
rect 2062 1058 2068 1059
rect 2143 1058 2149 1059
rect 2166 1058 2172 1059
rect 2246 1058 2253 1059
rect 2270 1058 2276 1059
rect 2343 1058 2349 1059
rect 2366 1058 2372 1059
rect 2438 1058 2445 1059
rect 2462 1058 2468 1059
rect 2519 1058 2525 1059
rect 2534 1059 2535 1060
rect 2539 1059 2540 1063
rect 2534 1058 2540 1059
rect 2542 1058 2548 1059
rect 1268 1056 1282 1058
rect 1268 1055 1269 1056
rect 1199 1054 1205 1055
rect 1222 1054 1228 1055
rect 1263 1054 1269 1055
rect 1286 1054 1292 1055
rect 310 1050 311 1054
rect 315 1050 316 1054
rect 310 1049 316 1050
rect 366 1050 367 1054
rect 371 1050 372 1054
rect 366 1049 372 1050
rect 438 1050 439 1054
rect 443 1050 444 1054
rect 438 1049 444 1050
rect 518 1050 519 1054
rect 523 1050 524 1054
rect 518 1049 524 1050
rect 606 1050 607 1054
rect 611 1050 612 1054
rect 606 1049 612 1050
rect 702 1050 703 1054
rect 707 1050 708 1054
rect 702 1049 708 1050
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 886 1050 887 1054
rect 891 1050 892 1054
rect 886 1049 892 1050
rect 974 1050 975 1054
rect 979 1050 980 1054
rect 974 1049 980 1050
rect 1054 1050 1055 1054
rect 1059 1050 1060 1054
rect 1054 1049 1060 1050
rect 1134 1050 1135 1054
rect 1139 1050 1140 1054
rect 1134 1049 1140 1050
rect 1222 1050 1223 1054
rect 1227 1050 1228 1054
rect 1222 1049 1228 1050
rect 1286 1050 1287 1054
rect 1291 1050 1292 1054
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1470 1054 1471 1058
rect 1475 1054 1476 1058
rect 1470 1053 1476 1054
rect 1534 1054 1535 1058
rect 1539 1054 1540 1058
rect 1534 1053 1540 1054
rect 1622 1054 1623 1058
rect 1627 1054 1628 1058
rect 1622 1053 1628 1054
rect 1726 1054 1727 1058
rect 1731 1054 1732 1058
rect 1726 1053 1732 1054
rect 1838 1054 1839 1058
rect 1843 1054 1844 1058
rect 1838 1053 1844 1054
rect 1950 1054 1951 1058
rect 1955 1054 1956 1058
rect 1950 1053 1956 1054
rect 2062 1054 2063 1058
rect 2067 1054 2068 1058
rect 2062 1053 2068 1054
rect 2166 1054 2167 1058
rect 2171 1054 2172 1058
rect 2166 1053 2172 1054
rect 2270 1054 2271 1058
rect 2275 1054 2276 1058
rect 2270 1053 2276 1054
rect 2366 1054 2367 1058
rect 2371 1054 2372 1058
rect 2366 1053 2372 1054
rect 2462 1054 2463 1058
rect 2467 1054 2468 1058
rect 2462 1053 2468 1054
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 1286 1049 1292 1050
rect 1366 1049 1372 1050
rect 110 1045 116 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 1326 1045 1332 1046
rect 1326 1041 1327 1045
rect 1331 1041 1332 1045
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 1326 1040 1332 1041
rect 1926 1039 1932 1040
rect 494 1035 500 1036
rect 494 1031 495 1035
rect 499 1034 500 1035
rect 1926 1035 1927 1039
rect 1931 1038 1932 1039
rect 2246 1039 2252 1040
rect 1931 1036 2074 1038
rect 1931 1035 1932 1036
rect 1926 1034 1932 1035
rect 499 1032 618 1034
rect 499 1031 500 1032
rect 494 1030 500 1031
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 294 1027 300 1028
rect 294 1023 295 1027
rect 299 1023 300 1027
rect 350 1027 356 1028
rect 294 1022 300 1023
rect 327 1023 333 1024
rect 327 1019 328 1023
rect 332 1022 333 1023
rect 335 1023 341 1024
rect 335 1022 336 1023
rect 332 1020 336 1022
rect 332 1019 333 1020
rect 327 1018 333 1019
rect 335 1019 336 1020
rect 340 1019 341 1023
rect 350 1023 351 1027
rect 355 1023 356 1027
rect 422 1027 428 1028
rect 350 1022 356 1023
rect 383 1023 392 1024
rect 335 1018 341 1019
rect 383 1019 384 1023
rect 391 1019 392 1023
rect 422 1023 423 1027
rect 427 1023 428 1027
rect 502 1027 508 1028
rect 422 1022 428 1023
rect 454 1023 461 1024
rect 383 1018 392 1019
rect 454 1019 455 1023
rect 460 1019 461 1023
rect 502 1023 503 1027
rect 507 1023 508 1027
rect 590 1027 596 1028
rect 502 1022 508 1023
rect 534 1023 541 1024
rect 454 1018 461 1019
rect 534 1019 535 1023
rect 540 1019 541 1023
rect 590 1023 591 1027
rect 595 1023 596 1027
rect 590 1022 596 1023
rect 616 1022 618 1032
rect 1366 1032 1372 1033
rect 1326 1028 1332 1029
rect 686 1027 692 1028
rect 623 1023 629 1024
rect 623 1022 624 1023
rect 616 1020 624 1022
rect 534 1018 541 1019
rect 623 1019 624 1020
rect 628 1019 629 1023
rect 686 1023 687 1027
rect 691 1023 692 1027
rect 782 1027 788 1028
rect 686 1022 692 1023
rect 719 1023 728 1024
rect 623 1018 629 1019
rect 719 1019 720 1023
rect 727 1019 728 1023
rect 782 1023 783 1027
rect 787 1023 788 1027
rect 870 1027 876 1028
rect 782 1022 788 1023
rect 815 1023 821 1024
rect 815 1022 816 1023
rect 792 1020 816 1022
rect 719 1018 728 1019
rect 754 1019 760 1020
rect 754 1015 755 1019
rect 759 1018 760 1019
rect 792 1018 794 1020
rect 815 1019 816 1020
rect 820 1019 821 1023
rect 870 1023 871 1027
rect 875 1023 876 1027
rect 958 1027 964 1028
rect 870 1022 876 1023
rect 903 1023 912 1024
rect 815 1018 821 1019
rect 903 1019 904 1023
rect 911 1019 912 1023
rect 958 1023 959 1027
rect 963 1023 964 1027
rect 1038 1027 1044 1028
rect 958 1022 964 1023
rect 991 1023 1000 1024
rect 903 1018 912 1019
rect 991 1019 992 1023
rect 999 1019 1000 1023
rect 1038 1023 1039 1027
rect 1043 1023 1044 1027
rect 1118 1027 1124 1028
rect 1038 1022 1044 1023
rect 1070 1023 1077 1024
rect 991 1018 1000 1019
rect 1070 1019 1071 1023
rect 1076 1019 1077 1023
rect 1118 1023 1119 1027
rect 1123 1023 1124 1027
rect 1206 1027 1212 1028
rect 1118 1022 1124 1023
rect 1151 1023 1160 1024
rect 1070 1018 1077 1019
rect 1151 1019 1152 1023
rect 1159 1019 1160 1023
rect 1206 1023 1207 1027
rect 1211 1023 1212 1027
rect 1270 1027 1276 1028
rect 1206 1022 1212 1023
rect 1234 1023 1245 1024
rect 1151 1018 1160 1019
rect 1234 1019 1235 1023
rect 1239 1019 1240 1023
rect 1244 1019 1245 1023
rect 1270 1023 1271 1027
rect 1275 1023 1276 1027
rect 1326 1024 1327 1028
rect 1331 1024 1332 1028
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1454 1031 1460 1032
rect 1398 1026 1404 1027
rect 1431 1027 1437 1028
rect 1431 1026 1432 1027
rect 1408 1024 1432 1026
rect 1270 1022 1276 1023
rect 1294 1023 1300 1024
rect 1234 1018 1245 1019
rect 1294 1019 1295 1023
rect 1299 1022 1300 1023
rect 1303 1023 1309 1024
rect 1326 1023 1332 1024
rect 1383 1023 1389 1024
rect 1303 1022 1304 1023
rect 1299 1020 1304 1022
rect 1299 1019 1300 1020
rect 1294 1018 1300 1019
rect 1303 1019 1304 1020
rect 1308 1019 1309 1023
rect 1303 1018 1309 1019
rect 1383 1019 1384 1023
rect 1388 1022 1389 1023
rect 1408 1022 1410 1024
rect 1431 1023 1432 1024
rect 1436 1023 1437 1027
rect 1454 1027 1455 1031
rect 1459 1027 1460 1031
rect 1518 1031 1524 1032
rect 1454 1026 1460 1027
rect 1487 1027 1493 1028
rect 1487 1026 1488 1027
rect 1464 1024 1488 1026
rect 1431 1022 1437 1023
rect 1439 1023 1445 1024
rect 1388 1020 1410 1022
rect 1388 1019 1389 1020
rect 1383 1018 1389 1019
rect 1439 1019 1440 1023
rect 1444 1022 1445 1023
rect 1464 1022 1466 1024
rect 1487 1023 1488 1024
rect 1492 1023 1493 1027
rect 1518 1027 1519 1031
rect 1523 1027 1524 1031
rect 1606 1031 1612 1032
rect 1518 1026 1524 1027
rect 1551 1027 1560 1028
rect 1487 1022 1493 1023
rect 1551 1023 1552 1027
rect 1559 1023 1560 1027
rect 1606 1027 1607 1031
rect 1611 1027 1612 1031
rect 1710 1031 1716 1032
rect 1606 1026 1612 1027
rect 1639 1027 1648 1028
rect 1551 1022 1560 1023
rect 1639 1023 1640 1027
rect 1647 1023 1648 1027
rect 1710 1027 1711 1031
rect 1715 1027 1716 1031
rect 1822 1031 1828 1032
rect 1710 1026 1716 1027
rect 1743 1027 1752 1028
rect 1639 1022 1648 1023
rect 1743 1023 1744 1027
rect 1751 1023 1752 1027
rect 1822 1027 1823 1031
rect 1827 1027 1828 1031
rect 1934 1031 1940 1032
rect 1822 1026 1828 1027
rect 1854 1027 1861 1028
rect 1743 1022 1752 1023
rect 1854 1023 1855 1027
rect 1860 1023 1861 1027
rect 1934 1027 1935 1031
rect 1939 1027 1940 1031
rect 2046 1031 2052 1032
rect 1934 1026 1940 1027
rect 1967 1027 1973 1028
rect 1967 1026 1968 1027
rect 1944 1024 1968 1026
rect 1854 1022 1861 1023
rect 1863 1023 1869 1024
rect 1444 1020 1466 1022
rect 1444 1019 1445 1020
rect 1439 1018 1445 1019
rect 1863 1019 1864 1023
rect 1868 1022 1869 1023
rect 1944 1022 1946 1024
rect 1967 1023 1968 1024
rect 1972 1023 1973 1027
rect 2046 1027 2047 1031
rect 2051 1027 2052 1031
rect 2046 1026 2052 1027
rect 2072 1026 2074 1036
rect 2246 1035 2247 1039
rect 2251 1038 2252 1039
rect 2438 1039 2444 1040
rect 2251 1036 2378 1038
rect 2251 1035 2252 1036
rect 2246 1034 2252 1035
rect 2150 1031 2156 1032
rect 2079 1027 2085 1028
rect 2079 1026 2080 1027
rect 2072 1024 2080 1026
rect 1967 1022 1973 1023
rect 2079 1023 2080 1024
rect 2084 1023 2085 1027
rect 2150 1027 2151 1031
rect 2155 1027 2156 1031
rect 2254 1031 2260 1032
rect 2150 1026 2156 1027
rect 2183 1027 2189 1028
rect 2183 1026 2184 1027
rect 2160 1024 2184 1026
rect 2079 1022 2085 1023
rect 2126 1023 2132 1024
rect 1868 1020 1946 1022
rect 1868 1019 1869 1020
rect 1863 1018 1869 1019
rect 2126 1019 2127 1023
rect 2131 1022 2132 1023
rect 2160 1022 2162 1024
rect 2183 1023 2184 1024
rect 2188 1023 2189 1027
rect 2254 1027 2255 1031
rect 2259 1027 2260 1031
rect 2350 1031 2356 1032
rect 2254 1026 2260 1027
rect 2286 1027 2293 1028
rect 2183 1022 2189 1023
rect 2286 1023 2287 1027
rect 2292 1023 2293 1027
rect 2350 1027 2351 1031
rect 2355 1027 2356 1031
rect 2350 1026 2356 1027
rect 2376 1026 2378 1036
rect 2438 1035 2439 1039
rect 2443 1038 2444 1039
rect 2443 1036 2563 1038
rect 2443 1035 2444 1036
rect 2438 1034 2444 1035
rect 2446 1031 2452 1032
rect 2383 1027 2389 1028
rect 2383 1026 2384 1027
rect 2376 1024 2384 1026
rect 2286 1022 2293 1023
rect 2383 1023 2384 1024
rect 2388 1023 2389 1027
rect 2446 1027 2447 1031
rect 2451 1027 2452 1031
rect 2526 1031 2532 1032
rect 2446 1026 2452 1027
rect 2478 1027 2485 1028
rect 2383 1022 2389 1023
rect 2478 1023 2479 1027
rect 2484 1023 2485 1027
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2561 1028 2563 1036
rect 2582 1032 2588 1033
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2526 1026 2532 1027
rect 2559 1027 2565 1028
rect 2582 1027 2588 1028
rect 2478 1022 2485 1023
rect 2559 1023 2560 1027
rect 2564 1023 2565 1027
rect 2559 1022 2565 1023
rect 2131 1020 2162 1022
rect 2131 1019 2132 1020
rect 2126 1018 2132 1019
rect 759 1016 794 1018
rect 759 1015 760 1016
rect 754 1014 760 1015
rect 946 1011 952 1012
rect 946 1007 947 1011
rect 951 1010 952 1011
rect 1062 1011 1068 1012
rect 1062 1010 1063 1011
rect 951 1008 1063 1010
rect 951 1007 952 1008
rect 946 1006 952 1007
rect 1062 1007 1063 1008
rect 1067 1007 1068 1011
rect 1062 1006 1068 1007
rect 438 999 444 1000
rect 438 995 439 999
rect 443 998 444 999
rect 806 999 812 1000
rect 443 996 618 998
rect 443 995 444 996
rect 438 994 444 995
rect 447 991 453 992
rect 414 989 420 990
rect 110 988 116 989
rect 110 984 111 988
rect 115 984 116 988
rect 414 985 415 989
rect 419 985 420 989
rect 447 987 448 991
rect 452 990 453 991
rect 462 991 468 992
rect 462 990 463 991
rect 452 988 463 990
rect 452 987 453 988
rect 447 986 453 987
rect 462 987 463 988
rect 467 987 468 991
rect 503 991 509 992
rect 462 986 468 987
rect 470 989 476 990
rect 414 984 420 985
rect 470 985 471 989
rect 475 985 476 989
rect 503 987 504 991
rect 508 990 509 991
rect 518 991 524 992
rect 518 990 519 991
rect 508 988 519 990
rect 508 987 509 988
rect 503 986 509 987
rect 518 987 519 988
rect 523 987 524 991
rect 559 991 568 992
rect 518 986 524 987
rect 526 989 532 990
rect 470 984 476 985
rect 526 985 527 989
rect 531 985 532 989
rect 559 987 560 991
rect 567 987 568 991
rect 616 990 618 996
rect 638 995 644 996
rect 623 991 629 992
rect 623 990 624 991
rect 559 986 568 987
rect 590 989 596 990
rect 526 984 532 985
rect 590 985 591 989
rect 595 985 596 989
rect 616 988 624 990
rect 623 987 624 988
rect 628 987 629 991
rect 638 991 639 995
rect 643 994 644 995
rect 806 995 807 999
rect 811 998 812 999
rect 811 996 1002 998
rect 811 995 812 996
rect 806 994 812 995
rect 643 992 682 994
rect 643 991 644 992
rect 638 990 644 991
rect 680 990 682 992
rect 687 991 693 992
rect 687 990 688 991
rect 623 986 629 987
rect 654 989 660 990
rect 590 984 596 985
rect 654 985 655 989
rect 659 985 660 989
rect 680 988 688 990
rect 687 987 688 988
rect 692 987 693 991
rect 746 991 757 992
rect 687 986 693 987
rect 718 989 724 990
rect 654 984 660 985
rect 718 985 719 989
rect 723 985 724 989
rect 746 987 747 991
rect 751 987 752 991
rect 756 987 757 991
rect 815 991 821 992
rect 746 986 757 987
rect 782 989 788 990
rect 718 984 724 985
rect 782 985 783 989
rect 787 985 788 989
rect 815 987 816 991
rect 820 990 821 991
rect 838 991 844 992
rect 838 990 839 991
rect 820 988 839 990
rect 820 987 821 988
rect 815 986 821 987
rect 838 987 839 988
rect 843 987 844 991
rect 879 991 885 992
rect 838 986 844 987
rect 846 989 852 990
rect 782 984 788 985
rect 846 985 847 989
rect 851 985 852 989
rect 879 987 880 991
rect 884 990 885 991
rect 902 991 908 992
rect 902 990 903 991
rect 884 988 903 990
rect 884 987 885 988
rect 879 986 885 987
rect 902 987 903 988
rect 907 987 908 991
rect 943 991 952 992
rect 902 986 908 987
rect 910 989 916 990
rect 846 984 852 985
rect 910 985 911 989
rect 915 985 916 989
rect 943 987 944 991
rect 951 987 952 991
rect 1000 990 1002 996
rect 1015 995 1021 996
rect 1007 991 1013 992
rect 1007 990 1008 991
rect 943 986 952 987
rect 974 989 980 990
rect 910 984 916 985
rect 974 985 975 989
rect 979 985 980 989
rect 1000 988 1008 990
rect 1007 987 1008 988
rect 1012 987 1013 991
rect 1015 991 1016 995
rect 1020 994 1021 995
rect 1079 995 1085 996
rect 1020 992 1066 994
rect 1020 991 1021 992
rect 1015 990 1021 991
rect 1064 990 1066 992
rect 1071 991 1077 992
rect 1071 990 1072 991
rect 1007 986 1013 987
rect 1038 989 1044 990
rect 974 984 980 985
rect 1038 985 1039 989
rect 1043 985 1044 989
rect 1064 988 1072 990
rect 1071 987 1072 988
rect 1076 987 1077 991
rect 1079 991 1080 995
rect 1084 994 1085 995
rect 1143 995 1149 996
rect 1084 992 1130 994
rect 1084 991 1085 992
rect 1079 990 1085 991
rect 1128 990 1130 992
rect 1135 991 1141 992
rect 1135 990 1136 991
rect 1071 986 1077 987
rect 1102 989 1108 990
rect 1038 984 1044 985
rect 1102 985 1103 989
rect 1107 985 1108 989
rect 1128 988 1136 990
rect 1135 987 1136 988
rect 1140 987 1141 991
rect 1143 991 1144 995
rect 1148 994 1149 995
rect 1199 995 1205 996
rect 1148 992 1186 994
rect 1148 991 1149 992
rect 1143 990 1149 991
rect 1184 990 1186 992
rect 1191 991 1197 992
rect 1191 990 1192 991
rect 1135 986 1141 987
rect 1158 989 1164 990
rect 1102 984 1108 985
rect 1158 985 1159 989
rect 1163 985 1164 989
rect 1184 988 1192 990
rect 1191 987 1192 988
rect 1196 987 1197 991
rect 1199 991 1200 995
rect 1204 994 1205 995
rect 1255 995 1261 996
rect 1204 992 1242 994
rect 1204 991 1205 992
rect 1199 990 1205 991
rect 1240 990 1242 992
rect 1247 991 1253 992
rect 1247 990 1248 991
rect 1191 986 1197 987
rect 1214 989 1220 990
rect 1158 984 1164 985
rect 1214 985 1215 989
rect 1219 985 1220 989
rect 1240 988 1248 990
rect 1247 987 1248 988
rect 1252 987 1253 991
rect 1255 991 1256 995
rect 1260 994 1261 995
rect 1260 992 1298 994
rect 1260 991 1261 992
rect 1255 990 1261 991
rect 1296 990 1298 992
rect 1303 991 1309 992
rect 1303 990 1304 991
rect 1247 986 1253 987
rect 1270 989 1276 990
rect 1214 984 1220 985
rect 1270 985 1271 989
rect 1275 985 1276 989
rect 1296 988 1304 990
rect 1303 987 1304 988
rect 1308 987 1309 991
rect 1526 991 1532 992
rect 1303 986 1309 987
rect 1326 988 1332 989
rect 1270 984 1276 985
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1526 987 1527 991
rect 1531 990 1532 991
rect 1531 988 1746 990
rect 1531 987 1532 988
rect 1526 986 1532 987
rect 110 983 116 984
rect 1326 983 1332 984
rect 1431 983 1437 984
rect 1398 981 1404 982
rect 1366 980 1372 981
rect 1366 976 1367 980
rect 1371 976 1372 980
rect 1398 977 1399 981
rect 1403 977 1404 981
rect 1431 979 1432 983
rect 1436 982 1437 983
rect 1446 983 1452 984
rect 1446 982 1447 983
rect 1436 980 1447 982
rect 1436 979 1437 980
rect 1431 978 1437 979
rect 1446 979 1447 980
rect 1451 979 1452 983
rect 1487 983 1493 984
rect 1446 978 1452 979
rect 1454 981 1460 982
rect 1398 976 1404 977
rect 1454 977 1455 981
rect 1459 977 1460 981
rect 1487 979 1488 983
rect 1492 982 1493 983
rect 1502 983 1508 984
rect 1502 982 1503 983
rect 1492 980 1503 982
rect 1492 979 1493 980
rect 1487 978 1493 979
rect 1502 979 1503 980
rect 1507 979 1508 983
rect 1543 983 1549 984
rect 1502 978 1508 979
rect 1510 981 1516 982
rect 1454 976 1460 977
rect 1510 977 1511 981
rect 1515 977 1516 981
rect 1543 979 1544 983
rect 1548 982 1549 983
rect 1558 983 1564 984
rect 1558 982 1559 983
rect 1548 980 1559 982
rect 1548 979 1549 980
rect 1543 978 1549 979
rect 1558 979 1559 980
rect 1563 979 1564 983
rect 1599 983 1605 984
rect 1558 978 1564 979
rect 1566 981 1572 982
rect 1510 976 1516 977
rect 1566 977 1567 981
rect 1571 977 1572 981
rect 1599 979 1600 983
rect 1604 982 1605 983
rect 1630 983 1636 984
rect 1630 982 1631 983
rect 1604 980 1631 982
rect 1604 979 1605 980
rect 1599 978 1605 979
rect 1630 979 1631 980
rect 1635 979 1636 983
rect 1671 983 1677 984
rect 1630 978 1636 979
rect 1638 981 1644 982
rect 1566 976 1572 977
rect 1638 977 1639 981
rect 1643 977 1644 981
rect 1671 979 1672 983
rect 1676 982 1677 983
rect 1710 983 1716 984
rect 1710 982 1711 983
rect 1676 980 1711 982
rect 1676 979 1677 980
rect 1671 978 1677 979
rect 1710 979 1711 980
rect 1715 979 1716 983
rect 1744 982 1746 988
rect 2534 987 2540 988
rect 1751 983 1757 984
rect 1751 982 1752 983
rect 1710 978 1716 979
rect 1718 981 1724 982
rect 1638 976 1644 977
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1744 980 1752 982
rect 1751 979 1752 980
rect 1756 979 1757 983
rect 1839 983 1845 984
rect 1751 978 1757 979
rect 1806 981 1812 982
rect 1718 976 1724 977
rect 1806 977 1807 981
rect 1811 977 1812 981
rect 1839 979 1840 983
rect 1844 982 1845 983
rect 1894 983 1900 984
rect 1894 982 1895 983
rect 1844 980 1895 982
rect 1844 979 1845 980
rect 1839 978 1845 979
rect 1894 979 1895 980
rect 1899 979 1900 983
rect 1935 983 1941 984
rect 1894 978 1900 979
rect 1902 981 1908 982
rect 1806 976 1812 977
rect 1902 977 1903 981
rect 1907 977 1908 981
rect 1935 979 1936 983
rect 1940 982 1941 983
rect 2006 983 2012 984
rect 2006 982 2007 983
rect 1940 980 2007 982
rect 1940 979 1941 980
rect 1935 978 1941 979
rect 2006 979 2007 980
rect 2011 979 2012 983
rect 2047 983 2053 984
rect 2006 978 2012 979
rect 2014 981 2020 982
rect 1902 976 1908 977
rect 2014 977 2015 981
rect 2019 977 2020 981
rect 2047 979 2048 983
rect 2052 982 2053 983
rect 2134 983 2140 984
rect 2134 982 2135 983
rect 2052 980 2135 982
rect 2052 979 2053 980
rect 2047 978 2053 979
rect 2134 979 2135 980
rect 2139 979 2140 983
rect 2175 983 2181 984
rect 2134 978 2140 979
rect 2142 981 2148 982
rect 2014 976 2020 977
rect 2142 977 2143 981
rect 2147 977 2148 981
rect 2175 979 2176 983
rect 2180 982 2181 983
rect 2262 983 2268 984
rect 2262 982 2263 983
rect 2180 980 2263 982
rect 2180 979 2181 980
rect 2175 978 2181 979
rect 2262 979 2263 980
rect 2267 979 2268 983
rect 2294 983 2300 984
rect 2262 978 2268 979
rect 2270 981 2276 982
rect 2142 976 2148 977
rect 2270 977 2271 981
rect 2275 977 2276 981
rect 2294 979 2295 983
rect 2299 982 2300 983
rect 2303 983 2309 984
rect 2303 982 2304 983
rect 2299 980 2304 982
rect 2299 979 2300 980
rect 2294 978 2300 979
rect 2303 979 2304 980
rect 2308 979 2309 983
rect 2439 983 2445 984
rect 2303 978 2309 979
rect 2406 981 2412 982
rect 2270 976 2276 977
rect 2406 977 2407 981
rect 2411 977 2412 981
rect 2439 979 2440 983
rect 2444 982 2445 983
rect 2518 983 2524 984
rect 2518 982 2519 983
rect 2444 980 2519 982
rect 2444 979 2445 980
rect 2439 978 2445 979
rect 2518 979 2519 980
rect 2523 979 2524 983
rect 2534 983 2535 987
rect 2539 986 2540 987
rect 2539 984 2563 986
rect 2539 983 2540 984
rect 2534 982 2540 983
rect 2559 983 2565 984
rect 2518 978 2524 979
rect 2526 981 2532 982
rect 2406 976 2412 977
rect 2526 977 2527 981
rect 2531 977 2532 981
rect 2559 979 2560 983
rect 2564 979 2565 983
rect 2559 978 2565 979
rect 2582 980 2588 981
rect 2526 976 2532 977
rect 2582 976 2583 980
rect 2587 976 2588 980
rect 1366 975 1372 976
rect 2582 975 2588 976
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 1326 971 1332 972
rect 1326 967 1327 971
rect 1331 967 1332 971
rect 1326 966 1332 967
rect 1366 963 1372 964
rect 430 962 436 963
rect 430 958 431 962
rect 435 958 436 962
rect 430 957 436 958
rect 486 962 492 963
rect 486 958 487 962
rect 491 958 492 962
rect 486 957 492 958
rect 542 962 548 963
rect 542 958 543 962
rect 547 958 548 962
rect 542 957 548 958
rect 606 962 612 963
rect 606 958 607 962
rect 611 958 612 962
rect 606 957 612 958
rect 670 962 676 963
rect 670 958 671 962
rect 675 958 676 962
rect 670 957 676 958
rect 734 962 740 963
rect 734 958 735 962
rect 739 958 740 962
rect 734 957 740 958
rect 798 962 804 963
rect 798 958 799 962
rect 803 958 804 962
rect 798 957 804 958
rect 862 962 868 963
rect 862 958 863 962
rect 867 958 868 962
rect 862 957 868 958
rect 926 962 932 963
rect 926 958 927 962
rect 931 958 932 962
rect 926 957 932 958
rect 990 962 996 963
rect 990 958 991 962
rect 995 958 996 962
rect 990 957 996 958
rect 1054 962 1060 963
rect 1054 958 1055 962
rect 1059 958 1060 962
rect 1054 957 1060 958
rect 1118 962 1124 963
rect 1118 958 1119 962
rect 1123 958 1124 962
rect 1118 957 1124 958
rect 1174 962 1180 963
rect 1174 958 1175 962
rect 1179 958 1180 962
rect 1174 957 1180 958
rect 1230 962 1236 963
rect 1230 958 1231 962
rect 1235 958 1236 962
rect 1230 957 1236 958
rect 1286 962 1292 963
rect 1286 958 1287 962
rect 1291 958 1292 962
rect 1366 959 1367 963
rect 1371 959 1372 963
rect 1366 958 1372 959
rect 2582 963 2588 964
rect 2582 959 2583 963
rect 2587 959 2588 963
rect 2582 958 2588 959
rect 1286 957 1292 958
rect 407 955 413 956
rect 407 951 408 955
rect 412 954 413 955
rect 438 955 444 956
rect 438 954 439 955
rect 412 952 439 954
rect 412 951 413 952
rect 407 950 413 951
rect 438 951 439 952
rect 443 951 444 955
rect 438 950 444 951
rect 462 955 469 956
rect 462 951 463 955
rect 468 951 469 955
rect 462 950 469 951
rect 518 955 525 956
rect 518 951 519 955
rect 524 951 525 955
rect 518 950 525 951
rect 583 955 589 956
rect 583 951 584 955
rect 588 954 589 955
rect 638 955 644 956
rect 638 954 639 955
rect 588 952 639 954
rect 588 951 589 952
rect 583 950 589 951
rect 638 951 639 952
rect 643 951 644 955
rect 638 950 644 951
rect 647 955 653 956
rect 647 951 648 955
rect 652 954 653 955
rect 662 955 668 956
rect 662 954 663 955
rect 652 952 663 954
rect 652 951 653 952
rect 647 950 653 951
rect 662 951 663 952
rect 667 951 668 955
rect 662 950 668 951
rect 711 955 717 956
rect 711 951 712 955
rect 716 954 717 955
rect 754 955 760 956
rect 754 954 755 955
rect 716 952 755 954
rect 716 951 717 952
rect 711 950 717 951
rect 754 951 755 952
rect 759 951 760 955
rect 754 950 760 951
rect 775 955 781 956
rect 775 951 776 955
rect 780 954 781 955
rect 806 955 812 956
rect 806 954 807 955
rect 780 952 807 954
rect 780 951 781 952
rect 775 950 781 951
rect 806 951 807 952
rect 811 951 812 955
rect 806 950 812 951
rect 838 955 845 956
rect 838 951 839 955
rect 844 951 845 955
rect 838 950 845 951
rect 902 955 909 956
rect 902 951 903 955
rect 908 951 909 955
rect 902 950 909 951
rect 967 955 973 956
rect 967 951 968 955
rect 972 954 973 955
rect 1015 955 1021 956
rect 1015 954 1016 955
rect 972 952 1016 954
rect 972 951 973 952
rect 967 950 973 951
rect 1015 951 1016 952
rect 1020 951 1021 955
rect 1015 950 1021 951
rect 1031 955 1037 956
rect 1031 951 1032 955
rect 1036 954 1037 955
rect 1079 955 1085 956
rect 1079 954 1080 955
rect 1036 952 1080 954
rect 1036 951 1037 952
rect 1031 950 1037 951
rect 1079 951 1080 952
rect 1084 951 1085 955
rect 1079 950 1085 951
rect 1095 955 1101 956
rect 1095 951 1096 955
rect 1100 954 1101 955
rect 1143 955 1149 956
rect 1143 954 1144 955
rect 1100 952 1144 954
rect 1100 951 1101 952
rect 1095 950 1101 951
rect 1143 951 1144 952
rect 1148 951 1149 955
rect 1143 950 1149 951
rect 1151 955 1157 956
rect 1151 951 1152 955
rect 1156 954 1157 955
rect 1199 955 1205 956
rect 1199 954 1200 955
rect 1156 952 1200 954
rect 1156 951 1157 952
rect 1151 950 1157 951
rect 1199 951 1200 952
rect 1204 951 1205 955
rect 1199 950 1205 951
rect 1207 955 1213 956
rect 1207 951 1208 955
rect 1212 954 1213 955
rect 1255 955 1261 956
rect 1255 954 1256 955
rect 1212 952 1256 954
rect 1212 951 1213 952
rect 1207 950 1213 951
rect 1255 951 1256 952
rect 1260 951 1261 955
rect 1255 950 1261 951
rect 1263 955 1269 956
rect 1263 951 1264 955
rect 1268 954 1269 955
rect 1294 955 1300 956
rect 1294 954 1295 955
rect 1268 952 1295 954
rect 1268 951 1269 952
rect 1263 950 1269 951
rect 1294 951 1295 952
rect 1299 951 1300 955
rect 1294 950 1300 951
rect 1414 954 1420 955
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1414 949 1420 950
rect 1470 954 1476 955
rect 1470 950 1471 954
rect 1475 950 1476 954
rect 1470 949 1476 950
rect 1526 954 1532 955
rect 1526 950 1527 954
rect 1531 950 1532 954
rect 1526 949 1532 950
rect 1582 954 1588 955
rect 1582 950 1583 954
rect 1587 950 1588 954
rect 1582 949 1588 950
rect 1654 954 1660 955
rect 1654 950 1655 954
rect 1659 950 1660 954
rect 1654 949 1660 950
rect 1734 954 1740 955
rect 1734 950 1735 954
rect 1739 950 1740 954
rect 1734 949 1740 950
rect 1822 954 1828 955
rect 1822 950 1823 954
rect 1827 950 1828 954
rect 1822 949 1828 950
rect 1918 954 1924 955
rect 1918 950 1919 954
rect 1923 950 1924 954
rect 1918 949 1924 950
rect 2030 954 2036 955
rect 2030 950 2031 954
rect 2035 950 2036 954
rect 2030 949 2036 950
rect 2158 954 2164 955
rect 2158 950 2159 954
rect 2163 950 2164 954
rect 2158 949 2164 950
rect 2286 954 2292 955
rect 2286 950 2287 954
rect 2291 950 2292 954
rect 2286 949 2292 950
rect 2422 954 2428 955
rect 2422 950 2423 954
rect 2427 950 2428 954
rect 2422 949 2428 950
rect 2542 954 2548 955
rect 2542 950 2543 954
rect 2547 950 2548 954
rect 2542 949 2548 950
rect 1391 947 1397 948
rect 746 943 752 944
rect 746 942 747 943
rect 735 941 747 942
rect 399 939 405 940
rect 399 935 400 939
rect 404 938 405 939
rect 414 939 420 940
rect 414 938 415 939
rect 404 936 415 938
rect 404 935 405 936
rect 399 934 405 935
rect 414 935 415 936
rect 419 935 420 939
rect 442 939 448 940
rect 442 935 443 939
rect 447 938 448 939
rect 455 939 461 940
rect 455 938 456 939
rect 447 936 456 938
rect 447 935 448 936
rect 414 934 420 935
rect 422 934 428 935
rect 442 934 448 935
rect 455 935 456 936
rect 460 935 461 939
rect 498 939 504 940
rect 498 935 499 939
rect 503 938 504 939
rect 511 939 517 940
rect 511 938 512 939
rect 503 936 512 938
rect 503 935 504 936
rect 455 934 461 935
rect 478 934 484 935
rect 498 934 504 935
rect 511 935 512 936
rect 516 935 517 939
rect 554 939 560 940
rect 554 935 555 939
rect 559 938 560 939
rect 567 939 573 940
rect 567 938 568 939
rect 559 936 568 938
rect 559 935 560 936
rect 511 934 517 935
rect 534 934 540 935
rect 554 934 560 935
rect 567 935 568 936
rect 572 935 573 939
rect 615 939 621 940
rect 615 935 616 939
rect 620 938 621 939
rect 623 939 629 940
rect 623 938 624 939
rect 620 936 624 938
rect 620 935 621 936
rect 567 934 573 935
rect 590 934 596 935
rect 615 934 621 935
rect 623 935 624 936
rect 628 935 629 939
rect 678 939 685 940
rect 678 935 679 939
rect 684 935 685 939
rect 735 937 736 941
rect 740 940 747 941
rect 740 937 741 940
rect 746 939 747 940
rect 751 939 752 943
rect 1391 943 1392 947
rect 1396 946 1397 947
rect 1430 947 1436 948
rect 1430 946 1431 947
rect 1396 944 1431 946
rect 1396 943 1397 944
rect 1391 942 1397 943
rect 1430 943 1431 944
rect 1435 943 1436 947
rect 1430 942 1436 943
rect 1446 947 1453 948
rect 1446 943 1447 947
rect 1452 943 1453 947
rect 1446 942 1453 943
rect 1502 947 1509 948
rect 1502 943 1503 947
rect 1508 943 1509 947
rect 1502 942 1509 943
rect 1558 947 1565 948
rect 1558 943 1559 947
rect 1564 943 1565 947
rect 1558 942 1565 943
rect 1630 947 1637 948
rect 1630 943 1631 947
rect 1636 943 1637 947
rect 1630 942 1637 943
rect 1710 947 1717 948
rect 1710 943 1711 947
rect 1716 943 1717 947
rect 1710 942 1717 943
rect 1799 947 1805 948
rect 1799 943 1800 947
rect 1804 946 1805 947
rect 1863 947 1869 948
rect 1863 946 1864 947
rect 1804 944 1864 946
rect 1804 943 1805 944
rect 1799 942 1805 943
rect 1863 943 1864 944
rect 1868 943 1869 947
rect 1863 942 1869 943
rect 1894 947 1901 948
rect 1894 943 1895 947
rect 1900 943 1901 947
rect 1894 942 1901 943
rect 2006 947 2013 948
rect 2006 943 2007 947
rect 2012 943 2013 947
rect 2006 942 2013 943
rect 2134 947 2141 948
rect 2134 943 2135 947
rect 2140 943 2141 947
rect 2134 942 2141 943
rect 2262 947 2269 948
rect 2262 943 2263 947
rect 2268 943 2269 947
rect 2262 942 2269 943
rect 2330 947 2336 948
rect 2330 943 2331 947
rect 2335 946 2336 947
rect 2399 947 2405 948
rect 2399 946 2400 947
rect 2335 944 2400 946
rect 2335 943 2336 944
rect 2330 942 2336 943
rect 2399 943 2400 944
rect 2404 943 2405 947
rect 2399 942 2405 943
rect 2518 947 2525 948
rect 2518 943 2519 947
rect 2524 943 2525 947
rect 2518 942 2525 943
rect 746 938 752 939
rect 778 939 784 940
rect 735 936 741 937
rect 778 935 779 939
rect 783 938 784 939
rect 791 939 797 940
rect 791 938 792 939
rect 783 936 792 938
rect 783 935 784 936
rect 623 934 629 935
rect 646 934 652 935
rect 678 934 685 935
rect 702 934 708 935
rect 422 930 423 934
rect 427 930 428 934
rect 422 929 428 930
rect 478 930 479 934
rect 483 930 484 934
rect 478 929 484 930
rect 534 930 535 934
rect 539 930 540 934
rect 534 929 540 930
rect 590 930 591 934
rect 595 930 596 934
rect 590 929 596 930
rect 646 930 647 934
rect 651 930 652 934
rect 646 929 652 930
rect 702 930 703 934
rect 707 930 708 934
rect 702 929 708 930
rect 758 934 764 935
rect 778 934 784 935
rect 791 935 792 936
rect 796 935 797 939
rect 1486 935 1492 936
rect 791 934 797 935
rect 814 934 820 935
rect 1486 934 1487 935
rect 758 930 759 934
rect 763 930 764 934
rect 758 929 764 930
rect 814 930 815 934
rect 819 930 820 934
rect 814 929 820 930
rect 1408 932 1487 934
rect 1391 927 1397 928
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1391 923 1392 927
rect 1396 926 1397 927
rect 1408 926 1410 932
rect 1486 931 1487 932
rect 1491 931 1492 935
rect 1630 935 1636 936
rect 1630 934 1631 935
rect 1486 930 1492 931
rect 1520 932 1631 934
rect 1396 924 1410 926
rect 1446 927 1453 928
rect 1396 923 1397 924
rect 1446 923 1447 927
rect 1452 923 1453 927
rect 1503 927 1509 928
rect 1503 923 1504 927
rect 1508 926 1509 927
rect 1520 926 1522 932
rect 1630 931 1631 932
rect 1635 931 1636 935
rect 2078 935 2084 936
rect 2078 934 2079 935
rect 1630 930 1636 931
rect 1999 932 2079 934
rect 1999 930 2001 932
rect 2078 931 2079 932
rect 2083 931 2084 935
rect 2294 935 2300 936
rect 2294 934 2295 935
rect 2078 930 2084 931
rect 2161 932 2295 934
rect 1936 928 2001 930
rect 2161 928 2163 932
rect 2294 931 2295 932
rect 2299 931 2300 935
rect 2454 935 2460 936
rect 2454 934 2455 935
rect 2294 930 2300 931
rect 2304 932 2455 934
rect 1508 924 1522 926
rect 1590 927 1597 928
rect 1508 923 1509 924
rect 1590 923 1591 927
rect 1596 923 1597 927
rect 1679 927 1685 928
rect 1679 923 1680 927
rect 1684 926 1685 927
rect 1687 927 1693 928
rect 1687 926 1688 927
rect 1684 924 1688 926
rect 1684 923 1685 924
rect 1391 922 1397 923
rect 1414 922 1420 923
rect 1446 922 1453 923
rect 1470 922 1476 923
rect 1503 922 1509 923
rect 1526 922 1532 923
rect 1590 922 1597 923
rect 1614 922 1620 923
rect 1679 922 1685 923
rect 1687 923 1688 924
rect 1692 923 1693 927
rect 1735 927 1741 928
rect 1735 923 1736 927
rect 1740 926 1741 927
rect 1799 927 1805 928
rect 1799 926 1800 927
rect 1740 924 1800 926
rect 1740 923 1741 924
rect 1687 922 1693 923
rect 1710 922 1716 923
rect 1735 922 1741 923
rect 1799 923 1800 924
rect 1804 923 1805 927
rect 1919 927 1925 928
rect 1919 923 1920 927
rect 1924 926 1925 927
rect 1936 926 1938 928
rect 1924 924 1938 926
rect 2038 927 2045 928
rect 1924 923 1925 924
rect 2038 923 2039 927
rect 2044 923 2045 927
rect 2159 927 2165 928
rect 2159 923 2160 927
rect 2164 923 2165 927
rect 2287 927 2293 928
rect 2287 923 2288 927
rect 2292 926 2293 927
rect 2304 926 2306 932
rect 2454 931 2455 932
rect 2459 931 2460 935
rect 2454 930 2460 931
rect 2292 924 2306 926
rect 2414 927 2421 928
rect 2292 923 2293 924
rect 2414 923 2415 927
rect 2420 923 2421 927
rect 2519 927 2525 928
rect 2519 923 2520 927
rect 2524 926 2525 927
rect 2534 927 2540 928
rect 2534 926 2535 927
rect 2524 924 2535 926
rect 2524 923 2525 924
rect 1799 922 1805 923
rect 1822 922 1828 923
rect 1919 922 1925 923
rect 1942 922 1948 923
rect 2038 922 2045 923
rect 2062 922 2068 923
rect 2159 922 2165 923
rect 2182 922 2188 923
rect 2287 922 2293 923
rect 2310 922 2316 923
rect 2414 922 2421 923
rect 2438 922 2444 923
rect 2519 922 2525 923
rect 2534 923 2535 924
rect 2539 923 2540 927
rect 2534 922 2540 923
rect 2542 922 2548 923
rect 1326 920 1332 921
rect 1414 918 1415 922
rect 1419 918 1420 922
rect 1414 917 1420 918
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1470 917 1476 918
rect 1526 918 1527 922
rect 1531 918 1532 922
rect 1526 917 1532 918
rect 1614 918 1615 922
rect 1619 918 1620 922
rect 1614 917 1620 918
rect 1710 918 1711 922
rect 1715 918 1716 922
rect 1710 917 1716 918
rect 1822 918 1823 922
rect 1827 918 1828 922
rect 1822 917 1828 918
rect 1942 918 1943 922
rect 1947 918 1948 922
rect 1942 917 1948 918
rect 2062 918 2063 922
rect 2067 918 2068 922
rect 2062 917 2068 918
rect 2182 918 2183 922
rect 2187 918 2188 922
rect 2182 917 2188 918
rect 2310 918 2311 922
rect 2315 918 2316 922
rect 2310 917 2316 918
rect 2438 918 2439 922
rect 2443 918 2444 922
rect 2438 917 2444 918
rect 2542 918 2543 922
rect 2547 918 2548 922
rect 2542 917 2548 918
rect 678 915 684 916
rect 678 911 679 915
rect 683 914 684 915
rect 683 912 826 914
rect 683 911 684 912
rect 678 910 684 911
rect 110 908 116 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 462 907 468 908
rect 406 902 412 903
rect 439 903 448 904
rect 439 899 440 903
rect 447 899 448 903
rect 462 903 463 907
rect 467 903 468 907
rect 518 907 524 908
rect 462 902 468 903
rect 495 903 504 904
rect 439 898 448 899
rect 495 899 496 903
rect 503 899 504 903
rect 518 903 519 907
rect 523 903 524 907
rect 574 907 580 908
rect 518 902 524 903
rect 551 903 560 904
rect 495 898 504 899
rect 551 899 552 903
rect 559 899 560 903
rect 574 903 575 907
rect 579 903 580 907
rect 630 907 636 908
rect 574 902 580 903
rect 607 903 613 904
rect 551 898 560 899
rect 607 899 608 903
rect 612 902 613 903
rect 615 903 621 904
rect 615 902 616 903
rect 612 900 616 902
rect 612 899 613 900
rect 607 898 613 899
rect 615 899 616 900
rect 620 899 621 903
rect 630 903 631 907
rect 635 903 636 907
rect 686 907 692 908
rect 630 902 636 903
rect 662 903 669 904
rect 615 898 621 899
rect 662 899 663 903
rect 668 899 669 903
rect 686 903 687 907
rect 691 903 692 907
rect 742 907 748 908
rect 686 902 692 903
rect 719 903 725 904
rect 719 902 720 903
rect 696 900 720 902
rect 662 898 669 899
rect 694 899 700 900
rect 694 895 695 899
rect 699 895 700 899
rect 719 899 720 900
rect 724 899 725 903
rect 742 903 743 907
rect 747 903 748 907
rect 798 907 804 908
rect 742 902 748 903
rect 775 903 784 904
rect 719 898 725 899
rect 775 899 776 903
rect 783 899 784 903
rect 798 903 799 907
rect 803 903 804 907
rect 798 902 804 903
rect 824 902 826 912
rect 1366 913 1372 914
rect 1366 909 1367 913
rect 1371 909 1372 913
rect 1326 908 1332 909
rect 1366 908 1372 909
rect 2582 913 2588 914
rect 2582 909 2583 913
rect 2587 909 2588 913
rect 2582 908 2588 909
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 831 903 837 904
rect 1326 903 1332 904
rect 1446 903 1452 904
rect 831 902 832 903
rect 824 900 832 902
rect 775 898 784 899
rect 831 899 832 900
rect 836 899 837 903
rect 831 898 837 899
rect 1446 899 1447 903
rect 1451 902 1452 903
rect 1590 903 1596 904
rect 1451 900 1538 902
rect 1451 899 1452 900
rect 1446 898 1452 899
rect 694 894 700 895
rect 1366 896 1372 897
rect 1366 892 1367 896
rect 1371 892 1372 896
rect 1366 891 1372 892
rect 1398 895 1404 896
rect 1398 891 1399 895
rect 1403 891 1404 895
rect 1454 895 1460 896
rect 1398 890 1404 891
rect 1430 891 1437 892
rect 1430 887 1431 891
rect 1436 887 1437 891
rect 1454 891 1455 895
rect 1459 891 1460 895
rect 1510 895 1516 896
rect 1454 890 1460 891
rect 1486 891 1493 892
rect 1430 886 1437 887
rect 1486 887 1487 891
rect 1492 887 1493 891
rect 1510 891 1511 895
rect 1515 891 1516 895
rect 1510 890 1516 891
rect 1536 890 1538 900
rect 1590 899 1591 903
rect 1595 902 1596 903
rect 2038 903 2044 904
rect 1595 900 1834 902
rect 1595 899 1596 900
rect 1590 898 1596 899
rect 1598 895 1604 896
rect 1543 891 1549 892
rect 1543 890 1544 891
rect 1536 888 1544 890
rect 1486 886 1493 887
rect 1543 887 1544 888
rect 1548 887 1549 891
rect 1598 891 1599 895
rect 1603 891 1604 895
rect 1694 895 1700 896
rect 1598 890 1604 891
rect 1630 891 1637 892
rect 1543 886 1549 887
rect 1630 887 1631 891
rect 1636 887 1637 891
rect 1694 891 1695 895
rect 1699 891 1700 895
rect 1806 895 1812 896
rect 1694 890 1700 891
rect 1727 891 1733 892
rect 1630 886 1637 887
rect 1727 887 1728 891
rect 1732 890 1733 891
rect 1735 891 1741 892
rect 1735 890 1736 891
rect 1732 888 1736 890
rect 1732 887 1733 888
rect 1727 886 1733 887
rect 1735 887 1736 888
rect 1740 887 1741 891
rect 1806 891 1807 895
rect 1811 891 1812 895
rect 1806 890 1812 891
rect 1832 890 1834 900
rect 2038 899 2039 903
rect 2043 902 2044 903
rect 2414 903 2420 904
rect 2043 900 2194 902
rect 2043 899 2044 900
rect 2038 898 2044 899
rect 1926 895 1932 896
rect 1839 891 1845 892
rect 1839 890 1840 891
rect 1832 888 1840 890
rect 1735 886 1741 887
rect 1839 887 1840 888
rect 1844 887 1845 891
rect 1926 891 1927 895
rect 1931 891 1932 895
rect 2046 895 2052 896
rect 1926 890 1932 891
rect 1950 891 1956 892
rect 1839 886 1845 887
rect 1950 887 1951 891
rect 1955 890 1956 891
rect 1959 891 1965 892
rect 1959 890 1960 891
rect 1955 888 1960 890
rect 1955 887 1956 888
rect 1950 886 1956 887
rect 1959 887 1960 888
rect 1964 887 1965 891
rect 2046 891 2047 895
rect 2051 891 2052 895
rect 2166 895 2172 896
rect 2046 890 2052 891
rect 2078 891 2085 892
rect 1959 886 1965 887
rect 2078 887 2079 891
rect 2084 887 2085 891
rect 2166 891 2167 895
rect 2171 891 2172 895
rect 2166 890 2172 891
rect 2192 890 2194 900
rect 2414 899 2415 903
rect 2419 902 2420 903
rect 2419 900 2563 902
rect 2419 899 2420 900
rect 2414 898 2420 899
rect 2294 895 2300 896
rect 2199 891 2205 892
rect 2199 890 2200 891
rect 2192 888 2200 890
rect 2078 886 2085 887
rect 2199 887 2200 888
rect 2204 887 2205 891
rect 2294 891 2295 895
rect 2299 891 2300 895
rect 2422 895 2428 896
rect 2294 890 2300 891
rect 2327 891 2336 892
rect 2199 886 2205 887
rect 2327 887 2328 891
rect 2335 887 2336 891
rect 2422 891 2423 895
rect 2427 891 2428 895
rect 2526 895 2532 896
rect 2422 890 2428 891
rect 2454 891 2461 892
rect 2327 886 2336 887
rect 2454 887 2455 891
rect 2460 887 2461 891
rect 2526 891 2527 895
rect 2531 891 2532 895
rect 2561 892 2563 900
rect 2582 896 2588 897
rect 2582 892 2583 896
rect 2587 892 2588 896
rect 2526 890 2532 891
rect 2559 891 2565 892
rect 2582 891 2588 892
rect 2454 886 2461 887
rect 2559 887 2560 891
rect 2564 887 2565 891
rect 2559 886 2565 887
rect 414 883 420 884
rect 414 879 415 883
rect 419 882 420 883
rect 419 880 610 882
rect 419 879 420 880
rect 414 878 420 879
rect 311 875 317 876
rect 278 873 284 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 278 869 279 873
rect 283 869 284 873
rect 311 871 312 875
rect 316 874 317 875
rect 326 875 332 876
rect 326 874 327 875
rect 316 872 327 874
rect 316 871 317 872
rect 311 870 317 871
rect 326 871 327 872
rect 331 871 332 875
rect 367 875 373 876
rect 326 870 332 871
rect 334 873 340 874
rect 278 868 284 869
rect 334 869 335 873
rect 339 869 340 873
rect 367 871 368 875
rect 372 874 373 875
rect 382 875 388 876
rect 382 874 383 875
rect 372 872 383 874
rect 372 871 373 872
rect 367 870 373 871
rect 382 871 383 872
rect 387 871 388 875
rect 423 875 429 876
rect 382 870 388 871
rect 390 873 396 874
rect 334 868 340 869
rect 390 869 391 873
rect 395 869 396 873
rect 423 871 424 875
rect 428 874 429 875
rect 446 875 452 876
rect 446 874 447 875
rect 428 872 447 874
rect 428 871 429 872
rect 423 870 429 871
rect 446 871 447 872
rect 451 871 452 875
rect 487 875 493 876
rect 446 870 452 871
rect 454 873 460 874
rect 390 868 396 869
rect 454 869 455 873
rect 459 869 460 873
rect 487 871 488 875
rect 492 874 493 875
rect 510 875 516 876
rect 510 874 511 875
rect 492 872 511 874
rect 492 871 493 872
rect 487 870 493 871
rect 510 871 511 872
rect 515 871 516 875
rect 551 875 557 876
rect 510 870 516 871
rect 518 873 524 874
rect 454 868 460 869
rect 518 869 519 873
rect 523 869 524 873
rect 551 871 552 875
rect 556 874 557 875
rect 574 875 580 876
rect 574 874 575 875
rect 556 872 575 874
rect 556 871 557 872
rect 551 870 557 871
rect 574 871 575 872
rect 579 871 580 875
rect 608 874 610 880
rect 615 875 621 876
rect 615 874 616 875
rect 574 870 580 871
rect 582 873 588 874
rect 518 868 524 869
rect 582 869 583 873
rect 587 869 588 873
rect 608 872 616 874
rect 615 871 616 872
rect 620 871 621 875
rect 679 875 685 876
rect 615 870 621 871
rect 646 873 652 874
rect 582 868 588 869
rect 646 869 647 873
rect 651 869 652 873
rect 679 871 680 875
rect 684 874 685 875
rect 702 875 708 876
rect 702 874 703 875
rect 684 872 703 874
rect 684 871 685 872
rect 679 870 685 871
rect 702 871 703 872
rect 707 871 708 875
rect 743 875 749 876
rect 702 870 708 871
rect 710 873 716 874
rect 646 868 652 869
rect 710 869 711 873
rect 715 869 716 873
rect 743 871 744 875
rect 748 874 749 875
rect 766 875 772 876
rect 766 874 767 875
rect 748 872 767 874
rect 748 871 749 872
rect 743 870 749 871
rect 766 871 767 872
rect 771 871 772 875
rect 807 875 813 876
rect 766 870 772 871
rect 774 873 780 874
rect 710 868 716 869
rect 774 869 775 873
rect 779 869 780 873
rect 807 871 808 875
rect 812 874 813 875
rect 838 875 844 876
rect 838 874 839 875
rect 812 872 839 874
rect 812 871 813 872
rect 807 870 813 871
rect 838 871 839 872
rect 843 871 844 875
rect 879 875 885 876
rect 838 870 844 871
rect 846 873 852 874
rect 774 868 780 869
rect 846 869 847 873
rect 851 869 852 873
rect 879 871 880 875
rect 884 874 885 875
rect 910 875 916 876
rect 910 874 911 875
rect 884 872 911 874
rect 884 871 885 872
rect 879 870 885 871
rect 910 871 911 872
rect 915 871 916 875
rect 942 875 948 876
rect 910 870 916 871
rect 918 873 924 874
rect 846 868 852 869
rect 918 869 919 873
rect 923 869 924 873
rect 942 871 943 875
rect 947 874 948 875
rect 951 875 957 876
rect 951 874 952 875
rect 947 872 952 874
rect 947 871 948 872
rect 942 870 948 871
rect 951 871 952 872
rect 956 871 957 875
rect 951 870 957 871
rect 1326 872 1332 873
rect 918 868 924 869
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 110 867 116 868
rect 1326 867 1332 868
rect 1750 871 1756 872
rect 1750 867 1751 871
rect 1755 870 1756 871
rect 1755 868 1842 870
rect 1755 867 1756 868
rect 1750 866 1756 867
rect 1503 863 1509 864
rect 1470 861 1476 862
rect 1366 860 1372 861
rect 1366 856 1367 860
rect 1371 856 1372 860
rect 1470 857 1471 861
rect 1475 857 1476 861
rect 1503 859 1504 863
rect 1508 862 1509 863
rect 1542 863 1548 864
rect 1542 862 1543 863
rect 1508 860 1543 862
rect 1508 859 1509 860
rect 1503 858 1509 859
rect 1542 859 1543 860
rect 1547 859 1548 863
rect 1583 863 1589 864
rect 1542 858 1548 859
rect 1550 861 1556 862
rect 1470 856 1476 857
rect 1550 857 1551 861
rect 1555 857 1556 861
rect 1583 859 1584 863
rect 1588 862 1589 863
rect 1630 863 1636 864
rect 1630 862 1631 863
rect 1588 860 1631 862
rect 1588 859 1589 860
rect 1583 858 1589 859
rect 1630 859 1631 860
rect 1635 859 1636 863
rect 1671 863 1677 864
rect 1630 858 1636 859
rect 1638 861 1644 862
rect 1550 856 1556 857
rect 1638 857 1639 861
rect 1643 857 1644 861
rect 1671 859 1672 863
rect 1676 862 1677 863
rect 1679 863 1685 864
rect 1679 862 1680 863
rect 1676 860 1680 862
rect 1676 859 1677 860
rect 1671 858 1677 859
rect 1679 859 1680 860
rect 1684 859 1685 863
rect 1758 863 1765 864
rect 1679 858 1685 859
rect 1726 861 1732 862
rect 1638 856 1644 857
rect 1726 857 1727 861
rect 1731 857 1732 861
rect 1758 859 1759 863
rect 1764 859 1765 863
rect 1840 862 1842 868
rect 2534 867 2540 868
rect 1847 863 1853 864
rect 1847 862 1848 863
rect 1758 858 1765 859
rect 1814 861 1820 862
rect 1726 856 1732 857
rect 1814 857 1815 861
rect 1819 857 1820 861
rect 1840 860 1848 862
rect 1847 859 1848 860
rect 1852 859 1853 863
rect 1935 863 1941 864
rect 1847 858 1853 859
rect 1902 861 1908 862
rect 1814 856 1820 857
rect 1902 857 1903 861
rect 1907 857 1908 861
rect 1935 859 1936 863
rect 1940 862 1941 863
rect 1982 863 1988 864
rect 1982 862 1983 863
rect 1940 860 1983 862
rect 1940 859 1941 860
rect 1935 858 1941 859
rect 1982 859 1983 860
rect 1987 859 1988 863
rect 2023 863 2029 864
rect 1982 858 1988 859
rect 1990 861 1996 862
rect 1902 856 1908 857
rect 1990 857 1991 861
rect 1995 857 1996 861
rect 2023 859 2024 863
rect 2028 862 2029 863
rect 2046 863 2052 864
rect 2046 862 2047 863
rect 2028 860 2047 862
rect 2028 859 2029 860
rect 2023 858 2029 859
rect 2046 859 2047 860
rect 2051 859 2052 863
rect 2103 863 2109 864
rect 2046 858 2052 859
rect 2070 861 2076 862
rect 1990 856 1996 857
rect 2070 857 2071 861
rect 2075 857 2076 861
rect 2103 859 2104 863
rect 2108 862 2109 863
rect 2134 863 2140 864
rect 2134 862 2135 863
rect 2108 860 2135 862
rect 2108 859 2109 860
rect 2103 858 2109 859
rect 2134 859 2135 860
rect 2139 859 2140 863
rect 2175 863 2181 864
rect 2134 858 2140 859
rect 2142 861 2148 862
rect 2070 856 2076 857
rect 2142 857 2143 861
rect 2147 857 2148 861
rect 2175 859 2176 863
rect 2180 862 2181 863
rect 2206 863 2212 864
rect 2206 862 2207 863
rect 2180 860 2207 862
rect 2180 859 2181 860
rect 2175 858 2181 859
rect 2206 859 2207 860
rect 2211 859 2212 863
rect 2247 863 2253 864
rect 2206 858 2212 859
rect 2214 861 2220 862
rect 2142 856 2148 857
rect 2214 857 2215 861
rect 2219 857 2220 861
rect 2247 859 2248 863
rect 2252 862 2253 863
rect 2270 863 2276 864
rect 2270 862 2271 863
rect 2252 860 2271 862
rect 2252 859 2253 860
rect 2247 858 2253 859
rect 2270 859 2271 860
rect 2275 859 2276 863
rect 2311 863 2317 864
rect 2270 858 2276 859
rect 2278 861 2284 862
rect 2214 856 2220 857
rect 2278 857 2279 861
rect 2283 857 2284 861
rect 2311 859 2312 863
rect 2316 862 2317 863
rect 2334 863 2340 864
rect 2334 862 2335 863
rect 2316 860 2335 862
rect 2316 859 2317 860
rect 2311 858 2317 859
rect 2334 859 2335 860
rect 2339 859 2340 863
rect 2375 863 2381 864
rect 2334 858 2340 859
rect 2342 861 2348 862
rect 2278 856 2284 857
rect 2342 857 2343 861
rect 2347 857 2348 861
rect 2375 859 2376 863
rect 2380 862 2381 863
rect 2398 863 2404 864
rect 2398 862 2399 863
rect 2380 860 2399 862
rect 2380 859 2381 860
rect 2375 858 2381 859
rect 2398 859 2399 860
rect 2403 859 2404 863
rect 2439 863 2445 864
rect 2398 858 2404 859
rect 2406 861 2412 862
rect 2342 856 2348 857
rect 2406 857 2407 861
rect 2411 857 2412 861
rect 2439 859 2440 863
rect 2444 862 2445 863
rect 2462 863 2468 864
rect 2462 862 2463 863
rect 2444 860 2463 862
rect 2444 859 2445 860
rect 2439 858 2445 859
rect 2462 859 2463 860
rect 2467 859 2468 863
rect 2503 863 2509 864
rect 2462 858 2468 859
rect 2470 861 2476 862
rect 2406 856 2412 857
rect 2470 857 2471 861
rect 2475 857 2476 861
rect 2503 859 2504 863
rect 2508 862 2509 863
rect 2518 863 2524 864
rect 2518 862 2519 863
rect 2508 860 2519 862
rect 2508 859 2509 860
rect 2503 858 2509 859
rect 2518 859 2519 860
rect 2523 859 2524 863
rect 2534 863 2535 867
rect 2539 866 2540 867
rect 2539 864 2563 866
rect 2539 863 2540 864
rect 2534 862 2540 863
rect 2559 863 2565 864
rect 2518 858 2524 859
rect 2526 861 2532 862
rect 2470 856 2476 857
rect 2526 857 2527 861
rect 2531 857 2532 861
rect 2559 859 2560 863
rect 2564 859 2565 863
rect 2559 858 2565 859
rect 2582 860 2588 861
rect 2526 856 2532 857
rect 2582 856 2583 860
rect 2587 856 2588 860
rect 110 855 116 856
rect 110 851 111 855
rect 115 851 116 855
rect 110 850 116 851
rect 1326 855 1332 856
rect 1366 855 1372 856
rect 2582 855 2588 856
rect 1326 851 1327 855
rect 1331 851 1332 855
rect 1326 850 1332 851
rect 294 846 300 847
rect 294 842 295 846
rect 299 842 300 846
rect 294 841 300 842
rect 350 846 356 847
rect 350 842 351 846
rect 355 842 356 846
rect 350 841 356 842
rect 406 846 412 847
rect 406 842 407 846
rect 411 842 412 846
rect 406 841 412 842
rect 470 846 476 847
rect 470 842 471 846
rect 475 842 476 846
rect 470 841 476 842
rect 534 846 540 847
rect 534 842 535 846
rect 539 842 540 846
rect 534 841 540 842
rect 598 846 604 847
rect 598 842 599 846
rect 603 842 604 846
rect 598 841 604 842
rect 662 846 668 847
rect 662 842 663 846
rect 667 842 668 846
rect 662 841 668 842
rect 726 846 732 847
rect 726 842 727 846
rect 731 842 732 846
rect 726 841 732 842
rect 790 846 796 847
rect 790 842 791 846
rect 795 842 796 846
rect 790 841 796 842
rect 862 846 868 847
rect 862 842 863 846
rect 867 842 868 846
rect 862 841 868 842
rect 934 846 940 847
rect 934 842 935 846
rect 939 842 940 846
rect 934 841 940 842
rect 1366 843 1372 844
rect 271 839 277 840
rect 271 835 272 839
rect 276 838 277 839
rect 326 839 333 840
rect 276 836 321 838
rect 276 835 277 836
rect 271 834 277 835
rect 319 830 321 836
rect 326 835 327 839
rect 332 835 333 839
rect 326 834 333 835
rect 382 839 389 840
rect 382 835 383 839
rect 388 835 389 839
rect 382 834 389 835
rect 446 839 453 840
rect 446 835 447 839
rect 452 835 453 839
rect 446 834 453 835
rect 510 839 517 840
rect 510 835 511 839
rect 516 835 517 839
rect 510 834 517 835
rect 574 839 581 840
rect 574 835 575 839
rect 580 835 581 839
rect 574 834 581 835
rect 639 839 645 840
rect 639 835 640 839
rect 644 838 645 839
rect 694 839 700 840
rect 694 838 695 839
rect 644 836 695 838
rect 644 835 645 836
rect 639 834 645 835
rect 694 835 695 836
rect 699 835 700 839
rect 694 834 700 835
rect 702 839 709 840
rect 702 835 703 839
rect 708 835 709 839
rect 702 834 709 835
rect 766 839 773 840
rect 766 835 767 839
rect 772 835 773 839
rect 766 834 773 835
rect 838 839 845 840
rect 838 835 839 839
rect 844 835 845 839
rect 838 834 845 835
rect 910 839 917 840
rect 910 835 911 839
rect 916 835 917 839
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 2582 843 2588 844
rect 2582 839 2583 843
rect 2587 839 2588 843
rect 2582 838 2588 839
rect 910 834 917 835
rect 1486 834 1492 835
rect 590 831 596 832
rect 590 830 591 831
rect 319 828 591 830
rect 590 827 591 828
rect 595 827 596 831
rect 1486 830 1487 834
rect 1491 830 1492 834
rect 1486 829 1492 830
rect 1566 834 1572 835
rect 1566 830 1567 834
rect 1571 830 1572 834
rect 1566 829 1572 830
rect 1654 834 1660 835
rect 1654 830 1655 834
rect 1659 830 1660 834
rect 1654 829 1660 830
rect 1742 834 1748 835
rect 1742 830 1743 834
rect 1747 830 1748 834
rect 1742 829 1748 830
rect 1830 834 1836 835
rect 1830 830 1831 834
rect 1835 830 1836 834
rect 1830 829 1836 830
rect 1918 834 1924 835
rect 1918 830 1919 834
rect 1923 830 1924 834
rect 1918 829 1924 830
rect 2006 834 2012 835
rect 2006 830 2007 834
rect 2011 830 2012 834
rect 2006 829 2012 830
rect 2086 834 2092 835
rect 2086 830 2087 834
rect 2091 830 2092 834
rect 2086 829 2092 830
rect 2158 834 2164 835
rect 2158 830 2159 834
rect 2163 830 2164 834
rect 2158 829 2164 830
rect 2230 834 2236 835
rect 2230 830 2231 834
rect 2235 830 2236 834
rect 2230 829 2236 830
rect 2294 834 2300 835
rect 2294 830 2295 834
rect 2299 830 2300 834
rect 2294 829 2300 830
rect 2358 834 2364 835
rect 2358 830 2359 834
rect 2363 830 2364 834
rect 2358 829 2364 830
rect 2422 834 2428 835
rect 2422 830 2423 834
rect 2427 830 2428 834
rect 2422 829 2428 830
rect 2486 834 2492 835
rect 2486 830 2487 834
rect 2491 830 2492 834
rect 2486 829 2492 830
rect 2542 834 2548 835
rect 2542 830 2543 834
rect 2547 830 2548 834
rect 2542 829 2548 830
rect 590 826 596 827
rect 942 827 948 828
rect 942 826 943 827
rect 649 824 943 826
rect 649 820 651 824
rect 942 823 943 824
rect 947 823 948 827
rect 942 822 948 823
rect 1463 827 1469 828
rect 1463 823 1464 827
rect 1468 826 1469 827
rect 1542 827 1549 828
rect 1468 824 1538 826
rect 1468 823 1469 824
rect 1463 822 1469 823
rect 143 819 149 820
rect 143 815 144 819
rect 148 818 149 819
rect 158 819 164 820
rect 158 818 159 819
rect 148 816 159 818
rect 148 815 149 816
rect 143 814 149 815
rect 158 815 159 816
rect 163 815 164 819
rect 186 819 192 820
rect 186 815 187 819
rect 191 818 192 819
rect 207 819 213 820
rect 207 818 208 819
rect 191 816 208 818
rect 191 815 192 816
rect 158 814 164 815
rect 166 814 172 815
rect 186 814 192 815
rect 207 815 208 816
rect 212 815 213 819
rect 250 819 256 820
rect 250 815 251 819
rect 255 818 256 819
rect 287 819 293 820
rect 287 818 288 819
rect 255 816 288 818
rect 255 815 256 816
rect 207 814 213 815
rect 230 814 236 815
rect 250 814 256 815
rect 287 815 288 816
rect 292 815 293 819
rect 330 819 336 820
rect 330 815 331 819
rect 335 818 336 819
rect 375 819 381 820
rect 375 818 376 819
rect 335 816 376 818
rect 335 815 336 816
rect 287 814 293 815
rect 310 814 316 815
rect 330 814 336 815
rect 375 815 376 816
rect 380 815 381 819
rect 418 819 424 820
rect 418 815 419 819
rect 423 818 424 819
rect 463 819 469 820
rect 463 818 464 819
rect 423 816 464 818
rect 423 815 424 816
rect 375 814 381 815
rect 398 814 404 815
rect 418 814 424 815
rect 463 815 464 816
rect 468 815 469 819
rect 506 819 512 820
rect 506 815 507 819
rect 511 818 512 819
rect 559 819 565 820
rect 559 818 560 819
rect 511 816 560 818
rect 511 815 512 816
rect 463 814 469 815
rect 486 814 492 815
rect 506 814 512 815
rect 559 815 560 816
rect 564 815 565 819
rect 647 819 653 820
rect 647 815 648 819
rect 652 815 653 819
rect 690 819 696 820
rect 690 815 691 819
rect 695 818 696 819
rect 735 819 741 820
rect 735 818 736 819
rect 695 816 736 818
rect 695 815 696 816
rect 559 814 565 815
rect 582 814 588 815
rect 647 814 653 815
rect 670 814 676 815
rect 690 814 696 815
rect 735 815 736 816
rect 740 815 741 819
rect 778 819 784 820
rect 778 815 779 819
rect 783 818 784 819
rect 815 819 821 820
rect 815 818 816 819
rect 783 816 816 818
rect 783 815 784 816
rect 735 814 741 815
rect 758 814 764 815
rect 778 814 784 815
rect 815 815 816 816
rect 820 815 821 819
rect 863 819 869 820
rect 863 815 864 819
rect 868 818 869 819
rect 895 819 901 820
rect 895 818 896 819
rect 868 816 896 818
rect 868 815 869 816
rect 815 814 821 815
rect 838 814 844 815
rect 863 814 869 815
rect 895 815 896 816
rect 900 815 901 819
rect 943 819 949 820
rect 943 815 944 819
rect 948 818 949 819
rect 983 819 989 820
rect 983 818 984 819
rect 948 816 984 818
rect 948 815 949 816
rect 895 814 901 815
rect 918 814 924 815
rect 943 814 949 815
rect 983 815 984 816
rect 988 815 989 819
rect 1026 819 1032 820
rect 1026 815 1027 819
rect 1031 818 1032 819
rect 1071 819 1077 820
rect 1071 818 1072 819
rect 1031 816 1072 818
rect 1031 815 1032 816
rect 983 814 989 815
rect 1006 814 1012 815
rect 1026 814 1032 815
rect 1071 815 1072 816
rect 1076 815 1077 819
rect 1536 818 1538 824
rect 1542 823 1543 827
rect 1548 823 1549 827
rect 1542 822 1549 823
rect 1630 827 1637 828
rect 1630 823 1631 827
rect 1636 823 1637 827
rect 1630 822 1637 823
rect 1719 827 1725 828
rect 1719 823 1720 827
rect 1724 826 1725 827
rect 1750 827 1756 828
rect 1750 826 1751 827
rect 1724 824 1751 826
rect 1724 823 1725 824
rect 1719 822 1725 823
rect 1750 823 1751 824
rect 1755 823 1756 827
rect 1770 827 1776 828
rect 1750 822 1756 823
rect 1758 823 1764 824
rect 1758 819 1759 823
rect 1763 819 1764 823
rect 1770 823 1771 827
rect 1775 826 1776 827
rect 1807 827 1813 828
rect 1807 826 1808 827
rect 1775 824 1808 826
rect 1775 823 1776 824
rect 1770 822 1776 823
rect 1807 823 1808 824
rect 1812 823 1813 827
rect 1807 822 1813 823
rect 1895 827 1901 828
rect 1895 823 1896 827
rect 1900 826 1901 827
rect 1950 827 1956 828
rect 1950 826 1951 827
rect 1900 824 1951 826
rect 1900 823 1901 824
rect 1895 822 1901 823
rect 1950 823 1951 824
rect 1955 823 1956 827
rect 1950 822 1956 823
rect 1982 827 1989 828
rect 1982 823 1983 827
rect 1988 823 1989 827
rect 1982 822 1989 823
rect 2063 827 2069 828
rect 2063 823 2064 827
rect 2068 826 2069 827
rect 2126 827 2132 828
rect 2126 826 2127 827
rect 2068 824 2127 826
rect 2068 823 2069 824
rect 2063 822 2069 823
rect 2126 823 2127 824
rect 2131 823 2132 827
rect 2126 822 2132 823
rect 2134 827 2141 828
rect 2134 823 2135 827
rect 2140 823 2141 827
rect 2134 822 2141 823
rect 2206 827 2213 828
rect 2206 823 2207 827
rect 2212 823 2213 827
rect 2206 822 2213 823
rect 2270 827 2277 828
rect 2270 823 2271 827
rect 2276 823 2277 827
rect 2270 822 2277 823
rect 2334 827 2341 828
rect 2334 823 2335 827
rect 2340 823 2341 827
rect 2334 822 2341 823
rect 2398 827 2405 828
rect 2398 823 2399 827
rect 2404 823 2405 827
rect 2398 822 2405 823
rect 2462 827 2469 828
rect 2462 823 2463 827
rect 2468 823 2469 827
rect 2462 822 2469 823
rect 2518 827 2525 828
rect 2518 823 2519 827
rect 2524 823 2525 827
rect 2518 822 2525 823
rect 1758 818 1764 819
rect 1536 816 1762 818
rect 1838 815 1844 816
rect 1071 814 1077 815
rect 1094 814 1100 815
rect 1838 814 1839 815
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 230 810 231 814
rect 235 810 236 814
rect 230 809 236 810
rect 310 810 311 814
rect 315 810 316 814
rect 310 809 316 810
rect 398 810 399 814
rect 403 810 404 814
rect 398 809 404 810
rect 486 810 487 814
rect 491 810 492 814
rect 486 809 492 810
rect 582 810 583 814
rect 587 810 588 814
rect 582 809 588 810
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 758 810 759 814
rect 763 810 764 814
rect 758 809 764 810
rect 838 810 839 814
rect 843 810 844 814
rect 838 809 844 810
rect 918 810 919 814
rect 923 810 924 814
rect 918 809 924 810
rect 1006 810 1007 814
rect 1011 810 1012 814
rect 1006 809 1012 810
rect 1094 810 1095 814
rect 1099 810 1100 814
rect 1094 809 1100 810
rect 1624 812 1839 814
rect 1607 807 1613 808
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 1326 805 1332 806
rect 1326 801 1327 805
rect 1331 801 1332 805
rect 1607 803 1608 807
rect 1612 806 1613 807
rect 1624 806 1626 812
rect 1838 811 1839 812
rect 1843 811 1844 815
rect 1998 815 2004 816
rect 1998 814 1999 815
rect 1838 810 1844 811
rect 1892 812 1999 814
rect 1612 804 1626 806
rect 1655 807 1661 808
rect 1612 803 1613 804
rect 1655 803 1656 807
rect 1660 806 1661 807
rect 1663 807 1669 808
rect 1663 806 1664 807
rect 1660 804 1664 806
rect 1660 803 1661 804
rect 1607 802 1613 803
rect 1630 802 1636 803
rect 1655 802 1661 803
rect 1663 803 1664 804
rect 1668 803 1669 807
rect 1706 807 1712 808
rect 1706 803 1707 807
rect 1711 806 1712 807
rect 1727 807 1733 808
rect 1727 806 1728 807
rect 1711 804 1728 806
rect 1711 803 1712 804
rect 1663 802 1669 803
rect 1686 802 1692 803
rect 1706 802 1712 803
rect 1727 803 1728 804
rect 1732 803 1733 807
rect 1798 807 1805 808
rect 1798 803 1799 807
rect 1804 803 1805 807
rect 1879 807 1885 808
rect 1879 803 1880 807
rect 1884 806 1885 807
rect 1892 806 1894 812
rect 1998 811 1999 812
rect 2003 811 2004 815
rect 1998 810 2004 811
rect 1884 804 1894 806
rect 1959 807 1965 808
rect 1884 803 1885 804
rect 1959 803 1960 807
rect 1964 806 1965 807
rect 1967 807 1973 808
rect 1967 806 1968 807
rect 1964 804 1968 806
rect 1964 803 1965 804
rect 1727 802 1733 803
rect 1750 802 1756 803
rect 1798 802 1805 803
rect 1822 802 1828 803
rect 1879 802 1885 803
rect 1902 802 1908 803
rect 1959 802 1965 803
rect 1967 803 1968 804
rect 1972 803 1973 807
rect 2046 807 2053 808
rect 2046 803 2047 807
rect 2052 803 2053 807
rect 2135 807 2141 808
rect 2135 803 2136 807
rect 2140 806 2141 807
rect 2150 807 2156 808
rect 2150 806 2151 807
rect 2140 804 2151 806
rect 2140 803 2141 804
rect 1967 802 1973 803
rect 1990 802 1996 803
rect 2046 802 2053 803
rect 2070 802 2076 803
rect 2135 802 2141 803
rect 2150 803 2151 804
rect 2155 803 2156 807
rect 2178 807 2184 808
rect 2178 803 2179 807
rect 2183 806 2184 807
rect 2223 807 2229 808
rect 2223 806 2224 807
rect 2183 804 2224 806
rect 2183 803 2184 804
rect 2150 802 2156 803
rect 2158 802 2164 803
rect 2178 802 2184 803
rect 2223 803 2224 804
rect 2228 803 2229 807
rect 2266 807 2272 808
rect 2266 803 2267 807
rect 2271 806 2272 807
rect 2311 807 2317 808
rect 2311 806 2312 807
rect 2271 804 2312 806
rect 2271 803 2272 804
rect 2223 802 2229 803
rect 2246 802 2252 803
rect 2266 802 2272 803
rect 2311 803 2312 804
rect 2316 803 2317 807
rect 2359 807 2365 808
rect 2359 803 2360 807
rect 2364 806 2365 807
rect 2399 807 2405 808
rect 2399 806 2400 807
rect 2364 804 2400 806
rect 2364 803 2365 804
rect 2311 802 2317 803
rect 2334 802 2340 803
rect 2359 802 2365 803
rect 2399 803 2400 804
rect 2404 803 2405 807
rect 2399 802 2405 803
rect 2422 802 2428 803
rect 1326 800 1332 801
rect 1630 798 1631 802
rect 1635 798 1636 802
rect 1630 797 1636 798
rect 1686 798 1687 802
rect 1691 798 1692 802
rect 1686 797 1692 798
rect 1750 798 1751 802
rect 1755 798 1756 802
rect 1750 797 1756 798
rect 1822 798 1823 802
rect 1827 798 1828 802
rect 1822 797 1828 798
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 1990 798 1991 802
rect 1995 798 1996 802
rect 1990 797 1996 798
rect 2070 798 2071 802
rect 2075 798 2076 802
rect 2070 797 2076 798
rect 2158 798 2159 802
rect 2163 798 2164 802
rect 2158 797 2164 798
rect 2246 798 2247 802
rect 2251 798 2252 802
rect 2246 797 2252 798
rect 2334 798 2335 802
rect 2339 798 2340 802
rect 2334 797 2340 798
rect 2422 798 2423 802
rect 2427 798 2428 802
rect 2422 797 2428 798
rect 1366 793 1372 794
rect 1366 789 1367 793
rect 1371 789 1372 793
rect 110 788 116 789
rect 1326 788 1332 789
rect 1366 788 1372 789
rect 2582 793 2588 794
rect 2582 789 2583 793
rect 2587 789 2588 793
rect 2582 788 2588 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 150 787 156 788
rect 150 783 151 787
rect 155 783 156 787
rect 214 787 220 788
rect 150 782 156 783
rect 183 783 192 784
rect 183 779 184 783
rect 191 779 192 783
rect 214 783 215 787
rect 219 783 220 787
rect 294 787 300 788
rect 214 782 220 783
rect 247 783 256 784
rect 183 778 192 779
rect 247 779 248 783
rect 255 779 256 783
rect 294 783 295 787
rect 299 783 300 787
rect 382 787 388 788
rect 294 782 300 783
rect 327 783 336 784
rect 247 778 256 779
rect 327 779 328 783
rect 335 779 336 783
rect 382 783 383 787
rect 387 783 388 787
rect 470 787 476 788
rect 382 782 388 783
rect 415 783 424 784
rect 327 778 336 779
rect 415 779 416 783
rect 423 779 424 783
rect 470 783 471 787
rect 475 783 476 787
rect 566 787 572 788
rect 470 782 476 783
rect 503 783 512 784
rect 415 778 424 779
rect 503 779 504 783
rect 511 779 512 783
rect 566 783 567 787
rect 571 783 572 787
rect 654 787 660 788
rect 566 782 572 783
rect 590 783 596 784
rect 503 778 512 779
rect 590 779 591 783
rect 595 782 596 783
rect 599 783 605 784
rect 599 782 600 783
rect 595 780 600 782
rect 595 779 596 780
rect 590 778 596 779
rect 599 779 600 780
rect 604 779 605 783
rect 654 783 655 787
rect 659 783 660 787
rect 742 787 748 788
rect 654 782 660 783
rect 687 783 696 784
rect 599 778 605 779
rect 687 779 688 783
rect 695 779 696 783
rect 742 783 743 787
rect 747 783 748 787
rect 822 787 828 788
rect 742 782 748 783
rect 775 783 784 784
rect 687 778 696 779
rect 775 779 776 783
rect 783 779 784 783
rect 822 783 823 787
rect 827 783 828 787
rect 902 787 908 788
rect 822 782 828 783
rect 855 783 861 784
rect 775 778 784 779
rect 855 779 856 783
rect 860 782 861 783
rect 863 783 869 784
rect 863 782 864 783
rect 860 780 864 782
rect 860 779 861 780
rect 855 778 861 779
rect 863 779 864 780
rect 868 779 869 783
rect 902 783 903 787
rect 907 783 908 787
rect 943 787 949 788
rect 943 786 944 787
rect 902 782 908 783
rect 935 785 944 786
rect 935 781 936 785
rect 940 784 944 785
rect 940 781 941 784
rect 943 783 944 784
rect 948 783 949 787
rect 943 782 949 783
rect 990 787 996 788
rect 990 783 991 787
rect 995 783 996 787
rect 1078 787 1084 788
rect 990 782 996 783
rect 1023 783 1032 784
rect 935 780 941 781
rect 863 778 869 779
rect 1023 779 1024 783
rect 1031 779 1032 783
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1326 784 1327 788
rect 1331 784 1332 788
rect 1078 782 1084 783
rect 1102 783 1108 784
rect 1023 778 1032 779
rect 1102 779 1103 783
rect 1107 782 1108 783
rect 1111 783 1117 784
rect 1326 783 1332 784
rect 1798 783 1804 784
rect 1111 782 1112 783
rect 1107 780 1112 782
rect 1107 779 1108 780
rect 1102 778 1108 779
rect 1111 779 1112 780
rect 1116 779 1117 783
rect 1111 778 1117 779
rect 1798 779 1799 783
rect 1803 782 1804 783
rect 1803 780 1914 782
rect 1803 779 1804 780
rect 1798 778 1804 779
rect 1366 776 1372 777
rect 1366 772 1367 776
rect 1371 772 1372 776
rect 1366 771 1372 772
rect 1614 775 1620 776
rect 1614 771 1615 775
rect 1619 771 1620 775
rect 1670 775 1676 776
rect 1614 770 1620 771
rect 1647 771 1653 772
rect 1647 767 1648 771
rect 1652 770 1653 771
rect 1655 771 1661 772
rect 1655 770 1656 771
rect 1652 768 1656 770
rect 1652 767 1653 768
rect 1647 766 1653 767
rect 1655 767 1656 768
rect 1660 767 1661 771
rect 1670 771 1671 775
rect 1675 771 1676 775
rect 1734 775 1740 776
rect 1670 770 1676 771
rect 1703 771 1712 772
rect 1655 766 1661 767
rect 1703 767 1704 771
rect 1711 767 1712 771
rect 1734 771 1735 775
rect 1739 771 1740 775
rect 1806 775 1812 776
rect 1734 770 1740 771
rect 1767 771 1776 772
rect 1703 766 1712 767
rect 1767 767 1768 771
rect 1775 767 1776 771
rect 1806 771 1807 775
rect 1811 771 1812 775
rect 1886 775 1892 776
rect 1806 770 1812 771
rect 1838 771 1845 772
rect 1767 766 1776 767
rect 1838 767 1839 771
rect 1844 767 1845 771
rect 1886 771 1887 775
rect 1891 771 1892 775
rect 1886 770 1892 771
rect 1912 770 1914 780
rect 2582 776 2588 777
rect 1974 775 1980 776
rect 1919 771 1925 772
rect 1919 770 1920 771
rect 1912 768 1920 770
rect 1838 766 1845 767
rect 1919 767 1920 768
rect 1924 767 1925 771
rect 1974 771 1975 775
rect 1979 771 1980 775
rect 2054 775 2060 776
rect 1974 770 1980 771
rect 1998 771 2004 772
rect 1919 766 1925 767
rect 1998 767 1999 771
rect 2003 770 2004 771
rect 2007 771 2013 772
rect 2007 770 2008 771
rect 2003 768 2008 770
rect 2003 767 2004 768
rect 1998 766 2004 767
rect 2007 767 2008 768
rect 2012 767 2013 771
rect 2054 771 2055 775
rect 2059 771 2060 775
rect 2142 775 2148 776
rect 2054 770 2060 771
rect 2086 771 2093 772
rect 2007 766 2013 767
rect 2086 767 2087 771
rect 2092 767 2093 771
rect 2142 771 2143 775
rect 2147 771 2148 775
rect 2230 775 2236 776
rect 2142 770 2148 771
rect 2175 771 2184 772
rect 2086 766 2093 767
rect 2175 767 2176 771
rect 2183 767 2184 771
rect 2230 771 2231 775
rect 2235 771 2236 775
rect 2318 775 2324 776
rect 2230 770 2236 771
rect 2263 771 2272 772
rect 2175 766 2184 767
rect 2263 767 2264 771
rect 2271 767 2272 771
rect 2318 771 2319 775
rect 2323 771 2324 775
rect 2406 775 2412 776
rect 2318 770 2324 771
rect 2351 771 2357 772
rect 2263 766 2272 767
rect 2351 767 2352 771
rect 2356 770 2357 771
rect 2359 771 2365 772
rect 2359 770 2360 771
rect 2356 768 2360 770
rect 2356 767 2357 768
rect 2351 766 2357 767
rect 2359 767 2360 768
rect 2364 767 2365 771
rect 2406 771 2407 775
rect 2411 771 2412 775
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2406 770 2412 771
rect 2438 771 2445 772
rect 2582 771 2588 772
rect 2359 766 2365 767
rect 2438 767 2439 771
rect 2444 767 2445 771
rect 2438 766 2445 767
rect 158 755 164 756
rect 158 751 159 755
rect 163 754 164 755
rect 163 752 626 754
rect 163 751 164 752
rect 158 750 164 751
rect 175 747 181 748
rect 142 745 148 746
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 142 741 143 745
rect 147 741 148 745
rect 175 743 176 747
rect 180 746 181 747
rect 190 747 196 748
rect 190 746 191 747
rect 180 744 191 746
rect 180 743 181 744
rect 175 742 181 743
rect 190 743 191 744
rect 195 743 196 747
rect 231 747 237 748
rect 190 742 196 743
rect 198 745 204 746
rect 142 740 148 741
rect 198 741 199 745
rect 203 741 204 745
rect 231 743 232 747
rect 236 746 237 747
rect 270 747 276 748
rect 270 746 271 747
rect 236 744 271 746
rect 236 743 237 744
rect 231 742 237 743
rect 270 743 271 744
rect 275 743 276 747
rect 311 747 317 748
rect 270 742 276 743
rect 278 745 284 746
rect 198 740 204 741
rect 278 741 279 745
rect 283 741 284 745
rect 311 743 312 747
rect 316 746 317 747
rect 374 747 380 748
rect 374 746 375 747
rect 316 744 375 746
rect 316 743 317 744
rect 311 742 317 743
rect 374 743 375 744
rect 379 743 380 747
rect 415 747 421 748
rect 374 742 380 743
rect 382 745 388 746
rect 278 740 284 741
rect 382 741 383 745
rect 387 741 388 745
rect 415 743 416 747
rect 420 746 421 747
rect 478 747 484 748
rect 478 746 479 747
rect 420 744 479 746
rect 420 743 421 744
rect 415 742 421 743
rect 478 743 479 744
rect 483 743 484 747
rect 519 747 525 748
rect 478 742 484 743
rect 486 745 492 746
rect 382 740 388 741
rect 486 741 487 745
rect 491 741 492 745
rect 519 743 520 747
rect 524 746 525 747
rect 590 747 596 748
rect 590 746 591 747
rect 524 744 591 746
rect 524 743 525 744
rect 519 742 525 743
rect 590 743 591 744
rect 595 743 596 747
rect 624 746 626 752
rect 631 747 637 748
rect 631 746 632 747
rect 590 742 596 743
rect 598 745 604 746
rect 486 740 492 741
rect 598 741 599 745
rect 603 741 604 745
rect 624 744 632 746
rect 631 743 632 744
rect 636 743 637 747
rect 735 747 741 748
rect 631 742 637 743
rect 702 745 708 746
rect 598 740 604 741
rect 702 741 703 745
rect 707 741 708 745
rect 735 743 736 747
rect 740 746 741 747
rect 798 747 804 748
rect 798 746 799 747
rect 740 744 799 746
rect 740 743 741 744
rect 735 742 741 743
rect 798 743 799 744
rect 803 743 804 747
rect 839 747 845 748
rect 798 742 804 743
rect 806 745 812 746
rect 702 740 708 741
rect 806 741 807 745
rect 811 741 812 745
rect 839 743 840 747
rect 844 746 845 747
rect 894 747 900 748
rect 894 746 895 747
rect 844 744 895 746
rect 844 743 845 744
rect 839 742 845 743
rect 894 743 895 744
rect 899 743 900 747
rect 935 747 941 748
rect 894 742 900 743
rect 902 745 908 746
rect 806 740 812 741
rect 902 741 903 745
rect 907 741 908 745
rect 935 743 936 747
rect 940 746 941 747
rect 982 747 988 748
rect 982 746 983 747
rect 940 744 983 746
rect 940 743 941 744
rect 935 742 941 743
rect 982 743 983 744
rect 987 743 988 747
rect 1023 747 1029 748
rect 982 742 988 743
rect 990 745 996 746
rect 902 740 908 741
rect 990 741 991 745
rect 995 741 996 745
rect 1023 743 1024 747
rect 1028 746 1029 747
rect 1070 747 1076 748
rect 1070 746 1071 747
rect 1028 744 1071 746
rect 1028 743 1029 744
rect 1023 742 1029 743
rect 1070 743 1071 744
rect 1075 743 1076 747
rect 1111 747 1117 748
rect 1070 742 1076 743
rect 1078 745 1084 746
rect 990 740 996 741
rect 1078 741 1079 745
rect 1083 741 1084 745
rect 1111 743 1112 747
rect 1116 746 1117 747
rect 1166 747 1172 748
rect 1166 746 1167 747
rect 1116 744 1167 746
rect 1116 743 1117 744
rect 1111 742 1117 743
rect 1166 743 1167 744
rect 1171 743 1172 747
rect 1198 747 1204 748
rect 1166 742 1172 743
rect 1174 745 1180 746
rect 1078 740 1084 741
rect 1174 741 1175 745
rect 1179 741 1180 745
rect 1198 743 1199 747
rect 1203 746 1204 747
rect 1207 747 1213 748
rect 1207 746 1208 747
rect 1203 744 1208 746
rect 1203 743 1204 744
rect 1198 742 1204 743
rect 1207 743 1208 744
rect 1212 743 1213 747
rect 2150 747 2156 748
rect 1207 742 1213 743
rect 1326 744 1332 745
rect 1174 740 1180 741
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 2054 743 2060 744
rect 110 739 116 740
rect 1326 739 1332 740
rect 1599 739 1605 740
rect 1566 737 1572 738
rect 1366 736 1372 737
rect 1366 732 1367 736
rect 1371 732 1372 736
rect 1566 733 1567 737
rect 1571 733 1572 737
rect 1599 735 1600 739
rect 1604 738 1605 739
rect 1614 739 1620 740
rect 1614 738 1615 739
rect 1604 736 1615 738
rect 1604 735 1605 736
rect 1599 734 1605 735
rect 1614 735 1615 736
rect 1619 735 1620 739
rect 1655 739 1661 740
rect 1614 734 1620 735
rect 1622 737 1628 738
rect 1566 732 1572 733
rect 1622 733 1623 737
rect 1627 733 1628 737
rect 1655 735 1656 739
rect 1660 738 1661 739
rect 1678 739 1684 740
rect 1678 738 1679 739
rect 1660 736 1679 738
rect 1660 735 1661 736
rect 1655 734 1661 735
rect 1678 735 1679 736
rect 1683 735 1684 739
rect 1719 739 1725 740
rect 1678 734 1684 735
rect 1686 737 1692 738
rect 1622 732 1628 733
rect 1686 733 1687 737
rect 1691 733 1692 737
rect 1719 735 1720 739
rect 1724 738 1725 739
rect 1750 739 1756 740
rect 1750 738 1751 739
rect 1724 736 1751 738
rect 1724 735 1725 736
rect 1719 734 1725 735
rect 1750 735 1751 736
rect 1755 735 1756 739
rect 1791 739 1797 740
rect 1750 734 1756 735
rect 1758 737 1764 738
rect 1686 732 1692 733
rect 1758 733 1759 737
rect 1763 733 1764 737
rect 1791 735 1792 739
rect 1796 738 1797 739
rect 1830 739 1836 740
rect 1830 738 1831 739
rect 1796 736 1831 738
rect 1796 735 1797 736
rect 1791 734 1797 735
rect 1830 735 1831 736
rect 1835 735 1836 739
rect 1871 739 1877 740
rect 1830 734 1836 735
rect 1838 737 1844 738
rect 1758 732 1764 733
rect 1838 733 1839 737
rect 1843 733 1844 737
rect 1871 735 1872 739
rect 1876 738 1877 739
rect 1910 739 1916 740
rect 1910 738 1911 739
rect 1876 736 1911 738
rect 1876 735 1877 736
rect 1871 734 1877 735
rect 1910 735 1911 736
rect 1915 735 1916 739
rect 1951 739 1957 740
rect 1910 734 1916 735
rect 1918 737 1924 738
rect 1838 732 1844 733
rect 1918 733 1919 737
rect 1923 733 1924 737
rect 1951 735 1952 739
rect 1956 738 1957 739
rect 1959 739 1965 740
rect 1959 738 1960 739
rect 1956 736 1960 738
rect 1956 735 1957 736
rect 1951 734 1957 735
rect 1959 735 1960 736
rect 1964 735 1965 739
rect 2030 739 2037 740
rect 1959 734 1965 735
rect 1998 737 2004 738
rect 1918 732 1924 733
rect 1998 733 1999 737
rect 2003 733 2004 737
rect 2030 735 2031 739
rect 2036 735 2037 739
rect 2054 739 2055 743
rect 2059 742 2060 743
rect 2150 743 2151 747
rect 2155 746 2156 747
rect 2155 744 2362 746
rect 2155 743 2156 744
rect 2150 742 2156 743
rect 2059 740 2106 742
rect 2059 739 2060 740
rect 2054 738 2060 739
rect 2104 738 2106 740
rect 2111 739 2117 740
rect 2111 738 2112 739
rect 2030 734 2037 735
rect 2078 737 2084 738
rect 1998 732 2004 733
rect 2078 733 2079 737
rect 2083 733 2084 737
rect 2104 736 2112 738
rect 2111 735 2112 736
rect 2116 735 2117 739
rect 2191 739 2197 740
rect 2111 734 2117 735
rect 2158 737 2164 738
rect 2078 732 2084 733
rect 2158 733 2159 737
rect 2163 733 2164 737
rect 2191 735 2192 739
rect 2196 738 2197 739
rect 2238 739 2244 740
rect 2238 738 2239 739
rect 2196 736 2239 738
rect 2196 735 2197 736
rect 2191 734 2197 735
rect 2238 735 2239 736
rect 2243 735 2244 739
rect 2279 739 2285 740
rect 2238 734 2244 735
rect 2246 737 2252 738
rect 2158 732 2164 733
rect 2246 733 2247 737
rect 2251 733 2252 737
rect 2279 735 2280 739
rect 2284 738 2285 739
rect 2326 739 2332 740
rect 2326 738 2327 739
rect 2284 736 2327 738
rect 2284 735 2285 736
rect 2279 734 2285 735
rect 2326 735 2327 736
rect 2331 735 2332 739
rect 2360 738 2362 744
rect 2367 739 2373 740
rect 2367 738 2368 739
rect 2326 734 2332 735
rect 2334 737 2340 738
rect 2246 732 2252 733
rect 2334 733 2335 737
rect 2339 733 2340 737
rect 2360 736 2368 738
rect 2367 735 2368 736
rect 2372 735 2373 739
rect 2367 734 2373 735
rect 2582 736 2588 737
rect 2334 732 2340 733
rect 2582 732 2583 736
rect 2587 732 2588 736
rect 1366 731 1372 732
rect 2582 731 2588 732
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 1326 727 1332 728
rect 1326 723 1327 727
rect 1331 723 1332 727
rect 1326 722 1332 723
rect 1366 719 1372 720
rect 158 718 164 719
rect 158 714 159 718
rect 163 714 164 718
rect 158 713 164 714
rect 214 718 220 719
rect 214 714 215 718
rect 219 714 220 718
rect 214 713 220 714
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 502 718 508 719
rect 502 714 503 718
rect 507 714 508 718
rect 502 713 508 714
rect 614 718 620 719
rect 614 714 615 718
rect 619 714 620 718
rect 614 713 620 714
rect 718 718 724 719
rect 718 714 719 718
rect 723 714 724 718
rect 718 713 724 714
rect 822 718 828 719
rect 822 714 823 718
rect 827 714 828 718
rect 822 713 828 714
rect 918 718 924 719
rect 918 714 919 718
rect 923 714 924 718
rect 918 713 924 714
rect 1006 718 1012 719
rect 1006 714 1007 718
rect 1011 714 1012 718
rect 1006 713 1012 714
rect 1094 718 1100 719
rect 1094 714 1095 718
rect 1099 714 1100 718
rect 1094 713 1100 714
rect 1190 718 1196 719
rect 1190 714 1191 718
rect 1195 714 1196 718
rect 1366 715 1367 719
rect 1371 715 1372 719
rect 1366 714 1372 715
rect 2582 719 2588 720
rect 2582 715 2583 719
rect 2587 715 2588 719
rect 2582 714 2588 715
rect 1190 713 1196 714
rect 135 711 141 712
rect 135 707 136 711
rect 140 710 141 711
rect 190 711 197 712
rect 140 708 186 710
rect 140 707 141 708
rect 135 706 141 707
rect 184 702 186 708
rect 190 707 191 711
rect 196 707 197 711
rect 190 706 197 707
rect 270 711 277 712
rect 270 707 271 711
rect 276 707 277 711
rect 270 706 277 707
rect 374 711 381 712
rect 374 707 375 711
rect 380 707 381 711
rect 374 706 381 707
rect 478 711 485 712
rect 478 707 479 711
rect 484 707 485 711
rect 478 706 485 707
rect 590 711 597 712
rect 590 707 591 711
rect 596 707 597 711
rect 590 706 597 707
rect 695 711 704 712
rect 695 707 696 711
rect 703 707 704 711
rect 695 706 704 707
rect 798 711 805 712
rect 798 707 799 711
rect 804 707 805 711
rect 798 706 805 707
rect 894 711 901 712
rect 894 707 895 711
rect 900 707 901 711
rect 894 706 901 707
rect 982 711 989 712
rect 982 707 983 711
rect 988 707 989 711
rect 982 706 989 707
rect 1070 711 1077 712
rect 1070 707 1071 711
rect 1076 707 1077 711
rect 1070 706 1077 707
rect 1166 711 1173 712
rect 1166 707 1167 711
rect 1172 707 1173 711
rect 1166 706 1173 707
rect 1582 710 1588 711
rect 1582 706 1583 710
rect 1587 706 1588 710
rect 1582 705 1588 706
rect 1638 710 1644 711
rect 1638 706 1639 710
rect 1643 706 1644 710
rect 1638 705 1644 706
rect 1702 710 1708 711
rect 1702 706 1703 710
rect 1707 706 1708 710
rect 1702 705 1708 706
rect 1774 710 1780 711
rect 1774 706 1775 710
rect 1779 706 1780 710
rect 1774 705 1780 706
rect 1854 710 1860 711
rect 1854 706 1855 710
rect 1859 706 1860 710
rect 1854 705 1860 706
rect 1934 710 1940 711
rect 1934 706 1935 710
rect 1939 706 1940 710
rect 1934 705 1940 706
rect 2014 710 2020 711
rect 2014 706 2015 710
rect 2019 706 2020 710
rect 2014 705 2020 706
rect 2094 710 2100 711
rect 2094 706 2095 710
rect 2099 706 2100 710
rect 2094 705 2100 706
rect 2174 710 2180 711
rect 2174 706 2175 710
rect 2179 706 2180 710
rect 2174 705 2180 706
rect 2262 710 2268 711
rect 2262 706 2263 710
rect 2267 706 2268 710
rect 2262 705 2268 706
rect 2350 710 2356 711
rect 2350 706 2351 710
rect 2355 706 2356 710
rect 2350 705 2356 706
rect 366 703 372 704
rect 366 702 367 703
rect 184 700 367 702
rect 366 699 367 700
rect 371 699 372 703
rect 726 703 732 704
rect 726 702 727 703
rect 366 698 372 699
rect 616 700 727 702
rect 134 695 141 696
rect 134 691 135 695
rect 140 691 141 695
rect 178 695 184 696
rect 178 691 179 695
rect 183 694 184 695
rect 191 695 197 696
rect 191 694 192 695
rect 183 692 192 694
rect 183 691 184 692
rect 134 690 141 691
rect 158 690 164 691
rect 178 690 184 691
rect 191 691 192 692
rect 196 691 197 695
rect 242 695 248 696
rect 242 691 243 695
rect 247 694 248 695
rect 255 695 261 696
rect 255 694 256 695
rect 247 692 256 694
rect 247 691 248 692
rect 191 690 197 691
rect 214 690 220 691
rect 242 690 248 691
rect 255 691 256 692
rect 260 691 261 695
rect 303 695 309 696
rect 303 691 304 695
rect 308 694 309 695
rect 335 695 341 696
rect 335 694 336 695
rect 308 692 336 694
rect 308 691 309 692
rect 255 690 261 691
rect 278 690 284 691
rect 303 690 309 691
rect 335 691 336 692
rect 340 691 341 695
rect 374 695 380 696
rect 374 691 375 695
rect 379 694 380 695
rect 423 695 429 696
rect 423 694 424 695
rect 379 692 424 694
rect 379 691 380 692
rect 335 690 341 691
rect 358 690 364 691
rect 374 690 380 691
rect 423 691 424 692
rect 428 691 429 695
rect 466 695 472 696
rect 466 691 467 695
rect 471 694 472 695
rect 511 695 517 696
rect 511 694 512 695
rect 471 692 512 694
rect 471 691 472 692
rect 423 690 429 691
rect 446 690 452 691
rect 466 690 472 691
rect 511 691 512 692
rect 516 691 517 695
rect 599 695 605 696
rect 599 691 600 695
rect 604 694 605 695
rect 616 694 618 700
rect 726 699 727 700
rect 731 699 732 703
rect 886 703 892 704
rect 886 702 887 703
rect 726 698 732 699
rect 785 700 887 702
rect 604 692 618 694
rect 686 695 693 696
rect 604 691 605 692
rect 686 691 687 695
rect 692 691 693 695
rect 767 695 773 696
rect 767 691 768 695
rect 772 694 773 695
rect 785 694 787 700
rect 886 699 887 700
rect 891 699 892 703
rect 1559 703 1565 704
rect 886 698 892 699
rect 1198 699 1204 700
rect 1198 698 1199 699
rect 1033 696 1199 698
rect 772 692 787 694
rect 846 695 853 696
rect 772 691 773 692
rect 846 691 847 695
rect 852 691 853 695
rect 927 695 933 696
rect 927 691 928 695
rect 932 694 933 695
rect 942 695 948 696
rect 942 694 943 695
rect 932 692 943 694
rect 932 691 933 692
rect 511 690 517 691
rect 534 690 540 691
rect 599 690 605 691
rect 622 690 628 691
rect 686 690 693 691
rect 710 690 716 691
rect 767 690 773 691
rect 790 690 796 691
rect 846 690 853 691
rect 870 690 876 691
rect 927 690 933 691
rect 942 691 943 692
rect 947 691 948 695
rect 1015 695 1021 696
rect 1015 691 1016 695
rect 1020 694 1021 695
rect 1033 694 1035 696
rect 1198 695 1199 696
rect 1203 695 1204 699
rect 1559 699 1560 703
rect 1564 702 1565 703
rect 1614 703 1621 704
rect 1564 700 1610 702
rect 1564 699 1565 700
rect 1559 698 1565 699
rect 1198 694 1204 695
rect 1608 694 1610 700
rect 1614 699 1615 703
rect 1620 699 1621 703
rect 1614 698 1621 699
rect 1678 703 1685 704
rect 1678 699 1679 703
rect 1684 699 1685 703
rect 1678 698 1685 699
rect 1750 703 1757 704
rect 1750 699 1751 703
rect 1756 699 1757 703
rect 1750 698 1757 699
rect 1830 703 1837 704
rect 1830 699 1831 703
rect 1836 699 1837 703
rect 1830 698 1837 699
rect 1910 703 1917 704
rect 1910 699 1911 703
rect 1916 699 1917 703
rect 1910 698 1917 699
rect 1991 703 1997 704
rect 1991 699 1992 703
rect 1996 702 1997 703
rect 2054 703 2060 704
rect 2054 702 2055 703
rect 1996 700 2055 702
rect 1996 699 1997 700
rect 1991 698 1997 699
rect 2054 699 2055 700
rect 2059 699 2060 703
rect 2054 698 2060 699
rect 2071 703 2077 704
rect 2071 699 2072 703
rect 2076 702 2077 703
rect 2086 703 2092 704
rect 2086 702 2087 703
rect 2076 700 2087 702
rect 2076 699 2077 700
rect 2071 698 2077 699
rect 2086 699 2087 700
rect 2091 699 2092 703
rect 2086 698 2092 699
rect 2138 703 2144 704
rect 2138 699 2139 703
rect 2143 702 2144 703
rect 2151 703 2157 704
rect 2151 702 2152 703
rect 2143 700 2152 702
rect 2143 699 2144 700
rect 2138 698 2144 699
rect 2151 699 2152 700
rect 2156 699 2157 703
rect 2151 698 2157 699
rect 2238 703 2245 704
rect 2238 699 2239 703
rect 2244 699 2245 703
rect 2238 698 2245 699
rect 2326 703 2333 704
rect 2326 699 2327 703
rect 2332 699 2333 703
rect 2326 698 2333 699
rect 1838 695 1844 696
rect 1838 694 1839 695
rect 1020 692 1035 694
rect 1608 692 1839 694
rect 1020 691 1021 692
rect 1838 691 1839 692
rect 1843 691 1844 695
rect 2030 695 2036 696
rect 2030 694 2031 695
rect 942 690 948 691
rect 950 690 956 691
rect 1015 690 1021 691
rect 1038 690 1044 691
rect 1838 690 1844 691
rect 1905 692 2031 694
rect 158 686 159 690
rect 163 686 164 690
rect 158 685 164 686
rect 214 686 215 690
rect 219 686 220 690
rect 214 685 220 686
rect 278 686 279 690
rect 283 686 284 690
rect 278 685 284 686
rect 358 686 359 690
rect 363 686 364 690
rect 358 685 364 686
rect 446 686 447 690
rect 451 686 452 690
rect 446 685 452 686
rect 534 686 535 690
rect 539 686 540 690
rect 534 685 540 686
rect 622 686 623 690
rect 627 686 628 690
rect 622 685 628 686
rect 710 686 711 690
rect 715 686 716 690
rect 710 685 716 686
rect 790 686 791 690
rect 795 686 796 690
rect 790 685 796 686
rect 870 686 871 690
rect 875 686 876 690
rect 870 685 876 686
rect 950 686 951 690
rect 955 686 956 690
rect 950 685 956 686
rect 1038 686 1039 690
rect 1043 686 1044 690
rect 1905 688 1907 692
rect 2030 691 2031 692
rect 2035 691 2036 695
rect 2222 695 2228 696
rect 2222 694 2223 695
rect 2030 690 2036 691
rect 2112 692 2223 694
rect 1038 685 1044 686
rect 1391 687 1397 688
rect 1391 683 1392 687
rect 1396 686 1397 687
rect 1406 687 1412 688
rect 1406 686 1407 687
rect 1396 684 1407 686
rect 1396 683 1397 684
rect 1391 682 1397 683
rect 1406 683 1407 684
rect 1411 683 1412 687
rect 1434 687 1440 688
rect 1434 683 1435 687
rect 1439 686 1440 687
rect 1487 687 1493 688
rect 1487 686 1488 687
rect 1439 684 1488 686
rect 1439 683 1440 684
rect 1406 682 1412 683
rect 1414 682 1420 683
rect 1434 682 1440 683
rect 1487 683 1488 684
rect 1492 683 1493 687
rect 1535 687 1541 688
rect 1535 683 1536 687
rect 1540 686 1541 687
rect 1591 687 1597 688
rect 1591 686 1592 687
rect 1540 684 1592 686
rect 1540 683 1541 684
rect 1487 682 1493 683
rect 1510 682 1516 683
rect 1535 682 1541 683
rect 1591 683 1592 684
rect 1596 683 1597 687
rect 1639 687 1645 688
rect 1639 683 1640 687
rect 1644 686 1645 687
rect 1695 687 1701 688
rect 1695 686 1696 687
rect 1644 684 1696 686
rect 1644 683 1645 684
rect 1591 682 1597 683
rect 1614 682 1620 683
rect 1639 682 1645 683
rect 1695 683 1696 684
rect 1700 683 1701 687
rect 1738 687 1744 688
rect 1738 683 1739 687
rect 1743 686 1744 687
rect 1799 687 1805 688
rect 1799 686 1800 687
rect 1743 684 1800 686
rect 1743 683 1744 684
rect 1695 682 1701 683
rect 1718 682 1724 683
rect 1738 682 1744 683
rect 1799 683 1800 684
rect 1804 683 1805 687
rect 1903 687 1909 688
rect 1903 683 1904 687
rect 1908 683 1909 687
rect 1946 687 1952 688
rect 1946 683 1947 687
rect 1951 686 1952 687
rect 1999 687 2005 688
rect 1999 686 2000 687
rect 1951 684 2000 686
rect 1951 683 1952 684
rect 1799 682 1805 683
rect 1822 682 1828 683
rect 1903 682 1909 683
rect 1926 682 1932 683
rect 1946 682 1952 683
rect 1999 683 2000 684
rect 2004 683 2005 687
rect 2095 687 2101 688
rect 2095 683 2096 687
rect 2100 686 2101 687
rect 2112 686 2114 692
rect 2222 691 2223 692
rect 2227 691 2228 695
rect 2222 690 2228 691
rect 2438 691 2444 692
rect 2438 690 2439 691
rect 2384 688 2439 690
rect 2100 684 2114 686
rect 2182 687 2189 688
rect 2100 683 2101 684
rect 2182 683 2183 687
rect 2188 683 2189 687
rect 2271 687 2277 688
rect 2271 683 2272 687
rect 2276 686 2277 687
rect 2286 687 2292 688
rect 2286 686 2287 687
rect 2276 684 2287 686
rect 2276 683 2277 684
rect 1999 682 2005 683
rect 2022 682 2028 683
rect 2095 682 2101 683
rect 2118 682 2124 683
rect 2182 682 2189 683
rect 2206 682 2212 683
rect 2271 682 2277 683
rect 2286 683 2287 684
rect 2291 683 2292 687
rect 2367 687 2373 688
rect 2367 683 2368 687
rect 2372 686 2373 687
rect 2384 686 2386 688
rect 2438 687 2439 688
rect 2443 687 2444 691
rect 2438 686 2444 687
rect 2372 684 2386 686
rect 2372 683 2373 684
rect 2286 682 2292 683
rect 2294 682 2300 683
rect 2367 682 2373 683
rect 2390 682 2396 683
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 1326 681 1332 682
rect 1326 677 1327 681
rect 1331 677 1332 681
rect 1414 678 1415 682
rect 1419 678 1420 682
rect 1414 677 1420 678
rect 1510 678 1511 682
rect 1515 678 1516 682
rect 1510 677 1516 678
rect 1614 678 1615 682
rect 1619 678 1620 682
rect 1614 677 1620 678
rect 1718 678 1719 682
rect 1723 678 1724 682
rect 1718 677 1724 678
rect 1822 678 1823 682
rect 1827 678 1828 682
rect 1822 677 1828 678
rect 1926 678 1927 682
rect 1931 678 1932 682
rect 1926 677 1932 678
rect 2022 678 2023 682
rect 2027 678 2028 682
rect 2022 677 2028 678
rect 2118 678 2119 682
rect 2123 678 2124 682
rect 2118 677 2124 678
rect 2206 678 2207 682
rect 2211 678 2212 682
rect 2206 677 2212 678
rect 2294 678 2295 682
rect 2299 678 2300 682
rect 2294 677 2300 678
rect 2390 678 2391 682
rect 2395 678 2396 682
rect 2390 677 2396 678
rect 1326 676 1332 677
rect 380 672 430 674
rect 1366 673 1372 674
rect 134 671 140 672
rect 134 667 135 671
rect 139 670 140 671
rect 380 670 382 672
rect 139 668 382 670
rect 428 670 430 672
rect 686 671 692 672
rect 428 668 546 670
rect 139 667 140 668
rect 134 666 140 667
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 142 663 148 664
rect 142 659 143 663
rect 147 659 148 663
rect 198 663 204 664
rect 142 658 148 659
rect 175 659 184 660
rect 175 655 176 659
rect 183 655 184 659
rect 198 659 199 663
rect 203 659 204 663
rect 262 663 268 664
rect 198 658 204 659
rect 231 659 237 660
rect 175 654 184 655
rect 231 655 232 659
rect 236 658 237 659
rect 242 659 248 660
rect 242 658 243 659
rect 236 656 243 658
rect 236 655 237 656
rect 231 654 237 655
rect 242 655 243 656
rect 247 655 248 659
rect 262 659 263 663
rect 267 659 268 663
rect 303 663 309 664
rect 303 662 304 663
rect 262 658 268 659
rect 295 661 304 662
rect 295 657 296 661
rect 300 660 304 661
rect 300 657 301 660
rect 303 659 304 660
rect 308 659 309 663
rect 303 658 309 659
rect 342 663 348 664
rect 342 659 343 663
rect 347 659 348 663
rect 430 663 436 664
rect 342 658 348 659
rect 366 659 372 660
rect 295 656 301 657
rect 242 654 248 655
rect 366 655 367 659
rect 371 658 372 659
rect 375 659 381 660
rect 375 658 376 659
rect 371 656 376 658
rect 371 655 372 656
rect 366 654 372 655
rect 375 655 376 656
rect 380 655 381 659
rect 430 659 431 663
rect 435 659 436 663
rect 518 663 524 664
rect 430 658 436 659
rect 463 659 472 660
rect 375 654 381 655
rect 463 655 464 659
rect 471 655 472 659
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 544 658 546 668
rect 686 667 687 671
rect 691 670 692 671
rect 846 671 852 672
rect 691 668 802 670
rect 691 667 692 668
rect 686 666 692 667
rect 606 663 612 664
rect 551 659 557 660
rect 551 658 552 659
rect 544 656 552 658
rect 463 654 472 655
rect 551 655 552 656
rect 556 655 557 659
rect 606 659 607 663
rect 611 659 612 663
rect 694 663 700 664
rect 606 658 612 659
rect 630 659 636 660
rect 551 654 557 655
rect 630 655 631 659
rect 635 658 636 659
rect 639 659 645 660
rect 639 658 640 659
rect 635 656 640 658
rect 635 655 636 656
rect 630 654 636 655
rect 639 655 640 656
rect 644 655 645 659
rect 694 659 695 663
rect 699 659 700 663
rect 774 663 780 664
rect 694 658 700 659
rect 726 659 733 660
rect 639 654 645 655
rect 726 655 727 659
rect 732 655 733 659
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 800 658 802 668
rect 846 667 847 671
rect 851 670 852 671
rect 851 668 962 670
rect 1366 669 1367 673
rect 1371 669 1372 673
rect 1366 668 1372 669
rect 2582 673 2588 674
rect 2582 669 2583 673
rect 2587 669 2588 673
rect 2582 668 2588 669
rect 851 667 852 668
rect 846 666 852 667
rect 854 663 860 664
rect 807 659 813 660
rect 807 658 808 659
rect 800 656 808 658
rect 726 654 733 655
rect 807 655 808 656
rect 812 655 813 659
rect 854 659 855 663
rect 859 659 860 663
rect 934 663 940 664
rect 854 658 860 659
rect 886 659 893 660
rect 807 654 813 655
rect 886 655 887 659
rect 892 655 893 659
rect 934 659 935 663
rect 939 659 940 663
rect 934 658 940 659
rect 960 658 962 668
rect 1326 664 1332 665
rect 1022 663 1028 664
rect 967 659 973 660
rect 967 658 968 659
rect 960 656 968 658
rect 886 654 893 655
rect 967 655 968 656
rect 972 655 973 659
rect 1022 659 1023 663
rect 1027 659 1028 663
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1022 658 1028 659
rect 1055 659 1061 660
rect 1326 659 1332 660
rect 2182 663 2188 664
rect 2182 659 2183 663
rect 2187 662 2188 663
rect 2187 660 2306 662
rect 2187 659 2188 660
rect 1055 658 1056 659
rect 967 654 973 655
rect 1032 656 1056 658
rect 942 651 948 652
rect 942 647 943 651
rect 947 650 948 651
rect 1032 650 1034 656
rect 1055 655 1056 656
rect 1060 655 1061 659
rect 2182 658 2188 659
rect 1055 654 1061 655
rect 1366 656 1372 657
rect 1366 652 1367 656
rect 1371 652 1372 656
rect 1366 651 1372 652
rect 1398 655 1404 656
rect 1398 651 1399 655
rect 1403 651 1404 655
rect 1494 655 1500 656
rect 1398 650 1404 651
rect 1431 651 1440 652
rect 947 648 1034 650
rect 947 647 948 648
rect 942 646 948 647
rect 1431 647 1432 651
rect 1439 647 1440 651
rect 1494 651 1495 655
rect 1499 651 1500 655
rect 1598 655 1604 656
rect 1494 650 1500 651
rect 1527 651 1533 652
rect 1431 646 1440 647
rect 1527 647 1528 651
rect 1532 650 1533 651
rect 1535 651 1541 652
rect 1535 650 1536 651
rect 1532 648 1536 650
rect 1532 647 1533 648
rect 1527 646 1533 647
rect 1535 647 1536 648
rect 1540 647 1541 651
rect 1598 651 1599 655
rect 1603 651 1604 655
rect 1702 655 1708 656
rect 1598 650 1604 651
rect 1631 651 1637 652
rect 1535 646 1541 647
rect 1631 647 1632 651
rect 1636 650 1637 651
rect 1639 651 1645 652
rect 1639 650 1640 651
rect 1636 648 1640 650
rect 1636 647 1637 648
rect 1631 646 1637 647
rect 1639 647 1640 648
rect 1644 647 1645 651
rect 1702 651 1703 655
rect 1707 651 1708 655
rect 1806 655 1812 656
rect 1702 650 1708 651
rect 1735 651 1744 652
rect 1639 646 1645 647
rect 1735 647 1736 651
rect 1743 647 1744 651
rect 1806 651 1807 655
rect 1811 651 1812 655
rect 1910 655 1916 656
rect 1806 650 1812 651
rect 1838 651 1845 652
rect 1735 646 1744 647
rect 1838 647 1839 651
rect 1844 647 1845 651
rect 1910 651 1911 655
rect 1915 651 1916 655
rect 2006 655 2012 656
rect 1910 650 1916 651
rect 1943 651 1952 652
rect 1838 646 1845 647
rect 1943 647 1944 651
rect 1951 647 1952 651
rect 2006 651 2007 655
rect 2011 651 2012 655
rect 2102 655 2108 656
rect 2006 650 2012 651
rect 2030 651 2036 652
rect 1943 646 1952 647
rect 2030 647 2031 651
rect 2035 650 2036 651
rect 2039 651 2045 652
rect 2039 650 2040 651
rect 2035 648 2040 650
rect 2035 647 2036 648
rect 2030 646 2036 647
rect 2039 647 2040 648
rect 2044 647 2045 651
rect 2102 651 2103 655
rect 2107 651 2108 655
rect 2190 655 2196 656
rect 2102 650 2108 651
rect 2135 651 2144 652
rect 2039 646 2045 647
rect 2135 647 2136 651
rect 2143 647 2144 651
rect 2190 651 2191 655
rect 2195 651 2196 655
rect 2278 655 2284 656
rect 2190 650 2196 651
rect 2222 651 2229 652
rect 2135 646 2144 647
rect 2222 647 2223 651
rect 2228 647 2229 651
rect 2278 651 2279 655
rect 2283 651 2284 655
rect 2278 650 2284 651
rect 2304 650 2306 660
rect 2582 656 2588 657
rect 2374 655 2380 656
rect 2311 651 2317 652
rect 2311 650 2312 651
rect 2304 648 2312 650
rect 2222 646 2229 647
rect 2311 647 2312 648
rect 2316 647 2317 651
rect 2374 651 2375 655
rect 2379 651 2380 655
rect 2582 652 2583 656
rect 2587 652 2588 656
rect 2374 650 2380 651
rect 2407 651 2413 652
rect 2582 651 2588 652
rect 2311 646 2317 647
rect 2407 647 2408 651
rect 2412 647 2413 651
rect 2407 646 2413 647
rect 2286 643 2292 644
rect 374 639 380 640
rect 374 638 375 639
rect 319 636 375 638
rect 319 626 321 636
rect 374 635 375 636
rect 379 635 380 639
rect 2286 639 2287 643
rect 2291 642 2292 643
rect 2409 642 2411 646
rect 2291 640 2411 642
rect 2291 639 2292 640
rect 2286 638 2292 639
rect 374 634 380 635
rect 1638 635 1644 636
rect 1638 634 1639 635
rect 1320 632 1639 634
rect 334 631 340 632
rect 334 627 335 631
rect 339 630 340 631
rect 339 628 506 630
rect 339 627 340 628
rect 334 626 340 627
rect 304 624 321 626
rect 175 623 181 624
rect 142 621 148 622
rect 110 620 116 621
rect 110 616 111 620
rect 115 616 116 620
rect 142 617 143 621
rect 147 617 148 621
rect 175 619 176 623
rect 180 622 181 623
rect 190 623 196 624
rect 190 622 191 623
rect 180 620 191 622
rect 180 619 181 620
rect 175 618 181 619
rect 190 619 191 620
rect 195 619 196 623
rect 231 623 237 624
rect 190 618 196 619
rect 198 621 204 622
rect 142 616 148 617
rect 198 617 199 621
rect 203 617 204 621
rect 231 619 232 623
rect 236 622 237 623
rect 246 623 252 624
rect 246 622 247 623
rect 236 620 247 622
rect 236 619 237 620
rect 231 618 237 619
rect 246 619 247 620
rect 251 619 252 623
rect 287 623 293 624
rect 246 618 252 619
rect 254 621 260 622
rect 198 616 204 617
rect 254 617 255 621
rect 259 617 260 621
rect 287 619 288 623
rect 292 622 293 623
rect 304 622 306 624
rect 342 623 349 624
rect 292 620 306 622
rect 310 621 316 622
rect 292 619 293 620
rect 287 618 293 619
rect 254 616 260 617
rect 310 617 311 621
rect 315 617 316 621
rect 342 619 343 623
rect 348 619 349 623
rect 423 623 429 624
rect 342 618 349 619
rect 390 621 396 622
rect 310 616 316 617
rect 390 617 391 621
rect 395 617 396 621
rect 423 619 424 623
rect 428 622 429 623
rect 470 623 476 624
rect 470 622 471 623
rect 428 620 471 622
rect 428 619 429 620
rect 423 618 429 619
rect 470 619 471 620
rect 475 619 476 623
rect 504 622 506 628
rect 511 623 517 624
rect 511 622 512 623
rect 470 618 476 619
rect 478 621 484 622
rect 390 616 396 617
rect 478 617 479 621
rect 483 617 484 621
rect 504 620 512 622
rect 511 619 512 620
rect 516 619 517 623
rect 607 623 613 624
rect 511 618 517 619
rect 574 621 580 622
rect 478 616 484 617
rect 574 617 575 621
rect 579 617 580 621
rect 607 619 608 623
rect 612 622 613 623
rect 670 623 676 624
rect 670 622 671 623
rect 612 620 671 622
rect 612 619 613 620
rect 607 618 613 619
rect 670 619 671 620
rect 675 619 676 623
rect 711 623 717 624
rect 670 618 676 619
rect 678 621 684 622
rect 574 616 580 617
rect 678 617 679 621
rect 683 617 684 621
rect 711 619 712 623
rect 716 622 717 623
rect 774 623 780 624
rect 774 622 775 623
rect 716 620 775 622
rect 716 619 717 620
rect 711 618 717 619
rect 774 619 775 620
rect 779 619 780 623
rect 815 623 821 624
rect 774 618 780 619
rect 782 621 788 622
rect 678 616 684 617
rect 782 617 783 621
rect 787 617 788 621
rect 815 619 816 623
rect 820 622 821 623
rect 878 623 884 624
rect 878 622 879 623
rect 820 620 879 622
rect 820 619 821 620
rect 815 618 821 619
rect 878 619 879 620
rect 883 619 884 623
rect 918 623 925 624
rect 878 618 884 619
rect 886 621 892 622
rect 782 616 788 617
rect 886 617 887 621
rect 891 617 892 621
rect 918 619 919 623
rect 924 619 925 623
rect 1023 623 1029 624
rect 918 618 925 619
rect 990 621 996 622
rect 886 616 892 617
rect 990 617 991 621
rect 995 617 996 621
rect 1023 619 1024 623
rect 1028 622 1029 623
rect 1078 623 1084 624
rect 1078 622 1079 623
rect 1028 620 1079 622
rect 1028 619 1029 620
rect 1023 618 1029 619
rect 1078 619 1079 620
rect 1083 619 1084 623
rect 1119 623 1125 624
rect 1078 618 1084 619
rect 1086 621 1092 622
rect 990 616 996 617
rect 1086 617 1087 621
rect 1091 617 1092 621
rect 1119 619 1120 623
rect 1124 622 1125 623
rect 1182 623 1188 624
rect 1182 622 1183 623
rect 1124 620 1183 622
rect 1124 619 1125 620
rect 1119 618 1125 619
rect 1182 619 1183 620
rect 1187 619 1188 623
rect 1223 623 1229 624
rect 1182 618 1188 619
rect 1190 621 1196 622
rect 1086 616 1092 617
rect 1190 617 1191 621
rect 1195 617 1196 621
rect 1223 619 1224 623
rect 1228 622 1229 623
rect 1262 623 1268 624
rect 1262 622 1263 623
rect 1228 620 1263 622
rect 1228 619 1229 620
rect 1223 618 1229 619
rect 1262 619 1263 620
rect 1267 619 1268 623
rect 1303 623 1309 624
rect 1262 618 1268 619
rect 1270 621 1276 622
rect 1190 616 1196 617
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1303 619 1304 623
rect 1308 622 1309 623
rect 1320 622 1322 632
rect 1638 631 1639 632
rect 1643 631 1644 635
rect 1638 630 1644 631
rect 1439 627 1445 628
rect 1422 623 1428 624
rect 1308 620 1322 622
rect 1398 621 1404 622
rect 1326 620 1332 621
rect 1308 619 1309 620
rect 1303 618 1309 619
rect 1270 616 1276 617
rect 1326 616 1327 620
rect 1331 616 1332 620
rect 110 615 116 616
rect 1326 615 1332 616
rect 1366 620 1372 621
rect 1366 616 1367 620
rect 1371 616 1372 620
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1422 619 1423 623
rect 1427 622 1428 623
rect 1431 623 1437 624
rect 1431 622 1432 623
rect 1427 620 1432 622
rect 1427 619 1428 620
rect 1422 618 1428 619
rect 1431 619 1432 620
rect 1436 619 1437 623
rect 1439 623 1440 627
rect 1444 626 1445 627
rect 1951 627 1957 628
rect 1444 624 1538 626
rect 1444 623 1445 624
rect 1439 622 1445 623
rect 1536 622 1538 624
rect 1543 623 1549 624
rect 1543 622 1544 623
rect 1431 618 1437 619
rect 1510 621 1516 622
rect 1398 616 1404 617
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1536 620 1544 622
rect 1543 619 1544 620
rect 1548 619 1549 623
rect 1679 623 1685 624
rect 1543 618 1549 619
rect 1646 621 1652 622
rect 1510 616 1516 617
rect 1646 617 1647 621
rect 1651 617 1652 621
rect 1679 619 1680 623
rect 1684 622 1685 623
rect 1774 623 1780 624
rect 1774 622 1775 623
rect 1684 620 1775 622
rect 1684 619 1685 620
rect 1679 618 1685 619
rect 1774 619 1775 620
rect 1779 619 1780 623
rect 1814 623 1821 624
rect 1774 618 1780 619
rect 1782 621 1788 622
rect 1646 616 1652 617
rect 1782 617 1783 621
rect 1787 617 1788 621
rect 1814 619 1815 623
rect 1820 619 1821 623
rect 1938 623 1949 624
rect 1814 618 1821 619
rect 1910 621 1916 622
rect 1782 616 1788 617
rect 1910 617 1911 621
rect 1915 617 1916 621
rect 1938 619 1939 623
rect 1943 619 1944 623
rect 1948 619 1949 623
rect 1951 623 1952 627
rect 1956 626 1957 627
rect 1956 624 2075 626
rect 1956 623 1957 624
rect 1951 622 1957 623
rect 2071 623 2077 624
rect 1938 618 1949 619
rect 2038 621 2044 622
rect 1910 616 1916 617
rect 2038 617 2039 621
rect 2043 617 2044 621
rect 2071 619 2072 623
rect 2076 619 2077 623
rect 2191 623 2197 624
rect 2071 618 2077 619
rect 2158 621 2164 622
rect 2038 616 2044 617
rect 2158 617 2159 621
rect 2163 617 2164 621
rect 2191 619 2192 623
rect 2196 622 2197 623
rect 2270 623 2276 624
rect 2270 622 2271 623
rect 2196 620 2271 622
rect 2196 619 2197 620
rect 2191 618 2197 619
rect 2270 619 2271 620
rect 2275 619 2276 623
rect 2311 623 2317 624
rect 2270 618 2276 619
rect 2278 621 2284 622
rect 2158 616 2164 617
rect 2278 617 2279 621
rect 2283 617 2284 621
rect 2311 619 2312 623
rect 2316 622 2317 623
rect 2398 623 2404 624
rect 2398 622 2399 623
rect 2316 620 2399 622
rect 2316 619 2317 620
rect 2311 618 2317 619
rect 2398 619 2399 620
rect 2403 619 2404 623
rect 2438 623 2445 624
rect 2398 618 2404 619
rect 2406 621 2412 622
rect 2278 616 2284 617
rect 2406 617 2407 621
rect 2411 617 2412 621
rect 2438 619 2439 623
rect 2444 619 2445 623
rect 2438 618 2445 619
rect 2582 620 2588 621
rect 2406 616 2412 617
rect 2582 616 2583 620
rect 2587 616 2588 620
rect 1366 615 1372 616
rect 2582 615 2588 616
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 1326 603 1332 604
rect 1326 599 1327 603
rect 1331 599 1332 603
rect 1326 598 1332 599
rect 1366 603 1372 604
rect 1366 599 1367 603
rect 1371 599 1372 603
rect 1366 598 1372 599
rect 2582 603 2588 604
rect 2582 599 2583 603
rect 2587 599 2588 603
rect 2582 598 2588 599
rect 158 594 164 595
rect 158 590 159 594
rect 163 590 164 594
rect 158 589 164 590
rect 214 594 220 595
rect 214 590 215 594
rect 219 590 220 594
rect 214 589 220 590
rect 270 594 276 595
rect 270 590 271 594
rect 275 590 276 594
rect 270 589 276 590
rect 326 594 332 595
rect 326 590 327 594
rect 331 590 332 594
rect 326 589 332 590
rect 406 594 412 595
rect 406 590 407 594
rect 411 590 412 594
rect 406 589 412 590
rect 494 594 500 595
rect 494 590 495 594
rect 499 590 500 594
rect 494 589 500 590
rect 590 594 596 595
rect 590 590 591 594
rect 595 590 596 594
rect 590 589 596 590
rect 694 594 700 595
rect 694 590 695 594
rect 699 590 700 594
rect 694 589 700 590
rect 798 594 804 595
rect 798 590 799 594
rect 803 590 804 594
rect 798 589 804 590
rect 902 594 908 595
rect 902 590 903 594
rect 907 590 908 594
rect 902 589 908 590
rect 1006 594 1012 595
rect 1006 590 1007 594
rect 1011 590 1012 594
rect 1006 589 1012 590
rect 1102 594 1108 595
rect 1102 590 1103 594
rect 1107 590 1108 594
rect 1102 589 1108 590
rect 1206 594 1212 595
rect 1206 590 1207 594
rect 1211 590 1212 594
rect 1206 589 1212 590
rect 1286 594 1292 595
rect 1286 590 1287 594
rect 1291 590 1292 594
rect 1286 589 1292 590
rect 1414 594 1420 595
rect 1414 590 1415 594
rect 1419 590 1420 594
rect 1414 589 1420 590
rect 1526 594 1532 595
rect 1526 590 1527 594
rect 1531 590 1532 594
rect 1526 589 1532 590
rect 1662 594 1668 595
rect 1662 590 1663 594
rect 1667 590 1668 594
rect 1662 589 1668 590
rect 1798 594 1804 595
rect 1798 590 1799 594
rect 1803 590 1804 594
rect 1798 589 1804 590
rect 1926 594 1932 595
rect 1926 590 1927 594
rect 1931 590 1932 594
rect 1926 589 1932 590
rect 2054 594 2060 595
rect 2054 590 2055 594
rect 2059 590 2060 594
rect 2054 589 2060 590
rect 2174 594 2180 595
rect 2174 590 2175 594
rect 2179 590 2180 594
rect 2174 589 2180 590
rect 2294 594 2300 595
rect 2294 590 2295 594
rect 2299 590 2300 594
rect 2294 589 2300 590
rect 2422 594 2428 595
rect 2422 590 2423 594
rect 2427 590 2428 594
rect 2422 589 2428 590
rect 135 587 141 588
rect 135 583 136 587
rect 140 586 141 587
rect 190 587 197 588
rect 140 584 186 586
rect 140 583 141 584
rect 135 582 141 583
rect 184 578 186 584
rect 190 583 191 587
rect 196 583 197 587
rect 190 582 197 583
rect 246 587 253 588
rect 246 583 247 587
rect 252 583 253 587
rect 246 582 253 583
rect 303 587 309 588
rect 303 583 304 587
rect 308 586 309 587
rect 334 587 340 588
rect 334 586 335 587
rect 308 584 335 586
rect 308 583 309 584
rect 303 582 309 583
rect 334 583 335 584
rect 339 583 340 587
rect 334 582 340 583
rect 354 587 360 588
rect 354 583 355 587
rect 359 586 360 587
rect 383 587 389 588
rect 383 586 384 587
rect 359 584 384 586
rect 359 583 360 584
rect 354 582 360 583
rect 383 583 384 584
rect 388 583 389 587
rect 383 582 389 583
rect 470 587 477 588
rect 470 583 471 587
rect 476 583 477 587
rect 470 582 477 583
rect 567 587 573 588
rect 567 583 568 587
rect 572 586 573 587
rect 630 587 636 588
rect 630 586 631 587
rect 572 584 631 586
rect 572 583 573 584
rect 567 582 573 583
rect 630 583 631 584
rect 635 583 636 587
rect 630 582 636 583
rect 670 587 677 588
rect 670 583 671 587
rect 676 583 677 587
rect 670 582 677 583
rect 774 587 781 588
rect 774 583 775 587
rect 780 583 781 587
rect 774 582 781 583
rect 878 587 885 588
rect 878 583 879 587
rect 884 583 885 587
rect 878 582 885 583
rect 983 587 989 588
rect 983 583 984 587
rect 988 586 989 587
rect 1070 587 1076 588
rect 1070 586 1071 587
rect 988 584 1071 586
rect 988 583 989 584
rect 983 582 989 583
rect 1070 583 1071 584
rect 1075 583 1076 587
rect 1070 582 1076 583
rect 1078 587 1085 588
rect 1078 583 1079 587
rect 1084 583 1085 587
rect 1078 582 1085 583
rect 1182 587 1189 588
rect 1182 583 1183 587
rect 1188 583 1189 587
rect 1182 582 1189 583
rect 1262 587 1269 588
rect 1262 583 1263 587
rect 1268 583 1269 587
rect 1262 582 1269 583
rect 1391 587 1397 588
rect 1391 583 1392 587
rect 1396 586 1397 587
rect 1439 587 1445 588
rect 1439 586 1440 587
rect 1396 584 1440 586
rect 1396 583 1397 584
rect 1391 582 1397 583
rect 1439 583 1440 584
rect 1444 583 1445 587
rect 1439 582 1445 583
rect 1490 587 1496 588
rect 1490 583 1491 587
rect 1495 586 1496 587
rect 1503 587 1509 588
rect 1503 586 1504 587
rect 1495 584 1504 586
rect 1495 583 1496 584
rect 1490 582 1496 583
rect 1503 583 1504 584
rect 1508 583 1509 587
rect 1503 582 1509 583
rect 1638 587 1645 588
rect 1638 583 1639 587
rect 1644 583 1645 587
rect 1638 582 1645 583
rect 1774 587 1781 588
rect 1774 583 1775 587
rect 1780 583 1781 587
rect 1774 582 1781 583
rect 1903 587 1909 588
rect 1903 583 1904 587
rect 1908 586 1909 587
rect 1951 587 1957 588
rect 1951 586 1952 587
rect 1908 584 1952 586
rect 1908 583 1909 584
rect 1903 582 1909 583
rect 1951 583 1952 584
rect 1956 583 1957 587
rect 1951 582 1957 583
rect 2030 587 2037 588
rect 2030 583 2031 587
rect 2036 583 2037 587
rect 2030 582 2037 583
rect 2151 587 2157 588
rect 2151 583 2152 587
rect 2156 586 2157 587
rect 2254 587 2260 588
rect 2254 586 2255 587
rect 2156 584 2255 586
rect 2156 583 2157 584
rect 2151 582 2157 583
rect 2254 583 2255 584
rect 2259 583 2260 587
rect 2254 582 2260 583
rect 2270 587 2277 588
rect 2270 583 2271 587
rect 2276 583 2277 587
rect 2270 582 2277 583
rect 2398 587 2405 588
rect 2398 583 2399 587
rect 2404 583 2405 587
rect 2398 582 2405 583
rect 342 579 348 580
rect 342 578 343 579
rect 184 576 343 578
rect 342 575 343 576
rect 347 575 348 579
rect 846 579 852 580
rect 846 578 847 579
rect 342 574 348 575
rect 713 576 847 578
rect 175 571 181 572
rect 175 567 176 571
rect 180 570 181 571
rect 190 571 196 572
rect 190 570 191 571
rect 180 568 191 570
rect 180 567 181 568
rect 175 566 181 567
rect 190 567 191 568
rect 195 567 196 571
rect 223 571 229 572
rect 223 567 224 571
rect 228 570 229 571
rect 239 571 245 572
rect 239 570 240 571
rect 228 568 240 570
rect 228 567 229 568
rect 190 566 196 567
rect 198 566 204 567
rect 223 566 229 567
rect 239 567 240 568
rect 244 567 245 571
rect 295 571 301 572
rect 295 567 296 571
rect 300 570 301 571
rect 311 571 317 572
rect 311 570 312 571
rect 300 568 312 570
rect 300 567 301 568
rect 239 566 245 567
rect 262 566 268 567
rect 295 566 301 567
rect 311 567 312 568
rect 316 567 317 571
rect 390 571 397 572
rect 390 567 391 571
rect 396 567 397 571
rect 471 571 477 572
rect 471 567 472 571
rect 476 570 477 571
rect 487 571 493 572
rect 487 570 488 571
rect 476 568 488 570
rect 476 567 477 568
rect 311 566 317 567
rect 334 566 340 567
rect 390 566 397 567
rect 414 566 420 567
rect 471 566 477 567
rect 487 567 488 568
rect 492 567 493 571
rect 530 571 536 572
rect 530 567 531 571
rect 535 570 536 571
rect 591 571 597 572
rect 591 570 592 571
rect 535 568 592 570
rect 535 567 536 568
rect 487 566 493 567
rect 510 566 516 567
rect 530 566 536 567
rect 591 567 592 568
rect 596 567 597 571
rect 695 571 701 572
rect 695 567 696 571
rect 700 570 701 571
rect 713 570 715 576
rect 846 575 847 576
rect 851 575 852 579
rect 1198 579 1204 580
rect 1198 578 1199 579
rect 846 574 852 575
rect 1056 576 1199 578
rect 700 568 715 570
rect 806 571 813 572
rect 700 567 701 568
rect 806 567 807 571
rect 812 567 813 571
rect 918 571 925 572
rect 918 567 919 571
rect 924 567 925 571
rect 1039 571 1045 572
rect 1039 567 1040 571
rect 1044 570 1045 571
rect 1056 570 1058 576
rect 1198 575 1199 576
rect 1203 575 1204 579
rect 1198 574 1204 575
rect 1422 575 1428 576
rect 1422 574 1423 575
rect 1280 572 1423 574
rect 1044 568 1058 570
rect 1158 571 1165 572
rect 1044 567 1045 568
rect 1158 567 1159 571
rect 1164 567 1165 571
rect 1263 571 1269 572
rect 1263 567 1264 571
rect 1268 570 1269 571
rect 1280 570 1282 572
rect 1422 571 1423 572
rect 1427 571 1428 575
rect 1654 575 1660 576
rect 1654 574 1655 575
rect 1422 570 1428 571
rect 1544 572 1655 574
rect 1268 568 1282 570
rect 1268 567 1269 568
rect 1390 567 1397 568
rect 591 566 597 567
rect 614 566 620 567
rect 695 566 701 567
rect 718 566 724 567
rect 806 566 813 567
rect 830 566 836 567
rect 918 566 925 567
rect 942 566 948 567
rect 1039 566 1045 567
rect 1062 566 1068 567
rect 1158 566 1165 567
rect 1182 566 1188 567
rect 1263 566 1269 567
rect 1286 566 1292 567
rect 198 562 199 566
rect 203 562 204 566
rect 198 561 204 562
rect 262 562 263 566
rect 267 562 268 566
rect 262 561 268 562
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 414 562 415 566
rect 419 562 420 566
rect 414 561 420 562
rect 510 562 511 566
rect 515 562 516 566
rect 510 561 516 562
rect 614 562 615 566
rect 619 562 620 566
rect 614 561 620 562
rect 718 562 719 566
rect 723 562 724 566
rect 718 561 724 562
rect 830 562 831 566
rect 835 562 836 566
rect 830 561 836 562
rect 942 562 943 566
rect 947 562 948 566
rect 942 561 948 562
rect 1062 562 1063 566
rect 1067 562 1068 566
rect 1062 561 1068 562
rect 1182 562 1183 566
rect 1187 562 1188 566
rect 1182 561 1188 562
rect 1286 562 1287 566
rect 1291 562 1292 566
rect 1390 563 1391 567
rect 1396 563 1397 567
rect 1434 567 1440 568
rect 1434 563 1435 567
rect 1439 566 1440 567
rect 1447 567 1453 568
rect 1447 566 1448 567
rect 1439 564 1448 566
rect 1439 563 1440 564
rect 1390 562 1397 563
rect 1414 562 1420 563
rect 1434 562 1440 563
rect 1447 563 1448 564
rect 1452 563 1453 567
rect 1527 567 1533 568
rect 1527 563 1528 567
rect 1532 566 1533 567
rect 1544 566 1546 572
rect 1654 571 1655 572
rect 1659 571 1660 575
rect 2414 575 2420 576
rect 2414 574 2415 575
rect 1654 570 1660 571
rect 2312 572 2415 574
rect 1532 564 1546 566
rect 1622 567 1629 568
rect 1532 563 1533 564
rect 1622 563 1623 567
rect 1628 563 1629 567
rect 1718 567 1724 568
rect 1718 563 1719 567
rect 1723 566 1724 567
rect 1727 567 1733 568
rect 1727 566 1728 567
rect 1723 564 1728 566
rect 1723 563 1724 564
rect 1447 562 1453 563
rect 1470 562 1476 563
rect 1527 562 1533 563
rect 1550 562 1556 563
rect 1622 562 1629 563
rect 1646 562 1652 563
rect 1718 562 1724 563
rect 1727 563 1728 564
rect 1732 563 1733 567
rect 1770 567 1776 568
rect 1770 563 1771 567
rect 1775 566 1776 567
rect 1831 567 1837 568
rect 1831 566 1832 567
rect 1775 564 1832 566
rect 1775 563 1776 564
rect 1727 562 1733 563
rect 1750 562 1756 563
rect 1770 562 1776 563
rect 1831 563 1832 564
rect 1836 563 1837 567
rect 1935 567 1944 568
rect 1935 563 1936 567
rect 1943 563 1944 567
rect 1983 567 1989 568
rect 1983 563 1984 567
rect 1988 566 1989 567
rect 2031 567 2037 568
rect 2031 566 2032 567
rect 1988 564 2032 566
rect 1988 563 1989 564
rect 1831 562 1837 563
rect 1854 562 1860 563
rect 1935 562 1944 563
rect 1958 562 1964 563
rect 1983 562 1989 563
rect 2031 563 2032 564
rect 2036 563 2037 567
rect 2074 567 2080 568
rect 2074 563 2075 567
rect 2079 566 2080 567
rect 2127 567 2133 568
rect 2127 566 2128 567
rect 2079 564 2128 566
rect 2079 563 2080 564
rect 2031 562 2037 563
rect 2054 562 2060 563
rect 2074 562 2080 563
rect 2127 563 2128 564
rect 2132 563 2133 567
rect 2214 567 2221 568
rect 2214 563 2215 567
rect 2220 563 2221 567
rect 2295 567 2301 568
rect 2295 563 2296 567
rect 2300 566 2301 567
rect 2312 566 2314 572
rect 2414 571 2415 572
rect 2419 571 2420 575
rect 2414 570 2420 571
rect 2300 564 2314 566
rect 2374 567 2381 568
rect 2300 563 2301 564
rect 2374 563 2375 567
rect 2380 563 2381 567
rect 2434 567 2440 568
rect 2434 563 2435 567
rect 2439 566 2440 567
rect 2455 567 2461 568
rect 2455 566 2456 567
rect 2439 564 2456 566
rect 2439 563 2440 564
rect 2127 562 2133 563
rect 2150 562 2156 563
rect 2214 562 2221 563
rect 2238 562 2244 563
rect 2295 562 2301 563
rect 2318 562 2324 563
rect 2374 562 2381 563
rect 2398 562 2404 563
rect 2434 562 2440 563
rect 2455 563 2456 564
rect 2460 563 2461 567
rect 2498 567 2504 568
rect 2498 563 2499 567
rect 2503 566 2504 567
rect 2519 567 2525 568
rect 2519 566 2520 567
rect 2503 564 2520 566
rect 2503 563 2504 564
rect 2455 562 2461 563
rect 2478 562 2484 563
rect 2498 562 2504 563
rect 2519 563 2520 564
rect 2524 563 2525 567
rect 2519 562 2525 563
rect 2542 562 2548 563
rect 1286 561 1292 562
rect 1414 558 1415 562
rect 1419 558 1420 562
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 110 552 116 553
rect 1326 557 1332 558
rect 1414 557 1420 558
rect 1470 558 1471 562
rect 1475 558 1476 562
rect 1470 557 1476 558
rect 1550 558 1551 562
rect 1555 558 1556 562
rect 1550 557 1556 558
rect 1646 558 1647 562
rect 1651 558 1652 562
rect 1646 557 1652 558
rect 1750 558 1751 562
rect 1755 558 1756 562
rect 1750 557 1756 558
rect 1854 558 1855 562
rect 1859 558 1860 562
rect 1854 557 1860 558
rect 1958 558 1959 562
rect 1963 558 1964 562
rect 1958 557 1964 558
rect 2054 558 2055 562
rect 2059 558 2060 562
rect 2054 557 2060 558
rect 2150 558 2151 562
rect 2155 558 2156 562
rect 2150 557 2156 558
rect 2238 558 2239 562
rect 2243 558 2244 562
rect 2238 557 2244 558
rect 2318 558 2319 562
rect 2323 558 2324 562
rect 2318 557 2324 558
rect 2398 558 2399 562
rect 2403 558 2404 562
rect 2398 557 2404 558
rect 2478 558 2479 562
rect 2483 558 2484 562
rect 2478 557 2484 558
rect 2542 558 2543 562
rect 2547 558 2548 562
rect 2542 557 2548 558
rect 1326 553 1327 557
rect 1331 553 1332 557
rect 1326 552 1332 553
rect 1366 553 1372 554
rect 1366 549 1367 553
rect 1371 549 1372 553
rect 1366 548 1372 549
rect 2582 553 2588 554
rect 2582 549 2583 553
rect 2587 549 2588 553
rect 2582 548 2588 549
rect 390 547 396 548
rect 390 543 391 547
rect 395 546 396 547
rect 806 547 812 548
rect 395 544 626 546
rect 395 543 396 544
rect 390 542 396 543
rect 110 540 116 541
rect 110 536 111 540
rect 115 536 116 540
rect 110 535 116 536
rect 182 539 188 540
rect 182 535 183 539
rect 187 535 188 539
rect 223 539 229 540
rect 223 538 224 539
rect 182 534 188 535
rect 215 537 224 538
rect 215 533 216 537
rect 220 536 224 537
rect 220 533 221 536
rect 223 535 224 536
rect 228 535 229 539
rect 223 534 229 535
rect 246 539 252 540
rect 246 535 247 539
rect 251 535 252 539
rect 318 539 324 540
rect 246 534 252 535
rect 279 535 285 536
rect 215 532 221 533
rect 279 531 280 535
rect 284 534 285 535
rect 295 535 301 536
rect 295 534 296 535
rect 284 532 296 534
rect 284 531 285 532
rect 279 530 285 531
rect 295 531 296 532
rect 300 531 301 535
rect 318 535 319 539
rect 323 535 324 539
rect 398 539 404 540
rect 318 534 324 535
rect 351 535 360 536
rect 295 530 301 531
rect 351 531 352 535
rect 359 531 360 535
rect 398 535 399 539
rect 403 535 404 539
rect 494 539 500 540
rect 398 534 404 535
rect 431 535 437 536
rect 431 534 432 535
rect 351 530 360 531
rect 408 532 432 534
rect 190 527 196 528
rect 190 523 191 527
rect 195 526 196 527
rect 408 526 410 532
rect 431 531 432 532
rect 436 531 437 535
rect 494 535 495 539
rect 499 535 500 539
rect 598 539 604 540
rect 494 534 500 535
rect 527 535 536 536
rect 431 530 437 531
rect 527 531 528 535
rect 535 531 536 535
rect 598 535 599 539
rect 603 535 604 539
rect 598 534 604 535
rect 624 534 626 544
rect 806 543 807 547
rect 811 546 812 547
rect 1158 547 1164 548
rect 811 544 954 546
rect 811 543 812 544
rect 806 542 812 543
rect 702 539 708 540
rect 631 535 637 536
rect 631 534 632 535
rect 624 532 632 534
rect 527 530 536 531
rect 631 531 632 532
rect 636 531 637 535
rect 702 535 703 539
rect 707 535 708 539
rect 814 539 820 540
rect 702 534 708 535
rect 726 535 732 536
rect 631 530 637 531
rect 726 531 727 535
rect 731 534 732 535
rect 735 535 741 536
rect 735 534 736 535
rect 731 532 736 534
rect 731 531 732 532
rect 726 530 732 531
rect 735 531 736 532
rect 740 531 741 535
rect 814 535 815 539
rect 819 535 820 539
rect 926 539 932 540
rect 814 534 820 535
rect 846 535 853 536
rect 735 530 741 531
rect 846 531 847 535
rect 852 531 853 535
rect 926 535 927 539
rect 931 535 932 539
rect 926 534 932 535
rect 952 534 954 544
rect 1158 543 1159 547
rect 1163 546 1164 547
rect 1163 544 1298 546
rect 1163 543 1164 544
rect 1158 542 1164 543
rect 1046 539 1052 540
rect 959 535 965 536
rect 959 534 960 535
rect 952 532 960 534
rect 846 530 853 531
rect 959 531 960 532
rect 964 531 965 535
rect 1046 535 1047 539
rect 1051 535 1052 539
rect 1166 539 1172 540
rect 1046 534 1052 535
rect 1070 535 1076 536
rect 959 530 965 531
rect 1070 531 1071 535
rect 1075 534 1076 535
rect 1079 535 1085 536
rect 1079 534 1080 535
rect 1075 532 1080 534
rect 1075 531 1076 532
rect 1070 530 1076 531
rect 1079 531 1080 532
rect 1084 531 1085 535
rect 1166 535 1167 539
rect 1171 535 1172 539
rect 1270 539 1276 540
rect 1166 534 1172 535
rect 1198 535 1205 536
rect 1079 530 1085 531
rect 1198 531 1199 535
rect 1204 531 1205 535
rect 1270 535 1271 539
rect 1275 535 1276 539
rect 1270 534 1276 535
rect 1296 534 1298 544
rect 1390 543 1396 544
rect 1326 540 1332 541
rect 1326 536 1327 540
rect 1331 536 1332 540
rect 1390 539 1391 543
rect 1395 542 1396 543
rect 1622 543 1628 544
rect 1395 540 1562 542
rect 1395 539 1396 540
rect 1390 538 1396 539
rect 1303 535 1309 536
rect 1326 535 1332 536
rect 1366 536 1372 537
rect 1303 534 1304 535
rect 1296 532 1304 534
rect 1198 530 1205 531
rect 1303 531 1304 532
rect 1308 531 1309 535
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1398 535 1404 536
rect 1398 531 1399 535
rect 1403 531 1404 535
rect 1454 535 1460 536
rect 1303 530 1309 531
rect 1398 530 1404 531
rect 1431 531 1440 532
rect 1431 527 1432 531
rect 1439 527 1440 531
rect 1454 531 1455 535
rect 1459 531 1460 535
rect 1534 535 1540 536
rect 1454 530 1460 531
rect 1487 531 1496 532
rect 1431 526 1440 527
rect 1487 527 1488 531
rect 1495 527 1496 531
rect 1534 531 1535 535
rect 1539 531 1540 535
rect 1534 530 1540 531
rect 1560 530 1562 540
rect 1622 539 1623 543
rect 1627 542 1628 543
rect 2214 543 2220 544
rect 1627 540 1866 542
rect 1627 539 1628 540
rect 1622 538 1628 539
rect 1630 535 1636 536
rect 1567 531 1573 532
rect 1567 530 1568 531
rect 1560 528 1568 530
rect 1487 526 1496 527
rect 1567 527 1568 528
rect 1572 527 1573 531
rect 1630 531 1631 535
rect 1635 531 1636 535
rect 1734 535 1740 536
rect 1630 530 1636 531
rect 1654 531 1660 532
rect 1567 526 1573 527
rect 1654 527 1655 531
rect 1659 530 1660 531
rect 1663 531 1669 532
rect 1663 530 1664 531
rect 1659 528 1664 530
rect 1659 527 1660 528
rect 1654 526 1660 527
rect 1663 527 1664 528
rect 1668 527 1669 531
rect 1734 531 1735 535
rect 1739 531 1740 535
rect 1838 535 1844 536
rect 1734 530 1740 531
rect 1767 531 1776 532
rect 1663 526 1669 527
rect 1767 527 1768 531
rect 1775 527 1776 531
rect 1838 531 1839 535
rect 1843 531 1844 535
rect 1838 530 1844 531
rect 1864 530 1866 540
rect 2214 539 2215 543
rect 2219 542 2220 543
rect 2374 543 2380 544
rect 2219 540 2330 542
rect 2219 539 2220 540
rect 2214 538 2220 539
rect 1942 535 1948 536
rect 1871 531 1877 532
rect 1871 530 1872 531
rect 1864 528 1872 530
rect 1767 526 1776 527
rect 1871 527 1872 528
rect 1876 527 1877 531
rect 1942 531 1943 535
rect 1947 531 1948 535
rect 2038 535 2044 536
rect 1942 530 1948 531
rect 1975 531 1981 532
rect 1871 526 1877 527
rect 1975 527 1976 531
rect 1980 530 1981 531
rect 1983 531 1989 532
rect 1983 530 1984 531
rect 1980 528 1984 530
rect 1980 527 1981 528
rect 1975 526 1981 527
rect 1983 527 1984 528
rect 1988 527 1989 531
rect 2038 531 2039 535
rect 2043 531 2044 535
rect 2134 535 2140 536
rect 2038 530 2044 531
rect 2071 531 2080 532
rect 1983 526 1989 527
rect 2071 527 2072 531
rect 2079 527 2080 531
rect 2134 531 2135 535
rect 2139 531 2140 535
rect 2222 535 2228 536
rect 2134 530 2140 531
rect 2167 531 2173 532
rect 2167 530 2168 531
rect 2071 526 2080 527
rect 2144 528 2168 530
rect 195 524 410 526
rect 195 523 196 524
rect 190 522 196 523
rect 2022 523 2028 524
rect 2022 519 2023 523
rect 2027 522 2028 523
rect 2144 522 2146 528
rect 2167 527 2168 528
rect 2172 527 2173 531
rect 2222 531 2223 535
rect 2227 531 2228 535
rect 2302 535 2308 536
rect 2222 530 2228 531
rect 2254 531 2261 532
rect 2167 526 2173 527
rect 2254 527 2255 531
rect 2260 527 2261 531
rect 2302 531 2303 535
rect 2307 531 2308 535
rect 2302 530 2308 531
rect 2328 530 2330 540
rect 2374 539 2375 543
rect 2379 542 2380 543
rect 2379 540 2563 542
rect 2379 539 2380 540
rect 2374 538 2380 539
rect 2382 535 2388 536
rect 2335 531 2341 532
rect 2335 530 2336 531
rect 2328 528 2336 530
rect 2254 526 2261 527
rect 2335 527 2336 528
rect 2340 527 2341 531
rect 2382 531 2383 535
rect 2387 531 2388 535
rect 2462 535 2468 536
rect 2382 530 2388 531
rect 2414 531 2421 532
rect 2335 526 2341 527
rect 2414 527 2415 531
rect 2420 527 2421 531
rect 2462 531 2463 535
rect 2467 531 2468 535
rect 2526 535 2532 536
rect 2462 530 2468 531
rect 2495 531 2504 532
rect 2414 526 2421 527
rect 2495 527 2496 531
rect 2503 527 2504 531
rect 2526 531 2527 535
rect 2531 531 2532 535
rect 2561 532 2563 540
rect 2582 536 2588 537
rect 2582 532 2583 536
rect 2587 532 2588 536
rect 2526 530 2532 531
rect 2559 531 2565 532
rect 2582 531 2588 532
rect 2495 526 2504 527
rect 2559 527 2560 531
rect 2564 527 2565 531
rect 2559 526 2565 527
rect 2027 520 2146 522
rect 2027 519 2028 520
rect 2022 518 2028 519
rect 1542 511 1548 512
rect 518 507 524 508
rect 518 503 519 507
rect 523 506 524 507
rect 1542 507 1543 511
rect 1547 510 1548 511
rect 1547 508 1954 510
rect 1547 507 1548 508
rect 1542 506 1548 507
rect 523 504 674 506
rect 523 503 524 504
rect 518 502 524 503
rect 335 499 341 500
rect 302 497 308 498
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 302 493 303 497
rect 307 493 308 497
rect 335 495 336 499
rect 340 498 341 499
rect 350 499 356 500
rect 350 498 351 499
rect 340 496 351 498
rect 340 495 341 496
rect 335 494 341 495
rect 350 495 351 496
rect 355 495 356 499
rect 391 499 397 500
rect 350 494 356 495
rect 358 497 364 498
rect 302 492 308 493
rect 358 493 359 497
rect 363 493 364 497
rect 391 495 392 499
rect 396 498 397 499
rect 414 499 420 500
rect 414 498 415 499
rect 396 496 415 498
rect 396 495 397 496
rect 391 494 397 495
rect 414 495 415 496
rect 419 495 420 499
rect 455 499 461 500
rect 414 494 420 495
rect 422 497 428 498
rect 358 492 364 493
rect 422 493 423 497
rect 427 493 428 497
rect 455 495 456 499
rect 460 498 461 499
rect 471 499 477 500
rect 471 498 472 499
rect 460 496 472 498
rect 460 495 461 496
rect 455 494 461 495
rect 471 495 472 496
rect 476 495 477 499
rect 526 499 533 500
rect 471 494 477 495
rect 494 497 500 498
rect 422 492 428 493
rect 494 493 495 497
rect 499 493 500 497
rect 526 495 527 499
rect 532 495 533 499
rect 607 499 613 500
rect 526 494 533 495
rect 574 497 580 498
rect 494 492 500 493
rect 574 493 575 497
rect 579 493 580 497
rect 607 495 608 499
rect 612 498 613 499
rect 638 499 644 500
rect 638 498 639 499
rect 612 496 639 498
rect 612 495 613 496
rect 607 494 613 495
rect 638 495 639 496
rect 643 495 644 499
rect 672 498 674 504
rect 1567 503 1573 504
rect 1534 501 1540 502
rect 1366 500 1372 501
rect 679 499 685 500
rect 679 498 680 499
rect 638 494 644 495
rect 646 497 652 498
rect 574 492 580 493
rect 646 493 647 497
rect 651 493 652 497
rect 672 496 680 498
rect 679 495 680 496
rect 684 495 685 499
rect 751 499 757 500
rect 679 494 685 495
rect 718 497 724 498
rect 646 492 652 493
rect 718 493 719 497
rect 723 493 724 497
rect 751 495 752 499
rect 756 498 757 499
rect 774 499 780 500
rect 774 498 775 499
rect 756 496 775 498
rect 756 495 757 496
rect 751 494 757 495
rect 774 495 775 496
rect 779 495 780 499
rect 823 499 829 500
rect 774 494 780 495
rect 790 497 796 498
rect 718 492 724 493
rect 790 493 791 497
rect 795 493 796 497
rect 823 495 824 499
rect 828 498 829 499
rect 854 499 860 500
rect 854 498 855 499
rect 828 496 855 498
rect 828 495 829 496
rect 823 494 829 495
rect 854 495 855 496
rect 859 495 860 499
rect 895 499 901 500
rect 854 494 860 495
rect 862 497 868 498
rect 790 492 796 493
rect 862 493 863 497
rect 867 493 868 497
rect 895 495 896 499
rect 900 498 901 499
rect 926 499 932 500
rect 926 498 927 499
rect 900 496 927 498
rect 900 495 901 496
rect 895 494 901 495
rect 926 495 927 496
rect 931 495 932 499
rect 967 499 973 500
rect 926 494 932 495
rect 934 497 940 498
rect 862 492 868 493
rect 934 493 935 497
rect 939 493 940 497
rect 967 495 968 499
rect 972 498 973 499
rect 998 499 1004 500
rect 998 498 999 499
rect 972 496 999 498
rect 972 495 973 496
rect 967 494 973 495
rect 998 495 999 496
rect 1003 495 1004 499
rect 1039 499 1045 500
rect 998 494 1004 495
rect 1006 497 1012 498
rect 934 492 940 493
rect 1006 493 1007 497
rect 1011 493 1012 497
rect 1039 495 1040 499
rect 1044 498 1045 499
rect 1078 499 1084 500
rect 1078 498 1079 499
rect 1044 496 1079 498
rect 1044 495 1045 496
rect 1039 494 1045 495
rect 1078 495 1079 496
rect 1083 495 1084 499
rect 1110 499 1116 500
rect 1078 494 1084 495
rect 1086 497 1092 498
rect 1006 492 1012 493
rect 1086 493 1087 497
rect 1091 493 1092 497
rect 1110 495 1111 499
rect 1115 498 1116 499
rect 1119 499 1125 500
rect 1119 498 1120 499
rect 1115 496 1120 498
rect 1115 495 1116 496
rect 1110 494 1116 495
rect 1119 495 1120 496
rect 1124 495 1125 499
rect 1119 494 1125 495
rect 1326 496 1332 497
rect 1086 492 1092 493
rect 1326 492 1327 496
rect 1331 492 1332 496
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1534 497 1535 501
rect 1539 497 1540 501
rect 1567 499 1568 503
rect 1572 502 1573 503
rect 1590 503 1596 504
rect 1590 502 1591 503
rect 1572 500 1591 502
rect 1572 499 1573 500
rect 1567 498 1573 499
rect 1590 499 1591 500
rect 1595 499 1596 503
rect 1631 503 1637 504
rect 1590 498 1596 499
rect 1598 501 1604 502
rect 1534 496 1540 497
rect 1598 497 1599 501
rect 1603 497 1604 501
rect 1631 499 1632 503
rect 1636 502 1637 503
rect 1662 503 1668 504
rect 1662 502 1663 503
rect 1636 500 1663 502
rect 1636 499 1637 500
rect 1631 498 1637 499
rect 1662 499 1663 500
rect 1667 499 1668 503
rect 1703 503 1709 504
rect 1662 498 1668 499
rect 1670 501 1676 502
rect 1598 496 1604 497
rect 1670 497 1671 501
rect 1675 497 1676 501
rect 1703 499 1704 503
rect 1708 502 1709 503
rect 1718 503 1724 504
rect 1718 502 1719 503
rect 1708 500 1719 502
rect 1708 499 1709 500
rect 1703 498 1709 499
rect 1718 499 1719 500
rect 1723 499 1724 503
rect 1783 503 1789 504
rect 1718 498 1724 499
rect 1750 501 1756 502
rect 1670 496 1676 497
rect 1750 497 1751 501
rect 1755 497 1756 501
rect 1783 499 1784 503
rect 1788 502 1789 503
rect 1830 503 1836 504
rect 1830 502 1831 503
rect 1788 500 1831 502
rect 1788 499 1789 500
rect 1783 498 1789 499
rect 1830 499 1831 500
rect 1835 499 1836 503
rect 1871 503 1877 504
rect 1830 498 1836 499
rect 1838 501 1844 502
rect 1750 496 1756 497
rect 1838 497 1839 501
rect 1843 497 1844 501
rect 1871 499 1872 503
rect 1876 502 1877 503
rect 1918 503 1924 504
rect 1918 502 1919 503
rect 1876 500 1919 502
rect 1876 499 1877 500
rect 1871 498 1877 499
rect 1918 499 1919 500
rect 1923 499 1924 503
rect 1952 502 1954 508
rect 2511 507 2517 508
rect 1959 503 1965 504
rect 1959 502 1960 503
rect 1918 498 1924 499
rect 1926 501 1932 502
rect 1838 496 1844 497
rect 1926 497 1927 501
rect 1931 497 1932 501
rect 1952 500 1960 502
rect 1959 499 1960 500
rect 1964 499 1965 503
rect 2047 503 2053 504
rect 1959 498 1965 499
rect 2014 501 2020 502
rect 1926 496 1932 497
rect 2014 497 2015 501
rect 2019 497 2020 501
rect 2047 499 2048 503
rect 2052 502 2053 503
rect 2086 503 2092 504
rect 2086 502 2087 503
rect 2052 500 2087 502
rect 2052 499 2053 500
rect 2047 498 2053 499
rect 2086 499 2087 500
rect 2091 499 2092 503
rect 2127 503 2133 504
rect 2086 498 2092 499
rect 2094 501 2100 502
rect 2014 496 2020 497
rect 2094 497 2095 501
rect 2099 497 2100 501
rect 2127 499 2128 503
rect 2132 502 2133 503
rect 2166 503 2172 504
rect 2166 502 2167 503
rect 2132 500 2167 502
rect 2132 499 2133 500
rect 2127 498 2133 499
rect 2166 499 2167 500
rect 2171 499 2172 503
rect 2198 503 2204 504
rect 2166 498 2172 499
rect 2174 501 2180 502
rect 2094 496 2100 497
rect 2174 497 2175 501
rect 2179 497 2180 501
rect 2198 499 2199 503
rect 2203 502 2204 503
rect 2207 503 2213 504
rect 2207 502 2208 503
rect 2203 500 2208 502
rect 2203 499 2204 500
rect 2198 498 2204 499
rect 2207 499 2208 500
rect 2212 499 2213 503
rect 2287 503 2293 504
rect 2207 498 2213 499
rect 2254 501 2260 502
rect 2174 496 2180 497
rect 2254 497 2255 501
rect 2259 497 2260 501
rect 2287 499 2288 503
rect 2292 502 2293 503
rect 2318 503 2324 504
rect 2318 502 2319 503
rect 2292 500 2319 502
rect 2292 499 2293 500
rect 2287 498 2293 499
rect 2318 499 2319 500
rect 2323 499 2324 503
rect 2359 503 2365 504
rect 2318 498 2324 499
rect 2326 501 2332 502
rect 2254 496 2260 497
rect 2326 497 2327 501
rect 2331 497 2332 501
rect 2359 499 2360 503
rect 2364 502 2365 503
rect 2390 503 2396 504
rect 2390 502 2391 503
rect 2364 500 2391 502
rect 2364 499 2365 500
rect 2359 498 2365 499
rect 2390 499 2391 500
rect 2395 499 2396 503
rect 2431 503 2440 504
rect 2390 498 2396 499
rect 2398 501 2404 502
rect 2326 496 2332 497
rect 2398 497 2399 501
rect 2403 497 2404 501
rect 2431 499 2432 503
rect 2439 499 2440 503
rect 2494 503 2500 504
rect 2431 498 2440 499
rect 2470 501 2476 502
rect 2398 496 2404 497
rect 2470 497 2471 501
rect 2475 497 2476 501
rect 2494 499 2495 503
rect 2499 502 2500 503
rect 2503 503 2509 504
rect 2503 502 2504 503
rect 2499 500 2504 502
rect 2499 499 2500 500
rect 2494 498 2500 499
rect 2503 499 2504 500
rect 2508 499 2509 503
rect 2511 503 2512 507
rect 2516 506 2517 507
rect 2516 504 2563 506
rect 2516 503 2517 504
rect 2511 502 2517 503
rect 2559 503 2565 504
rect 2503 498 2509 499
rect 2526 501 2532 502
rect 2470 496 2476 497
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2559 499 2560 503
rect 2564 499 2565 503
rect 2559 498 2565 499
rect 2582 500 2588 501
rect 2526 496 2532 497
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 1366 495 1372 496
rect 2582 495 2588 496
rect 110 491 116 492
rect 1326 491 1332 492
rect 1366 483 1372 484
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 1326 479 1332 480
rect 1326 475 1327 479
rect 1331 475 1332 479
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 1326 474 1332 475
rect 1550 474 1556 475
rect 318 470 324 471
rect 318 466 319 470
rect 323 466 324 470
rect 318 465 324 466
rect 374 470 380 471
rect 374 466 375 470
rect 379 466 380 470
rect 374 465 380 466
rect 438 470 444 471
rect 438 466 439 470
rect 443 466 444 470
rect 438 465 444 466
rect 510 470 516 471
rect 510 466 511 470
rect 515 466 516 470
rect 510 465 516 466
rect 590 470 596 471
rect 590 466 591 470
rect 595 466 596 470
rect 590 465 596 466
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 662 465 668 466
rect 734 470 740 471
rect 734 466 735 470
rect 739 466 740 470
rect 734 465 740 466
rect 806 470 812 471
rect 806 466 807 470
rect 811 466 812 470
rect 806 465 812 466
rect 878 470 884 471
rect 878 466 879 470
rect 883 466 884 470
rect 878 465 884 466
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 950 465 956 466
rect 1022 470 1028 471
rect 1022 466 1023 470
rect 1027 466 1028 470
rect 1022 465 1028 466
rect 1102 470 1108 471
rect 1102 466 1103 470
rect 1107 466 1108 470
rect 1550 470 1551 474
rect 1555 470 1556 474
rect 1550 469 1556 470
rect 1614 474 1620 475
rect 1614 470 1615 474
rect 1619 470 1620 474
rect 1614 469 1620 470
rect 1686 474 1692 475
rect 1686 470 1687 474
rect 1691 470 1692 474
rect 1686 469 1692 470
rect 1766 474 1772 475
rect 1766 470 1767 474
rect 1771 470 1772 474
rect 1766 469 1772 470
rect 1854 474 1860 475
rect 1854 470 1855 474
rect 1859 470 1860 474
rect 1854 469 1860 470
rect 1942 474 1948 475
rect 1942 470 1943 474
rect 1947 470 1948 474
rect 1942 469 1948 470
rect 2030 474 2036 475
rect 2030 470 2031 474
rect 2035 470 2036 474
rect 2030 469 2036 470
rect 2110 474 2116 475
rect 2110 470 2111 474
rect 2115 470 2116 474
rect 2110 469 2116 470
rect 2190 474 2196 475
rect 2190 470 2191 474
rect 2195 470 2196 474
rect 2190 469 2196 470
rect 2270 474 2276 475
rect 2270 470 2271 474
rect 2275 470 2276 474
rect 2270 469 2276 470
rect 2342 474 2348 475
rect 2342 470 2343 474
rect 2347 470 2348 474
rect 2342 469 2348 470
rect 2414 474 2420 475
rect 2414 470 2415 474
rect 2419 470 2420 474
rect 2414 469 2420 470
rect 2486 474 2492 475
rect 2486 470 2487 474
rect 2491 470 2492 474
rect 2486 469 2492 470
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 1102 465 1108 466
rect 1527 467 1533 468
rect 295 463 301 464
rect 295 459 296 463
rect 300 462 301 463
rect 350 463 357 464
rect 300 460 321 462
rect 300 459 301 460
rect 295 458 301 459
rect 319 454 321 460
rect 350 459 351 463
rect 356 459 357 463
rect 350 458 357 459
rect 414 463 421 464
rect 414 459 415 463
rect 420 459 421 463
rect 414 458 421 459
rect 487 463 493 464
rect 487 459 488 463
rect 492 462 493 463
rect 518 463 524 464
rect 518 462 519 463
rect 492 460 519 462
rect 492 459 493 460
rect 487 458 493 459
rect 518 459 519 460
rect 523 459 524 463
rect 518 458 524 459
rect 567 463 573 464
rect 567 459 568 463
rect 572 462 573 463
rect 582 463 588 464
rect 582 462 583 463
rect 572 460 583 462
rect 572 459 573 460
rect 567 458 573 459
rect 582 459 583 460
rect 587 459 588 463
rect 582 458 588 459
rect 638 463 645 464
rect 638 459 639 463
rect 644 459 645 463
rect 638 458 645 459
rect 711 463 717 464
rect 711 459 712 463
rect 716 462 717 463
rect 726 463 732 464
rect 726 462 727 463
rect 716 460 727 462
rect 716 459 717 460
rect 711 458 717 459
rect 726 459 727 460
rect 731 459 732 463
rect 726 458 732 459
rect 774 463 780 464
rect 774 459 775 463
rect 779 462 780 463
rect 783 463 789 464
rect 783 462 784 463
rect 779 460 784 462
rect 779 459 780 460
rect 774 458 780 459
rect 783 459 784 460
rect 788 459 789 463
rect 783 458 789 459
rect 854 463 861 464
rect 854 459 855 463
rect 860 459 861 463
rect 854 458 861 459
rect 926 463 933 464
rect 926 459 927 463
rect 932 459 933 463
rect 926 458 933 459
rect 998 463 1005 464
rect 998 459 999 463
rect 1004 459 1005 463
rect 998 458 1005 459
rect 1078 463 1085 464
rect 1078 459 1079 463
rect 1084 459 1085 463
rect 1527 463 1528 467
rect 1532 466 1533 467
rect 1542 467 1548 468
rect 1542 466 1543 467
rect 1532 464 1543 466
rect 1532 463 1533 464
rect 1527 462 1533 463
rect 1542 463 1543 464
rect 1547 463 1548 467
rect 1542 462 1548 463
rect 1590 467 1597 468
rect 1590 463 1591 467
rect 1596 463 1597 467
rect 1590 462 1597 463
rect 1662 467 1669 468
rect 1662 463 1663 467
rect 1668 463 1669 467
rect 1662 462 1669 463
rect 1743 467 1749 468
rect 1743 463 1744 467
rect 1748 466 1749 467
rect 1774 467 1780 468
rect 1774 466 1775 467
rect 1748 464 1775 466
rect 1748 463 1749 464
rect 1743 462 1749 463
rect 1774 463 1775 464
rect 1779 463 1780 467
rect 1774 462 1780 463
rect 1830 467 1837 468
rect 1830 463 1831 467
rect 1836 463 1837 467
rect 1830 462 1837 463
rect 1918 467 1925 468
rect 1918 463 1919 467
rect 1924 463 1925 467
rect 1918 462 1925 463
rect 2007 467 2013 468
rect 2007 463 2008 467
rect 2012 466 2013 467
rect 2022 467 2028 468
rect 2022 466 2023 467
rect 2012 464 2023 466
rect 2012 463 2013 464
rect 2007 462 2013 463
rect 2022 463 2023 464
rect 2027 463 2028 467
rect 2022 462 2028 463
rect 2086 467 2093 468
rect 2086 463 2087 467
rect 2092 463 2093 467
rect 2086 462 2093 463
rect 2166 467 2173 468
rect 2166 463 2167 467
rect 2172 463 2173 467
rect 2166 462 2173 463
rect 2247 467 2253 468
rect 2247 463 2248 467
rect 2252 463 2253 467
rect 2247 462 2253 463
rect 2318 467 2325 468
rect 2318 463 2319 467
rect 2324 463 2325 467
rect 2318 462 2325 463
rect 2390 467 2397 468
rect 2390 463 2391 467
rect 2396 463 2397 467
rect 2390 462 2397 463
rect 2463 467 2469 468
rect 2463 463 2464 467
rect 2468 466 2469 467
rect 2511 467 2517 468
rect 2511 466 2512 467
rect 2468 464 2512 466
rect 2468 463 2469 464
rect 2463 462 2469 463
rect 2511 463 2512 464
rect 2516 463 2517 467
rect 2511 462 2517 463
rect 2519 467 2525 468
rect 2519 463 2520 467
rect 2524 466 2525 467
rect 2558 467 2564 468
rect 2558 466 2559 467
rect 2524 464 2559 466
rect 2524 463 2525 464
rect 2519 462 2525 463
rect 2558 463 2559 464
rect 2563 463 2564 467
rect 2558 462 2564 463
rect 1078 458 1085 459
rect 2249 458 2251 462
rect 2494 459 2500 460
rect 2494 458 2495 459
rect 2249 456 2495 458
rect 526 455 532 456
rect 526 454 527 455
rect 319 452 527 454
rect 526 451 527 452
rect 531 451 532 455
rect 742 455 748 456
rect 742 454 743 455
rect 526 450 532 451
rect 640 452 743 454
rect 430 447 437 448
rect 430 443 431 447
rect 436 443 437 447
rect 470 447 476 448
rect 470 443 471 447
rect 475 446 476 447
rect 487 447 493 448
rect 487 446 488 447
rect 475 444 488 446
rect 475 443 476 444
rect 430 442 437 443
rect 454 442 460 443
rect 470 442 476 443
rect 487 443 488 444
rect 492 443 493 447
rect 530 447 536 448
rect 530 443 531 447
rect 535 446 536 447
rect 551 447 557 448
rect 551 446 552 447
rect 535 444 552 446
rect 535 443 536 444
rect 487 442 493 443
rect 510 442 516 443
rect 530 442 536 443
rect 551 443 552 444
rect 556 443 557 447
rect 623 447 629 448
rect 623 443 624 447
rect 628 446 629 447
rect 640 446 642 452
rect 742 451 743 452
rect 747 451 748 455
rect 1110 455 1116 456
rect 1110 454 1111 455
rect 742 450 748 451
rect 865 452 1111 454
rect 628 444 642 446
rect 702 447 709 448
rect 628 443 629 444
rect 702 443 703 447
rect 708 443 709 447
rect 775 447 781 448
rect 775 443 776 447
rect 780 446 781 447
rect 790 447 796 448
rect 790 446 791 447
rect 780 444 791 446
rect 780 443 781 444
rect 551 442 557 443
rect 574 442 580 443
rect 623 442 629 443
rect 646 442 652 443
rect 702 442 709 443
rect 726 442 732 443
rect 775 442 781 443
rect 790 443 791 444
rect 795 443 796 447
rect 847 447 853 448
rect 847 443 848 447
rect 852 446 853 447
rect 865 446 867 452
rect 1110 451 1111 452
rect 1115 451 1116 455
rect 1886 455 1892 456
rect 1886 454 1887 455
rect 1110 450 1116 451
rect 1808 452 1887 454
rect 852 444 867 446
rect 890 447 896 448
rect 852 443 853 444
rect 890 443 891 447
rect 895 446 896 447
rect 919 447 925 448
rect 919 446 920 447
rect 895 444 920 446
rect 895 443 896 444
rect 790 442 796 443
rect 798 442 804 443
rect 847 442 853 443
rect 870 442 876 443
rect 890 442 896 443
rect 919 443 920 444
rect 924 443 925 447
rect 962 447 968 448
rect 962 443 963 447
rect 967 446 968 447
rect 991 447 997 448
rect 991 446 992 447
rect 967 444 992 446
rect 967 443 968 444
rect 919 442 925 443
rect 942 442 948 443
rect 962 442 968 443
rect 991 443 992 444
rect 996 443 997 447
rect 1034 447 1040 448
rect 1034 443 1035 447
rect 1039 446 1040 447
rect 1063 447 1069 448
rect 1063 446 1064 447
rect 1039 444 1064 446
rect 1039 443 1040 444
rect 991 442 997 443
rect 1014 442 1020 443
rect 1034 442 1040 443
rect 1063 443 1064 444
rect 1068 443 1069 447
rect 1122 447 1128 448
rect 1122 443 1123 447
rect 1127 446 1128 447
rect 1135 447 1141 448
rect 1135 446 1136 447
rect 1127 444 1136 446
rect 1127 443 1128 444
rect 1063 442 1069 443
rect 1086 442 1092 443
rect 1122 442 1128 443
rect 1135 443 1136 444
rect 1140 443 1141 447
rect 1178 447 1184 448
rect 1178 443 1179 447
rect 1183 446 1184 447
rect 1215 447 1221 448
rect 1215 446 1216 447
rect 1183 444 1216 446
rect 1183 443 1184 444
rect 1135 442 1141 443
rect 1158 442 1164 443
rect 1178 442 1184 443
rect 1215 443 1216 444
rect 1220 443 1221 447
rect 1622 447 1629 448
rect 1622 443 1623 447
rect 1628 443 1629 447
rect 1666 447 1672 448
rect 1666 443 1667 447
rect 1671 446 1672 447
rect 1679 447 1685 448
rect 1679 446 1680 447
rect 1671 444 1680 446
rect 1671 443 1672 444
rect 1215 442 1221 443
rect 1238 442 1244 443
rect 1622 442 1629 443
rect 1646 442 1652 443
rect 1666 442 1672 443
rect 1679 443 1680 444
rect 1684 443 1685 447
rect 1722 447 1728 448
rect 1722 443 1723 447
rect 1727 446 1728 447
rect 1735 447 1741 448
rect 1735 446 1736 447
rect 1727 444 1736 446
rect 1727 443 1728 444
rect 1679 442 1685 443
rect 1702 442 1708 443
rect 1722 442 1728 443
rect 1735 443 1736 444
rect 1740 443 1741 447
rect 1791 447 1797 448
rect 1791 443 1792 447
rect 1796 446 1797 447
rect 1808 446 1810 452
rect 1886 451 1887 452
rect 1891 451 1892 455
rect 2494 455 2495 456
rect 2499 455 2500 459
rect 2494 454 2500 455
rect 1886 450 1892 451
rect 2198 451 2204 452
rect 2198 450 2199 451
rect 2184 448 2199 450
rect 1796 444 1810 446
rect 1846 447 1853 448
rect 1796 443 1797 444
rect 1846 443 1847 447
rect 1852 443 1853 447
rect 1903 447 1909 448
rect 1903 443 1904 447
rect 1908 446 1909 447
rect 1918 447 1924 448
rect 1918 446 1919 447
rect 1908 444 1919 446
rect 1908 443 1909 444
rect 1735 442 1741 443
rect 1758 442 1764 443
rect 1791 442 1797 443
rect 1814 442 1820 443
rect 1846 442 1853 443
rect 1870 442 1876 443
rect 1903 442 1909 443
rect 1918 443 1919 444
rect 1923 443 1924 447
rect 1974 447 1981 448
rect 1974 443 1975 447
rect 1980 443 1981 447
rect 2063 447 2069 448
rect 2063 443 2064 447
rect 2068 446 2069 447
rect 2078 447 2084 448
rect 2078 446 2079 447
rect 2068 444 2079 446
rect 2068 443 2069 444
rect 1918 442 1924 443
rect 1926 442 1932 443
rect 1974 442 1981 443
rect 1998 442 2004 443
rect 2063 442 2069 443
rect 2078 443 2079 444
rect 2083 443 2084 447
rect 2167 447 2173 448
rect 2167 443 2168 447
rect 2172 446 2173 447
rect 2184 446 2186 448
rect 2198 447 2199 448
rect 2203 447 2204 451
rect 2198 446 2204 447
rect 2210 447 2216 448
rect 2172 444 2186 446
rect 2172 443 2173 444
rect 2210 443 2211 447
rect 2215 446 2216 447
rect 2287 447 2293 448
rect 2287 446 2288 447
rect 2215 444 2288 446
rect 2215 443 2216 444
rect 2078 442 2084 443
rect 2086 442 2092 443
rect 2167 442 2173 443
rect 2190 442 2196 443
rect 2210 442 2216 443
rect 2287 443 2288 444
rect 2292 443 2293 447
rect 2330 447 2336 448
rect 2330 443 2331 447
rect 2335 446 2336 447
rect 2415 447 2421 448
rect 2415 446 2416 447
rect 2335 444 2416 446
rect 2335 443 2336 444
rect 2287 442 2293 443
rect 2310 442 2316 443
rect 2330 442 2336 443
rect 2415 443 2416 444
rect 2420 443 2421 447
rect 2519 447 2525 448
rect 2519 443 2520 447
rect 2524 446 2525 447
rect 2534 447 2540 448
rect 2534 446 2535 447
rect 2524 444 2535 446
rect 2524 443 2525 444
rect 2415 442 2421 443
rect 2438 442 2444 443
rect 2519 442 2525 443
rect 2534 443 2535 444
rect 2539 443 2540 447
rect 2534 442 2540 443
rect 2542 442 2548 443
rect 454 438 455 442
rect 459 438 460 442
rect 454 437 460 438
rect 510 438 511 442
rect 515 438 516 442
rect 510 437 516 438
rect 574 438 575 442
rect 579 438 580 442
rect 574 437 580 438
rect 646 438 647 442
rect 651 438 652 442
rect 646 437 652 438
rect 726 438 727 442
rect 731 438 732 442
rect 726 437 732 438
rect 798 438 799 442
rect 803 438 804 442
rect 798 437 804 438
rect 870 438 871 442
rect 875 438 876 442
rect 870 437 876 438
rect 942 438 943 442
rect 947 438 948 442
rect 942 437 948 438
rect 1014 438 1015 442
rect 1019 438 1020 442
rect 1014 437 1020 438
rect 1086 438 1087 442
rect 1091 438 1092 442
rect 1086 437 1092 438
rect 1158 438 1159 442
rect 1163 438 1164 442
rect 1158 437 1164 438
rect 1238 438 1239 442
rect 1243 438 1244 442
rect 1238 437 1244 438
rect 1646 438 1647 442
rect 1651 438 1652 442
rect 1646 437 1652 438
rect 1702 438 1703 442
rect 1707 438 1708 442
rect 1702 437 1708 438
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1814 438 1815 442
rect 1819 438 1820 442
rect 1814 437 1820 438
rect 1870 438 1871 442
rect 1875 438 1876 442
rect 1870 437 1876 438
rect 1926 438 1927 442
rect 1931 438 1932 442
rect 1926 437 1932 438
rect 1998 438 1999 442
rect 2003 438 2004 442
rect 1998 437 2004 438
rect 2086 438 2087 442
rect 2091 438 2092 442
rect 2086 437 2092 438
rect 2190 438 2191 442
rect 2195 438 2196 442
rect 2190 437 2196 438
rect 2310 438 2311 442
rect 2315 438 2316 442
rect 2310 437 2316 438
rect 2438 438 2439 442
rect 2443 438 2444 442
rect 2438 437 2444 438
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 110 428 116 429
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1326 428 1332 429
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 1366 428 1372 429
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 430 423 436 424
rect 430 419 431 423
rect 435 422 436 423
rect 702 423 708 424
rect 435 420 658 422
rect 435 419 436 420
rect 430 418 436 419
rect 110 416 116 417
rect 110 412 111 416
rect 115 412 116 416
rect 110 411 116 412
rect 438 415 444 416
rect 438 411 439 415
rect 443 411 444 415
rect 494 415 500 416
rect 438 410 444 411
rect 470 411 477 412
rect 470 407 471 411
rect 476 407 477 411
rect 494 411 495 415
rect 499 411 500 415
rect 558 415 564 416
rect 494 410 500 411
rect 527 411 536 412
rect 470 406 477 407
rect 527 407 528 411
rect 535 407 536 411
rect 558 411 559 415
rect 563 411 564 415
rect 630 415 636 416
rect 558 410 564 411
rect 582 411 588 412
rect 527 406 536 407
rect 582 407 583 411
rect 587 410 588 411
rect 591 411 597 412
rect 591 410 592 411
rect 587 408 592 410
rect 587 407 588 408
rect 582 406 588 407
rect 591 407 592 408
rect 596 407 597 411
rect 630 411 631 415
rect 635 411 636 415
rect 630 410 636 411
rect 656 410 658 420
rect 702 419 703 423
rect 707 422 708 423
rect 1622 423 1628 424
rect 707 420 810 422
rect 707 419 708 420
rect 702 418 708 419
rect 710 415 716 416
rect 663 411 669 412
rect 663 410 664 411
rect 656 408 664 410
rect 591 406 597 407
rect 663 407 664 408
rect 668 407 669 411
rect 710 411 711 415
rect 715 411 716 415
rect 782 415 788 416
rect 710 410 716 411
rect 742 411 749 412
rect 663 406 669 407
rect 742 407 743 411
rect 748 407 749 411
rect 782 411 783 415
rect 787 411 788 415
rect 782 410 788 411
rect 808 410 810 420
rect 1622 419 1623 423
rect 1627 422 1628 423
rect 1846 423 1852 424
rect 1627 420 1826 422
rect 1627 419 1628 420
rect 1622 418 1628 419
rect 1326 416 1332 417
rect 854 415 860 416
rect 815 411 821 412
rect 815 410 816 411
rect 808 408 816 410
rect 742 406 749 407
rect 815 407 816 408
rect 820 407 821 411
rect 854 411 855 415
rect 859 411 860 415
rect 926 415 932 416
rect 854 410 860 411
rect 887 411 896 412
rect 815 406 821 407
rect 887 407 888 411
rect 895 407 896 411
rect 926 411 927 415
rect 931 411 932 415
rect 998 415 1004 416
rect 926 410 932 411
rect 959 411 968 412
rect 887 406 896 407
rect 959 407 960 411
rect 967 407 968 411
rect 998 411 999 415
rect 1003 411 1004 415
rect 1070 415 1076 416
rect 998 410 1004 411
rect 1031 411 1040 412
rect 959 406 968 407
rect 1031 407 1032 411
rect 1039 407 1040 411
rect 1070 411 1071 415
rect 1075 411 1076 415
rect 1122 415 1128 416
rect 1122 414 1123 415
rect 1070 410 1076 411
rect 1103 413 1123 414
rect 1103 409 1104 413
rect 1108 412 1123 413
rect 1108 409 1109 412
rect 1122 411 1123 412
rect 1127 411 1128 415
rect 1122 410 1128 411
rect 1142 415 1148 416
rect 1142 411 1143 415
rect 1147 411 1148 415
rect 1222 415 1228 416
rect 1142 410 1148 411
rect 1175 411 1184 412
rect 1103 408 1109 409
rect 1031 406 1040 407
rect 1175 407 1176 411
rect 1183 407 1184 411
rect 1222 411 1223 415
rect 1227 411 1228 415
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1222 410 1228 411
rect 1254 411 1261 412
rect 1326 411 1332 412
rect 1366 416 1372 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1630 415 1636 416
rect 1630 411 1631 415
rect 1635 411 1636 415
rect 1686 415 1692 416
rect 1175 406 1184 407
rect 1254 407 1255 411
rect 1260 407 1261 411
rect 1630 410 1636 411
rect 1663 411 1672 412
rect 1254 406 1261 407
rect 1663 407 1664 411
rect 1671 407 1672 411
rect 1686 411 1687 415
rect 1691 411 1692 415
rect 1742 415 1748 416
rect 1686 410 1692 411
rect 1719 411 1728 412
rect 1663 406 1672 407
rect 1719 407 1720 411
rect 1727 407 1728 411
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1798 415 1804 416
rect 1742 410 1748 411
rect 1774 411 1781 412
rect 1719 406 1728 407
rect 1774 407 1775 411
rect 1780 407 1781 411
rect 1798 411 1799 415
rect 1803 411 1804 415
rect 1798 410 1804 411
rect 1824 410 1826 420
rect 1846 419 1847 423
rect 1851 422 1852 423
rect 1974 423 1980 424
rect 1851 420 1938 422
rect 1851 419 1852 420
rect 1846 418 1852 419
rect 1854 415 1860 416
rect 1831 411 1837 412
rect 1831 410 1832 411
rect 1824 408 1832 410
rect 1774 406 1781 407
rect 1831 407 1832 408
rect 1836 407 1837 411
rect 1854 411 1855 415
rect 1859 411 1860 415
rect 1910 415 1916 416
rect 1854 410 1860 411
rect 1886 411 1893 412
rect 1831 406 1837 407
rect 1886 407 1887 411
rect 1892 407 1893 411
rect 1910 411 1911 415
rect 1915 411 1916 415
rect 1910 410 1916 411
rect 1936 410 1938 420
rect 1974 419 1975 423
rect 1979 422 1980 423
rect 1979 420 2098 422
rect 1979 419 1980 420
rect 1974 418 1980 419
rect 1982 415 1988 416
rect 1943 411 1949 412
rect 1943 410 1944 411
rect 1936 408 1944 410
rect 1886 406 1893 407
rect 1943 407 1944 408
rect 1948 407 1949 411
rect 1982 411 1983 415
rect 1987 411 1988 415
rect 2070 415 2076 416
rect 1982 410 1988 411
rect 2015 411 2024 412
rect 1943 406 1949 407
rect 2015 407 2016 411
rect 2023 407 2024 411
rect 2070 411 2071 415
rect 2075 411 2076 415
rect 2070 410 2076 411
rect 2096 410 2098 420
rect 2582 416 2588 417
rect 2174 415 2180 416
rect 2103 411 2109 412
rect 2103 410 2104 411
rect 2096 408 2104 410
rect 2015 406 2024 407
rect 2103 407 2104 408
rect 2108 407 2109 411
rect 2174 411 2175 415
rect 2179 411 2180 415
rect 2294 415 2300 416
rect 2174 410 2180 411
rect 2207 411 2216 412
rect 2103 406 2109 407
rect 2207 407 2208 411
rect 2215 407 2216 411
rect 2294 411 2295 415
rect 2299 411 2300 415
rect 2422 415 2428 416
rect 2294 410 2300 411
rect 2327 411 2336 412
rect 2207 406 2216 407
rect 2327 407 2328 411
rect 2335 407 2336 411
rect 2422 411 2423 415
rect 2427 411 2428 415
rect 2526 415 2532 416
rect 2422 410 2428 411
rect 2454 411 2461 412
rect 2327 406 2336 407
rect 2454 407 2455 411
rect 2460 407 2461 411
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2526 410 2532 411
rect 2558 411 2565 412
rect 2582 411 2588 412
rect 2454 406 2461 407
rect 2558 407 2559 411
rect 2564 407 2565 411
rect 2558 406 2565 407
rect 1918 391 1924 392
rect 934 387 940 388
rect 807 383 813 384
rect 447 379 453 380
rect 414 377 420 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 414 373 415 377
rect 419 373 420 377
rect 447 375 448 379
rect 452 378 453 379
rect 462 379 468 380
rect 462 378 463 379
rect 452 376 463 378
rect 452 375 453 376
rect 447 374 453 375
rect 462 375 463 376
rect 467 375 468 379
rect 503 379 509 380
rect 462 374 468 375
rect 470 377 476 378
rect 414 372 420 373
rect 470 373 471 377
rect 475 373 476 377
rect 503 375 504 379
rect 508 378 509 379
rect 526 379 532 380
rect 526 378 527 379
rect 508 376 527 378
rect 508 375 509 376
rect 503 374 509 375
rect 526 375 527 376
rect 531 375 532 379
rect 567 379 573 380
rect 526 374 532 375
rect 534 377 540 378
rect 470 372 476 373
rect 534 373 535 377
rect 539 373 540 377
rect 567 375 568 379
rect 572 378 573 379
rect 598 379 604 380
rect 598 378 599 379
rect 572 376 599 378
rect 572 375 573 376
rect 567 374 573 375
rect 598 375 599 376
rect 603 375 604 379
rect 639 379 645 380
rect 598 374 604 375
rect 606 377 612 378
rect 534 372 540 373
rect 606 373 607 377
rect 611 373 612 377
rect 639 375 640 379
rect 644 378 645 379
rect 678 379 684 380
rect 678 378 679 379
rect 644 376 679 378
rect 644 375 645 376
rect 639 374 645 375
rect 678 375 679 376
rect 683 375 684 379
rect 710 379 716 380
rect 678 374 684 375
rect 686 377 692 378
rect 606 372 612 373
rect 686 373 687 377
rect 691 373 692 377
rect 710 375 711 379
rect 715 378 716 379
rect 719 379 725 380
rect 719 378 720 379
rect 715 376 720 378
rect 715 375 716 376
rect 710 374 716 375
rect 719 375 720 376
rect 724 375 725 379
rect 790 379 796 380
rect 719 374 725 375
rect 766 377 772 378
rect 686 372 692 373
rect 766 373 767 377
rect 771 373 772 377
rect 790 375 791 379
rect 795 378 796 379
rect 799 379 805 380
rect 799 378 800 379
rect 795 376 800 378
rect 795 375 796 376
rect 790 374 796 375
rect 799 375 800 376
rect 804 375 805 379
rect 807 379 808 383
rect 812 382 813 383
rect 934 383 935 387
rect 939 386 940 387
rect 1918 387 1919 391
rect 1923 390 1924 391
rect 1923 388 1987 390
rect 1923 387 1924 388
rect 1918 386 1924 387
rect 939 384 1114 386
rect 1985 384 1987 388
rect 2534 387 2540 388
rect 939 383 940 384
rect 934 382 940 383
rect 812 380 874 382
rect 812 379 813 380
rect 807 378 813 379
rect 872 378 874 380
rect 879 379 885 380
rect 879 378 880 379
rect 799 374 805 375
rect 846 377 852 378
rect 766 372 772 373
rect 846 373 847 377
rect 851 373 852 377
rect 872 376 880 378
rect 879 375 880 376
rect 884 375 885 379
rect 959 379 965 380
rect 879 374 885 375
rect 926 377 932 378
rect 846 372 852 373
rect 926 373 927 377
rect 931 373 932 377
rect 959 375 960 379
rect 964 378 965 379
rect 998 379 1004 380
rect 998 378 999 379
rect 964 376 999 378
rect 964 375 965 376
rect 959 374 965 375
rect 998 375 999 376
rect 1003 375 1004 379
rect 1039 379 1045 380
rect 998 374 1004 375
rect 1006 377 1012 378
rect 926 372 932 373
rect 1006 373 1007 377
rect 1011 373 1012 377
rect 1039 375 1040 379
rect 1044 378 1045 379
rect 1078 379 1084 380
rect 1078 378 1079 379
rect 1044 376 1079 378
rect 1044 375 1045 376
rect 1039 374 1045 375
rect 1078 375 1079 376
rect 1083 375 1084 379
rect 1112 378 1114 384
rect 1127 383 1133 384
rect 1119 379 1125 380
rect 1119 378 1120 379
rect 1078 374 1084 375
rect 1086 377 1092 378
rect 1006 372 1012 373
rect 1086 373 1087 377
rect 1091 373 1092 377
rect 1112 376 1120 378
rect 1119 375 1120 376
rect 1124 375 1125 379
rect 1127 379 1128 383
rect 1132 382 1133 383
rect 1215 383 1221 384
rect 1132 380 1202 382
rect 1132 379 1133 380
rect 1127 378 1133 379
rect 1200 378 1202 380
rect 1207 379 1213 380
rect 1207 378 1208 379
rect 1119 374 1125 375
rect 1174 377 1180 378
rect 1086 372 1092 373
rect 1174 373 1175 377
rect 1179 373 1180 377
rect 1200 376 1208 378
rect 1207 375 1208 376
rect 1212 375 1213 379
rect 1215 379 1216 383
rect 1220 382 1221 383
rect 1687 383 1693 384
rect 1220 380 1290 382
rect 1654 381 1660 382
rect 1366 380 1372 381
rect 1220 379 1221 380
rect 1215 378 1221 379
rect 1288 378 1290 380
rect 1295 379 1301 380
rect 1295 378 1296 379
rect 1207 374 1213 375
rect 1262 377 1268 378
rect 1174 372 1180 373
rect 1262 373 1263 377
rect 1267 373 1268 377
rect 1288 376 1296 378
rect 1295 375 1296 376
rect 1300 375 1301 379
rect 1295 374 1301 375
rect 1326 376 1332 377
rect 1262 372 1268 373
rect 1326 372 1327 376
rect 1331 372 1332 376
rect 1366 376 1367 380
rect 1371 376 1372 380
rect 1654 377 1655 381
rect 1659 377 1660 381
rect 1687 379 1688 383
rect 1692 382 1693 383
rect 1702 383 1708 384
rect 1702 382 1703 383
rect 1692 380 1703 382
rect 1692 379 1693 380
rect 1687 378 1693 379
rect 1702 379 1703 380
rect 1707 379 1708 383
rect 1743 383 1749 384
rect 1702 378 1708 379
rect 1710 381 1716 382
rect 1654 376 1660 377
rect 1710 377 1711 381
rect 1715 377 1716 381
rect 1743 379 1744 383
rect 1748 382 1749 383
rect 1758 383 1764 384
rect 1758 382 1759 383
rect 1748 380 1759 382
rect 1748 379 1749 380
rect 1743 378 1749 379
rect 1758 379 1759 380
rect 1763 379 1764 383
rect 1799 383 1805 384
rect 1758 378 1764 379
rect 1766 381 1772 382
rect 1710 376 1716 377
rect 1766 377 1767 381
rect 1771 377 1772 381
rect 1799 379 1800 383
rect 1804 382 1805 383
rect 1814 383 1820 384
rect 1814 382 1815 383
rect 1804 380 1815 382
rect 1804 379 1805 380
rect 1799 378 1805 379
rect 1814 379 1815 380
rect 1819 379 1820 383
rect 1855 383 1861 384
rect 1814 378 1820 379
rect 1822 381 1828 382
rect 1766 376 1772 377
rect 1822 377 1823 381
rect 1827 377 1828 381
rect 1855 379 1856 383
rect 1860 382 1861 383
rect 1870 383 1876 384
rect 1870 382 1871 383
rect 1860 380 1871 382
rect 1860 379 1861 380
rect 1855 378 1861 379
rect 1870 379 1871 380
rect 1875 379 1876 383
rect 1911 383 1917 384
rect 1870 378 1876 379
rect 1878 381 1884 382
rect 1822 376 1828 377
rect 1878 377 1879 381
rect 1883 377 1884 381
rect 1911 379 1912 383
rect 1916 382 1917 383
rect 1942 383 1948 384
rect 1942 382 1943 383
rect 1916 380 1943 382
rect 1916 379 1917 380
rect 1911 378 1917 379
rect 1942 379 1943 380
rect 1947 379 1948 383
rect 1983 383 1989 384
rect 1942 378 1948 379
rect 1950 381 1956 382
rect 1878 376 1884 377
rect 1950 377 1951 381
rect 1955 377 1956 381
rect 1983 379 1984 383
rect 1988 379 1989 383
rect 2071 383 2077 384
rect 1983 378 1989 379
rect 2038 381 2044 382
rect 1950 376 1956 377
rect 2038 377 2039 381
rect 2043 377 2044 381
rect 2071 379 2072 383
rect 2076 382 2077 383
rect 2142 383 2148 384
rect 2142 382 2143 383
rect 2076 380 2143 382
rect 2076 379 2077 380
rect 2071 378 2077 379
rect 2142 379 2143 380
rect 2147 379 2148 383
rect 2183 383 2189 384
rect 2142 378 2148 379
rect 2150 381 2156 382
rect 2038 376 2044 377
rect 2150 377 2151 381
rect 2155 377 2156 381
rect 2183 379 2184 383
rect 2188 382 2189 383
rect 2270 383 2276 384
rect 2270 382 2271 383
rect 2188 380 2271 382
rect 2188 379 2189 380
rect 2183 378 2189 379
rect 2270 379 2271 380
rect 2275 379 2276 383
rect 2311 383 2317 384
rect 2270 378 2276 379
rect 2278 381 2284 382
rect 2150 376 2156 377
rect 2278 377 2279 381
rect 2283 377 2284 381
rect 2311 379 2312 383
rect 2316 382 2317 383
rect 2406 383 2412 384
rect 2406 382 2407 383
rect 2316 380 2407 382
rect 2316 379 2317 380
rect 2311 378 2317 379
rect 2406 379 2407 380
rect 2411 379 2412 383
rect 2438 383 2444 384
rect 2406 378 2412 379
rect 2414 381 2420 382
rect 2278 376 2284 377
rect 2414 377 2415 381
rect 2419 377 2420 381
rect 2438 379 2439 383
rect 2443 382 2444 383
rect 2447 383 2453 384
rect 2447 382 2448 383
rect 2443 380 2448 382
rect 2443 379 2444 380
rect 2438 378 2444 379
rect 2447 379 2448 380
rect 2452 379 2453 383
rect 2534 383 2535 387
rect 2539 386 2540 387
rect 2539 384 2563 386
rect 2539 383 2540 384
rect 2534 382 2540 383
rect 2559 383 2565 384
rect 2447 378 2453 379
rect 2526 381 2532 382
rect 2414 376 2420 377
rect 2526 377 2527 381
rect 2531 377 2532 381
rect 2559 379 2560 383
rect 2564 379 2565 383
rect 2559 378 2565 379
rect 2582 380 2588 381
rect 2526 376 2532 377
rect 2582 376 2583 380
rect 2587 376 2588 380
rect 1366 375 1372 376
rect 2582 375 2588 376
rect 110 371 116 372
rect 1326 371 1332 372
rect 1366 363 1372 364
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 1326 359 1332 360
rect 1326 355 1327 359
rect 1331 355 1332 359
rect 1366 359 1367 363
rect 1371 359 1372 363
rect 1366 358 1372 359
rect 2582 363 2588 364
rect 2582 359 2583 363
rect 2587 359 2588 363
rect 2582 358 2588 359
rect 1326 354 1332 355
rect 1670 354 1676 355
rect 430 350 436 351
rect 430 346 431 350
rect 435 346 436 350
rect 430 345 436 346
rect 486 350 492 351
rect 486 346 487 350
rect 491 346 492 350
rect 486 345 492 346
rect 550 350 556 351
rect 550 346 551 350
rect 555 346 556 350
rect 550 345 556 346
rect 622 350 628 351
rect 622 346 623 350
rect 627 346 628 350
rect 622 345 628 346
rect 702 350 708 351
rect 702 346 703 350
rect 707 346 708 350
rect 702 345 708 346
rect 782 350 788 351
rect 782 346 783 350
rect 787 346 788 350
rect 782 345 788 346
rect 862 350 868 351
rect 862 346 863 350
rect 867 346 868 350
rect 862 345 868 346
rect 942 350 948 351
rect 942 346 943 350
rect 947 346 948 350
rect 942 345 948 346
rect 1022 350 1028 351
rect 1022 346 1023 350
rect 1027 346 1028 350
rect 1022 345 1028 346
rect 1102 350 1108 351
rect 1102 346 1103 350
rect 1107 346 1108 350
rect 1102 345 1108 346
rect 1190 350 1196 351
rect 1190 346 1191 350
rect 1195 346 1196 350
rect 1190 345 1196 346
rect 1278 350 1284 351
rect 1278 346 1279 350
rect 1283 346 1284 350
rect 1670 350 1671 354
rect 1675 350 1676 354
rect 1670 349 1676 350
rect 1726 354 1732 355
rect 1726 350 1727 354
rect 1731 350 1732 354
rect 1726 349 1732 350
rect 1782 354 1788 355
rect 1782 350 1783 354
rect 1787 350 1788 354
rect 1782 349 1788 350
rect 1838 354 1844 355
rect 1838 350 1839 354
rect 1843 350 1844 354
rect 1838 349 1844 350
rect 1894 354 1900 355
rect 1894 350 1895 354
rect 1899 350 1900 354
rect 1894 349 1900 350
rect 1966 354 1972 355
rect 1966 350 1967 354
rect 1971 350 1972 354
rect 1966 349 1972 350
rect 2054 354 2060 355
rect 2054 350 2055 354
rect 2059 350 2060 354
rect 2054 349 2060 350
rect 2166 354 2172 355
rect 2166 350 2167 354
rect 2171 350 2172 354
rect 2166 349 2172 350
rect 2294 354 2300 355
rect 2294 350 2295 354
rect 2299 350 2300 354
rect 2294 349 2300 350
rect 2430 354 2436 355
rect 2430 350 2431 354
rect 2435 350 2436 354
rect 2430 349 2436 350
rect 2542 354 2548 355
rect 2542 350 2543 354
rect 2547 350 2548 354
rect 2542 349 2548 350
rect 1278 345 1284 346
rect 1647 347 1653 348
rect 407 343 413 344
rect 407 339 408 343
rect 412 342 413 343
rect 454 343 460 344
rect 454 342 455 343
rect 412 340 455 342
rect 412 339 413 340
rect 407 338 413 339
rect 454 339 455 340
rect 459 339 460 343
rect 454 338 460 339
rect 462 343 469 344
rect 462 339 463 343
rect 468 339 469 343
rect 462 338 469 339
rect 526 343 533 344
rect 526 339 527 343
rect 532 339 533 343
rect 526 338 533 339
rect 598 343 605 344
rect 598 339 599 343
rect 604 339 605 343
rect 598 338 605 339
rect 678 343 685 344
rect 678 339 679 343
rect 684 339 685 343
rect 678 338 685 339
rect 759 343 765 344
rect 759 339 760 343
rect 764 342 765 343
rect 807 343 813 344
rect 807 342 808 343
rect 764 340 808 342
rect 764 339 765 340
rect 759 338 765 339
rect 807 339 808 340
rect 812 339 813 343
rect 807 338 813 339
rect 839 343 845 344
rect 839 339 840 343
rect 844 342 845 343
rect 854 343 860 344
rect 854 342 855 343
rect 844 340 855 342
rect 844 339 845 340
rect 839 338 845 339
rect 854 339 855 340
rect 859 339 860 343
rect 854 338 860 339
rect 919 343 925 344
rect 919 339 920 343
rect 924 342 925 343
rect 934 343 940 344
rect 934 342 935 343
rect 924 340 935 342
rect 924 339 925 340
rect 919 338 925 339
rect 934 339 935 340
rect 939 339 940 343
rect 934 338 940 339
rect 998 343 1005 344
rect 998 339 999 343
rect 1004 339 1005 343
rect 998 338 1005 339
rect 1079 343 1085 344
rect 1079 339 1080 343
rect 1084 342 1085 343
rect 1127 343 1133 344
rect 1127 342 1128 343
rect 1084 340 1128 342
rect 1084 339 1085 340
rect 1079 338 1085 339
rect 1127 339 1128 340
rect 1132 339 1133 343
rect 1127 338 1133 339
rect 1167 343 1173 344
rect 1167 339 1168 343
rect 1172 342 1173 343
rect 1215 343 1221 344
rect 1215 342 1216 343
rect 1172 340 1216 342
rect 1172 339 1173 340
rect 1167 338 1173 339
rect 1215 339 1216 340
rect 1220 339 1221 343
rect 1215 338 1221 339
rect 1254 343 1261 344
rect 1254 339 1255 343
rect 1260 339 1261 343
rect 1647 343 1648 347
rect 1652 343 1653 347
rect 1647 342 1653 343
rect 1702 347 1709 348
rect 1702 343 1703 347
rect 1708 343 1709 347
rect 1702 342 1709 343
rect 1758 347 1765 348
rect 1758 343 1759 347
rect 1764 343 1765 347
rect 1758 342 1765 343
rect 1814 347 1821 348
rect 1814 343 1815 347
rect 1820 343 1821 347
rect 1814 342 1821 343
rect 1870 347 1877 348
rect 1870 343 1871 347
rect 1876 343 1877 347
rect 1870 342 1877 343
rect 1942 347 1949 348
rect 1942 343 1943 347
rect 1948 343 1949 347
rect 1942 342 1949 343
rect 2018 347 2024 348
rect 2018 343 2019 347
rect 2023 346 2024 347
rect 2031 347 2037 348
rect 2031 346 2032 347
rect 2023 344 2032 346
rect 2023 343 2024 344
rect 2018 342 2024 343
rect 2031 343 2032 344
rect 2036 343 2037 347
rect 2031 342 2037 343
rect 2142 347 2149 348
rect 2142 343 2143 347
rect 2148 343 2149 347
rect 2142 342 2149 343
rect 2270 347 2277 348
rect 2270 343 2271 347
rect 2276 343 2277 347
rect 2270 342 2277 343
rect 2406 347 2413 348
rect 2406 343 2407 347
rect 2412 343 2413 347
rect 2406 342 2413 343
rect 2519 347 2525 348
rect 2519 343 2520 347
rect 2524 346 2525 347
rect 2558 347 2564 348
rect 2558 346 2559 347
rect 2524 344 2559 346
rect 2524 343 2525 344
rect 2519 342 2525 343
rect 2558 343 2559 344
rect 2563 343 2564 347
rect 2558 342 2564 343
rect 1254 338 1261 339
rect 1649 338 1651 342
rect 1982 339 1988 340
rect 1982 338 1983 339
rect 1649 336 1983 338
rect 710 335 716 336
rect 710 334 711 335
rect 568 332 711 334
rect 438 327 445 328
rect 438 323 439 327
rect 444 323 445 327
rect 495 327 501 328
rect 495 323 496 327
rect 500 326 501 327
rect 510 327 516 328
rect 510 326 511 327
rect 500 324 511 326
rect 500 323 501 324
rect 438 322 445 323
rect 462 322 468 323
rect 495 322 501 323
rect 510 323 511 324
rect 515 323 516 327
rect 551 327 557 328
rect 551 323 552 327
rect 556 326 557 327
rect 568 326 570 332
rect 710 331 711 332
rect 715 331 716 335
rect 934 335 940 336
rect 934 334 935 335
rect 710 330 716 331
rect 760 332 935 334
rect 556 324 570 326
rect 594 327 600 328
rect 556 323 557 324
rect 594 323 595 327
rect 599 326 600 327
rect 607 327 613 328
rect 607 326 608 327
rect 599 324 608 326
rect 599 323 600 324
rect 510 322 516 323
rect 518 322 524 323
rect 551 322 557 323
rect 574 322 580 323
rect 594 322 600 323
rect 607 323 608 324
rect 612 323 613 327
rect 650 327 656 328
rect 650 323 651 327
rect 655 326 656 327
rect 671 327 677 328
rect 671 326 672 327
rect 655 324 672 326
rect 655 323 656 324
rect 607 322 613 323
rect 630 322 636 323
rect 650 322 656 323
rect 671 323 672 324
rect 676 323 677 327
rect 743 327 749 328
rect 743 323 744 327
rect 748 326 749 327
rect 760 326 762 332
rect 934 331 935 332
rect 939 331 940 335
rect 1982 335 1983 336
rect 1987 335 1988 339
rect 1982 334 1988 335
rect 934 330 940 331
rect 748 324 762 326
rect 791 327 797 328
rect 748 323 749 324
rect 791 323 792 327
rect 796 326 797 327
rect 823 327 829 328
rect 823 326 824 327
rect 796 324 824 326
rect 796 323 797 324
rect 671 322 677 323
rect 694 322 700 323
rect 743 322 749 323
rect 766 322 772 323
rect 791 322 797 323
rect 823 323 824 324
rect 828 323 829 327
rect 902 327 909 328
rect 902 323 903 327
rect 908 323 909 327
rect 962 327 968 328
rect 962 323 963 327
rect 967 326 968 327
rect 991 327 997 328
rect 991 326 992 327
rect 967 324 992 326
rect 967 323 968 324
rect 823 322 829 323
rect 846 322 852 323
rect 902 322 909 323
rect 926 322 932 323
rect 962 322 968 323
rect 991 323 992 324
rect 996 323 997 327
rect 1078 327 1084 328
rect 1078 323 1079 327
rect 1083 326 1084 327
rect 1087 327 1093 328
rect 1087 326 1088 327
rect 1083 324 1088 326
rect 1083 323 1084 324
rect 991 322 997 323
rect 1014 322 1020 323
rect 1078 322 1084 323
rect 1087 323 1088 324
rect 1092 323 1093 327
rect 1130 327 1136 328
rect 1130 323 1131 327
rect 1135 326 1136 327
rect 1191 327 1197 328
rect 1191 326 1192 327
rect 1135 324 1192 326
rect 1135 323 1136 324
rect 1087 322 1093 323
rect 1110 322 1116 323
rect 1130 322 1136 323
rect 1191 323 1192 324
rect 1196 323 1197 327
rect 1607 327 1613 328
rect 1607 323 1608 327
rect 1612 326 1613 327
rect 1622 327 1628 328
rect 1622 326 1623 327
rect 1612 324 1623 326
rect 1612 323 1613 324
rect 1191 322 1197 323
rect 1214 322 1220 323
rect 1607 322 1613 323
rect 1622 323 1623 324
rect 1627 323 1628 327
rect 1650 327 1656 328
rect 1650 323 1651 327
rect 1655 326 1656 327
rect 1663 327 1669 328
rect 1663 326 1664 327
rect 1655 324 1664 326
rect 1655 323 1656 324
rect 1622 322 1628 323
rect 1630 322 1636 323
rect 1650 322 1656 323
rect 1663 323 1664 324
rect 1668 323 1669 327
rect 1706 327 1712 328
rect 1706 323 1707 327
rect 1711 326 1712 327
rect 1719 327 1725 328
rect 1719 326 1720 327
rect 1711 324 1720 326
rect 1711 323 1712 324
rect 1663 322 1669 323
rect 1686 322 1692 323
rect 1706 322 1712 323
rect 1719 323 1720 324
rect 1724 323 1725 327
rect 1762 327 1768 328
rect 1762 323 1763 327
rect 1767 326 1768 327
rect 1783 327 1789 328
rect 1783 326 1784 327
rect 1767 324 1784 326
rect 1767 323 1768 324
rect 1719 322 1725 323
rect 1742 322 1748 323
rect 1762 322 1768 323
rect 1783 323 1784 324
rect 1788 323 1789 327
rect 1826 327 1832 328
rect 1826 323 1827 327
rect 1831 326 1832 327
rect 1863 327 1869 328
rect 1863 326 1864 327
rect 1831 324 1864 326
rect 1831 323 1832 324
rect 1783 322 1789 323
rect 1806 322 1812 323
rect 1826 322 1832 323
rect 1863 323 1864 324
rect 1868 323 1869 327
rect 1906 327 1912 328
rect 1906 323 1907 327
rect 1911 326 1912 327
rect 1943 327 1949 328
rect 1943 326 1944 327
rect 1911 324 1944 326
rect 1911 323 1912 324
rect 1863 322 1869 323
rect 1886 322 1892 323
rect 1906 322 1912 323
rect 1943 323 1944 324
rect 1948 323 1949 327
rect 2030 327 2037 328
rect 2030 323 2031 327
rect 2036 323 2037 327
rect 2119 327 2128 328
rect 2119 323 2120 327
rect 2127 323 2128 327
rect 2207 327 2213 328
rect 2207 323 2208 327
rect 2212 326 2213 327
rect 2222 327 2228 328
rect 2222 326 2223 327
rect 2212 324 2223 326
rect 2212 323 2213 324
rect 1943 322 1949 323
rect 1966 322 1972 323
rect 2030 322 2037 323
rect 2054 322 2060 323
rect 2119 322 2128 323
rect 2142 322 2148 323
rect 2207 322 2213 323
rect 2222 323 2223 324
rect 2227 323 2228 327
rect 2250 327 2256 328
rect 2250 323 2251 327
rect 2255 326 2256 327
rect 2287 327 2293 328
rect 2287 326 2288 327
rect 2255 324 2288 326
rect 2255 323 2256 324
rect 2222 322 2228 323
rect 2230 322 2236 323
rect 2250 322 2256 323
rect 2287 323 2288 324
rect 2292 323 2293 327
rect 2330 327 2336 328
rect 2330 323 2331 327
rect 2335 326 2336 327
rect 2367 327 2373 328
rect 2367 326 2368 327
rect 2335 324 2368 326
rect 2335 323 2336 324
rect 2287 322 2293 323
rect 2310 322 2316 323
rect 2330 322 2336 323
rect 2367 323 2368 324
rect 2372 323 2373 327
rect 2454 327 2461 328
rect 2454 323 2455 327
rect 2460 323 2461 327
rect 2498 327 2504 328
rect 2498 323 2499 327
rect 2503 326 2504 327
rect 2519 327 2525 328
rect 2519 326 2520 327
rect 2503 324 2520 326
rect 2503 323 2504 324
rect 2367 322 2373 323
rect 2390 322 2396 323
rect 2454 322 2461 323
rect 2478 322 2484 323
rect 2498 322 2504 323
rect 2519 323 2520 324
rect 2524 323 2525 327
rect 2519 322 2525 323
rect 2542 322 2548 323
rect 462 318 463 322
rect 467 318 468 322
rect 462 317 468 318
rect 518 318 519 322
rect 523 318 524 322
rect 518 317 524 318
rect 574 318 575 322
rect 579 318 580 322
rect 574 317 580 318
rect 630 318 631 322
rect 635 318 636 322
rect 630 317 636 318
rect 694 318 695 322
rect 699 318 700 322
rect 694 317 700 318
rect 766 318 767 322
rect 771 318 772 322
rect 766 317 772 318
rect 846 318 847 322
rect 851 318 852 322
rect 846 317 852 318
rect 926 318 927 322
rect 931 318 932 322
rect 926 317 932 318
rect 1014 318 1015 322
rect 1019 318 1020 322
rect 1014 317 1020 318
rect 1110 318 1111 322
rect 1115 318 1116 322
rect 1110 317 1116 318
rect 1214 318 1215 322
rect 1219 318 1220 322
rect 1214 317 1220 318
rect 1630 318 1631 322
rect 1635 318 1636 322
rect 1630 317 1636 318
rect 1686 318 1687 322
rect 1691 318 1692 322
rect 1686 317 1692 318
rect 1742 318 1743 322
rect 1747 318 1748 322
rect 1742 317 1748 318
rect 1806 318 1807 322
rect 1811 318 1812 322
rect 1806 317 1812 318
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1966 318 1967 322
rect 1971 318 1972 322
rect 1966 317 1972 318
rect 2054 318 2055 322
rect 2059 318 2060 322
rect 2054 317 2060 318
rect 2142 318 2143 322
rect 2147 318 2148 322
rect 2142 317 2148 318
rect 2230 318 2231 322
rect 2235 318 2236 322
rect 2230 317 2236 318
rect 2310 318 2311 322
rect 2315 318 2316 322
rect 2310 317 2316 318
rect 2390 318 2391 322
rect 2395 318 2396 322
rect 2390 317 2396 318
rect 2478 318 2479 322
rect 2483 318 2484 322
rect 2478 317 2484 318
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1326 308 1332 309
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 438 303 444 304
rect 438 299 439 303
rect 443 302 444 303
rect 902 303 908 304
rect 443 300 530 302
rect 443 299 444 300
rect 438 298 444 299
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 446 295 452 296
rect 446 291 447 295
rect 451 291 452 295
rect 502 295 508 296
rect 446 290 452 291
rect 479 291 485 292
rect 479 290 480 291
rect 456 288 480 290
rect 454 287 460 288
rect 454 283 455 287
rect 459 283 460 287
rect 479 287 480 288
rect 484 287 485 291
rect 502 291 503 295
rect 507 291 508 295
rect 502 290 508 291
rect 528 290 530 300
rect 902 299 903 303
rect 907 302 908 303
rect 2030 303 2036 304
rect 907 300 1026 302
rect 907 299 908 300
rect 902 298 908 299
rect 558 295 564 296
rect 535 291 541 292
rect 535 290 536 291
rect 528 288 536 290
rect 479 286 485 287
rect 535 287 536 288
rect 540 287 541 291
rect 558 291 559 295
rect 563 291 564 295
rect 614 295 620 296
rect 558 290 564 291
rect 591 291 600 292
rect 535 286 541 287
rect 591 287 592 291
rect 599 287 600 291
rect 614 291 615 295
rect 619 291 620 295
rect 678 295 684 296
rect 614 290 620 291
rect 647 291 656 292
rect 591 286 600 287
rect 647 287 648 291
rect 655 287 656 291
rect 678 291 679 295
rect 683 291 684 295
rect 750 295 756 296
rect 678 290 684 291
rect 710 291 717 292
rect 647 286 656 287
rect 710 287 711 291
rect 716 287 717 291
rect 750 291 751 295
rect 755 291 756 295
rect 791 295 797 296
rect 791 294 792 295
rect 750 290 756 291
rect 783 293 792 294
rect 783 289 784 293
rect 788 292 792 293
rect 788 289 789 292
rect 791 291 792 292
rect 796 291 797 295
rect 791 290 797 291
rect 830 295 836 296
rect 830 291 831 295
rect 835 291 836 295
rect 910 295 916 296
rect 830 290 836 291
rect 854 291 860 292
rect 783 288 789 289
rect 710 286 717 287
rect 854 287 855 291
rect 859 290 860 291
rect 863 291 869 292
rect 863 290 864 291
rect 859 288 864 290
rect 859 287 860 288
rect 854 286 860 287
rect 863 287 864 288
rect 868 287 869 291
rect 910 291 911 295
rect 915 291 916 295
rect 998 295 1004 296
rect 910 290 916 291
rect 934 291 940 292
rect 863 286 869 287
rect 934 287 935 291
rect 939 290 940 291
rect 943 291 949 292
rect 943 290 944 291
rect 939 288 944 290
rect 939 287 940 288
rect 934 286 940 287
rect 943 287 944 288
rect 948 287 949 291
rect 998 291 999 295
rect 1003 291 1004 295
rect 998 290 1004 291
rect 1024 290 1026 300
rect 2030 299 2031 303
rect 2035 302 2036 303
rect 2035 300 2154 302
rect 2035 299 2036 300
rect 2030 298 2036 299
rect 1326 296 1332 297
rect 1094 295 1100 296
rect 1031 291 1037 292
rect 1031 290 1032 291
rect 1024 288 1032 290
rect 943 286 949 287
rect 1031 287 1032 288
rect 1036 287 1037 291
rect 1094 291 1095 295
rect 1099 291 1100 295
rect 1198 295 1204 296
rect 1094 290 1100 291
rect 1127 291 1136 292
rect 1031 286 1037 287
rect 1127 287 1128 291
rect 1135 287 1136 291
rect 1198 291 1199 295
rect 1203 291 1204 295
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1198 290 1204 291
rect 1222 291 1228 292
rect 1127 286 1136 287
rect 1222 287 1223 291
rect 1227 290 1228 291
rect 1231 291 1237 292
rect 1326 291 1332 292
rect 1366 296 1372 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1614 295 1620 296
rect 1614 291 1615 295
rect 1619 291 1620 295
rect 1670 295 1676 296
rect 1231 290 1232 291
rect 1227 288 1232 290
rect 1227 287 1228 288
rect 1222 286 1228 287
rect 1231 287 1232 288
rect 1236 287 1237 291
rect 1614 290 1620 291
rect 1647 291 1656 292
rect 1231 286 1237 287
rect 1647 287 1648 291
rect 1655 287 1656 291
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1726 295 1732 296
rect 1670 290 1676 291
rect 1703 291 1712 292
rect 1647 286 1656 287
rect 1703 287 1704 291
rect 1711 287 1712 291
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1790 295 1796 296
rect 1726 290 1732 291
rect 1759 291 1768 292
rect 1703 286 1712 287
rect 1759 287 1760 291
rect 1767 287 1768 291
rect 1790 291 1791 295
rect 1795 291 1796 295
rect 1870 295 1876 296
rect 1790 290 1796 291
rect 1823 291 1832 292
rect 1759 286 1768 287
rect 1823 287 1824 291
rect 1831 287 1832 291
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1950 295 1956 296
rect 1870 290 1876 291
rect 1903 291 1912 292
rect 1823 286 1832 287
rect 1903 287 1904 291
rect 1911 287 1912 291
rect 1950 291 1951 295
rect 1955 291 1956 295
rect 2038 295 2044 296
rect 1950 290 1956 291
rect 1982 291 1989 292
rect 1903 286 1912 287
rect 1982 287 1983 291
rect 1988 287 1989 291
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2126 295 2132 296
rect 2038 290 2044 291
rect 2071 291 2077 292
rect 2071 290 2072 291
rect 2048 288 2072 290
rect 1982 286 1989 287
rect 1991 287 1997 288
rect 454 282 460 283
rect 1991 283 1992 287
rect 1996 286 1997 287
rect 2048 286 2050 288
rect 2071 287 2072 288
rect 2076 287 2077 291
rect 2126 291 2127 295
rect 2131 291 2132 295
rect 2126 290 2132 291
rect 2152 290 2154 300
rect 2582 296 2588 297
rect 2214 295 2220 296
rect 2159 291 2165 292
rect 2159 290 2160 291
rect 2152 288 2160 290
rect 2071 286 2077 287
rect 2159 287 2160 288
rect 2164 287 2165 291
rect 2214 291 2215 295
rect 2219 291 2220 295
rect 2294 295 2300 296
rect 2214 290 2220 291
rect 2247 291 2256 292
rect 2159 286 2165 287
rect 2247 287 2248 291
rect 2255 287 2256 291
rect 2294 291 2295 295
rect 2299 291 2300 295
rect 2374 295 2380 296
rect 2294 290 2300 291
rect 2327 291 2336 292
rect 2247 286 2256 287
rect 2327 287 2328 291
rect 2335 287 2336 291
rect 2374 291 2375 295
rect 2379 291 2380 295
rect 2462 295 2468 296
rect 2374 290 2380 291
rect 2398 291 2404 292
rect 2327 286 2336 287
rect 2398 287 2399 291
rect 2403 290 2404 291
rect 2407 291 2413 292
rect 2407 290 2408 291
rect 2403 288 2408 290
rect 2403 287 2404 288
rect 2398 286 2404 287
rect 2407 287 2408 288
rect 2412 287 2413 291
rect 2462 291 2463 295
rect 2467 291 2468 295
rect 2526 295 2532 296
rect 2462 290 2468 291
rect 2495 291 2504 292
rect 2407 286 2413 287
rect 2495 287 2496 291
rect 2503 287 2504 291
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2526 290 2532 291
rect 2558 291 2565 292
rect 2582 291 2588 292
rect 2495 286 2504 287
rect 2558 287 2559 291
rect 2564 287 2565 291
rect 2558 286 2565 287
rect 1996 284 2050 286
rect 1996 283 1997 284
rect 1991 282 1997 283
rect 1622 271 1628 272
rect 510 267 516 268
rect 510 263 511 267
rect 515 266 516 267
rect 846 267 852 268
rect 515 264 650 266
rect 515 263 516 264
rect 510 262 516 263
rect 319 259 325 260
rect 286 257 292 258
rect 110 256 116 257
rect 110 252 111 256
rect 115 252 116 256
rect 286 253 287 257
rect 291 253 292 257
rect 319 255 320 259
rect 324 258 325 259
rect 342 259 348 260
rect 342 258 343 259
rect 324 256 343 258
rect 324 255 325 256
rect 319 254 325 255
rect 342 255 343 256
rect 347 255 348 259
rect 391 259 397 260
rect 342 254 348 255
rect 358 257 364 258
rect 286 252 292 253
rect 358 253 359 257
rect 363 253 364 257
rect 391 255 392 259
rect 396 258 397 259
rect 430 259 436 260
rect 430 258 431 259
rect 396 256 431 258
rect 396 255 397 256
rect 391 254 397 255
rect 430 255 431 256
rect 435 255 436 259
rect 471 259 477 260
rect 430 254 436 255
rect 438 257 444 258
rect 358 252 364 253
rect 438 253 439 257
rect 443 253 444 257
rect 471 255 472 259
rect 476 258 477 259
rect 518 259 524 260
rect 518 258 519 259
rect 476 256 519 258
rect 476 255 477 256
rect 471 254 477 255
rect 518 255 519 256
rect 523 255 524 259
rect 559 259 565 260
rect 518 254 524 255
rect 526 257 532 258
rect 438 252 444 253
rect 526 253 527 257
rect 531 253 532 257
rect 559 255 560 259
rect 564 258 565 259
rect 614 259 620 260
rect 614 258 615 259
rect 564 256 615 258
rect 564 255 565 256
rect 559 254 565 255
rect 614 255 615 256
rect 619 255 620 259
rect 648 258 650 264
rect 846 263 847 267
rect 851 266 852 267
rect 1622 267 1623 271
rect 1627 270 1628 271
rect 2222 271 2228 272
rect 1627 268 1890 270
rect 1627 267 1628 268
rect 1622 266 1628 267
rect 851 264 1058 266
rect 851 263 852 264
rect 846 262 852 263
rect 655 259 661 260
rect 655 258 656 259
rect 614 254 620 255
rect 622 257 628 258
rect 526 252 532 253
rect 622 253 623 257
rect 627 253 628 257
rect 648 256 656 258
rect 655 255 656 256
rect 660 255 661 259
rect 751 259 757 260
rect 655 254 661 255
rect 718 257 724 258
rect 622 252 628 253
rect 718 253 719 257
rect 723 253 724 257
rect 751 255 752 259
rect 756 258 757 259
rect 766 259 772 260
rect 766 258 767 259
rect 756 256 767 258
rect 756 255 757 256
rect 751 254 757 255
rect 766 255 767 256
rect 771 255 772 259
rect 855 259 861 260
rect 766 254 772 255
rect 822 257 828 258
rect 718 252 724 253
rect 822 253 823 257
rect 827 253 828 257
rect 855 255 856 259
rect 860 258 861 259
rect 918 259 924 260
rect 918 258 919 259
rect 860 256 919 258
rect 860 255 861 256
rect 855 254 861 255
rect 918 255 919 256
rect 923 255 924 259
rect 959 259 968 260
rect 918 254 924 255
rect 926 257 932 258
rect 822 252 828 253
rect 926 253 927 257
rect 931 253 932 257
rect 959 255 960 259
rect 967 255 968 259
rect 1056 258 1058 264
rect 1567 263 1573 264
rect 1534 261 1540 262
rect 1366 260 1372 261
rect 1063 259 1069 260
rect 1063 258 1064 259
rect 959 254 968 255
rect 1030 257 1036 258
rect 926 252 932 253
rect 1030 253 1031 257
rect 1035 253 1036 257
rect 1056 256 1064 258
rect 1063 255 1064 256
rect 1068 255 1069 259
rect 1175 259 1181 260
rect 1063 254 1069 255
rect 1142 257 1148 258
rect 1030 252 1036 253
rect 1142 253 1143 257
rect 1147 253 1148 257
rect 1175 255 1176 259
rect 1180 258 1181 259
rect 1246 259 1252 260
rect 1246 258 1247 259
rect 1180 256 1247 258
rect 1180 255 1181 256
rect 1175 254 1181 255
rect 1246 255 1247 256
rect 1251 255 1252 259
rect 1278 259 1284 260
rect 1246 254 1252 255
rect 1254 257 1260 258
rect 1142 252 1148 253
rect 1254 253 1255 257
rect 1259 253 1260 257
rect 1278 255 1279 259
rect 1283 258 1284 259
rect 1287 259 1293 260
rect 1287 258 1288 259
rect 1283 256 1288 258
rect 1283 255 1284 256
rect 1278 254 1284 255
rect 1287 255 1288 256
rect 1292 255 1293 259
rect 1287 254 1293 255
rect 1326 256 1332 257
rect 1254 252 1260 253
rect 1326 252 1327 256
rect 1331 252 1332 256
rect 1366 256 1367 260
rect 1371 256 1372 260
rect 1534 257 1535 261
rect 1539 257 1540 261
rect 1567 259 1568 263
rect 1572 262 1573 263
rect 1598 263 1604 264
rect 1598 262 1599 263
rect 1572 260 1599 262
rect 1572 259 1573 260
rect 1567 258 1573 259
rect 1598 259 1599 260
rect 1603 259 1604 263
rect 1639 263 1645 264
rect 1598 258 1604 259
rect 1606 261 1612 262
rect 1534 256 1540 257
rect 1606 257 1607 261
rect 1611 257 1612 261
rect 1639 259 1640 263
rect 1644 262 1645 263
rect 1678 263 1684 264
rect 1678 262 1679 263
rect 1644 260 1679 262
rect 1644 259 1645 260
rect 1639 258 1645 259
rect 1678 259 1679 260
rect 1683 259 1684 263
rect 1719 263 1725 264
rect 1678 258 1684 259
rect 1686 261 1692 262
rect 1606 256 1612 257
rect 1686 257 1687 261
rect 1691 257 1692 261
rect 1719 259 1720 263
rect 1724 262 1725 263
rect 1766 263 1772 264
rect 1766 262 1767 263
rect 1724 260 1767 262
rect 1724 259 1725 260
rect 1719 258 1725 259
rect 1766 259 1767 260
rect 1771 259 1772 263
rect 1807 263 1813 264
rect 1766 258 1772 259
rect 1774 261 1780 262
rect 1686 256 1692 257
rect 1774 257 1775 261
rect 1779 257 1780 261
rect 1807 259 1808 263
rect 1812 262 1813 263
rect 1846 263 1852 264
rect 1846 262 1847 263
rect 1812 260 1847 262
rect 1812 259 1813 260
rect 1807 258 1813 259
rect 1846 259 1847 260
rect 1851 259 1852 263
rect 1888 262 1890 268
rect 2222 267 2223 271
rect 2227 270 2228 271
rect 2454 271 2460 272
rect 2227 268 2371 270
rect 2227 267 2228 268
rect 2222 266 2228 267
rect 2369 264 2371 268
rect 2454 267 2455 271
rect 2459 270 2460 271
rect 2459 268 2554 270
rect 2459 267 2460 268
rect 2454 266 2460 267
rect 1895 263 1901 264
rect 1895 262 1896 263
rect 1846 258 1852 259
rect 1862 261 1868 262
rect 1774 256 1780 257
rect 1862 257 1863 261
rect 1867 257 1868 261
rect 1888 260 1896 262
rect 1895 259 1896 260
rect 1900 259 1901 263
rect 1983 263 1989 264
rect 1895 258 1901 259
rect 1950 261 1956 262
rect 1862 256 1868 257
rect 1950 257 1951 261
rect 1955 257 1956 261
rect 1983 259 1984 263
rect 1988 262 1989 263
rect 2030 263 2036 264
rect 2030 262 2031 263
rect 1988 260 2031 262
rect 1988 259 1989 260
rect 1983 258 1989 259
rect 2030 259 2031 260
rect 2035 259 2036 263
rect 2070 263 2077 264
rect 2030 258 2036 259
rect 2038 261 2044 262
rect 1950 256 1956 257
rect 2038 257 2039 261
rect 2043 257 2044 261
rect 2070 259 2071 263
rect 2076 259 2077 263
rect 2151 263 2157 264
rect 2070 258 2077 259
rect 2118 261 2124 262
rect 2038 256 2044 257
rect 2118 257 2119 261
rect 2123 257 2124 261
rect 2151 259 2152 263
rect 2156 262 2157 263
rect 2190 263 2196 264
rect 2190 262 2191 263
rect 2156 260 2191 262
rect 2156 259 2157 260
rect 2151 258 2157 259
rect 2190 259 2191 260
rect 2195 259 2196 263
rect 2231 263 2237 264
rect 2190 258 2196 259
rect 2198 261 2204 262
rect 2118 256 2124 257
rect 2198 257 2199 261
rect 2203 257 2204 261
rect 2231 259 2232 263
rect 2236 262 2237 263
rect 2254 263 2260 264
rect 2254 262 2255 263
rect 2236 260 2255 262
rect 2236 259 2237 260
rect 2231 258 2237 259
rect 2254 259 2255 260
rect 2259 259 2260 263
rect 2303 263 2309 264
rect 2254 258 2260 259
rect 2270 261 2276 262
rect 2198 256 2204 257
rect 2270 257 2271 261
rect 2275 257 2276 261
rect 2303 259 2304 263
rect 2308 262 2309 263
rect 2326 263 2332 264
rect 2326 262 2327 263
rect 2308 260 2327 262
rect 2308 259 2309 260
rect 2303 258 2309 259
rect 2326 259 2327 260
rect 2331 259 2332 263
rect 2367 263 2373 264
rect 2326 258 2332 259
rect 2334 261 2340 262
rect 2270 256 2276 257
rect 2334 257 2335 261
rect 2339 257 2340 261
rect 2367 259 2368 263
rect 2372 259 2373 263
rect 2439 263 2445 264
rect 2367 258 2373 259
rect 2406 261 2412 262
rect 2334 256 2340 257
rect 2406 257 2407 261
rect 2411 257 2412 261
rect 2439 259 2440 263
rect 2444 262 2445 263
rect 2455 263 2461 264
rect 2455 262 2456 263
rect 2444 260 2456 262
rect 2444 259 2445 260
rect 2439 258 2445 259
rect 2455 259 2456 260
rect 2460 259 2461 263
rect 2494 263 2500 264
rect 2455 258 2461 259
rect 2470 261 2476 262
rect 2406 256 2412 257
rect 2470 257 2471 261
rect 2475 257 2476 261
rect 2494 259 2495 263
rect 2499 262 2500 263
rect 2503 263 2509 264
rect 2503 262 2504 263
rect 2499 260 2504 262
rect 2499 259 2500 260
rect 2494 258 2500 259
rect 2503 259 2504 260
rect 2508 259 2509 263
rect 2552 262 2554 268
rect 2559 263 2565 264
rect 2559 262 2560 263
rect 2503 258 2509 259
rect 2526 261 2532 262
rect 2470 256 2476 257
rect 2526 257 2527 261
rect 2531 257 2532 261
rect 2552 260 2560 262
rect 2559 259 2560 260
rect 2564 259 2565 263
rect 2559 258 2565 259
rect 2582 260 2588 261
rect 2526 256 2532 257
rect 2582 256 2583 260
rect 2587 256 2588 260
rect 1366 255 1372 256
rect 2582 255 2588 256
rect 110 251 116 252
rect 1326 251 1332 252
rect 1366 243 1372 244
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1366 239 1367 243
rect 1371 239 1372 243
rect 1366 238 1372 239
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 1326 234 1332 235
rect 1550 234 1556 235
rect 302 230 308 231
rect 302 226 303 230
rect 307 226 308 230
rect 302 225 308 226
rect 374 230 380 231
rect 374 226 375 230
rect 379 226 380 230
rect 374 225 380 226
rect 454 230 460 231
rect 454 226 455 230
rect 459 226 460 230
rect 454 225 460 226
rect 542 230 548 231
rect 542 226 543 230
rect 547 226 548 230
rect 542 225 548 226
rect 638 230 644 231
rect 638 226 639 230
rect 643 226 644 230
rect 638 225 644 226
rect 734 230 740 231
rect 734 226 735 230
rect 739 226 740 230
rect 734 225 740 226
rect 838 230 844 231
rect 838 226 839 230
rect 843 226 844 230
rect 838 225 844 226
rect 942 230 948 231
rect 942 226 943 230
rect 947 226 948 230
rect 942 225 948 226
rect 1046 230 1052 231
rect 1046 226 1047 230
rect 1051 226 1052 230
rect 1046 225 1052 226
rect 1158 230 1164 231
rect 1158 226 1159 230
rect 1163 226 1164 230
rect 1158 225 1164 226
rect 1270 230 1276 231
rect 1270 226 1271 230
rect 1275 226 1276 230
rect 1550 230 1551 234
rect 1555 230 1556 234
rect 1550 229 1556 230
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1702 234 1708 235
rect 1702 230 1703 234
rect 1707 230 1708 234
rect 1702 229 1708 230
rect 1790 234 1796 235
rect 1790 230 1791 234
rect 1795 230 1796 234
rect 1790 229 1796 230
rect 1878 234 1884 235
rect 1878 230 1879 234
rect 1883 230 1884 234
rect 1878 229 1884 230
rect 1966 234 1972 235
rect 1966 230 1967 234
rect 1971 230 1972 234
rect 1966 229 1972 230
rect 2054 234 2060 235
rect 2054 230 2055 234
rect 2059 230 2060 234
rect 2054 229 2060 230
rect 2134 234 2140 235
rect 2134 230 2135 234
rect 2139 230 2140 234
rect 2134 229 2140 230
rect 2214 234 2220 235
rect 2214 230 2215 234
rect 2219 230 2220 234
rect 2214 229 2220 230
rect 2286 234 2292 235
rect 2286 230 2287 234
rect 2291 230 2292 234
rect 2286 229 2292 230
rect 2350 234 2356 235
rect 2350 230 2351 234
rect 2355 230 2356 234
rect 2350 229 2356 230
rect 2422 234 2428 235
rect 2422 230 2423 234
rect 2427 230 2428 234
rect 2422 229 2428 230
rect 2486 234 2492 235
rect 2486 230 2487 234
rect 2491 230 2492 234
rect 2486 229 2492 230
rect 2542 234 2548 235
rect 2542 230 2543 234
rect 2547 230 2548 234
rect 2542 229 2548 230
rect 1270 225 1276 226
rect 1527 227 1533 228
rect 279 223 285 224
rect 279 219 280 223
rect 284 222 285 223
rect 334 223 340 224
rect 334 222 335 223
rect 284 220 335 222
rect 284 219 285 220
rect 279 218 285 219
rect 334 219 335 220
rect 339 219 340 223
rect 334 218 340 219
rect 342 223 348 224
rect 342 219 343 223
rect 347 222 348 223
rect 351 223 357 224
rect 351 222 352 223
rect 347 220 352 222
rect 347 219 348 220
rect 342 218 348 219
rect 351 219 352 220
rect 356 219 357 223
rect 351 218 357 219
rect 430 223 437 224
rect 430 219 431 223
rect 436 219 437 223
rect 430 218 437 219
rect 518 223 525 224
rect 518 219 519 223
rect 524 219 525 223
rect 518 218 525 219
rect 614 223 621 224
rect 614 219 615 223
rect 620 219 621 223
rect 614 218 621 219
rect 710 223 717 224
rect 710 219 711 223
rect 716 219 717 223
rect 710 218 717 219
rect 815 223 821 224
rect 815 219 816 223
rect 820 222 821 223
rect 846 223 852 224
rect 846 222 847 223
rect 820 220 847 222
rect 820 219 821 220
rect 815 218 821 219
rect 846 219 847 220
rect 851 219 852 223
rect 846 218 852 219
rect 918 223 925 224
rect 918 219 919 223
rect 924 219 925 223
rect 918 218 925 219
rect 1023 223 1029 224
rect 1023 219 1024 223
rect 1028 222 1029 223
rect 1038 223 1044 224
rect 1038 222 1039 223
rect 1028 220 1039 222
rect 1028 219 1029 220
rect 1023 218 1029 219
rect 1038 219 1039 220
rect 1043 219 1044 223
rect 1038 218 1044 219
rect 1135 223 1141 224
rect 1135 219 1136 223
rect 1140 222 1141 223
rect 1222 223 1228 224
rect 1222 222 1223 223
rect 1140 220 1223 222
rect 1140 219 1141 220
rect 1135 218 1141 219
rect 1222 219 1223 220
rect 1227 219 1228 223
rect 1222 218 1228 219
rect 1246 223 1253 224
rect 1246 219 1247 223
rect 1252 219 1253 223
rect 1527 223 1528 227
rect 1532 226 1533 227
rect 1590 227 1596 228
rect 1590 226 1591 227
rect 1532 224 1591 226
rect 1532 223 1533 224
rect 1527 222 1533 223
rect 1590 223 1591 224
rect 1595 223 1596 227
rect 1590 222 1596 223
rect 1598 227 1605 228
rect 1598 223 1599 227
rect 1604 223 1605 227
rect 1598 222 1605 223
rect 1678 227 1685 228
rect 1678 223 1679 227
rect 1684 223 1685 227
rect 1678 222 1685 223
rect 1766 227 1773 228
rect 1766 223 1767 227
rect 1772 223 1773 227
rect 1766 222 1773 223
rect 1846 227 1852 228
rect 1846 223 1847 227
rect 1851 226 1852 227
rect 1855 227 1861 228
rect 1855 226 1856 227
rect 1851 224 1856 226
rect 1851 223 1852 224
rect 1846 222 1852 223
rect 1855 223 1856 224
rect 1860 223 1861 227
rect 1855 222 1861 223
rect 1943 227 1949 228
rect 1943 223 1944 227
rect 1948 226 1949 227
rect 1991 227 1997 228
rect 1991 226 1992 227
rect 1948 224 1992 226
rect 1948 223 1949 224
rect 1943 222 1949 223
rect 1991 223 1992 224
rect 1996 223 1997 227
rect 1991 222 1997 223
rect 2030 227 2037 228
rect 2030 223 2031 227
rect 2036 223 2037 227
rect 2030 222 2037 223
rect 2111 227 2117 228
rect 2111 223 2112 227
rect 2116 226 2117 227
rect 2182 227 2188 228
rect 2182 226 2183 227
rect 2116 224 2183 226
rect 2116 223 2117 224
rect 2111 222 2117 223
rect 2182 223 2183 224
rect 2187 223 2188 227
rect 2182 222 2188 223
rect 2190 227 2197 228
rect 2190 223 2191 227
rect 2196 223 2197 227
rect 2190 222 2197 223
rect 2254 227 2260 228
rect 2254 223 2255 227
rect 2259 226 2260 227
rect 2263 227 2269 228
rect 2263 226 2264 227
rect 2259 224 2264 226
rect 2259 223 2260 224
rect 2254 222 2260 223
rect 2263 223 2264 224
rect 2268 223 2269 227
rect 2263 222 2269 223
rect 2326 227 2333 228
rect 2326 223 2327 227
rect 2332 223 2333 227
rect 2326 222 2333 223
rect 2398 227 2405 228
rect 2398 223 2399 227
rect 2404 223 2405 227
rect 2398 222 2405 223
rect 2455 227 2461 228
rect 2455 223 2456 227
rect 2460 226 2461 227
rect 2463 227 2469 228
rect 2463 226 2464 227
rect 2460 224 2464 226
rect 2460 223 2461 224
rect 2455 222 2461 223
rect 2463 223 2464 224
rect 2468 223 2469 227
rect 2519 227 2525 228
rect 2463 222 2469 223
rect 2494 223 2500 224
rect 2494 222 2495 223
rect 2472 220 2495 222
rect 1246 218 1253 219
rect 2070 219 2076 220
rect 2070 218 2071 219
rect 2048 216 2071 218
rect 1278 215 1284 216
rect 1278 214 1279 215
rect 1264 212 1279 214
rect 175 211 181 212
rect 175 207 176 211
rect 180 210 181 211
rect 190 211 196 212
rect 190 210 191 211
rect 180 208 191 210
rect 180 207 181 208
rect 175 206 181 207
rect 190 207 191 208
rect 195 207 196 211
rect 218 211 224 212
rect 218 207 219 211
rect 223 210 224 211
rect 247 211 253 212
rect 247 210 248 211
rect 223 208 248 210
rect 223 207 224 208
rect 190 206 196 207
rect 198 206 204 207
rect 218 206 224 207
rect 247 207 248 208
rect 252 207 253 211
rect 290 211 296 212
rect 290 207 291 211
rect 295 210 296 211
rect 335 211 341 212
rect 335 210 336 211
rect 295 208 336 210
rect 295 207 296 208
rect 247 206 253 207
rect 270 206 276 207
rect 290 206 296 207
rect 335 207 336 208
rect 340 207 341 211
rect 383 211 389 212
rect 383 207 384 211
rect 388 210 389 211
rect 439 211 445 212
rect 439 210 440 211
rect 388 208 440 210
rect 388 207 389 208
rect 335 206 341 207
rect 358 206 364 207
rect 383 206 389 207
rect 439 207 440 208
rect 444 207 445 211
rect 482 211 488 212
rect 482 207 483 211
rect 487 210 488 211
rect 543 211 549 212
rect 543 210 544 211
rect 487 208 544 210
rect 487 207 488 208
rect 439 206 445 207
rect 462 206 468 207
rect 482 206 488 207
rect 543 207 544 208
rect 548 207 549 211
rect 654 211 661 212
rect 654 207 655 211
rect 660 207 661 211
rect 766 211 773 212
rect 766 207 767 211
rect 772 207 773 211
rect 886 211 893 212
rect 886 207 887 211
rect 892 207 893 211
rect 930 211 936 212
rect 930 207 931 211
rect 935 210 936 211
rect 1007 211 1013 212
rect 1007 210 1008 211
rect 935 208 1008 210
rect 935 207 936 208
rect 543 206 549 207
rect 566 206 572 207
rect 654 206 661 207
rect 678 206 684 207
rect 766 206 773 207
rect 790 206 796 207
rect 886 206 893 207
rect 910 206 916 207
rect 930 206 936 207
rect 1007 207 1008 208
rect 1012 207 1013 211
rect 1114 211 1120 212
rect 1114 207 1115 211
rect 1119 210 1120 211
rect 1127 211 1133 212
rect 1127 210 1128 211
rect 1119 208 1128 210
rect 1119 207 1120 208
rect 1007 206 1013 207
rect 1030 206 1036 207
rect 1114 206 1120 207
rect 1127 207 1128 208
rect 1132 207 1133 211
rect 1247 211 1253 212
rect 1247 207 1248 211
rect 1252 210 1253 211
rect 1264 210 1266 212
rect 1278 211 1279 212
rect 1283 211 1284 215
rect 1278 210 1284 211
rect 1391 215 1397 216
rect 1391 211 1392 215
rect 1396 214 1397 215
rect 1406 215 1412 216
rect 1406 214 1407 215
rect 1396 212 1407 214
rect 1396 211 1397 212
rect 1391 210 1397 211
rect 1406 211 1407 212
rect 1411 211 1412 215
rect 1434 215 1440 216
rect 1434 211 1435 215
rect 1439 214 1440 215
rect 1455 215 1461 216
rect 1455 214 1456 215
rect 1439 212 1456 214
rect 1439 211 1440 212
rect 1406 210 1412 211
rect 1414 210 1420 211
rect 1434 210 1440 211
rect 1455 211 1456 212
rect 1460 211 1461 215
rect 1498 215 1504 216
rect 1498 211 1499 215
rect 1503 214 1504 215
rect 1535 215 1541 216
rect 1535 214 1536 215
rect 1503 212 1536 214
rect 1503 211 1504 212
rect 1455 210 1461 211
rect 1478 210 1484 211
rect 1498 210 1504 211
rect 1535 211 1536 212
rect 1540 211 1541 215
rect 1578 215 1584 216
rect 1578 211 1579 215
rect 1583 214 1584 215
rect 1631 215 1637 216
rect 1631 214 1632 215
rect 1583 212 1632 214
rect 1583 211 1584 212
rect 1535 210 1541 211
rect 1558 210 1564 211
rect 1578 210 1584 211
rect 1631 211 1632 212
rect 1636 211 1637 215
rect 1674 215 1680 216
rect 1674 211 1675 215
rect 1679 214 1680 215
rect 1727 215 1733 216
rect 1727 214 1728 215
rect 1679 212 1728 214
rect 1679 211 1680 212
rect 1631 210 1637 211
rect 1654 210 1660 211
rect 1674 210 1680 211
rect 1727 211 1728 212
rect 1732 211 1733 215
rect 1770 215 1776 216
rect 1770 211 1771 215
rect 1775 214 1776 215
rect 1831 215 1837 216
rect 1831 214 1832 215
rect 1775 212 1832 214
rect 1775 211 1776 212
rect 1727 210 1733 211
rect 1750 210 1756 211
rect 1770 210 1776 211
rect 1831 211 1832 212
rect 1836 211 1837 215
rect 1934 215 1941 216
rect 1934 211 1935 215
rect 1940 211 1941 215
rect 2039 215 2045 216
rect 2039 211 2040 215
rect 2044 214 2045 215
rect 2048 214 2050 216
rect 2070 215 2071 216
rect 2075 215 2076 219
rect 2472 218 2474 220
rect 2494 219 2495 220
rect 2499 219 2500 223
rect 2519 223 2520 227
rect 2524 226 2525 227
rect 2558 227 2564 228
rect 2558 226 2559 227
rect 2524 224 2559 226
rect 2524 223 2525 224
rect 2519 222 2525 223
rect 2558 223 2559 224
rect 2563 223 2564 227
rect 2558 222 2564 223
rect 2494 218 2500 219
rect 2457 216 2474 218
rect 2070 214 2076 215
rect 2143 215 2149 216
rect 2044 212 2050 214
rect 2044 211 2045 212
rect 2143 211 2144 215
rect 2148 214 2149 215
rect 2158 215 2164 216
rect 2158 214 2159 215
rect 2148 212 2159 214
rect 2148 211 2149 212
rect 1831 210 1837 211
rect 1854 210 1860 211
rect 1934 210 1941 211
rect 1958 210 1964 211
rect 2039 210 2045 211
rect 2062 210 2068 211
rect 2143 210 2149 211
rect 2158 211 2159 212
rect 2163 211 2164 215
rect 2238 215 2245 216
rect 2238 211 2239 215
rect 2244 211 2245 215
rect 2334 215 2341 216
rect 2334 211 2335 215
rect 2340 211 2341 215
rect 2439 215 2445 216
rect 2439 211 2440 215
rect 2444 214 2445 215
rect 2457 214 2459 216
rect 2444 212 2459 214
rect 2487 215 2493 216
rect 2444 211 2445 212
rect 2487 211 2488 215
rect 2492 214 2493 215
rect 2519 215 2525 216
rect 2519 214 2520 215
rect 2492 212 2520 214
rect 2492 211 2493 212
rect 2158 210 2164 211
rect 2166 210 2172 211
rect 2238 210 2245 211
rect 2262 210 2268 211
rect 2334 210 2341 211
rect 2358 210 2364 211
rect 2439 210 2445 211
rect 2462 210 2468 211
rect 2487 210 2493 211
rect 2519 211 2520 212
rect 2524 211 2525 215
rect 2519 210 2525 211
rect 2542 210 2548 211
rect 1252 208 1266 210
rect 1252 207 1253 208
rect 1127 206 1133 207
rect 1150 206 1156 207
rect 1247 206 1253 207
rect 1270 206 1276 207
rect 198 202 199 206
rect 203 202 204 206
rect 198 201 204 202
rect 270 202 271 206
rect 275 202 276 206
rect 270 201 276 202
rect 358 202 359 206
rect 363 202 364 206
rect 358 201 364 202
rect 462 202 463 206
rect 467 202 468 206
rect 462 201 468 202
rect 566 202 567 206
rect 571 202 572 206
rect 566 201 572 202
rect 678 202 679 206
rect 683 202 684 206
rect 678 201 684 202
rect 790 202 791 206
rect 795 202 796 206
rect 790 201 796 202
rect 910 202 911 206
rect 915 202 916 206
rect 910 201 916 202
rect 1030 202 1031 206
rect 1035 202 1036 206
rect 1030 201 1036 202
rect 1150 202 1151 206
rect 1155 202 1156 206
rect 1150 201 1156 202
rect 1270 202 1271 206
rect 1275 202 1276 206
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1414 205 1420 206
rect 1478 206 1479 210
rect 1483 206 1484 210
rect 1478 205 1484 206
rect 1558 206 1559 210
rect 1563 206 1564 210
rect 1558 205 1564 206
rect 1654 206 1655 210
rect 1659 206 1660 210
rect 1654 205 1660 206
rect 1750 206 1751 210
rect 1755 206 1756 210
rect 1750 205 1756 206
rect 1854 206 1855 210
rect 1859 206 1860 210
rect 1854 205 1860 206
rect 1958 206 1959 210
rect 1963 206 1964 210
rect 1958 205 1964 206
rect 2062 206 2063 210
rect 2067 206 2068 210
rect 2062 205 2068 206
rect 2166 206 2167 210
rect 2171 206 2172 210
rect 2166 205 2172 206
rect 2262 206 2263 210
rect 2267 206 2268 210
rect 2262 205 2268 206
rect 2358 206 2359 210
rect 2363 206 2364 210
rect 2358 205 2364 206
rect 2462 206 2463 210
rect 2467 206 2468 210
rect 2462 205 2468 206
rect 2542 206 2543 210
rect 2547 206 2548 210
rect 2542 205 2548 206
rect 1270 201 1276 202
rect 1366 201 1372 202
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1366 197 1367 201
rect 1371 197 1372 201
rect 1366 196 1372 197
rect 2582 201 2588 202
rect 2582 197 2583 201
rect 2587 197 2588 201
rect 2582 196 2588 197
rect 1326 192 1332 193
rect 1934 191 1940 192
rect 334 187 340 188
rect 334 183 335 187
rect 339 186 340 187
rect 654 187 660 188
rect 339 184 578 186
rect 339 183 340 184
rect 334 182 340 183
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 182 179 188 180
rect 182 175 183 179
rect 187 175 188 179
rect 254 179 260 180
rect 182 174 188 175
rect 215 175 224 176
rect 215 171 216 175
rect 223 171 224 175
rect 254 175 255 179
rect 259 175 260 179
rect 342 179 348 180
rect 254 174 260 175
rect 287 175 296 176
rect 215 170 224 171
rect 287 171 288 175
rect 295 171 296 175
rect 342 175 343 179
rect 347 175 348 179
rect 446 179 452 180
rect 342 174 348 175
rect 375 175 381 176
rect 287 170 296 171
rect 375 171 376 175
rect 380 174 381 175
rect 383 175 389 176
rect 383 174 384 175
rect 380 172 384 174
rect 380 171 381 172
rect 375 170 381 171
rect 383 171 384 172
rect 388 171 389 175
rect 446 175 447 179
rect 451 175 452 179
rect 550 179 556 180
rect 446 174 452 175
rect 479 175 488 176
rect 383 170 389 171
rect 479 171 480 175
rect 487 171 488 175
rect 550 175 551 179
rect 555 175 556 179
rect 550 174 556 175
rect 576 174 578 184
rect 654 183 655 187
rect 659 186 660 187
rect 886 187 892 188
rect 659 184 802 186
rect 659 183 660 184
rect 654 182 660 183
rect 662 179 668 180
rect 583 175 589 176
rect 583 174 584 175
rect 576 172 584 174
rect 479 170 488 171
rect 583 171 584 172
rect 588 171 589 175
rect 662 175 663 179
rect 667 175 668 179
rect 774 179 780 180
rect 662 174 668 175
rect 686 175 692 176
rect 583 170 589 171
rect 686 171 687 175
rect 691 174 692 175
rect 695 175 701 176
rect 695 174 696 175
rect 691 172 696 174
rect 691 171 692 172
rect 686 170 692 171
rect 695 171 696 172
rect 700 171 701 175
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 800 174 802 184
rect 886 183 887 187
rect 891 186 892 187
rect 1934 187 1935 191
rect 1939 190 1940 191
rect 2238 191 2244 192
rect 1939 188 2074 190
rect 1939 187 1940 188
rect 1934 186 1940 187
rect 891 184 1161 186
rect 891 183 892 184
rect 886 182 892 183
rect 894 179 900 180
rect 807 175 813 176
rect 807 174 808 175
rect 800 172 808 174
rect 695 170 701 171
rect 807 171 808 172
rect 812 171 813 175
rect 894 175 895 179
rect 899 175 900 179
rect 1014 179 1020 180
rect 894 174 900 175
rect 927 175 936 176
rect 807 170 813 171
rect 927 171 928 175
rect 935 171 936 175
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1134 179 1140 180
rect 1014 174 1020 175
rect 1038 175 1044 176
rect 927 170 936 171
rect 1038 171 1039 175
rect 1043 174 1044 175
rect 1047 175 1053 176
rect 1047 174 1048 175
rect 1043 172 1048 174
rect 1043 171 1044 172
rect 1038 170 1044 171
rect 1047 171 1048 172
rect 1052 171 1053 175
rect 1134 175 1135 179
rect 1139 175 1140 179
rect 1134 174 1140 175
rect 1159 174 1161 184
rect 1366 184 1372 185
rect 1326 180 1332 181
rect 1254 179 1260 180
rect 1167 175 1173 176
rect 1167 174 1168 175
rect 1159 172 1168 174
rect 1047 170 1053 171
rect 1167 171 1168 172
rect 1172 171 1173 175
rect 1254 175 1255 179
rect 1259 175 1260 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1366 180 1367 184
rect 1371 180 1372 184
rect 1366 179 1372 180
rect 1398 183 1404 184
rect 1398 179 1399 183
rect 1403 179 1404 183
rect 1462 183 1468 184
rect 1398 178 1404 179
rect 1431 179 1440 180
rect 1254 174 1260 175
rect 1287 175 1293 176
rect 1326 175 1332 176
rect 1431 175 1432 179
rect 1439 175 1440 179
rect 1462 179 1463 183
rect 1467 179 1468 183
rect 1542 183 1548 184
rect 1462 178 1468 179
rect 1495 179 1504 180
rect 1287 174 1288 175
rect 1264 172 1288 174
rect 1167 170 1173 171
rect 1198 171 1204 172
rect 1198 167 1199 171
rect 1203 170 1204 171
rect 1264 170 1266 172
rect 1287 171 1288 172
rect 1292 171 1293 175
rect 1431 174 1440 175
rect 1495 175 1496 179
rect 1503 175 1504 179
rect 1542 179 1543 183
rect 1547 179 1548 183
rect 1638 183 1644 184
rect 1542 178 1548 179
rect 1575 179 1584 180
rect 1495 174 1504 175
rect 1575 175 1576 179
rect 1583 175 1584 179
rect 1638 179 1639 183
rect 1643 179 1644 183
rect 1734 183 1740 184
rect 1638 178 1644 179
rect 1671 179 1680 180
rect 1575 174 1584 175
rect 1671 175 1672 179
rect 1679 175 1680 179
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1838 183 1844 184
rect 1734 178 1740 179
rect 1767 179 1776 180
rect 1671 174 1680 175
rect 1767 175 1768 179
rect 1775 175 1776 179
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1942 183 1948 184
rect 1838 178 1844 179
rect 1870 179 1877 180
rect 1767 174 1776 175
rect 1870 175 1871 179
rect 1876 175 1877 179
rect 1942 179 1943 183
rect 1947 179 1948 183
rect 2046 183 2052 184
rect 1942 178 1948 179
rect 1975 179 1981 180
rect 1975 178 1976 179
rect 1952 176 1976 178
rect 1870 174 1877 175
rect 1894 175 1900 176
rect 1287 170 1293 171
rect 1894 171 1895 175
rect 1899 174 1900 175
rect 1952 174 1954 176
rect 1975 175 1976 176
rect 1980 175 1981 179
rect 2046 179 2047 183
rect 2051 179 2052 183
rect 2046 178 2052 179
rect 2072 178 2074 188
rect 2238 187 2239 191
rect 2243 190 2244 191
rect 2243 188 2370 190
rect 2243 187 2244 188
rect 2238 186 2244 187
rect 2150 183 2156 184
rect 2079 179 2085 180
rect 2079 178 2080 179
rect 2072 176 2080 178
rect 1975 174 1981 175
rect 2079 175 2080 176
rect 2084 175 2085 179
rect 2150 179 2151 183
rect 2155 179 2156 183
rect 2246 183 2252 184
rect 2150 178 2156 179
rect 2182 179 2189 180
rect 2079 174 2085 175
rect 2182 175 2183 179
rect 2188 175 2189 179
rect 2246 179 2247 183
rect 2251 179 2252 183
rect 2342 183 2348 184
rect 2246 178 2252 179
rect 2279 179 2285 180
rect 2279 178 2280 179
rect 2182 174 2189 175
rect 2256 176 2280 178
rect 1899 172 1954 174
rect 1899 171 1900 172
rect 1894 170 1900 171
rect 2158 171 2164 172
rect 1203 168 1266 170
rect 1203 167 1204 168
rect 1198 166 1204 167
rect 2158 167 2159 171
rect 2163 170 2164 171
rect 2256 170 2258 176
rect 2279 175 2280 176
rect 2284 175 2285 179
rect 2342 179 2343 183
rect 2347 179 2348 183
rect 2342 178 2348 179
rect 2368 178 2370 188
rect 2582 184 2588 185
rect 2446 183 2452 184
rect 2375 179 2381 180
rect 2375 178 2376 179
rect 2368 176 2376 178
rect 2279 174 2285 175
rect 2375 175 2376 176
rect 2380 175 2381 179
rect 2446 179 2447 183
rect 2451 179 2452 183
rect 2526 183 2532 184
rect 2446 178 2452 179
rect 2479 179 2485 180
rect 2375 174 2381 175
rect 2479 175 2480 179
rect 2484 178 2485 179
rect 2487 179 2493 180
rect 2487 178 2488 179
rect 2484 176 2488 178
rect 2484 175 2485 176
rect 2479 174 2485 175
rect 2487 175 2488 176
rect 2492 175 2493 179
rect 2526 179 2527 183
rect 2531 179 2532 183
rect 2582 180 2583 184
rect 2587 180 2588 184
rect 2526 178 2532 179
rect 2558 179 2565 180
rect 2582 179 2588 180
rect 2487 174 2493 175
rect 2558 175 2559 179
rect 2564 175 2565 179
rect 2558 174 2565 175
rect 2163 168 2258 170
rect 2163 167 2164 168
rect 2158 166 2164 167
rect 2334 143 2340 144
rect 2334 139 2335 143
rect 2339 142 2340 143
rect 2339 140 2442 142
rect 2339 139 2340 140
rect 2334 138 2340 139
rect 1431 135 1437 136
rect 1398 133 1404 134
rect 1366 132 1372 133
rect 1366 128 1367 132
rect 1371 128 1372 132
rect 1398 129 1399 133
rect 1403 129 1404 133
rect 1431 131 1432 135
rect 1436 134 1437 135
rect 1446 135 1452 136
rect 1446 134 1447 135
rect 1436 132 1447 134
rect 1436 131 1437 132
rect 1431 130 1437 131
rect 1446 131 1447 132
rect 1451 131 1452 135
rect 1487 135 1493 136
rect 1446 130 1452 131
rect 1454 133 1460 134
rect 1398 128 1404 129
rect 1454 129 1455 133
rect 1459 129 1460 133
rect 1487 131 1488 135
rect 1492 134 1493 135
rect 1502 135 1508 136
rect 1502 134 1503 135
rect 1492 132 1503 134
rect 1492 131 1493 132
rect 1487 130 1493 131
rect 1502 131 1503 132
rect 1507 131 1508 135
rect 1543 135 1549 136
rect 1502 130 1508 131
rect 1510 133 1516 134
rect 1454 128 1460 129
rect 1510 129 1511 133
rect 1515 129 1516 133
rect 1543 131 1544 135
rect 1548 134 1549 135
rect 1558 135 1564 136
rect 1558 134 1559 135
rect 1548 132 1559 134
rect 1548 131 1549 132
rect 1543 130 1549 131
rect 1558 131 1559 132
rect 1563 131 1564 135
rect 1599 135 1605 136
rect 1558 130 1564 131
rect 1566 133 1572 134
rect 1510 128 1516 129
rect 1566 129 1567 133
rect 1571 129 1572 133
rect 1599 131 1600 135
rect 1604 134 1605 135
rect 1622 135 1628 136
rect 1622 134 1623 135
rect 1604 132 1623 134
rect 1604 131 1605 132
rect 1599 130 1605 131
rect 1622 131 1623 132
rect 1627 131 1628 135
rect 1663 135 1669 136
rect 1622 130 1628 131
rect 1630 133 1636 134
rect 1566 128 1572 129
rect 1630 129 1631 133
rect 1635 129 1636 133
rect 1663 131 1664 135
rect 1668 134 1669 135
rect 1702 135 1708 136
rect 1702 134 1703 135
rect 1668 132 1703 134
rect 1668 131 1669 132
rect 1663 130 1669 131
rect 1702 131 1703 132
rect 1707 131 1708 135
rect 1743 135 1749 136
rect 1702 130 1708 131
rect 1710 133 1716 134
rect 1630 128 1636 129
rect 1710 129 1711 133
rect 1715 129 1716 133
rect 1743 131 1744 135
rect 1748 134 1749 135
rect 1782 135 1788 136
rect 1782 134 1783 135
rect 1748 132 1783 134
rect 1748 131 1749 132
rect 1743 130 1749 131
rect 1782 131 1783 132
rect 1787 131 1788 135
rect 1822 135 1829 136
rect 1782 130 1788 131
rect 1790 133 1796 134
rect 1710 128 1716 129
rect 1790 129 1791 133
rect 1795 129 1796 133
rect 1822 131 1823 135
rect 1828 131 1829 135
rect 1903 135 1909 136
rect 1822 130 1829 131
rect 1870 133 1876 134
rect 1790 128 1796 129
rect 1870 129 1871 133
rect 1875 129 1876 133
rect 1903 131 1904 135
rect 1908 134 1909 135
rect 1934 135 1940 136
rect 1934 134 1935 135
rect 1908 132 1935 134
rect 1908 131 1909 132
rect 1903 130 1909 131
rect 1934 131 1935 132
rect 1939 131 1940 135
rect 1975 135 1981 136
rect 1934 130 1940 131
rect 1942 133 1948 134
rect 1870 128 1876 129
rect 1942 129 1943 133
rect 1947 129 1948 133
rect 1975 131 1976 135
rect 1980 134 1981 135
rect 2006 135 2012 136
rect 2006 134 2007 135
rect 1980 132 2007 134
rect 1980 131 1981 132
rect 1975 130 1981 131
rect 2006 131 2007 132
rect 2011 131 2012 135
rect 2047 135 2053 136
rect 2006 130 2012 131
rect 2014 133 2020 134
rect 1942 128 1948 129
rect 2014 129 2015 133
rect 2019 129 2020 133
rect 2047 131 2048 135
rect 2052 134 2053 135
rect 2070 135 2076 136
rect 2070 134 2071 135
rect 2052 132 2071 134
rect 2052 131 2053 132
rect 2047 130 2053 131
rect 2070 131 2071 132
rect 2075 131 2076 135
rect 2111 135 2117 136
rect 2070 130 2076 131
rect 2078 133 2084 134
rect 2014 128 2020 129
rect 2078 129 2079 133
rect 2083 129 2084 133
rect 2111 131 2112 135
rect 2116 134 2117 135
rect 2134 135 2140 136
rect 2134 134 2135 135
rect 2116 132 2135 134
rect 2116 131 2117 132
rect 2111 130 2117 131
rect 2134 131 2135 132
rect 2139 131 2140 135
rect 2175 135 2181 136
rect 2134 130 2140 131
rect 2142 133 2148 134
rect 2078 128 2084 129
rect 2142 129 2143 133
rect 2147 129 2148 133
rect 2175 131 2176 135
rect 2180 134 2181 135
rect 2198 135 2204 136
rect 2198 134 2199 135
rect 2180 132 2199 134
rect 2180 131 2181 132
rect 2175 130 2181 131
rect 2198 131 2199 132
rect 2203 131 2204 135
rect 2239 135 2245 136
rect 2198 130 2204 131
rect 2206 133 2212 134
rect 2142 128 2148 129
rect 2206 129 2207 133
rect 2211 129 2212 133
rect 2239 131 2240 135
rect 2244 134 2245 135
rect 2262 135 2268 136
rect 2262 134 2263 135
rect 2244 132 2263 134
rect 2244 131 2245 132
rect 2239 130 2245 131
rect 2262 131 2263 132
rect 2267 131 2268 135
rect 2303 135 2309 136
rect 2262 130 2268 131
rect 2270 133 2276 134
rect 2206 128 2212 129
rect 2270 129 2271 133
rect 2275 129 2276 133
rect 2303 131 2304 135
rect 2308 134 2309 135
rect 2334 135 2340 136
rect 2334 134 2335 135
rect 2308 132 2335 134
rect 2308 131 2309 132
rect 2303 130 2309 131
rect 2334 131 2335 132
rect 2339 131 2340 135
rect 2375 135 2381 136
rect 2334 130 2340 131
rect 2342 133 2348 134
rect 2270 128 2276 129
rect 2342 129 2343 133
rect 2347 129 2348 133
rect 2375 131 2376 135
rect 2380 134 2381 135
rect 2406 135 2412 136
rect 2406 134 2407 135
rect 2380 132 2407 134
rect 2380 131 2381 132
rect 2375 130 2381 131
rect 2406 131 2407 132
rect 2411 131 2412 135
rect 2440 134 2442 140
rect 2447 135 2453 136
rect 2447 134 2448 135
rect 2406 130 2412 131
rect 2414 133 2420 134
rect 2342 128 2348 129
rect 2414 129 2415 133
rect 2419 129 2420 133
rect 2440 132 2448 134
rect 2447 131 2448 132
rect 2452 131 2453 135
rect 2447 130 2453 131
rect 2582 132 2588 133
rect 2414 128 2420 129
rect 2582 128 2583 132
rect 2587 128 2588 132
rect 1366 127 1372 128
rect 2582 127 2588 128
rect 175 123 181 124
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 175 119 176 123
rect 180 122 181 123
rect 190 123 196 124
rect 190 122 191 123
rect 180 120 191 122
rect 180 119 181 120
rect 175 118 181 119
rect 190 119 191 120
rect 195 119 196 123
rect 231 123 237 124
rect 190 118 196 119
rect 198 121 204 122
rect 142 116 148 117
rect 198 117 199 121
rect 203 117 204 121
rect 231 119 232 123
rect 236 122 237 123
rect 246 123 252 124
rect 246 122 247 123
rect 236 120 247 122
rect 236 119 237 120
rect 231 118 237 119
rect 246 119 247 120
rect 251 119 252 123
rect 287 123 293 124
rect 246 118 252 119
rect 254 121 260 122
rect 198 116 204 117
rect 254 117 255 121
rect 259 117 260 121
rect 287 119 288 123
rect 292 122 293 123
rect 302 123 308 124
rect 302 122 303 123
rect 292 120 303 122
rect 292 119 293 120
rect 287 118 293 119
rect 302 119 303 120
rect 307 119 308 123
rect 343 123 349 124
rect 302 118 308 119
rect 310 121 316 122
rect 254 116 260 117
rect 310 117 311 121
rect 315 117 316 121
rect 343 119 344 123
rect 348 122 349 123
rect 358 123 364 124
rect 358 122 359 123
rect 348 120 359 122
rect 348 119 349 120
rect 343 118 349 119
rect 358 119 359 120
rect 363 119 364 123
rect 399 123 405 124
rect 358 118 364 119
rect 366 121 372 122
rect 310 116 316 117
rect 366 117 367 121
rect 371 117 372 121
rect 399 119 400 123
rect 404 122 405 123
rect 414 123 420 124
rect 414 122 415 123
rect 404 120 415 122
rect 404 119 405 120
rect 399 118 405 119
rect 414 119 415 120
rect 419 119 420 123
rect 455 123 461 124
rect 414 118 420 119
rect 422 121 428 122
rect 366 116 372 117
rect 422 117 423 121
rect 427 117 428 121
rect 455 119 456 123
rect 460 122 461 123
rect 470 123 476 124
rect 470 122 471 123
rect 460 120 471 122
rect 460 119 461 120
rect 455 118 461 119
rect 470 119 471 120
rect 475 119 476 123
rect 511 123 517 124
rect 470 118 476 119
rect 478 121 484 122
rect 422 116 428 117
rect 478 117 479 121
rect 483 117 484 121
rect 511 119 512 123
rect 516 122 517 123
rect 526 123 532 124
rect 526 122 527 123
rect 516 120 527 122
rect 516 119 517 120
rect 511 118 517 119
rect 526 119 527 120
rect 531 119 532 123
rect 567 123 573 124
rect 526 118 532 119
rect 534 121 540 122
rect 478 116 484 117
rect 534 117 535 121
rect 539 117 540 121
rect 567 119 568 123
rect 572 122 573 123
rect 582 123 588 124
rect 582 122 583 123
rect 572 120 583 122
rect 572 119 573 120
rect 567 118 573 119
rect 582 119 583 120
rect 587 119 588 123
rect 622 123 629 124
rect 582 118 588 119
rect 590 121 596 122
rect 534 116 540 117
rect 590 117 591 121
rect 595 117 596 121
rect 622 119 623 123
rect 628 119 629 123
rect 679 123 685 124
rect 622 118 629 119
rect 646 121 652 122
rect 590 116 596 117
rect 646 117 647 121
rect 651 117 652 121
rect 679 119 680 123
rect 684 122 685 123
rect 694 123 700 124
rect 694 122 695 123
rect 684 120 695 122
rect 684 119 685 120
rect 679 118 685 119
rect 694 119 695 120
rect 699 119 700 123
rect 735 123 741 124
rect 694 118 700 119
rect 702 121 708 122
rect 646 116 652 117
rect 702 117 703 121
rect 707 117 708 121
rect 735 119 736 123
rect 740 122 741 123
rect 750 123 756 124
rect 750 122 751 123
rect 740 120 751 122
rect 740 119 741 120
rect 735 118 741 119
rect 750 119 751 120
rect 755 119 756 123
rect 791 123 797 124
rect 750 118 756 119
rect 758 121 764 122
rect 702 116 708 117
rect 758 117 759 121
rect 763 117 764 121
rect 791 119 792 123
rect 796 122 797 123
rect 814 123 820 124
rect 814 122 815 123
rect 796 120 815 122
rect 796 119 797 120
rect 791 118 797 119
rect 814 119 815 120
rect 819 119 820 123
rect 855 123 861 124
rect 814 118 820 119
rect 822 121 828 122
rect 758 116 764 117
rect 822 117 823 121
rect 827 117 828 121
rect 855 119 856 123
rect 860 122 861 123
rect 878 123 884 124
rect 878 122 879 123
rect 860 120 879 122
rect 860 119 861 120
rect 855 118 861 119
rect 878 119 879 120
rect 883 119 884 123
rect 919 123 925 124
rect 878 118 884 119
rect 886 121 892 122
rect 822 116 828 117
rect 886 117 887 121
rect 891 117 892 121
rect 919 119 920 123
rect 924 122 925 123
rect 942 123 948 124
rect 942 122 943 123
rect 924 120 943 122
rect 924 119 925 120
rect 919 118 925 119
rect 942 119 943 120
rect 947 119 948 123
rect 983 123 989 124
rect 942 118 948 119
rect 950 121 956 122
rect 886 116 892 117
rect 950 117 951 121
rect 955 117 956 121
rect 983 119 984 123
rect 988 122 989 123
rect 1006 123 1012 124
rect 1006 122 1007 123
rect 988 120 1007 122
rect 988 119 989 120
rect 983 118 989 119
rect 1006 119 1007 120
rect 1011 119 1012 123
rect 1047 123 1053 124
rect 1006 118 1012 119
rect 1014 121 1020 122
rect 950 116 956 117
rect 1014 117 1015 121
rect 1019 117 1020 121
rect 1047 119 1048 123
rect 1052 122 1053 123
rect 1070 123 1076 124
rect 1070 122 1071 123
rect 1052 120 1071 122
rect 1052 119 1053 120
rect 1047 118 1053 119
rect 1070 119 1071 120
rect 1075 119 1076 123
rect 1111 123 1120 124
rect 1070 118 1076 119
rect 1078 121 1084 122
rect 1014 116 1020 117
rect 1078 117 1079 121
rect 1083 117 1084 121
rect 1111 119 1112 123
rect 1119 119 1120 123
rect 1183 123 1189 124
rect 1111 118 1120 119
rect 1150 121 1156 122
rect 1078 116 1084 117
rect 1150 117 1151 121
rect 1155 117 1156 121
rect 1183 119 1184 123
rect 1188 122 1189 123
rect 1206 123 1212 124
rect 1206 122 1207 123
rect 1188 120 1207 122
rect 1188 119 1189 120
rect 1183 118 1189 119
rect 1206 119 1207 120
rect 1211 119 1212 123
rect 1247 123 1253 124
rect 1206 118 1212 119
rect 1214 121 1220 122
rect 1150 116 1156 117
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1247 119 1248 123
rect 1252 122 1253 123
rect 1262 123 1268 124
rect 1262 122 1263 123
rect 1252 120 1263 122
rect 1252 119 1253 120
rect 1247 118 1253 119
rect 1262 119 1263 120
rect 1267 119 1268 123
rect 1303 123 1309 124
rect 1262 118 1268 119
rect 1270 121 1276 122
rect 1214 116 1220 117
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1303 119 1304 123
rect 1308 122 1309 123
rect 1308 120 1322 122
rect 1308 119 1309 120
rect 1303 118 1309 119
rect 1270 116 1276 117
rect 110 115 116 116
rect 1320 110 1322 120
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 1326 115 1332 116
rect 1366 115 1372 116
rect 1366 111 1367 115
rect 1371 111 1372 115
rect 1366 110 1372 111
rect 2582 115 2588 116
rect 2582 111 2583 115
rect 2587 111 2588 115
rect 2582 110 2588 111
rect 1320 108 1350 110
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1326 98 1332 99
rect 1348 98 1350 108
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1470 106 1476 107
rect 1470 102 1471 106
rect 1475 102 1476 106
rect 1470 101 1476 102
rect 1526 106 1532 107
rect 1526 102 1527 106
rect 1531 102 1532 106
rect 1526 101 1532 102
rect 1582 106 1588 107
rect 1582 102 1583 106
rect 1587 102 1588 106
rect 1582 101 1588 102
rect 1646 106 1652 107
rect 1646 102 1647 106
rect 1651 102 1652 106
rect 1646 101 1652 102
rect 1726 106 1732 107
rect 1726 102 1727 106
rect 1731 102 1732 106
rect 1726 101 1732 102
rect 1806 106 1812 107
rect 1806 102 1807 106
rect 1811 102 1812 106
rect 1806 101 1812 102
rect 1886 106 1892 107
rect 1886 102 1887 106
rect 1891 102 1892 106
rect 1886 101 1892 102
rect 1958 106 1964 107
rect 1958 102 1959 106
rect 1963 102 1964 106
rect 1958 101 1964 102
rect 2030 106 2036 107
rect 2030 102 2031 106
rect 2035 102 2036 106
rect 2030 101 2036 102
rect 2094 106 2100 107
rect 2094 102 2095 106
rect 2099 102 2100 106
rect 2094 101 2100 102
rect 2158 106 2164 107
rect 2158 102 2159 106
rect 2163 102 2164 106
rect 2158 101 2164 102
rect 2222 106 2228 107
rect 2222 102 2223 106
rect 2227 102 2228 106
rect 2222 101 2228 102
rect 2286 106 2292 107
rect 2286 102 2287 106
rect 2291 102 2292 106
rect 2286 101 2292 102
rect 2358 106 2364 107
rect 2358 102 2359 106
rect 2363 102 2364 106
rect 2358 101 2364 102
rect 2430 106 2436 107
rect 2430 102 2431 106
rect 2435 102 2436 106
rect 2430 101 2436 102
rect 1391 99 1397 100
rect 1391 98 1392 99
rect 1348 96 1392 98
rect 1391 95 1392 96
rect 1396 95 1397 99
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 606 94 612 95
rect 606 90 607 94
rect 611 90 612 94
rect 606 89 612 90
rect 662 94 668 95
rect 662 90 663 94
rect 667 90 668 94
rect 662 89 668 90
rect 718 94 724 95
rect 718 90 719 94
rect 723 90 724 94
rect 718 89 724 90
rect 774 94 780 95
rect 774 90 775 94
rect 779 90 780 94
rect 774 89 780 90
rect 838 94 844 95
rect 838 90 839 94
rect 843 90 844 94
rect 838 89 844 90
rect 902 94 908 95
rect 902 90 903 94
rect 907 90 908 94
rect 902 89 908 90
rect 966 94 972 95
rect 966 90 967 94
rect 971 90 972 94
rect 966 89 972 90
rect 1030 94 1036 95
rect 1030 90 1031 94
rect 1035 90 1036 94
rect 1030 89 1036 90
rect 1094 94 1100 95
rect 1094 90 1095 94
rect 1099 90 1100 94
rect 1094 89 1100 90
rect 1166 94 1172 95
rect 1166 90 1167 94
rect 1171 90 1172 94
rect 1166 89 1172 90
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1286 94 1292 95
rect 1391 94 1397 95
rect 1446 99 1453 100
rect 1446 95 1447 99
rect 1452 95 1453 99
rect 1446 94 1453 95
rect 1502 99 1509 100
rect 1502 95 1503 99
rect 1508 95 1509 99
rect 1502 94 1509 95
rect 1558 99 1565 100
rect 1558 95 1559 99
rect 1564 95 1565 99
rect 1558 94 1565 95
rect 1622 99 1629 100
rect 1622 95 1623 99
rect 1628 95 1629 99
rect 1622 94 1629 95
rect 1702 99 1709 100
rect 1702 95 1703 99
rect 1708 95 1709 99
rect 1702 94 1709 95
rect 1782 99 1789 100
rect 1782 95 1783 99
rect 1788 95 1789 99
rect 1782 94 1789 95
rect 1863 99 1869 100
rect 1863 95 1864 99
rect 1868 98 1869 99
rect 1894 99 1900 100
rect 1894 98 1895 99
rect 1868 96 1895 98
rect 1868 95 1869 96
rect 1863 94 1869 95
rect 1894 95 1895 96
rect 1899 95 1900 99
rect 1894 94 1900 95
rect 1934 99 1941 100
rect 1934 95 1935 99
rect 1940 95 1941 99
rect 1934 94 1941 95
rect 2006 99 2013 100
rect 2006 95 2007 99
rect 2012 95 2013 99
rect 2006 94 2013 95
rect 2070 99 2077 100
rect 2070 95 2071 99
rect 2076 95 2077 99
rect 2070 94 2077 95
rect 2134 99 2141 100
rect 2134 95 2135 99
rect 2140 95 2141 99
rect 2134 94 2141 95
rect 2198 99 2205 100
rect 2198 95 2199 99
rect 2204 95 2205 99
rect 2198 94 2205 95
rect 2262 99 2269 100
rect 2262 95 2263 99
rect 2268 95 2269 99
rect 2262 94 2269 95
rect 2334 99 2341 100
rect 2334 95 2335 99
rect 2340 95 2341 99
rect 2334 94 2341 95
rect 2406 99 2413 100
rect 2406 95 2407 99
rect 2412 95 2413 99
rect 2406 94 2413 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
rect 190 87 197 88
rect 190 83 191 87
rect 196 83 197 87
rect 190 82 197 83
rect 246 87 253 88
rect 246 83 247 87
rect 252 83 253 87
rect 246 82 253 83
rect 302 87 309 88
rect 302 83 303 87
rect 308 83 309 87
rect 302 82 309 83
rect 358 87 365 88
rect 358 83 359 87
rect 364 83 365 87
rect 358 82 365 83
rect 414 87 421 88
rect 414 83 415 87
rect 420 83 421 87
rect 414 82 421 83
rect 470 87 477 88
rect 470 83 471 87
rect 476 83 477 87
rect 470 82 477 83
rect 526 87 533 88
rect 526 83 527 87
rect 532 83 533 87
rect 526 82 533 83
rect 582 87 589 88
rect 582 83 583 87
rect 588 83 589 87
rect 582 82 589 83
rect 639 87 645 88
rect 639 83 640 87
rect 644 86 645 87
rect 686 87 692 88
rect 686 86 687 87
rect 644 84 687 86
rect 644 83 645 84
rect 639 82 645 83
rect 686 83 687 84
rect 691 83 692 87
rect 686 82 692 83
rect 694 87 701 88
rect 694 83 695 87
rect 700 83 701 87
rect 694 82 701 83
rect 750 87 757 88
rect 750 83 751 87
rect 756 83 757 87
rect 750 82 757 83
rect 814 87 821 88
rect 814 83 815 87
rect 820 83 821 87
rect 814 82 821 83
rect 878 87 885 88
rect 878 83 879 87
rect 884 83 885 87
rect 878 82 885 83
rect 942 87 949 88
rect 942 83 943 87
rect 948 83 949 87
rect 942 82 949 83
rect 1006 87 1013 88
rect 1006 83 1007 87
rect 1012 83 1013 87
rect 1006 82 1013 83
rect 1070 87 1077 88
rect 1070 83 1071 87
rect 1076 83 1077 87
rect 1070 82 1077 83
rect 1143 87 1149 88
rect 1143 83 1144 87
rect 1148 86 1149 87
rect 1198 87 1204 88
rect 1198 86 1199 87
rect 1148 84 1199 86
rect 1148 83 1149 84
rect 1143 82 1149 83
rect 1198 83 1199 84
rect 1203 83 1204 87
rect 1198 82 1204 83
rect 1206 87 1213 88
rect 1206 83 1207 87
rect 1212 83 1213 87
rect 1206 82 1213 83
rect 1262 87 1269 88
rect 1262 83 1263 87
rect 1268 83 1269 87
rect 1262 82 1269 83
<< m3c >>
rect 623 2639 627 2643
rect 583 2631 584 2635
rect 584 2631 587 2635
rect 735 2639 739 2643
rect 695 2631 696 2635
rect 696 2631 699 2635
rect 751 2631 752 2635
rect 752 2631 755 2635
rect 551 2626 555 2630
rect 607 2626 611 2630
rect 663 2626 667 2630
rect 719 2626 723 2630
rect 775 2626 779 2630
rect 1623 2635 1627 2639
rect 1583 2627 1584 2631
rect 1584 2627 1587 2631
rect 1735 2635 1739 2639
rect 1695 2627 1696 2631
rect 1696 2627 1699 2631
rect 1839 2635 1843 2639
rect 1807 2627 1808 2631
rect 1808 2627 1811 2631
rect 1959 2635 1963 2639
rect 2183 2635 2187 2639
rect 1919 2627 1920 2631
rect 1920 2627 1923 2631
rect 2027 2627 2031 2631
rect 2075 2627 2079 2631
rect 2131 2627 2135 2631
rect 1551 2622 1555 2626
rect 111 2617 115 2621
rect 1607 2622 1611 2626
rect 1663 2622 1667 2626
rect 1719 2622 1723 2626
rect 1775 2622 1779 2626
rect 1831 2622 1835 2626
rect 1887 2622 1891 2626
rect 1943 2622 1947 2626
rect 1999 2622 2003 2626
rect 2055 2622 2059 2626
rect 2111 2622 2115 2626
rect 2167 2622 2171 2626
rect 1327 2617 1331 2621
rect 1367 2613 1371 2617
rect 2583 2613 2587 2617
rect 583 2607 587 2611
rect 111 2600 115 2604
rect 535 2599 539 2603
rect 559 2595 563 2599
rect 591 2599 595 2603
rect 623 2595 624 2599
rect 624 2595 627 2599
rect 647 2599 651 2603
rect 695 2607 699 2611
rect 703 2599 707 2603
rect 735 2595 736 2599
rect 736 2595 739 2599
rect 759 2599 763 2603
rect 1327 2600 1331 2604
rect 1583 2603 1587 2607
rect 1367 2596 1371 2600
rect 1535 2595 1539 2599
rect 1447 2587 1451 2591
rect 1591 2595 1595 2599
rect 1623 2591 1624 2595
rect 1624 2591 1627 2595
rect 1647 2595 1651 2599
rect 1695 2603 1699 2607
rect 1703 2595 1707 2599
rect 1735 2591 1736 2595
rect 1736 2591 1739 2595
rect 1759 2595 1763 2599
rect 1807 2603 1811 2607
rect 1815 2595 1819 2599
rect 1839 2591 1843 2595
rect 1871 2595 1875 2599
rect 1919 2603 1923 2607
rect 1927 2595 1931 2599
rect 1959 2591 1960 2595
rect 1960 2591 1963 2595
rect 1983 2595 1987 2599
rect 2039 2595 2043 2599
rect 2075 2591 2076 2595
rect 2076 2591 2079 2595
rect 2095 2595 2099 2599
rect 2131 2591 2132 2595
rect 2132 2591 2135 2595
rect 2151 2595 2155 2599
rect 2583 2596 2587 2600
rect 2183 2591 2184 2595
rect 2184 2591 2187 2595
rect 239 2575 243 2579
rect 111 2564 115 2568
rect 215 2565 219 2569
rect 263 2567 267 2571
rect 271 2565 275 2569
rect 319 2567 323 2571
rect 327 2565 331 2569
rect 355 2567 359 2571
rect 383 2565 387 2569
rect 439 2565 443 2569
rect 527 2575 531 2579
rect 495 2565 499 2569
rect 551 2565 555 2569
rect 599 2567 603 2571
rect 687 2575 691 2579
rect 607 2565 611 2569
rect 663 2565 667 2569
rect 711 2567 715 2571
rect 719 2565 723 2569
rect 751 2567 752 2571
rect 752 2567 755 2571
rect 775 2565 779 2569
rect 831 2565 835 2569
rect 887 2565 891 2569
rect 975 2575 979 2579
rect 943 2565 947 2569
rect 999 2565 1003 2569
rect 1047 2567 1051 2571
rect 1055 2565 1059 2569
rect 1103 2567 1107 2571
rect 1111 2565 1115 2569
rect 1327 2564 1331 2568
rect 1367 2560 1371 2564
rect 1439 2561 1443 2565
rect 1535 2563 1539 2567
rect 1543 2561 1547 2565
rect 1647 2563 1651 2567
rect 1655 2561 1659 2565
rect 1759 2563 1763 2567
rect 1767 2561 1771 2565
rect 1871 2563 1875 2567
rect 1879 2561 1883 2565
rect 1903 2563 1907 2567
rect 1991 2561 1995 2565
rect 2027 2563 2028 2567
rect 2028 2563 2031 2567
rect 2071 2567 2075 2571
rect 2111 2561 2115 2565
rect 2231 2561 2235 2565
rect 2351 2561 2355 2565
rect 2583 2560 2587 2564
rect 111 2547 115 2551
rect 1327 2547 1331 2551
rect 1367 2543 1371 2547
rect 231 2538 235 2542
rect 287 2538 291 2542
rect 343 2538 347 2542
rect 399 2538 403 2542
rect 455 2538 459 2542
rect 511 2538 515 2542
rect 567 2538 571 2542
rect 623 2538 627 2542
rect 679 2538 683 2542
rect 735 2538 739 2542
rect 791 2538 795 2542
rect 847 2538 851 2542
rect 903 2538 907 2542
rect 959 2538 963 2542
rect 1015 2538 1019 2542
rect 1071 2538 1075 2542
rect 2583 2543 2587 2547
rect 1127 2538 1131 2542
rect 239 2531 243 2535
rect 263 2531 264 2535
rect 264 2531 267 2535
rect 319 2531 320 2535
rect 320 2531 323 2535
rect 527 2531 531 2535
rect 559 2531 563 2535
rect 599 2531 600 2535
rect 600 2531 603 2535
rect 687 2531 691 2535
rect 711 2531 712 2535
rect 712 2531 715 2535
rect 975 2531 979 2535
rect 1047 2531 1048 2535
rect 1048 2531 1051 2535
rect 1103 2531 1104 2535
rect 1104 2531 1107 2535
rect 1455 2534 1459 2538
rect 1559 2534 1563 2538
rect 1671 2534 1675 2538
rect 1783 2534 1787 2538
rect 1895 2534 1899 2538
rect 2007 2534 2011 2538
rect 2127 2534 2131 2538
rect 2247 2534 2251 2538
rect 2367 2534 2371 2538
rect 355 2519 359 2523
rect 387 2515 391 2519
rect 443 2515 447 2519
rect 655 2515 656 2519
rect 656 2515 659 2519
rect 707 2515 711 2519
rect 759 2515 763 2519
rect 1023 2523 1027 2527
rect 1447 2527 1451 2531
rect 1535 2527 1536 2531
rect 1536 2527 1539 2531
rect 1647 2527 1648 2531
rect 1648 2527 1651 2531
rect 1759 2527 1760 2531
rect 1760 2527 1763 2531
rect 1871 2527 1872 2531
rect 1872 2527 1875 2531
rect 2071 2527 2075 2531
rect 2315 2527 2319 2531
rect 979 2515 983 2519
rect 367 2510 371 2514
rect 423 2510 427 2514
rect 487 2510 491 2514
rect 551 2510 555 2514
rect 615 2510 619 2514
rect 679 2510 683 2514
rect 743 2510 747 2514
rect 807 2510 811 2514
rect 871 2510 875 2514
rect 943 2510 947 2514
rect 1015 2510 1019 2514
rect 1543 2507 1547 2511
rect 1571 2507 1575 2511
rect 1651 2507 1655 2511
rect 1739 2507 1743 2511
rect 1827 2507 1831 2511
rect 1975 2507 1976 2511
rect 1976 2507 1979 2511
rect 2019 2507 2023 2511
rect 2115 2507 2119 2511
rect 2271 2507 2272 2511
rect 2272 2507 2275 2511
rect 2391 2507 2395 2511
rect 111 2501 115 2505
rect 1327 2501 1331 2505
rect 1551 2502 1555 2506
rect 1631 2502 1635 2506
rect 1719 2502 1723 2506
rect 1807 2502 1811 2506
rect 1903 2502 1907 2506
rect 1999 2502 2003 2506
rect 2095 2502 2099 2506
rect 2191 2502 2195 2506
rect 2295 2502 2299 2506
rect 2399 2502 2403 2506
rect 655 2491 659 2495
rect 1367 2493 1371 2497
rect 2583 2493 2587 2497
rect 111 2484 115 2488
rect 351 2483 355 2487
rect 387 2479 388 2483
rect 388 2479 391 2483
rect 407 2483 411 2487
rect 443 2479 444 2483
rect 444 2479 447 2483
rect 471 2483 475 2487
rect 535 2483 539 2487
rect 599 2483 603 2487
rect 623 2479 627 2483
rect 663 2483 667 2487
rect 707 2479 711 2483
rect 727 2483 731 2487
rect 759 2479 760 2483
rect 760 2479 763 2483
rect 791 2483 795 2487
rect 855 2483 859 2487
rect 927 2483 931 2487
rect 979 2483 983 2487
rect 999 2483 1003 2487
rect 1327 2484 1331 2488
rect 1023 2479 1027 2483
rect 2271 2483 2275 2487
rect 1367 2476 1371 2480
rect 1535 2475 1539 2479
rect 1571 2471 1572 2475
rect 1572 2471 1575 2475
rect 1615 2475 1619 2479
rect 1651 2471 1652 2475
rect 1652 2471 1655 2475
rect 1703 2475 1707 2479
rect 1739 2471 1740 2475
rect 1740 2471 1743 2475
rect 1791 2475 1795 2479
rect 1827 2471 1828 2475
rect 1828 2471 1831 2475
rect 1887 2475 1891 2479
rect 1655 2463 1659 2467
rect 1983 2475 1987 2479
rect 2019 2471 2020 2475
rect 2020 2471 2023 2475
rect 2079 2475 2083 2479
rect 2115 2471 2116 2475
rect 2116 2471 2119 2475
rect 2175 2475 2179 2479
rect 2255 2471 2259 2475
rect 2279 2475 2283 2479
rect 2315 2471 2316 2475
rect 2316 2471 2319 2475
rect 2383 2475 2387 2479
rect 2583 2476 2587 2480
rect 279 2455 283 2459
rect 111 2444 115 2448
rect 271 2445 275 2449
rect 327 2447 331 2451
rect 335 2445 339 2449
rect 391 2447 395 2451
rect 399 2445 403 2449
rect 423 2447 427 2451
rect 471 2445 475 2449
rect 551 2445 555 2449
rect 719 2455 723 2459
rect 631 2445 635 2449
rect 711 2445 715 2449
rect 775 2447 779 2451
rect 783 2445 787 2449
rect 855 2447 859 2451
rect 863 2445 867 2449
rect 943 2445 947 2449
rect 1015 2447 1019 2451
rect 1023 2445 1027 2449
rect 1975 2451 1979 2455
rect 1327 2444 1331 2448
rect 1367 2440 1371 2444
rect 1647 2441 1651 2445
rect 1695 2443 1699 2447
rect 1703 2441 1707 2445
rect 1759 2443 1763 2447
rect 1767 2441 1771 2445
rect 1831 2443 1835 2447
rect 1839 2441 1843 2445
rect 1903 2443 1907 2447
rect 1911 2441 1915 2445
rect 1935 2443 1939 2447
rect 1991 2441 1995 2445
rect 2071 2443 2075 2447
rect 2079 2441 2083 2445
rect 2159 2443 2163 2447
rect 2167 2441 2171 2445
rect 2211 2447 2215 2451
rect 2263 2441 2267 2445
rect 2359 2441 2363 2445
rect 2391 2443 2392 2447
rect 2392 2443 2395 2447
rect 2463 2447 2467 2451
rect 2455 2441 2459 2445
rect 2527 2441 2531 2445
rect 2583 2440 2587 2444
rect 111 2427 115 2431
rect 1327 2427 1331 2431
rect 1367 2423 1371 2427
rect 287 2418 291 2422
rect 351 2418 355 2422
rect 415 2418 419 2422
rect 487 2418 491 2422
rect 567 2418 571 2422
rect 647 2418 651 2422
rect 727 2418 731 2422
rect 799 2418 803 2422
rect 879 2418 883 2422
rect 959 2418 963 2422
rect 2583 2423 2587 2427
rect 1039 2418 1043 2422
rect 279 2411 283 2415
rect 327 2411 328 2415
rect 328 2411 331 2415
rect 391 2411 392 2415
rect 392 2411 395 2415
rect 623 2411 624 2415
rect 624 2411 627 2415
rect 719 2411 723 2415
rect 775 2411 776 2415
rect 776 2411 779 2415
rect 855 2411 856 2415
rect 856 2411 859 2415
rect 935 2411 936 2415
rect 936 2411 939 2415
rect 1015 2411 1016 2415
rect 1016 2411 1019 2415
rect 1663 2414 1667 2418
rect 1719 2414 1723 2418
rect 1783 2414 1787 2418
rect 1855 2414 1859 2418
rect 1927 2414 1931 2418
rect 2007 2414 2011 2418
rect 2095 2414 2099 2418
rect 2183 2414 2187 2418
rect 2279 2414 2283 2418
rect 2375 2414 2379 2418
rect 2471 2414 2475 2418
rect 2543 2414 2547 2418
rect 1655 2407 1659 2411
rect 1695 2407 1696 2411
rect 1696 2407 1699 2411
rect 1759 2407 1760 2411
rect 1760 2407 1763 2411
rect 1831 2407 1832 2411
rect 1832 2407 1835 2411
rect 1903 2407 1904 2411
rect 1904 2407 1907 2411
rect 1935 2403 1939 2407
rect 1963 2407 1967 2411
rect 2071 2407 2072 2411
rect 2072 2407 2075 2411
rect 2159 2407 2160 2411
rect 2160 2407 2163 2411
rect 2255 2407 2256 2411
rect 2256 2407 2259 2411
rect 2439 2407 2443 2411
rect 2463 2407 2467 2411
rect 2559 2407 2563 2411
rect 239 2395 243 2399
rect 267 2395 271 2399
rect 423 2395 427 2399
rect 451 2395 455 2399
rect 547 2395 551 2399
rect 703 2395 704 2399
rect 704 2395 707 2399
rect 747 2395 751 2399
rect 843 2395 847 2399
rect 247 2390 251 2394
rect 335 2390 339 2394
rect 431 2390 435 2394
rect 527 2390 531 2394
rect 631 2390 635 2394
rect 727 2390 731 2394
rect 823 2390 827 2394
rect 919 2390 923 2394
rect 1015 2390 1019 2394
rect 1111 2390 1115 2394
rect 1447 2391 1451 2395
rect 2055 2399 2059 2403
rect 1579 2391 1583 2395
rect 1683 2391 1687 2395
rect 2015 2391 2016 2395
rect 2016 2391 2019 2395
rect 2127 2391 2131 2395
rect 2211 2391 2212 2395
rect 2212 2391 2215 2395
rect 2247 2391 2251 2395
rect 2423 2391 2424 2395
rect 2424 2391 2427 2395
rect 2535 2391 2539 2395
rect 1455 2386 1459 2390
rect 111 2381 115 2385
rect 1559 2386 1563 2390
rect 1663 2386 1667 2390
rect 1759 2386 1763 2390
rect 1855 2386 1859 2390
rect 1943 2386 1947 2390
rect 2039 2386 2043 2390
rect 2135 2386 2139 2390
rect 2231 2386 2235 2390
rect 2335 2386 2339 2390
rect 2447 2386 2451 2390
rect 2543 2386 2547 2390
rect 1327 2381 1331 2385
rect 1367 2377 1371 2381
rect 2583 2377 2587 2381
rect 703 2371 707 2375
rect 111 2364 115 2368
rect 231 2363 235 2367
rect 267 2359 268 2363
rect 268 2359 271 2363
rect 319 2363 323 2367
rect 355 2359 356 2363
rect 356 2359 359 2363
rect 415 2363 419 2367
rect 451 2359 452 2363
rect 452 2359 455 2363
rect 511 2363 515 2367
rect 547 2359 548 2363
rect 548 2359 551 2363
rect 615 2363 619 2367
rect 647 2359 648 2363
rect 648 2359 651 2363
rect 711 2363 715 2367
rect 747 2359 748 2363
rect 748 2359 751 2363
rect 807 2363 811 2367
rect 843 2359 844 2363
rect 844 2359 847 2363
rect 903 2363 907 2367
rect 935 2359 936 2363
rect 936 2359 939 2363
rect 999 2363 1003 2367
rect 1095 2363 1099 2367
rect 1327 2364 1331 2368
rect 2015 2367 2019 2371
rect 1367 2360 1371 2364
rect 1439 2359 1443 2363
rect 1535 2355 1539 2359
rect 1543 2359 1547 2363
rect 1579 2355 1580 2359
rect 1580 2355 1583 2359
rect 1647 2359 1651 2363
rect 1683 2355 1684 2359
rect 1684 2355 1687 2359
rect 1743 2359 1747 2363
rect 1839 2359 1843 2363
rect 1863 2355 1867 2359
rect 1927 2359 1931 2363
rect 1963 2355 1964 2359
rect 1964 2355 1967 2359
rect 2023 2359 2027 2363
rect 2055 2355 2056 2359
rect 2056 2355 2059 2359
rect 2119 2359 2123 2363
rect 2215 2359 2219 2363
rect 2247 2355 2248 2359
rect 2248 2355 2251 2359
rect 2319 2359 2323 2363
rect 2375 2355 2379 2359
rect 2431 2359 2435 2363
rect 2439 2351 2443 2355
rect 2527 2359 2531 2363
rect 2583 2360 2587 2364
rect 2559 2355 2560 2359
rect 2560 2355 2563 2359
rect 167 2339 171 2343
rect 111 2328 115 2332
rect 159 2329 163 2333
rect 255 2331 259 2335
rect 263 2329 267 2333
rect 347 2331 351 2335
rect 375 2329 379 2333
rect 479 2331 483 2335
rect 487 2329 491 2333
rect 591 2331 595 2335
rect 735 2339 739 2343
rect 599 2329 603 2333
rect 711 2329 715 2333
rect 807 2331 811 2335
rect 815 2329 819 2333
rect 903 2331 907 2335
rect 911 2329 915 2333
rect 1007 2329 1011 2333
rect 1095 2331 1099 2335
rect 1103 2329 1107 2333
rect 1191 2331 1195 2335
rect 1199 2329 1203 2333
rect 1447 2335 1451 2339
rect 1327 2328 1331 2332
rect 1367 2324 1371 2328
rect 1399 2325 1403 2329
rect 1447 2327 1451 2331
rect 1455 2325 1459 2329
rect 1503 2327 1507 2331
rect 2127 2335 2131 2339
rect 1511 2325 1515 2329
rect 1567 2325 1571 2329
rect 1631 2327 1635 2331
rect 1639 2325 1643 2329
rect 1719 2327 1723 2331
rect 1727 2325 1731 2329
rect 1815 2327 1819 2331
rect 1823 2325 1827 2329
rect 1935 2327 1939 2331
rect 1943 2325 1947 2329
rect 2071 2327 2075 2331
rect 2079 2325 2083 2329
rect 2215 2327 2219 2331
rect 2223 2325 2227 2329
rect 2383 2325 2387 2329
rect 2415 2327 2416 2331
rect 2416 2327 2419 2331
rect 2535 2331 2539 2335
rect 2527 2325 2531 2329
rect 2583 2324 2587 2328
rect 111 2311 115 2315
rect 1327 2311 1331 2315
rect 1367 2307 1371 2311
rect 175 2302 179 2306
rect 279 2302 283 2306
rect 391 2302 395 2306
rect 503 2302 507 2306
rect 615 2302 619 2306
rect 727 2302 731 2306
rect 831 2302 835 2306
rect 927 2302 931 2306
rect 1023 2302 1027 2306
rect 1119 2302 1123 2306
rect 2583 2307 2587 2311
rect 1215 2302 1219 2306
rect 167 2295 171 2299
rect 255 2295 256 2299
rect 256 2295 259 2299
rect 355 2295 359 2299
rect 479 2295 480 2299
rect 480 2295 483 2299
rect 591 2295 592 2299
rect 592 2295 595 2299
rect 735 2295 739 2299
rect 807 2295 808 2299
rect 808 2295 811 2299
rect 903 2295 904 2299
rect 904 2295 907 2299
rect 1015 2295 1019 2299
rect 1095 2295 1096 2299
rect 1096 2295 1099 2299
rect 1191 2295 1192 2299
rect 1192 2295 1195 2299
rect 1415 2298 1419 2302
rect 1471 2298 1475 2302
rect 1527 2298 1531 2302
rect 1583 2298 1587 2302
rect 1655 2298 1659 2302
rect 1743 2298 1747 2302
rect 1839 2298 1843 2302
rect 1959 2298 1963 2302
rect 2095 2298 2099 2302
rect 2239 2298 2243 2302
rect 2399 2298 2403 2302
rect 2543 2298 2547 2302
rect 647 2287 651 2291
rect 135 2279 136 2283
rect 136 2279 139 2283
rect 347 2279 351 2283
rect 443 2279 447 2283
rect 531 2279 535 2283
rect 1111 2287 1115 2291
rect 1307 2291 1311 2295
rect 1447 2291 1448 2295
rect 1448 2291 1451 2295
rect 1503 2291 1504 2295
rect 1504 2291 1507 2295
rect 1535 2291 1539 2295
rect 1631 2291 1632 2295
rect 1632 2291 1635 2295
rect 1719 2291 1720 2295
rect 1720 2291 1723 2295
rect 1863 2291 1867 2295
rect 1935 2291 1936 2295
rect 1936 2291 1939 2295
rect 2071 2291 2072 2295
rect 2072 2291 2075 2295
rect 2215 2291 2216 2295
rect 2216 2291 2219 2295
rect 2375 2291 2376 2295
rect 2376 2291 2379 2295
rect 2559 2291 2563 2295
rect 823 2279 827 2283
rect 907 2279 911 2283
rect 1079 2279 1080 2283
rect 1080 2279 1083 2283
rect 1199 2279 1203 2283
rect 1279 2279 1283 2283
rect 159 2274 163 2278
rect 247 2274 251 2278
rect 375 2274 379 2278
rect 511 2274 515 2278
rect 639 2274 643 2278
rect 767 2274 771 2278
rect 887 2274 891 2278
rect 999 2274 1003 2278
rect 1103 2274 1107 2278
rect 1207 2274 1211 2278
rect 1287 2274 1291 2278
rect 1391 2271 1392 2275
rect 1392 2271 1395 2275
rect 1487 2271 1491 2275
rect 1663 2275 1667 2279
rect 1711 2271 1712 2275
rect 1712 2271 1715 2275
rect 1815 2271 1819 2275
rect 2415 2279 2419 2283
rect 1987 2271 1991 2275
rect 2187 2271 2191 2275
rect 2275 2271 2279 2275
rect 2383 2271 2384 2275
rect 2384 2271 2387 2275
rect 2415 2271 2419 2275
rect 2507 2271 2511 2275
rect 111 2265 115 2269
rect 1327 2265 1331 2269
rect 1415 2266 1419 2270
rect 1495 2266 1499 2270
rect 1615 2266 1619 2270
rect 1735 2266 1739 2270
rect 1855 2266 1859 2270
rect 1967 2266 1971 2270
rect 2071 2266 2075 2270
rect 2167 2266 2171 2270
rect 2255 2266 2259 2270
rect 2335 2266 2339 2270
rect 2407 2266 2411 2270
rect 2487 2266 2491 2270
rect 2543 2266 2547 2270
rect 135 2255 139 2259
rect 111 2248 115 2252
rect 143 2247 147 2251
rect 167 2243 171 2247
rect 231 2247 235 2251
rect 1079 2255 1083 2259
rect 1367 2257 1371 2261
rect 2583 2257 2587 2261
rect 359 2247 363 2251
rect 443 2247 447 2251
rect 495 2247 499 2251
rect 531 2243 532 2247
rect 532 2243 535 2247
rect 623 2247 627 2251
rect 647 2243 651 2247
rect 751 2247 755 2251
rect 823 2243 827 2247
rect 871 2247 875 2251
rect 907 2243 908 2247
rect 908 2243 911 2247
rect 983 2247 987 2251
rect 1015 2243 1016 2247
rect 1016 2243 1019 2247
rect 1087 2247 1091 2251
rect 1111 2243 1115 2247
rect 1191 2247 1195 2251
rect 1271 2247 1275 2251
rect 1327 2248 1331 2252
rect 1391 2247 1395 2251
rect 1307 2243 1308 2247
rect 1308 2243 1311 2247
rect 1367 2240 1371 2244
rect 1399 2239 1403 2243
rect 1279 2231 1283 2235
rect 1479 2239 1483 2243
rect 1711 2247 1715 2251
rect 1599 2239 1603 2243
rect 1487 2227 1491 2231
rect 1719 2239 1723 2243
rect 1751 2235 1752 2239
rect 1752 2235 1755 2239
rect 1839 2239 1843 2243
rect 1951 2239 1955 2243
rect 1987 2235 1988 2239
rect 1988 2235 1991 2239
rect 2055 2239 2059 2243
rect 2151 2239 2155 2243
rect 2187 2235 2188 2239
rect 2188 2235 2191 2239
rect 2239 2239 2243 2243
rect 2275 2235 2276 2239
rect 2276 2235 2279 2239
rect 2319 2239 2323 2243
rect 2391 2239 2395 2243
rect 2415 2231 2419 2235
rect 2423 2235 2424 2239
rect 2424 2235 2427 2239
rect 2471 2239 2475 2243
rect 2507 2235 2508 2239
rect 2508 2235 2511 2239
rect 2527 2239 2531 2243
rect 2583 2240 2587 2244
rect 2559 2235 2560 2239
rect 2560 2235 2563 2239
rect 1199 2215 1203 2219
rect 111 2204 115 2208
rect 143 2205 147 2209
rect 223 2207 227 2211
rect 231 2205 235 2209
rect 351 2207 355 2211
rect 359 2205 363 2209
rect 487 2207 491 2211
rect 495 2205 499 2209
rect 615 2207 619 2211
rect 623 2205 627 2209
rect 647 2207 651 2211
rect 751 2205 755 2209
rect 863 2207 867 2211
rect 871 2205 875 2209
rect 975 2207 979 2211
rect 983 2205 987 2209
rect 1079 2207 1083 2211
rect 1087 2205 1091 2209
rect 1183 2207 1187 2211
rect 1191 2205 1195 2209
rect 1263 2207 1267 2211
rect 1271 2205 1275 2209
rect 1327 2204 1331 2208
rect 1367 2192 1371 2196
rect 1455 2193 1459 2197
rect 1527 2195 1531 2199
rect 1535 2193 1539 2197
rect 1623 2195 1627 2199
rect 1631 2193 1635 2197
rect 1663 2195 1664 2199
rect 1664 2195 1667 2199
rect 1743 2193 1747 2197
rect 1855 2195 1859 2199
rect 1863 2193 1867 2197
rect 1975 2195 1979 2199
rect 1983 2193 1987 2197
rect 2007 2195 2011 2199
rect 2095 2193 2099 2197
rect 2199 2195 2203 2199
rect 2207 2193 2211 2197
rect 2303 2195 2307 2199
rect 2311 2193 2315 2197
rect 2339 2195 2343 2199
rect 2383 2199 2387 2203
rect 2423 2193 2427 2197
rect 2527 2193 2531 2197
rect 2583 2192 2587 2196
rect 111 2187 115 2191
rect 1327 2187 1331 2191
rect 159 2178 163 2182
rect 247 2178 251 2182
rect 375 2178 379 2182
rect 511 2178 515 2182
rect 639 2178 643 2182
rect 767 2178 771 2182
rect 887 2178 891 2182
rect 999 2178 1003 2182
rect 1103 2178 1107 2182
rect 1207 2178 1211 2182
rect 1287 2178 1291 2182
rect 167 2171 171 2175
rect 223 2171 224 2175
rect 224 2171 227 2175
rect 351 2171 352 2175
rect 352 2171 355 2175
rect 487 2171 488 2175
rect 488 2171 491 2175
rect 615 2171 616 2175
rect 616 2171 619 2175
rect 855 2171 859 2175
rect 863 2171 864 2175
rect 864 2171 867 2175
rect 975 2171 976 2175
rect 976 2171 979 2175
rect 1079 2171 1080 2175
rect 1080 2171 1083 2175
rect 1183 2171 1184 2175
rect 1184 2171 1187 2175
rect 1263 2171 1264 2175
rect 1264 2171 1267 2175
rect 1367 2175 1371 2179
rect 2583 2175 2587 2179
rect 1471 2166 1475 2170
rect 1551 2166 1555 2170
rect 1647 2166 1651 2170
rect 1759 2166 1763 2170
rect 1879 2166 1883 2170
rect 1999 2166 2003 2170
rect 2111 2166 2115 2170
rect 2223 2166 2227 2170
rect 2327 2166 2331 2170
rect 2439 2166 2443 2170
rect 2543 2166 2547 2170
rect 139 2155 140 2159
rect 140 2155 143 2159
rect 179 2155 183 2159
rect 235 2155 239 2159
rect 331 2155 335 2159
rect 563 2155 567 2159
rect 751 2155 752 2159
rect 752 2155 755 2159
rect 795 2155 799 2159
rect 899 2155 903 2159
rect 1091 2155 1095 2159
rect 159 2150 163 2154
rect 215 2150 219 2154
rect 311 2150 315 2154
rect 423 2150 427 2154
rect 543 2150 547 2154
rect 663 2150 667 2154
rect 775 2150 779 2154
rect 879 2150 883 2154
rect 975 2150 979 2154
rect 1071 2150 1075 2154
rect 1167 2150 1171 2154
rect 1271 2150 1275 2154
rect 1527 2159 1528 2163
rect 1528 2159 1531 2163
rect 1623 2159 1624 2163
rect 1624 2159 1627 2163
rect 1751 2159 1755 2163
rect 1855 2159 1856 2163
rect 1856 2159 1859 2163
rect 1975 2159 1976 2163
rect 1976 2159 1979 2163
rect 2075 2159 2079 2163
rect 2199 2159 2200 2163
rect 2200 2159 2203 2163
rect 2303 2159 2304 2163
rect 2304 2159 2307 2163
rect 2559 2159 2563 2163
rect 1511 2147 1512 2151
rect 1512 2147 1515 2151
rect 1543 2151 1547 2155
rect 1623 2147 1627 2151
rect 1683 2147 1687 2151
rect 1815 2147 1816 2151
rect 1816 2147 1819 2151
rect 2007 2151 2011 2155
rect 2047 2147 2051 2151
rect 2135 2147 2136 2151
rect 2136 2147 2139 2151
rect 2295 2151 2299 2155
rect 2339 2147 2340 2151
rect 2340 2147 2343 2151
rect 2535 2147 2539 2151
rect 111 2141 115 2145
rect 1327 2141 1331 2145
rect 1535 2142 1539 2146
rect 1631 2142 1635 2146
rect 1735 2142 1739 2146
rect 1839 2142 1843 2146
rect 1951 2142 1955 2146
rect 2055 2142 2059 2146
rect 2159 2142 2163 2146
rect 2263 2142 2267 2146
rect 2359 2142 2363 2146
rect 2463 2142 2467 2146
rect 2543 2142 2547 2146
rect 1367 2133 1371 2137
rect 2583 2133 2587 2137
rect 111 2124 115 2128
rect 143 2123 147 2127
rect 179 2119 180 2123
rect 180 2119 183 2123
rect 199 2123 203 2127
rect 235 2119 236 2123
rect 236 2119 239 2123
rect 295 2123 299 2127
rect 331 2119 332 2123
rect 332 2119 335 2123
rect 407 2123 411 2127
rect 527 2123 531 2127
rect 563 2119 564 2123
rect 564 2119 567 2123
rect 647 2123 651 2127
rect 671 2119 675 2123
rect 759 2123 763 2127
rect 795 2119 796 2123
rect 796 2119 799 2123
rect 863 2123 867 2127
rect 899 2119 900 2123
rect 900 2119 903 2123
rect 959 2123 963 2127
rect 1055 2123 1059 2127
rect 1091 2119 1092 2123
rect 1092 2119 1095 2123
rect 1151 2123 1155 2127
rect 1255 2123 1259 2127
rect 1327 2124 1331 2128
rect 1511 2123 1515 2127
rect 1287 2119 1288 2123
rect 1288 2119 1291 2123
rect 1367 2116 1371 2120
rect 1519 2115 1523 2119
rect 1543 2111 1547 2115
rect 1615 2115 1619 2119
rect 1815 2123 1819 2127
rect 1719 2115 1723 2119
rect 1623 2103 1627 2107
rect 1823 2115 1827 2119
rect 1855 2111 1856 2115
rect 1856 2111 1859 2115
rect 1935 2115 1939 2119
rect 2135 2123 2139 2127
rect 2039 2115 2043 2119
rect 2075 2111 2076 2115
rect 2076 2111 2079 2115
rect 2143 2115 2147 2119
rect 2047 2103 2051 2107
rect 2247 2115 2251 2119
rect 2343 2115 2347 2119
rect 2447 2115 2451 2119
rect 2479 2111 2480 2115
rect 2480 2111 2483 2115
rect 2527 2115 2531 2119
rect 2583 2116 2587 2120
rect 2559 2111 2560 2115
rect 2560 2111 2563 2115
rect 751 2091 755 2095
rect 111 2080 115 2084
rect 263 2081 267 2085
rect 319 2083 323 2087
rect 327 2081 331 2085
rect 391 2083 395 2087
rect 399 2081 403 2085
rect 471 2083 475 2087
rect 479 2081 483 2085
rect 559 2083 563 2087
rect 567 2081 571 2085
rect 647 2083 651 2087
rect 655 2081 659 2085
rect 679 2083 683 2087
rect 735 2081 739 2085
rect 807 2083 811 2087
rect 815 2081 819 2085
rect 879 2083 883 2087
rect 887 2081 891 2085
rect 959 2083 963 2087
rect 967 2081 971 2085
rect 1039 2083 1043 2087
rect 1047 2081 1051 2085
rect 1119 2083 1123 2087
rect 1127 2081 1131 2085
rect 1327 2080 1331 2084
rect 1367 2080 1371 2084
rect 1431 2081 1435 2085
rect 1527 2083 1531 2087
rect 1535 2081 1539 2085
rect 1639 2083 1643 2087
rect 1647 2081 1651 2085
rect 1683 2083 1684 2087
rect 1684 2083 1687 2087
rect 1759 2081 1763 2085
rect 1787 2083 1791 2087
rect 1863 2081 1867 2085
rect 1967 2081 1971 2085
rect 2063 2083 2067 2087
rect 2071 2081 2075 2085
rect 2167 2083 2171 2087
rect 2175 2081 2179 2085
rect 2263 2083 2267 2087
rect 2271 2081 2275 2085
rect 2295 2083 2299 2087
rect 2359 2081 2363 2085
rect 2423 2083 2427 2087
rect 2431 2087 2435 2091
rect 2455 2081 2459 2085
rect 2535 2087 2539 2091
rect 2527 2081 2531 2085
rect 2583 2080 2587 2084
rect 111 2063 115 2067
rect 1327 2063 1331 2067
rect 1367 2063 1371 2067
rect 2583 2063 2587 2067
rect 279 2054 283 2058
rect 343 2054 347 2058
rect 415 2054 419 2058
rect 495 2054 499 2058
rect 583 2054 587 2058
rect 671 2054 675 2058
rect 751 2054 755 2058
rect 831 2054 835 2058
rect 903 2054 907 2058
rect 983 2054 987 2058
rect 1063 2054 1067 2058
rect 1143 2054 1147 2058
rect 1447 2054 1451 2058
rect 1551 2054 1555 2058
rect 1663 2054 1667 2058
rect 1775 2054 1779 2058
rect 1879 2054 1883 2058
rect 1983 2054 1987 2058
rect 2087 2054 2091 2058
rect 2191 2054 2195 2058
rect 2287 2054 2291 2058
rect 2375 2054 2379 2058
rect 2471 2054 2475 2058
rect 2543 2054 2547 2058
rect 259 2047 260 2051
rect 260 2047 263 2051
rect 319 2047 320 2051
rect 320 2047 323 2051
rect 391 2047 392 2051
rect 392 2047 395 2051
rect 471 2047 472 2051
rect 472 2047 475 2051
rect 559 2047 560 2051
rect 560 2047 563 2051
rect 647 2047 648 2051
rect 648 2047 651 2051
rect 807 2047 808 2051
rect 808 2047 811 2051
rect 879 2047 880 2051
rect 880 2047 883 2051
rect 959 2047 960 2051
rect 960 2047 963 2051
rect 1039 2047 1040 2051
rect 1040 2047 1043 2051
rect 1119 2047 1120 2051
rect 1120 2047 1123 2051
rect 1427 2047 1428 2051
rect 1428 2047 1431 2051
rect 1527 2047 1528 2051
rect 1528 2047 1531 2051
rect 1639 2047 1640 2051
rect 1640 2047 1643 2051
rect 1855 2047 1856 2051
rect 1856 2047 1859 2051
rect 2055 2047 2059 2051
rect 2063 2047 2064 2051
rect 2064 2047 2067 2051
rect 2167 2047 2168 2051
rect 2168 2047 2171 2051
rect 2263 2047 2264 2051
rect 2264 2047 2267 2051
rect 2431 2047 2435 2051
rect 2479 2047 2483 2051
rect 2559 2047 2563 2051
rect 679 2035 683 2039
rect 1047 2039 1051 2043
rect 1391 2035 1392 2039
rect 1392 2035 1395 2039
rect 1495 2035 1499 2039
rect 1523 2035 1527 2039
rect 1687 2035 1688 2039
rect 1688 2035 1691 2039
rect 1787 2035 1788 2039
rect 1788 2035 1791 2039
rect 1895 2035 1899 2039
rect 1919 2035 1923 2039
rect 2131 2035 2135 2039
rect 2235 2035 2239 2039
rect 2423 2035 2424 2039
rect 2424 2035 2427 2039
rect 547 2027 551 2031
rect 603 2027 607 2031
rect 659 2027 663 2031
rect 743 2027 747 2031
rect 1415 2030 1419 2034
rect 1503 2030 1507 2034
rect 1607 2030 1611 2034
rect 1711 2030 1715 2034
rect 1807 2030 1811 2034
rect 1903 2030 1907 2034
rect 2007 2030 2011 2034
rect 2111 2030 2115 2034
rect 2215 2030 2219 2034
rect 2327 2030 2331 2034
rect 2447 2030 2451 2034
rect 2543 2030 2547 2034
rect 415 2022 419 2026
rect 471 2022 475 2026
rect 527 2022 531 2026
rect 583 2022 587 2026
rect 639 2022 643 2026
rect 695 2022 699 2026
rect 751 2022 755 2026
rect 807 2022 811 2026
rect 863 2022 867 2026
rect 919 2022 923 2026
rect 975 2022 979 2026
rect 1031 2022 1035 2026
rect 1367 2021 1371 2025
rect 2583 2021 2587 2025
rect 111 2013 115 2017
rect 1327 2013 1331 2017
rect 1391 2011 1395 2015
rect 1367 2004 1371 2008
rect 1399 2003 1403 2007
rect 111 1996 115 2000
rect 399 1995 403 1999
rect 455 1995 459 1999
rect 511 1995 515 1999
rect 547 1991 548 1995
rect 548 1991 551 1995
rect 567 1995 571 1999
rect 603 1991 604 1995
rect 604 1991 607 1995
rect 623 1995 627 1999
rect 659 1991 660 1995
rect 660 1991 663 1995
rect 679 1995 683 1999
rect 591 1983 595 1987
rect 735 1995 739 1999
rect 791 1995 795 1999
rect 847 1995 851 1999
rect 903 1995 907 1999
rect 959 1995 963 1999
rect 1015 1995 1019 1999
rect 1327 1996 1331 2000
rect 1427 1999 1431 2003
rect 1487 2003 1491 2007
rect 1523 1999 1524 2003
rect 1524 1999 1527 2003
rect 1591 2003 1595 2007
rect 1687 2011 1691 2015
rect 1695 2003 1699 2007
rect 1759 1999 1763 2003
rect 1791 2003 1795 2007
rect 2055 2011 2059 2015
rect 1887 2003 1891 2007
rect 1919 1999 1920 2003
rect 1920 1999 1923 2003
rect 1991 2003 1995 2007
rect 2095 2003 2099 2007
rect 2131 1999 2132 2003
rect 2132 1999 2135 2003
rect 2199 2003 2203 2007
rect 2235 1999 2236 2003
rect 2236 1999 2239 2003
rect 2311 2003 2315 2007
rect 2431 2003 2435 2007
rect 2527 2003 2531 2007
rect 2583 2004 2587 2008
rect 2559 1999 2560 2003
rect 2560 1999 2563 2003
rect 1047 1991 1048 1995
rect 1048 1991 1051 1995
rect 359 1967 363 1971
rect 1367 1968 1371 1972
rect 1399 1969 1403 1973
rect 1471 1971 1475 1975
rect 1495 1975 1499 1979
rect 1607 1979 1611 1983
rect 1479 1969 1483 1973
rect 1583 1969 1587 1973
rect 1671 1971 1675 1975
rect 1679 1969 1683 1973
rect 1707 1971 1711 1975
rect 1895 1979 1899 1983
rect 1767 1969 1771 1973
rect 1847 1969 1851 1973
rect 1919 1971 1923 1975
rect 1927 1969 1931 1973
rect 1999 1971 2003 1975
rect 2007 1969 2011 1973
rect 2079 1971 2083 1975
rect 2087 1969 2091 1973
rect 2583 1968 2587 1972
rect 111 1956 115 1960
rect 335 1957 339 1961
rect 383 1959 387 1963
rect 391 1957 395 1961
rect 439 1959 443 1963
rect 447 1957 451 1961
rect 495 1959 499 1963
rect 503 1957 507 1961
rect 567 1957 571 1961
rect 647 1957 651 1961
rect 735 1959 739 1963
rect 743 1957 747 1961
rect 855 1959 859 1963
rect 863 1957 867 1961
rect 991 1959 995 1963
rect 999 1957 1003 1961
rect 1135 1959 1139 1963
rect 1143 1957 1147 1961
rect 1175 1959 1176 1963
rect 1176 1959 1179 1963
rect 1271 1957 1275 1961
rect 1327 1956 1331 1960
rect 1367 1951 1371 1955
rect 2583 1951 2587 1955
rect 111 1939 115 1943
rect 1327 1939 1331 1943
rect 1415 1942 1419 1946
rect 1495 1942 1499 1946
rect 1599 1942 1603 1946
rect 1695 1942 1699 1946
rect 1783 1942 1787 1946
rect 1863 1942 1867 1946
rect 1943 1942 1947 1946
rect 2023 1942 2027 1946
rect 2103 1942 2107 1946
rect 351 1930 355 1934
rect 407 1930 411 1934
rect 463 1930 467 1934
rect 519 1930 523 1934
rect 583 1930 587 1934
rect 663 1930 667 1934
rect 759 1930 763 1934
rect 879 1930 883 1934
rect 1015 1930 1019 1934
rect 1159 1930 1163 1934
rect 1471 1935 1472 1939
rect 1472 1935 1475 1939
rect 1607 1935 1611 1939
rect 1671 1935 1672 1939
rect 1672 1935 1675 1939
rect 1759 1935 1760 1939
rect 1760 1935 1763 1939
rect 1843 1935 1844 1939
rect 1844 1935 1847 1939
rect 1919 1935 1920 1939
rect 1920 1935 1923 1939
rect 1999 1935 2000 1939
rect 2000 1935 2003 1939
rect 2079 1935 2080 1939
rect 2080 1935 2083 1939
rect 1287 1930 1291 1934
rect 359 1923 363 1927
rect 383 1923 384 1927
rect 384 1923 387 1927
rect 439 1923 440 1927
rect 440 1923 443 1927
rect 591 1923 595 1927
rect 671 1923 675 1927
rect 735 1923 736 1927
rect 736 1923 739 1927
rect 855 1923 856 1927
rect 856 1923 859 1927
rect 991 1923 992 1927
rect 992 1923 995 1927
rect 1135 1923 1136 1927
rect 1136 1923 1139 1927
rect 1219 1923 1223 1927
rect 1707 1923 1711 1927
rect 1739 1919 1743 1923
rect 135 1911 136 1915
rect 136 1911 139 1915
rect 223 1911 227 1915
rect 303 1911 304 1915
rect 304 1911 307 1915
rect 423 1911 427 1915
rect 495 1911 499 1915
rect 631 1911 632 1915
rect 632 1911 635 1915
rect 847 1915 851 1919
rect 1807 1919 1808 1923
rect 1808 1919 1811 1923
rect 1959 1927 1963 1931
rect 2135 1927 2139 1931
rect 1919 1919 1920 1923
rect 1920 1919 1923 1923
rect 2031 1919 2032 1923
rect 2032 1919 2035 1923
rect 855 1911 856 1915
rect 856 1911 859 1915
rect 975 1911 979 1915
rect 1063 1911 1064 1915
rect 1064 1911 1067 1915
rect 1107 1911 1111 1915
rect 1279 1911 1283 1915
rect 1719 1914 1723 1918
rect 1775 1914 1779 1918
rect 1831 1914 1835 1918
rect 1887 1914 1891 1918
rect 1943 1914 1947 1918
rect 1999 1914 2003 1918
rect 2055 1914 2059 1918
rect 2119 1914 2123 1918
rect 159 1906 163 1910
rect 231 1906 235 1910
rect 327 1906 331 1910
rect 431 1906 435 1910
rect 543 1906 547 1910
rect 655 1906 659 1910
rect 767 1906 771 1910
rect 879 1906 883 1910
rect 983 1906 987 1910
rect 1087 1906 1091 1910
rect 1199 1906 1203 1910
rect 1287 1906 1291 1910
rect 1367 1905 1371 1909
rect 2583 1905 2587 1909
rect 111 1897 115 1901
rect 1327 1897 1331 1901
rect 1807 1895 1811 1899
rect 135 1887 139 1891
rect 111 1880 115 1884
rect 143 1879 147 1883
rect 167 1875 171 1879
rect 215 1879 219 1883
rect 303 1887 307 1891
rect 311 1879 315 1883
rect 223 1867 227 1871
rect 415 1879 419 1883
rect 631 1887 635 1891
rect 527 1879 531 1883
rect 423 1867 427 1871
rect 639 1879 643 1883
rect 671 1875 672 1879
rect 672 1875 675 1879
rect 751 1879 755 1883
rect 855 1887 859 1891
rect 863 1879 867 1883
rect 847 1871 851 1875
rect 967 1879 971 1883
rect 1063 1887 1067 1891
rect 1071 1879 1075 1883
rect 1107 1875 1108 1879
rect 1108 1875 1111 1879
rect 1183 1879 1187 1883
rect 1219 1875 1220 1879
rect 1220 1875 1223 1879
rect 1271 1879 1275 1883
rect 1367 1888 1371 1892
rect 1703 1887 1707 1891
rect 1327 1880 1331 1884
rect 1739 1883 1740 1887
rect 1740 1883 1743 1887
rect 1759 1887 1763 1891
rect 1783 1883 1787 1887
rect 1815 1887 1819 1891
rect 1843 1883 1847 1887
rect 1871 1887 1875 1891
rect 1919 1895 1923 1899
rect 1927 1887 1931 1891
rect 1959 1883 1960 1887
rect 1960 1883 1963 1887
rect 1983 1887 1987 1891
rect 2039 1887 2043 1891
rect 2103 1887 2107 1891
rect 2583 1888 2587 1892
rect 2135 1883 2136 1887
rect 2136 1883 2139 1887
rect 1279 1855 1283 1859
rect 975 1847 979 1851
rect 111 1836 115 1840
rect 143 1837 147 1841
rect 191 1839 195 1843
rect 199 1837 203 1841
rect 255 1839 259 1843
rect 263 1837 267 1841
rect 343 1839 347 1843
rect 351 1837 355 1841
rect 431 1839 435 1843
rect 439 1837 443 1841
rect 527 1839 531 1843
rect 535 1837 539 1841
rect 559 1839 563 1843
rect 623 1837 627 1841
rect 703 1839 707 1843
rect 711 1837 715 1841
rect 783 1839 787 1843
rect 791 1837 795 1841
rect 863 1839 867 1843
rect 871 1837 875 1841
rect 943 1839 947 1843
rect 951 1837 955 1841
rect 1031 1839 1035 1843
rect 1367 1848 1371 1852
rect 1399 1849 1403 1853
rect 1463 1849 1467 1853
rect 1559 1849 1563 1853
rect 1655 1849 1659 1853
rect 1715 1855 1719 1859
rect 1743 1849 1747 1853
rect 1831 1849 1835 1853
rect 1911 1851 1915 1855
rect 1919 1849 1923 1853
rect 1999 1851 2003 1855
rect 2007 1849 2011 1853
rect 2031 1851 2035 1855
rect 2095 1849 2099 1853
rect 2175 1851 2179 1855
rect 2183 1849 2187 1853
rect 2207 1851 2211 1855
rect 2583 1848 2587 1852
rect 1039 1837 1043 1841
rect 1327 1836 1331 1840
rect 1367 1831 1371 1835
rect 2583 1831 2587 1835
rect 111 1819 115 1823
rect 1327 1819 1331 1823
rect 1415 1822 1419 1826
rect 1479 1822 1483 1826
rect 1575 1822 1579 1826
rect 1671 1822 1675 1826
rect 1759 1822 1763 1826
rect 1847 1822 1851 1826
rect 1935 1822 1939 1826
rect 2023 1822 2027 1826
rect 2111 1822 2115 1826
rect 2199 1822 2203 1826
rect 159 1810 163 1814
rect 215 1810 219 1814
rect 279 1810 283 1814
rect 367 1810 371 1814
rect 455 1810 459 1814
rect 551 1810 555 1814
rect 639 1810 643 1814
rect 727 1810 731 1814
rect 807 1810 811 1814
rect 887 1810 891 1814
rect 967 1810 971 1814
rect 1643 1815 1647 1819
rect 1783 1815 1787 1819
rect 1827 1815 1828 1819
rect 1828 1815 1831 1819
rect 1911 1815 1912 1819
rect 1912 1815 1915 1819
rect 1999 1815 2000 1819
rect 2000 1815 2003 1819
rect 2083 1815 2087 1819
rect 2175 1815 2176 1819
rect 2176 1815 2179 1819
rect 1055 1810 1059 1814
rect 167 1803 171 1807
rect 191 1803 192 1807
rect 192 1803 195 1807
rect 255 1803 256 1807
rect 256 1803 259 1807
rect 343 1803 344 1807
rect 344 1803 347 1807
rect 431 1803 432 1807
rect 432 1803 435 1807
rect 527 1803 528 1807
rect 528 1803 531 1807
rect 631 1803 635 1807
rect 703 1803 704 1807
rect 704 1803 707 1807
rect 783 1803 784 1807
rect 784 1803 787 1807
rect 863 1803 864 1807
rect 864 1803 867 1807
rect 959 1803 963 1807
rect 1031 1803 1032 1807
rect 1032 1803 1035 1807
rect 1407 1803 1411 1807
rect 1435 1803 1439 1807
rect 1531 1803 1535 1807
rect 1715 1803 1716 1807
rect 1716 1803 1719 1807
rect 1927 1803 1928 1807
rect 1928 1803 1931 1807
rect 1971 1803 1975 1807
rect 2155 1803 2159 1807
rect 2235 1803 2239 1807
rect 2323 1803 2327 1807
rect 2535 1803 2539 1807
rect 559 1795 563 1799
rect 1415 1798 1419 1802
rect 1511 1798 1515 1802
rect 1623 1798 1627 1802
rect 1735 1798 1739 1802
rect 1839 1798 1843 1802
rect 1951 1798 1955 1802
rect 2063 1798 2067 1802
rect 2183 1798 2187 1802
rect 2303 1798 2307 1802
rect 2431 1798 2435 1802
rect 2543 1798 2547 1802
rect 251 1787 255 1791
rect 315 1787 319 1791
rect 387 1787 391 1791
rect 467 1787 471 1791
rect 599 1787 600 1791
rect 600 1787 603 1791
rect 231 1782 235 1786
rect 295 1782 299 1786
rect 367 1782 371 1786
rect 447 1782 451 1786
rect 535 1782 539 1786
rect 623 1782 627 1786
rect 711 1782 715 1786
rect 727 1783 731 1787
rect 863 1787 867 1791
rect 911 1787 915 1791
rect 943 1791 947 1795
rect 1367 1789 1371 1793
rect 2583 1789 2587 1793
rect 791 1782 795 1786
rect 871 1782 875 1786
rect 951 1782 955 1786
rect 1031 1782 1035 1786
rect 1119 1782 1123 1786
rect 1927 1779 1931 1783
rect 111 1773 115 1777
rect 1327 1773 1331 1777
rect 1367 1772 1371 1776
rect 1399 1771 1403 1775
rect 599 1763 603 1767
rect 1435 1767 1436 1771
rect 1436 1767 1439 1771
rect 1495 1771 1499 1775
rect 1531 1767 1532 1771
rect 1532 1767 1535 1771
rect 1607 1771 1611 1775
rect 1643 1767 1644 1771
rect 1644 1767 1647 1771
rect 1719 1771 1723 1775
rect 1823 1771 1827 1775
rect 1919 1767 1923 1771
rect 1935 1771 1939 1775
rect 1971 1767 1972 1771
rect 1972 1767 1975 1771
rect 2047 1771 2051 1775
rect 2083 1767 2084 1771
rect 2084 1767 2087 1771
rect 2167 1771 2171 1775
rect 2235 1767 2239 1771
rect 2287 1771 2291 1775
rect 2323 1767 2324 1771
rect 2324 1767 2327 1771
rect 2415 1771 2419 1775
rect 2527 1771 2531 1775
rect 2583 1772 2587 1776
rect 111 1756 115 1760
rect 215 1755 219 1759
rect 251 1751 252 1755
rect 252 1751 255 1755
rect 279 1755 283 1759
rect 315 1751 316 1755
rect 316 1751 319 1755
rect 351 1755 355 1759
rect 387 1751 388 1755
rect 388 1751 391 1755
rect 431 1755 435 1759
rect 467 1751 468 1755
rect 468 1751 471 1755
rect 519 1755 523 1759
rect 359 1743 363 1747
rect 607 1755 611 1759
rect 631 1751 635 1755
rect 695 1755 699 1759
rect 727 1751 728 1755
rect 728 1751 731 1755
rect 775 1755 779 1759
rect 2471 1763 2475 1767
rect 855 1755 859 1759
rect 911 1755 915 1759
rect 935 1755 939 1759
rect 959 1751 963 1755
rect 1015 1755 1019 1759
rect 1103 1755 1107 1759
rect 1327 1756 1331 1760
rect 1407 1743 1411 1747
rect 1367 1736 1371 1740
rect 1439 1737 1443 1741
rect 1519 1737 1523 1741
rect 1615 1737 1619 1741
rect 1719 1737 1723 1741
rect 1775 1743 1779 1747
rect 1823 1737 1827 1741
rect 1927 1737 1931 1741
rect 2023 1737 2027 1741
rect 2111 1739 2115 1743
rect 2119 1737 2123 1741
rect 2155 1739 2156 1743
rect 2156 1739 2159 1743
rect 2207 1737 2211 1741
rect 2279 1739 2283 1743
rect 2287 1737 2291 1741
rect 2367 1739 2371 1743
rect 2375 1737 2379 1741
rect 2399 1739 2403 1743
rect 2463 1737 2467 1741
rect 2495 1739 2496 1743
rect 2496 1739 2499 1743
rect 2535 1743 2539 1747
rect 2527 1737 2531 1741
rect 2583 1736 2587 1740
rect 111 1716 115 1720
rect 351 1717 355 1721
rect 399 1719 403 1723
rect 407 1717 411 1721
rect 463 1719 467 1723
rect 471 1717 475 1721
rect 543 1719 547 1723
rect 551 1717 555 1721
rect 583 1719 584 1723
rect 584 1719 587 1723
rect 639 1717 643 1721
rect 727 1717 731 1721
rect 863 1727 867 1731
rect 823 1717 827 1721
rect 919 1717 923 1721
rect 1015 1717 1019 1721
rect 1103 1719 1107 1723
rect 1111 1717 1115 1721
rect 1199 1719 1203 1723
rect 1207 1717 1211 1721
rect 1231 1719 1235 1723
rect 1327 1716 1331 1720
rect 1367 1719 1371 1723
rect 2583 1719 2587 1723
rect 1455 1710 1459 1714
rect 1535 1710 1539 1714
rect 1631 1710 1635 1714
rect 1735 1710 1739 1714
rect 1839 1710 1843 1714
rect 1943 1710 1947 1714
rect 2039 1710 2043 1714
rect 2135 1710 2139 1714
rect 2223 1710 2227 1714
rect 2303 1710 2307 1714
rect 2391 1710 2395 1714
rect 2479 1710 2483 1714
rect 2543 1710 2547 1714
rect 111 1699 115 1703
rect 1327 1699 1331 1703
rect 1723 1703 1727 1707
rect 1919 1703 1920 1707
rect 1920 1703 1923 1707
rect 2019 1703 2020 1707
rect 2020 1703 2023 1707
rect 2111 1703 2112 1707
rect 2112 1703 2115 1707
rect 2231 1703 2235 1707
rect 2279 1703 2280 1707
rect 2280 1703 2283 1707
rect 2367 1703 2368 1707
rect 2368 1703 2371 1707
rect 2471 1703 2475 1707
rect 2559 1703 2563 1707
rect 367 1690 371 1694
rect 423 1690 427 1694
rect 487 1690 491 1694
rect 567 1690 571 1694
rect 655 1690 659 1694
rect 743 1690 747 1694
rect 839 1690 843 1694
rect 935 1690 939 1694
rect 1031 1690 1035 1694
rect 1127 1690 1131 1694
rect 1223 1690 1227 1694
rect 359 1683 363 1687
rect 399 1683 400 1687
rect 400 1683 403 1687
rect 463 1683 464 1687
rect 464 1683 467 1687
rect 543 1683 544 1687
rect 544 1683 547 1687
rect 819 1683 820 1687
rect 820 1683 823 1687
rect 983 1683 987 1687
rect 1103 1683 1104 1687
rect 1104 1683 1107 1687
rect 1199 1683 1200 1687
rect 1200 1683 1203 1687
rect 583 1675 587 1679
rect 1551 1679 1555 1683
rect 1579 1679 1583 1683
rect 1651 1679 1655 1683
rect 1775 1679 1776 1683
rect 1776 1679 1779 1683
rect 1819 1679 1823 1683
rect 1903 1679 1907 1683
rect 2295 1687 2299 1691
rect 2083 1679 2087 1683
rect 2163 1679 2167 1683
rect 2263 1679 2264 1683
rect 2264 1679 2267 1683
rect 2435 1687 2439 1691
rect 2399 1679 2400 1683
rect 2400 1679 2403 1683
rect 2495 1683 2499 1687
rect 2535 1679 2539 1683
rect 471 1667 475 1671
rect 531 1667 535 1671
rect 595 1667 599 1671
rect 667 1667 671 1671
rect 767 1667 771 1671
rect 855 1667 859 1671
rect 1023 1667 1024 1671
rect 1024 1667 1027 1671
rect 1067 1667 1071 1671
rect 1231 1671 1235 1675
rect 1559 1674 1563 1678
rect 1631 1674 1635 1678
rect 1711 1674 1715 1678
rect 1799 1674 1803 1678
rect 1887 1674 1891 1678
rect 1975 1674 1979 1678
rect 2063 1674 2067 1678
rect 2143 1674 2147 1678
rect 2215 1674 2219 1678
rect 2287 1674 2291 1678
rect 2351 1674 2355 1678
rect 2423 1674 2427 1678
rect 2487 1674 2491 1678
rect 2543 1674 2547 1678
rect 1243 1667 1247 1671
rect 399 1662 403 1666
rect 455 1662 459 1666
rect 511 1662 515 1666
rect 575 1662 579 1666
rect 647 1662 651 1666
rect 727 1662 731 1666
rect 807 1662 811 1666
rect 887 1662 891 1666
rect 967 1662 971 1666
rect 1047 1662 1051 1666
rect 1135 1662 1139 1666
rect 1223 1662 1227 1666
rect 1287 1662 1291 1666
rect 1367 1665 1371 1669
rect 2583 1665 2587 1669
rect 111 1653 115 1657
rect 1327 1653 1331 1657
rect 2263 1655 2267 1659
rect 1367 1648 1371 1652
rect 1543 1647 1547 1651
rect 1023 1643 1027 1647
rect 111 1636 115 1640
rect 383 1635 387 1639
rect 439 1635 443 1639
rect 471 1631 472 1635
rect 472 1631 475 1635
rect 495 1635 499 1639
rect 531 1631 532 1635
rect 532 1631 535 1635
rect 559 1635 563 1639
rect 595 1631 596 1635
rect 596 1631 599 1635
rect 631 1635 635 1639
rect 667 1631 668 1635
rect 668 1631 671 1635
rect 711 1635 715 1639
rect 767 1635 771 1639
rect 791 1635 795 1639
rect 819 1631 823 1635
rect 871 1635 875 1639
rect 951 1635 955 1639
rect 983 1631 984 1635
rect 984 1631 987 1635
rect 1031 1635 1035 1639
rect 1067 1631 1068 1635
rect 1068 1631 1071 1635
rect 1119 1635 1123 1639
rect 1143 1631 1147 1635
rect 1207 1635 1211 1639
rect 1243 1631 1244 1635
rect 1244 1631 1247 1635
rect 1271 1635 1275 1639
rect 1579 1643 1580 1647
rect 1580 1643 1583 1647
rect 1615 1647 1619 1651
rect 1651 1643 1652 1647
rect 1652 1643 1655 1647
rect 1695 1647 1699 1651
rect 1723 1643 1727 1647
rect 1783 1647 1787 1651
rect 1819 1643 1820 1647
rect 1820 1643 1823 1647
rect 1871 1647 1875 1651
rect 1903 1643 1904 1647
rect 1904 1643 1907 1647
rect 1959 1647 1963 1651
rect 1983 1643 1987 1647
rect 2047 1647 2051 1651
rect 2083 1643 2084 1647
rect 2084 1643 2087 1647
rect 2127 1647 2131 1651
rect 2163 1643 2164 1647
rect 2164 1643 2167 1647
rect 2199 1647 2203 1651
rect 2231 1643 2232 1647
rect 2232 1643 2235 1647
rect 2271 1647 2275 1651
rect 2295 1643 2299 1647
rect 2335 1647 2339 1651
rect 2399 1655 2403 1659
rect 2407 1647 2411 1651
rect 2435 1643 2439 1647
rect 2471 1647 2475 1651
rect 2527 1647 2531 1651
rect 2583 1648 2587 1652
rect 2559 1643 2560 1647
rect 2560 1643 2563 1647
rect 1327 1636 1331 1640
rect 1551 1607 1555 1611
rect 1367 1600 1371 1604
rect 1575 1601 1579 1605
rect 1631 1601 1635 1605
rect 1687 1601 1691 1605
rect 1751 1601 1755 1605
rect 1831 1601 1835 1605
rect 1919 1601 1923 1605
rect 1999 1603 2003 1607
rect 2007 1601 2011 1605
rect 2095 1603 2099 1607
rect 2103 1601 2107 1605
rect 2127 1603 2131 1607
rect 2207 1601 2211 1605
rect 2311 1603 2315 1607
rect 2319 1601 2323 1605
rect 2423 1603 2427 1607
rect 2431 1601 2435 1605
rect 2463 1603 2464 1607
rect 2464 1603 2467 1607
rect 2535 1607 2539 1611
rect 2527 1601 2531 1605
rect 2583 1600 2587 1604
rect 911 1595 915 1599
rect 111 1584 115 1588
rect 287 1585 291 1589
rect 359 1587 363 1591
rect 367 1585 371 1589
rect 447 1587 451 1591
rect 455 1585 459 1589
rect 535 1587 539 1591
rect 551 1585 555 1589
rect 639 1587 643 1591
rect 647 1585 651 1589
rect 671 1587 675 1591
rect 735 1585 739 1589
rect 815 1587 819 1591
rect 823 1585 827 1589
rect 855 1587 856 1591
rect 856 1587 859 1591
rect 903 1585 907 1589
rect 983 1585 987 1589
rect 1031 1587 1035 1591
rect 1063 1585 1067 1589
rect 1151 1585 1155 1589
rect 1327 1584 1331 1588
rect 1367 1583 1371 1587
rect 2583 1583 2587 1587
rect 1591 1574 1595 1578
rect 1647 1574 1651 1578
rect 1703 1574 1707 1578
rect 1767 1574 1771 1578
rect 1847 1574 1851 1578
rect 1935 1574 1939 1578
rect 2023 1574 2027 1578
rect 2119 1574 2123 1578
rect 2223 1574 2227 1578
rect 2335 1574 2339 1578
rect 2447 1574 2451 1578
rect 2543 1574 2547 1578
rect 111 1567 115 1571
rect 1327 1567 1331 1571
rect 1903 1567 1907 1571
rect 1983 1567 1987 1571
rect 1999 1567 2000 1571
rect 2000 1567 2003 1571
rect 2095 1567 2096 1571
rect 2096 1567 2099 1571
rect 2311 1567 2312 1571
rect 2312 1567 2315 1571
rect 2423 1567 2424 1571
rect 2424 1567 2427 1571
rect 2559 1567 2563 1571
rect 303 1558 307 1562
rect 383 1558 387 1562
rect 471 1558 475 1562
rect 567 1558 571 1562
rect 663 1558 667 1562
rect 751 1558 755 1562
rect 839 1558 843 1562
rect 919 1558 923 1562
rect 999 1558 1003 1562
rect 1079 1558 1083 1562
rect 1167 1558 1171 1562
rect 295 1551 299 1555
rect 359 1551 360 1555
rect 360 1551 363 1555
rect 415 1547 419 1551
rect 447 1551 448 1555
rect 448 1551 451 1555
rect 535 1551 539 1555
rect 639 1551 640 1555
rect 640 1551 643 1555
rect 671 1547 675 1551
rect 707 1551 711 1555
rect 815 1551 816 1555
rect 816 1551 819 1555
rect 911 1551 915 1555
rect 1143 1551 1144 1555
rect 1144 1551 1147 1555
rect 1671 1551 1675 1555
rect 1755 1551 1759 1555
rect 1811 1551 1815 1555
rect 1875 1551 1879 1555
rect 1947 1551 1951 1555
rect 2127 1555 2131 1559
rect 2343 1559 2347 1563
rect 2143 1551 2144 1555
rect 2144 1551 2147 1555
rect 2267 1551 2271 1555
rect 2383 1551 2384 1555
rect 2384 1551 2387 1555
rect 2463 1551 2464 1555
rect 2464 1551 2467 1555
rect 2535 1551 2539 1555
rect 1679 1546 1683 1550
rect 1735 1546 1739 1550
rect 1791 1546 1795 1550
rect 1855 1546 1859 1550
rect 1927 1546 1931 1550
rect 2007 1546 2011 1550
rect 2087 1546 2091 1550
rect 2167 1546 2171 1550
rect 2247 1546 2251 1550
rect 2327 1546 2331 1550
rect 2407 1546 2411 1550
rect 2487 1546 2491 1550
rect 2543 1546 2547 1550
rect 255 1539 256 1543
rect 256 1539 259 1543
rect 391 1539 395 1543
rect 447 1539 448 1543
rect 448 1539 451 1543
rect 491 1539 495 1543
rect 679 1539 683 1543
rect 735 1539 736 1543
rect 736 1539 739 1543
rect 807 1539 808 1543
rect 808 1539 811 1543
rect 879 1539 880 1543
rect 880 1539 883 1543
rect 967 1539 971 1543
rect 1031 1539 1032 1543
rect 1032 1539 1035 1543
rect 279 1534 283 1538
rect 335 1534 339 1538
rect 399 1534 403 1538
rect 471 1534 475 1538
rect 543 1534 547 1538
rect 615 1534 619 1538
rect 687 1534 691 1538
rect 759 1534 763 1538
rect 831 1534 835 1538
rect 903 1534 907 1538
rect 975 1534 979 1538
rect 1055 1534 1059 1538
rect 1367 1537 1371 1541
rect 2583 1537 2587 1541
rect 111 1525 115 1529
rect 1327 1525 1331 1529
rect 1903 1527 1907 1531
rect 1367 1520 1371 1524
rect 255 1515 259 1519
rect 111 1508 115 1512
rect 263 1507 267 1511
rect 295 1503 296 1507
rect 296 1503 299 1507
rect 319 1507 323 1511
rect 447 1515 451 1519
rect 383 1507 387 1511
rect 415 1503 416 1507
rect 416 1503 419 1507
rect 455 1507 459 1511
rect 491 1503 492 1507
rect 492 1503 495 1507
rect 527 1507 531 1511
rect 575 1503 579 1507
rect 599 1507 603 1511
rect 735 1515 739 1519
rect 1663 1519 1667 1523
rect 671 1507 675 1511
rect 707 1503 708 1507
rect 708 1503 711 1507
rect 743 1507 747 1511
rect 679 1495 683 1499
rect 815 1507 819 1511
rect 879 1515 883 1519
rect 887 1507 891 1511
rect 911 1503 915 1507
rect 959 1507 963 1511
rect 1719 1519 1723 1523
rect 1755 1515 1756 1519
rect 1756 1515 1759 1519
rect 1775 1519 1779 1523
rect 1811 1515 1812 1519
rect 1812 1515 1815 1519
rect 1839 1519 1843 1523
rect 1875 1515 1876 1519
rect 1876 1515 1879 1519
rect 1911 1519 1915 1523
rect 1947 1515 1948 1519
rect 1948 1515 1951 1519
rect 1991 1519 1995 1523
rect 2143 1527 2147 1531
rect 2071 1519 2075 1523
rect 1039 1507 1043 1511
rect 1327 1508 1331 1512
rect 2035 1511 2039 1515
rect 2151 1519 2155 1523
rect 2231 1519 2235 1523
rect 2383 1527 2387 1531
rect 2311 1519 2315 1523
rect 2343 1515 2344 1519
rect 2344 1515 2347 1519
rect 2391 1519 2395 1523
rect 2415 1515 2419 1519
rect 2471 1519 2475 1523
rect 2527 1519 2531 1523
rect 2583 1520 2587 1524
rect 2559 1515 2560 1519
rect 2560 1515 2563 1519
rect 967 1495 971 1499
rect 1671 1487 1675 1491
rect 111 1468 115 1472
rect 199 1469 203 1473
rect 279 1471 283 1475
rect 287 1469 291 1473
rect 375 1471 379 1475
rect 391 1475 395 1479
rect 383 1469 387 1473
rect 487 1469 491 1473
rect 511 1471 515 1475
rect 1367 1476 1371 1480
rect 1519 1477 1523 1481
rect 1567 1479 1571 1483
rect 1575 1477 1579 1481
rect 1639 1479 1643 1483
rect 1647 1477 1651 1481
rect 1719 1479 1723 1483
rect 1727 1477 1731 1481
rect 1799 1479 1803 1483
rect 1807 1477 1811 1481
rect 1887 1479 1891 1483
rect 1895 1477 1899 1481
rect 1983 1477 1987 1481
rect 2007 1479 2011 1483
rect 2071 1477 2075 1481
rect 2143 1479 2147 1483
rect 2151 1477 2155 1481
rect 2223 1479 2227 1483
rect 2231 1477 2235 1481
rect 2267 1479 2268 1483
rect 2268 1479 2271 1483
rect 2283 1483 2287 1487
rect 2311 1477 2315 1481
rect 2355 1483 2359 1487
rect 2391 1477 2395 1481
rect 2471 1477 2475 1481
rect 2519 1479 2523 1483
rect 2535 1483 2539 1487
rect 2527 1477 2531 1481
rect 2583 1476 2587 1480
rect 583 1469 587 1473
rect 679 1469 683 1473
rect 767 1471 771 1475
rect 775 1469 779 1473
rect 807 1471 808 1475
rect 808 1471 811 1475
rect 863 1469 867 1473
rect 943 1471 947 1475
rect 951 1469 955 1473
rect 1031 1471 1035 1475
rect 1039 1469 1043 1473
rect 1127 1471 1131 1475
rect 1135 1469 1139 1473
rect 1191 1471 1195 1475
rect 1327 1468 1331 1472
rect 1367 1459 1371 1463
rect 2583 1459 2587 1463
rect 111 1451 115 1455
rect 1327 1451 1331 1455
rect 1535 1450 1539 1454
rect 1591 1450 1595 1454
rect 1663 1450 1667 1454
rect 1743 1450 1747 1454
rect 1823 1450 1827 1454
rect 1911 1450 1915 1454
rect 1999 1450 2003 1454
rect 2087 1450 2091 1454
rect 2167 1450 2171 1454
rect 2247 1450 2251 1454
rect 2327 1450 2331 1454
rect 2407 1450 2411 1454
rect 2487 1450 2491 1454
rect 2543 1450 2547 1454
rect 215 1442 219 1446
rect 303 1442 307 1446
rect 399 1442 403 1446
rect 503 1442 507 1446
rect 599 1442 603 1446
rect 695 1442 699 1446
rect 791 1442 795 1446
rect 879 1442 883 1446
rect 967 1442 971 1446
rect 1055 1442 1059 1446
rect 1151 1442 1155 1446
rect 175 1435 179 1439
rect 279 1435 280 1439
rect 280 1435 283 1439
rect 375 1435 376 1439
rect 376 1435 379 1439
rect 575 1435 576 1439
rect 576 1435 579 1439
rect 759 1435 763 1439
rect 767 1435 768 1439
rect 768 1435 771 1439
rect 911 1435 915 1439
rect 943 1435 944 1439
rect 944 1435 947 1439
rect 1031 1435 1032 1439
rect 1032 1435 1035 1439
rect 1127 1435 1128 1439
rect 1128 1435 1131 1439
rect 1567 1443 1568 1447
rect 1568 1443 1571 1447
rect 1639 1443 1640 1447
rect 1640 1443 1643 1447
rect 1719 1443 1720 1447
rect 1720 1443 1723 1447
rect 1799 1443 1800 1447
rect 1800 1443 1803 1447
rect 1887 1443 1888 1447
rect 1888 1443 1891 1447
rect 2035 1443 2039 1447
rect 2043 1443 2047 1447
rect 2143 1443 2144 1447
rect 2144 1443 2147 1447
rect 2223 1443 2224 1447
rect 2224 1443 2227 1447
rect 2355 1443 2359 1447
rect 2415 1443 2419 1447
rect 2519 1443 2520 1447
rect 2520 1443 2523 1447
rect 1839 1435 1843 1439
rect 135 1419 136 1423
rect 136 1419 139 1423
rect 359 1427 363 1431
rect 335 1419 339 1423
rect 511 1427 515 1431
rect 467 1419 471 1423
rect 571 1419 575 1423
rect 743 1419 744 1423
rect 744 1419 747 1423
rect 871 1419 875 1423
rect 1119 1427 1123 1431
rect 1079 1419 1080 1423
rect 1080 1419 1083 1423
rect 1191 1419 1192 1423
rect 1192 1419 1195 1423
rect 1407 1423 1411 1427
rect 1435 1423 1439 1427
rect 1503 1423 1507 1427
rect 1555 1423 1559 1427
rect 1643 1423 1647 1427
rect 2007 1431 2011 1435
rect 2135 1431 2139 1435
rect 2559 1435 2563 1439
rect 2095 1423 2096 1427
rect 2096 1423 2099 1427
rect 2239 1427 2243 1431
rect 2283 1423 2284 1427
rect 2284 1423 2287 1427
rect 2507 1423 2511 1427
rect 159 1414 163 1418
rect 247 1414 251 1418
rect 343 1414 347 1418
rect 447 1414 451 1418
rect 551 1414 555 1418
rect 663 1414 667 1418
rect 767 1414 771 1418
rect 879 1414 883 1418
rect 991 1414 995 1418
rect 1103 1414 1107 1418
rect 1215 1414 1219 1418
rect 1415 1418 1419 1422
rect 1471 1418 1475 1422
rect 1535 1418 1539 1422
rect 1623 1418 1627 1422
rect 1719 1418 1723 1422
rect 1823 1418 1827 1422
rect 1927 1418 1931 1422
rect 2023 1418 2027 1422
rect 2119 1418 2123 1422
rect 2215 1418 2219 1422
rect 2303 1418 2307 1422
rect 2391 1418 2395 1422
rect 2479 1418 2483 1422
rect 2543 1418 2547 1422
rect 111 1405 115 1409
rect 1327 1405 1331 1409
rect 1367 1409 1371 1413
rect 2583 1409 2587 1413
rect 135 1395 139 1399
rect 111 1388 115 1392
rect 143 1387 147 1391
rect 175 1383 176 1387
rect 176 1383 179 1387
rect 231 1387 235 1391
rect 743 1395 747 1399
rect 327 1387 331 1391
rect 359 1383 360 1387
rect 360 1383 363 1387
rect 431 1387 435 1391
rect 467 1383 468 1387
rect 468 1383 471 1387
rect 535 1387 539 1391
rect 571 1383 572 1387
rect 572 1383 575 1387
rect 647 1387 651 1391
rect 671 1383 675 1387
rect 751 1387 755 1391
rect 759 1379 763 1383
rect 863 1387 867 1391
rect 1079 1395 1083 1399
rect 2095 1399 2099 1403
rect 975 1387 979 1391
rect 999 1383 1003 1387
rect 1087 1387 1091 1391
rect 1119 1383 1120 1387
rect 1120 1383 1123 1387
rect 1199 1387 1203 1391
rect 1327 1388 1331 1392
rect 1367 1392 1371 1396
rect 1399 1391 1403 1395
rect 1435 1387 1436 1391
rect 1436 1387 1439 1391
rect 1455 1391 1459 1395
rect 1503 1387 1507 1391
rect 1519 1391 1523 1395
rect 1555 1387 1556 1391
rect 1556 1387 1559 1391
rect 1607 1391 1611 1395
rect 1643 1387 1644 1391
rect 1644 1387 1647 1391
rect 1703 1391 1707 1395
rect 1807 1391 1811 1395
rect 1839 1387 1840 1391
rect 1840 1387 1843 1391
rect 1911 1391 1915 1395
rect 1935 1387 1939 1391
rect 2007 1391 2011 1395
rect 2043 1387 2044 1391
rect 2044 1387 2047 1391
rect 2103 1391 2107 1395
rect 2135 1387 2136 1391
rect 2136 1387 2139 1391
rect 2199 1391 2203 1395
rect 2287 1391 2291 1395
rect 2375 1391 2379 1395
rect 2463 1391 2467 1395
rect 2507 1387 2511 1391
rect 2527 1391 2531 1395
rect 2583 1392 2587 1396
rect 2559 1387 2560 1391
rect 2560 1387 2563 1391
rect 335 1363 339 1367
rect 111 1352 115 1356
rect 143 1353 147 1357
rect 199 1355 203 1359
rect 207 1353 211 1357
rect 287 1355 291 1359
rect 295 1353 299 1357
rect 391 1355 395 1359
rect 399 1353 403 1357
rect 475 1359 479 1363
rect 511 1353 515 1357
rect 623 1353 627 1357
rect 735 1353 739 1357
rect 839 1355 843 1359
rect 847 1353 851 1357
rect 871 1355 875 1359
rect 959 1353 963 1357
rect 1063 1355 1067 1359
rect 1071 1353 1075 1357
rect 1175 1355 1179 1359
rect 1183 1353 1187 1357
rect 1263 1355 1267 1359
rect 1271 1353 1275 1357
rect 1295 1355 1299 1359
rect 1327 1352 1331 1356
rect 1367 1348 1371 1352
rect 1399 1349 1403 1353
rect 1447 1351 1451 1355
rect 1455 1349 1459 1353
rect 1535 1351 1539 1355
rect 1543 1349 1547 1353
rect 1623 1351 1627 1355
rect 1631 1349 1635 1353
rect 1711 1351 1715 1355
rect 1719 1349 1723 1353
rect 1751 1351 1752 1355
rect 1752 1351 1755 1355
rect 1807 1349 1811 1353
rect 1839 1351 1840 1355
rect 1840 1351 1843 1355
rect 1887 1349 1891 1353
rect 1967 1349 1971 1353
rect 2039 1351 2043 1355
rect 2047 1349 2051 1353
rect 2119 1351 2123 1355
rect 2127 1349 2131 1353
rect 2199 1351 2203 1355
rect 2207 1349 2211 1353
rect 2239 1351 2240 1355
rect 2240 1351 2243 1355
rect 2583 1348 2587 1352
rect 111 1335 115 1339
rect 1327 1335 1331 1339
rect 1367 1331 1371 1335
rect 159 1326 163 1330
rect 223 1326 227 1330
rect 311 1326 315 1330
rect 415 1326 419 1330
rect 527 1326 531 1330
rect 639 1326 643 1330
rect 751 1326 755 1330
rect 863 1326 867 1330
rect 975 1326 979 1330
rect 1087 1326 1091 1330
rect 1199 1326 1203 1330
rect 2583 1331 2587 1335
rect 1287 1326 1291 1330
rect 175 1319 179 1323
rect 199 1319 200 1323
rect 200 1319 203 1323
rect 287 1319 288 1323
rect 288 1319 291 1323
rect 343 1315 347 1319
rect 391 1319 392 1323
rect 392 1319 395 1323
rect 671 1319 675 1323
rect 743 1319 747 1323
rect 839 1319 840 1323
rect 840 1319 843 1323
rect 999 1319 1003 1323
rect 1063 1319 1064 1323
rect 1064 1319 1067 1323
rect 1175 1319 1176 1323
rect 1176 1319 1179 1323
rect 1263 1319 1264 1323
rect 1264 1319 1267 1323
rect 1415 1322 1419 1326
rect 1471 1322 1475 1326
rect 1559 1322 1563 1326
rect 1647 1322 1651 1326
rect 1735 1322 1739 1326
rect 1823 1322 1827 1326
rect 1903 1322 1907 1326
rect 1983 1322 1987 1326
rect 2063 1322 2067 1326
rect 2143 1322 2147 1326
rect 2223 1322 2227 1326
rect 135 1307 136 1311
rect 136 1307 139 1311
rect 303 1307 304 1311
rect 304 1307 307 1311
rect 475 1311 479 1315
rect 1307 1315 1311 1319
rect 1447 1315 1448 1319
rect 1448 1315 1451 1319
rect 1535 1315 1536 1319
rect 1536 1315 1539 1319
rect 1623 1315 1624 1319
rect 1624 1315 1627 1319
rect 1711 1315 1712 1319
rect 1712 1315 1715 1319
rect 1935 1315 1939 1319
rect 1975 1315 1979 1319
rect 2039 1315 2040 1319
rect 2040 1315 2043 1319
rect 2119 1315 2120 1319
rect 2120 1315 2123 1319
rect 2199 1315 2200 1319
rect 2200 1315 2203 1319
rect 483 1307 487 1311
rect 607 1307 608 1311
rect 608 1307 611 1311
rect 651 1307 655 1311
rect 779 1307 783 1311
rect 891 1307 892 1311
rect 892 1307 895 1311
rect 931 1307 935 1311
rect 1011 1307 1015 1311
rect 1111 1307 1115 1311
rect 1171 1307 1175 1311
rect 1251 1307 1255 1311
rect 159 1302 163 1306
rect 231 1302 235 1306
rect 327 1302 331 1306
rect 431 1302 435 1306
rect 535 1302 539 1306
rect 631 1302 635 1306
rect 727 1302 731 1306
rect 823 1302 827 1306
rect 911 1302 915 1306
rect 991 1302 995 1306
rect 1071 1302 1075 1306
rect 1151 1302 1155 1306
rect 1231 1302 1235 1306
rect 1287 1302 1291 1306
rect 1791 1303 1795 1307
rect 2055 1307 2059 1311
rect 1839 1299 1840 1303
rect 1840 1299 1843 1303
rect 2023 1299 2024 1303
rect 2024 1299 2027 1303
rect 2247 1307 2251 1311
rect 2187 1299 2191 1303
rect 111 1293 115 1297
rect 1327 1293 1331 1297
rect 1671 1294 1675 1298
rect 1767 1294 1771 1298
rect 1863 1294 1867 1298
rect 1959 1294 1963 1298
rect 2047 1294 2051 1298
rect 2135 1294 2139 1298
rect 2231 1294 2235 1298
rect 135 1283 139 1287
rect 111 1276 115 1280
rect 143 1275 147 1279
rect 175 1271 176 1275
rect 176 1271 179 1275
rect 215 1275 219 1279
rect 607 1283 611 1287
rect 1367 1285 1371 1289
rect 2583 1285 2587 1289
rect 311 1275 315 1279
rect 343 1271 344 1275
rect 344 1271 347 1275
rect 415 1275 419 1279
rect 483 1271 487 1275
rect 519 1275 523 1279
rect 543 1271 547 1275
rect 615 1275 619 1279
rect 651 1271 652 1275
rect 652 1271 655 1275
rect 711 1275 715 1279
rect 743 1271 744 1275
rect 744 1271 747 1275
rect 807 1275 811 1279
rect 895 1275 899 1279
rect 931 1271 932 1275
rect 932 1271 935 1275
rect 975 1275 979 1279
rect 1011 1271 1012 1275
rect 1012 1271 1015 1275
rect 1055 1275 1059 1279
rect 1111 1275 1115 1279
rect 1135 1275 1139 1279
rect 1171 1271 1172 1275
rect 1172 1271 1175 1275
rect 1215 1275 1219 1279
rect 1251 1271 1252 1275
rect 1252 1271 1255 1275
rect 1271 1275 1275 1279
rect 1327 1276 1331 1280
rect 2023 1275 2027 1279
rect 1307 1271 1308 1275
rect 1308 1271 1311 1275
rect 1367 1268 1371 1272
rect 1655 1267 1659 1271
rect 1663 1259 1667 1263
rect 1751 1267 1755 1271
rect 1847 1267 1851 1271
rect 1935 1263 1939 1267
rect 1943 1267 1947 1271
rect 1975 1263 1976 1267
rect 1976 1263 1979 1267
rect 2031 1267 2035 1271
rect 2055 1263 2059 1267
rect 2119 1267 2123 1271
rect 2215 1267 2219 1271
rect 2583 1268 2587 1272
rect 2247 1263 2248 1267
rect 2248 1263 2251 1267
rect 151 1239 155 1243
rect 111 1228 115 1232
rect 143 1229 147 1233
rect 191 1231 195 1235
rect 199 1229 203 1233
rect 271 1231 275 1235
rect 279 1229 283 1233
rect 303 1231 307 1235
rect 359 1229 363 1233
rect 439 1229 443 1233
rect 487 1231 491 1235
rect 495 1235 499 1239
rect 823 1239 827 1243
rect 1519 1243 1523 1247
rect 519 1229 523 1233
rect 599 1229 603 1233
rect 663 1231 667 1235
rect 671 1229 675 1233
rect 735 1231 739 1235
rect 743 1229 747 1233
rect 779 1231 780 1235
rect 780 1231 783 1235
rect 815 1229 819 1233
rect 847 1231 848 1235
rect 848 1231 851 1235
rect 895 1229 899 1233
rect 1327 1228 1331 1232
rect 1367 1232 1371 1236
rect 1495 1233 1499 1237
rect 1551 1235 1555 1239
rect 1559 1233 1563 1237
rect 1587 1235 1591 1239
rect 1695 1243 1699 1247
rect 1623 1233 1627 1237
rect 1687 1233 1691 1237
rect 1751 1235 1755 1239
rect 1759 1233 1763 1237
rect 1791 1235 1792 1239
rect 1792 1235 1795 1239
rect 1823 1233 1827 1237
rect 2087 1243 2091 1247
rect 1887 1233 1891 1237
rect 1951 1233 1955 1237
rect 2007 1235 2011 1239
rect 2015 1233 2019 1237
rect 2039 1235 2043 1239
rect 2079 1233 2083 1237
rect 2139 1235 2143 1239
rect 2151 1233 2155 1237
rect 2187 1235 2188 1239
rect 2188 1235 2191 1239
rect 2223 1233 2227 1237
rect 2287 1235 2291 1239
rect 2295 1233 2299 1237
rect 2583 1232 2587 1236
rect 111 1211 115 1215
rect 1327 1211 1331 1215
rect 1367 1215 1371 1219
rect 2583 1215 2587 1219
rect 159 1202 163 1206
rect 215 1202 219 1206
rect 295 1202 299 1206
rect 375 1202 379 1206
rect 455 1202 459 1206
rect 535 1202 539 1206
rect 615 1202 619 1206
rect 687 1202 691 1206
rect 759 1202 763 1206
rect 831 1202 835 1206
rect 911 1202 915 1206
rect 1511 1206 1515 1210
rect 1575 1206 1579 1210
rect 1639 1206 1643 1210
rect 1703 1206 1707 1210
rect 1775 1206 1779 1210
rect 1839 1206 1843 1210
rect 1903 1206 1907 1210
rect 1967 1206 1971 1210
rect 2031 1206 2035 1210
rect 2095 1206 2099 1210
rect 2167 1206 2171 1210
rect 2239 1206 2243 1210
rect 2311 1206 2315 1210
rect 151 1195 155 1199
rect 191 1195 192 1199
rect 192 1195 195 1199
rect 271 1195 272 1199
rect 272 1195 275 1199
rect 347 1195 351 1199
rect 495 1195 499 1199
rect 543 1195 547 1199
rect 663 1195 664 1199
rect 664 1195 667 1199
rect 735 1195 736 1199
rect 736 1195 739 1199
rect 823 1195 827 1199
rect 859 1195 863 1199
rect 1519 1199 1523 1203
rect 1551 1199 1552 1203
rect 1552 1199 1555 1203
rect 1663 1199 1667 1203
rect 1695 1199 1699 1203
rect 1751 1199 1752 1203
rect 1752 1199 1755 1203
rect 1927 1199 1931 1203
rect 1935 1199 1939 1203
rect 2007 1199 2008 1203
rect 2008 1199 2011 1203
rect 2087 1199 2091 1203
rect 2139 1199 2143 1203
rect 2219 1199 2220 1203
rect 2220 1199 2223 1203
rect 2287 1199 2288 1203
rect 2288 1199 2291 1203
rect 847 1187 851 1191
rect 135 1179 136 1183
rect 136 1179 139 1183
rect 259 1179 263 1183
rect 355 1179 359 1183
rect 487 1179 488 1183
rect 488 1179 491 1183
rect 679 1179 683 1183
rect 707 1179 711 1183
rect 787 1179 791 1183
rect 887 1179 888 1183
rect 888 1179 891 1183
rect 1003 1179 1007 1183
rect 1391 1179 1392 1183
rect 1392 1179 1395 1183
rect 1495 1179 1499 1183
rect 1587 1183 1591 1187
rect 1619 1179 1623 1183
rect 159 1174 163 1178
rect 239 1174 243 1178
rect 327 1174 331 1178
rect 423 1174 427 1178
rect 511 1174 515 1178
rect 599 1174 603 1178
rect 687 1174 691 1178
rect 767 1174 771 1178
rect 839 1174 843 1178
rect 911 1174 915 1178
rect 983 1174 987 1178
rect 1063 1174 1067 1178
rect 1415 1174 1419 1178
rect 1503 1174 1507 1178
rect 1723 1179 1727 1183
rect 1827 1179 1831 1183
rect 2039 1183 2043 1187
rect 2087 1179 2088 1183
rect 2088 1179 2091 1183
rect 2131 1179 2135 1183
rect 2295 1179 2299 1183
rect 2323 1179 2327 1183
rect 1599 1174 1603 1178
rect 1703 1174 1707 1178
rect 1807 1174 1811 1178
rect 1911 1174 1915 1178
rect 2015 1174 2019 1178
rect 2111 1174 2115 1178
rect 2207 1174 2211 1178
rect 2303 1174 2307 1178
rect 2399 1174 2403 1178
rect 111 1165 115 1169
rect 1327 1165 1331 1169
rect 1367 1165 1371 1169
rect 2583 1165 2587 1169
rect 135 1155 139 1159
rect 111 1148 115 1152
rect 143 1147 147 1151
rect 223 1147 227 1151
rect 259 1143 260 1147
rect 260 1143 263 1147
rect 311 1147 315 1151
rect 347 1143 348 1147
rect 348 1143 351 1147
rect 407 1147 411 1151
rect 887 1155 891 1159
rect 495 1147 499 1151
rect 583 1147 587 1151
rect 619 1143 620 1147
rect 620 1143 623 1147
rect 671 1147 675 1151
rect 707 1143 708 1147
rect 708 1143 711 1147
rect 751 1147 755 1151
rect 787 1143 788 1147
rect 788 1143 791 1147
rect 823 1147 827 1151
rect 859 1143 860 1147
rect 860 1143 863 1147
rect 895 1147 899 1151
rect 679 1135 683 1139
rect 967 1147 971 1151
rect 1003 1143 1004 1147
rect 1004 1143 1007 1147
rect 1047 1147 1051 1151
rect 1391 1155 1395 1159
rect 1327 1148 1331 1152
rect 1367 1148 1371 1152
rect 1399 1147 1403 1151
rect 1423 1143 1427 1147
rect 1487 1147 1491 1151
rect 2087 1155 2091 1159
rect 1583 1147 1587 1151
rect 1495 1135 1499 1139
rect 1687 1147 1691 1151
rect 1723 1143 1724 1147
rect 1724 1143 1727 1147
rect 1791 1147 1795 1151
rect 1827 1143 1828 1147
rect 1828 1143 1831 1147
rect 1895 1147 1899 1151
rect 1927 1143 1928 1147
rect 1928 1143 1931 1147
rect 1999 1147 2003 1151
rect 2095 1147 2099 1151
rect 2131 1143 2132 1147
rect 2132 1143 2135 1147
rect 2191 1147 2195 1151
rect 2219 1143 2223 1147
rect 2287 1147 2291 1151
rect 2323 1143 2324 1147
rect 2324 1143 2327 1147
rect 2383 1147 2387 1151
rect 2583 1148 2587 1152
rect 1015 1115 1019 1119
rect 111 1104 115 1108
rect 223 1105 227 1109
rect 311 1107 315 1111
rect 319 1105 323 1109
rect 355 1107 356 1111
rect 356 1107 359 1111
rect 423 1105 427 1109
rect 519 1107 523 1111
rect 527 1105 531 1109
rect 551 1107 555 1111
rect 631 1105 635 1109
rect 679 1107 683 1111
rect 727 1105 731 1109
rect 815 1107 819 1111
rect 823 1105 827 1109
rect 903 1107 907 1111
rect 911 1105 915 1109
rect 991 1105 995 1109
rect 1023 1107 1024 1111
rect 1024 1107 1027 1111
rect 1079 1105 1083 1109
rect 1159 1107 1163 1111
rect 1167 1105 1171 1109
rect 1327 1104 1331 1108
rect 1367 1108 1371 1112
rect 1399 1109 1403 1113
rect 1471 1111 1475 1115
rect 1479 1109 1483 1113
rect 1503 1111 1507 1115
rect 1583 1109 1587 1113
rect 1619 1111 1620 1115
rect 1620 1111 1623 1115
rect 1627 1115 1631 1119
rect 1687 1109 1691 1113
rect 1791 1109 1795 1113
rect 1887 1109 1891 1113
rect 1967 1111 1971 1115
rect 1975 1109 1979 1113
rect 2039 1111 2043 1115
rect 2063 1109 2067 1113
rect 2135 1111 2139 1115
rect 2143 1109 2147 1113
rect 2207 1111 2211 1115
rect 2215 1109 2219 1113
rect 2271 1111 2275 1115
rect 2295 1115 2299 1119
rect 2279 1109 2283 1113
rect 2343 1109 2347 1113
rect 2375 1111 2376 1115
rect 2376 1111 2379 1115
rect 2439 1119 2443 1123
rect 2407 1109 2411 1113
rect 2471 1109 2475 1113
rect 2519 1111 2523 1115
rect 2527 1109 2531 1113
rect 2583 1108 2587 1112
rect 111 1087 115 1091
rect 1327 1087 1331 1091
rect 1367 1091 1371 1095
rect 2583 1091 2587 1095
rect 239 1078 243 1082
rect 335 1078 339 1082
rect 439 1078 443 1082
rect 543 1078 547 1082
rect 647 1078 651 1082
rect 743 1078 747 1082
rect 839 1078 843 1082
rect 927 1078 931 1082
rect 1007 1078 1011 1082
rect 1095 1078 1099 1082
rect 1183 1078 1187 1082
rect 1415 1082 1419 1086
rect 1495 1082 1499 1086
rect 1599 1082 1603 1086
rect 1703 1082 1707 1086
rect 1807 1082 1811 1086
rect 1903 1082 1907 1086
rect 1991 1082 1995 1086
rect 2079 1082 2083 1086
rect 2159 1082 2163 1086
rect 2231 1082 2235 1086
rect 2295 1082 2299 1086
rect 2359 1082 2363 1086
rect 2423 1082 2427 1086
rect 2487 1082 2491 1086
rect 2543 1082 2547 1086
rect 219 1071 220 1075
rect 220 1071 223 1075
rect 311 1071 312 1075
rect 312 1071 315 1075
rect 455 1071 459 1075
rect 519 1071 520 1075
rect 520 1071 523 1075
rect 619 1071 623 1075
rect 535 1063 539 1067
rect 815 1071 816 1075
rect 816 1071 819 1075
rect 903 1071 904 1075
rect 904 1071 907 1075
rect 1015 1071 1019 1075
rect 1071 1071 1072 1075
rect 1072 1071 1075 1075
rect 1159 1071 1160 1075
rect 1160 1071 1163 1075
rect 1423 1075 1427 1079
rect 1471 1075 1472 1079
rect 1472 1075 1475 1079
rect 1627 1075 1631 1079
rect 1855 1075 1859 1079
rect 1967 1075 1968 1079
rect 1968 1075 1971 1079
rect 2127 1075 2131 1079
rect 2135 1075 2136 1079
rect 2136 1075 2139 1079
rect 2207 1075 2208 1079
rect 2208 1075 2211 1079
rect 2271 1075 2272 1079
rect 2272 1075 2275 1079
rect 2439 1075 2443 1079
rect 2479 1075 2483 1079
rect 2519 1075 2520 1079
rect 2520 1075 2523 1079
rect 1023 1063 1027 1067
rect 387 1055 391 1059
rect 495 1055 496 1059
rect 496 1055 499 1059
rect 563 1055 567 1059
rect 679 1055 680 1059
rect 680 1055 683 1059
rect 723 1055 727 1059
rect 879 1055 883 1059
rect 907 1055 911 1059
rect 995 1055 999 1059
rect 1063 1055 1067 1059
rect 1155 1055 1159 1059
rect 1503 1063 1507 1067
rect 1527 1059 1531 1063
rect 1555 1059 1559 1063
rect 1643 1059 1647 1063
rect 1747 1059 1751 1063
rect 1927 1059 1928 1063
rect 1928 1059 1931 1063
rect 2039 1059 2040 1063
rect 2040 1059 2043 1063
rect 2287 1067 2291 1071
rect 2247 1059 2248 1063
rect 2248 1059 2251 1063
rect 2375 1063 2379 1067
rect 2439 1059 2440 1063
rect 2440 1059 2443 1063
rect 2535 1059 2539 1063
rect 311 1050 315 1054
rect 367 1050 371 1054
rect 439 1050 443 1054
rect 519 1050 523 1054
rect 607 1050 611 1054
rect 703 1050 707 1054
rect 799 1050 803 1054
rect 887 1050 891 1054
rect 975 1050 979 1054
rect 1055 1050 1059 1054
rect 1135 1050 1139 1054
rect 1223 1050 1227 1054
rect 1287 1050 1291 1054
rect 1415 1054 1419 1058
rect 1471 1054 1475 1058
rect 1535 1054 1539 1058
rect 1623 1054 1627 1058
rect 1727 1054 1731 1058
rect 1839 1054 1843 1058
rect 1951 1054 1955 1058
rect 2063 1054 2067 1058
rect 2167 1054 2171 1058
rect 2271 1054 2275 1058
rect 2367 1054 2371 1058
rect 2463 1054 2467 1058
rect 2543 1054 2547 1058
rect 111 1041 115 1045
rect 1327 1041 1331 1045
rect 1367 1045 1371 1049
rect 2583 1045 2587 1049
rect 495 1031 499 1035
rect 1927 1035 1931 1039
rect 111 1024 115 1028
rect 295 1023 299 1027
rect 351 1023 355 1027
rect 387 1019 388 1023
rect 388 1019 391 1023
rect 423 1023 427 1027
rect 455 1019 456 1023
rect 456 1019 459 1023
rect 503 1023 507 1027
rect 535 1019 536 1023
rect 536 1019 539 1023
rect 591 1023 595 1027
rect 687 1023 691 1027
rect 723 1019 724 1023
rect 724 1019 727 1023
rect 783 1023 787 1027
rect 755 1015 759 1019
rect 871 1023 875 1027
rect 907 1019 908 1023
rect 908 1019 911 1023
rect 959 1023 963 1027
rect 995 1019 996 1023
rect 996 1019 999 1023
rect 1039 1023 1043 1027
rect 1071 1019 1072 1023
rect 1072 1019 1075 1023
rect 1119 1023 1123 1027
rect 1155 1019 1156 1023
rect 1156 1019 1159 1023
rect 1207 1023 1211 1027
rect 1235 1019 1239 1023
rect 1271 1023 1275 1027
rect 1327 1024 1331 1028
rect 1367 1028 1371 1032
rect 1399 1027 1403 1031
rect 1295 1019 1299 1023
rect 1455 1027 1459 1031
rect 1519 1027 1523 1031
rect 1555 1023 1556 1027
rect 1556 1023 1559 1027
rect 1607 1027 1611 1031
rect 1643 1023 1644 1027
rect 1644 1023 1647 1027
rect 1711 1027 1715 1031
rect 1747 1023 1748 1027
rect 1748 1023 1751 1027
rect 1823 1027 1827 1031
rect 1855 1023 1856 1027
rect 1856 1023 1859 1027
rect 1935 1027 1939 1031
rect 2047 1027 2051 1031
rect 2247 1035 2251 1039
rect 2151 1027 2155 1031
rect 2127 1019 2131 1023
rect 2255 1027 2259 1031
rect 2287 1023 2288 1027
rect 2288 1023 2291 1027
rect 2351 1027 2355 1031
rect 2439 1035 2443 1039
rect 2447 1027 2451 1031
rect 2479 1023 2480 1027
rect 2480 1023 2483 1027
rect 2527 1027 2531 1031
rect 2583 1028 2587 1032
rect 947 1007 951 1011
rect 1063 1007 1067 1011
rect 439 995 443 999
rect 111 984 115 988
rect 415 985 419 989
rect 463 987 467 991
rect 471 985 475 989
rect 519 987 523 991
rect 527 985 531 989
rect 563 987 564 991
rect 564 987 567 991
rect 591 985 595 989
rect 639 991 643 995
rect 807 995 811 999
rect 655 985 659 989
rect 719 985 723 989
rect 747 987 751 991
rect 783 985 787 989
rect 839 987 843 991
rect 847 985 851 989
rect 903 987 907 991
rect 911 985 915 989
rect 947 987 948 991
rect 948 987 951 991
rect 975 985 979 989
rect 1039 985 1043 989
rect 1103 985 1107 989
rect 1159 985 1163 989
rect 1215 985 1219 989
rect 1271 985 1275 989
rect 1327 984 1331 988
rect 1527 987 1531 991
rect 1367 976 1371 980
rect 1399 977 1403 981
rect 1447 979 1451 983
rect 1455 977 1459 981
rect 1503 979 1507 983
rect 1511 977 1515 981
rect 1559 979 1563 983
rect 1567 977 1571 981
rect 1631 979 1635 983
rect 1639 977 1643 981
rect 1711 979 1715 983
rect 1719 977 1723 981
rect 1807 977 1811 981
rect 1895 979 1899 983
rect 1903 977 1907 981
rect 2007 979 2011 983
rect 2015 977 2019 981
rect 2135 979 2139 983
rect 2143 977 2147 981
rect 2263 979 2267 983
rect 2271 977 2275 981
rect 2295 979 2299 983
rect 2407 977 2411 981
rect 2519 979 2523 983
rect 2535 983 2539 987
rect 2527 977 2531 981
rect 2583 976 2587 980
rect 111 967 115 971
rect 1327 967 1331 971
rect 431 958 435 962
rect 487 958 491 962
rect 543 958 547 962
rect 607 958 611 962
rect 671 958 675 962
rect 735 958 739 962
rect 799 958 803 962
rect 863 958 867 962
rect 927 958 931 962
rect 991 958 995 962
rect 1055 958 1059 962
rect 1119 958 1123 962
rect 1175 958 1179 962
rect 1231 958 1235 962
rect 1287 958 1291 962
rect 1367 959 1371 963
rect 2583 959 2587 963
rect 439 951 443 955
rect 463 951 464 955
rect 464 951 467 955
rect 519 951 520 955
rect 520 951 523 955
rect 639 951 643 955
rect 663 951 667 955
rect 755 951 759 955
rect 807 951 811 955
rect 839 951 840 955
rect 840 951 843 955
rect 903 951 904 955
rect 904 951 907 955
rect 1295 951 1299 955
rect 1415 950 1419 954
rect 1471 950 1475 954
rect 1527 950 1531 954
rect 1583 950 1587 954
rect 1655 950 1659 954
rect 1735 950 1739 954
rect 1823 950 1827 954
rect 1919 950 1923 954
rect 2031 950 2035 954
rect 2159 950 2163 954
rect 2287 950 2291 954
rect 2423 950 2427 954
rect 2543 950 2547 954
rect 415 935 419 939
rect 443 935 447 939
rect 499 935 503 939
rect 555 935 559 939
rect 679 935 680 939
rect 680 935 683 939
rect 747 939 751 943
rect 1431 943 1435 947
rect 1447 943 1448 947
rect 1448 943 1451 947
rect 1503 943 1504 947
rect 1504 943 1507 947
rect 1559 943 1560 947
rect 1560 943 1563 947
rect 1631 943 1632 947
rect 1632 943 1635 947
rect 1711 943 1712 947
rect 1712 943 1715 947
rect 1895 943 1896 947
rect 1896 943 1899 947
rect 2007 943 2008 947
rect 2008 943 2011 947
rect 2135 943 2136 947
rect 2136 943 2139 947
rect 2263 943 2264 947
rect 2264 943 2267 947
rect 2331 943 2335 947
rect 2519 943 2520 947
rect 2520 943 2523 947
rect 779 935 783 939
rect 423 930 427 934
rect 479 930 483 934
rect 535 930 539 934
rect 591 930 595 934
rect 647 930 651 934
rect 703 930 707 934
rect 759 930 763 934
rect 815 930 819 934
rect 111 921 115 925
rect 1327 921 1331 925
rect 1487 931 1491 935
rect 1447 923 1448 927
rect 1448 923 1451 927
rect 1631 931 1635 935
rect 2079 931 2083 935
rect 2295 931 2299 935
rect 1591 923 1592 927
rect 1592 923 1595 927
rect 2039 923 2040 927
rect 2040 923 2043 927
rect 2455 931 2459 935
rect 2415 923 2416 927
rect 2416 923 2419 927
rect 2535 923 2539 927
rect 1415 918 1419 922
rect 1471 918 1475 922
rect 1527 918 1531 922
rect 1615 918 1619 922
rect 1711 918 1715 922
rect 1823 918 1827 922
rect 1943 918 1947 922
rect 2063 918 2067 922
rect 2183 918 2187 922
rect 2311 918 2315 922
rect 2439 918 2443 922
rect 2543 918 2547 922
rect 679 911 683 915
rect 111 904 115 908
rect 407 903 411 907
rect 443 899 444 903
rect 444 899 447 903
rect 463 903 467 907
rect 499 899 500 903
rect 500 899 503 903
rect 519 903 523 907
rect 555 899 556 903
rect 556 899 559 903
rect 575 903 579 907
rect 631 903 635 907
rect 663 899 664 903
rect 664 899 667 903
rect 687 903 691 907
rect 695 895 699 899
rect 743 903 747 907
rect 779 899 780 903
rect 780 899 783 903
rect 799 903 803 907
rect 1367 909 1371 913
rect 2583 909 2587 913
rect 1327 904 1331 908
rect 1447 899 1451 903
rect 1367 892 1371 896
rect 1399 891 1403 895
rect 1431 887 1432 891
rect 1432 887 1435 891
rect 1455 891 1459 895
rect 1487 887 1488 891
rect 1488 887 1491 891
rect 1511 891 1515 895
rect 1591 899 1595 903
rect 1599 891 1603 895
rect 1631 887 1632 891
rect 1632 887 1635 891
rect 1695 891 1699 895
rect 1807 891 1811 895
rect 2039 899 2043 903
rect 1927 891 1931 895
rect 1951 887 1955 891
rect 2047 891 2051 895
rect 2079 887 2080 891
rect 2080 887 2083 891
rect 2167 891 2171 895
rect 2415 899 2419 903
rect 2295 891 2299 895
rect 2331 887 2332 891
rect 2332 887 2335 891
rect 2423 891 2427 895
rect 2455 887 2456 891
rect 2456 887 2459 891
rect 2527 891 2531 895
rect 2583 892 2587 896
rect 415 879 419 883
rect 111 868 115 872
rect 279 869 283 873
rect 327 871 331 875
rect 335 869 339 873
rect 383 871 387 875
rect 391 869 395 873
rect 447 871 451 875
rect 455 869 459 873
rect 511 871 515 875
rect 519 869 523 873
rect 575 871 579 875
rect 583 869 587 873
rect 647 869 651 873
rect 703 871 707 875
rect 711 869 715 873
rect 767 871 771 875
rect 775 869 779 873
rect 839 871 843 875
rect 847 869 851 873
rect 911 871 915 875
rect 919 869 923 873
rect 943 871 947 875
rect 1327 868 1331 872
rect 1751 867 1755 871
rect 1367 856 1371 860
rect 1471 857 1475 861
rect 1543 859 1547 863
rect 1551 857 1555 861
rect 1631 859 1635 863
rect 1639 857 1643 861
rect 1727 857 1731 861
rect 1759 859 1760 863
rect 1760 859 1763 863
rect 1815 857 1819 861
rect 1903 857 1907 861
rect 1983 859 1987 863
rect 1991 857 1995 861
rect 2047 859 2051 863
rect 2071 857 2075 861
rect 2135 859 2139 863
rect 2143 857 2147 861
rect 2207 859 2211 863
rect 2215 857 2219 861
rect 2271 859 2275 863
rect 2279 857 2283 861
rect 2335 859 2339 863
rect 2343 857 2347 861
rect 2399 859 2403 863
rect 2407 857 2411 861
rect 2463 859 2467 863
rect 2471 857 2475 861
rect 2519 859 2523 863
rect 2535 863 2539 867
rect 2527 857 2531 861
rect 2583 856 2587 860
rect 111 851 115 855
rect 1327 851 1331 855
rect 295 842 299 846
rect 351 842 355 846
rect 407 842 411 846
rect 471 842 475 846
rect 535 842 539 846
rect 599 842 603 846
rect 663 842 667 846
rect 727 842 731 846
rect 791 842 795 846
rect 863 842 867 846
rect 935 842 939 846
rect 327 835 328 839
rect 328 835 331 839
rect 383 835 384 839
rect 384 835 387 839
rect 447 835 448 839
rect 448 835 451 839
rect 511 835 512 839
rect 512 835 515 839
rect 575 835 576 839
rect 576 835 579 839
rect 695 835 699 839
rect 703 835 704 839
rect 704 835 707 839
rect 767 835 768 839
rect 768 835 771 839
rect 839 835 840 839
rect 840 835 843 839
rect 911 835 912 839
rect 912 835 915 839
rect 1367 839 1371 843
rect 2583 839 2587 843
rect 591 827 595 831
rect 1487 830 1491 834
rect 1567 830 1571 834
rect 1655 830 1659 834
rect 1743 830 1747 834
rect 1831 830 1835 834
rect 1919 830 1923 834
rect 2007 830 2011 834
rect 2087 830 2091 834
rect 2159 830 2163 834
rect 2231 830 2235 834
rect 2295 830 2299 834
rect 2359 830 2363 834
rect 2423 830 2427 834
rect 2487 830 2491 834
rect 2543 830 2547 834
rect 943 823 947 827
rect 159 815 163 819
rect 187 815 191 819
rect 251 815 255 819
rect 331 815 335 819
rect 419 815 423 819
rect 507 815 511 819
rect 691 815 695 819
rect 779 815 783 819
rect 1027 815 1031 819
rect 1543 823 1544 827
rect 1544 823 1547 827
rect 1631 823 1632 827
rect 1632 823 1635 827
rect 1751 823 1755 827
rect 1759 819 1763 823
rect 1771 823 1775 827
rect 1951 823 1955 827
rect 1983 823 1984 827
rect 1984 823 1987 827
rect 2127 823 2131 827
rect 2135 823 2136 827
rect 2136 823 2139 827
rect 2207 823 2208 827
rect 2208 823 2211 827
rect 2271 823 2272 827
rect 2272 823 2275 827
rect 2335 823 2336 827
rect 2336 823 2339 827
rect 2399 823 2400 827
rect 2400 823 2403 827
rect 2463 823 2464 827
rect 2464 823 2467 827
rect 2519 823 2520 827
rect 2520 823 2523 827
rect 167 810 171 814
rect 231 810 235 814
rect 311 810 315 814
rect 399 810 403 814
rect 487 810 491 814
rect 583 810 587 814
rect 671 810 675 814
rect 759 810 763 814
rect 839 810 843 814
rect 919 810 923 814
rect 1007 810 1011 814
rect 1095 810 1099 814
rect 111 801 115 805
rect 1327 801 1331 805
rect 1839 811 1843 815
rect 1707 803 1711 807
rect 1799 803 1800 807
rect 1800 803 1803 807
rect 1999 811 2003 815
rect 2047 803 2048 807
rect 2048 803 2051 807
rect 2151 803 2155 807
rect 2179 803 2183 807
rect 2267 803 2271 807
rect 1631 798 1635 802
rect 1687 798 1691 802
rect 1751 798 1755 802
rect 1823 798 1827 802
rect 1903 798 1907 802
rect 1991 798 1995 802
rect 2071 798 2075 802
rect 2159 798 2163 802
rect 2247 798 2251 802
rect 2335 798 2339 802
rect 2423 798 2427 802
rect 1367 789 1371 793
rect 2583 789 2587 793
rect 111 784 115 788
rect 151 783 155 787
rect 187 779 188 783
rect 188 779 191 783
rect 215 783 219 787
rect 251 779 252 783
rect 252 779 255 783
rect 295 783 299 787
rect 331 779 332 783
rect 332 779 335 783
rect 383 783 387 787
rect 419 779 420 783
rect 420 779 423 783
rect 471 783 475 787
rect 507 779 508 783
rect 508 779 511 783
rect 567 783 571 787
rect 591 779 595 783
rect 655 783 659 787
rect 691 779 692 783
rect 692 779 695 783
rect 743 783 747 787
rect 779 779 780 783
rect 780 779 783 783
rect 823 783 827 787
rect 903 783 907 787
rect 991 783 995 787
rect 1027 779 1028 783
rect 1028 779 1031 783
rect 1079 783 1083 787
rect 1327 784 1331 788
rect 1103 779 1107 783
rect 1799 779 1803 783
rect 1367 772 1371 776
rect 1615 771 1619 775
rect 1671 771 1675 775
rect 1707 767 1708 771
rect 1708 767 1711 771
rect 1735 771 1739 775
rect 1771 767 1772 771
rect 1772 767 1775 771
rect 1807 771 1811 775
rect 1839 767 1840 771
rect 1840 767 1843 771
rect 1887 771 1891 775
rect 1975 771 1979 775
rect 1999 767 2003 771
rect 2055 771 2059 775
rect 2087 767 2088 771
rect 2088 767 2091 771
rect 2143 771 2147 775
rect 2179 767 2180 771
rect 2180 767 2183 771
rect 2231 771 2235 775
rect 2267 767 2268 771
rect 2268 767 2271 771
rect 2319 771 2323 775
rect 2407 771 2411 775
rect 2583 772 2587 776
rect 2439 767 2440 771
rect 2440 767 2443 771
rect 159 751 163 755
rect 111 740 115 744
rect 143 741 147 745
rect 191 743 195 747
rect 199 741 203 745
rect 271 743 275 747
rect 279 741 283 745
rect 375 743 379 747
rect 383 741 387 745
rect 479 743 483 747
rect 487 741 491 745
rect 591 743 595 747
rect 599 741 603 745
rect 703 741 707 745
rect 799 743 803 747
rect 807 741 811 745
rect 895 743 899 747
rect 903 741 907 745
rect 983 743 987 747
rect 991 741 995 745
rect 1071 743 1075 747
rect 1079 741 1083 745
rect 1167 743 1171 747
rect 1175 741 1179 745
rect 1199 743 1203 747
rect 1327 740 1331 744
rect 1367 732 1371 736
rect 1567 733 1571 737
rect 1615 735 1619 739
rect 1623 733 1627 737
rect 1679 735 1683 739
rect 1687 733 1691 737
rect 1751 735 1755 739
rect 1759 733 1763 737
rect 1831 735 1835 739
rect 1839 733 1843 737
rect 1911 735 1915 739
rect 1919 733 1923 737
rect 1999 733 2003 737
rect 2031 735 2032 739
rect 2032 735 2035 739
rect 2055 739 2059 743
rect 2151 743 2155 747
rect 2079 733 2083 737
rect 2159 733 2163 737
rect 2239 735 2243 739
rect 2247 733 2251 737
rect 2327 735 2331 739
rect 2335 733 2339 737
rect 2583 732 2587 736
rect 111 723 115 727
rect 1327 723 1331 727
rect 159 714 163 718
rect 215 714 219 718
rect 295 714 299 718
rect 399 714 403 718
rect 503 714 507 718
rect 615 714 619 718
rect 719 714 723 718
rect 823 714 827 718
rect 919 714 923 718
rect 1007 714 1011 718
rect 1095 714 1099 718
rect 1191 714 1195 718
rect 1367 715 1371 719
rect 2583 715 2587 719
rect 191 707 192 711
rect 192 707 195 711
rect 271 707 272 711
rect 272 707 275 711
rect 375 707 376 711
rect 376 707 379 711
rect 479 707 480 711
rect 480 707 483 711
rect 591 707 592 711
rect 592 707 595 711
rect 699 707 700 711
rect 700 707 703 711
rect 799 707 800 711
rect 800 707 803 711
rect 895 707 896 711
rect 896 707 899 711
rect 983 707 984 711
rect 984 707 987 711
rect 1071 707 1072 711
rect 1072 707 1075 711
rect 1167 707 1168 711
rect 1168 707 1171 711
rect 1583 706 1587 710
rect 1639 706 1643 710
rect 1703 706 1707 710
rect 1775 706 1779 710
rect 1855 706 1859 710
rect 1935 706 1939 710
rect 2015 706 2019 710
rect 2095 706 2099 710
rect 2175 706 2179 710
rect 2263 706 2267 710
rect 2351 706 2355 710
rect 367 699 371 703
rect 135 691 136 695
rect 136 691 139 695
rect 179 691 183 695
rect 243 691 247 695
rect 375 691 379 695
rect 467 691 471 695
rect 727 699 731 703
rect 687 691 688 695
rect 688 691 691 695
rect 887 699 891 703
rect 847 691 848 695
rect 848 691 851 695
rect 943 691 947 695
rect 1199 695 1203 699
rect 1615 699 1616 703
rect 1616 699 1619 703
rect 1679 699 1680 703
rect 1680 699 1683 703
rect 1751 699 1752 703
rect 1752 699 1755 703
rect 1831 699 1832 703
rect 1832 699 1835 703
rect 1911 699 1912 703
rect 1912 699 1915 703
rect 2055 699 2059 703
rect 2087 699 2091 703
rect 2139 699 2143 703
rect 2239 699 2240 703
rect 2240 699 2243 703
rect 2327 699 2328 703
rect 2328 699 2331 703
rect 1839 691 1843 695
rect 159 686 163 690
rect 215 686 219 690
rect 279 686 283 690
rect 359 686 363 690
rect 447 686 451 690
rect 535 686 539 690
rect 623 686 627 690
rect 711 686 715 690
rect 791 686 795 690
rect 871 686 875 690
rect 951 686 955 690
rect 1039 686 1043 690
rect 2031 691 2035 695
rect 1407 683 1411 687
rect 1435 683 1439 687
rect 1739 683 1743 687
rect 1947 683 1951 687
rect 2223 691 2227 695
rect 2183 683 2184 687
rect 2184 683 2187 687
rect 2287 683 2291 687
rect 2439 687 2443 691
rect 111 677 115 681
rect 1327 677 1331 681
rect 1415 678 1419 682
rect 1511 678 1515 682
rect 1615 678 1619 682
rect 1719 678 1723 682
rect 1823 678 1827 682
rect 1927 678 1931 682
rect 2023 678 2027 682
rect 2119 678 2123 682
rect 2207 678 2211 682
rect 2295 678 2299 682
rect 2391 678 2395 682
rect 135 667 139 671
rect 111 660 115 664
rect 143 659 147 663
rect 179 655 180 659
rect 180 655 183 659
rect 199 659 203 663
rect 243 655 247 659
rect 263 659 267 663
rect 343 659 347 663
rect 367 655 371 659
rect 431 659 435 663
rect 467 655 468 659
rect 468 655 471 659
rect 519 659 523 663
rect 687 667 691 671
rect 607 659 611 663
rect 631 655 635 659
rect 695 659 699 663
rect 727 655 728 659
rect 728 655 731 659
rect 775 659 779 663
rect 847 667 851 671
rect 1367 669 1371 673
rect 2583 669 2587 673
rect 855 659 859 663
rect 887 655 888 659
rect 888 655 891 659
rect 935 659 939 663
rect 1023 659 1027 663
rect 1327 660 1331 664
rect 2183 659 2187 663
rect 943 647 947 651
rect 1367 652 1371 656
rect 1399 651 1403 655
rect 1435 647 1436 651
rect 1436 647 1439 651
rect 1495 651 1499 655
rect 1599 651 1603 655
rect 1703 651 1707 655
rect 1739 647 1740 651
rect 1740 647 1743 651
rect 1807 651 1811 655
rect 1839 647 1840 651
rect 1840 647 1843 651
rect 1911 651 1915 655
rect 1947 647 1948 651
rect 1948 647 1951 651
rect 2007 651 2011 655
rect 2031 647 2035 651
rect 2103 651 2107 655
rect 2139 647 2140 651
rect 2140 647 2143 651
rect 2191 651 2195 655
rect 2223 647 2224 651
rect 2224 647 2227 651
rect 2279 651 2283 655
rect 2375 651 2379 655
rect 2583 652 2587 656
rect 375 635 379 639
rect 2287 639 2291 643
rect 335 627 339 631
rect 111 616 115 620
rect 143 617 147 621
rect 191 619 195 623
rect 199 617 203 621
rect 247 619 251 623
rect 255 617 259 621
rect 311 617 315 621
rect 343 619 344 623
rect 344 619 347 623
rect 391 617 395 621
rect 471 619 475 623
rect 479 617 483 621
rect 575 617 579 621
rect 671 619 675 623
rect 679 617 683 621
rect 775 619 779 623
rect 783 617 787 621
rect 879 619 883 623
rect 887 617 891 621
rect 919 619 920 623
rect 920 619 923 623
rect 991 617 995 621
rect 1079 619 1083 623
rect 1087 617 1091 621
rect 1183 619 1187 623
rect 1191 617 1195 621
rect 1263 619 1267 623
rect 1271 617 1275 621
rect 1639 631 1643 635
rect 1327 616 1331 620
rect 1367 616 1371 620
rect 1399 617 1403 621
rect 1423 619 1427 623
rect 1511 617 1515 621
rect 1647 617 1651 621
rect 1775 619 1779 623
rect 1783 617 1787 621
rect 1815 619 1816 623
rect 1816 619 1819 623
rect 1911 617 1915 621
rect 1939 619 1943 623
rect 2039 617 2043 621
rect 2159 617 2163 621
rect 2271 619 2275 623
rect 2279 617 2283 621
rect 2399 619 2403 623
rect 2407 617 2411 621
rect 2439 619 2440 623
rect 2440 619 2443 623
rect 2583 616 2587 620
rect 111 599 115 603
rect 1327 599 1331 603
rect 1367 599 1371 603
rect 2583 599 2587 603
rect 159 590 163 594
rect 215 590 219 594
rect 271 590 275 594
rect 327 590 331 594
rect 407 590 411 594
rect 495 590 499 594
rect 591 590 595 594
rect 695 590 699 594
rect 799 590 803 594
rect 903 590 907 594
rect 1007 590 1011 594
rect 1103 590 1107 594
rect 1207 590 1211 594
rect 1287 590 1291 594
rect 1415 590 1419 594
rect 1527 590 1531 594
rect 1663 590 1667 594
rect 1799 590 1803 594
rect 1927 590 1931 594
rect 2055 590 2059 594
rect 2175 590 2179 594
rect 2295 590 2299 594
rect 2423 590 2427 594
rect 191 583 192 587
rect 192 583 195 587
rect 247 583 248 587
rect 248 583 251 587
rect 335 583 339 587
rect 355 583 359 587
rect 471 583 472 587
rect 472 583 475 587
rect 631 583 635 587
rect 671 583 672 587
rect 672 583 675 587
rect 775 583 776 587
rect 776 583 779 587
rect 879 583 880 587
rect 880 583 883 587
rect 1071 583 1075 587
rect 1079 583 1080 587
rect 1080 583 1083 587
rect 1183 583 1184 587
rect 1184 583 1187 587
rect 1263 583 1264 587
rect 1264 583 1267 587
rect 1491 583 1495 587
rect 1639 583 1640 587
rect 1640 583 1643 587
rect 1775 583 1776 587
rect 1776 583 1779 587
rect 2031 583 2032 587
rect 2032 583 2035 587
rect 2255 583 2259 587
rect 2271 583 2272 587
rect 2272 583 2275 587
rect 2399 583 2400 587
rect 2400 583 2403 587
rect 343 575 347 579
rect 191 567 195 571
rect 391 567 392 571
rect 392 567 395 571
rect 531 567 535 571
rect 847 575 851 579
rect 807 567 808 571
rect 808 567 811 571
rect 919 567 920 571
rect 920 567 923 571
rect 1199 575 1203 579
rect 1159 567 1160 571
rect 1160 567 1163 571
rect 1423 571 1427 575
rect 199 562 203 566
rect 263 562 267 566
rect 335 562 339 566
rect 415 562 419 566
rect 511 562 515 566
rect 615 562 619 566
rect 719 562 723 566
rect 831 562 835 566
rect 943 562 947 566
rect 1063 562 1067 566
rect 1183 562 1187 566
rect 1287 562 1291 566
rect 1391 563 1392 567
rect 1392 563 1395 567
rect 1435 563 1439 567
rect 1655 571 1659 575
rect 1623 563 1624 567
rect 1624 563 1627 567
rect 1719 563 1723 567
rect 1771 563 1775 567
rect 1939 563 1940 567
rect 1940 563 1943 567
rect 2075 563 2079 567
rect 2215 563 2216 567
rect 2216 563 2219 567
rect 2415 571 2419 575
rect 2375 563 2376 567
rect 2376 563 2379 567
rect 2435 563 2439 567
rect 2499 563 2503 567
rect 1415 558 1419 562
rect 111 553 115 557
rect 1471 558 1475 562
rect 1551 558 1555 562
rect 1647 558 1651 562
rect 1751 558 1755 562
rect 1855 558 1859 562
rect 1959 558 1963 562
rect 2055 558 2059 562
rect 2151 558 2155 562
rect 2239 558 2243 562
rect 2319 558 2323 562
rect 2399 558 2403 562
rect 2479 558 2483 562
rect 2543 558 2547 562
rect 1327 553 1331 557
rect 1367 549 1371 553
rect 2583 549 2587 553
rect 391 543 395 547
rect 111 536 115 540
rect 183 535 187 539
rect 247 535 251 539
rect 319 535 323 539
rect 355 531 356 535
rect 356 531 359 535
rect 399 535 403 539
rect 191 523 195 527
rect 495 535 499 539
rect 531 531 532 535
rect 532 531 535 535
rect 599 535 603 539
rect 807 543 811 547
rect 703 535 707 539
rect 727 531 731 535
rect 815 535 819 539
rect 847 531 848 535
rect 848 531 851 535
rect 927 535 931 539
rect 1159 543 1163 547
rect 1047 535 1051 539
rect 1071 531 1075 535
rect 1167 535 1171 539
rect 1199 531 1200 535
rect 1200 531 1203 535
rect 1271 535 1275 539
rect 1327 536 1331 540
rect 1391 539 1395 543
rect 1367 532 1371 536
rect 1399 531 1403 535
rect 1435 527 1436 531
rect 1436 527 1439 531
rect 1455 531 1459 535
rect 1491 527 1492 531
rect 1492 527 1495 531
rect 1535 531 1539 535
rect 1623 539 1627 543
rect 1631 531 1635 535
rect 1655 527 1659 531
rect 1735 531 1739 535
rect 1771 527 1772 531
rect 1772 527 1775 531
rect 1839 531 1843 535
rect 2215 539 2219 543
rect 1943 531 1947 535
rect 2039 531 2043 535
rect 2075 527 2076 531
rect 2076 527 2079 531
rect 2135 531 2139 535
rect 2023 519 2027 523
rect 2223 531 2227 535
rect 2255 527 2256 531
rect 2256 527 2259 531
rect 2303 531 2307 535
rect 2375 539 2379 543
rect 2383 531 2387 535
rect 2415 527 2416 531
rect 2416 527 2419 531
rect 2463 531 2467 535
rect 2499 527 2500 531
rect 2500 527 2503 531
rect 2527 531 2531 535
rect 2583 532 2587 536
rect 519 503 523 507
rect 1543 507 1547 511
rect 111 492 115 496
rect 303 493 307 497
rect 351 495 355 499
rect 359 493 363 497
rect 415 495 419 499
rect 423 493 427 497
rect 495 493 499 497
rect 527 495 528 499
rect 528 495 531 499
rect 575 493 579 497
rect 639 495 643 499
rect 647 493 651 497
rect 719 493 723 497
rect 775 495 779 499
rect 791 493 795 497
rect 855 495 859 499
rect 863 493 867 497
rect 927 495 931 499
rect 935 493 939 497
rect 999 495 1003 499
rect 1007 493 1011 497
rect 1079 495 1083 499
rect 1087 493 1091 497
rect 1111 495 1115 499
rect 1327 492 1331 496
rect 1367 496 1371 500
rect 1535 497 1539 501
rect 1591 499 1595 503
rect 1599 497 1603 501
rect 1663 499 1667 503
rect 1671 497 1675 501
rect 1719 499 1723 503
rect 1751 497 1755 501
rect 1831 499 1835 503
rect 1839 497 1843 501
rect 1919 499 1923 503
rect 1927 497 1931 501
rect 2015 497 2019 501
rect 2087 499 2091 503
rect 2095 497 2099 501
rect 2167 499 2171 503
rect 2175 497 2179 501
rect 2199 499 2203 503
rect 2255 497 2259 501
rect 2319 499 2323 503
rect 2327 497 2331 501
rect 2391 499 2395 503
rect 2399 497 2403 501
rect 2435 499 2436 503
rect 2436 499 2439 503
rect 2471 497 2475 501
rect 2495 499 2499 503
rect 2527 497 2531 501
rect 2583 496 2587 500
rect 111 475 115 479
rect 1327 475 1331 479
rect 1367 479 1371 483
rect 2583 479 2587 483
rect 319 466 323 470
rect 375 466 379 470
rect 439 466 443 470
rect 511 466 515 470
rect 591 466 595 470
rect 663 466 667 470
rect 735 466 739 470
rect 807 466 811 470
rect 879 466 883 470
rect 951 466 955 470
rect 1023 466 1027 470
rect 1103 466 1107 470
rect 1551 470 1555 474
rect 1615 470 1619 474
rect 1687 470 1691 474
rect 1767 470 1771 474
rect 1855 470 1859 474
rect 1943 470 1947 474
rect 2031 470 2035 474
rect 2111 470 2115 474
rect 2191 470 2195 474
rect 2271 470 2275 474
rect 2343 470 2347 474
rect 2415 470 2419 474
rect 2487 470 2491 474
rect 2543 470 2547 474
rect 351 459 352 463
rect 352 459 355 463
rect 415 459 416 463
rect 416 459 419 463
rect 519 459 523 463
rect 583 459 587 463
rect 639 459 640 463
rect 640 459 643 463
rect 727 459 731 463
rect 775 459 779 463
rect 855 459 856 463
rect 856 459 859 463
rect 927 459 928 463
rect 928 459 931 463
rect 999 459 1000 463
rect 1000 459 1003 463
rect 1079 459 1080 463
rect 1080 459 1083 463
rect 1543 463 1547 467
rect 1591 463 1592 467
rect 1592 463 1595 467
rect 1663 463 1664 467
rect 1664 463 1667 467
rect 1775 463 1779 467
rect 1831 463 1832 467
rect 1832 463 1835 467
rect 1919 463 1920 467
rect 1920 463 1923 467
rect 2023 463 2027 467
rect 2087 463 2088 467
rect 2088 463 2091 467
rect 2167 463 2168 467
rect 2168 463 2171 467
rect 2319 463 2320 467
rect 2320 463 2323 467
rect 2391 463 2392 467
rect 2392 463 2395 467
rect 2559 463 2563 467
rect 527 451 531 455
rect 431 443 432 447
rect 432 443 435 447
rect 471 443 475 447
rect 531 443 535 447
rect 743 451 747 455
rect 703 443 704 447
rect 704 443 707 447
rect 791 443 795 447
rect 1111 451 1115 455
rect 891 443 895 447
rect 963 443 967 447
rect 1035 443 1039 447
rect 1123 443 1127 447
rect 1179 443 1183 447
rect 1623 443 1624 447
rect 1624 443 1627 447
rect 1667 443 1671 447
rect 1723 443 1727 447
rect 1887 451 1891 455
rect 2495 455 2499 459
rect 1847 443 1848 447
rect 1848 443 1851 447
rect 1919 443 1923 447
rect 1975 443 1976 447
rect 1976 443 1979 447
rect 2079 443 2083 447
rect 2199 447 2203 451
rect 2211 443 2215 447
rect 2331 443 2335 447
rect 2535 443 2539 447
rect 455 438 459 442
rect 511 438 515 442
rect 575 438 579 442
rect 647 438 651 442
rect 727 438 731 442
rect 799 438 803 442
rect 871 438 875 442
rect 943 438 947 442
rect 1015 438 1019 442
rect 1087 438 1091 442
rect 1159 438 1163 442
rect 1239 438 1243 442
rect 1647 438 1651 442
rect 1703 438 1707 442
rect 1759 438 1763 442
rect 1815 438 1819 442
rect 1871 438 1875 442
rect 1927 438 1931 442
rect 1999 438 2003 442
rect 2087 438 2091 442
rect 2191 438 2195 442
rect 2311 438 2315 442
rect 2439 438 2443 442
rect 2543 438 2547 442
rect 111 429 115 433
rect 1327 429 1331 433
rect 1367 429 1371 433
rect 2583 429 2587 433
rect 431 419 435 423
rect 111 412 115 416
rect 439 411 443 415
rect 471 407 472 411
rect 472 407 475 411
rect 495 411 499 415
rect 531 407 532 411
rect 532 407 535 411
rect 559 411 563 415
rect 583 407 587 411
rect 631 411 635 415
rect 703 419 707 423
rect 711 411 715 415
rect 743 407 744 411
rect 744 407 747 411
rect 783 411 787 415
rect 1623 419 1627 423
rect 855 411 859 415
rect 891 407 892 411
rect 892 407 895 411
rect 927 411 931 415
rect 963 407 964 411
rect 964 407 967 411
rect 999 411 1003 415
rect 1035 407 1036 411
rect 1036 407 1039 411
rect 1071 411 1075 415
rect 1123 411 1127 415
rect 1143 411 1147 415
rect 1179 407 1180 411
rect 1180 407 1183 411
rect 1223 411 1227 415
rect 1327 412 1331 416
rect 1367 412 1371 416
rect 1631 411 1635 415
rect 1255 407 1256 411
rect 1256 407 1259 411
rect 1667 407 1668 411
rect 1668 407 1671 411
rect 1687 411 1691 415
rect 1723 407 1724 411
rect 1724 407 1727 411
rect 1743 411 1747 415
rect 1775 407 1776 411
rect 1776 407 1779 411
rect 1799 411 1803 415
rect 1847 419 1851 423
rect 1855 411 1859 415
rect 1887 407 1888 411
rect 1888 407 1891 411
rect 1911 411 1915 415
rect 1975 419 1979 423
rect 1983 411 1987 415
rect 2019 407 2020 411
rect 2020 407 2023 411
rect 2071 411 2075 415
rect 2175 411 2179 415
rect 2211 407 2212 411
rect 2212 407 2215 411
rect 2295 411 2299 415
rect 2331 407 2332 411
rect 2332 407 2335 411
rect 2423 411 2427 415
rect 2455 407 2456 411
rect 2456 407 2459 411
rect 2527 411 2531 415
rect 2583 412 2587 416
rect 2559 407 2560 411
rect 2560 407 2563 411
rect 111 372 115 376
rect 415 373 419 377
rect 463 375 467 379
rect 471 373 475 377
rect 527 375 531 379
rect 535 373 539 377
rect 599 375 603 379
rect 607 373 611 377
rect 679 375 683 379
rect 687 373 691 377
rect 711 375 715 379
rect 767 373 771 377
rect 791 375 795 379
rect 935 383 939 387
rect 1919 387 1923 391
rect 847 373 851 377
rect 927 373 931 377
rect 999 375 1003 379
rect 1007 373 1011 377
rect 1079 375 1083 379
rect 1087 373 1091 377
rect 1175 373 1179 377
rect 1263 373 1267 377
rect 1327 372 1331 376
rect 1367 376 1371 380
rect 1655 377 1659 381
rect 1703 379 1707 383
rect 1711 377 1715 381
rect 1759 379 1763 383
rect 1767 377 1771 381
rect 1815 379 1819 383
rect 1823 377 1827 381
rect 1871 379 1875 383
rect 1879 377 1883 381
rect 1943 379 1947 383
rect 1951 377 1955 381
rect 2039 377 2043 381
rect 2143 379 2147 383
rect 2151 377 2155 381
rect 2271 379 2275 383
rect 2279 377 2283 381
rect 2407 379 2411 383
rect 2415 377 2419 381
rect 2439 379 2443 383
rect 2535 383 2539 387
rect 2527 377 2531 381
rect 2583 376 2587 380
rect 111 355 115 359
rect 1327 355 1331 359
rect 1367 359 1371 363
rect 2583 359 2587 363
rect 431 346 435 350
rect 487 346 491 350
rect 551 346 555 350
rect 623 346 627 350
rect 703 346 707 350
rect 783 346 787 350
rect 863 346 867 350
rect 943 346 947 350
rect 1023 346 1027 350
rect 1103 346 1107 350
rect 1191 346 1195 350
rect 1279 346 1283 350
rect 1671 350 1675 354
rect 1727 350 1731 354
rect 1783 350 1787 354
rect 1839 350 1843 354
rect 1895 350 1899 354
rect 1967 350 1971 354
rect 2055 350 2059 354
rect 2167 350 2171 354
rect 2295 350 2299 354
rect 2431 350 2435 354
rect 2543 350 2547 354
rect 455 339 459 343
rect 463 339 464 343
rect 464 339 467 343
rect 527 339 528 343
rect 528 339 531 343
rect 599 339 600 343
rect 600 339 603 343
rect 679 339 680 343
rect 680 339 683 343
rect 855 339 859 343
rect 935 339 939 343
rect 999 339 1000 343
rect 1000 339 1003 343
rect 1255 339 1256 343
rect 1256 339 1259 343
rect 1703 343 1704 347
rect 1704 343 1707 347
rect 1759 343 1760 347
rect 1760 343 1763 347
rect 1815 343 1816 347
rect 1816 343 1819 347
rect 1871 343 1872 347
rect 1872 343 1875 347
rect 1943 343 1944 347
rect 1944 343 1947 347
rect 2019 343 2023 347
rect 2143 343 2144 347
rect 2144 343 2147 347
rect 2271 343 2272 347
rect 2272 343 2275 347
rect 2407 343 2408 347
rect 2408 343 2411 347
rect 2559 343 2563 347
rect 439 323 440 327
rect 440 323 443 327
rect 511 323 515 327
rect 711 331 715 335
rect 595 323 599 327
rect 651 323 655 327
rect 935 331 939 335
rect 1983 335 1987 339
rect 903 323 904 327
rect 904 323 907 327
rect 963 323 967 327
rect 1079 323 1083 327
rect 1131 323 1135 327
rect 1623 323 1627 327
rect 1651 323 1655 327
rect 1707 323 1711 327
rect 1763 323 1767 327
rect 1827 323 1831 327
rect 1907 323 1911 327
rect 2031 323 2032 327
rect 2032 323 2035 327
rect 2123 323 2124 327
rect 2124 323 2127 327
rect 2223 323 2227 327
rect 2251 323 2255 327
rect 2331 323 2335 327
rect 2455 323 2456 327
rect 2456 323 2459 327
rect 2499 323 2503 327
rect 463 318 467 322
rect 519 318 523 322
rect 575 318 579 322
rect 631 318 635 322
rect 695 318 699 322
rect 767 318 771 322
rect 847 318 851 322
rect 927 318 931 322
rect 1015 318 1019 322
rect 1111 318 1115 322
rect 1215 318 1219 322
rect 1631 318 1635 322
rect 1687 318 1691 322
rect 1743 318 1747 322
rect 1807 318 1811 322
rect 1887 318 1891 322
rect 1967 318 1971 322
rect 2055 318 2059 322
rect 2143 318 2147 322
rect 2231 318 2235 322
rect 2311 318 2315 322
rect 2391 318 2395 322
rect 2479 318 2483 322
rect 2543 318 2547 322
rect 111 309 115 313
rect 1327 309 1331 313
rect 1367 309 1371 313
rect 2583 309 2587 313
rect 439 299 443 303
rect 111 292 115 296
rect 447 291 451 295
rect 455 283 459 287
rect 503 291 507 295
rect 903 299 907 303
rect 559 291 563 295
rect 595 287 596 291
rect 596 287 599 291
rect 615 291 619 295
rect 651 287 652 291
rect 652 287 655 291
rect 679 291 683 295
rect 711 287 712 291
rect 712 287 715 291
rect 751 291 755 295
rect 831 291 835 295
rect 855 287 859 291
rect 911 291 915 295
rect 935 287 939 291
rect 999 291 1003 295
rect 2031 299 2035 303
rect 1095 291 1099 295
rect 1131 287 1132 291
rect 1132 287 1135 291
rect 1199 291 1203 295
rect 1327 292 1331 296
rect 1223 287 1227 291
rect 1367 292 1371 296
rect 1615 291 1619 295
rect 1651 287 1652 291
rect 1652 287 1655 291
rect 1671 291 1675 295
rect 1707 287 1708 291
rect 1708 287 1711 291
rect 1727 291 1731 295
rect 1763 287 1764 291
rect 1764 287 1767 291
rect 1791 291 1795 295
rect 1827 287 1828 291
rect 1828 287 1831 291
rect 1871 291 1875 295
rect 1907 287 1908 291
rect 1908 287 1911 291
rect 1951 291 1955 295
rect 1983 287 1984 291
rect 1984 287 1987 291
rect 2039 291 2043 295
rect 2127 291 2131 295
rect 2215 291 2219 295
rect 2251 287 2252 291
rect 2252 287 2255 291
rect 2295 291 2299 295
rect 2331 287 2332 291
rect 2332 287 2335 291
rect 2375 291 2379 295
rect 2399 287 2403 291
rect 2463 291 2467 295
rect 2499 287 2500 291
rect 2500 287 2503 291
rect 2527 291 2531 295
rect 2583 292 2587 296
rect 2559 287 2560 291
rect 2560 287 2563 291
rect 511 263 515 267
rect 111 252 115 256
rect 287 253 291 257
rect 343 255 347 259
rect 359 253 363 257
rect 431 255 435 259
rect 439 253 443 257
rect 519 255 523 259
rect 527 253 531 257
rect 615 255 619 259
rect 847 263 851 267
rect 1623 267 1627 271
rect 623 253 627 257
rect 719 253 723 257
rect 767 255 771 259
rect 823 253 827 257
rect 919 255 923 259
rect 927 253 931 257
rect 963 255 964 259
rect 964 255 967 259
rect 1031 253 1035 257
rect 1143 253 1147 257
rect 1247 255 1251 259
rect 1255 253 1259 257
rect 1279 255 1283 259
rect 1327 252 1331 256
rect 1367 256 1371 260
rect 1535 257 1539 261
rect 1599 259 1603 263
rect 1607 257 1611 261
rect 1679 259 1683 263
rect 1687 257 1691 261
rect 1767 259 1771 263
rect 1775 257 1779 261
rect 1847 259 1851 263
rect 2223 267 2227 271
rect 2455 267 2459 271
rect 1863 257 1867 261
rect 1951 257 1955 261
rect 2031 259 2035 263
rect 2039 257 2043 261
rect 2071 259 2072 263
rect 2072 259 2075 263
rect 2119 257 2123 261
rect 2191 259 2195 263
rect 2199 257 2203 261
rect 2255 259 2259 263
rect 2271 257 2275 261
rect 2327 259 2331 263
rect 2335 257 2339 261
rect 2407 257 2411 261
rect 2471 257 2475 261
rect 2495 259 2499 263
rect 2527 257 2531 261
rect 2583 256 2587 260
rect 111 235 115 239
rect 1327 235 1331 239
rect 1367 239 1371 243
rect 2583 239 2587 243
rect 303 226 307 230
rect 375 226 379 230
rect 455 226 459 230
rect 543 226 547 230
rect 639 226 643 230
rect 735 226 739 230
rect 839 226 843 230
rect 943 226 947 230
rect 1047 226 1051 230
rect 1159 226 1163 230
rect 1271 226 1275 230
rect 1551 230 1555 234
rect 1623 230 1627 234
rect 1703 230 1707 234
rect 1791 230 1795 234
rect 1879 230 1883 234
rect 1967 230 1971 234
rect 2055 230 2059 234
rect 2135 230 2139 234
rect 2215 230 2219 234
rect 2287 230 2291 234
rect 2351 230 2355 234
rect 2423 230 2427 234
rect 2487 230 2491 234
rect 2543 230 2547 234
rect 335 219 339 223
rect 343 219 347 223
rect 431 219 432 223
rect 432 219 435 223
rect 519 219 520 223
rect 520 219 523 223
rect 615 219 616 223
rect 616 219 619 223
rect 711 219 712 223
rect 712 219 715 223
rect 847 219 851 223
rect 919 219 920 223
rect 920 219 923 223
rect 1039 219 1043 223
rect 1223 219 1227 223
rect 1247 219 1248 223
rect 1248 219 1251 223
rect 1591 223 1595 227
rect 1599 223 1600 227
rect 1600 223 1603 227
rect 1679 223 1680 227
rect 1680 223 1683 227
rect 1767 223 1768 227
rect 1768 223 1771 227
rect 1847 223 1851 227
rect 2031 223 2032 227
rect 2032 223 2035 227
rect 2183 223 2187 227
rect 2191 223 2192 227
rect 2192 223 2195 227
rect 2255 223 2259 227
rect 2327 223 2328 227
rect 2328 223 2331 227
rect 2399 223 2400 227
rect 2400 223 2403 227
rect 191 207 195 211
rect 219 207 223 211
rect 291 207 295 211
rect 483 207 487 211
rect 655 207 656 211
rect 656 207 659 211
rect 767 207 768 211
rect 768 207 771 211
rect 887 207 888 211
rect 888 207 891 211
rect 931 207 935 211
rect 1115 207 1119 211
rect 1279 211 1283 215
rect 1407 211 1411 215
rect 1435 211 1439 215
rect 1499 211 1503 215
rect 1579 211 1583 215
rect 1675 211 1679 215
rect 1771 211 1775 215
rect 1935 211 1936 215
rect 1936 211 1939 215
rect 2071 215 2075 219
rect 2495 219 2499 223
rect 2559 223 2563 227
rect 2159 211 2163 215
rect 2239 211 2240 215
rect 2240 211 2243 215
rect 2335 211 2336 215
rect 2336 211 2339 215
rect 199 202 203 206
rect 271 202 275 206
rect 359 202 363 206
rect 463 202 467 206
rect 567 202 571 206
rect 679 202 683 206
rect 791 202 795 206
rect 911 202 915 206
rect 1031 202 1035 206
rect 1151 202 1155 206
rect 1271 202 1275 206
rect 1415 206 1419 210
rect 1479 206 1483 210
rect 1559 206 1563 210
rect 1655 206 1659 210
rect 1751 206 1755 210
rect 1855 206 1859 210
rect 1959 206 1963 210
rect 2063 206 2067 210
rect 2167 206 2171 210
rect 2263 206 2267 210
rect 2359 206 2363 210
rect 2463 206 2467 210
rect 2543 206 2547 210
rect 111 193 115 197
rect 1327 193 1331 197
rect 1367 197 1371 201
rect 2583 197 2587 201
rect 335 183 339 187
rect 111 176 115 180
rect 183 175 187 179
rect 219 171 220 175
rect 220 171 223 175
rect 255 175 259 179
rect 291 171 292 175
rect 292 171 295 175
rect 343 175 347 179
rect 447 175 451 179
rect 483 171 484 175
rect 484 171 487 175
rect 551 175 555 179
rect 655 183 659 187
rect 663 175 667 179
rect 687 171 691 175
rect 775 175 779 179
rect 887 183 891 187
rect 1935 187 1939 191
rect 895 175 899 179
rect 931 171 932 175
rect 932 171 935 175
rect 1015 175 1019 179
rect 1039 171 1043 175
rect 1135 175 1139 179
rect 1255 175 1259 179
rect 1327 176 1331 180
rect 1367 180 1371 184
rect 1399 179 1403 183
rect 1435 175 1436 179
rect 1436 175 1439 179
rect 1463 179 1467 183
rect 1199 167 1203 171
rect 1499 175 1500 179
rect 1500 175 1503 179
rect 1543 179 1547 183
rect 1579 175 1580 179
rect 1580 175 1583 179
rect 1639 179 1643 183
rect 1675 175 1676 179
rect 1676 175 1679 179
rect 1735 179 1739 183
rect 1771 175 1772 179
rect 1772 175 1775 179
rect 1839 179 1843 183
rect 1871 175 1872 179
rect 1872 175 1875 179
rect 1943 179 1947 183
rect 1895 171 1899 175
rect 2047 179 2051 183
rect 2239 187 2243 191
rect 2151 179 2155 183
rect 2183 175 2184 179
rect 2184 175 2187 179
rect 2247 179 2251 183
rect 2159 167 2163 171
rect 2343 179 2347 183
rect 2447 179 2451 183
rect 2527 179 2531 183
rect 2583 180 2587 184
rect 2559 175 2560 179
rect 2560 175 2563 179
rect 2335 139 2339 143
rect 1367 128 1371 132
rect 1399 129 1403 133
rect 1447 131 1451 135
rect 1455 129 1459 133
rect 1503 131 1507 135
rect 1511 129 1515 133
rect 1559 131 1563 135
rect 1567 129 1571 133
rect 1623 131 1627 135
rect 1631 129 1635 133
rect 1703 131 1707 135
rect 1711 129 1715 133
rect 1783 131 1787 135
rect 1791 129 1795 133
rect 1823 131 1824 135
rect 1824 131 1827 135
rect 1871 129 1875 133
rect 1935 131 1939 135
rect 1943 129 1947 133
rect 2007 131 2011 135
rect 2015 129 2019 133
rect 2071 131 2075 135
rect 2079 129 2083 133
rect 2135 131 2139 135
rect 2143 129 2147 133
rect 2199 131 2203 135
rect 2207 129 2211 133
rect 2263 131 2267 135
rect 2271 129 2275 133
rect 2335 131 2339 135
rect 2343 129 2347 133
rect 2407 131 2411 135
rect 2415 129 2419 133
rect 2583 128 2587 132
rect 111 116 115 120
rect 143 117 147 121
rect 191 119 195 123
rect 199 117 203 121
rect 247 119 251 123
rect 255 117 259 121
rect 303 119 307 123
rect 311 117 315 121
rect 359 119 363 123
rect 367 117 371 121
rect 415 119 419 123
rect 423 117 427 121
rect 471 119 475 123
rect 479 117 483 121
rect 527 119 531 123
rect 535 117 539 121
rect 583 119 587 123
rect 591 117 595 121
rect 623 119 624 123
rect 624 119 627 123
rect 647 117 651 121
rect 695 119 699 123
rect 703 117 707 121
rect 751 119 755 123
rect 759 117 763 121
rect 815 119 819 123
rect 823 117 827 121
rect 879 119 883 123
rect 887 117 891 121
rect 943 119 947 123
rect 951 117 955 121
rect 1007 119 1011 123
rect 1015 117 1019 121
rect 1071 119 1075 123
rect 1079 117 1083 121
rect 1115 119 1116 123
rect 1116 119 1119 123
rect 1151 117 1155 121
rect 1207 119 1211 123
rect 1215 117 1219 121
rect 1263 119 1267 123
rect 1271 117 1275 121
rect 1327 116 1331 120
rect 1367 111 1371 115
rect 2583 111 2587 115
rect 111 99 115 103
rect 1327 99 1331 103
rect 1415 102 1419 106
rect 1471 102 1475 106
rect 1527 102 1531 106
rect 1583 102 1587 106
rect 1647 102 1651 106
rect 1727 102 1731 106
rect 1807 102 1811 106
rect 1887 102 1891 106
rect 1959 102 1963 106
rect 2031 102 2035 106
rect 2095 102 2099 106
rect 2159 102 2163 106
rect 2223 102 2227 106
rect 2287 102 2291 106
rect 2359 102 2363 106
rect 2431 102 2435 106
rect 159 90 163 94
rect 215 90 219 94
rect 271 90 275 94
rect 327 90 331 94
rect 383 90 387 94
rect 439 90 443 94
rect 495 90 499 94
rect 551 90 555 94
rect 607 90 611 94
rect 663 90 667 94
rect 719 90 723 94
rect 775 90 779 94
rect 839 90 843 94
rect 903 90 907 94
rect 967 90 971 94
rect 1031 90 1035 94
rect 1095 90 1099 94
rect 1167 90 1171 94
rect 1231 90 1235 94
rect 1447 95 1448 99
rect 1448 95 1451 99
rect 1503 95 1504 99
rect 1504 95 1507 99
rect 1559 95 1560 99
rect 1560 95 1563 99
rect 1623 95 1624 99
rect 1624 95 1627 99
rect 1703 95 1704 99
rect 1704 95 1707 99
rect 1783 95 1784 99
rect 1784 95 1787 99
rect 1895 95 1899 99
rect 1935 95 1936 99
rect 1936 95 1939 99
rect 2007 95 2008 99
rect 2008 95 2011 99
rect 2071 95 2072 99
rect 2072 95 2075 99
rect 2135 95 2136 99
rect 2136 95 2139 99
rect 2199 95 2200 99
rect 2200 95 2203 99
rect 2263 95 2264 99
rect 2264 95 2267 99
rect 2335 95 2336 99
rect 2336 95 2339 99
rect 2407 95 2408 99
rect 2408 95 2411 99
rect 1287 90 1291 94
rect 191 83 192 87
rect 192 83 195 87
rect 247 83 248 87
rect 248 83 251 87
rect 303 83 304 87
rect 304 83 307 87
rect 359 83 360 87
rect 360 83 363 87
rect 415 83 416 87
rect 416 83 419 87
rect 471 83 472 87
rect 472 83 475 87
rect 527 83 528 87
rect 528 83 531 87
rect 583 83 584 87
rect 584 83 587 87
rect 687 83 691 87
rect 695 83 696 87
rect 696 83 699 87
rect 751 83 752 87
rect 752 83 755 87
rect 815 83 816 87
rect 816 83 819 87
rect 879 83 880 87
rect 880 83 883 87
rect 943 83 944 87
rect 944 83 947 87
rect 1007 83 1008 87
rect 1008 83 1011 87
rect 1071 83 1072 87
rect 1072 83 1075 87
rect 1199 83 1203 87
rect 1207 83 1208 87
rect 1208 83 1211 87
rect 1263 83 1264 87
rect 1264 83 1267 87
<< m3 >>
rect 622 2643 628 2644
rect 734 2643 740 2644
rect 111 2642 115 2643
rect 111 2637 115 2638
rect 551 2642 555 2643
rect 551 2637 555 2638
rect 607 2642 611 2643
rect 622 2639 623 2643
rect 627 2639 628 2643
rect 622 2638 628 2639
rect 663 2642 667 2643
rect 607 2637 611 2638
rect 112 2622 114 2637
rect 552 2631 554 2637
rect 582 2635 588 2636
rect 582 2631 583 2635
rect 587 2631 588 2635
rect 608 2631 610 2637
rect 550 2630 556 2631
rect 582 2630 588 2631
rect 606 2630 612 2631
rect 550 2626 551 2630
rect 555 2626 556 2630
rect 550 2625 556 2626
rect 110 2621 116 2622
rect 110 2617 111 2621
rect 115 2617 116 2621
rect 110 2616 116 2617
rect 584 2612 586 2630
rect 606 2626 607 2630
rect 611 2626 612 2630
rect 606 2625 612 2626
rect 582 2611 588 2612
rect 582 2607 583 2611
rect 587 2607 588 2611
rect 582 2606 588 2607
rect 110 2604 116 2605
rect 110 2600 111 2604
rect 115 2600 116 2604
rect 110 2599 116 2600
rect 534 2603 540 2604
rect 534 2599 535 2603
rect 539 2599 540 2603
rect 590 2603 596 2604
rect 112 2587 114 2599
rect 534 2598 540 2599
rect 558 2599 564 2600
rect 536 2587 538 2598
rect 558 2595 559 2599
rect 563 2595 564 2599
rect 590 2599 591 2603
rect 595 2599 596 2603
rect 624 2600 626 2638
rect 663 2637 667 2638
rect 719 2642 723 2643
rect 734 2639 735 2643
rect 739 2639 740 2643
rect 734 2638 740 2639
rect 775 2642 779 2643
rect 719 2637 723 2638
rect 664 2631 666 2637
rect 694 2635 700 2636
rect 694 2631 695 2635
rect 699 2631 700 2635
rect 720 2631 722 2637
rect 662 2630 668 2631
rect 694 2630 700 2631
rect 718 2630 724 2631
rect 662 2626 663 2630
rect 667 2626 668 2630
rect 662 2625 668 2626
rect 696 2612 698 2630
rect 718 2626 719 2630
rect 723 2626 724 2630
rect 718 2625 724 2626
rect 694 2611 700 2612
rect 694 2607 695 2611
rect 699 2607 700 2611
rect 694 2606 700 2607
rect 646 2603 652 2604
rect 590 2598 596 2599
rect 622 2599 628 2600
rect 558 2594 564 2595
rect 111 2586 115 2587
rect 111 2581 115 2582
rect 215 2586 219 2587
rect 215 2581 219 2582
rect 271 2586 275 2587
rect 271 2581 275 2582
rect 327 2586 331 2587
rect 327 2581 331 2582
rect 383 2586 387 2587
rect 383 2581 387 2582
rect 439 2586 443 2587
rect 439 2581 443 2582
rect 495 2586 499 2587
rect 495 2581 499 2582
rect 535 2586 539 2587
rect 535 2581 539 2582
rect 551 2586 555 2587
rect 551 2581 555 2582
rect 112 2569 114 2581
rect 216 2570 218 2581
rect 238 2579 244 2580
rect 238 2575 239 2579
rect 243 2575 244 2579
rect 238 2574 244 2575
rect 214 2569 220 2570
rect 110 2568 116 2569
rect 110 2564 111 2568
rect 115 2564 116 2568
rect 214 2565 215 2569
rect 219 2565 220 2569
rect 214 2564 220 2565
rect 110 2563 116 2564
rect 110 2551 116 2552
rect 110 2547 111 2551
rect 115 2547 116 2551
rect 110 2546 116 2547
rect 112 2527 114 2546
rect 230 2542 236 2543
rect 230 2538 231 2542
rect 235 2538 236 2542
rect 230 2537 236 2538
rect 232 2527 234 2537
rect 240 2536 242 2574
rect 262 2571 268 2572
rect 262 2567 263 2571
rect 267 2567 268 2571
rect 272 2570 274 2581
rect 318 2571 324 2572
rect 262 2566 268 2567
rect 270 2569 276 2570
rect 264 2536 266 2566
rect 270 2565 271 2569
rect 275 2565 276 2569
rect 318 2567 319 2571
rect 323 2567 324 2571
rect 328 2570 330 2581
rect 354 2571 360 2572
rect 318 2566 324 2567
rect 326 2569 332 2570
rect 270 2564 276 2565
rect 286 2542 292 2543
rect 286 2538 287 2542
rect 291 2538 292 2542
rect 286 2537 292 2538
rect 238 2535 244 2536
rect 238 2531 239 2535
rect 243 2531 244 2535
rect 238 2530 244 2531
rect 262 2535 268 2536
rect 262 2531 263 2535
rect 267 2531 268 2535
rect 262 2530 268 2531
rect 288 2527 290 2537
rect 320 2536 322 2566
rect 326 2565 327 2569
rect 331 2565 332 2569
rect 354 2567 355 2571
rect 359 2567 360 2571
rect 384 2570 386 2581
rect 440 2570 442 2581
rect 496 2570 498 2581
rect 526 2579 532 2580
rect 526 2575 527 2579
rect 531 2575 532 2579
rect 526 2574 532 2575
rect 354 2566 360 2567
rect 382 2569 388 2570
rect 326 2564 332 2565
rect 342 2542 348 2543
rect 342 2538 343 2542
rect 347 2538 348 2542
rect 342 2537 348 2538
rect 318 2535 324 2536
rect 318 2531 319 2535
rect 323 2531 324 2535
rect 318 2530 324 2531
rect 344 2527 346 2537
rect 111 2526 115 2527
rect 111 2521 115 2522
rect 231 2526 235 2527
rect 231 2521 235 2522
rect 287 2526 291 2527
rect 287 2521 291 2522
rect 343 2526 347 2527
rect 356 2524 358 2566
rect 382 2565 383 2569
rect 387 2565 388 2569
rect 382 2564 388 2565
rect 438 2569 444 2570
rect 438 2565 439 2569
rect 443 2565 444 2569
rect 438 2564 444 2565
rect 494 2569 500 2570
rect 494 2565 495 2569
rect 499 2565 500 2569
rect 494 2564 500 2565
rect 398 2542 404 2543
rect 398 2538 399 2542
rect 403 2538 404 2542
rect 398 2537 404 2538
rect 454 2542 460 2543
rect 454 2538 455 2542
rect 459 2538 460 2542
rect 454 2537 460 2538
rect 510 2542 516 2543
rect 510 2538 511 2542
rect 515 2538 516 2542
rect 510 2537 516 2538
rect 400 2527 402 2537
rect 456 2527 458 2537
rect 512 2527 514 2537
rect 528 2536 530 2574
rect 552 2570 554 2581
rect 550 2569 556 2570
rect 550 2565 551 2569
rect 555 2565 556 2569
rect 550 2564 556 2565
rect 560 2536 562 2594
rect 592 2587 594 2598
rect 622 2595 623 2599
rect 627 2595 628 2599
rect 646 2599 647 2603
rect 651 2599 652 2603
rect 646 2598 652 2599
rect 702 2603 708 2604
rect 702 2599 703 2603
rect 707 2599 708 2603
rect 736 2600 738 2638
rect 775 2637 779 2638
rect 1327 2642 1331 2643
rect 1622 2639 1628 2640
rect 1734 2639 1740 2640
rect 1838 2639 1844 2640
rect 1958 2639 1964 2640
rect 2182 2639 2188 2640
rect 1327 2637 1331 2638
rect 1367 2638 1371 2639
rect 750 2635 756 2636
rect 750 2631 751 2635
rect 755 2631 756 2635
rect 776 2631 778 2637
rect 750 2630 756 2631
rect 774 2630 780 2631
rect 702 2598 708 2599
rect 734 2599 740 2600
rect 622 2594 628 2595
rect 648 2587 650 2598
rect 704 2587 706 2598
rect 734 2595 735 2599
rect 739 2595 740 2599
rect 734 2594 740 2595
rect 591 2586 595 2587
rect 591 2581 595 2582
rect 607 2586 611 2587
rect 607 2581 611 2582
rect 647 2586 651 2587
rect 647 2581 651 2582
rect 663 2586 667 2587
rect 663 2581 667 2582
rect 703 2586 707 2587
rect 703 2581 707 2582
rect 719 2586 723 2587
rect 719 2581 723 2582
rect 598 2571 604 2572
rect 598 2567 599 2571
rect 603 2567 604 2571
rect 608 2570 610 2581
rect 664 2570 666 2581
rect 686 2579 692 2580
rect 686 2575 687 2579
rect 691 2575 692 2579
rect 686 2574 692 2575
rect 598 2566 604 2567
rect 606 2569 612 2570
rect 566 2542 572 2543
rect 566 2538 567 2542
rect 571 2538 572 2542
rect 566 2537 572 2538
rect 526 2535 532 2536
rect 526 2531 527 2535
rect 531 2531 532 2535
rect 526 2530 532 2531
rect 558 2535 564 2536
rect 558 2531 559 2535
rect 563 2531 564 2535
rect 558 2530 564 2531
rect 568 2527 570 2537
rect 600 2536 602 2566
rect 606 2565 607 2569
rect 611 2565 612 2569
rect 606 2564 612 2565
rect 662 2569 668 2570
rect 662 2565 663 2569
rect 667 2565 668 2569
rect 662 2564 668 2565
rect 622 2542 628 2543
rect 622 2538 623 2542
rect 627 2538 628 2542
rect 622 2537 628 2538
rect 678 2542 684 2543
rect 678 2538 679 2542
rect 683 2538 684 2542
rect 678 2537 684 2538
rect 598 2535 604 2536
rect 598 2531 599 2535
rect 603 2531 604 2535
rect 598 2530 604 2531
rect 624 2527 626 2537
rect 680 2527 682 2537
rect 688 2536 690 2574
rect 710 2571 716 2572
rect 710 2567 711 2571
rect 715 2567 716 2571
rect 720 2570 722 2581
rect 752 2572 754 2630
rect 774 2626 775 2630
rect 779 2626 780 2630
rect 774 2625 780 2626
rect 1328 2622 1330 2637
rect 1367 2633 1371 2634
rect 1551 2638 1555 2639
rect 1551 2633 1555 2634
rect 1607 2638 1611 2639
rect 1622 2635 1623 2639
rect 1627 2635 1628 2639
rect 1622 2634 1628 2635
rect 1663 2638 1667 2639
rect 1607 2633 1611 2634
rect 1326 2621 1332 2622
rect 1326 2617 1327 2621
rect 1331 2617 1332 2621
rect 1368 2618 1370 2633
rect 1552 2627 1554 2633
rect 1582 2631 1588 2632
rect 1582 2627 1583 2631
rect 1587 2627 1588 2631
rect 1608 2627 1610 2633
rect 1550 2626 1556 2627
rect 1582 2626 1588 2627
rect 1606 2626 1612 2627
rect 1550 2622 1551 2626
rect 1555 2622 1556 2626
rect 1550 2621 1556 2622
rect 1326 2616 1332 2617
rect 1366 2617 1372 2618
rect 1366 2613 1367 2617
rect 1371 2613 1372 2617
rect 1366 2612 1372 2613
rect 1584 2608 1586 2626
rect 1606 2622 1607 2626
rect 1611 2622 1612 2626
rect 1606 2621 1612 2622
rect 1582 2607 1588 2608
rect 1326 2604 1332 2605
rect 758 2603 764 2604
rect 758 2599 759 2603
rect 763 2599 764 2603
rect 1326 2600 1327 2604
rect 1331 2600 1332 2604
rect 1582 2603 1583 2607
rect 1587 2603 1588 2607
rect 1582 2602 1588 2603
rect 1326 2599 1332 2600
rect 1366 2600 1372 2601
rect 758 2598 764 2599
rect 760 2587 762 2598
rect 1328 2587 1330 2599
rect 1366 2596 1367 2600
rect 1371 2596 1372 2600
rect 1366 2595 1372 2596
rect 1534 2599 1540 2600
rect 1534 2595 1535 2599
rect 1539 2595 1540 2599
rect 759 2586 763 2587
rect 759 2581 763 2582
rect 775 2586 779 2587
rect 775 2581 779 2582
rect 831 2586 835 2587
rect 831 2581 835 2582
rect 887 2586 891 2587
rect 887 2581 891 2582
rect 943 2586 947 2587
rect 943 2581 947 2582
rect 999 2586 1003 2587
rect 999 2581 1003 2582
rect 1055 2586 1059 2587
rect 1055 2581 1059 2582
rect 1111 2586 1115 2587
rect 1111 2581 1115 2582
rect 1327 2586 1331 2587
rect 1368 2583 1370 2595
rect 1534 2594 1540 2595
rect 1590 2599 1596 2600
rect 1590 2595 1591 2599
rect 1595 2595 1596 2599
rect 1624 2596 1626 2634
rect 1663 2633 1667 2634
rect 1719 2638 1723 2639
rect 1734 2635 1735 2639
rect 1739 2635 1740 2639
rect 1734 2634 1740 2635
rect 1775 2638 1779 2639
rect 1719 2633 1723 2634
rect 1664 2627 1666 2633
rect 1694 2631 1700 2632
rect 1694 2627 1695 2631
rect 1699 2627 1700 2631
rect 1720 2627 1722 2633
rect 1662 2626 1668 2627
rect 1694 2626 1700 2627
rect 1718 2626 1724 2627
rect 1662 2622 1663 2626
rect 1667 2622 1668 2626
rect 1662 2621 1668 2622
rect 1696 2608 1698 2626
rect 1718 2622 1719 2626
rect 1723 2622 1724 2626
rect 1718 2621 1724 2622
rect 1694 2607 1700 2608
rect 1694 2603 1695 2607
rect 1699 2603 1700 2607
rect 1694 2602 1700 2603
rect 1646 2599 1652 2600
rect 1590 2594 1596 2595
rect 1622 2595 1628 2596
rect 1446 2591 1452 2592
rect 1446 2587 1447 2591
rect 1451 2587 1452 2591
rect 1446 2586 1452 2587
rect 1327 2581 1331 2582
rect 1367 2582 1371 2583
rect 750 2571 756 2572
rect 710 2566 716 2567
rect 718 2569 724 2570
rect 712 2536 714 2566
rect 718 2565 719 2569
rect 723 2565 724 2569
rect 750 2567 751 2571
rect 755 2567 756 2571
rect 776 2570 778 2581
rect 832 2570 834 2581
rect 888 2570 890 2581
rect 944 2570 946 2581
rect 974 2579 980 2580
rect 974 2575 975 2579
rect 979 2575 980 2579
rect 974 2574 980 2575
rect 750 2566 756 2567
rect 774 2569 780 2570
rect 718 2564 724 2565
rect 774 2565 775 2569
rect 779 2565 780 2569
rect 774 2564 780 2565
rect 830 2569 836 2570
rect 830 2565 831 2569
rect 835 2565 836 2569
rect 830 2564 836 2565
rect 886 2569 892 2570
rect 886 2565 887 2569
rect 891 2565 892 2569
rect 886 2564 892 2565
rect 942 2569 948 2570
rect 942 2565 943 2569
rect 947 2565 948 2569
rect 942 2564 948 2565
rect 734 2542 740 2543
rect 734 2538 735 2542
rect 739 2538 740 2542
rect 734 2537 740 2538
rect 790 2542 796 2543
rect 790 2538 791 2542
rect 795 2538 796 2542
rect 790 2537 796 2538
rect 846 2542 852 2543
rect 846 2538 847 2542
rect 851 2538 852 2542
rect 846 2537 852 2538
rect 902 2542 908 2543
rect 902 2538 903 2542
rect 907 2538 908 2542
rect 902 2537 908 2538
rect 958 2542 964 2543
rect 958 2538 959 2542
rect 963 2538 964 2542
rect 958 2537 964 2538
rect 686 2535 692 2536
rect 686 2531 687 2535
rect 691 2531 692 2535
rect 686 2530 692 2531
rect 710 2535 716 2536
rect 710 2531 711 2535
rect 715 2531 716 2535
rect 710 2530 716 2531
rect 736 2527 738 2537
rect 792 2527 794 2537
rect 848 2527 850 2537
rect 904 2527 906 2537
rect 960 2527 962 2537
rect 976 2536 978 2574
rect 1000 2570 1002 2581
rect 1046 2571 1052 2572
rect 998 2569 1004 2570
rect 998 2565 999 2569
rect 1003 2565 1004 2569
rect 1046 2567 1047 2571
rect 1051 2567 1052 2571
rect 1056 2570 1058 2581
rect 1102 2571 1108 2572
rect 1046 2566 1052 2567
rect 1054 2569 1060 2570
rect 998 2564 1004 2565
rect 1014 2542 1020 2543
rect 1014 2538 1015 2542
rect 1019 2538 1020 2542
rect 1014 2537 1020 2538
rect 974 2535 980 2536
rect 974 2531 975 2535
rect 979 2531 980 2535
rect 974 2530 980 2531
rect 1016 2527 1018 2537
rect 1048 2536 1050 2566
rect 1054 2565 1055 2569
rect 1059 2565 1060 2569
rect 1102 2567 1103 2571
rect 1107 2567 1108 2571
rect 1112 2570 1114 2581
rect 1102 2566 1108 2567
rect 1110 2569 1116 2570
rect 1328 2569 1330 2581
rect 1367 2577 1371 2578
rect 1439 2582 1443 2583
rect 1439 2577 1443 2578
rect 1054 2564 1060 2565
rect 1070 2542 1076 2543
rect 1070 2538 1071 2542
rect 1075 2538 1076 2542
rect 1070 2537 1076 2538
rect 1046 2535 1052 2536
rect 1046 2531 1047 2535
rect 1051 2531 1052 2535
rect 1046 2530 1052 2531
rect 1022 2527 1028 2528
rect 1072 2527 1074 2537
rect 1104 2536 1106 2566
rect 1110 2565 1111 2569
rect 1115 2565 1116 2569
rect 1110 2564 1116 2565
rect 1326 2568 1332 2569
rect 1326 2564 1327 2568
rect 1331 2564 1332 2568
rect 1368 2565 1370 2577
rect 1440 2566 1442 2577
rect 1438 2565 1444 2566
rect 1326 2563 1332 2564
rect 1366 2564 1372 2565
rect 1366 2560 1367 2564
rect 1371 2560 1372 2564
rect 1438 2561 1439 2565
rect 1443 2561 1444 2565
rect 1438 2560 1444 2561
rect 1366 2559 1372 2560
rect 1326 2551 1332 2552
rect 1326 2547 1327 2551
rect 1331 2547 1332 2551
rect 1326 2546 1332 2547
rect 1366 2547 1372 2548
rect 1126 2542 1132 2543
rect 1126 2538 1127 2542
rect 1131 2538 1132 2542
rect 1126 2537 1132 2538
rect 1102 2535 1108 2536
rect 1102 2531 1103 2535
rect 1107 2531 1108 2535
rect 1102 2530 1108 2531
rect 1128 2527 1130 2537
rect 1328 2527 1330 2546
rect 1366 2543 1367 2547
rect 1371 2543 1372 2547
rect 1366 2542 1372 2543
rect 367 2526 371 2527
rect 343 2521 347 2522
rect 354 2523 360 2524
rect 112 2506 114 2521
rect 354 2519 355 2523
rect 359 2519 360 2523
rect 367 2521 371 2522
rect 399 2526 403 2527
rect 399 2521 403 2522
rect 423 2526 427 2527
rect 423 2521 427 2522
rect 455 2526 459 2527
rect 455 2521 459 2522
rect 487 2526 491 2527
rect 487 2521 491 2522
rect 511 2526 515 2527
rect 511 2521 515 2522
rect 551 2526 555 2527
rect 551 2521 555 2522
rect 567 2526 571 2527
rect 567 2521 571 2522
rect 615 2526 619 2527
rect 615 2521 619 2522
rect 623 2526 627 2527
rect 623 2521 627 2522
rect 679 2526 683 2527
rect 679 2521 683 2522
rect 735 2526 739 2527
rect 735 2521 739 2522
rect 743 2526 747 2527
rect 743 2521 747 2522
rect 791 2526 795 2527
rect 791 2521 795 2522
rect 807 2526 811 2527
rect 807 2521 811 2522
rect 847 2526 851 2527
rect 847 2521 851 2522
rect 871 2526 875 2527
rect 871 2521 875 2522
rect 903 2526 907 2527
rect 903 2521 907 2522
rect 943 2526 947 2527
rect 943 2521 947 2522
rect 959 2526 963 2527
rect 959 2521 963 2522
rect 1015 2526 1019 2527
rect 1022 2523 1023 2527
rect 1027 2523 1028 2527
rect 1022 2522 1028 2523
rect 1071 2526 1075 2527
rect 1015 2521 1019 2522
rect 354 2518 360 2519
rect 368 2515 370 2521
rect 386 2519 392 2520
rect 386 2515 387 2519
rect 391 2515 392 2519
rect 424 2515 426 2521
rect 442 2519 448 2520
rect 442 2515 443 2519
rect 447 2515 448 2519
rect 488 2515 490 2521
rect 552 2515 554 2521
rect 616 2515 618 2521
rect 654 2519 660 2520
rect 654 2515 655 2519
rect 659 2515 660 2519
rect 680 2515 682 2521
rect 706 2519 712 2520
rect 706 2515 707 2519
rect 711 2515 712 2519
rect 744 2515 746 2521
rect 758 2519 764 2520
rect 758 2515 759 2519
rect 763 2515 764 2519
rect 808 2515 810 2521
rect 872 2515 874 2521
rect 944 2515 946 2521
rect 978 2519 984 2520
rect 978 2515 979 2519
rect 983 2515 984 2519
rect 1016 2515 1018 2521
rect 366 2514 372 2515
rect 386 2514 392 2515
rect 422 2514 428 2515
rect 442 2514 448 2515
rect 486 2514 492 2515
rect 366 2510 367 2514
rect 371 2510 372 2514
rect 366 2509 372 2510
rect 110 2505 116 2506
rect 110 2501 111 2505
rect 115 2501 116 2505
rect 110 2500 116 2501
rect 110 2488 116 2489
rect 110 2484 111 2488
rect 115 2484 116 2488
rect 110 2483 116 2484
rect 350 2487 356 2488
rect 350 2483 351 2487
rect 355 2483 356 2487
rect 388 2484 390 2514
rect 422 2510 423 2514
rect 427 2510 428 2514
rect 422 2509 428 2510
rect 406 2487 412 2488
rect 112 2467 114 2483
rect 350 2482 356 2483
rect 386 2483 392 2484
rect 352 2467 354 2482
rect 386 2479 387 2483
rect 391 2479 392 2483
rect 406 2483 407 2487
rect 411 2483 412 2487
rect 444 2484 446 2514
rect 486 2510 487 2514
rect 491 2510 492 2514
rect 486 2509 492 2510
rect 550 2514 556 2515
rect 550 2510 551 2514
rect 555 2510 556 2514
rect 550 2509 556 2510
rect 614 2514 620 2515
rect 654 2514 660 2515
rect 678 2514 684 2515
rect 706 2514 712 2515
rect 742 2514 748 2515
rect 758 2514 764 2515
rect 806 2514 812 2515
rect 614 2510 615 2514
rect 619 2510 620 2514
rect 614 2509 620 2510
rect 656 2496 658 2514
rect 678 2510 679 2514
rect 683 2510 684 2514
rect 678 2509 684 2510
rect 654 2495 660 2496
rect 654 2491 655 2495
rect 659 2491 660 2495
rect 654 2490 660 2491
rect 470 2487 476 2488
rect 406 2482 412 2483
rect 442 2483 448 2484
rect 386 2478 392 2479
rect 408 2467 410 2482
rect 442 2479 443 2483
rect 447 2479 448 2483
rect 470 2483 471 2487
rect 475 2483 476 2487
rect 470 2482 476 2483
rect 534 2487 540 2488
rect 534 2483 535 2487
rect 539 2483 540 2487
rect 534 2482 540 2483
rect 598 2487 604 2488
rect 598 2483 599 2487
rect 603 2483 604 2487
rect 662 2487 668 2488
rect 598 2482 604 2483
rect 622 2483 628 2484
rect 442 2478 448 2479
rect 472 2467 474 2482
rect 536 2467 538 2482
rect 600 2467 602 2482
rect 622 2479 623 2483
rect 627 2479 628 2483
rect 662 2483 663 2487
rect 667 2483 668 2487
rect 708 2484 710 2514
rect 742 2510 743 2514
rect 747 2510 748 2514
rect 742 2509 748 2510
rect 726 2487 732 2488
rect 662 2482 668 2483
rect 706 2483 712 2484
rect 622 2478 628 2479
rect 111 2466 115 2467
rect 111 2461 115 2462
rect 271 2466 275 2467
rect 271 2461 275 2462
rect 335 2466 339 2467
rect 335 2461 339 2462
rect 351 2466 355 2467
rect 351 2461 355 2462
rect 399 2466 403 2467
rect 399 2461 403 2462
rect 407 2466 411 2467
rect 407 2461 411 2462
rect 471 2466 475 2467
rect 471 2461 475 2462
rect 535 2466 539 2467
rect 535 2461 539 2462
rect 551 2466 555 2467
rect 551 2461 555 2462
rect 599 2466 603 2467
rect 599 2461 603 2462
rect 112 2449 114 2461
rect 272 2450 274 2461
rect 278 2459 284 2460
rect 278 2455 279 2459
rect 283 2455 284 2459
rect 278 2454 284 2455
rect 270 2449 276 2450
rect 110 2448 116 2449
rect 110 2444 111 2448
rect 115 2444 116 2448
rect 270 2445 271 2449
rect 275 2445 276 2449
rect 270 2444 276 2445
rect 110 2443 116 2444
rect 110 2431 116 2432
rect 110 2427 111 2431
rect 115 2427 116 2431
rect 110 2426 116 2427
rect 112 2407 114 2426
rect 280 2416 282 2454
rect 326 2451 332 2452
rect 326 2447 327 2451
rect 331 2447 332 2451
rect 336 2450 338 2461
rect 390 2451 396 2452
rect 326 2446 332 2447
rect 334 2449 340 2450
rect 286 2422 292 2423
rect 286 2418 287 2422
rect 291 2418 292 2422
rect 286 2417 292 2418
rect 278 2415 284 2416
rect 278 2411 279 2415
rect 283 2411 284 2415
rect 278 2410 284 2411
rect 288 2407 290 2417
rect 328 2416 330 2446
rect 334 2445 335 2449
rect 339 2445 340 2449
rect 390 2447 391 2451
rect 395 2447 396 2451
rect 400 2450 402 2461
rect 422 2451 428 2452
rect 390 2446 396 2447
rect 398 2449 404 2450
rect 334 2444 340 2445
rect 350 2422 356 2423
rect 350 2418 351 2422
rect 355 2418 356 2422
rect 350 2417 356 2418
rect 326 2415 332 2416
rect 326 2411 327 2415
rect 331 2411 332 2415
rect 326 2410 332 2411
rect 352 2407 354 2417
rect 392 2416 394 2446
rect 398 2445 399 2449
rect 403 2445 404 2449
rect 422 2447 423 2451
rect 427 2447 428 2451
rect 472 2450 474 2461
rect 552 2450 554 2461
rect 422 2446 428 2447
rect 470 2449 476 2450
rect 398 2444 404 2445
rect 414 2422 420 2423
rect 414 2418 415 2422
rect 419 2418 420 2422
rect 414 2417 420 2418
rect 390 2415 396 2416
rect 390 2411 391 2415
rect 395 2411 396 2415
rect 390 2410 396 2411
rect 416 2407 418 2417
rect 111 2406 115 2407
rect 111 2401 115 2402
rect 247 2406 251 2407
rect 247 2401 251 2402
rect 287 2406 291 2407
rect 287 2401 291 2402
rect 335 2406 339 2407
rect 335 2401 339 2402
rect 351 2406 355 2407
rect 351 2401 355 2402
rect 415 2406 419 2407
rect 415 2401 419 2402
rect 112 2386 114 2401
rect 238 2399 244 2400
rect 238 2395 239 2399
rect 243 2395 244 2399
rect 248 2395 250 2401
rect 266 2399 272 2400
rect 266 2395 267 2399
rect 271 2395 272 2399
rect 336 2395 338 2401
rect 424 2400 426 2446
rect 470 2445 471 2449
rect 475 2445 476 2449
rect 470 2444 476 2445
rect 550 2449 556 2450
rect 550 2445 551 2449
rect 555 2445 556 2449
rect 550 2444 556 2445
rect 486 2422 492 2423
rect 486 2418 487 2422
rect 491 2418 492 2422
rect 486 2417 492 2418
rect 566 2422 572 2423
rect 566 2418 567 2422
rect 571 2418 572 2422
rect 566 2417 572 2418
rect 488 2407 490 2417
rect 568 2407 570 2417
rect 624 2416 626 2478
rect 664 2467 666 2482
rect 706 2479 707 2483
rect 711 2479 712 2483
rect 726 2483 727 2487
rect 731 2483 732 2487
rect 760 2484 762 2514
rect 806 2510 807 2514
rect 811 2510 812 2514
rect 806 2509 812 2510
rect 870 2514 876 2515
rect 870 2510 871 2514
rect 875 2510 876 2514
rect 870 2509 876 2510
rect 942 2514 948 2515
rect 978 2514 984 2515
rect 1014 2514 1020 2515
rect 942 2510 943 2514
rect 947 2510 948 2514
rect 942 2509 948 2510
rect 980 2488 982 2514
rect 1014 2510 1015 2514
rect 1019 2510 1020 2514
rect 1014 2509 1020 2510
rect 790 2487 796 2488
rect 726 2482 732 2483
rect 758 2483 764 2484
rect 706 2478 712 2479
rect 728 2467 730 2482
rect 758 2479 759 2483
rect 763 2479 764 2483
rect 790 2483 791 2487
rect 795 2483 796 2487
rect 790 2482 796 2483
rect 854 2487 860 2488
rect 854 2483 855 2487
rect 859 2483 860 2487
rect 854 2482 860 2483
rect 926 2487 932 2488
rect 926 2483 927 2487
rect 931 2483 932 2487
rect 926 2482 932 2483
rect 978 2487 984 2488
rect 978 2483 979 2487
rect 983 2483 984 2487
rect 978 2482 984 2483
rect 998 2487 1004 2488
rect 998 2483 999 2487
rect 1003 2483 1004 2487
rect 1024 2484 1026 2522
rect 1071 2521 1075 2522
rect 1127 2526 1131 2527
rect 1127 2521 1131 2522
rect 1327 2526 1331 2527
rect 1327 2521 1331 2522
rect 1328 2506 1330 2521
rect 1368 2519 1370 2542
rect 1448 2532 1450 2586
rect 1536 2583 1538 2594
rect 1592 2583 1594 2594
rect 1622 2591 1623 2595
rect 1627 2591 1628 2595
rect 1646 2595 1647 2599
rect 1651 2595 1652 2599
rect 1646 2594 1652 2595
rect 1702 2599 1708 2600
rect 1702 2595 1703 2599
rect 1707 2595 1708 2599
rect 1736 2596 1738 2634
rect 1775 2633 1779 2634
rect 1831 2638 1835 2639
rect 1838 2635 1839 2639
rect 1843 2635 1844 2639
rect 1838 2634 1844 2635
rect 1887 2638 1891 2639
rect 1831 2633 1835 2634
rect 1776 2627 1778 2633
rect 1806 2631 1812 2632
rect 1806 2627 1807 2631
rect 1811 2627 1812 2631
rect 1832 2627 1834 2633
rect 1774 2626 1780 2627
rect 1806 2626 1812 2627
rect 1830 2626 1836 2627
rect 1774 2622 1775 2626
rect 1779 2622 1780 2626
rect 1774 2621 1780 2622
rect 1808 2608 1810 2626
rect 1830 2622 1831 2626
rect 1835 2622 1836 2626
rect 1830 2621 1836 2622
rect 1806 2607 1812 2608
rect 1806 2603 1807 2607
rect 1811 2603 1812 2607
rect 1806 2602 1812 2603
rect 1758 2599 1764 2600
rect 1702 2594 1708 2595
rect 1734 2595 1740 2596
rect 1622 2590 1628 2591
rect 1648 2583 1650 2594
rect 1704 2583 1706 2594
rect 1734 2591 1735 2595
rect 1739 2591 1740 2595
rect 1758 2595 1759 2599
rect 1763 2595 1764 2599
rect 1758 2594 1764 2595
rect 1814 2599 1820 2600
rect 1814 2595 1815 2599
rect 1819 2595 1820 2599
rect 1840 2596 1842 2634
rect 1887 2633 1891 2634
rect 1943 2638 1947 2639
rect 1958 2635 1959 2639
rect 1963 2635 1964 2639
rect 1958 2634 1964 2635
rect 1999 2638 2003 2639
rect 1943 2633 1947 2634
rect 1888 2627 1890 2633
rect 1918 2631 1924 2632
rect 1918 2627 1919 2631
rect 1923 2627 1924 2631
rect 1944 2627 1946 2633
rect 1886 2626 1892 2627
rect 1918 2626 1924 2627
rect 1942 2626 1948 2627
rect 1886 2622 1887 2626
rect 1891 2622 1892 2626
rect 1886 2621 1892 2622
rect 1920 2608 1922 2626
rect 1942 2622 1943 2626
rect 1947 2622 1948 2626
rect 1942 2621 1948 2622
rect 1918 2607 1924 2608
rect 1918 2603 1919 2607
rect 1923 2603 1924 2607
rect 1918 2602 1924 2603
rect 1870 2599 1876 2600
rect 1814 2594 1820 2595
rect 1838 2595 1844 2596
rect 1734 2590 1740 2591
rect 1760 2583 1762 2594
rect 1816 2583 1818 2594
rect 1838 2591 1839 2595
rect 1843 2591 1844 2595
rect 1870 2595 1871 2599
rect 1875 2595 1876 2599
rect 1870 2594 1876 2595
rect 1926 2599 1932 2600
rect 1926 2595 1927 2599
rect 1931 2595 1932 2599
rect 1960 2596 1962 2634
rect 1999 2633 2003 2634
rect 2055 2638 2059 2639
rect 2055 2633 2059 2634
rect 2111 2638 2115 2639
rect 2111 2633 2115 2634
rect 2167 2638 2171 2639
rect 2182 2635 2183 2639
rect 2187 2635 2188 2639
rect 2182 2634 2188 2635
rect 2583 2638 2587 2639
rect 2167 2633 2171 2634
rect 2000 2627 2002 2633
rect 2026 2631 2032 2632
rect 2026 2627 2027 2631
rect 2031 2627 2032 2631
rect 2056 2627 2058 2633
rect 2074 2631 2080 2632
rect 2074 2627 2075 2631
rect 2079 2627 2080 2631
rect 2112 2627 2114 2633
rect 2130 2631 2136 2632
rect 2130 2627 2131 2631
rect 2135 2627 2136 2631
rect 2168 2627 2170 2633
rect 1998 2626 2004 2627
rect 2026 2626 2032 2627
rect 2054 2626 2060 2627
rect 2074 2626 2080 2627
rect 2110 2626 2116 2627
rect 2130 2626 2136 2627
rect 2166 2626 2172 2627
rect 1998 2622 1999 2626
rect 2003 2622 2004 2626
rect 1998 2621 2004 2622
rect 1982 2599 1988 2600
rect 1926 2594 1932 2595
rect 1958 2595 1964 2596
rect 1838 2590 1844 2591
rect 1872 2583 1874 2594
rect 1928 2583 1930 2594
rect 1958 2591 1959 2595
rect 1963 2591 1964 2595
rect 1982 2595 1983 2599
rect 1987 2595 1988 2599
rect 1982 2594 1988 2595
rect 1958 2590 1964 2591
rect 1984 2583 1986 2594
rect 1535 2582 1539 2583
rect 1535 2577 1539 2578
rect 1543 2582 1547 2583
rect 1543 2577 1547 2578
rect 1591 2582 1595 2583
rect 1591 2577 1595 2578
rect 1647 2582 1651 2583
rect 1647 2577 1651 2578
rect 1655 2582 1659 2583
rect 1655 2577 1659 2578
rect 1703 2582 1707 2583
rect 1703 2577 1707 2578
rect 1759 2582 1763 2583
rect 1759 2577 1763 2578
rect 1767 2582 1771 2583
rect 1767 2577 1771 2578
rect 1815 2582 1819 2583
rect 1815 2577 1819 2578
rect 1871 2582 1875 2583
rect 1871 2577 1875 2578
rect 1879 2582 1883 2583
rect 1879 2577 1883 2578
rect 1927 2582 1931 2583
rect 1927 2577 1931 2578
rect 1983 2582 1987 2583
rect 1983 2577 1987 2578
rect 1991 2582 1995 2583
rect 1991 2577 1995 2578
rect 1534 2567 1540 2568
rect 1534 2563 1535 2567
rect 1539 2563 1540 2567
rect 1544 2566 1546 2577
rect 1646 2567 1652 2568
rect 1534 2562 1540 2563
rect 1542 2565 1548 2566
rect 1454 2538 1460 2539
rect 1454 2534 1455 2538
rect 1459 2534 1460 2538
rect 1454 2533 1460 2534
rect 1446 2531 1452 2532
rect 1446 2527 1447 2531
rect 1451 2527 1452 2531
rect 1446 2526 1452 2527
rect 1456 2519 1458 2533
rect 1536 2532 1538 2562
rect 1542 2561 1543 2565
rect 1547 2561 1548 2565
rect 1646 2563 1647 2567
rect 1651 2563 1652 2567
rect 1656 2566 1658 2577
rect 1758 2567 1764 2568
rect 1646 2562 1652 2563
rect 1654 2565 1660 2566
rect 1542 2560 1548 2561
rect 1558 2538 1564 2539
rect 1558 2534 1559 2538
rect 1563 2534 1564 2538
rect 1558 2533 1564 2534
rect 1543 2532 1547 2533
rect 1534 2531 1540 2532
rect 1534 2527 1535 2531
rect 1539 2527 1540 2531
rect 1543 2527 1547 2528
rect 1534 2526 1540 2527
rect 1367 2518 1371 2519
rect 1367 2513 1371 2514
rect 1455 2518 1459 2519
rect 1455 2513 1459 2514
rect 1326 2505 1332 2506
rect 1326 2501 1327 2505
rect 1331 2501 1332 2505
rect 1326 2500 1332 2501
rect 1368 2498 1370 2513
rect 1544 2512 1546 2527
rect 1560 2519 1562 2533
rect 1648 2532 1650 2562
rect 1654 2561 1655 2565
rect 1659 2561 1660 2565
rect 1758 2563 1759 2567
rect 1763 2563 1764 2567
rect 1768 2566 1770 2577
rect 1870 2567 1876 2568
rect 1758 2562 1764 2563
rect 1766 2565 1772 2566
rect 1654 2560 1660 2561
rect 1670 2538 1676 2539
rect 1670 2534 1671 2538
rect 1675 2534 1676 2538
rect 1670 2533 1676 2534
rect 1646 2531 1652 2532
rect 1646 2527 1647 2531
rect 1651 2527 1652 2531
rect 1646 2526 1652 2527
rect 1672 2519 1674 2533
rect 1760 2532 1762 2562
rect 1766 2561 1767 2565
rect 1771 2561 1772 2565
rect 1870 2563 1871 2567
rect 1875 2563 1876 2567
rect 1880 2566 1882 2577
rect 1902 2567 1908 2568
rect 1870 2562 1876 2563
rect 1878 2565 1884 2566
rect 1766 2560 1772 2561
rect 1782 2538 1788 2539
rect 1782 2534 1783 2538
rect 1787 2534 1788 2538
rect 1782 2533 1788 2534
rect 1758 2531 1764 2532
rect 1758 2527 1759 2531
rect 1763 2527 1764 2531
rect 1758 2526 1764 2527
rect 1784 2519 1786 2533
rect 1872 2532 1874 2562
rect 1878 2561 1879 2565
rect 1883 2561 1884 2565
rect 1902 2563 1903 2567
rect 1907 2563 1908 2567
rect 1992 2566 1994 2577
rect 2028 2568 2030 2626
rect 2054 2622 2055 2626
rect 2059 2622 2060 2626
rect 2054 2621 2060 2622
rect 2038 2599 2044 2600
rect 2038 2595 2039 2599
rect 2043 2595 2044 2599
rect 2076 2596 2078 2626
rect 2110 2622 2111 2626
rect 2115 2622 2116 2626
rect 2110 2621 2116 2622
rect 2094 2599 2100 2600
rect 2038 2594 2044 2595
rect 2074 2595 2080 2596
rect 2040 2583 2042 2594
rect 2074 2591 2075 2595
rect 2079 2591 2080 2595
rect 2094 2595 2095 2599
rect 2099 2595 2100 2599
rect 2132 2596 2134 2626
rect 2166 2622 2167 2626
rect 2171 2622 2172 2626
rect 2166 2621 2172 2622
rect 2150 2599 2156 2600
rect 2094 2594 2100 2595
rect 2130 2595 2136 2596
rect 2074 2590 2080 2591
rect 2096 2583 2098 2594
rect 2130 2591 2131 2595
rect 2135 2591 2136 2595
rect 2150 2595 2151 2599
rect 2155 2595 2156 2599
rect 2184 2596 2186 2634
rect 2583 2633 2587 2634
rect 2584 2618 2586 2633
rect 2582 2617 2588 2618
rect 2582 2613 2583 2617
rect 2587 2613 2588 2617
rect 2582 2612 2588 2613
rect 2582 2600 2588 2601
rect 2582 2596 2583 2600
rect 2587 2596 2588 2600
rect 2150 2594 2156 2595
rect 2182 2595 2188 2596
rect 2582 2595 2588 2596
rect 2130 2590 2136 2591
rect 2152 2583 2154 2594
rect 2182 2591 2183 2595
rect 2187 2591 2188 2595
rect 2182 2590 2188 2591
rect 2584 2583 2586 2595
rect 2039 2582 2043 2583
rect 2039 2577 2043 2578
rect 2095 2582 2099 2583
rect 2095 2577 2099 2578
rect 2111 2582 2115 2583
rect 2111 2577 2115 2578
rect 2151 2582 2155 2583
rect 2151 2577 2155 2578
rect 2231 2582 2235 2583
rect 2231 2577 2235 2578
rect 2351 2582 2355 2583
rect 2351 2577 2355 2578
rect 2583 2582 2587 2583
rect 2583 2577 2587 2578
rect 2070 2571 2076 2572
rect 2026 2567 2032 2568
rect 1902 2562 1908 2563
rect 1990 2565 1996 2566
rect 1878 2560 1884 2561
rect 1894 2538 1900 2539
rect 1894 2534 1895 2538
rect 1899 2534 1900 2538
rect 1894 2533 1900 2534
rect 1904 2533 1906 2562
rect 1990 2561 1991 2565
rect 1995 2561 1996 2565
rect 2026 2563 2027 2567
rect 2031 2563 2032 2567
rect 2070 2567 2071 2571
rect 2075 2567 2076 2571
rect 2070 2566 2076 2567
rect 2112 2566 2114 2577
rect 2232 2566 2234 2577
rect 2352 2566 2354 2577
rect 2026 2562 2032 2563
rect 1990 2560 1996 2561
rect 2006 2538 2012 2539
rect 2006 2534 2007 2538
rect 2011 2534 2012 2538
rect 2006 2533 2012 2534
rect 1870 2531 1876 2532
rect 1870 2527 1871 2531
rect 1875 2527 1876 2531
rect 1870 2526 1876 2527
rect 1896 2519 1898 2533
rect 1903 2532 1907 2533
rect 1903 2527 1907 2528
rect 2008 2519 2010 2533
rect 2072 2532 2074 2566
rect 2110 2565 2116 2566
rect 2110 2561 2111 2565
rect 2115 2561 2116 2565
rect 2110 2560 2116 2561
rect 2230 2565 2236 2566
rect 2230 2561 2231 2565
rect 2235 2561 2236 2565
rect 2230 2560 2236 2561
rect 2350 2565 2356 2566
rect 2584 2565 2586 2577
rect 2350 2561 2351 2565
rect 2355 2561 2356 2565
rect 2350 2560 2356 2561
rect 2582 2564 2588 2565
rect 2582 2560 2583 2564
rect 2587 2560 2588 2564
rect 2582 2559 2588 2560
rect 2582 2547 2588 2548
rect 2582 2543 2583 2547
rect 2587 2543 2588 2547
rect 2582 2542 2588 2543
rect 2126 2538 2132 2539
rect 2126 2534 2127 2538
rect 2131 2534 2132 2538
rect 2126 2533 2132 2534
rect 2246 2538 2252 2539
rect 2246 2534 2247 2538
rect 2251 2534 2252 2538
rect 2246 2533 2252 2534
rect 2366 2538 2372 2539
rect 2366 2534 2367 2538
rect 2371 2534 2372 2538
rect 2366 2533 2372 2534
rect 2070 2531 2076 2532
rect 2070 2527 2071 2531
rect 2075 2527 2076 2531
rect 2070 2526 2076 2527
rect 2128 2519 2130 2533
rect 2248 2519 2250 2533
rect 2314 2531 2320 2532
rect 2314 2527 2315 2531
rect 2319 2527 2320 2531
rect 2314 2526 2320 2527
rect 1551 2518 1555 2519
rect 1551 2513 1555 2514
rect 1559 2518 1563 2519
rect 1559 2513 1563 2514
rect 1631 2518 1635 2519
rect 1631 2513 1635 2514
rect 1671 2518 1675 2519
rect 1671 2513 1675 2514
rect 1719 2518 1723 2519
rect 1719 2513 1723 2514
rect 1783 2518 1787 2519
rect 1783 2513 1787 2514
rect 1807 2518 1811 2519
rect 1807 2513 1811 2514
rect 1895 2518 1899 2519
rect 1895 2513 1899 2514
rect 1903 2518 1907 2519
rect 1903 2513 1907 2514
rect 1999 2518 2003 2519
rect 1999 2513 2003 2514
rect 2007 2518 2011 2519
rect 2007 2513 2011 2514
rect 2095 2518 2099 2519
rect 2095 2513 2099 2514
rect 2127 2518 2131 2519
rect 2127 2513 2131 2514
rect 2191 2518 2195 2519
rect 2191 2513 2195 2514
rect 2247 2518 2251 2519
rect 2247 2513 2251 2514
rect 2295 2518 2299 2519
rect 2295 2513 2299 2514
rect 1542 2511 1548 2512
rect 1542 2507 1543 2511
rect 1547 2507 1548 2511
rect 1552 2507 1554 2513
rect 1570 2511 1576 2512
rect 1570 2507 1571 2511
rect 1575 2507 1576 2511
rect 1632 2507 1634 2513
rect 1650 2511 1656 2512
rect 1650 2507 1651 2511
rect 1655 2507 1656 2511
rect 1720 2507 1722 2513
rect 1738 2511 1744 2512
rect 1738 2507 1739 2511
rect 1743 2507 1744 2511
rect 1808 2507 1810 2513
rect 1826 2511 1832 2512
rect 1826 2507 1827 2511
rect 1831 2507 1832 2511
rect 1904 2507 1906 2513
rect 1974 2511 1980 2512
rect 1974 2507 1975 2511
rect 1979 2507 1980 2511
rect 2000 2507 2002 2513
rect 2018 2511 2024 2512
rect 2018 2507 2019 2511
rect 2023 2507 2024 2511
rect 2096 2507 2098 2513
rect 2114 2511 2120 2512
rect 2114 2507 2115 2511
rect 2119 2507 2120 2511
rect 2192 2507 2194 2513
rect 2270 2511 2276 2512
rect 2270 2507 2271 2511
rect 2275 2507 2276 2511
rect 2296 2507 2298 2513
rect 1542 2506 1548 2507
rect 1550 2506 1556 2507
rect 1570 2506 1576 2507
rect 1630 2506 1636 2507
rect 1650 2506 1656 2507
rect 1718 2506 1724 2507
rect 1738 2506 1744 2507
rect 1806 2506 1812 2507
rect 1826 2506 1832 2507
rect 1902 2506 1908 2507
rect 1974 2506 1980 2507
rect 1998 2506 2004 2507
rect 2018 2506 2024 2507
rect 2094 2506 2100 2507
rect 2114 2506 2120 2507
rect 2190 2506 2196 2507
rect 2270 2506 2276 2507
rect 2294 2506 2300 2507
rect 1550 2502 1551 2506
rect 1555 2502 1556 2506
rect 1550 2501 1556 2502
rect 1366 2497 1372 2498
rect 1366 2493 1367 2497
rect 1371 2493 1372 2497
rect 1366 2492 1372 2493
rect 1326 2488 1332 2489
rect 1326 2484 1327 2488
rect 1331 2484 1332 2488
rect 998 2482 1004 2483
rect 1022 2483 1028 2484
rect 1326 2483 1332 2484
rect 758 2478 764 2479
rect 792 2467 794 2482
rect 856 2467 858 2482
rect 928 2467 930 2482
rect 1000 2467 1002 2482
rect 1022 2479 1023 2483
rect 1027 2479 1028 2483
rect 1022 2478 1028 2479
rect 1328 2467 1330 2483
rect 1366 2480 1372 2481
rect 1366 2476 1367 2480
rect 1371 2476 1372 2480
rect 1366 2475 1372 2476
rect 1534 2479 1540 2480
rect 1534 2475 1535 2479
rect 1539 2475 1540 2479
rect 1572 2476 1574 2506
rect 1630 2502 1631 2506
rect 1635 2502 1636 2506
rect 1630 2501 1636 2502
rect 1614 2479 1620 2480
rect 631 2466 635 2467
rect 631 2461 635 2462
rect 663 2466 667 2467
rect 663 2461 667 2462
rect 711 2466 715 2467
rect 711 2461 715 2462
rect 727 2466 731 2467
rect 727 2461 731 2462
rect 783 2466 787 2467
rect 783 2461 787 2462
rect 791 2466 795 2467
rect 791 2461 795 2462
rect 855 2466 859 2467
rect 855 2461 859 2462
rect 863 2466 867 2467
rect 863 2461 867 2462
rect 927 2466 931 2467
rect 927 2461 931 2462
rect 943 2466 947 2467
rect 943 2461 947 2462
rect 999 2466 1003 2467
rect 999 2461 1003 2462
rect 1023 2466 1027 2467
rect 1023 2461 1027 2462
rect 1327 2466 1331 2467
rect 1368 2463 1370 2475
rect 1534 2474 1540 2475
rect 1570 2475 1576 2476
rect 1536 2463 1538 2474
rect 1570 2471 1571 2475
rect 1575 2471 1576 2475
rect 1614 2475 1615 2479
rect 1619 2475 1620 2479
rect 1652 2476 1654 2506
rect 1718 2502 1719 2506
rect 1723 2502 1724 2506
rect 1718 2501 1724 2502
rect 1702 2479 1708 2480
rect 1614 2474 1620 2475
rect 1650 2475 1656 2476
rect 1570 2470 1576 2471
rect 1616 2463 1618 2474
rect 1650 2471 1651 2475
rect 1655 2471 1656 2475
rect 1702 2475 1703 2479
rect 1707 2475 1708 2479
rect 1740 2476 1742 2506
rect 1806 2502 1807 2506
rect 1811 2502 1812 2506
rect 1806 2501 1812 2502
rect 1790 2479 1796 2480
rect 1702 2474 1708 2475
rect 1738 2475 1744 2476
rect 1650 2470 1656 2471
rect 1654 2467 1660 2468
rect 1654 2463 1655 2467
rect 1659 2463 1660 2467
rect 1704 2463 1706 2474
rect 1738 2471 1739 2475
rect 1743 2471 1744 2475
rect 1790 2475 1791 2479
rect 1795 2475 1796 2479
rect 1828 2476 1830 2506
rect 1902 2502 1903 2506
rect 1907 2502 1908 2506
rect 1902 2501 1908 2502
rect 1886 2479 1892 2480
rect 1790 2474 1796 2475
rect 1826 2475 1832 2476
rect 1738 2470 1744 2471
rect 1792 2463 1794 2474
rect 1826 2471 1827 2475
rect 1831 2471 1832 2475
rect 1886 2475 1887 2479
rect 1891 2475 1892 2479
rect 1886 2474 1892 2475
rect 1826 2470 1832 2471
rect 1888 2463 1890 2474
rect 1327 2461 1331 2462
rect 1367 2462 1371 2463
rect 632 2450 634 2461
rect 712 2450 714 2461
rect 718 2459 724 2460
rect 718 2455 719 2459
rect 723 2455 724 2459
rect 718 2454 724 2455
rect 630 2449 636 2450
rect 630 2445 631 2449
rect 635 2445 636 2449
rect 630 2444 636 2445
rect 710 2449 716 2450
rect 710 2445 711 2449
rect 715 2445 716 2449
rect 710 2444 716 2445
rect 646 2422 652 2423
rect 646 2418 647 2422
rect 651 2418 652 2422
rect 646 2417 652 2418
rect 622 2415 628 2416
rect 622 2411 623 2415
rect 627 2411 628 2415
rect 622 2410 628 2411
rect 648 2407 650 2417
rect 720 2416 722 2454
rect 774 2451 780 2452
rect 774 2447 775 2451
rect 779 2447 780 2451
rect 784 2450 786 2461
rect 854 2451 860 2452
rect 774 2446 780 2447
rect 782 2449 788 2450
rect 726 2422 732 2423
rect 726 2418 727 2422
rect 731 2418 732 2422
rect 726 2417 732 2418
rect 718 2415 724 2416
rect 718 2411 719 2415
rect 723 2411 724 2415
rect 718 2410 724 2411
rect 728 2407 730 2417
rect 776 2416 778 2446
rect 782 2445 783 2449
rect 787 2445 788 2449
rect 854 2447 855 2451
rect 859 2447 860 2451
rect 864 2450 866 2461
rect 944 2450 946 2461
rect 1014 2451 1020 2452
rect 854 2446 860 2447
rect 862 2449 868 2450
rect 782 2444 788 2445
rect 798 2422 804 2423
rect 798 2418 799 2422
rect 803 2418 804 2422
rect 798 2417 804 2418
rect 774 2415 780 2416
rect 774 2411 775 2415
rect 779 2411 780 2415
rect 774 2410 780 2411
rect 800 2407 802 2417
rect 856 2416 858 2446
rect 862 2445 863 2449
rect 867 2445 868 2449
rect 862 2444 868 2445
rect 942 2449 948 2450
rect 942 2445 943 2449
rect 947 2445 948 2449
rect 1014 2447 1015 2451
rect 1019 2447 1020 2451
rect 1024 2450 1026 2461
rect 1014 2446 1020 2447
rect 1022 2449 1028 2450
rect 1328 2449 1330 2461
rect 1367 2457 1371 2458
rect 1535 2462 1539 2463
rect 1535 2457 1539 2458
rect 1615 2462 1619 2463
rect 1615 2457 1619 2458
rect 1647 2462 1651 2463
rect 1654 2462 1660 2463
rect 1703 2462 1707 2463
rect 1647 2457 1651 2458
rect 942 2444 948 2445
rect 878 2422 884 2423
rect 878 2418 879 2422
rect 883 2418 884 2422
rect 878 2417 884 2418
rect 958 2422 964 2423
rect 958 2418 959 2422
rect 963 2418 964 2422
rect 958 2417 964 2418
rect 854 2415 860 2416
rect 854 2411 855 2415
rect 859 2411 860 2415
rect 854 2410 860 2411
rect 880 2407 882 2417
rect 934 2415 940 2416
rect 934 2411 935 2415
rect 939 2411 940 2415
rect 934 2410 940 2411
rect 431 2406 435 2407
rect 431 2401 435 2402
rect 487 2406 491 2407
rect 487 2401 491 2402
rect 527 2406 531 2407
rect 527 2401 531 2402
rect 567 2406 571 2407
rect 567 2401 571 2402
rect 631 2406 635 2407
rect 631 2401 635 2402
rect 647 2406 651 2407
rect 647 2401 651 2402
rect 727 2406 731 2407
rect 727 2401 731 2402
rect 799 2406 803 2407
rect 799 2401 803 2402
rect 823 2406 827 2407
rect 823 2401 827 2402
rect 879 2406 883 2407
rect 879 2401 883 2402
rect 919 2406 923 2407
rect 919 2401 923 2402
rect 422 2399 428 2400
rect 422 2395 423 2399
rect 427 2395 428 2399
rect 432 2395 434 2401
rect 450 2399 456 2400
rect 450 2395 451 2399
rect 455 2395 456 2399
rect 528 2395 530 2401
rect 546 2399 552 2400
rect 546 2395 547 2399
rect 551 2395 552 2399
rect 632 2395 634 2401
rect 702 2399 708 2400
rect 702 2395 703 2399
rect 707 2395 708 2399
rect 728 2395 730 2401
rect 746 2399 752 2400
rect 746 2395 747 2399
rect 751 2395 752 2399
rect 824 2395 826 2401
rect 842 2399 848 2400
rect 842 2395 843 2399
rect 847 2395 848 2399
rect 920 2395 922 2401
rect 238 2394 244 2395
rect 246 2394 252 2395
rect 266 2394 272 2395
rect 334 2394 340 2395
rect 422 2394 428 2395
rect 430 2394 436 2395
rect 450 2394 456 2395
rect 526 2394 532 2395
rect 546 2394 552 2395
rect 630 2394 636 2395
rect 702 2394 708 2395
rect 726 2394 732 2395
rect 746 2394 752 2395
rect 822 2394 828 2395
rect 842 2394 848 2395
rect 918 2394 924 2395
rect 110 2385 116 2386
rect 110 2381 111 2385
rect 115 2381 116 2385
rect 110 2380 116 2381
rect 240 2373 242 2394
rect 246 2390 247 2394
rect 251 2390 252 2394
rect 246 2389 252 2390
rect 239 2372 243 2373
rect 110 2368 116 2369
rect 110 2364 111 2368
rect 115 2364 116 2368
rect 110 2363 116 2364
rect 230 2367 236 2368
rect 239 2367 243 2368
rect 230 2363 231 2367
rect 235 2363 236 2367
rect 268 2364 270 2394
rect 334 2390 335 2394
rect 339 2390 340 2394
rect 334 2389 340 2390
rect 430 2390 431 2394
rect 435 2390 436 2394
rect 430 2389 436 2390
rect 318 2367 324 2368
rect 112 2351 114 2363
rect 230 2362 236 2363
rect 266 2363 272 2364
rect 232 2351 234 2362
rect 266 2359 267 2363
rect 271 2359 272 2363
rect 318 2363 319 2367
rect 323 2363 324 2367
rect 414 2367 420 2368
rect 318 2362 324 2363
rect 354 2363 360 2364
rect 266 2358 272 2359
rect 320 2351 322 2362
rect 354 2359 355 2363
rect 359 2359 360 2363
rect 414 2363 415 2367
rect 419 2363 420 2367
rect 452 2364 454 2394
rect 526 2390 527 2394
rect 531 2390 532 2394
rect 526 2389 532 2390
rect 510 2367 516 2368
rect 414 2362 420 2363
rect 450 2363 456 2364
rect 354 2358 360 2359
rect 111 2350 115 2351
rect 111 2345 115 2346
rect 159 2350 163 2351
rect 159 2345 163 2346
rect 231 2350 235 2351
rect 231 2345 235 2346
rect 263 2350 267 2351
rect 263 2345 267 2346
rect 319 2350 323 2351
rect 319 2345 323 2346
rect 112 2333 114 2345
rect 160 2334 162 2345
rect 166 2343 172 2344
rect 166 2339 167 2343
rect 171 2339 172 2343
rect 166 2338 172 2339
rect 158 2333 164 2334
rect 110 2332 116 2333
rect 110 2328 111 2332
rect 115 2328 116 2332
rect 158 2329 159 2333
rect 163 2329 164 2333
rect 158 2328 164 2329
rect 110 2327 116 2328
rect 110 2315 116 2316
rect 110 2311 111 2315
rect 115 2311 116 2315
rect 110 2310 116 2311
rect 112 2291 114 2310
rect 168 2300 170 2338
rect 254 2335 260 2336
rect 254 2331 255 2335
rect 259 2331 260 2335
rect 264 2334 266 2345
rect 346 2335 352 2336
rect 254 2330 260 2331
rect 262 2333 268 2334
rect 174 2306 180 2307
rect 174 2302 175 2306
rect 179 2302 180 2306
rect 174 2301 180 2302
rect 166 2299 172 2300
rect 166 2295 167 2299
rect 171 2295 172 2299
rect 166 2294 172 2295
rect 176 2291 178 2301
rect 256 2300 258 2330
rect 262 2329 263 2333
rect 267 2329 268 2333
rect 346 2331 347 2335
rect 351 2331 352 2335
rect 346 2330 352 2331
rect 262 2328 268 2329
rect 278 2306 284 2307
rect 278 2302 279 2306
rect 283 2302 284 2306
rect 278 2301 284 2302
rect 254 2299 260 2300
rect 254 2295 255 2299
rect 259 2295 260 2299
rect 254 2294 260 2295
rect 280 2291 282 2301
rect 111 2290 115 2291
rect 111 2285 115 2286
rect 159 2290 163 2291
rect 159 2285 163 2286
rect 175 2290 179 2291
rect 175 2285 179 2286
rect 247 2290 251 2291
rect 247 2285 251 2286
rect 279 2290 283 2291
rect 279 2285 283 2286
rect 112 2270 114 2285
rect 134 2283 140 2284
rect 134 2279 135 2283
rect 139 2279 140 2283
rect 160 2279 162 2285
rect 248 2279 250 2285
rect 348 2284 350 2330
rect 356 2300 358 2358
rect 416 2351 418 2362
rect 450 2359 451 2363
rect 455 2359 456 2363
rect 510 2363 511 2367
rect 515 2363 516 2367
rect 548 2364 550 2394
rect 630 2390 631 2394
rect 635 2390 636 2394
rect 630 2389 636 2390
rect 704 2376 706 2394
rect 726 2390 727 2394
rect 731 2390 732 2394
rect 726 2389 732 2390
rect 702 2375 708 2376
rect 647 2372 651 2373
rect 702 2371 703 2375
rect 707 2371 708 2375
rect 702 2370 708 2371
rect 614 2367 620 2368
rect 647 2367 651 2368
rect 710 2367 716 2368
rect 510 2362 516 2363
rect 546 2363 552 2364
rect 450 2358 456 2359
rect 512 2351 514 2362
rect 546 2359 547 2363
rect 551 2359 552 2363
rect 614 2363 615 2367
rect 619 2363 620 2367
rect 648 2364 650 2367
rect 614 2362 620 2363
rect 646 2363 652 2364
rect 546 2358 552 2359
rect 616 2351 618 2362
rect 646 2359 647 2363
rect 651 2359 652 2363
rect 710 2363 711 2367
rect 715 2363 716 2367
rect 748 2364 750 2394
rect 822 2390 823 2394
rect 827 2390 828 2394
rect 822 2389 828 2390
rect 806 2367 812 2368
rect 710 2362 716 2363
rect 746 2363 752 2364
rect 646 2358 652 2359
rect 712 2351 714 2362
rect 746 2359 747 2363
rect 751 2359 752 2363
rect 806 2363 807 2367
rect 811 2363 812 2367
rect 844 2364 846 2394
rect 918 2390 919 2394
rect 923 2390 924 2394
rect 918 2389 924 2390
rect 902 2367 908 2368
rect 806 2362 812 2363
rect 842 2363 848 2364
rect 746 2358 752 2359
rect 808 2351 810 2362
rect 842 2359 843 2363
rect 847 2359 848 2363
rect 902 2363 903 2367
rect 907 2363 908 2367
rect 936 2364 938 2410
rect 960 2407 962 2417
rect 1016 2416 1018 2446
rect 1022 2445 1023 2449
rect 1027 2445 1028 2449
rect 1022 2444 1028 2445
rect 1326 2448 1332 2449
rect 1326 2444 1327 2448
rect 1331 2444 1332 2448
rect 1368 2445 1370 2457
rect 1648 2446 1650 2457
rect 1646 2445 1652 2446
rect 1326 2443 1332 2444
rect 1366 2444 1372 2445
rect 1366 2440 1367 2444
rect 1371 2440 1372 2444
rect 1646 2441 1647 2445
rect 1651 2441 1652 2445
rect 1646 2440 1652 2441
rect 1366 2439 1372 2440
rect 1326 2431 1332 2432
rect 1326 2427 1327 2431
rect 1331 2427 1332 2431
rect 1326 2426 1332 2427
rect 1366 2427 1372 2428
rect 1038 2422 1044 2423
rect 1038 2418 1039 2422
rect 1043 2418 1044 2422
rect 1038 2417 1044 2418
rect 1014 2415 1020 2416
rect 1014 2411 1015 2415
rect 1019 2411 1020 2415
rect 1014 2410 1020 2411
rect 1040 2407 1042 2417
rect 1328 2407 1330 2426
rect 1366 2423 1367 2427
rect 1371 2423 1372 2427
rect 1366 2422 1372 2423
rect 959 2406 963 2407
rect 959 2401 963 2402
rect 1015 2406 1019 2407
rect 1015 2401 1019 2402
rect 1039 2406 1043 2407
rect 1039 2401 1043 2402
rect 1111 2406 1115 2407
rect 1111 2401 1115 2402
rect 1327 2406 1331 2407
rect 1368 2403 1370 2422
rect 1656 2412 1658 2462
rect 1703 2457 1707 2458
rect 1767 2462 1771 2463
rect 1767 2457 1771 2458
rect 1791 2462 1795 2463
rect 1791 2457 1795 2458
rect 1839 2462 1843 2463
rect 1839 2457 1843 2458
rect 1887 2462 1891 2463
rect 1887 2457 1891 2458
rect 1911 2462 1915 2463
rect 1911 2457 1915 2458
rect 1694 2447 1700 2448
rect 1694 2443 1695 2447
rect 1699 2443 1700 2447
rect 1704 2446 1706 2457
rect 1758 2447 1764 2448
rect 1694 2442 1700 2443
rect 1702 2445 1708 2446
rect 1662 2418 1668 2419
rect 1662 2414 1663 2418
rect 1667 2414 1668 2418
rect 1662 2413 1668 2414
rect 1654 2411 1660 2412
rect 1654 2407 1655 2411
rect 1659 2407 1660 2411
rect 1654 2406 1660 2407
rect 1664 2403 1666 2413
rect 1696 2412 1698 2442
rect 1702 2441 1703 2445
rect 1707 2441 1708 2445
rect 1758 2443 1759 2447
rect 1763 2443 1764 2447
rect 1768 2446 1770 2457
rect 1830 2447 1836 2448
rect 1758 2442 1764 2443
rect 1766 2445 1772 2446
rect 1702 2440 1708 2441
rect 1718 2418 1724 2419
rect 1718 2414 1719 2418
rect 1723 2414 1724 2418
rect 1718 2413 1724 2414
rect 1694 2411 1700 2412
rect 1694 2407 1695 2411
rect 1699 2407 1700 2411
rect 1694 2406 1700 2407
rect 1720 2403 1722 2413
rect 1760 2412 1762 2442
rect 1766 2441 1767 2445
rect 1771 2441 1772 2445
rect 1830 2443 1831 2447
rect 1835 2443 1836 2447
rect 1840 2446 1842 2457
rect 1902 2447 1908 2448
rect 1830 2442 1836 2443
rect 1838 2445 1844 2446
rect 1766 2440 1772 2441
rect 1782 2418 1788 2419
rect 1782 2414 1783 2418
rect 1787 2414 1788 2418
rect 1782 2413 1788 2414
rect 1758 2411 1764 2412
rect 1758 2407 1759 2411
rect 1763 2407 1764 2411
rect 1758 2406 1764 2407
rect 1784 2403 1786 2413
rect 1832 2412 1834 2442
rect 1838 2441 1839 2445
rect 1843 2441 1844 2445
rect 1902 2443 1903 2447
rect 1907 2443 1908 2447
rect 1912 2446 1914 2457
rect 1976 2456 1978 2506
rect 1998 2502 1999 2506
rect 2003 2502 2004 2506
rect 1998 2501 2004 2502
rect 1982 2479 1988 2480
rect 1982 2475 1983 2479
rect 1987 2475 1988 2479
rect 2020 2476 2022 2506
rect 2094 2502 2095 2506
rect 2099 2502 2100 2506
rect 2094 2501 2100 2502
rect 2078 2479 2084 2480
rect 1982 2474 1988 2475
rect 2018 2475 2024 2476
rect 1984 2463 1986 2474
rect 2018 2471 2019 2475
rect 2023 2471 2024 2475
rect 2078 2475 2079 2479
rect 2083 2475 2084 2479
rect 2116 2476 2118 2506
rect 2190 2502 2191 2506
rect 2195 2502 2196 2506
rect 2190 2501 2196 2502
rect 2272 2488 2274 2506
rect 2294 2502 2295 2506
rect 2299 2502 2300 2506
rect 2294 2501 2300 2502
rect 2270 2487 2276 2488
rect 2270 2483 2271 2487
rect 2275 2483 2276 2487
rect 2270 2482 2276 2483
rect 2174 2479 2180 2480
rect 2078 2474 2084 2475
rect 2114 2475 2120 2476
rect 2018 2470 2024 2471
rect 2080 2463 2082 2474
rect 2114 2471 2115 2475
rect 2119 2471 2120 2475
rect 2174 2475 2175 2479
rect 2179 2475 2180 2479
rect 2278 2479 2284 2480
rect 2174 2474 2180 2475
rect 2254 2475 2260 2476
rect 2114 2470 2120 2471
rect 2176 2463 2178 2474
rect 2254 2471 2255 2475
rect 2259 2471 2260 2475
rect 2278 2475 2279 2479
rect 2283 2475 2284 2479
rect 2316 2476 2318 2526
rect 2368 2519 2370 2533
rect 2584 2519 2586 2542
rect 2367 2518 2371 2519
rect 2367 2513 2371 2514
rect 2399 2518 2403 2519
rect 2399 2513 2403 2514
rect 2583 2518 2587 2519
rect 2583 2513 2587 2514
rect 2390 2511 2396 2512
rect 2390 2507 2391 2511
rect 2395 2507 2396 2511
rect 2400 2507 2402 2513
rect 2390 2506 2396 2507
rect 2398 2506 2404 2507
rect 2382 2479 2388 2480
rect 2278 2474 2284 2475
rect 2314 2475 2320 2476
rect 2254 2470 2260 2471
rect 1983 2462 1987 2463
rect 1983 2457 1987 2458
rect 1991 2462 1995 2463
rect 1991 2457 1995 2458
rect 2079 2462 2083 2463
rect 2079 2457 2083 2458
rect 2167 2462 2171 2463
rect 2167 2457 2171 2458
rect 2175 2462 2179 2463
rect 2175 2457 2179 2458
rect 1974 2455 1980 2456
rect 1974 2451 1975 2455
rect 1979 2451 1980 2455
rect 1974 2450 1980 2451
rect 1934 2447 1940 2448
rect 1902 2442 1908 2443
rect 1910 2445 1916 2446
rect 1838 2440 1844 2441
rect 1854 2418 1860 2419
rect 1854 2414 1855 2418
rect 1859 2414 1860 2418
rect 1854 2413 1860 2414
rect 1830 2411 1836 2412
rect 1830 2407 1831 2411
rect 1835 2407 1836 2411
rect 1830 2406 1836 2407
rect 1856 2403 1858 2413
rect 1904 2412 1906 2442
rect 1910 2441 1911 2445
rect 1915 2441 1916 2445
rect 1934 2443 1935 2447
rect 1939 2443 1940 2447
rect 1992 2446 1994 2457
rect 2070 2447 2076 2448
rect 1934 2442 1940 2443
rect 1990 2445 1996 2446
rect 1910 2440 1916 2441
rect 1926 2418 1932 2419
rect 1926 2414 1927 2418
rect 1931 2414 1932 2418
rect 1926 2413 1932 2414
rect 1902 2411 1908 2412
rect 1902 2407 1903 2411
rect 1907 2407 1908 2411
rect 1902 2406 1908 2407
rect 1928 2403 1930 2413
rect 1936 2408 1938 2442
rect 1990 2441 1991 2445
rect 1995 2441 1996 2445
rect 2070 2443 2071 2447
rect 2075 2443 2076 2447
rect 2080 2446 2082 2457
rect 2158 2447 2164 2448
rect 2070 2442 2076 2443
rect 2078 2445 2084 2446
rect 1990 2440 1996 2441
rect 2006 2418 2012 2419
rect 2006 2414 2007 2418
rect 2011 2414 2012 2418
rect 2006 2413 2012 2414
rect 1962 2411 1968 2412
rect 1934 2407 1940 2408
rect 1934 2403 1935 2407
rect 1939 2403 1940 2407
rect 1962 2407 1963 2411
rect 1967 2407 1968 2411
rect 1962 2406 1968 2407
rect 1327 2401 1331 2402
rect 1367 2402 1371 2403
rect 1016 2395 1018 2401
rect 1112 2395 1114 2401
rect 1014 2394 1020 2395
rect 1014 2390 1015 2394
rect 1019 2390 1020 2394
rect 1014 2389 1020 2390
rect 1110 2394 1116 2395
rect 1110 2390 1111 2394
rect 1115 2390 1116 2394
rect 1110 2389 1116 2390
rect 1328 2386 1330 2401
rect 1367 2397 1371 2398
rect 1455 2402 1459 2403
rect 1455 2397 1459 2398
rect 1559 2402 1563 2403
rect 1559 2397 1563 2398
rect 1663 2402 1667 2403
rect 1663 2397 1667 2398
rect 1719 2402 1723 2403
rect 1719 2397 1723 2398
rect 1759 2402 1763 2403
rect 1759 2397 1763 2398
rect 1783 2402 1787 2403
rect 1783 2397 1787 2398
rect 1855 2402 1859 2403
rect 1855 2397 1859 2398
rect 1927 2402 1931 2403
rect 1934 2402 1940 2403
rect 1943 2402 1947 2403
rect 1927 2397 1931 2398
rect 1943 2397 1947 2398
rect 1326 2385 1332 2386
rect 1326 2381 1327 2385
rect 1331 2381 1332 2385
rect 1368 2382 1370 2397
rect 1446 2395 1452 2396
rect 1446 2391 1447 2395
rect 1451 2391 1452 2395
rect 1456 2391 1458 2397
rect 1560 2391 1562 2397
rect 1578 2395 1584 2396
rect 1578 2391 1579 2395
rect 1583 2391 1584 2395
rect 1664 2391 1666 2397
rect 1682 2395 1688 2396
rect 1682 2391 1683 2395
rect 1687 2391 1688 2395
rect 1760 2391 1762 2397
rect 1856 2391 1858 2397
rect 1944 2391 1946 2397
rect 1446 2390 1452 2391
rect 1454 2390 1460 2391
rect 1326 2380 1332 2381
rect 1366 2381 1372 2382
rect 1366 2377 1367 2381
rect 1371 2377 1372 2381
rect 1366 2376 1372 2377
rect 1326 2368 1332 2369
rect 998 2367 1004 2368
rect 902 2362 908 2363
rect 934 2363 940 2364
rect 842 2358 848 2359
rect 904 2351 906 2362
rect 934 2359 935 2363
rect 939 2359 940 2363
rect 998 2363 999 2367
rect 1003 2363 1004 2367
rect 998 2362 1004 2363
rect 1094 2367 1100 2368
rect 1094 2363 1095 2367
rect 1099 2363 1100 2367
rect 1326 2364 1327 2368
rect 1331 2364 1332 2368
rect 1326 2363 1332 2364
rect 1366 2364 1372 2365
rect 1094 2362 1100 2363
rect 934 2358 940 2359
rect 1000 2351 1002 2362
rect 1096 2351 1098 2362
rect 1328 2351 1330 2363
rect 1366 2360 1367 2364
rect 1371 2360 1372 2364
rect 1366 2359 1372 2360
rect 1438 2363 1444 2364
rect 1438 2359 1439 2363
rect 1443 2359 1444 2363
rect 375 2350 379 2351
rect 375 2345 379 2346
rect 415 2350 419 2351
rect 415 2345 419 2346
rect 487 2350 491 2351
rect 487 2345 491 2346
rect 511 2350 515 2351
rect 511 2345 515 2346
rect 599 2350 603 2351
rect 599 2345 603 2346
rect 615 2350 619 2351
rect 615 2345 619 2346
rect 711 2350 715 2351
rect 711 2345 715 2346
rect 807 2350 811 2351
rect 807 2345 811 2346
rect 815 2350 819 2351
rect 815 2345 819 2346
rect 903 2350 907 2351
rect 903 2345 907 2346
rect 911 2350 915 2351
rect 911 2345 915 2346
rect 999 2350 1003 2351
rect 999 2345 1003 2346
rect 1007 2350 1011 2351
rect 1007 2345 1011 2346
rect 1095 2350 1099 2351
rect 1095 2345 1099 2346
rect 1103 2350 1107 2351
rect 1103 2345 1107 2346
rect 1199 2350 1203 2351
rect 1199 2345 1203 2346
rect 1327 2350 1331 2351
rect 1368 2347 1370 2359
rect 1438 2358 1444 2359
rect 1440 2347 1442 2358
rect 1327 2345 1331 2346
rect 1367 2346 1371 2347
rect 376 2334 378 2345
rect 478 2335 484 2336
rect 374 2333 380 2334
rect 374 2329 375 2333
rect 379 2329 380 2333
rect 478 2331 479 2335
rect 483 2331 484 2335
rect 488 2334 490 2345
rect 590 2335 596 2336
rect 478 2330 484 2331
rect 486 2333 492 2334
rect 374 2328 380 2329
rect 390 2306 396 2307
rect 390 2302 391 2306
rect 395 2302 396 2306
rect 390 2301 396 2302
rect 354 2299 360 2300
rect 354 2295 355 2299
rect 359 2295 360 2299
rect 354 2294 360 2295
rect 392 2291 394 2301
rect 480 2300 482 2330
rect 486 2329 487 2333
rect 491 2329 492 2333
rect 590 2331 591 2335
rect 595 2331 596 2335
rect 600 2334 602 2345
rect 712 2334 714 2345
rect 734 2343 740 2344
rect 734 2339 735 2343
rect 739 2339 740 2343
rect 734 2338 740 2339
rect 590 2330 596 2331
rect 598 2333 604 2334
rect 486 2328 492 2329
rect 502 2306 508 2307
rect 502 2302 503 2306
rect 507 2302 508 2306
rect 502 2301 508 2302
rect 478 2299 484 2300
rect 478 2295 479 2299
rect 483 2295 484 2299
rect 478 2294 484 2295
rect 504 2291 506 2301
rect 592 2300 594 2330
rect 598 2329 599 2333
rect 603 2329 604 2333
rect 598 2328 604 2329
rect 710 2333 716 2334
rect 710 2329 711 2333
rect 715 2329 716 2333
rect 710 2328 716 2329
rect 614 2306 620 2307
rect 614 2302 615 2306
rect 619 2302 620 2306
rect 614 2301 620 2302
rect 726 2306 732 2307
rect 726 2302 727 2306
rect 731 2302 732 2306
rect 726 2301 732 2302
rect 590 2299 596 2300
rect 590 2295 591 2299
rect 595 2295 596 2299
rect 590 2294 596 2295
rect 616 2291 618 2301
rect 646 2291 652 2292
rect 728 2291 730 2301
rect 736 2300 738 2338
rect 806 2335 812 2336
rect 806 2331 807 2335
rect 811 2331 812 2335
rect 816 2334 818 2345
rect 902 2335 908 2336
rect 806 2330 812 2331
rect 814 2333 820 2334
rect 808 2300 810 2330
rect 814 2329 815 2333
rect 819 2329 820 2333
rect 902 2331 903 2335
rect 907 2331 908 2335
rect 912 2334 914 2345
rect 1008 2334 1010 2345
rect 1094 2335 1100 2336
rect 902 2330 908 2331
rect 910 2333 916 2334
rect 814 2328 820 2329
rect 830 2306 836 2307
rect 830 2302 831 2306
rect 835 2302 836 2306
rect 830 2301 836 2302
rect 734 2299 740 2300
rect 734 2295 735 2299
rect 739 2295 740 2299
rect 734 2294 740 2295
rect 806 2299 812 2300
rect 806 2295 807 2299
rect 811 2295 812 2299
rect 806 2294 812 2295
rect 832 2291 834 2301
rect 904 2300 906 2330
rect 910 2329 911 2333
rect 915 2329 916 2333
rect 910 2328 916 2329
rect 1006 2333 1012 2334
rect 1006 2329 1007 2333
rect 1011 2329 1012 2333
rect 1094 2331 1095 2335
rect 1099 2331 1100 2335
rect 1104 2334 1106 2345
rect 1190 2335 1196 2336
rect 1094 2330 1100 2331
rect 1102 2333 1108 2334
rect 1006 2328 1012 2329
rect 926 2306 932 2307
rect 926 2302 927 2306
rect 931 2302 932 2306
rect 926 2301 932 2302
rect 1022 2306 1028 2307
rect 1022 2302 1023 2306
rect 1027 2302 1028 2306
rect 1022 2301 1028 2302
rect 902 2299 908 2300
rect 902 2295 903 2299
rect 907 2295 908 2299
rect 902 2294 908 2295
rect 928 2291 930 2301
rect 1014 2299 1020 2300
rect 1014 2295 1015 2299
rect 1019 2295 1020 2299
rect 1014 2294 1020 2295
rect 375 2290 379 2291
rect 375 2285 379 2286
rect 391 2290 395 2291
rect 391 2285 395 2286
rect 503 2290 507 2291
rect 503 2285 507 2286
rect 511 2290 515 2291
rect 511 2285 515 2286
rect 615 2290 619 2291
rect 615 2285 619 2286
rect 639 2290 643 2291
rect 646 2287 647 2291
rect 651 2287 652 2291
rect 646 2286 652 2287
rect 727 2290 731 2291
rect 639 2285 643 2286
rect 346 2283 352 2284
rect 346 2279 347 2283
rect 351 2279 352 2283
rect 376 2279 378 2285
rect 442 2283 448 2284
rect 442 2279 443 2283
rect 447 2279 448 2283
rect 512 2279 514 2285
rect 530 2283 536 2284
rect 530 2279 531 2283
rect 535 2279 536 2283
rect 640 2279 642 2285
rect 134 2278 140 2279
rect 158 2278 164 2279
rect 110 2269 116 2270
rect 110 2265 111 2269
rect 115 2265 116 2269
rect 110 2264 116 2265
rect 136 2260 138 2278
rect 158 2274 159 2278
rect 163 2274 164 2278
rect 158 2273 164 2274
rect 246 2278 252 2279
rect 346 2278 352 2279
rect 374 2278 380 2279
rect 442 2278 448 2279
rect 510 2278 516 2279
rect 530 2278 536 2279
rect 638 2278 644 2279
rect 246 2274 247 2278
rect 251 2274 252 2278
rect 246 2273 252 2274
rect 374 2274 375 2278
rect 379 2274 380 2278
rect 374 2273 380 2274
rect 134 2259 140 2260
rect 134 2255 135 2259
rect 139 2255 140 2259
rect 134 2254 140 2255
rect 110 2252 116 2253
rect 444 2252 446 2278
rect 510 2274 511 2278
rect 515 2274 516 2278
rect 510 2273 516 2274
rect 110 2248 111 2252
rect 115 2248 116 2252
rect 110 2247 116 2248
rect 142 2251 148 2252
rect 142 2247 143 2251
rect 147 2247 148 2251
rect 230 2251 236 2252
rect 112 2227 114 2247
rect 142 2246 148 2247
rect 166 2247 172 2248
rect 144 2227 146 2246
rect 166 2243 167 2247
rect 171 2243 172 2247
rect 230 2247 231 2251
rect 235 2247 236 2251
rect 230 2246 236 2247
rect 358 2251 364 2252
rect 358 2247 359 2251
rect 363 2247 364 2251
rect 358 2246 364 2247
rect 442 2251 448 2252
rect 442 2247 443 2251
rect 447 2247 448 2251
rect 442 2246 448 2247
rect 494 2251 500 2252
rect 494 2247 495 2251
rect 499 2247 500 2251
rect 532 2248 534 2278
rect 638 2274 639 2278
rect 643 2274 644 2278
rect 638 2273 644 2274
rect 622 2251 628 2252
rect 494 2246 500 2247
rect 530 2247 536 2248
rect 166 2242 172 2243
rect 111 2226 115 2227
rect 111 2221 115 2222
rect 143 2226 147 2227
rect 143 2221 147 2222
rect 112 2209 114 2221
rect 144 2210 146 2221
rect 142 2209 148 2210
rect 110 2208 116 2209
rect 110 2204 111 2208
rect 115 2204 116 2208
rect 142 2205 143 2209
rect 147 2205 148 2209
rect 142 2204 148 2205
rect 110 2203 116 2204
rect 110 2191 116 2192
rect 110 2187 111 2191
rect 115 2187 116 2191
rect 110 2186 116 2187
rect 139 2188 143 2189
rect 112 2167 114 2186
rect 139 2183 143 2184
rect 111 2166 115 2167
rect 111 2161 115 2162
rect 112 2146 114 2161
rect 140 2160 142 2183
rect 158 2182 164 2183
rect 158 2178 159 2182
rect 163 2178 164 2182
rect 158 2177 164 2178
rect 160 2167 162 2177
rect 168 2176 170 2242
rect 232 2227 234 2246
rect 360 2227 362 2246
rect 496 2227 498 2246
rect 530 2243 531 2247
rect 535 2243 536 2247
rect 622 2247 623 2251
rect 627 2247 628 2251
rect 648 2248 650 2286
rect 727 2285 731 2286
rect 767 2290 771 2291
rect 767 2285 771 2286
rect 831 2290 835 2291
rect 831 2285 835 2286
rect 887 2290 891 2291
rect 887 2285 891 2286
rect 927 2290 931 2291
rect 927 2285 931 2286
rect 999 2290 1003 2291
rect 999 2285 1003 2286
rect 768 2279 770 2285
rect 822 2283 828 2284
rect 822 2279 823 2283
rect 827 2279 828 2283
rect 888 2279 890 2285
rect 906 2283 912 2284
rect 906 2279 907 2283
rect 911 2279 912 2283
rect 1000 2279 1002 2285
rect 766 2278 772 2279
rect 822 2278 828 2279
rect 886 2278 892 2279
rect 906 2278 912 2279
rect 998 2278 1004 2279
rect 766 2274 767 2278
rect 771 2274 772 2278
rect 766 2273 772 2274
rect 750 2251 756 2252
rect 622 2246 628 2247
rect 646 2247 652 2248
rect 530 2242 536 2243
rect 624 2227 626 2246
rect 646 2243 647 2247
rect 651 2243 652 2247
rect 750 2247 751 2251
rect 755 2247 756 2251
rect 824 2248 826 2278
rect 886 2274 887 2278
rect 891 2274 892 2278
rect 886 2273 892 2274
rect 870 2251 876 2252
rect 750 2246 756 2247
rect 822 2247 828 2248
rect 646 2242 652 2243
rect 752 2227 754 2246
rect 822 2243 823 2247
rect 827 2243 828 2247
rect 870 2247 871 2251
rect 875 2247 876 2251
rect 908 2248 910 2278
rect 998 2274 999 2278
rect 1003 2274 1004 2278
rect 998 2273 1004 2274
rect 982 2251 988 2252
rect 870 2246 876 2247
rect 906 2247 912 2248
rect 822 2242 828 2243
rect 872 2227 874 2246
rect 906 2243 907 2247
rect 911 2243 912 2247
rect 982 2247 983 2251
rect 987 2247 988 2251
rect 1016 2248 1018 2294
rect 1024 2291 1026 2301
rect 1096 2300 1098 2330
rect 1102 2329 1103 2333
rect 1107 2329 1108 2333
rect 1190 2331 1191 2335
rect 1195 2331 1196 2335
rect 1200 2334 1202 2345
rect 1190 2330 1196 2331
rect 1198 2333 1204 2334
rect 1328 2333 1330 2345
rect 1367 2341 1371 2342
rect 1399 2346 1403 2347
rect 1399 2341 1403 2342
rect 1439 2346 1443 2347
rect 1439 2341 1443 2342
rect 1102 2328 1108 2329
rect 1118 2306 1124 2307
rect 1118 2302 1119 2306
rect 1123 2302 1124 2306
rect 1118 2301 1124 2302
rect 1094 2299 1100 2300
rect 1094 2295 1095 2299
rect 1099 2295 1100 2299
rect 1094 2294 1100 2295
rect 1110 2291 1116 2292
rect 1120 2291 1122 2301
rect 1192 2300 1194 2330
rect 1198 2329 1199 2333
rect 1203 2329 1204 2333
rect 1198 2328 1204 2329
rect 1326 2332 1332 2333
rect 1326 2328 1327 2332
rect 1331 2328 1332 2332
rect 1368 2329 1370 2341
rect 1400 2330 1402 2341
rect 1448 2340 1450 2390
rect 1454 2386 1455 2390
rect 1459 2386 1460 2390
rect 1454 2385 1460 2386
rect 1558 2390 1564 2391
rect 1578 2390 1584 2391
rect 1662 2390 1668 2391
rect 1682 2390 1688 2391
rect 1758 2390 1764 2391
rect 1558 2386 1559 2390
rect 1563 2386 1564 2390
rect 1558 2385 1564 2386
rect 1542 2363 1548 2364
rect 1534 2359 1540 2360
rect 1534 2355 1535 2359
rect 1539 2355 1540 2359
rect 1542 2359 1543 2363
rect 1547 2359 1548 2363
rect 1580 2360 1582 2390
rect 1662 2386 1663 2390
rect 1667 2386 1668 2390
rect 1662 2385 1668 2386
rect 1646 2363 1652 2364
rect 1542 2358 1548 2359
rect 1578 2359 1584 2360
rect 1534 2354 1540 2355
rect 1455 2346 1459 2347
rect 1455 2341 1459 2342
rect 1511 2346 1515 2347
rect 1511 2341 1515 2342
rect 1446 2339 1452 2340
rect 1446 2335 1447 2339
rect 1451 2335 1452 2339
rect 1446 2334 1452 2335
rect 1446 2331 1452 2332
rect 1398 2329 1404 2330
rect 1326 2327 1332 2328
rect 1366 2328 1372 2329
rect 1366 2324 1367 2328
rect 1371 2324 1372 2328
rect 1398 2325 1399 2329
rect 1403 2325 1404 2329
rect 1446 2327 1447 2331
rect 1451 2327 1452 2331
rect 1456 2330 1458 2341
rect 1502 2331 1508 2332
rect 1446 2326 1452 2327
rect 1454 2329 1460 2330
rect 1398 2324 1404 2325
rect 1366 2323 1372 2324
rect 1326 2315 1332 2316
rect 1326 2311 1327 2315
rect 1331 2311 1332 2315
rect 1326 2310 1332 2311
rect 1366 2311 1372 2312
rect 1214 2306 1220 2307
rect 1214 2302 1215 2306
rect 1219 2302 1220 2306
rect 1214 2301 1220 2302
rect 1190 2299 1196 2300
rect 1190 2295 1191 2299
rect 1195 2295 1196 2299
rect 1190 2294 1196 2295
rect 1216 2291 1218 2301
rect 1306 2295 1312 2296
rect 1306 2291 1307 2295
rect 1311 2291 1312 2295
rect 1328 2291 1330 2310
rect 1366 2307 1367 2311
rect 1371 2307 1372 2311
rect 1366 2306 1372 2307
rect 1023 2290 1027 2291
rect 1023 2285 1027 2286
rect 1103 2290 1107 2291
rect 1110 2287 1111 2291
rect 1115 2287 1116 2291
rect 1110 2286 1116 2287
rect 1119 2290 1123 2291
rect 1103 2285 1107 2286
rect 1078 2283 1084 2284
rect 1078 2279 1079 2283
rect 1083 2279 1084 2283
rect 1104 2279 1106 2285
rect 1078 2278 1084 2279
rect 1102 2278 1108 2279
rect 1080 2260 1082 2278
rect 1102 2274 1103 2278
rect 1107 2274 1108 2278
rect 1102 2273 1108 2274
rect 1078 2259 1084 2260
rect 1078 2255 1079 2259
rect 1083 2255 1084 2259
rect 1078 2254 1084 2255
rect 1086 2251 1092 2252
rect 982 2246 988 2247
rect 1014 2247 1020 2248
rect 906 2242 912 2243
rect 984 2227 986 2246
rect 1014 2243 1015 2247
rect 1019 2243 1020 2247
rect 1086 2247 1087 2251
rect 1091 2247 1092 2251
rect 1112 2248 1114 2286
rect 1119 2285 1123 2286
rect 1207 2290 1211 2291
rect 1207 2285 1211 2286
rect 1215 2290 1219 2291
rect 1215 2285 1219 2286
rect 1287 2290 1291 2291
rect 1306 2290 1312 2291
rect 1327 2290 1331 2291
rect 1287 2285 1291 2286
rect 1198 2283 1204 2284
rect 1198 2279 1199 2283
rect 1203 2279 1204 2283
rect 1208 2279 1210 2285
rect 1278 2283 1284 2284
rect 1278 2279 1279 2283
rect 1283 2279 1284 2283
rect 1288 2279 1290 2285
rect 1198 2278 1204 2279
rect 1206 2278 1212 2279
rect 1278 2278 1284 2279
rect 1286 2278 1292 2279
rect 1190 2251 1196 2252
rect 1086 2246 1092 2247
rect 1110 2247 1116 2248
rect 1014 2242 1020 2243
rect 1088 2227 1090 2246
rect 1110 2243 1111 2247
rect 1115 2243 1116 2247
rect 1190 2247 1191 2251
rect 1195 2247 1196 2251
rect 1190 2246 1196 2247
rect 1110 2242 1116 2243
rect 1192 2227 1194 2246
rect 231 2226 235 2227
rect 231 2221 235 2222
rect 359 2226 363 2227
rect 359 2221 363 2222
rect 495 2226 499 2227
rect 495 2221 499 2222
rect 623 2226 627 2227
rect 623 2221 627 2222
rect 751 2226 755 2227
rect 751 2221 755 2222
rect 871 2226 875 2227
rect 871 2221 875 2222
rect 983 2226 987 2227
rect 983 2221 987 2222
rect 1087 2226 1091 2227
rect 1087 2221 1091 2222
rect 1191 2226 1195 2227
rect 1191 2221 1195 2222
rect 222 2211 228 2212
rect 222 2207 223 2211
rect 227 2207 228 2211
rect 232 2210 234 2221
rect 350 2211 356 2212
rect 222 2206 228 2207
rect 230 2209 236 2210
rect 224 2176 226 2206
rect 230 2205 231 2209
rect 235 2205 236 2209
rect 350 2207 351 2211
rect 355 2207 356 2211
rect 360 2210 362 2221
rect 486 2211 492 2212
rect 350 2206 356 2207
rect 358 2209 364 2210
rect 230 2204 236 2205
rect 246 2182 252 2183
rect 246 2178 247 2182
rect 251 2178 252 2182
rect 246 2177 252 2178
rect 166 2175 172 2176
rect 166 2171 167 2175
rect 171 2171 172 2175
rect 166 2170 172 2171
rect 222 2175 228 2176
rect 222 2171 223 2175
rect 227 2171 228 2175
rect 222 2170 228 2171
rect 248 2167 250 2177
rect 352 2176 354 2206
rect 358 2205 359 2209
rect 363 2205 364 2209
rect 486 2207 487 2211
rect 491 2207 492 2211
rect 496 2210 498 2221
rect 614 2211 620 2212
rect 486 2206 492 2207
rect 494 2209 500 2210
rect 358 2204 364 2205
rect 374 2182 380 2183
rect 374 2178 375 2182
rect 379 2178 380 2182
rect 374 2177 380 2178
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 350 2170 356 2171
rect 376 2167 378 2177
rect 488 2176 490 2206
rect 494 2205 495 2209
rect 499 2205 500 2209
rect 614 2207 615 2211
rect 619 2207 620 2211
rect 624 2210 626 2221
rect 646 2211 652 2212
rect 614 2206 620 2207
rect 622 2209 628 2210
rect 494 2204 500 2205
rect 510 2182 516 2183
rect 510 2178 511 2182
rect 515 2178 516 2182
rect 510 2177 516 2178
rect 486 2175 492 2176
rect 486 2171 487 2175
rect 491 2171 492 2175
rect 486 2170 492 2171
rect 512 2167 514 2177
rect 616 2176 618 2206
rect 622 2205 623 2209
rect 627 2205 628 2209
rect 646 2207 647 2211
rect 651 2207 652 2211
rect 752 2210 754 2221
rect 862 2211 868 2212
rect 646 2206 652 2207
rect 750 2209 756 2210
rect 622 2204 628 2205
rect 648 2189 650 2206
rect 750 2205 751 2209
rect 755 2205 756 2209
rect 862 2207 863 2211
rect 867 2207 868 2211
rect 872 2210 874 2221
rect 974 2211 980 2212
rect 862 2206 868 2207
rect 870 2209 876 2210
rect 750 2204 756 2205
rect 647 2188 651 2189
rect 647 2183 651 2184
rect 638 2182 644 2183
rect 638 2178 639 2182
rect 643 2178 644 2182
rect 638 2177 644 2178
rect 766 2182 772 2183
rect 766 2178 767 2182
rect 771 2178 772 2182
rect 766 2177 772 2178
rect 614 2175 620 2176
rect 614 2171 615 2175
rect 619 2171 620 2175
rect 614 2170 620 2171
rect 640 2167 642 2177
rect 768 2167 770 2177
rect 864 2176 866 2206
rect 870 2205 871 2209
rect 875 2205 876 2209
rect 974 2207 975 2211
rect 979 2207 980 2211
rect 984 2210 986 2221
rect 1078 2211 1084 2212
rect 974 2206 980 2207
rect 982 2209 988 2210
rect 870 2204 876 2205
rect 886 2182 892 2183
rect 886 2178 887 2182
rect 891 2178 892 2182
rect 886 2177 892 2178
rect 854 2175 860 2176
rect 854 2171 855 2175
rect 859 2171 860 2175
rect 854 2170 860 2171
rect 862 2175 868 2176
rect 862 2171 863 2175
rect 867 2171 868 2175
rect 862 2170 868 2171
rect 159 2166 163 2167
rect 159 2161 163 2162
rect 215 2166 219 2167
rect 215 2161 219 2162
rect 247 2166 251 2167
rect 247 2161 251 2162
rect 311 2166 315 2167
rect 311 2161 315 2162
rect 375 2166 379 2167
rect 375 2161 379 2162
rect 423 2166 427 2167
rect 423 2161 427 2162
rect 511 2166 515 2167
rect 511 2161 515 2162
rect 543 2166 547 2167
rect 543 2161 547 2162
rect 639 2166 643 2167
rect 639 2161 643 2162
rect 663 2166 667 2167
rect 663 2161 667 2162
rect 767 2166 771 2167
rect 767 2161 771 2162
rect 775 2166 779 2167
rect 775 2161 779 2162
rect 138 2159 144 2160
rect 138 2155 139 2159
rect 143 2155 144 2159
rect 160 2155 162 2161
rect 178 2159 184 2160
rect 178 2155 179 2159
rect 183 2155 184 2159
rect 216 2155 218 2161
rect 234 2159 240 2160
rect 234 2155 235 2159
rect 239 2155 240 2159
rect 312 2155 314 2161
rect 330 2159 336 2160
rect 330 2155 331 2159
rect 335 2155 336 2159
rect 424 2155 426 2161
rect 544 2155 546 2161
rect 562 2159 568 2160
rect 562 2155 563 2159
rect 567 2155 568 2159
rect 664 2155 666 2161
rect 750 2159 756 2160
rect 750 2155 751 2159
rect 755 2155 756 2159
rect 776 2155 778 2161
rect 794 2159 800 2160
rect 794 2155 795 2159
rect 799 2155 800 2159
rect 138 2154 144 2155
rect 158 2154 164 2155
rect 178 2154 184 2155
rect 214 2154 220 2155
rect 234 2154 240 2155
rect 310 2154 316 2155
rect 330 2154 336 2155
rect 422 2154 428 2155
rect 158 2150 159 2154
rect 163 2150 164 2154
rect 158 2149 164 2150
rect 110 2145 116 2146
rect 110 2141 111 2145
rect 115 2141 116 2145
rect 110 2140 116 2141
rect 110 2128 116 2129
rect 110 2124 111 2128
rect 115 2124 116 2128
rect 110 2123 116 2124
rect 142 2127 148 2128
rect 142 2123 143 2127
rect 147 2123 148 2127
rect 180 2124 182 2154
rect 214 2150 215 2154
rect 219 2150 220 2154
rect 214 2149 220 2150
rect 198 2127 204 2128
rect 112 2103 114 2123
rect 142 2122 148 2123
rect 178 2123 184 2124
rect 144 2103 146 2122
rect 178 2119 179 2123
rect 183 2119 184 2123
rect 198 2123 199 2127
rect 203 2123 204 2127
rect 236 2124 238 2154
rect 310 2150 311 2154
rect 315 2150 316 2154
rect 310 2149 316 2150
rect 294 2127 300 2128
rect 198 2122 204 2123
rect 234 2123 240 2124
rect 178 2118 184 2119
rect 200 2103 202 2122
rect 234 2119 235 2123
rect 239 2119 240 2123
rect 294 2123 295 2127
rect 299 2123 300 2127
rect 332 2124 334 2154
rect 422 2150 423 2154
rect 427 2150 428 2154
rect 422 2149 428 2150
rect 542 2154 548 2155
rect 562 2154 568 2155
rect 662 2154 668 2155
rect 750 2154 756 2155
rect 774 2154 780 2155
rect 794 2154 800 2155
rect 542 2150 543 2154
rect 547 2150 548 2154
rect 542 2149 548 2150
rect 406 2127 412 2128
rect 294 2122 300 2123
rect 330 2123 336 2124
rect 234 2118 240 2119
rect 296 2103 298 2122
rect 330 2119 331 2123
rect 335 2119 336 2123
rect 406 2123 407 2127
rect 411 2123 412 2127
rect 406 2122 412 2123
rect 526 2127 532 2128
rect 526 2123 527 2127
rect 531 2123 532 2127
rect 564 2124 566 2154
rect 662 2150 663 2154
rect 667 2150 668 2154
rect 662 2149 668 2150
rect 646 2127 652 2128
rect 526 2122 532 2123
rect 562 2123 568 2124
rect 330 2118 336 2119
rect 408 2103 410 2122
rect 528 2103 530 2122
rect 562 2119 563 2123
rect 567 2119 568 2123
rect 646 2123 647 2127
rect 651 2123 652 2127
rect 646 2122 652 2123
rect 670 2123 676 2124
rect 562 2118 568 2119
rect 648 2103 650 2122
rect 670 2119 671 2123
rect 675 2119 676 2123
rect 670 2118 676 2119
rect 111 2102 115 2103
rect 111 2097 115 2098
rect 143 2102 147 2103
rect 143 2097 147 2098
rect 199 2102 203 2103
rect 199 2097 203 2098
rect 263 2102 267 2103
rect 263 2097 267 2098
rect 295 2102 299 2103
rect 295 2097 299 2098
rect 327 2102 331 2103
rect 327 2097 331 2098
rect 399 2102 403 2103
rect 399 2097 403 2098
rect 407 2102 411 2103
rect 407 2097 411 2098
rect 479 2102 483 2103
rect 479 2097 483 2098
rect 527 2102 531 2103
rect 527 2097 531 2098
rect 567 2102 571 2103
rect 567 2097 571 2098
rect 647 2102 651 2103
rect 647 2097 651 2098
rect 655 2102 659 2103
rect 655 2097 659 2098
rect 112 2085 114 2097
rect 264 2086 266 2097
rect 318 2087 324 2088
rect 262 2085 268 2086
rect 110 2084 116 2085
rect 110 2080 111 2084
rect 115 2080 116 2084
rect 262 2081 263 2085
rect 267 2081 268 2085
rect 318 2083 319 2087
rect 323 2083 324 2087
rect 328 2086 330 2097
rect 390 2087 396 2088
rect 318 2082 324 2083
rect 326 2085 332 2086
rect 262 2080 268 2081
rect 110 2079 116 2080
rect 259 2076 263 2077
rect 259 2071 263 2072
rect 110 2067 116 2068
rect 110 2063 111 2067
rect 115 2063 116 2067
rect 110 2062 116 2063
rect 112 2039 114 2062
rect 260 2052 262 2071
rect 278 2058 284 2059
rect 278 2054 279 2058
rect 283 2054 284 2058
rect 278 2053 284 2054
rect 258 2051 264 2052
rect 258 2047 259 2051
rect 263 2047 264 2051
rect 258 2046 264 2047
rect 280 2039 282 2053
rect 320 2052 322 2082
rect 326 2081 327 2085
rect 331 2081 332 2085
rect 390 2083 391 2087
rect 395 2083 396 2087
rect 400 2086 402 2097
rect 470 2087 476 2088
rect 390 2082 396 2083
rect 398 2085 404 2086
rect 326 2080 332 2081
rect 342 2058 348 2059
rect 342 2054 343 2058
rect 347 2054 348 2058
rect 342 2053 348 2054
rect 318 2051 324 2052
rect 318 2047 319 2051
rect 323 2047 324 2051
rect 318 2046 324 2047
rect 344 2039 346 2053
rect 392 2052 394 2082
rect 398 2081 399 2085
rect 403 2081 404 2085
rect 470 2083 471 2087
rect 475 2083 476 2087
rect 480 2086 482 2097
rect 558 2087 564 2088
rect 470 2082 476 2083
rect 478 2085 484 2086
rect 398 2080 404 2081
rect 414 2058 420 2059
rect 414 2054 415 2058
rect 419 2054 420 2058
rect 414 2053 420 2054
rect 390 2051 396 2052
rect 390 2047 391 2051
rect 395 2047 396 2051
rect 390 2046 396 2047
rect 416 2039 418 2053
rect 472 2052 474 2082
rect 478 2081 479 2085
rect 483 2081 484 2085
rect 558 2083 559 2087
rect 563 2083 564 2087
rect 568 2086 570 2097
rect 646 2087 652 2088
rect 558 2082 564 2083
rect 566 2085 572 2086
rect 478 2080 484 2081
rect 494 2058 500 2059
rect 494 2054 495 2058
rect 499 2054 500 2058
rect 494 2053 500 2054
rect 470 2051 476 2052
rect 470 2047 471 2051
rect 475 2047 476 2051
rect 470 2046 476 2047
rect 496 2039 498 2053
rect 560 2052 562 2082
rect 566 2081 567 2085
rect 571 2081 572 2085
rect 646 2083 647 2087
rect 651 2083 652 2087
rect 656 2086 658 2097
rect 646 2082 652 2083
rect 654 2085 660 2086
rect 566 2080 572 2081
rect 582 2058 588 2059
rect 582 2054 583 2058
rect 587 2054 588 2058
rect 582 2053 588 2054
rect 558 2051 564 2052
rect 558 2047 559 2051
rect 563 2047 564 2051
rect 558 2046 564 2047
rect 584 2039 586 2053
rect 648 2052 650 2082
rect 654 2081 655 2085
rect 659 2081 660 2085
rect 654 2080 660 2081
rect 672 2077 674 2118
rect 735 2102 739 2103
rect 735 2097 739 2098
rect 678 2087 684 2088
rect 678 2083 679 2087
rect 683 2083 684 2087
rect 736 2086 738 2097
rect 752 2096 754 2154
rect 774 2150 775 2154
rect 779 2150 780 2154
rect 774 2149 780 2150
rect 758 2127 764 2128
rect 758 2123 759 2127
rect 763 2123 764 2127
rect 796 2124 798 2154
rect 856 2133 858 2170
rect 888 2167 890 2177
rect 976 2176 978 2206
rect 982 2205 983 2209
rect 987 2205 988 2209
rect 1078 2207 1079 2211
rect 1083 2207 1084 2211
rect 1088 2210 1090 2221
rect 1182 2211 1188 2212
rect 1078 2206 1084 2207
rect 1086 2209 1092 2210
rect 982 2204 988 2205
rect 998 2182 1004 2183
rect 998 2178 999 2182
rect 1003 2178 1004 2182
rect 998 2177 1004 2178
rect 974 2175 980 2176
rect 974 2171 975 2175
rect 979 2171 980 2175
rect 974 2170 980 2171
rect 1000 2167 1002 2177
rect 1080 2176 1082 2206
rect 1086 2205 1087 2209
rect 1091 2205 1092 2209
rect 1182 2207 1183 2211
rect 1187 2207 1188 2211
rect 1192 2210 1194 2221
rect 1200 2220 1202 2278
rect 1206 2274 1207 2278
rect 1211 2274 1212 2278
rect 1206 2273 1212 2274
rect 1270 2251 1276 2252
rect 1270 2247 1271 2251
rect 1275 2247 1276 2251
rect 1270 2246 1276 2247
rect 1272 2227 1274 2246
rect 1280 2236 1282 2278
rect 1286 2274 1287 2278
rect 1291 2274 1292 2278
rect 1286 2273 1292 2274
rect 1308 2248 1310 2290
rect 1327 2285 1331 2286
rect 1328 2270 1330 2285
rect 1368 2283 1370 2306
rect 1414 2302 1420 2303
rect 1414 2298 1415 2302
rect 1419 2298 1420 2302
rect 1414 2297 1420 2298
rect 1416 2283 1418 2297
rect 1448 2296 1450 2326
rect 1454 2325 1455 2329
rect 1459 2325 1460 2329
rect 1502 2327 1503 2331
rect 1507 2327 1508 2331
rect 1512 2330 1514 2341
rect 1502 2326 1508 2327
rect 1510 2329 1516 2330
rect 1454 2324 1460 2325
rect 1470 2302 1476 2303
rect 1470 2298 1471 2302
rect 1475 2298 1476 2302
rect 1470 2297 1476 2298
rect 1446 2295 1452 2296
rect 1446 2291 1447 2295
rect 1451 2291 1452 2295
rect 1446 2290 1452 2291
rect 1472 2283 1474 2297
rect 1504 2296 1506 2326
rect 1510 2325 1511 2329
rect 1515 2325 1516 2329
rect 1510 2324 1516 2325
rect 1526 2302 1532 2303
rect 1526 2298 1527 2302
rect 1531 2298 1532 2302
rect 1526 2297 1532 2298
rect 1502 2295 1508 2296
rect 1502 2291 1503 2295
rect 1507 2291 1508 2295
rect 1502 2290 1508 2291
rect 1528 2283 1530 2297
rect 1536 2296 1538 2354
rect 1544 2347 1546 2358
rect 1578 2355 1579 2359
rect 1583 2355 1584 2359
rect 1646 2359 1647 2363
rect 1651 2359 1652 2363
rect 1684 2360 1686 2390
rect 1758 2386 1759 2390
rect 1763 2386 1764 2390
rect 1758 2385 1764 2386
rect 1854 2390 1860 2391
rect 1854 2386 1855 2390
rect 1859 2386 1860 2390
rect 1854 2385 1860 2386
rect 1942 2390 1948 2391
rect 1942 2386 1943 2390
rect 1947 2386 1948 2390
rect 1942 2385 1948 2386
rect 1742 2363 1748 2364
rect 1646 2358 1652 2359
rect 1682 2359 1688 2360
rect 1578 2354 1584 2355
rect 1648 2347 1650 2358
rect 1682 2355 1683 2359
rect 1687 2355 1688 2359
rect 1742 2359 1743 2363
rect 1747 2359 1748 2363
rect 1742 2358 1748 2359
rect 1838 2363 1844 2364
rect 1838 2359 1839 2363
rect 1843 2359 1844 2363
rect 1926 2363 1932 2364
rect 1838 2358 1844 2359
rect 1862 2359 1868 2360
rect 1682 2354 1688 2355
rect 1744 2347 1746 2358
rect 1840 2347 1842 2358
rect 1862 2355 1863 2359
rect 1867 2355 1868 2359
rect 1926 2359 1927 2363
rect 1931 2359 1932 2363
rect 1964 2360 1966 2406
rect 2008 2403 2010 2413
rect 2072 2412 2074 2442
rect 2078 2441 2079 2445
rect 2083 2441 2084 2445
rect 2158 2443 2159 2447
rect 2163 2443 2164 2447
rect 2168 2446 2170 2457
rect 2210 2451 2216 2452
rect 2210 2447 2211 2451
rect 2215 2447 2216 2451
rect 2210 2446 2216 2447
rect 2158 2442 2164 2443
rect 2166 2445 2172 2446
rect 2078 2440 2084 2441
rect 2094 2418 2100 2419
rect 2094 2414 2095 2418
rect 2099 2414 2100 2418
rect 2094 2413 2100 2414
rect 2070 2411 2076 2412
rect 2070 2407 2071 2411
rect 2075 2407 2076 2411
rect 2070 2406 2076 2407
rect 2054 2403 2060 2404
rect 2096 2403 2098 2413
rect 2160 2412 2162 2442
rect 2166 2441 2167 2445
rect 2171 2441 2172 2445
rect 2166 2440 2172 2441
rect 2182 2418 2188 2419
rect 2182 2414 2183 2418
rect 2187 2414 2188 2418
rect 2182 2413 2188 2414
rect 2158 2411 2164 2412
rect 2158 2407 2159 2411
rect 2163 2407 2164 2411
rect 2158 2406 2164 2407
rect 2184 2403 2186 2413
rect 2007 2402 2011 2403
rect 2007 2397 2011 2398
rect 2039 2402 2043 2403
rect 2054 2399 2055 2403
rect 2059 2399 2060 2403
rect 2054 2398 2060 2399
rect 2095 2402 2099 2403
rect 2039 2397 2043 2398
rect 2014 2395 2020 2396
rect 2014 2391 2015 2395
rect 2019 2391 2020 2395
rect 2040 2391 2042 2397
rect 2014 2390 2020 2391
rect 2038 2390 2044 2391
rect 2016 2372 2018 2390
rect 2038 2386 2039 2390
rect 2043 2386 2044 2390
rect 2038 2385 2044 2386
rect 2014 2371 2020 2372
rect 2014 2367 2015 2371
rect 2019 2367 2020 2371
rect 2014 2366 2020 2367
rect 2022 2363 2028 2364
rect 1926 2358 1932 2359
rect 1962 2359 1968 2360
rect 1862 2354 1868 2355
rect 1543 2346 1547 2347
rect 1543 2341 1547 2342
rect 1567 2346 1571 2347
rect 1567 2341 1571 2342
rect 1639 2346 1643 2347
rect 1639 2341 1643 2342
rect 1647 2346 1651 2347
rect 1647 2341 1651 2342
rect 1727 2346 1731 2347
rect 1727 2341 1731 2342
rect 1743 2346 1747 2347
rect 1743 2341 1747 2342
rect 1823 2346 1827 2347
rect 1823 2341 1827 2342
rect 1839 2346 1843 2347
rect 1839 2341 1843 2342
rect 1568 2330 1570 2341
rect 1630 2331 1636 2332
rect 1566 2329 1572 2330
rect 1566 2325 1567 2329
rect 1571 2325 1572 2329
rect 1630 2327 1631 2331
rect 1635 2327 1636 2331
rect 1640 2330 1642 2341
rect 1718 2331 1724 2332
rect 1630 2326 1636 2327
rect 1638 2329 1644 2330
rect 1566 2324 1572 2325
rect 1582 2302 1588 2303
rect 1582 2298 1583 2302
rect 1587 2298 1588 2302
rect 1582 2297 1588 2298
rect 1534 2295 1540 2296
rect 1534 2291 1535 2295
rect 1539 2291 1540 2295
rect 1534 2290 1540 2291
rect 1584 2283 1586 2297
rect 1632 2296 1634 2326
rect 1638 2325 1639 2329
rect 1643 2325 1644 2329
rect 1718 2327 1719 2331
rect 1723 2327 1724 2331
rect 1728 2330 1730 2341
rect 1814 2331 1820 2332
rect 1718 2326 1724 2327
rect 1726 2329 1732 2330
rect 1638 2324 1644 2325
rect 1654 2302 1660 2303
rect 1654 2298 1655 2302
rect 1659 2298 1660 2302
rect 1654 2297 1660 2298
rect 1630 2295 1636 2296
rect 1630 2291 1631 2295
rect 1635 2291 1636 2295
rect 1630 2290 1636 2291
rect 1656 2283 1658 2297
rect 1720 2296 1722 2326
rect 1726 2325 1727 2329
rect 1731 2325 1732 2329
rect 1814 2327 1815 2331
rect 1819 2327 1820 2331
rect 1824 2330 1826 2341
rect 1814 2326 1820 2327
rect 1822 2329 1828 2330
rect 1726 2324 1732 2325
rect 1742 2302 1748 2303
rect 1742 2298 1743 2302
rect 1747 2298 1748 2302
rect 1742 2297 1748 2298
rect 1718 2295 1724 2296
rect 1718 2291 1719 2295
rect 1723 2291 1724 2295
rect 1718 2290 1724 2291
rect 1744 2283 1746 2297
rect 1367 2282 1371 2283
rect 1367 2277 1371 2278
rect 1415 2282 1419 2283
rect 1415 2277 1419 2278
rect 1471 2282 1475 2283
rect 1471 2277 1475 2278
rect 1495 2282 1499 2283
rect 1495 2277 1499 2278
rect 1527 2282 1531 2283
rect 1527 2277 1531 2278
rect 1583 2282 1587 2283
rect 1583 2277 1587 2278
rect 1615 2282 1619 2283
rect 1615 2277 1619 2278
rect 1655 2282 1659 2283
rect 1735 2282 1739 2283
rect 1655 2277 1659 2278
rect 1662 2279 1668 2280
rect 1326 2269 1332 2270
rect 1326 2265 1327 2269
rect 1331 2265 1332 2269
rect 1326 2264 1332 2265
rect 1368 2262 1370 2277
rect 1390 2275 1396 2276
rect 1390 2271 1391 2275
rect 1395 2271 1396 2275
rect 1416 2271 1418 2277
rect 1486 2275 1492 2276
rect 1486 2271 1487 2275
rect 1491 2271 1492 2275
rect 1496 2271 1498 2277
rect 1616 2271 1618 2277
rect 1662 2275 1663 2279
rect 1667 2275 1668 2279
rect 1735 2277 1739 2278
rect 1743 2282 1747 2283
rect 1743 2277 1747 2278
rect 1662 2274 1668 2275
rect 1710 2275 1716 2276
rect 1390 2270 1396 2271
rect 1414 2270 1420 2271
rect 1486 2270 1492 2271
rect 1494 2270 1500 2271
rect 1366 2261 1372 2262
rect 1366 2257 1367 2261
rect 1371 2257 1372 2261
rect 1366 2256 1372 2257
rect 1326 2252 1332 2253
rect 1392 2252 1394 2270
rect 1414 2266 1415 2270
rect 1419 2266 1420 2270
rect 1414 2265 1420 2266
rect 1326 2248 1327 2252
rect 1331 2248 1332 2252
rect 1306 2247 1312 2248
rect 1326 2247 1332 2248
rect 1390 2251 1396 2252
rect 1390 2247 1391 2251
rect 1395 2247 1396 2251
rect 1306 2243 1307 2247
rect 1311 2243 1312 2247
rect 1306 2242 1312 2243
rect 1278 2235 1284 2236
rect 1278 2231 1279 2235
rect 1283 2231 1284 2235
rect 1278 2230 1284 2231
rect 1328 2227 1330 2247
rect 1390 2246 1396 2247
rect 1366 2244 1372 2245
rect 1366 2240 1367 2244
rect 1371 2240 1372 2244
rect 1366 2239 1372 2240
rect 1398 2243 1404 2244
rect 1398 2239 1399 2243
rect 1403 2239 1404 2243
rect 1271 2226 1275 2227
rect 1271 2221 1275 2222
rect 1327 2226 1331 2227
rect 1327 2221 1331 2222
rect 1198 2219 1204 2220
rect 1198 2215 1199 2219
rect 1203 2215 1204 2219
rect 1198 2214 1204 2215
rect 1262 2211 1268 2212
rect 1182 2206 1188 2207
rect 1190 2209 1196 2210
rect 1086 2204 1092 2205
rect 1102 2182 1108 2183
rect 1102 2178 1103 2182
rect 1107 2178 1108 2182
rect 1102 2177 1108 2178
rect 1078 2175 1084 2176
rect 1078 2171 1079 2175
rect 1083 2171 1084 2175
rect 1078 2170 1084 2171
rect 1104 2167 1106 2177
rect 1184 2176 1186 2206
rect 1190 2205 1191 2209
rect 1195 2205 1196 2209
rect 1262 2207 1263 2211
rect 1267 2207 1268 2211
rect 1272 2210 1274 2221
rect 1262 2206 1268 2207
rect 1270 2209 1276 2210
rect 1328 2209 1330 2221
rect 1368 2215 1370 2239
rect 1398 2238 1404 2239
rect 1478 2243 1484 2244
rect 1478 2239 1479 2243
rect 1483 2239 1484 2243
rect 1478 2238 1484 2239
rect 1400 2215 1402 2238
rect 1480 2215 1482 2238
rect 1488 2232 1490 2270
rect 1494 2266 1495 2270
rect 1499 2266 1500 2270
rect 1494 2265 1500 2266
rect 1614 2270 1620 2271
rect 1614 2266 1615 2270
rect 1619 2266 1620 2270
rect 1614 2265 1620 2266
rect 1598 2243 1604 2244
rect 1598 2239 1599 2243
rect 1603 2239 1604 2243
rect 1598 2238 1604 2239
rect 1486 2231 1492 2232
rect 1486 2227 1487 2231
rect 1491 2227 1492 2231
rect 1486 2226 1492 2227
rect 1600 2215 1602 2238
rect 1367 2214 1371 2215
rect 1367 2209 1371 2210
rect 1399 2214 1403 2215
rect 1399 2209 1403 2210
rect 1455 2214 1459 2215
rect 1455 2209 1459 2210
rect 1479 2214 1483 2215
rect 1479 2209 1483 2210
rect 1535 2214 1539 2215
rect 1535 2209 1539 2210
rect 1599 2214 1603 2215
rect 1599 2209 1603 2210
rect 1631 2214 1635 2215
rect 1631 2209 1635 2210
rect 1190 2204 1196 2205
rect 1206 2182 1212 2183
rect 1206 2178 1207 2182
rect 1211 2178 1212 2182
rect 1206 2177 1212 2178
rect 1182 2175 1188 2176
rect 1182 2171 1183 2175
rect 1187 2171 1188 2175
rect 1182 2170 1188 2171
rect 1208 2167 1210 2177
rect 1264 2176 1266 2206
rect 1270 2205 1271 2209
rect 1275 2205 1276 2209
rect 1270 2204 1276 2205
rect 1326 2208 1332 2209
rect 1326 2204 1327 2208
rect 1331 2204 1332 2208
rect 1326 2203 1332 2204
rect 1368 2197 1370 2209
rect 1456 2198 1458 2209
rect 1526 2199 1532 2200
rect 1454 2197 1460 2198
rect 1366 2196 1372 2197
rect 1366 2192 1367 2196
rect 1371 2192 1372 2196
rect 1454 2193 1455 2197
rect 1459 2193 1460 2197
rect 1526 2195 1527 2199
rect 1531 2195 1532 2199
rect 1536 2198 1538 2209
rect 1622 2199 1628 2200
rect 1526 2194 1532 2195
rect 1534 2197 1540 2198
rect 1454 2192 1460 2193
rect 1326 2191 1332 2192
rect 1366 2191 1372 2192
rect 1326 2187 1327 2191
rect 1331 2187 1332 2191
rect 1326 2186 1332 2187
rect 1286 2182 1292 2183
rect 1286 2178 1287 2182
rect 1291 2178 1292 2182
rect 1286 2177 1292 2178
rect 1262 2175 1268 2176
rect 1262 2171 1263 2175
rect 1267 2171 1268 2175
rect 1262 2170 1268 2171
rect 1288 2167 1290 2177
rect 1328 2167 1330 2186
rect 1366 2179 1372 2180
rect 1366 2175 1367 2179
rect 1371 2175 1372 2179
rect 1366 2174 1372 2175
rect 879 2166 883 2167
rect 879 2161 883 2162
rect 887 2166 891 2167
rect 887 2161 891 2162
rect 975 2166 979 2167
rect 975 2161 979 2162
rect 999 2166 1003 2167
rect 999 2161 1003 2162
rect 1071 2166 1075 2167
rect 1071 2161 1075 2162
rect 1103 2166 1107 2167
rect 1103 2161 1107 2162
rect 1167 2166 1171 2167
rect 1167 2161 1171 2162
rect 1207 2166 1211 2167
rect 1207 2161 1211 2162
rect 1271 2166 1275 2167
rect 1271 2161 1275 2162
rect 1287 2166 1291 2167
rect 1287 2161 1291 2162
rect 1327 2166 1331 2167
rect 1327 2161 1331 2162
rect 880 2155 882 2161
rect 898 2159 904 2160
rect 898 2155 899 2159
rect 903 2155 904 2159
rect 976 2155 978 2161
rect 1072 2155 1074 2161
rect 1090 2159 1096 2160
rect 1090 2155 1091 2159
rect 1095 2155 1096 2159
rect 1168 2155 1170 2161
rect 1272 2155 1274 2161
rect 878 2154 884 2155
rect 898 2154 904 2155
rect 974 2154 980 2155
rect 878 2150 879 2154
rect 883 2150 884 2154
rect 878 2149 884 2150
rect 855 2132 859 2133
rect 855 2127 859 2128
rect 862 2127 868 2128
rect 758 2122 764 2123
rect 794 2123 800 2124
rect 760 2103 762 2122
rect 794 2119 795 2123
rect 799 2119 800 2123
rect 862 2123 863 2127
rect 867 2123 868 2127
rect 900 2124 902 2154
rect 974 2150 975 2154
rect 979 2150 980 2154
rect 974 2149 980 2150
rect 1070 2154 1076 2155
rect 1090 2154 1096 2155
rect 1166 2154 1172 2155
rect 1070 2150 1071 2154
rect 1075 2150 1076 2154
rect 1070 2149 1076 2150
rect 958 2127 964 2128
rect 862 2122 868 2123
rect 898 2123 904 2124
rect 794 2118 800 2119
rect 864 2103 866 2122
rect 898 2119 899 2123
rect 903 2119 904 2123
rect 958 2123 959 2127
rect 963 2123 964 2127
rect 958 2122 964 2123
rect 1054 2127 1060 2128
rect 1054 2123 1055 2127
rect 1059 2123 1060 2127
rect 1092 2124 1094 2154
rect 1166 2150 1167 2154
rect 1171 2150 1172 2154
rect 1166 2149 1172 2150
rect 1270 2154 1276 2155
rect 1270 2150 1271 2154
rect 1275 2150 1276 2154
rect 1270 2149 1276 2150
rect 1328 2146 1330 2161
rect 1368 2159 1370 2174
rect 1470 2170 1476 2171
rect 1470 2166 1471 2170
rect 1475 2166 1476 2170
rect 1470 2165 1476 2166
rect 1472 2159 1474 2165
rect 1528 2164 1530 2194
rect 1534 2193 1535 2197
rect 1539 2193 1540 2197
rect 1622 2195 1623 2199
rect 1627 2195 1628 2199
rect 1632 2198 1634 2209
rect 1664 2200 1666 2274
rect 1710 2271 1711 2275
rect 1715 2271 1716 2275
rect 1736 2271 1738 2277
rect 1816 2276 1818 2326
rect 1822 2325 1823 2329
rect 1827 2325 1828 2329
rect 1822 2324 1828 2325
rect 1838 2302 1844 2303
rect 1838 2298 1839 2302
rect 1843 2298 1844 2302
rect 1838 2297 1844 2298
rect 1840 2283 1842 2297
rect 1864 2296 1866 2354
rect 1928 2347 1930 2358
rect 1962 2355 1963 2359
rect 1967 2355 1968 2359
rect 2022 2359 2023 2363
rect 2027 2359 2028 2363
rect 2056 2360 2058 2398
rect 2095 2397 2099 2398
rect 2135 2402 2139 2403
rect 2135 2397 2139 2398
rect 2183 2402 2187 2403
rect 2183 2397 2187 2398
rect 2126 2395 2132 2396
rect 2126 2391 2127 2395
rect 2131 2391 2132 2395
rect 2136 2391 2138 2397
rect 2212 2396 2214 2446
rect 2256 2412 2258 2470
rect 2280 2463 2282 2474
rect 2314 2471 2315 2475
rect 2319 2471 2320 2475
rect 2382 2475 2383 2479
rect 2387 2475 2388 2479
rect 2382 2474 2388 2475
rect 2314 2470 2320 2471
rect 2384 2463 2386 2474
rect 2263 2462 2267 2463
rect 2263 2457 2267 2458
rect 2279 2462 2283 2463
rect 2279 2457 2283 2458
rect 2359 2462 2363 2463
rect 2359 2457 2363 2458
rect 2383 2462 2387 2463
rect 2383 2457 2387 2458
rect 2264 2446 2266 2457
rect 2360 2446 2362 2457
rect 2392 2448 2394 2506
rect 2398 2502 2399 2506
rect 2403 2502 2404 2506
rect 2398 2501 2404 2502
rect 2584 2498 2586 2513
rect 2582 2497 2588 2498
rect 2582 2493 2583 2497
rect 2587 2493 2588 2497
rect 2582 2492 2588 2493
rect 2582 2480 2588 2481
rect 2582 2476 2583 2480
rect 2587 2476 2588 2480
rect 2582 2475 2588 2476
rect 2584 2463 2586 2475
rect 2455 2462 2459 2463
rect 2455 2457 2459 2458
rect 2527 2462 2531 2463
rect 2527 2457 2531 2458
rect 2583 2462 2587 2463
rect 2583 2457 2587 2458
rect 2390 2447 2396 2448
rect 2262 2445 2268 2446
rect 2262 2441 2263 2445
rect 2267 2441 2268 2445
rect 2262 2440 2268 2441
rect 2358 2445 2364 2446
rect 2358 2441 2359 2445
rect 2363 2441 2364 2445
rect 2390 2443 2391 2447
rect 2395 2443 2396 2447
rect 2456 2446 2458 2457
rect 2462 2451 2468 2452
rect 2462 2447 2463 2451
rect 2467 2447 2468 2451
rect 2462 2446 2468 2447
rect 2528 2446 2530 2457
rect 2390 2442 2396 2443
rect 2454 2445 2460 2446
rect 2358 2440 2364 2441
rect 2454 2441 2455 2445
rect 2459 2441 2460 2445
rect 2454 2440 2460 2441
rect 2278 2418 2284 2419
rect 2278 2414 2279 2418
rect 2283 2414 2284 2418
rect 2278 2413 2284 2414
rect 2374 2418 2380 2419
rect 2374 2414 2375 2418
rect 2379 2414 2380 2418
rect 2374 2413 2380 2414
rect 2254 2411 2260 2412
rect 2254 2407 2255 2411
rect 2259 2407 2260 2411
rect 2254 2406 2260 2407
rect 2280 2403 2282 2413
rect 2376 2403 2378 2413
rect 2464 2412 2466 2446
rect 2526 2445 2532 2446
rect 2584 2445 2586 2457
rect 2526 2441 2527 2445
rect 2531 2441 2532 2445
rect 2526 2440 2532 2441
rect 2582 2444 2588 2445
rect 2582 2440 2583 2444
rect 2587 2440 2588 2444
rect 2582 2439 2588 2440
rect 2582 2427 2588 2428
rect 2582 2423 2583 2427
rect 2587 2423 2588 2427
rect 2582 2422 2588 2423
rect 2470 2418 2476 2419
rect 2470 2414 2471 2418
rect 2475 2414 2476 2418
rect 2470 2413 2476 2414
rect 2542 2418 2548 2419
rect 2542 2414 2543 2418
rect 2547 2414 2548 2418
rect 2542 2413 2548 2414
rect 2438 2411 2444 2412
rect 2438 2407 2439 2411
rect 2443 2407 2444 2411
rect 2438 2406 2444 2407
rect 2462 2411 2468 2412
rect 2462 2407 2463 2411
rect 2467 2407 2468 2411
rect 2462 2406 2468 2407
rect 2231 2402 2235 2403
rect 2231 2397 2235 2398
rect 2279 2402 2283 2403
rect 2279 2397 2283 2398
rect 2335 2402 2339 2403
rect 2335 2397 2339 2398
rect 2375 2402 2379 2403
rect 2375 2397 2379 2398
rect 2210 2395 2216 2396
rect 2210 2391 2211 2395
rect 2215 2391 2216 2395
rect 2232 2391 2234 2397
rect 2246 2395 2252 2396
rect 2246 2391 2247 2395
rect 2251 2391 2252 2395
rect 2336 2391 2338 2397
rect 2422 2395 2428 2396
rect 2422 2391 2423 2395
rect 2427 2391 2428 2395
rect 2126 2390 2132 2391
rect 2134 2390 2140 2391
rect 2210 2390 2216 2391
rect 2230 2390 2236 2391
rect 2246 2390 2252 2391
rect 2334 2390 2340 2391
rect 2422 2390 2428 2391
rect 2118 2363 2124 2364
rect 2022 2358 2028 2359
rect 2054 2359 2060 2360
rect 1962 2354 1968 2355
rect 2024 2347 2026 2358
rect 2054 2355 2055 2359
rect 2059 2355 2060 2359
rect 2118 2359 2119 2363
rect 2123 2359 2124 2363
rect 2118 2358 2124 2359
rect 2054 2354 2060 2355
rect 2120 2347 2122 2358
rect 1927 2346 1931 2347
rect 1927 2341 1931 2342
rect 1943 2346 1947 2347
rect 1943 2341 1947 2342
rect 2023 2346 2027 2347
rect 2023 2341 2027 2342
rect 2079 2346 2083 2347
rect 2079 2341 2083 2342
rect 2119 2346 2123 2347
rect 2119 2341 2123 2342
rect 1934 2331 1940 2332
rect 1934 2327 1935 2331
rect 1939 2327 1940 2331
rect 1944 2330 1946 2341
rect 2070 2331 2076 2332
rect 1934 2326 1940 2327
rect 1942 2329 1948 2330
rect 1936 2296 1938 2326
rect 1942 2325 1943 2329
rect 1947 2325 1948 2329
rect 2070 2327 2071 2331
rect 2075 2327 2076 2331
rect 2080 2330 2082 2341
rect 2128 2340 2130 2390
rect 2134 2386 2135 2390
rect 2139 2386 2140 2390
rect 2134 2385 2140 2386
rect 2230 2386 2231 2390
rect 2235 2386 2236 2390
rect 2230 2385 2236 2386
rect 2214 2363 2220 2364
rect 2214 2359 2215 2363
rect 2219 2359 2220 2363
rect 2248 2360 2250 2390
rect 2334 2386 2335 2390
rect 2339 2386 2340 2390
rect 2334 2385 2340 2386
rect 2318 2363 2324 2364
rect 2214 2358 2220 2359
rect 2246 2359 2252 2360
rect 2216 2347 2218 2358
rect 2246 2355 2247 2359
rect 2251 2355 2252 2359
rect 2318 2359 2319 2363
rect 2323 2359 2324 2363
rect 2318 2358 2324 2359
rect 2374 2359 2380 2360
rect 2246 2354 2252 2355
rect 2320 2347 2322 2358
rect 2374 2355 2375 2359
rect 2379 2355 2380 2359
rect 2374 2354 2380 2355
rect 2215 2346 2219 2347
rect 2215 2341 2219 2342
rect 2223 2346 2227 2347
rect 2223 2341 2227 2342
rect 2319 2346 2323 2347
rect 2319 2341 2323 2342
rect 2126 2339 2132 2340
rect 2126 2335 2127 2339
rect 2131 2335 2132 2339
rect 2126 2334 2132 2335
rect 2214 2331 2220 2332
rect 2070 2326 2076 2327
rect 2078 2329 2084 2330
rect 1942 2324 1948 2325
rect 1958 2302 1964 2303
rect 1958 2298 1959 2302
rect 1963 2298 1964 2302
rect 1958 2297 1964 2298
rect 1862 2295 1868 2296
rect 1862 2291 1863 2295
rect 1867 2291 1868 2295
rect 1862 2290 1868 2291
rect 1934 2295 1940 2296
rect 1934 2291 1935 2295
rect 1939 2291 1940 2295
rect 1934 2290 1940 2291
rect 1960 2283 1962 2297
rect 2072 2296 2074 2326
rect 2078 2325 2079 2329
rect 2083 2325 2084 2329
rect 2214 2327 2215 2331
rect 2219 2327 2220 2331
rect 2224 2330 2226 2341
rect 2214 2326 2220 2327
rect 2222 2329 2228 2330
rect 2078 2324 2084 2325
rect 2094 2302 2100 2303
rect 2094 2298 2095 2302
rect 2099 2298 2100 2302
rect 2094 2297 2100 2298
rect 2070 2295 2076 2296
rect 2070 2291 2071 2295
rect 2075 2291 2076 2295
rect 2070 2290 2076 2291
rect 2096 2283 2098 2297
rect 2216 2296 2218 2326
rect 2222 2325 2223 2329
rect 2227 2325 2228 2329
rect 2222 2324 2228 2325
rect 2238 2302 2244 2303
rect 2238 2298 2239 2302
rect 2243 2298 2244 2302
rect 2238 2297 2244 2298
rect 2214 2295 2220 2296
rect 2214 2291 2215 2295
rect 2219 2291 2220 2295
rect 2214 2290 2220 2291
rect 2240 2283 2242 2297
rect 2376 2296 2378 2354
rect 2383 2346 2387 2347
rect 2383 2341 2387 2342
rect 2384 2330 2386 2341
rect 2414 2331 2420 2332
rect 2382 2329 2388 2330
rect 2382 2325 2383 2329
rect 2387 2325 2388 2329
rect 2414 2327 2415 2331
rect 2419 2327 2420 2331
rect 2414 2326 2420 2327
rect 2382 2324 2388 2325
rect 2398 2302 2404 2303
rect 2398 2298 2399 2302
rect 2403 2298 2404 2302
rect 2398 2297 2404 2298
rect 2374 2295 2380 2296
rect 2374 2291 2375 2295
rect 2379 2291 2380 2295
rect 2374 2290 2380 2291
rect 2400 2283 2402 2297
rect 2416 2284 2418 2326
rect 2414 2283 2420 2284
rect 1839 2282 1843 2283
rect 1839 2277 1843 2278
rect 1855 2282 1859 2283
rect 1855 2277 1859 2278
rect 1959 2282 1963 2283
rect 1959 2277 1963 2278
rect 1967 2282 1971 2283
rect 1967 2277 1971 2278
rect 2071 2282 2075 2283
rect 2071 2277 2075 2278
rect 2095 2282 2099 2283
rect 2095 2277 2099 2278
rect 2167 2282 2171 2283
rect 2167 2277 2171 2278
rect 2239 2282 2243 2283
rect 2239 2277 2243 2278
rect 2255 2282 2259 2283
rect 2255 2277 2259 2278
rect 2335 2282 2339 2283
rect 2335 2277 2339 2278
rect 2399 2282 2403 2283
rect 2399 2277 2403 2278
rect 2407 2282 2411 2283
rect 2414 2279 2415 2283
rect 2419 2279 2420 2283
rect 2414 2278 2420 2279
rect 2407 2277 2411 2278
rect 1814 2275 1820 2276
rect 1814 2271 1815 2275
rect 1819 2271 1820 2275
rect 1856 2271 1858 2277
rect 1968 2271 1970 2277
rect 1986 2275 1992 2276
rect 1986 2271 1987 2275
rect 1991 2271 1992 2275
rect 2072 2271 2074 2277
rect 2168 2271 2170 2277
rect 2186 2275 2192 2276
rect 2186 2271 2187 2275
rect 2191 2271 2192 2275
rect 2256 2271 2258 2277
rect 2274 2275 2280 2276
rect 2274 2271 2275 2275
rect 2279 2271 2280 2275
rect 2336 2271 2338 2277
rect 2382 2275 2388 2276
rect 2382 2271 2383 2275
rect 2387 2271 2388 2275
rect 2408 2271 2410 2277
rect 2414 2275 2420 2276
rect 2414 2271 2415 2275
rect 2419 2271 2420 2275
rect 1710 2270 1716 2271
rect 1734 2270 1740 2271
rect 1814 2270 1820 2271
rect 1854 2270 1860 2271
rect 1712 2252 1714 2270
rect 1734 2266 1735 2270
rect 1739 2266 1740 2270
rect 1734 2265 1740 2266
rect 1854 2266 1855 2270
rect 1859 2266 1860 2270
rect 1854 2265 1860 2266
rect 1966 2270 1972 2271
rect 1986 2270 1992 2271
rect 2070 2270 2076 2271
rect 1966 2266 1967 2270
rect 1971 2266 1972 2270
rect 1966 2265 1972 2266
rect 1710 2251 1716 2252
rect 1710 2247 1711 2251
rect 1715 2247 1716 2251
rect 1710 2246 1716 2247
rect 1718 2243 1724 2244
rect 1718 2239 1719 2243
rect 1723 2239 1724 2243
rect 1838 2243 1844 2244
rect 1718 2238 1724 2239
rect 1750 2239 1756 2240
rect 1720 2215 1722 2238
rect 1750 2235 1751 2239
rect 1755 2235 1756 2239
rect 1838 2239 1839 2243
rect 1843 2239 1844 2243
rect 1838 2238 1844 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1988 2240 1990 2270
rect 2070 2266 2071 2270
rect 2075 2266 2076 2270
rect 2070 2265 2076 2266
rect 2166 2270 2172 2271
rect 2186 2270 2192 2271
rect 2254 2270 2260 2271
rect 2274 2270 2280 2271
rect 2334 2270 2340 2271
rect 2382 2270 2388 2271
rect 2406 2270 2412 2271
rect 2414 2270 2420 2271
rect 2166 2266 2167 2270
rect 2171 2266 2172 2270
rect 2166 2265 2172 2266
rect 2054 2243 2060 2244
rect 1950 2238 1956 2239
rect 1986 2239 1992 2240
rect 1750 2234 1756 2235
rect 1719 2214 1723 2215
rect 1719 2209 1723 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1662 2199 1668 2200
rect 1622 2194 1628 2195
rect 1630 2197 1636 2198
rect 1534 2192 1540 2193
rect 1550 2170 1556 2171
rect 1550 2166 1551 2170
rect 1555 2166 1556 2170
rect 1550 2165 1556 2166
rect 1526 2163 1532 2164
rect 1526 2159 1527 2163
rect 1531 2159 1532 2163
rect 1552 2159 1554 2165
rect 1624 2164 1626 2194
rect 1630 2193 1631 2197
rect 1635 2193 1636 2197
rect 1662 2195 1663 2199
rect 1667 2195 1668 2199
rect 1744 2198 1746 2209
rect 1662 2194 1668 2195
rect 1742 2197 1748 2198
rect 1630 2192 1636 2193
rect 1742 2193 1743 2197
rect 1747 2193 1748 2197
rect 1742 2192 1748 2193
rect 1646 2170 1652 2171
rect 1646 2166 1647 2170
rect 1651 2166 1652 2170
rect 1646 2165 1652 2166
rect 1622 2163 1628 2164
rect 1622 2159 1623 2163
rect 1627 2159 1628 2163
rect 1648 2159 1650 2165
rect 1752 2164 1754 2234
rect 1840 2215 1842 2238
rect 1952 2215 1954 2238
rect 1986 2235 1987 2239
rect 1991 2235 1992 2239
rect 2054 2239 2055 2243
rect 2059 2239 2060 2243
rect 2054 2238 2060 2239
rect 2150 2243 2156 2244
rect 2150 2239 2151 2243
rect 2155 2239 2156 2243
rect 2188 2240 2190 2270
rect 2254 2266 2255 2270
rect 2259 2266 2260 2270
rect 2254 2265 2260 2266
rect 2238 2243 2244 2244
rect 2150 2238 2156 2239
rect 2186 2239 2192 2240
rect 1986 2234 1992 2235
rect 2056 2215 2058 2238
rect 2152 2215 2154 2238
rect 2186 2235 2187 2239
rect 2191 2235 2192 2239
rect 2238 2239 2239 2243
rect 2243 2239 2244 2243
rect 2276 2240 2278 2270
rect 2334 2266 2335 2270
rect 2339 2266 2340 2270
rect 2334 2265 2340 2266
rect 2318 2243 2324 2244
rect 2238 2238 2244 2239
rect 2274 2239 2280 2240
rect 2186 2234 2192 2235
rect 2240 2215 2242 2238
rect 2274 2235 2275 2239
rect 2279 2235 2280 2239
rect 2318 2239 2319 2243
rect 2323 2239 2324 2243
rect 2318 2238 2324 2239
rect 2274 2234 2280 2235
rect 2320 2215 2322 2238
rect 1839 2214 1843 2215
rect 1839 2209 1843 2210
rect 1863 2214 1867 2215
rect 1863 2209 1867 2210
rect 1951 2214 1955 2215
rect 1951 2209 1955 2210
rect 1983 2214 1987 2215
rect 1983 2209 1987 2210
rect 2055 2214 2059 2215
rect 2055 2209 2059 2210
rect 2095 2214 2099 2215
rect 2095 2209 2099 2210
rect 2151 2214 2155 2215
rect 2151 2209 2155 2210
rect 2207 2214 2211 2215
rect 2207 2209 2211 2210
rect 2239 2214 2243 2215
rect 2239 2209 2243 2210
rect 2311 2214 2315 2215
rect 2311 2209 2315 2210
rect 2319 2214 2323 2215
rect 2319 2209 2323 2210
rect 1854 2199 1860 2200
rect 1854 2195 1855 2199
rect 1859 2195 1860 2199
rect 1864 2198 1866 2209
rect 1974 2199 1980 2200
rect 1854 2194 1860 2195
rect 1862 2197 1868 2198
rect 1758 2170 1764 2171
rect 1758 2166 1759 2170
rect 1763 2166 1764 2170
rect 1758 2165 1764 2166
rect 1750 2163 1756 2164
rect 1750 2159 1751 2163
rect 1755 2159 1756 2163
rect 1760 2159 1762 2165
rect 1856 2164 1858 2194
rect 1862 2193 1863 2197
rect 1867 2193 1868 2197
rect 1974 2195 1975 2199
rect 1979 2195 1980 2199
rect 1984 2198 1986 2209
rect 2006 2199 2012 2200
rect 1974 2194 1980 2195
rect 1982 2197 1988 2198
rect 1862 2192 1868 2193
rect 1878 2170 1884 2171
rect 1878 2166 1879 2170
rect 1883 2166 1884 2170
rect 1878 2165 1884 2166
rect 1854 2163 1860 2164
rect 1854 2159 1855 2163
rect 1859 2159 1860 2163
rect 1880 2159 1882 2165
rect 1976 2164 1978 2194
rect 1982 2193 1983 2197
rect 1987 2193 1988 2197
rect 2006 2195 2007 2199
rect 2011 2195 2012 2199
rect 2096 2198 2098 2209
rect 2198 2199 2204 2200
rect 2006 2194 2012 2195
rect 2094 2197 2100 2198
rect 1982 2192 1988 2193
rect 1998 2170 2004 2171
rect 1998 2166 1999 2170
rect 2003 2166 2004 2170
rect 1998 2165 2004 2166
rect 1974 2163 1980 2164
rect 1974 2159 1975 2163
rect 1979 2159 1980 2163
rect 2000 2159 2002 2165
rect 1367 2158 1371 2159
rect 1367 2153 1371 2154
rect 1471 2158 1475 2159
rect 1526 2158 1532 2159
rect 1535 2158 1539 2159
rect 1471 2153 1475 2154
rect 1551 2158 1555 2159
rect 1622 2158 1628 2159
rect 1631 2158 1635 2159
rect 1535 2153 1539 2154
rect 1542 2155 1548 2156
rect 1326 2145 1332 2146
rect 1326 2141 1327 2145
rect 1331 2141 1332 2145
rect 1326 2140 1332 2141
rect 1368 2138 1370 2153
rect 1510 2151 1516 2152
rect 1510 2147 1511 2151
rect 1515 2147 1516 2151
rect 1536 2147 1538 2153
rect 1542 2151 1543 2155
rect 1547 2151 1548 2155
rect 1551 2153 1555 2154
rect 1631 2153 1635 2154
rect 1647 2158 1651 2159
rect 1647 2153 1651 2154
rect 1735 2158 1739 2159
rect 1750 2158 1756 2159
rect 1759 2158 1763 2159
rect 1735 2153 1739 2154
rect 1759 2153 1763 2154
rect 1839 2158 1843 2159
rect 1854 2158 1860 2159
rect 1879 2158 1883 2159
rect 1839 2153 1843 2154
rect 1879 2153 1883 2154
rect 1951 2158 1955 2159
rect 1974 2158 1980 2159
rect 1999 2158 2003 2159
rect 1951 2153 1955 2154
rect 2008 2156 2010 2194
rect 2094 2193 2095 2197
rect 2099 2193 2100 2197
rect 2198 2195 2199 2199
rect 2203 2195 2204 2199
rect 2208 2198 2210 2209
rect 2302 2199 2308 2200
rect 2198 2194 2204 2195
rect 2206 2197 2212 2198
rect 2094 2192 2100 2193
rect 2110 2170 2116 2171
rect 2110 2166 2111 2170
rect 2115 2166 2116 2170
rect 2110 2165 2116 2166
rect 2074 2163 2080 2164
rect 2074 2159 2075 2163
rect 2079 2159 2080 2163
rect 2112 2159 2114 2165
rect 2200 2164 2202 2194
rect 2206 2193 2207 2197
rect 2211 2193 2212 2197
rect 2302 2195 2303 2199
rect 2307 2195 2308 2199
rect 2312 2198 2314 2209
rect 2384 2204 2386 2270
rect 2406 2266 2407 2270
rect 2411 2266 2412 2270
rect 2406 2265 2412 2266
rect 2390 2243 2396 2244
rect 2390 2239 2391 2243
rect 2395 2239 2396 2243
rect 2390 2238 2396 2239
rect 2392 2215 2394 2238
rect 2416 2236 2418 2270
rect 2424 2240 2426 2390
rect 2430 2363 2436 2364
rect 2430 2359 2431 2363
rect 2435 2359 2436 2363
rect 2430 2358 2436 2359
rect 2432 2347 2434 2358
rect 2440 2356 2442 2406
rect 2472 2403 2474 2413
rect 2544 2403 2546 2413
rect 2558 2411 2564 2412
rect 2558 2407 2559 2411
rect 2563 2407 2564 2411
rect 2558 2406 2564 2407
rect 2447 2402 2451 2403
rect 2447 2397 2451 2398
rect 2471 2402 2475 2403
rect 2471 2397 2475 2398
rect 2543 2402 2547 2403
rect 2543 2397 2547 2398
rect 2448 2391 2450 2397
rect 2534 2395 2540 2396
rect 2534 2391 2535 2395
rect 2539 2391 2540 2395
rect 2544 2391 2546 2397
rect 2446 2390 2452 2391
rect 2534 2390 2540 2391
rect 2542 2390 2548 2391
rect 2446 2386 2447 2390
rect 2451 2386 2452 2390
rect 2446 2385 2452 2386
rect 2526 2363 2532 2364
rect 2526 2359 2527 2363
rect 2531 2359 2532 2363
rect 2526 2358 2532 2359
rect 2438 2355 2444 2356
rect 2438 2351 2439 2355
rect 2443 2351 2444 2355
rect 2438 2350 2444 2351
rect 2528 2347 2530 2358
rect 2431 2346 2435 2347
rect 2431 2341 2435 2342
rect 2527 2346 2531 2347
rect 2527 2341 2531 2342
rect 2528 2330 2530 2341
rect 2536 2336 2538 2390
rect 2542 2386 2543 2390
rect 2547 2386 2548 2390
rect 2542 2385 2548 2386
rect 2560 2360 2562 2406
rect 2584 2403 2586 2422
rect 2583 2402 2587 2403
rect 2583 2397 2587 2398
rect 2584 2382 2586 2397
rect 2582 2381 2588 2382
rect 2582 2377 2583 2381
rect 2587 2377 2588 2381
rect 2582 2376 2588 2377
rect 2582 2364 2588 2365
rect 2582 2360 2583 2364
rect 2587 2360 2588 2364
rect 2558 2359 2564 2360
rect 2582 2359 2588 2360
rect 2558 2355 2559 2359
rect 2563 2355 2564 2359
rect 2558 2354 2564 2355
rect 2584 2347 2586 2359
rect 2583 2346 2587 2347
rect 2583 2341 2587 2342
rect 2534 2335 2540 2336
rect 2534 2331 2535 2335
rect 2539 2331 2540 2335
rect 2534 2330 2540 2331
rect 2526 2329 2532 2330
rect 2584 2329 2586 2341
rect 2526 2325 2527 2329
rect 2531 2325 2532 2329
rect 2526 2324 2532 2325
rect 2582 2328 2588 2329
rect 2582 2324 2583 2328
rect 2587 2324 2588 2328
rect 2582 2323 2588 2324
rect 2582 2311 2588 2312
rect 2582 2307 2583 2311
rect 2587 2307 2588 2311
rect 2582 2306 2588 2307
rect 2542 2302 2548 2303
rect 2542 2298 2543 2302
rect 2547 2298 2548 2302
rect 2542 2297 2548 2298
rect 2544 2283 2546 2297
rect 2558 2295 2564 2296
rect 2558 2291 2559 2295
rect 2563 2291 2564 2295
rect 2558 2290 2564 2291
rect 2487 2282 2491 2283
rect 2487 2277 2491 2278
rect 2543 2282 2547 2283
rect 2543 2277 2547 2278
rect 2488 2271 2490 2277
rect 2506 2275 2512 2276
rect 2506 2271 2507 2275
rect 2511 2271 2512 2275
rect 2544 2271 2546 2277
rect 2486 2270 2492 2271
rect 2506 2270 2512 2271
rect 2542 2270 2548 2271
rect 2486 2266 2487 2270
rect 2491 2266 2492 2270
rect 2486 2265 2492 2266
rect 2470 2243 2476 2244
rect 2422 2239 2428 2240
rect 2414 2235 2420 2236
rect 2414 2231 2415 2235
rect 2419 2231 2420 2235
rect 2422 2235 2423 2239
rect 2427 2235 2428 2239
rect 2470 2239 2471 2243
rect 2475 2239 2476 2243
rect 2508 2240 2510 2270
rect 2542 2266 2543 2270
rect 2547 2266 2548 2270
rect 2542 2265 2548 2266
rect 2526 2243 2532 2244
rect 2470 2238 2476 2239
rect 2506 2239 2512 2240
rect 2422 2234 2428 2235
rect 2414 2230 2420 2231
rect 2472 2215 2474 2238
rect 2506 2235 2507 2239
rect 2511 2235 2512 2239
rect 2526 2239 2527 2243
rect 2531 2239 2532 2243
rect 2560 2240 2562 2290
rect 2584 2283 2586 2306
rect 2583 2282 2587 2283
rect 2583 2277 2587 2278
rect 2584 2262 2586 2277
rect 2582 2261 2588 2262
rect 2582 2257 2583 2261
rect 2587 2257 2588 2261
rect 2582 2256 2588 2257
rect 2582 2244 2588 2245
rect 2582 2240 2583 2244
rect 2587 2240 2588 2244
rect 2526 2238 2532 2239
rect 2558 2239 2564 2240
rect 2582 2239 2588 2240
rect 2506 2234 2512 2235
rect 2528 2215 2530 2238
rect 2558 2235 2559 2239
rect 2563 2235 2564 2239
rect 2558 2234 2564 2235
rect 2584 2215 2586 2239
rect 2391 2214 2395 2215
rect 2391 2209 2395 2210
rect 2423 2214 2427 2215
rect 2423 2209 2427 2210
rect 2471 2214 2475 2215
rect 2471 2209 2475 2210
rect 2527 2214 2531 2215
rect 2527 2209 2531 2210
rect 2583 2214 2587 2215
rect 2583 2209 2587 2210
rect 2382 2203 2388 2204
rect 2338 2199 2344 2200
rect 2302 2194 2308 2195
rect 2310 2197 2316 2198
rect 2206 2192 2212 2193
rect 2222 2170 2228 2171
rect 2222 2166 2223 2170
rect 2227 2166 2228 2170
rect 2222 2165 2228 2166
rect 2198 2163 2204 2164
rect 2198 2159 2199 2163
rect 2203 2159 2204 2163
rect 2224 2159 2226 2165
rect 2304 2164 2306 2194
rect 2310 2193 2311 2197
rect 2315 2193 2316 2197
rect 2338 2195 2339 2199
rect 2343 2195 2344 2199
rect 2382 2199 2383 2203
rect 2387 2199 2388 2203
rect 2382 2198 2388 2199
rect 2424 2198 2426 2209
rect 2528 2198 2530 2209
rect 2338 2194 2344 2195
rect 2422 2197 2428 2198
rect 2310 2192 2316 2193
rect 2326 2170 2332 2171
rect 2326 2166 2327 2170
rect 2331 2166 2332 2170
rect 2326 2165 2332 2166
rect 2302 2163 2308 2164
rect 2302 2159 2303 2163
rect 2307 2159 2308 2163
rect 2328 2159 2330 2165
rect 2055 2158 2059 2159
rect 2074 2158 2080 2159
rect 2111 2158 2115 2159
rect 1999 2153 2003 2154
rect 2006 2155 2012 2156
rect 1542 2150 1548 2151
rect 1622 2151 1628 2152
rect 1510 2146 1516 2147
rect 1534 2146 1540 2147
rect 1366 2137 1372 2138
rect 1366 2133 1367 2137
rect 1371 2133 1372 2137
rect 1287 2132 1291 2133
rect 1366 2132 1372 2133
rect 1150 2127 1156 2128
rect 1054 2122 1060 2123
rect 1090 2123 1096 2124
rect 898 2118 904 2119
rect 960 2103 962 2122
rect 1056 2103 1058 2122
rect 1090 2119 1091 2123
rect 1095 2119 1096 2123
rect 1150 2123 1151 2127
rect 1155 2123 1156 2127
rect 1150 2122 1156 2123
rect 1254 2127 1260 2128
rect 1287 2127 1291 2128
rect 1326 2128 1332 2129
rect 1512 2128 1514 2146
rect 1534 2142 1535 2146
rect 1539 2142 1540 2146
rect 1534 2141 1540 2142
rect 1254 2123 1255 2127
rect 1259 2123 1260 2127
rect 1288 2124 1290 2127
rect 1326 2124 1327 2128
rect 1331 2124 1332 2128
rect 1254 2122 1260 2123
rect 1286 2123 1292 2124
rect 1326 2123 1332 2124
rect 1510 2127 1516 2128
rect 1510 2123 1511 2127
rect 1515 2123 1516 2127
rect 1090 2118 1096 2119
rect 1152 2103 1154 2122
rect 1256 2103 1258 2122
rect 1286 2119 1287 2123
rect 1291 2119 1292 2123
rect 1286 2118 1292 2119
rect 1328 2103 1330 2123
rect 1510 2122 1516 2123
rect 1366 2120 1372 2121
rect 1366 2116 1367 2120
rect 1371 2116 1372 2120
rect 1366 2115 1372 2116
rect 1518 2119 1524 2120
rect 1518 2115 1519 2119
rect 1523 2115 1524 2119
rect 1544 2116 1546 2150
rect 1622 2147 1623 2151
rect 1627 2147 1628 2151
rect 1632 2147 1634 2153
rect 1682 2151 1688 2152
rect 1682 2147 1683 2151
rect 1687 2147 1688 2151
rect 1736 2147 1738 2153
rect 1814 2151 1820 2152
rect 1814 2147 1815 2151
rect 1819 2147 1820 2151
rect 1840 2147 1842 2153
rect 1952 2147 1954 2153
rect 2006 2151 2007 2155
rect 2011 2151 2012 2155
rect 2055 2153 2059 2154
rect 2006 2150 2012 2151
rect 2046 2151 2052 2152
rect 2046 2147 2047 2151
rect 2051 2147 2052 2151
rect 2056 2147 2058 2153
rect 1622 2146 1628 2147
rect 1630 2146 1636 2147
rect 1682 2146 1688 2147
rect 1734 2146 1740 2147
rect 1814 2146 1820 2147
rect 1838 2146 1844 2147
rect 1614 2119 1620 2120
rect 1368 2103 1370 2115
rect 1518 2114 1524 2115
rect 1542 2115 1548 2116
rect 1520 2103 1522 2114
rect 1542 2111 1543 2115
rect 1547 2111 1548 2115
rect 1614 2115 1615 2119
rect 1619 2115 1620 2119
rect 1614 2114 1620 2115
rect 1542 2110 1548 2111
rect 1616 2103 1618 2114
rect 1624 2108 1626 2146
rect 1630 2142 1631 2146
rect 1635 2142 1636 2146
rect 1630 2141 1636 2142
rect 1622 2107 1628 2108
rect 1622 2103 1623 2107
rect 1627 2103 1628 2107
rect 759 2102 763 2103
rect 759 2097 763 2098
rect 815 2102 819 2103
rect 815 2097 819 2098
rect 863 2102 867 2103
rect 863 2097 867 2098
rect 887 2102 891 2103
rect 887 2097 891 2098
rect 959 2102 963 2103
rect 959 2097 963 2098
rect 967 2102 971 2103
rect 967 2097 971 2098
rect 1047 2102 1051 2103
rect 1047 2097 1051 2098
rect 1055 2102 1059 2103
rect 1055 2097 1059 2098
rect 1127 2102 1131 2103
rect 1127 2097 1131 2098
rect 1151 2102 1155 2103
rect 1151 2097 1155 2098
rect 1255 2102 1259 2103
rect 1255 2097 1259 2098
rect 1327 2102 1331 2103
rect 1327 2097 1331 2098
rect 1367 2102 1371 2103
rect 1367 2097 1371 2098
rect 1431 2102 1435 2103
rect 1431 2097 1435 2098
rect 1519 2102 1523 2103
rect 1519 2097 1523 2098
rect 1535 2102 1539 2103
rect 1535 2097 1539 2098
rect 1615 2102 1619 2103
rect 1622 2102 1628 2103
rect 1647 2102 1651 2103
rect 1615 2097 1619 2098
rect 1647 2097 1651 2098
rect 750 2095 756 2096
rect 750 2091 751 2095
rect 755 2091 756 2095
rect 750 2090 756 2091
rect 806 2087 812 2088
rect 678 2082 684 2083
rect 734 2085 740 2086
rect 671 2076 675 2077
rect 671 2071 675 2072
rect 670 2058 676 2059
rect 670 2054 671 2058
rect 675 2054 676 2058
rect 670 2053 676 2054
rect 646 2051 652 2052
rect 646 2047 647 2051
rect 651 2047 652 2051
rect 646 2046 652 2047
rect 672 2039 674 2053
rect 680 2040 682 2082
rect 734 2081 735 2085
rect 739 2081 740 2085
rect 806 2083 807 2087
rect 811 2083 812 2087
rect 816 2086 818 2097
rect 878 2087 884 2088
rect 806 2082 812 2083
rect 814 2085 820 2086
rect 734 2080 740 2081
rect 750 2058 756 2059
rect 750 2054 751 2058
rect 755 2054 756 2058
rect 750 2053 756 2054
rect 678 2039 684 2040
rect 752 2039 754 2053
rect 808 2052 810 2082
rect 814 2081 815 2085
rect 819 2081 820 2085
rect 878 2083 879 2087
rect 883 2083 884 2087
rect 888 2086 890 2097
rect 958 2087 964 2088
rect 878 2082 884 2083
rect 886 2085 892 2086
rect 814 2080 820 2081
rect 830 2058 836 2059
rect 830 2054 831 2058
rect 835 2054 836 2058
rect 830 2053 836 2054
rect 806 2051 812 2052
rect 806 2047 807 2051
rect 811 2047 812 2051
rect 806 2046 812 2047
rect 832 2039 834 2053
rect 880 2052 882 2082
rect 886 2081 887 2085
rect 891 2081 892 2085
rect 958 2083 959 2087
rect 963 2083 964 2087
rect 968 2086 970 2097
rect 1038 2087 1044 2088
rect 958 2082 964 2083
rect 966 2085 972 2086
rect 886 2080 892 2081
rect 902 2058 908 2059
rect 902 2054 903 2058
rect 907 2054 908 2058
rect 902 2053 908 2054
rect 878 2051 884 2052
rect 878 2047 879 2051
rect 883 2047 884 2051
rect 878 2046 884 2047
rect 904 2039 906 2053
rect 960 2052 962 2082
rect 966 2081 967 2085
rect 971 2081 972 2085
rect 1038 2083 1039 2087
rect 1043 2083 1044 2087
rect 1048 2086 1050 2097
rect 1118 2087 1124 2088
rect 1038 2082 1044 2083
rect 1046 2085 1052 2086
rect 966 2080 972 2081
rect 982 2058 988 2059
rect 982 2054 983 2058
rect 987 2054 988 2058
rect 982 2053 988 2054
rect 958 2051 964 2052
rect 958 2047 959 2051
rect 963 2047 964 2051
rect 958 2046 964 2047
rect 984 2039 986 2053
rect 1040 2052 1042 2082
rect 1046 2081 1047 2085
rect 1051 2081 1052 2085
rect 1118 2083 1119 2087
rect 1123 2083 1124 2087
rect 1128 2086 1130 2097
rect 1118 2082 1124 2083
rect 1126 2085 1132 2086
rect 1328 2085 1330 2097
rect 1368 2085 1370 2097
rect 1432 2086 1434 2097
rect 1526 2087 1532 2088
rect 1430 2085 1436 2086
rect 1046 2080 1052 2081
rect 1062 2058 1068 2059
rect 1062 2054 1063 2058
rect 1067 2054 1068 2058
rect 1062 2053 1068 2054
rect 1038 2051 1044 2052
rect 1038 2047 1039 2051
rect 1043 2047 1044 2051
rect 1038 2046 1044 2047
rect 1046 2043 1052 2044
rect 1046 2039 1047 2043
rect 1051 2039 1052 2043
rect 1064 2039 1066 2053
rect 1120 2052 1122 2082
rect 1126 2081 1127 2085
rect 1131 2081 1132 2085
rect 1126 2080 1132 2081
rect 1326 2084 1332 2085
rect 1326 2080 1327 2084
rect 1331 2080 1332 2084
rect 1326 2079 1332 2080
rect 1366 2084 1372 2085
rect 1366 2080 1367 2084
rect 1371 2080 1372 2084
rect 1430 2081 1431 2085
rect 1435 2081 1436 2085
rect 1526 2083 1527 2087
rect 1531 2083 1532 2087
rect 1536 2086 1538 2097
rect 1638 2087 1644 2088
rect 1526 2082 1532 2083
rect 1534 2085 1540 2086
rect 1430 2080 1436 2081
rect 1366 2079 1372 2080
rect 1326 2067 1332 2068
rect 1326 2063 1327 2067
rect 1331 2063 1332 2067
rect 1326 2062 1332 2063
rect 1366 2067 1372 2068
rect 1366 2063 1367 2067
rect 1371 2063 1372 2067
rect 1366 2062 1372 2063
rect 1142 2058 1148 2059
rect 1142 2054 1143 2058
rect 1147 2054 1148 2058
rect 1142 2053 1148 2054
rect 1118 2051 1124 2052
rect 1118 2047 1119 2051
rect 1123 2047 1124 2051
rect 1118 2046 1124 2047
rect 1144 2039 1146 2053
rect 1328 2039 1330 2062
rect 1368 2047 1370 2062
rect 1446 2058 1452 2059
rect 1446 2054 1447 2058
rect 1451 2054 1452 2058
rect 1446 2053 1452 2054
rect 1426 2051 1432 2052
rect 1426 2047 1427 2051
rect 1431 2047 1432 2051
rect 1448 2047 1450 2053
rect 1528 2052 1530 2082
rect 1534 2081 1535 2085
rect 1539 2081 1540 2085
rect 1638 2083 1639 2087
rect 1643 2083 1644 2087
rect 1648 2086 1650 2097
rect 1684 2088 1686 2146
rect 1734 2142 1735 2146
rect 1739 2142 1740 2146
rect 1734 2141 1740 2142
rect 1816 2128 1818 2146
rect 1838 2142 1839 2146
rect 1843 2142 1844 2146
rect 1838 2141 1844 2142
rect 1950 2146 1956 2147
rect 2046 2146 2052 2147
rect 2054 2146 2060 2147
rect 1950 2142 1951 2146
rect 1955 2142 1956 2146
rect 1950 2141 1956 2142
rect 1814 2127 1820 2128
rect 1814 2123 1815 2127
rect 1819 2123 1820 2127
rect 1814 2122 1820 2123
rect 1718 2119 1724 2120
rect 1718 2115 1719 2119
rect 1723 2115 1724 2119
rect 1718 2114 1724 2115
rect 1822 2119 1828 2120
rect 1822 2115 1823 2119
rect 1827 2115 1828 2119
rect 1934 2119 1940 2120
rect 1822 2114 1828 2115
rect 1854 2115 1860 2116
rect 1720 2103 1722 2114
rect 1824 2103 1826 2114
rect 1854 2111 1855 2115
rect 1859 2111 1860 2115
rect 1934 2115 1935 2119
rect 1939 2115 1940 2119
rect 1934 2114 1940 2115
rect 2038 2119 2044 2120
rect 2038 2115 2039 2119
rect 2043 2115 2044 2119
rect 2038 2114 2044 2115
rect 1854 2110 1860 2111
rect 1719 2102 1723 2103
rect 1719 2097 1723 2098
rect 1759 2102 1763 2103
rect 1759 2097 1763 2098
rect 1823 2102 1827 2103
rect 1823 2097 1827 2098
rect 1682 2087 1688 2088
rect 1638 2082 1644 2083
rect 1646 2085 1652 2086
rect 1534 2080 1540 2081
rect 1550 2058 1556 2059
rect 1550 2054 1551 2058
rect 1555 2054 1556 2058
rect 1550 2053 1556 2054
rect 1526 2051 1532 2052
rect 1526 2047 1527 2051
rect 1531 2047 1532 2051
rect 1552 2047 1554 2053
rect 1640 2052 1642 2082
rect 1646 2081 1647 2085
rect 1651 2081 1652 2085
rect 1682 2083 1683 2087
rect 1687 2083 1688 2087
rect 1760 2086 1762 2097
rect 1786 2087 1792 2088
rect 1682 2082 1688 2083
rect 1758 2085 1764 2086
rect 1646 2080 1652 2081
rect 1758 2081 1759 2085
rect 1763 2081 1764 2085
rect 1786 2083 1787 2087
rect 1791 2083 1792 2087
rect 1786 2082 1792 2083
rect 1758 2080 1764 2081
rect 1662 2058 1668 2059
rect 1662 2054 1663 2058
rect 1667 2054 1668 2058
rect 1662 2053 1668 2054
rect 1774 2058 1780 2059
rect 1774 2054 1775 2058
rect 1779 2054 1780 2058
rect 1774 2053 1780 2054
rect 1638 2051 1644 2052
rect 1638 2047 1639 2051
rect 1643 2047 1644 2051
rect 1664 2047 1666 2053
rect 1776 2047 1778 2053
rect 1367 2046 1371 2047
rect 1367 2041 1371 2042
rect 1415 2046 1419 2047
rect 1426 2046 1432 2047
rect 1447 2046 1451 2047
rect 1415 2041 1419 2042
rect 111 2038 115 2039
rect 111 2033 115 2034
rect 279 2038 283 2039
rect 279 2033 283 2034
rect 343 2038 347 2039
rect 343 2033 347 2034
rect 415 2038 419 2039
rect 415 2033 419 2034
rect 471 2038 475 2039
rect 471 2033 475 2034
rect 495 2038 499 2039
rect 495 2033 499 2034
rect 527 2038 531 2039
rect 527 2033 531 2034
rect 583 2038 587 2039
rect 583 2033 587 2034
rect 639 2038 643 2039
rect 639 2033 643 2034
rect 671 2038 675 2039
rect 678 2035 679 2039
rect 683 2035 684 2039
rect 678 2034 684 2035
rect 695 2038 699 2039
rect 671 2033 675 2034
rect 695 2033 699 2034
rect 751 2038 755 2039
rect 751 2033 755 2034
rect 807 2038 811 2039
rect 807 2033 811 2034
rect 831 2038 835 2039
rect 831 2033 835 2034
rect 863 2038 867 2039
rect 863 2033 867 2034
rect 903 2038 907 2039
rect 903 2033 907 2034
rect 919 2038 923 2039
rect 919 2033 923 2034
rect 975 2038 979 2039
rect 975 2033 979 2034
rect 983 2038 987 2039
rect 983 2033 987 2034
rect 1031 2038 1035 2039
rect 1046 2038 1052 2039
rect 1063 2038 1067 2039
rect 1031 2033 1035 2034
rect 112 2018 114 2033
rect 416 2027 418 2033
rect 472 2027 474 2033
rect 528 2027 530 2033
rect 546 2031 552 2032
rect 546 2027 547 2031
rect 551 2027 552 2031
rect 584 2027 586 2033
rect 602 2031 608 2032
rect 602 2027 603 2031
rect 607 2027 608 2031
rect 640 2027 642 2033
rect 658 2031 664 2032
rect 658 2027 659 2031
rect 663 2027 664 2031
rect 696 2027 698 2033
rect 742 2031 748 2032
rect 742 2027 743 2031
rect 747 2027 748 2031
rect 752 2027 754 2033
rect 808 2027 810 2033
rect 864 2027 866 2033
rect 920 2027 922 2033
rect 976 2027 978 2033
rect 1032 2027 1034 2033
rect 414 2026 420 2027
rect 414 2022 415 2026
rect 419 2022 420 2026
rect 414 2021 420 2022
rect 470 2026 476 2027
rect 470 2022 471 2026
rect 475 2022 476 2026
rect 470 2021 476 2022
rect 526 2026 532 2027
rect 546 2026 552 2027
rect 582 2026 588 2027
rect 602 2026 608 2027
rect 638 2026 644 2027
rect 658 2026 664 2027
rect 694 2026 700 2027
rect 742 2026 748 2027
rect 750 2026 756 2027
rect 526 2022 527 2026
rect 531 2022 532 2026
rect 526 2021 532 2022
rect 110 2017 116 2018
rect 110 2013 111 2017
rect 115 2013 116 2017
rect 110 2012 116 2013
rect 110 2000 116 2001
rect 110 1996 111 2000
rect 115 1996 116 2000
rect 110 1995 116 1996
rect 398 1999 404 2000
rect 398 1995 399 1999
rect 403 1995 404 1999
rect 112 1979 114 1995
rect 398 1994 404 1995
rect 454 1999 460 2000
rect 454 1995 455 1999
rect 459 1995 460 1999
rect 454 1994 460 1995
rect 510 1999 516 2000
rect 510 1995 511 1999
rect 515 1995 516 1999
rect 548 1996 550 2026
rect 582 2022 583 2026
rect 587 2022 588 2026
rect 582 2021 588 2022
rect 566 1999 572 2000
rect 510 1994 516 1995
rect 546 1995 552 1996
rect 400 1979 402 1994
rect 456 1979 458 1994
rect 512 1979 514 1994
rect 546 1991 547 1995
rect 551 1991 552 1995
rect 566 1995 567 1999
rect 571 1995 572 1999
rect 604 1996 606 2026
rect 638 2022 639 2026
rect 643 2022 644 2026
rect 638 2021 644 2022
rect 622 1999 628 2000
rect 566 1994 572 1995
rect 602 1995 608 1996
rect 546 1990 552 1991
rect 568 1979 570 1994
rect 602 1991 603 1995
rect 607 1991 608 1995
rect 622 1995 623 1999
rect 627 1995 628 1999
rect 660 1996 662 2026
rect 694 2022 695 2026
rect 699 2022 700 2026
rect 694 2021 700 2022
rect 678 1999 684 2000
rect 622 1994 628 1995
rect 658 1995 664 1996
rect 602 1990 608 1991
rect 590 1987 596 1988
rect 590 1983 591 1987
rect 595 1983 596 1987
rect 590 1982 596 1983
rect 111 1978 115 1979
rect 111 1973 115 1974
rect 335 1978 339 1979
rect 335 1973 339 1974
rect 391 1978 395 1979
rect 391 1973 395 1974
rect 399 1978 403 1979
rect 399 1973 403 1974
rect 447 1978 451 1979
rect 447 1973 451 1974
rect 455 1978 459 1979
rect 455 1973 459 1974
rect 503 1978 507 1979
rect 503 1973 507 1974
rect 511 1978 515 1979
rect 511 1973 515 1974
rect 567 1978 571 1979
rect 567 1973 571 1974
rect 112 1961 114 1973
rect 336 1962 338 1973
rect 358 1971 364 1972
rect 358 1967 359 1971
rect 363 1967 364 1971
rect 358 1966 364 1967
rect 334 1961 340 1962
rect 110 1960 116 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 334 1957 335 1961
rect 339 1957 340 1961
rect 334 1956 340 1957
rect 110 1955 116 1956
rect 110 1943 116 1944
rect 110 1939 111 1943
rect 115 1939 116 1943
rect 110 1938 116 1939
rect 112 1923 114 1938
rect 350 1934 356 1935
rect 350 1930 351 1934
rect 355 1930 356 1934
rect 350 1929 356 1930
rect 352 1923 354 1929
rect 360 1928 362 1966
rect 382 1963 388 1964
rect 382 1959 383 1963
rect 387 1959 388 1963
rect 392 1962 394 1973
rect 438 1963 444 1964
rect 382 1958 388 1959
rect 390 1961 396 1962
rect 384 1928 386 1958
rect 390 1957 391 1961
rect 395 1957 396 1961
rect 438 1959 439 1963
rect 443 1959 444 1963
rect 448 1962 450 1973
rect 494 1963 500 1964
rect 438 1958 444 1959
rect 446 1961 452 1962
rect 390 1956 396 1957
rect 406 1934 412 1935
rect 406 1930 407 1934
rect 411 1930 412 1934
rect 406 1929 412 1930
rect 358 1927 364 1928
rect 358 1923 359 1927
rect 363 1923 364 1927
rect 111 1922 115 1923
rect 111 1917 115 1918
rect 159 1922 163 1923
rect 159 1917 163 1918
rect 231 1922 235 1923
rect 231 1917 235 1918
rect 327 1922 331 1923
rect 327 1917 331 1918
rect 351 1922 355 1923
rect 358 1922 364 1923
rect 382 1927 388 1928
rect 382 1923 383 1927
rect 387 1923 388 1927
rect 408 1923 410 1929
rect 440 1928 442 1958
rect 446 1957 447 1961
rect 451 1957 452 1961
rect 494 1959 495 1963
rect 499 1959 500 1963
rect 504 1962 506 1973
rect 568 1962 570 1973
rect 494 1958 500 1959
rect 502 1961 508 1962
rect 446 1956 452 1957
rect 462 1934 468 1935
rect 462 1930 463 1934
rect 467 1930 468 1934
rect 462 1929 468 1930
rect 438 1927 444 1928
rect 438 1923 439 1927
rect 443 1923 444 1927
rect 464 1923 466 1929
rect 382 1922 388 1923
rect 407 1922 411 1923
rect 351 1917 355 1918
rect 407 1917 411 1918
rect 431 1922 435 1923
rect 438 1922 444 1923
rect 463 1922 467 1923
rect 431 1917 435 1918
rect 463 1917 467 1918
rect 112 1902 114 1917
rect 134 1915 140 1916
rect 134 1911 135 1915
rect 139 1911 140 1915
rect 160 1911 162 1917
rect 222 1915 228 1916
rect 222 1911 223 1915
rect 227 1911 228 1915
rect 232 1911 234 1917
rect 302 1915 308 1916
rect 302 1911 303 1915
rect 307 1911 308 1915
rect 328 1911 330 1917
rect 422 1915 428 1916
rect 422 1911 423 1915
rect 427 1911 428 1915
rect 432 1911 434 1917
rect 496 1916 498 1958
rect 502 1957 503 1961
rect 507 1957 508 1961
rect 502 1956 508 1957
rect 566 1961 572 1962
rect 566 1957 567 1961
rect 571 1957 572 1961
rect 566 1956 572 1957
rect 518 1934 524 1935
rect 518 1930 519 1934
rect 523 1930 524 1934
rect 518 1929 524 1930
rect 582 1934 588 1935
rect 582 1930 583 1934
rect 587 1930 588 1934
rect 582 1929 588 1930
rect 520 1923 522 1929
rect 584 1923 586 1929
rect 592 1928 594 1982
rect 624 1979 626 1994
rect 658 1991 659 1995
rect 663 1991 664 1995
rect 678 1995 679 1999
rect 683 1995 684 1999
rect 678 1994 684 1995
rect 734 1999 740 2000
rect 734 1995 735 1999
rect 739 1995 740 1999
rect 744 1997 746 2026
rect 750 2022 751 2026
rect 755 2022 756 2026
rect 750 2021 756 2022
rect 806 2026 812 2027
rect 806 2022 807 2026
rect 811 2022 812 2026
rect 806 2021 812 2022
rect 862 2026 868 2027
rect 862 2022 863 2026
rect 867 2022 868 2026
rect 862 2021 868 2022
rect 918 2026 924 2027
rect 918 2022 919 2026
rect 923 2022 924 2026
rect 918 2021 924 2022
rect 974 2026 980 2027
rect 974 2022 975 2026
rect 979 2022 980 2026
rect 974 2021 980 2022
rect 1030 2026 1036 2027
rect 1030 2022 1031 2026
rect 1035 2022 1036 2026
rect 1030 2021 1036 2022
rect 790 1999 796 2000
rect 734 1994 740 1995
rect 743 1996 747 1997
rect 658 1990 664 1991
rect 680 1979 682 1994
rect 736 1979 738 1994
rect 790 1995 791 1999
rect 795 1995 796 1999
rect 790 1994 796 1995
rect 846 1999 852 2000
rect 846 1995 847 1999
rect 851 1995 852 1999
rect 846 1994 852 1995
rect 902 1999 908 2000
rect 902 1995 903 1999
rect 907 1995 908 1999
rect 902 1994 908 1995
rect 958 1999 964 2000
rect 958 1995 959 1999
rect 963 1995 964 1999
rect 958 1994 964 1995
rect 1014 1999 1020 2000
rect 1014 1995 1015 1999
rect 1019 1995 1020 1999
rect 1048 1996 1050 2038
rect 1063 2033 1067 2034
rect 1143 2038 1147 2039
rect 1143 2033 1147 2034
rect 1327 2038 1331 2039
rect 1327 2033 1331 2034
rect 1328 2018 1330 2033
rect 1368 2026 1370 2041
rect 1390 2039 1396 2040
rect 1390 2035 1391 2039
rect 1395 2035 1396 2039
rect 1416 2035 1418 2041
rect 1390 2034 1396 2035
rect 1414 2034 1420 2035
rect 1366 2025 1372 2026
rect 1366 2021 1367 2025
rect 1371 2021 1372 2025
rect 1366 2020 1372 2021
rect 1326 2017 1332 2018
rect 1326 2013 1327 2017
rect 1331 2013 1332 2017
rect 1392 2016 1394 2034
rect 1414 2030 1415 2034
rect 1419 2030 1420 2034
rect 1414 2029 1420 2030
rect 1326 2012 1332 2013
rect 1390 2015 1396 2016
rect 1390 2011 1391 2015
rect 1395 2011 1396 2015
rect 1390 2010 1396 2011
rect 1366 2008 1372 2009
rect 1366 2004 1367 2008
rect 1371 2004 1372 2008
rect 1366 2003 1372 2004
rect 1398 2007 1404 2008
rect 1398 2003 1399 2007
rect 1403 2003 1404 2007
rect 1428 2004 1430 2046
rect 1447 2041 1451 2042
rect 1503 2046 1507 2047
rect 1526 2046 1532 2047
rect 1551 2046 1555 2047
rect 1503 2041 1507 2042
rect 1551 2041 1555 2042
rect 1607 2046 1611 2047
rect 1638 2046 1644 2047
rect 1663 2046 1667 2047
rect 1607 2041 1611 2042
rect 1663 2041 1667 2042
rect 1711 2046 1715 2047
rect 1711 2041 1715 2042
rect 1775 2046 1779 2047
rect 1775 2041 1779 2042
rect 1494 2039 1500 2040
rect 1494 2035 1495 2039
rect 1499 2035 1500 2039
rect 1504 2035 1506 2041
rect 1522 2039 1528 2040
rect 1522 2035 1523 2039
rect 1527 2035 1528 2039
rect 1608 2035 1610 2041
rect 1686 2039 1692 2040
rect 1686 2035 1687 2039
rect 1691 2035 1692 2039
rect 1712 2035 1714 2041
rect 1788 2040 1790 2082
rect 1856 2052 1858 2110
rect 1936 2103 1938 2114
rect 2040 2103 2042 2114
rect 2048 2108 2050 2146
rect 2054 2142 2055 2146
rect 2059 2142 2060 2146
rect 2054 2141 2060 2142
rect 2076 2116 2078 2158
rect 2111 2153 2115 2154
rect 2159 2158 2163 2159
rect 2198 2158 2204 2159
rect 2223 2158 2227 2159
rect 2159 2153 2163 2154
rect 2223 2153 2227 2154
rect 2263 2158 2267 2159
rect 2302 2158 2308 2159
rect 2327 2158 2331 2159
rect 2263 2153 2267 2154
rect 2294 2155 2300 2156
rect 2134 2151 2140 2152
rect 2134 2147 2135 2151
rect 2139 2147 2140 2151
rect 2160 2147 2162 2153
rect 2264 2147 2266 2153
rect 2294 2151 2295 2155
rect 2299 2151 2300 2155
rect 2327 2153 2331 2154
rect 2340 2152 2342 2194
rect 2422 2193 2423 2197
rect 2427 2193 2428 2197
rect 2422 2192 2428 2193
rect 2526 2197 2532 2198
rect 2584 2197 2586 2209
rect 2526 2193 2527 2197
rect 2531 2193 2532 2197
rect 2526 2192 2532 2193
rect 2582 2196 2588 2197
rect 2582 2192 2583 2196
rect 2587 2192 2588 2196
rect 2582 2191 2588 2192
rect 2582 2179 2588 2180
rect 2582 2175 2583 2179
rect 2587 2175 2588 2179
rect 2582 2174 2588 2175
rect 2438 2170 2444 2171
rect 2438 2166 2439 2170
rect 2443 2166 2444 2170
rect 2438 2165 2444 2166
rect 2542 2170 2548 2171
rect 2542 2166 2543 2170
rect 2547 2166 2548 2170
rect 2542 2165 2548 2166
rect 2440 2159 2442 2165
rect 2544 2159 2546 2165
rect 2558 2163 2564 2164
rect 2558 2159 2559 2163
rect 2563 2159 2564 2163
rect 2584 2159 2586 2174
rect 2359 2158 2363 2159
rect 2359 2153 2363 2154
rect 2439 2158 2443 2159
rect 2439 2153 2443 2154
rect 2463 2158 2467 2159
rect 2463 2153 2467 2154
rect 2543 2158 2547 2159
rect 2558 2158 2564 2159
rect 2583 2158 2587 2159
rect 2543 2153 2547 2154
rect 2294 2150 2300 2151
rect 2338 2151 2344 2152
rect 2134 2146 2140 2147
rect 2158 2146 2164 2147
rect 2136 2128 2138 2146
rect 2158 2142 2159 2146
rect 2163 2142 2164 2146
rect 2158 2141 2164 2142
rect 2262 2146 2268 2147
rect 2262 2142 2263 2146
rect 2267 2142 2268 2146
rect 2262 2141 2268 2142
rect 2134 2127 2140 2128
rect 2134 2123 2135 2127
rect 2139 2123 2140 2127
rect 2134 2122 2140 2123
rect 2142 2119 2148 2120
rect 2074 2115 2080 2116
rect 2074 2111 2075 2115
rect 2079 2111 2080 2115
rect 2142 2115 2143 2119
rect 2147 2115 2148 2119
rect 2142 2114 2148 2115
rect 2246 2119 2252 2120
rect 2246 2115 2247 2119
rect 2251 2115 2252 2119
rect 2246 2114 2252 2115
rect 2074 2110 2080 2111
rect 2046 2107 2052 2108
rect 2046 2103 2047 2107
rect 2051 2103 2052 2107
rect 2144 2103 2146 2114
rect 2248 2103 2250 2114
rect 1863 2102 1867 2103
rect 1863 2097 1867 2098
rect 1935 2102 1939 2103
rect 1935 2097 1939 2098
rect 1967 2102 1971 2103
rect 1967 2097 1971 2098
rect 2039 2102 2043 2103
rect 2046 2102 2052 2103
rect 2071 2102 2075 2103
rect 2039 2097 2043 2098
rect 2071 2097 2075 2098
rect 2143 2102 2147 2103
rect 2143 2097 2147 2098
rect 2175 2102 2179 2103
rect 2175 2097 2179 2098
rect 2247 2102 2251 2103
rect 2247 2097 2251 2098
rect 2271 2102 2275 2103
rect 2271 2097 2275 2098
rect 1864 2086 1866 2097
rect 1968 2086 1970 2097
rect 2062 2087 2068 2088
rect 1862 2085 1868 2086
rect 1862 2081 1863 2085
rect 1867 2081 1868 2085
rect 1862 2080 1868 2081
rect 1966 2085 1972 2086
rect 1966 2081 1967 2085
rect 1971 2081 1972 2085
rect 2062 2083 2063 2087
rect 2067 2083 2068 2087
rect 2072 2086 2074 2097
rect 2166 2087 2172 2088
rect 2062 2082 2068 2083
rect 2070 2085 2076 2086
rect 1966 2080 1972 2081
rect 1878 2058 1884 2059
rect 1878 2054 1879 2058
rect 1883 2054 1884 2058
rect 1878 2053 1884 2054
rect 1982 2058 1988 2059
rect 1982 2054 1983 2058
rect 1987 2054 1988 2058
rect 1982 2053 1988 2054
rect 1854 2051 1860 2052
rect 1854 2047 1855 2051
rect 1859 2047 1860 2051
rect 1880 2047 1882 2053
rect 1984 2047 1986 2053
rect 2064 2052 2066 2082
rect 2070 2081 2071 2085
rect 2075 2081 2076 2085
rect 2166 2083 2167 2087
rect 2171 2083 2172 2087
rect 2176 2086 2178 2097
rect 2262 2087 2268 2088
rect 2166 2082 2172 2083
rect 2174 2085 2180 2086
rect 2070 2080 2076 2081
rect 2086 2058 2092 2059
rect 2086 2054 2087 2058
rect 2091 2054 2092 2058
rect 2086 2053 2092 2054
rect 2054 2051 2060 2052
rect 2054 2047 2055 2051
rect 2059 2047 2060 2051
rect 1807 2046 1811 2047
rect 1854 2046 1860 2047
rect 1879 2046 1883 2047
rect 1807 2041 1811 2042
rect 1879 2041 1883 2042
rect 1903 2046 1907 2047
rect 1903 2041 1907 2042
rect 1983 2046 1987 2047
rect 1983 2041 1987 2042
rect 2007 2046 2011 2047
rect 2054 2046 2060 2047
rect 2062 2051 2068 2052
rect 2062 2047 2063 2051
rect 2067 2047 2068 2051
rect 2088 2047 2090 2053
rect 2168 2052 2170 2082
rect 2174 2081 2175 2085
rect 2179 2081 2180 2085
rect 2262 2083 2263 2087
rect 2267 2083 2268 2087
rect 2272 2086 2274 2097
rect 2296 2088 2298 2150
rect 2338 2147 2339 2151
rect 2343 2147 2344 2151
rect 2360 2147 2362 2153
rect 2464 2147 2466 2153
rect 2534 2151 2540 2152
rect 2534 2147 2535 2151
rect 2539 2147 2540 2151
rect 2544 2147 2546 2153
rect 2338 2146 2344 2147
rect 2358 2146 2364 2147
rect 2358 2142 2359 2146
rect 2363 2142 2364 2146
rect 2358 2141 2364 2142
rect 2462 2146 2468 2147
rect 2534 2146 2540 2147
rect 2542 2146 2548 2147
rect 2462 2142 2463 2146
rect 2467 2142 2468 2146
rect 2462 2141 2468 2142
rect 2342 2119 2348 2120
rect 2342 2115 2343 2119
rect 2347 2115 2348 2119
rect 2342 2114 2348 2115
rect 2446 2119 2452 2120
rect 2446 2115 2447 2119
rect 2451 2115 2452 2119
rect 2526 2119 2532 2120
rect 2446 2114 2452 2115
rect 2478 2115 2484 2116
rect 2344 2103 2346 2114
rect 2448 2103 2450 2114
rect 2478 2111 2479 2115
rect 2483 2111 2484 2115
rect 2526 2115 2527 2119
rect 2531 2115 2532 2119
rect 2526 2114 2532 2115
rect 2478 2110 2484 2111
rect 2343 2102 2347 2103
rect 2343 2097 2347 2098
rect 2359 2102 2363 2103
rect 2359 2097 2363 2098
rect 2447 2102 2451 2103
rect 2447 2097 2451 2098
rect 2455 2102 2459 2103
rect 2455 2097 2459 2098
rect 2294 2087 2300 2088
rect 2262 2082 2268 2083
rect 2270 2085 2276 2086
rect 2174 2080 2180 2081
rect 2190 2058 2196 2059
rect 2190 2054 2191 2058
rect 2195 2054 2196 2058
rect 2190 2053 2196 2054
rect 2166 2051 2172 2052
rect 2166 2047 2167 2051
rect 2171 2047 2172 2051
rect 2192 2047 2194 2053
rect 2264 2052 2266 2082
rect 2270 2081 2271 2085
rect 2275 2081 2276 2085
rect 2294 2083 2295 2087
rect 2299 2083 2300 2087
rect 2360 2086 2362 2097
rect 2430 2091 2436 2092
rect 2422 2087 2428 2088
rect 2294 2082 2300 2083
rect 2358 2085 2364 2086
rect 2270 2080 2276 2081
rect 2358 2081 2359 2085
rect 2363 2081 2364 2085
rect 2422 2083 2423 2087
rect 2427 2083 2428 2087
rect 2430 2087 2431 2091
rect 2435 2087 2436 2091
rect 2430 2086 2436 2087
rect 2456 2086 2458 2097
rect 2422 2082 2428 2083
rect 2358 2080 2364 2081
rect 2286 2058 2292 2059
rect 2286 2054 2287 2058
rect 2291 2054 2292 2058
rect 2286 2053 2292 2054
rect 2374 2058 2380 2059
rect 2374 2054 2375 2058
rect 2379 2054 2380 2058
rect 2374 2053 2380 2054
rect 2262 2051 2268 2052
rect 2262 2047 2263 2051
rect 2267 2047 2268 2051
rect 2288 2047 2290 2053
rect 2376 2047 2378 2053
rect 2062 2046 2068 2047
rect 2087 2046 2091 2047
rect 2007 2041 2011 2042
rect 1786 2039 1792 2040
rect 1786 2035 1787 2039
rect 1791 2035 1792 2039
rect 1808 2035 1810 2041
rect 1894 2039 1900 2040
rect 1894 2035 1895 2039
rect 1899 2035 1900 2039
rect 1904 2035 1906 2041
rect 1918 2039 1924 2040
rect 1918 2035 1919 2039
rect 1923 2035 1924 2039
rect 2008 2035 2010 2041
rect 1494 2034 1500 2035
rect 1502 2034 1508 2035
rect 1522 2034 1528 2035
rect 1606 2034 1612 2035
rect 1686 2034 1692 2035
rect 1710 2034 1716 2035
rect 1786 2034 1792 2035
rect 1806 2034 1812 2035
rect 1894 2034 1900 2035
rect 1902 2034 1908 2035
rect 1918 2034 1924 2035
rect 2006 2034 2012 2035
rect 1486 2007 1492 2008
rect 1326 2000 1332 2001
rect 1175 1996 1179 1997
rect 1014 1994 1020 1995
rect 1046 1995 1052 1996
rect 743 1991 747 1992
rect 792 1979 794 1994
rect 848 1979 850 1994
rect 904 1979 906 1994
rect 960 1979 962 1994
rect 1016 1979 1018 1994
rect 1046 1991 1047 1995
rect 1051 1991 1052 1995
rect 1326 1996 1327 2000
rect 1331 1996 1332 2000
rect 1326 1995 1332 1996
rect 1175 1991 1179 1992
rect 1046 1990 1052 1991
rect 623 1978 627 1979
rect 623 1973 627 1974
rect 647 1978 651 1979
rect 647 1973 651 1974
rect 679 1978 683 1979
rect 679 1973 683 1974
rect 735 1978 739 1979
rect 735 1973 739 1974
rect 743 1978 747 1979
rect 743 1973 747 1974
rect 791 1978 795 1979
rect 791 1973 795 1974
rect 847 1978 851 1979
rect 847 1973 851 1974
rect 863 1978 867 1979
rect 863 1973 867 1974
rect 903 1978 907 1979
rect 903 1973 907 1974
rect 959 1978 963 1979
rect 959 1973 963 1974
rect 999 1978 1003 1979
rect 999 1973 1003 1974
rect 1015 1978 1019 1979
rect 1015 1973 1019 1974
rect 1143 1978 1147 1979
rect 1143 1973 1147 1974
rect 648 1962 650 1973
rect 734 1963 740 1964
rect 646 1961 652 1962
rect 646 1957 647 1961
rect 651 1957 652 1961
rect 734 1959 735 1963
rect 739 1959 740 1963
rect 744 1962 746 1973
rect 854 1963 860 1964
rect 734 1958 740 1959
rect 742 1961 748 1962
rect 646 1956 652 1957
rect 662 1934 668 1935
rect 662 1930 663 1934
rect 667 1930 668 1934
rect 662 1929 668 1930
rect 590 1927 596 1928
rect 590 1923 591 1927
rect 595 1923 596 1927
rect 664 1923 666 1929
rect 736 1928 738 1958
rect 742 1957 743 1961
rect 747 1957 748 1961
rect 854 1959 855 1963
rect 859 1959 860 1963
rect 864 1962 866 1973
rect 990 1963 996 1964
rect 854 1958 860 1959
rect 862 1961 868 1962
rect 742 1956 748 1957
rect 758 1934 764 1935
rect 758 1930 759 1934
rect 763 1930 764 1934
rect 758 1929 764 1930
rect 670 1927 676 1928
rect 670 1923 671 1927
rect 675 1923 676 1927
rect 519 1922 523 1923
rect 519 1917 523 1918
rect 543 1922 547 1923
rect 543 1917 547 1918
rect 583 1922 587 1923
rect 590 1922 596 1923
rect 655 1922 659 1923
rect 583 1917 587 1918
rect 655 1917 659 1918
rect 663 1922 667 1923
rect 670 1922 676 1923
rect 734 1927 740 1928
rect 734 1923 735 1927
rect 739 1923 740 1927
rect 760 1923 762 1929
rect 856 1928 858 1958
rect 862 1957 863 1961
rect 867 1957 868 1961
rect 990 1959 991 1963
rect 995 1959 996 1963
rect 1000 1962 1002 1973
rect 1134 1963 1140 1964
rect 990 1958 996 1959
rect 998 1961 1004 1962
rect 862 1956 868 1957
rect 878 1934 884 1935
rect 878 1930 879 1934
rect 883 1930 884 1934
rect 878 1929 884 1930
rect 854 1927 860 1928
rect 854 1923 855 1927
rect 859 1923 860 1927
rect 880 1923 882 1929
rect 992 1928 994 1958
rect 998 1957 999 1961
rect 1003 1957 1004 1961
rect 1134 1959 1135 1963
rect 1139 1959 1140 1963
rect 1144 1962 1146 1973
rect 1176 1964 1178 1991
rect 1328 1979 1330 1995
rect 1368 1991 1370 2003
rect 1398 2002 1404 2003
rect 1426 2003 1432 2004
rect 1400 1991 1402 2002
rect 1426 1999 1427 2003
rect 1431 1999 1432 2003
rect 1486 2003 1487 2007
rect 1491 2003 1492 2007
rect 1486 2002 1492 2003
rect 1426 1998 1432 1999
rect 1488 1991 1490 2002
rect 1367 1990 1371 1991
rect 1367 1985 1371 1986
rect 1399 1990 1403 1991
rect 1399 1985 1403 1986
rect 1479 1990 1483 1991
rect 1479 1985 1483 1986
rect 1487 1990 1491 1991
rect 1487 1985 1491 1986
rect 1271 1978 1275 1979
rect 1271 1973 1275 1974
rect 1327 1978 1331 1979
rect 1327 1973 1331 1974
rect 1368 1973 1370 1985
rect 1400 1974 1402 1985
rect 1470 1975 1476 1976
rect 1398 1973 1404 1974
rect 1174 1963 1180 1964
rect 1134 1958 1140 1959
rect 1142 1961 1148 1962
rect 998 1956 1004 1957
rect 1014 1934 1020 1935
rect 1014 1930 1015 1934
rect 1019 1930 1020 1934
rect 1014 1929 1020 1930
rect 990 1927 996 1928
rect 990 1923 991 1927
rect 995 1923 996 1927
rect 1016 1923 1018 1929
rect 1136 1928 1138 1958
rect 1142 1957 1143 1961
rect 1147 1957 1148 1961
rect 1174 1959 1175 1963
rect 1179 1959 1180 1963
rect 1272 1962 1274 1973
rect 1174 1958 1180 1959
rect 1270 1961 1276 1962
rect 1328 1961 1330 1973
rect 1366 1972 1372 1973
rect 1366 1968 1367 1972
rect 1371 1968 1372 1972
rect 1398 1969 1399 1973
rect 1403 1969 1404 1973
rect 1470 1971 1471 1975
rect 1475 1971 1476 1975
rect 1480 1974 1482 1985
rect 1496 1980 1498 2034
rect 1502 2030 1503 2034
rect 1507 2030 1508 2034
rect 1502 2029 1508 2030
rect 1524 2004 1526 2034
rect 1606 2030 1607 2034
rect 1611 2030 1612 2034
rect 1606 2029 1612 2030
rect 1688 2016 1690 2034
rect 1710 2030 1711 2034
rect 1715 2030 1716 2034
rect 1710 2029 1716 2030
rect 1806 2030 1807 2034
rect 1811 2030 1812 2034
rect 1806 2029 1812 2030
rect 1686 2015 1692 2016
rect 1686 2011 1687 2015
rect 1691 2011 1692 2015
rect 1686 2010 1692 2011
rect 1590 2007 1596 2008
rect 1522 2003 1528 2004
rect 1522 1999 1523 2003
rect 1527 1999 1528 2003
rect 1590 2003 1591 2007
rect 1595 2003 1596 2007
rect 1590 2002 1596 2003
rect 1694 2007 1700 2008
rect 1694 2003 1695 2007
rect 1699 2003 1700 2007
rect 1790 2007 1796 2008
rect 1694 2002 1700 2003
rect 1758 2003 1764 2004
rect 1522 1998 1528 1999
rect 1592 1991 1594 2002
rect 1696 1991 1698 2002
rect 1758 1999 1759 2003
rect 1763 1999 1764 2003
rect 1790 2003 1791 2007
rect 1795 2003 1796 2007
rect 1790 2002 1796 2003
rect 1886 2007 1892 2008
rect 1886 2003 1887 2007
rect 1891 2003 1892 2007
rect 1886 2002 1892 2003
rect 1758 1998 1764 1999
rect 1583 1990 1587 1991
rect 1583 1985 1587 1986
rect 1591 1990 1595 1991
rect 1591 1985 1595 1986
rect 1679 1990 1683 1991
rect 1679 1985 1683 1986
rect 1695 1990 1699 1991
rect 1695 1985 1699 1986
rect 1494 1979 1500 1980
rect 1494 1975 1495 1979
rect 1499 1975 1500 1979
rect 1494 1974 1500 1975
rect 1584 1974 1586 1985
rect 1606 1983 1612 1984
rect 1606 1979 1607 1983
rect 1611 1979 1612 1983
rect 1606 1978 1612 1979
rect 1470 1970 1476 1971
rect 1478 1973 1484 1974
rect 1398 1968 1404 1969
rect 1366 1967 1372 1968
rect 1142 1956 1148 1957
rect 1270 1957 1271 1961
rect 1275 1957 1276 1961
rect 1270 1956 1276 1957
rect 1326 1960 1332 1961
rect 1326 1956 1327 1960
rect 1331 1956 1332 1960
rect 1326 1955 1332 1956
rect 1366 1955 1372 1956
rect 1366 1951 1367 1955
rect 1371 1951 1372 1955
rect 1366 1950 1372 1951
rect 1326 1943 1332 1944
rect 1326 1939 1327 1943
rect 1331 1939 1332 1943
rect 1326 1938 1332 1939
rect 1158 1934 1164 1935
rect 1158 1930 1159 1934
rect 1163 1930 1164 1934
rect 1158 1929 1164 1930
rect 1286 1934 1292 1935
rect 1286 1930 1287 1934
rect 1291 1930 1292 1934
rect 1286 1929 1292 1930
rect 1134 1927 1140 1928
rect 1134 1923 1135 1927
rect 1139 1923 1140 1927
rect 1160 1923 1162 1929
rect 1218 1927 1224 1928
rect 1218 1923 1219 1927
rect 1223 1923 1224 1927
rect 1288 1923 1290 1929
rect 1328 1923 1330 1938
rect 1368 1931 1370 1950
rect 1414 1946 1420 1947
rect 1414 1942 1415 1946
rect 1419 1942 1420 1946
rect 1414 1941 1420 1942
rect 1416 1931 1418 1941
rect 1472 1940 1474 1970
rect 1478 1969 1479 1973
rect 1483 1969 1484 1973
rect 1478 1968 1484 1969
rect 1582 1973 1588 1974
rect 1582 1969 1583 1973
rect 1587 1969 1588 1973
rect 1582 1968 1588 1969
rect 1494 1946 1500 1947
rect 1494 1942 1495 1946
rect 1499 1942 1500 1946
rect 1494 1941 1500 1942
rect 1598 1946 1604 1947
rect 1598 1942 1599 1946
rect 1603 1942 1604 1946
rect 1598 1941 1604 1942
rect 1470 1939 1476 1940
rect 1470 1935 1471 1939
rect 1475 1935 1476 1939
rect 1470 1934 1476 1935
rect 1496 1931 1498 1941
rect 1600 1931 1602 1941
rect 1608 1940 1610 1978
rect 1670 1975 1676 1976
rect 1670 1971 1671 1975
rect 1675 1971 1676 1975
rect 1680 1974 1682 1985
rect 1706 1975 1712 1976
rect 1670 1970 1676 1971
rect 1678 1973 1684 1974
rect 1672 1940 1674 1970
rect 1678 1969 1679 1973
rect 1683 1969 1684 1973
rect 1706 1971 1707 1975
rect 1711 1971 1712 1975
rect 1706 1970 1712 1971
rect 1678 1968 1684 1969
rect 1694 1946 1700 1947
rect 1694 1942 1695 1946
rect 1699 1942 1700 1946
rect 1694 1941 1700 1942
rect 1606 1939 1612 1940
rect 1606 1935 1607 1939
rect 1611 1935 1612 1939
rect 1606 1934 1612 1935
rect 1670 1939 1676 1940
rect 1670 1935 1671 1939
rect 1675 1935 1676 1939
rect 1670 1934 1676 1935
rect 1696 1931 1698 1941
rect 1367 1930 1371 1931
rect 1367 1925 1371 1926
rect 1415 1930 1419 1931
rect 1415 1925 1419 1926
rect 1495 1930 1499 1931
rect 1495 1925 1499 1926
rect 1599 1930 1603 1931
rect 1599 1925 1603 1926
rect 1695 1930 1699 1931
rect 1708 1928 1710 1970
rect 1760 1940 1762 1998
rect 1792 1991 1794 2002
rect 1888 1991 1890 2002
rect 1767 1990 1771 1991
rect 1767 1985 1771 1986
rect 1791 1990 1795 1991
rect 1791 1985 1795 1986
rect 1847 1990 1851 1991
rect 1847 1985 1851 1986
rect 1887 1990 1891 1991
rect 1887 1985 1891 1986
rect 1768 1974 1770 1985
rect 1848 1974 1850 1985
rect 1896 1984 1898 2034
rect 1902 2030 1903 2034
rect 1907 2030 1908 2034
rect 1902 2029 1908 2030
rect 1920 2004 1922 2034
rect 2006 2030 2007 2034
rect 2011 2030 2012 2034
rect 2006 2029 2012 2030
rect 2056 2016 2058 2046
rect 2087 2041 2091 2042
rect 2111 2046 2115 2047
rect 2166 2046 2172 2047
rect 2191 2046 2195 2047
rect 2111 2041 2115 2042
rect 2191 2041 2195 2042
rect 2215 2046 2219 2047
rect 2262 2046 2268 2047
rect 2287 2046 2291 2047
rect 2215 2041 2219 2042
rect 2287 2041 2291 2042
rect 2327 2046 2331 2047
rect 2327 2041 2331 2042
rect 2375 2046 2379 2047
rect 2375 2041 2379 2042
rect 2112 2035 2114 2041
rect 2130 2039 2136 2040
rect 2130 2035 2131 2039
rect 2135 2035 2136 2039
rect 2216 2035 2218 2041
rect 2234 2039 2240 2040
rect 2234 2035 2235 2039
rect 2239 2035 2240 2039
rect 2328 2035 2330 2041
rect 2424 2040 2426 2082
rect 2432 2052 2434 2086
rect 2454 2085 2460 2086
rect 2454 2081 2455 2085
rect 2459 2081 2460 2085
rect 2454 2080 2460 2081
rect 2470 2058 2476 2059
rect 2470 2054 2471 2058
rect 2475 2054 2476 2058
rect 2470 2053 2476 2054
rect 2430 2051 2436 2052
rect 2430 2047 2431 2051
rect 2435 2047 2436 2051
rect 2472 2047 2474 2053
rect 2480 2052 2482 2110
rect 2528 2103 2530 2114
rect 2527 2102 2531 2103
rect 2527 2097 2531 2098
rect 2528 2086 2530 2097
rect 2536 2092 2538 2146
rect 2542 2142 2543 2146
rect 2547 2142 2548 2146
rect 2542 2141 2548 2142
rect 2560 2116 2562 2158
rect 2583 2153 2587 2154
rect 2584 2138 2586 2153
rect 2582 2137 2588 2138
rect 2582 2133 2583 2137
rect 2587 2133 2588 2137
rect 2582 2132 2588 2133
rect 2582 2120 2588 2121
rect 2582 2116 2583 2120
rect 2587 2116 2588 2120
rect 2558 2115 2564 2116
rect 2582 2115 2588 2116
rect 2558 2111 2559 2115
rect 2563 2111 2564 2115
rect 2558 2110 2564 2111
rect 2584 2103 2586 2115
rect 2583 2102 2587 2103
rect 2583 2097 2587 2098
rect 2534 2091 2540 2092
rect 2534 2087 2535 2091
rect 2539 2087 2540 2091
rect 2534 2086 2540 2087
rect 2526 2085 2532 2086
rect 2584 2085 2586 2097
rect 2526 2081 2527 2085
rect 2531 2081 2532 2085
rect 2526 2080 2532 2081
rect 2582 2084 2588 2085
rect 2582 2080 2583 2084
rect 2587 2080 2588 2084
rect 2582 2079 2588 2080
rect 2582 2067 2588 2068
rect 2582 2063 2583 2067
rect 2587 2063 2588 2067
rect 2582 2062 2588 2063
rect 2542 2058 2548 2059
rect 2542 2054 2543 2058
rect 2547 2054 2548 2058
rect 2542 2053 2548 2054
rect 2478 2051 2484 2052
rect 2478 2047 2479 2051
rect 2483 2047 2484 2051
rect 2544 2047 2546 2053
rect 2558 2051 2564 2052
rect 2558 2047 2559 2051
rect 2563 2047 2564 2051
rect 2584 2047 2586 2062
rect 2430 2046 2436 2047
rect 2447 2046 2451 2047
rect 2447 2041 2451 2042
rect 2471 2046 2475 2047
rect 2478 2046 2484 2047
rect 2543 2046 2547 2047
rect 2558 2046 2564 2047
rect 2583 2046 2587 2047
rect 2471 2041 2475 2042
rect 2543 2041 2547 2042
rect 2422 2039 2428 2040
rect 2422 2035 2423 2039
rect 2427 2035 2428 2039
rect 2448 2035 2450 2041
rect 2544 2035 2546 2041
rect 2110 2034 2116 2035
rect 2130 2034 2136 2035
rect 2214 2034 2220 2035
rect 2234 2034 2240 2035
rect 2326 2034 2332 2035
rect 2422 2034 2428 2035
rect 2446 2034 2452 2035
rect 2110 2030 2111 2034
rect 2115 2030 2116 2034
rect 2110 2029 2116 2030
rect 2054 2015 2060 2016
rect 2054 2011 2055 2015
rect 2059 2011 2060 2015
rect 2054 2010 2060 2011
rect 1990 2007 1996 2008
rect 1918 2003 1924 2004
rect 1918 1999 1919 2003
rect 1923 1999 1924 2003
rect 1990 2003 1991 2007
rect 1995 2003 1996 2007
rect 1990 2002 1996 2003
rect 2094 2007 2100 2008
rect 2094 2003 2095 2007
rect 2099 2003 2100 2007
rect 2132 2004 2134 2034
rect 2214 2030 2215 2034
rect 2219 2030 2220 2034
rect 2214 2029 2220 2030
rect 2198 2007 2204 2008
rect 2094 2002 2100 2003
rect 2130 2003 2136 2004
rect 1918 1998 1924 1999
rect 1992 1991 1994 2002
rect 2096 1991 2098 2002
rect 2130 1999 2131 2003
rect 2135 1999 2136 2003
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2236 2004 2238 2034
rect 2326 2030 2327 2034
rect 2331 2030 2332 2034
rect 2326 2029 2332 2030
rect 2446 2030 2447 2034
rect 2451 2030 2452 2034
rect 2446 2029 2452 2030
rect 2542 2034 2548 2035
rect 2542 2030 2543 2034
rect 2547 2030 2548 2034
rect 2542 2029 2548 2030
rect 2310 2007 2316 2008
rect 2198 2002 2204 2003
rect 2234 2003 2240 2004
rect 2130 1998 2136 1999
rect 2200 1991 2202 2002
rect 2234 1999 2235 2003
rect 2239 1999 2240 2003
rect 2310 2003 2311 2007
rect 2315 2003 2316 2007
rect 2310 2002 2316 2003
rect 2430 2007 2436 2008
rect 2430 2003 2431 2007
rect 2435 2003 2436 2007
rect 2430 2002 2436 2003
rect 2526 2007 2532 2008
rect 2526 2003 2527 2007
rect 2531 2003 2532 2007
rect 2560 2004 2562 2046
rect 2583 2041 2587 2042
rect 2584 2026 2586 2041
rect 2582 2025 2588 2026
rect 2582 2021 2583 2025
rect 2587 2021 2588 2025
rect 2582 2020 2588 2021
rect 2582 2008 2588 2009
rect 2582 2004 2583 2008
rect 2587 2004 2588 2008
rect 2526 2002 2532 2003
rect 2558 2003 2564 2004
rect 2582 2003 2588 2004
rect 2234 1998 2240 1999
rect 2312 1991 2314 2002
rect 2432 1991 2434 2002
rect 2528 1991 2530 2002
rect 2558 1999 2559 2003
rect 2563 1999 2564 2003
rect 2558 1998 2564 1999
rect 2584 1991 2586 2003
rect 1927 1990 1931 1991
rect 1927 1985 1931 1986
rect 1991 1990 1995 1991
rect 1991 1985 1995 1986
rect 2007 1990 2011 1991
rect 2007 1985 2011 1986
rect 2087 1990 2091 1991
rect 2087 1985 2091 1986
rect 2095 1990 2099 1991
rect 2095 1985 2099 1986
rect 2199 1990 2203 1991
rect 2199 1985 2203 1986
rect 2311 1990 2315 1991
rect 2311 1985 2315 1986
rect 2431 1990 2435 1991
rect 2431 1985 2435 1986
rect 2527 1990 2531 1991
rect 2527 1985 2531 1986
rect 2583 1990 2587 1991
rect 2583 1985 2587 1986
rect 1894 1983 1900 1984
rect 1894 1979 1895 1983
rect 1899 1979 1900 1983
rect 1894 1978 1900 1979
rect 1918 1975 1924 1976
rect 1766 1973 1772 1974
rect 1766 1969 1767 1973
rect 1771 1969 1772 1973
rect 1766 1968 1772 1969
rect 1846 1973 1852 1974
rect 1846 1969 1847 1973
rect 1851 1969 1852 1973
rect 1918 1971 1919 1975
rect 1923 1971 1924 1975
rect 1928 1974 1930 1985
rect 1998 1975 2004 1976
rect 1918 1970 1924 1971
rect 1926 1973 1932 1974
rect 1846 1968 1852 1969
rect 1782 1946 1788 1947
rect 1782 1942 1783 1946
rect 1787 1942 1788 1946
rect 1782 1941 1788 1942
rect 1862 1946 1868 1947
rect 1862 1942 1863 1946
rect 1867 1942 1868 1946
rect 1862 1941 1868 1942
rect 1758 1939 1764 1940
rect 1758 1935 1759 1939
rect 1763 1935 1764 1939
rect 1758 1934 1764 1935
rect 1784 1931 1786 1941
rect 1842 1939 1848 1940
rect 1842 1935 1843 1939
rect 1847 1935 1848 1939
rect 1842 1934 1848 1935
rect 1719 1930 1723 1931
rect 1695 1925 1699 1926
rect 1706 1927 1712 1928
rect 734 1922 740 1923
rect 759 1922 763 1923
rect 663 1917 667 1918
rect 494 1915 500 1916
rect 494 1911 495 1915
rect 499 1911 500 1915
rect 544 1911 546 1917
rect 630 1915 636 1916
rect 630 1911 631 1915
rect 635 1911 636 1915
rect 656 1911 658 1917
rect 134 1910 140 1911
rect 158 1910 164 1911
rect 222 1910 228 1911
rect 230 1910 236 1911
rect 302 1910 308 1911
rect 326 1910 332 1911
rect 422 1910 428 1911
rect 430 1910 436 1911
rect 494 1910 500 1911
rect 542 1910 548 1911
rect 630 1910 636 1911
rect 654 1910 660 1911
rect 110 1901 116 1902
rect 110 1897 111 1901
rect 115 1897 116 1901
rect 110 1896 116 1897
rect 136 1892 138 1910
rect 158 1906 159 1910
rect 163 1906 164 1910
rect 158 1905 164 1906
rect 134 1891 140 1892
rect 134 1887 135 1891
rect 139 1887 140 1891
rect 134 1886 140 1887
rect 110 1884 116 1885
rect 110 1880 111 1884
rect 115 1880 116 1884
rect 110 1879 116 1880
rect 142 1883 148 1884
rect 142 1879 143 1883
rect 147 1879 148 1883
rect 214 1883 220 1884
rect 112 1859 114 1879
rect 142 1878 148 1879
rect 166 1879 172 1880
rect 144 1859 146 1878
rect 166 1875 167 1879
rect 171 1875 172 1879
rect 214 1879 215 1883
rect 219 1879 220 1883
rect 214 1878 220 1879
rect 166 1874 172 1875
rect 111 1858 115 1859
rect 111 1853 115 1854
rect 143 1858 147 1859
rect 143 1853 147 1854
rect 112 1841 114 1853
rect 144 1842 146 1853
rect 142 1841 148 1842
rect 110 1840 116 1841
rect 110 1836 111 1840
rect 115 1836 116 1840
rect 142 1837 143 1841
rect 147 1837 148 1841
rect 142 1836 148 1837
rect 110 1835 116 1836
rect 110 1823 116 1824
rect 110 1819 111 1823
rect 115 1819 116 1823
rect 110 1818 116 1819
rect 112 1799 114 1818
rect 158 1814 164 1815
rect 158 1810 159 1814
rect 163 1810 164 1814
rect 158 1809 164 1810
rect 160 1799 162 1809
rect 168 1808 170 1874
rect 216 1859 218 1878
rect 224 1872 226 1910
rect 230 1906 231 1910
rect 235 1906 236 1910
rect 230 1905 236 1906
rect 304 1892 306 1910
rect 326 1906 327 1910
rect 331 1906 332 1910
rect 326 1905 332 1906
rect 302 1891 308 1892
rect 302 1887 303 1891
rect 307 1887 308 1891
rect 302 1886 308 1887
rect 310 1883 316 1884
rect 310 1879 311 1883
rect 315 1879 316 1883
rect 310 1878 316 1879
rect 414 1883 420 1884
rect 414 1879 415 1883
rect 419 1879 420 1883
rect 414 1878 420 1879
rect 222 1871 228 1872
rect 222 1867 223 1871
rect 227 1867 228 1871
rect 222 1866 228 1867
rect 312 1859 314 1878
rect 416 1859 418 1878
rect 424 1872 426 1910
rect 430 1906 431 1910
rect 435 1906 436 1910
rect 430 1905 436 1906
rect 542 1906 543 1910
rect 547 1906 548 1910
rect 542 1905 548 1906
rect 632 1892 634 1910
rect 654 1906 655 1910
rect 659 1906 660 1910
rect 654 1905 660 1906
rect 630 1891 636 1892
rect 630 1887 631 1891
rect 635 1887 636 1891
rect 630 1886 636 1887
rect 526 1883 532 1884
rect 526 1879 527 1883
rect 531 1879 532 1883
rect 526 1878 532 1879
rect 638 1883 644 1884
rect 638 1879 639 1883
rect 643 1879 644 1883
rect 672 1880 674 1922
rect 759 1917 763 1918
rect 767 1922 771 1923
rect 854 1922 860 1923
rect 879 1922 883 1923
rect 767 1917 771 1918
rect 846 1919 852 1920
rect 768 1911 770 1917
rect 846 1915 847 1919
rect 851 1915 852 1919
rect 879 1917 883 1918
rect 983 1922 987 1923
rect 990 1922 996 1923
rect 1015 1922 1019 1923
rect 983 1917 987 1918
rect 1015 1917 1019 1918
rect 1087 1922 1091 1923
rect 1134 1922 1140 1923
rect 1159 1922 1163 1923
rect 1087 1917 1091 1918
rect 1159 1917 1163 1918
rect 1199 1922 1203 1923
rect 1218 1922 1224 1923
rect 1287 1922 1291 1923
rect 1199 1917 1203 1918
rect 846 1914 852 1915
rect 854 1915 860 1916
rect 766 1910 772 1911
rect 766 1906 767 1910
rect 771 1906 772 1910
rect 766 1905 772 1906
rect 750 1883 756 1884
rect 638 1878 644 1879
rect 670 1879 676 1880
rect 422 1871 428 1872
rect 422 1867 423 1871
rect 427 1867 428 1871
rect 422 1866 428 1867
rect 528 1859 530 1878
rect 640 1859 642 1878
rect 670 1875 671 1879
rect 675 1875 676 1879
rect 750 1879 751 1883
rect 755 1879 756 1883
rect 750 1878 756 1879
rect 670 1874 676 1875
rect 752 1859 754 1878
rect 848 1876 850 1914
rect 854 1911 855 1915
rect 859 1911 860 1915
rect 880 1911 882 1917
rect 974 1915 980 1916
rect 974 1911 975 1915
rect 979 1911 980 1915
rect 984 1911 986 1917
rect 1062 1915 1068 1916
rect 1062 1911 1063 1915
rect 1067 1911 1068 1915
rect 1088 1911 1090 1917
rect 1106 1915 1112 1916
rect 1106 1911 1107 1915
rect 1111 1911 1112 1915
rect 1200 1911 1202 1917
rect 854 1910 860 1911
rect 878 1910 884 1911
rect 974 1910 980 1911
rect 982 1910 988 1911
rect 1062 1910 1068 1911
rect 1086 1910 1092 1911
rect 1106 1910 1112 1911
rect 1198 1910 1204 1911
rect 856 1892 858 1910
rect 878 1906 879 1910
rect 883 1906 884 1910
rect 878 1905 884 1906
rect 854 1891 860 1892
rect 854 1887 855 1891
rect 859 1887 860 1891
rect 854 1886 860 1887
rect 862 1883 868 1884
rect 862 1879 863 1883
rect 867 1879 868 1883
rect 862 1878 868 1879
rect 966 1883 972 1884
rect 966 1879 967 1883
rect 971 1879 972 1883
rect 966 1878 972 1879
rect 846 1875 852 1876
rect 846 1871 847 1875
rect 851 1871 852 1875
rect 846 1870 852 1871
rect 864 1859 866 1878
rect 968 1859 970 1878
rect 199 1858 203 1859
rect 199 1853 203 1854
rect 215 1858 219 1859
rect 215 1853 219 1854
rect 263 1858 267 1859
rect 263 1853 267 1854
rect 311 1858 315 1859
rect 311 1853 315 1854
rect 351 1858 355 1859
rect 351 1853 355 1854
rect 415 1858 419 1859
rect 415 1853 419 1854
rect 439 1858 443 1859
rect 439 1853 443 1854
rect 527 1858 531 1859
rect 527 1853 531 1854
rect 535 1858 539 1859
rect 535 1853 539 1854
rect 623 1858 627 1859
rect 623 1853 627 1854
rect 639 1858 643 1859
rect 639 1853 643 1854
rect 711 1858 715 1859
rect 711 1853 715 1854
rect 751 1858 755 1859
rect 751 1853 755 1854
rect 791 1858 795 1859
rect 791 1853 795 1854
rect 863 1858 867 1859
rect 863 1853 867 1854
rect 871 1858 875 1859
rect 871 1853 875 1854
rect 951 1858 955 1859
rect 951 1853 955 1854
rect 967 1858 971 1859
rect 967 1853 971 1854
rect 190 1843 196 1844
rect 190 1839 191 1843
rect 195 1839 196 1843
rect 200 1842 202 1853
rect 254 1843 260 1844
rect 190 1838 196 1839
rect 198 1841 204 1842
rect 192 1808 194 1838
rect 198 1837 199 1841
rect 203 1837 204 1841
rect 254 1839 255 1843
rect 259 1839 260 1843
rect 264 1842 266 1853
rect 342 1843 348 1844
rect 254 1838 260 1839
rect 262 1841 268 1842
rect 198 1836 204 1837
rect 214 1814 220 1815
rect 214 1810 215 1814
rect 219 1810 220 1814
rect 214 1809 220 1810
rect 166 1807 172 1808
rect 166 1803 167 1807
rect 171 1803 172 1807
rect 166 1802 172 1803
rect 190 1807 196 1808
rect 190 1803 191 1807
rect 195 1803 196 1807
rect 190 1802 196 1803
rect 216 1799 218 1809
rect 256 1808 258 1838
rect 262 1837 263 1841
rect 267 1837 268 1841
rect 342 1839 343 1843
rect 347 1839 348 1843
rect 352 1842 354 1853
rect 430 1843 436 1844
rect 342 1838 348 1839
rect 350 1841 356 1842
rect 262 1836 268 1837
rect 278 1814 284 1815
rect 278 1810 279 1814
rect 283 1810 284 1814
rect 278 1809 284 1810
rect 254 1807 260 1808
rect 254 1803 255 1807
rect 259 1803 260 1807
rect 254 1802 260 1803
rect 280 1799 282 1809
rect 344 1808 346 1838
rect 350 1837 351 1841
rect 355 1837 356 1841
rect 430 1839 431 1843
rect 435 1839 436 1843
rect 440 1842 442 1853
rect 526 1843 532 1844
rect 430 1838 436 1839
rect 438 1841 444 1842
rect 350 1836 356 1837
rect 366 1814 372 1815
rect 366 1810 367 1814
rect 371 1810 372 1814
rect 366 1809 372 1810
rect 342 1807 348 1808
rect 342 1803 343 1807
rect 347 1803 348 1807
rect 342 1802 348 1803
rect 368 1799 370 1809
rect 432 1808 434 1838
rect 438 1837 439 1841
rect 443 1837 444 1841
rect 526 1839 527 1843
rect 531 1839 532 1843
rect 536 1842 538 1853
rect 558 1843 564 1844
rect 526 1838 532 1839
rect 534 1841 540 1842
rect 438 1836 444 1837
rect 454 1814 460 1815
rect 454 1810 455 1814
rect 459 1810 460 1814
rect 454 1809 460 1810
rect 430 1807 436 1808
rect 430 1803 431 1807
rect 435 1803 436 1807
rect 430 1802 436 1803
rect 456 1799 458 1809
rect 528 1808 530 1838
rect 534 1837 535 1841
rect 539 1837 540 1841
rect 558 1839 559 1843
rect 563 1839 564 1843
rect 624 1842 626 1853
rect 702 1843 708 1844
rect 558 1838 564 1839
rect 622 1841 628 1842
rect 534 1836 540 1837
rect 550 1814 556 1815
rect 550 1810 551 1814
rect 555 1810 556 1814
rect 550 1809 556 1810
rect 526 1807 532 1808
rect 526 1803 527 1807
rect 531 1803 532 1807
rect 526 1802 532 1803
rect 552 1799 554 1809
rect 560 1800 562 1838
rect 622 1837 623 1841
rect 627 1837 628 1841
rect 702 1839 703 1843
rect 707 1839 708 1843
rect 712 1842 714 1853
rect 782 1843 788 1844
rect 702 1838 708 1839
rect 710 1841 716 1842
rect 622 1836 628 1837
rect 638 1814 644 1815
rect 638 1810 639 1814
rect 643 1810 644 1814
rect 638 1809 644 1810
rect 630 1807 636 1808
rect 630 1803 631 1807
rect 635 1803 636 1807
rect 630 1802 636 1803
rect 558 1799 564 1800
rect 111 1798 115 1799
rect 111 1793 115 1794
rect 159 1798 163 1799
rect 159 1793 163 1794
rect 215 1798 219 1799
rect 215 1793 219 1794
rect 231 1798 235 1799
rect 231 1793 235 1794
rect 279 1798 283 1799
rect 279 1793 283 1794
rect 295 1798 299 1799
rect 295 1793 299 1794
rect 367 1798 371 1799
rect 367 1793 371 1794
rect 447 1798 451 1799
rect 447 1793 451 1794
rect 455 1798 459 1799
rect 455 1793 459 1794
rect 535 1798 539 1799
rect 535 1793 539 1794
rect 551 1798 555 1799
rect 558 1795 559 1799
rect 563 1795 564 1799
rect 558 1794 564 1795
rect 623 1798 627 1799
rect 551 1793 555 1794
rect 623 1793 627 1794
rect 112 1778 114 1793
rect 232 1787 234 1793
rect 250 1791 256 1792
rect 250 1787 251 1791
rect 255 1787 256 1791
rect 296 1787 298 1793
rect 314 1791 320 1792
rect 314 1787 315 1791
rect 319 1787 320 1791
rect 368 1787 370 1793
rect 386 1791 392 1792
rect 386 1787 387 1791
rect 391 1787 392 1791
rect 448 1787 450 1793
rect 466 1791 472 1792
rect 466 1787 467 1791
rect 471 1787 472 1791
rect 536 1787 538 1793
rect 598 1791 604 1792
rect 598 1787 599 1791
rect 603 1787 604 1791
rect 624 1787 626 1793
rect 230 1786 236 1787
rect 250 1786 256 1787
rect 294 1786 300 1787
rect 314 1786 320 1787
rect 366 1786 372 1787
rect 386 1786 392 1787
rect 446 1786 452 1787
rect 466 1786 472 1787
rect 534 1786 540 1787
rect 598 1786 604 1787
rect 622 1786 628 1787
rect 230 1782 231 1786
rect 235 1782 236 1786
rect 230 1781 236 1782
rect 110 1777 116 1778
rect 110 1773 111 1777
rect 115 1773 116 1777
rect 110 1772 116 1773
rect 110 1760 116 1761
rect 110 1756 111 1760
rect 115 1756 116 1760
rect 110 1755 116 1756
rect 214 1759 220 1760
rect 214 1755 215 1759
rect 219 1755 220 1759
rect 252 1756 254 1786
rect 294 1782 295 1786
rect 299 1782 300 1786
rect 294 1781 300 1782
rect 278 1759 284 1760
rect 112 1739 114 1755
rect 214 1754 220 1755
rect 250 1755 256 1756
rect 216 1739 218 1754
rect 250 1751 251 1755
rect 255 1751 256 1755
rect 278 1755 279 1759
rect 283 1755 284 1759
rect 316 1756 318 1786
rect 366 1782 367 1786
rect 371 1782 372 1786
rect 366 1781 372 1782
rect 350 1759 356 1760
rect 278 1754 284 1755
rect 314 1755 320 1756
rect 250 1750 256 1751
rect 280 1739 282 1754
rect 314 1751 315 1755
rect 319 1751 320 1755
rect 350 1755 351 1759
rect 355 1755 356 1759
rect 388 1756 390 1786
rect 446 1782 447 1786
rect 451 1782 452 1786
rect 446 1781 452 1782
rect 430 1759 436 1760
rect 350 1754 356 1755
rect 386 1755 392 1756
rect 314 1750 320 1751
rect 352 1739 354 1754
rect 386 1751 387 1755
rect 391 1751 392 1755
rect 430 1755 431 1759
rect 435 1755 436 1759
rect 468 1756 470 1786
rect 534 1782 535 1786
rect 539 1782 540 1786
rect 534 1781 540 1782
rect 600 1768 602 1786
rect 622 1782 623 1786
rect 627 1782 628 1786
rect 622 1781 628 1782
rect 598 1767 604 1768
rect 598 1763 599 1767
rect 603 1763 604 1767
rect 598 1762 604 1763
rect 518 1759 524 1760
rect 430 1754 436 1755
rect 466 1755 472 1756
rect 386 1750 392 1751
rect 358 1747 364 1748
rect 358 1743 359 1747
rect 363 1743 364 1747
rect 358 1742 364 1743
rect 111 1738 115 1739
rect 111 1733 115 1734
rect 215 1738 219 1739
rect 215 1733 219 1734
rect 279 1738 283 1739
rect 279 1733 283 1734
rect 351 1738 355 1739
rect 351 1733 355 1734
rect 112 1721 114 1733
rect 352 1722 354 1733
rect 350 1721 356 1722
rect 110 1720 116 1721
rect 110 1716 111 1720
rect 115 1716 116 1720
rect 350 1717 351 1721
rect 355 1717 356 1721
rect 350 1716 356 1717
rect 110 1715 116 1716
rect 110 1703 116 1704
rect 110 1699 111 1703
rect 115 1699 116 1703
rect 110 1698 116 1699
rect 112 1679 114 1698
rect 360 1688 362 1742
rect 432 1739 434 1754
rect 466 1751 467 1755
rect 471 1751 472 1755
rect 518 1755 519 1759
rect 523 1755 524 1759
rect 518 1754 524 1755
rect 606 1759 612 1760
rect 606 1755 607 1759
rect 611 1755 612 1759
rect 632 1756 634 1802
rect 640 1799 642 1809
rect 704 1808 706 1838
rect 710 1837 711 1841
rect 715 1837 716 1841
rect 782 1839 783 1843
rect 787 1839 788 1843
rect 792 1842 794 1853
rect 862 1843 868 1844
rect 782 1838 788 1839
rect 790 1841 796 1842
rect 710 1836 716 1837
rect 726 1814 732 1815
rect 726 1810 727 1814
rect 731 1810 732 1814
rect 726 1809 732 1810
rect 702 1807 708 1808
rect 702 1803 703 1807
rect 707 1803 708 1807
rect 702 1802 708 1803
rect 728 1799 730 1809
rect 784 1808 786 1838
rect 790 1837 791 1841
rect 795 1837 796 1841
rect 862 1839 863 1843
rect 867 1839 868 1843
rect 872 1842 874 1853
rect 942 1843 948 1844
rect 862 1838 868 1839
rect 870 1841 876 1842
rect 790 1836 796 1837
rect 806 1814 812 1815
rect 806 1810 807 1814
rect 811 1810 812 1814
rect 806 1809 812 1810
rect 782 1807 788 1808
rect 782 1803 783 1807
rect 787 1803 788 1807
rect 782 1802 788 1803
rect 808 1799 810 1809
rect 864 1808 866 1838
rect 870 1837 871 1841
rect 875 1837 876 1841
rect 942 1839 943 1843
rect 947 1839 948 1843
rect 952 1842 954 1853
rect 976 1852 978 1910
rect 982 1906 983 1910
rect 987 1906 988 1910
rect 982 1905 988 1906
rect 1064 1892 1066 1910
rect 1086 1906 1087 1910
rect 1091 1906 1092 1910
rect 1086 1905 1092 1906
rect 1062 1891 1068 1892
rect 1062 1887 1063 1891
rect 1067 1887 1068 1891
rect 1062 1886 1068 1887
rect 1070 1883 1076 1884
rect 1070 1879 1071 1883
rect 1075 1879 1076 1883
rect 1108 1880 1110 1910
rect 1198 1906 1199 1910
rect 1203 1906 1204 1910
rect 1198 1905 1204 1906
rect 1182 1883 1188 1884
rect 1070 1878 1076 1879
rect 1106 1879 1112 1880
rect 1072 1859 1074 1878
rect 1106 1875 1107 1879
rect 1111 1875 1112 1879
rect 1182 1879 1183 1883
rect 1187 1879 1188 1883
rect 1220 1880 1222 1922
rect 1287 1917 1291 1918
rect 1327 1922 1331 1923
rect 1327 1917 1331 1918
rect 1278 1915 1284 1916
rect 1278 1911 1279 1915
rect 1283 1911 1284 1915
rect 1288 1911 1290 1917
rect 1278 1910 1284 1911
rect 1286 1910 1292 1911
rect 1270 1883 1276 1884
rect 1182 1878 1188 1879
rect 1218 1879 1224 1880
rect 1106 1874 1112 1875
rect 1184 1859 1186 1878
rect 1218 1875 1219 1879
rect 1223 1875 1224 1879
rect 1270 1879 1271 1883
rect 1275 1879 1276 1883
rect 1270 1878 1276 1879
rect 1218 1874 1224 1875
rect 1272 1859 1274 1878
rect 1280 1860 1282 1910
rect 1286 1906 1287 1910
rect 1291 1906 1292 1910
rect 1286 1905 1292 1906
rect 1328 1902 1330 1917
rect 1368 1910 1370 1925
rect 1706 1923 1707 1927
rect 1711 1923 1712 1927
rect 1719 1925 1723 1926
rect 1775 1930 1779 1931
rect 1775 1925 1779 1926
rect 1783 1930 1787 1931
rect 1783 1925 1787 1926
rect 1831 1930 1835 1931
rect 1831 1925 1835 1926
rect 1706 1922 1712 1923
rect 1720 1919 1722 1925
rect 1738 1923 1744 1924
rect 1738 1919 1739 1923
rect 1743 1919 1744 1923
rect 1776 1919 1778 1925
rect 1806 1923 1812 1924
rect 1806 1919 1807 1923
rect 1811 1919 1812 1923
rect 1832 1919 1834 1925
rect 1718 1918 1724 1919
rect 1738 1918 1744 1919
rect 1774 1918 1780 1919
rect 1806 1918 1812 1919
rect 1830 1918 1836 1919
rect 1718 1914 1719 1918
rect 1723 1914 1724 1918
rect 1718 1913 1724 1914
rect 1366 1909 1372 1910
rect 1366 1905 1367 1909
rect 1371 1905 1372 1909
rect 1366 1904 1372 1905
rect 1326 1901 1332 1902
rect 1326 1897 1327 1901
rect 1331 1897 1332 1901
rect 1326 1896 1332 1897
rect 1366 1892 1372 1893
rect 1366 1888 1367 1892
rect 1371 1888 1372 1892
rect 1366 1887 1372 1888
rect 1702 1891 1708 1892
rect 1702 1887 1703 1891
rect 1707 1887 1708 1891
rect 1740 1888 1742 1918
rect 1774 1914 1775 1918
rect 1779 1914 1780 1918
rect 1774 1913 1780 1914
rect 1808 1900 1810 1918
rect 1830 1914 1831 1918
rect 1835 1914 1836 1918
rect 1830 1913 1836 1914
rect 1806 1899 1812 1900
rect 1806 1895 1807 1899
rect 1811 1895 1812 1899
rect 1806 1894 1812 1895
rect 1758 1891 1764 1892
rect 1326 1884 1332 1885
rect 1326 1880 1327 1884
rect 1331 1880 1332 1884
rect 1326 1879 1332 1880
rect 1278 1859 1284 1860
rect 1328 1859 1330 1879
rect 1368 1871 1370 1887
rect 1702 1886 1708 1887
rect 1738 1887 1744 1888
rect 1704 1871 1706 1886
rect 1738 1883 1739 1887
rect 1743 1883 1744 1887
rect 1758 1887 1759 1891
rect 1763 1887 1764 1891
rect 1814 1891 1820 1892
rect 1758 1886 1764 1887
rect 1782 1887 1788 1888
rect 1738 1882 1744 1883
rect 1760 1871 1762 1886
rect 1782 1883 1783 1887
rect 1787 1883 1788 1887
rect 1814 1887 1815 1891
rect 1819 1887 1820 1891
rect 1844 1888 1846 1934
rect 1864 1931 1866 1941
rect 1920 1940 1922 1970
rect 1926 1969 1927 1973
rect 1931 1969 1932 1973
rect 1998 1971 1999 1975
rect 2003 1971 2004 1975
rect 2008 1974 2010 1985
rect 2078 1975 2084 1976
rect 1998 1970 2004 1971
rect 2006 1973 2012 1974
rect 1926 1968 1932 1969
rect 1942 1946 1948 1947
rect 1942 1942 1943 1946
rect 1947 1942 1948 1946
rect 1942 1941 1948 1942
rect 1918 1939 1924 1940
rect 1918 1935 1919 1939
rect 1923 1935 1924 1939
rect 1918 1934 1924 1935
rect 1944 1931 1946 1941
rect 2000 1940 2002 1970
rect 2006 1969 2007 1973
rect 2011 1969 2012 1973
rect 2078 1971 2079 1975
rect 2083 1971 2084 1975
rect 2088 1974 2090 1985
rect 2078 1970 2084 1971
rect 2086 1973 2092 1974
rect 2584 1973 2586 1985
rect 2006 1968 2012 1969
rect 2022 1946 2028 1947
rect 2022 1942 2023 1946
rect 2027 1942 2028 1946
rect 2022 1941 2028 1942
rect 1998 1939 2004 1940
rect 1998 1935 1999 1939
rect 2003 1935 2004 1939
rect 1998 1934 2004 1935
rect 1958 1931 1964 1932
rect 2024 1931 2026 1941
rect 2080 1940 2082 1970
rect 2086 1969 2087 1973
rect 2091 1969 2092 1973
rect 2086 1968 2092 1969
rect 2582 1972 2588 1973
rect 2582 1968 2583 1972
rect 2587 1968 2588 1972
rect 2582 1967 2588 1968
rect 2582 1955 2588 1956
rect 2582 1951 2583 1955
rect 2587 1951 2588 1955
rect 2582 1950 2588 1951
rect 2102 1946 2108 1947
rect 2102 1942 2103 1946
rect 2107 1942 2108 1946
rect 2102 1941 2108 1942
rect 2078 1939 2084 1940
rect 2078 1935 2079 1939
rect 2083 1935 2084 1939
rect 2078 1934 2084 1935
rect 2104 1931 2106 1941
rect 2134 1931 2140 1932
rect 2584 1931 2586 1950
rect 1863 1930 1867 1931
rect 1863 1925 1867 1926
rect 1887 1930 1891 1931
rect 1887 1925 1891 1926
rect 1943 1930 1947 1931
rect 1958 1927 1959 1931
rect 1963 1927 1964 1931
rect 1958 1926 1964 1927
rect 1999 1930 2003 1931
rect 1943 1925 1947 1926
rect 1888 1919 1890 1925
rect 1918 1923 1924 1924
rect 1918 1919 1919 1923
rect 1923 1919 1924 1923
rect 1944 1919 1946 1925
rect 1886 1918 1892 1919
rect 1918 1918 1924 1919
rect 1942 1918 1948 1919
rect 1886 1914 1887 1918
rect 1891 1914 1892 1918
rect 1886 1913 1892 1914
rect 1920 1900 1922 1918
rect 1942 1914 1943 1918
rect 1947 1914 1948 1918
rect 1942 1913 1948 1914
rect 1918 1899 1924 1900
rect 1918 1895 1919 1899
rect 1923 1895 1924 1899
rect 1918 1894 1924 1895
rect 1870 1891 1876 1892
rect 1814 1886 1820 1887
rect 1842 1887 1848 1888
rect 1782 1882 1788 1883
rect 1367 1870 1371 1871
rect 1367 1865 1371 1866
rect 1399 1870 1403 1871
rect 1399 1865 1403 1866
rect 1463 1870 1467 1871
rect 1463 1865 1467 1866
rect 1559 1870 1563 1871
rect 1559 1865 1563 1866
rect 1655 1870 1659 1871
rect 1655 1865 1659 1866
rect 1703 1870 1707 1871
rect 1703 1865 1707 1866
rect 1743 1870 1747 1871
rect 1743 1865 1747 1866
rect 1759 1870 1763 1871
rect 1759 1865 1763 1866
rect 1039 1858 1043 1859
rect 1039 1853 1043 1854
rect 1071 1858 1075 1859
rect 1071 1853 1075 1854
rect 1183 1858 1187 1859
rect 1183 1853 1187 1854
rect 1271 1858 1275 1859
rect 1278 1855 1279 1859
rect 1283 1855 1284 1859
rect 1278 1854 1284 1855
rect 1327 1858 1331 1859
rect 1271 1853 1275 1854
rect 1327 1853 1331 1854
rect 1368 1853 1370 1865
rect 1400 1854 1402 1865
rect 1464 1854 1466 1865
rect 1560 1854 1562 1865
rect 1656 1854 1658 1865
rect 1714 1859 1720 1860
rect 1714 1855 1715 1859
rect 1719 1855 1720 1859
rect 1714 1854 1720 1855
rect 1744 1854 1746 1865
rect 1398 1853 1404 1854
rect 974 1851 980 1852
rect 974 1847 975 1851
rect 979 1847 980 1851
rect 974 1846 980 1847
rect 1030 1843 1036 1844
rect 942 1838 948 1839
rect 950 1841 956 1842
rect 870 1836 876 1837
rect 886 1814 892 1815
rect 886 1810 887 1814
rect 891 1810 892 1814
rect 886 1809 892 1810
rect 862 1807 868 1808
rect 862 1803 863 1807
rect 867 1803 868 1807
rect 862 1802 868 1803
rect 888 1799 890 1809
rect 639 1798 643 1799
rect 639 1793 643 1794
rect 711 1798 715 1799
rect 711 1793 715 1794
rect 727 1798 731 1799
rect 727 1793 731 1794
rect 791 1798 795 1799
rect 791 1793 795 1794
rect 807 1798 811 1799
rect 807 1793 811 1794
rect 871 1798 875 1799
rect 871 1793 875 1794
rect 887 1798 891 1799
rect 944 1796 946 1838
rect 950 1837 951 1841
rect 955 1837 956 1841
rect 1030 1839 1031 1843
rect 1035 1839 1036 1843
rect 1040 1842 1042 1853
rect 1030 1838 1036 1839
rect 1038 1841 1044 1842
rect 1328 1841 1330 1853
rect 1366 1852 1372 1853
rect 1366 1848 1367 1852
rect 1371 1848 1372 1852
rect 1398 1849 1399 1853
rect 1403 1849 1404 1853
rect 1398 1848 1404 1849
rect 1462 1853 1468 1854
rect 1462 1849 1463 1853
rect 1467 1849 1468 1853
rect 1462 1848 1468 1849
rect 1558 1853 1564 1854
rect 1558 1849 1559 1853
rect 1563 1849 1564 1853
rect 1558 1848 1564 1849
rect 1654 1853 1660 1854
rect 1654 1849 1655 1853
rect 1659 1849 1660 1853
rect 1654 1848 1660 1849
rect 1366 1847 1372 1848
rect 950 1836 956 1837
rect 966 1814 972 1815
rect 966 1810 967 1814
rect 971 1810 972 1814
rect 966 1809 972 1810
rect 958 1807 964 1808
rect 958 1803 959 1807
rect 963 1803 964 1807
rect 958 1802 964 1803
rect 951 1798 955 1799
rect 887 1793 891 1794
rect 942 1795 948 1796
rect 712 1787 714 1793
rect 726 1787 732 1788
rect 792 1787 794 1793
rect 862 1791 868 1792
rect 862 1787 863 1791
rect 867 1787 868 1791
rect 872 1787 874 1793
rect 910 1791 916 1792
rect 910 1787 911 1791
rect 915 1787 916 1791
rect 942 1791 943 1795
rect 947 1791 948 1795
rect 951 1793 955 1794
rect 942 1790 948 1791
rect 952 1787 954 1793
rect 710 1786 716 1787
rect 710 1782 711 1786
rect 715 1782 716 1786
rect 726 1783 727 1787
rect 731 1783 732 1787
rect 726 1782 732 1783
rect 790 1786 796 1787
rect 862 1786 868 1787
rect 870 1786 876 1787
rect 910 1786 916 1787
rect 950 1786 956 1787
rect 790 1782 791 1786
rect 795 1782 796 1786
rect 710 1781 716 1782
rect 694 1759 700 1760
rect 606 1754 612 1755
rect 630 1755 636 1756
rect 466 1750 472 1751
rect 520 1739 522 1754
rect 608 1739 610 1754
rect 630 1751 631 1755
rect 635 1751 636 1755
rect 694 1755 695 1759
rect 699 1755 700 1759
rect 728 1756 730 1782
rect 790 1781 796 1782
rect 774 1759 780 1760
rect 694 1754 700 1755
rect 726 1755 732 1756
rect 630 1750 636 1751
rect 696 1739 698 1754
rect 726 1751 727 1755
rect 731 1751 732 1755
rect 774 1755 775 1759
rect 779 1755 780 1759
rect 774 1754 780 1755
rect 854 1759 860 1760
rect 854 1755 855 1759
rect 859 1755 860 1759
rect 854 1754 860 1755
rect 726 1750 732 1751
rect 776 1739 778 1754
rect 856 1739 858 1754
rect 407 1738 411 1739
rect 407 1733 411 1734
rect 431 1738 435 1739
rect 431 1733 435 1734
rect 471 1738 475 1739
rect 471 1733 475 1734
rect 519 1738 523 1739
rect 519 1733 523 1734
rect 551 1738 555 1739
rect 551 1733 555 1734
rect 607 1738 611 1739
rect 607 1733 611 1734
rect 639 1738 643 1739
rect 639 1733 643 1734
rect 695 1738 699 1739
rect 695 1733 699 1734
rect 727 1738 731 1739
rect 727 1733 731 1734
rect 775 1738 779 1739
rect 775 1733 779 1734
rect 823 1738 827 1739
rect 823 1733 827 1734
rect 855 1738 859 1739
rect 855 1733 859 1734
rect 398 1723 404 1724
rect 398 1719 399 1723
rect 403 1719 404 1723
rect 408 1722 410 1733
rect 462 1723 468 1724
rect 398 1718 404 1719
rect 406 1721 412 1722
rect 366 1694 372 1695
rect 366 1690 367 1694
rect 371 1690 372 1694
rect 366 1689 372 1690
rect 358 1687 364 1688
rect 358 1683 359 1687
rect 363 1683 364 1687
rect 358 1682 364 1683
rect 368 1679 370 1689
rect 400 1688 402 1718
rect 406 1717 407 1721
rect 411 1717 412 1721
rect 462 1719 463 1723
rect 467 1719 468 1723
rect 472 1722 474 1733
rect 542 1723 548 1724
rect 462 1718 468 1719
rect 470 1721 476 1722
rect 406 1716 412 1717
rect 422 1694 428 1695
rect 422 1690 423 1694
rect 427 1690 428 1694
rect 422 1689 428 1690
rect 398 1687 404 1688
rect 398 1683 399 1687
rect 403 1683 404 1687
rect 398 1682 404 1683
rect 424 1679 426 1689
rect 464 1688 466 1718
rect 470 1717 471 1721
rect 475 1717 476 1721
rect 542 1719 543 1723
rect 547 1719 548 1723
rect 552 1722 554 1733
rect 582 1723 588 1724
rect 542 1718 548 1719
rect 550 1721 556 1722
rect 470 1716 476 1717
rect 486 1694 492 1695
rect 486 1690 487 1694
rect 491 1690 492 1694
rect 486 1689 492 1690
rect 462 1687 468 1688
rect 462 1683 463 1687
rect 467 1683 468 1687
rect 462 1682 468 1683
rect 488 1679 490 1689
rect 544 1688 546 1718
rect 550 1717 551 1721
rect 555 1717 556 1721
rect 582 1719 583 1723
rect 587 1719 588 1723
rect 640 1722 642 1733
rect 728 1722 730 1733
rect 824 1722 826 1733
rect 864 1732 866 1786
rect 870 1782 871 1786
rect 875 1782 876 1786
rect 870 1781 876 1782
rect 912 1760 914 1786
rect 950 1782 951 1786
rect 955 1782 956 1786
rect 950 1781 956 1782
rect 910 1759 916 1760
rect 910 1755 911 1759
rect 915 1755 916 1759
rect 910 1754 916 1755
rect 934 1759 940 1760
rect 934 1755 935 1759
rect 939 1755 940 1759
rect 960 1756 962 1802
rect 968 1799 970 1809
rect 1032 1808 1034 1838
rect 1038 1837 1039 1841
rect 1043 1837 1044 1841
rect 1038 1836 1044 1837
rect 1326 1840 1332 1841
rect 1326 1836 1327 1840
rect 1331 1836 1332 1840
rect 1326 1835 1332 1836
rect 1366 1835 1372 1836
rect 1366 1831 1367 1835
rect 1371 1831 1372 1835
rect 1366 1830 1372 1831
rect 1326 1823 1332 1824
rect 1326 1819 1327 1823
rect 1331 1819 1332 1823
rect 1326 1818 1332 1819
rect 1054 1814 1060 1815
rect 1054 1810 1055 1814
rect 1059 1810 1060 1814
rect 1054 1809 1060 1810
rect 1030 1807 1036 1808
rect 1030 1803 1031 1807
rect 1035 1803 1036 1807
rect 1030 1802 1036 1803
rect 1056 1799 1058 1809
rect 1328 1799 1330 1818
rect 1368 1815 1370 1830
rect 1414 1826 1420 1827
rect 1414 1822 1415 1826
rect 1419 1822 1420 1826
rect 1414 1821 1420 1822
rect 1478 1826 1484 1827
rect 1478 1822 1479 1826
rect 1483 1822 1484 1826
rect 1478 1821 1484 1822
rect 1574 1826 1580 1827
rect 1574 1822 1575 1826
rect 1579 1822 1580 1826
rect 1574 1821 1580 1822
rect 1670 1826 1676 1827
rect 1670 1822 1671 1826
rect 1675 1822 1676 1826
rect 1670 1821 1676 1822
rect 1416 1815 1418 1821
rect 1480 1815 1482 1821
rect 1576 1815 1578 1821
rect 1642 1819 1648 1820
rect 1642 1815 1643 1819
rect 1647 1815 1648 1819
rect 1672 1815 1674 1821
rect 1367 1814 1371 1815
rect 1367 1809 1371 1810
rect 1415 1814 1419 1815
rect 1415 1809 1419 1810
rect 1479 1814 1483 1815
rect 1479 1809 1483 1810
rect 1511 1814 1515 1815
rect 1511 1809 1515 1810
rect 1575 1814 1579 1815
rect 1575 1809 1579 1810
rect 1623 1814 1627 1815
rect 1642 1814 1648 1815
rect 1671 1814 1675 1815
rect 1623 1809 1627 1810
rect 967 1798 971 1799
rect 967 1793 971 1794
rect 1031 1798 1035 1799
rect 1031 1793 1035 1794
rect 1055 1798 1059 1799
rect 1055 1793 1059 1794
rect 1119 1798 1123 1799
rect 1119 1793 1123 1794
rect 1327 1798 1331 1799
rect 1368 1794 1370 1809
rect 1406 1807 1412 1808
rect 1406 1803 1407 1807
rect 1411 1803 1412 1807
rect 1416 1803 1418 1809
rect 1434 1807 1440 1808
rect 1434 1803 1435 1807
rect 1439 1803 1440 1807
rect 1512 1803 1514 1809
rect 1530 1807 1536 1808
rect 1530 1803 1531 1807
rect 1535 1803 1536 1807
rect 1624 1803 1626 1809
rect 1406 1802 1412 1803
rect 1414 1802 1420 1803
rect 1434 1802 1440 1803
rect 1510 1802 1516 1803
rect 1530 1802 1536 1803
rect 1622 1802 1628 1803
rect 1327 1793 1331 1794
rect 1366 1793 1372 1794
rect 1032 1787 1034 1793
rect 1120 1787 1122 1793
rect 1030 1786 1036 1787
rect 1030 1782 1031 1786
rect 1035 1782 1036 1786
rect 1030 1781 1036 1782
rect 1118 1786 1124 1787
rect 1118 1782 1119 1786
rect 1123 1782 1124 1786
rect 1118 1781 1124 1782
rect 1328 1778 1330 1793
rect 1366 1789 1367 1793
rect 1371 1789 1372 1793
rect 1366 1788 1372 1789
rect 1326 1777 1332 1778
rect 1326 1773 1327 1777
rect 1331 1773 1332 1777
rect 1326 1772 1332 1773
rect 1366 1776 1372 1777
rect 1366 1772 1367 1776
rect 1371 1772 1372 1776
rect 1366 1771 1372 1772
rect 1398 1775 1404 1776
rect 1398 1771 1399 1775
rect 1403 1771 1404 1775
rect 1326 1760 1332 1761
rect 1014 1759 1020 1760
rect 934 1754 940 1755
rect 958 1755 964 1756
rect 936 1739 938 1754
rect 958 1751 959 1755
rect 963 1751 964 1755
rect 1014 1755 1015 1759
rect 1019 1755 1020 1759
rect 1014 1754 1020 1755
rect 1102 1759 1108 1760
rect 1102 1755 1103 1759
rect 1107 1755 1108 1759
rect 1326 1756 1327 1760
rect 1331 1756 1332 1760
rect 1368 1759 1370 1771
rect 1398 1770 1404 1771
rect 1400 1759 1402 1770
rect 1326 1755 1332 1756
rect 1367 1758 1371 1759
rect 1102 1754 1108 1755
rect 958 1750 964 1751
rect 1016 1739 1018 1754
rect 1104 1739 1106 1754
rect 1328 1739 1330 1755
rect 1367 1753 1371 1754
rect 1399 1758 1403 1759
rect 1399 1753 1403 1754
rect 1368 1741 1370 1753
rect 1408 1748 1410 1802
rect 1414 1798 1415 1802
rect 1419 1798 1420 1802
rect 1414 1797 1420 1798
rect 1436 1772 1438 1802
rect 1510 1798 1511 1802
rect 1515 1798 1516 1802
rect 1510 1797 1516 1798
rect 1494 1775 1500 1776
rect 1434 1771 1440 1772
rect 1434 1767 1435 1771
rect 1439 1767 1440 1771
rect 1494 1771 1495 1775
rect 1499 1771 1500 1775
rect 1532 1772 1534 1802
rect 1622 1798 1623 1802
rect 1627 1798 1628 1802
rect 1622 1797 1628 1798
rect 1606 1775 1612 1776
rect 1494 1770 1500 1771
rect 1530 1771 1536 1772
rect 1434 1766 1440 1767
rect 1496 1759 1498 1770
rect 1530 1767 1531 1771
rect 1535 1767 1536 1771
rect 1606 1771 1607 1775
rect 1611 1771 1612 1775
rect 1644 1772 1646 1814
rect 1671 1809 1675 1810
rect 1716 1808 1718 1854
rect 1742 1853 1748 1854
rect 1742 1849 1743 1853
rect 1747 1849 1748 1853
rect 1742 1848 1748 1849
rect 1758 1826 1764 1827
rect 1758 1822 1759 1826
rect 1763 1822 1764 1826
rect 1758 1821 1764 1822
rect 1760 1815 1762 1821
rect 1784 1820 1786 1882
rect 1816 1871 1818 1886
rect 1842 1883 1843 1887
rect 1847 1883 1848 1887
rect 1870 1887 1871 1891
rect 1875 1887 1876 1891
rect 1870 1886 1876 1887
rect 1926 1891 1932 1892
rect 1926 1887 1927 1891
rect 1931 1887 1932 1891
rect 1960 1888 1962 1926
rect 1999 1925 2003 1926
rect 2023 1930 2027 1931
rect 2023 1925 2027 1926
rect 2055 1930 2059 1931
rect 2055 1925 2059 1926
rect 2103 1930 2107 1931
rect 2103 1925 2107 1926
rect 2119 1930 2123 1931
rect 2134 1927 2135 1931
rect 2139 1927 2140 1931
rect 2134 1926 2140 1927
rect 2583 1930 2587 1931
rect 2119 1925 2123 1926
rect 2000 1919 2002 1925
rect 2030 1923 2036 1924
rect 2030 1919 2031 1923
rect 2035 1919 2036 1923
rect 2056 1919 2058 1925
rect 2120 1919 2122 1925
rect 1998 1918 2004 1919
rect 2030 1918 2036 1919
rect 2054 1918 2060 1919
rect 1998 1914 1999 1918
rect 2003 1914 2004 1918
rect 1998 1913 2004 1914
rect 1982 1891 1988 1892
rect 1926 1886 1932 1887
rect 1958 1887 1964 1888
rect 1842 1882 1848 1883
rect 1872 1871 1874 1886
rect 1928 1871 1930 1886
rect 1958 1883 1959 1887
rect 1963 1883 1964 1887
rect 1982 1887 1983 1891
rect 1987 1887 1988 1891
rect 1982 1886 1988 1887
rect 1958 1882 1964 1883
rect 1984 1871 1986 1886
rect 1815 1870 1819 1871
rect 1815 1865 1819 1866
rect 1831 1870 1835 1871
rect 1831 1865 1835 1866
rect 1871 1870 1875 1871
rect 1871 1865 1875 1866
rect 1919 1870 1923 1871
rect 1919 1865 1923 1866
rect 1927 1870 1931 1871
rect 1927 1865 1931 1866
rect 1983 1870 1987 1871
rect 1983 1865 1987 1866
rect 2007 1870 2011 1871
rect 2007 1865 2011 1866
rect 1832 1854 1834 1865
rect 1910 1855 1916 1856
rect 1830 1853 1836 1854
rect 1830 1849 1831 1853
rect 1835 1849 1836 1853
rect 1910 1851 1911 1855
rect 1915 1851 1916 1855
rect 1920 1854 1922 1865
rect 1998 1855 2004 1856
rect 1910 1850 1916 1851
rect 1918 1853 1924 1854
rect 1830 1848 1836 1849
rect 1827 1828 1831 1829
rect 1827 1823 1831 1824
rect 1846 1826 1852 1827
rect 1828 1820 1830 1823
rect 1846 1822 1847 1826
rect 1851 1822 1852 1826
rect 1846 1821 1852 1822
rect 1782 1819 1788 1820
rect 1782 1815 1783 1819
rect 1787 1815 1788 1819
rect 1735 1814 1739 1815
rect 1735 1809 1739 1810
rect 1759 1814 1763 1815
rect 1782 1814 1788 1815
rect 1826 1819 1832 1820
rect 1826 1815 1827 1819
rect 1831 1815 1832 1819
rect 1848 1815 1850 1821
rect 1912 1820 1914 1850
rect 1918 1849 1919 1853
rect 1923 1849 1924 1853
rect 1998 1851 1999 1855
rect 2003 1851 2004 1855
rect 2008 1854 2010 1865
rect 2032 1856 2034 1918
rect 2054 1914 2055 1918
rect 2059 1914 2060 1918
rect 2054 1913 2060 1914
rect 2118 1918 2124 1919
rect 2118 1914 2119 1918
rect 2123 1914 2124 1918
rect 2118 1913 2124 1914
rect 2038 1891 2044 1892
rect 2038 1887 2039 1891
rect 2043 1887 2044 1891
rect 2038 1886 2044 1887
rect 2102 1891 2108 1892
rect 2102 1887 2103 1891
rect 2107 1887 2108 1891
rect 2136 1888 2138 1926
rect 2583 1925 2587 1926
rect 2584 1910 2586 1925
rect 2582 1909 2588 1910
rect 2582 1905 2583 1909
rect 2587 1905 2588 1909
rect 2582 1904 2588 1905
rect 2582 1892 2588 1893
rect 2582 1888 2583 1892
rect 2587 1888 2588 1892
rect 2102 1886 2108 1887
rect 2134 1887 2140 1888
rect 2582 1887 2588 1888
rect 2040 1871 2042 1886
rect 2104 1871 2106 1886
rect 2134 1883 2135 1887
rect 2139 1883 2140 1887
rect 2134 1882 2140 1883
rect 2584 1871 2586 1887
rect 2039 1870 2043 1871
rect 2039 1865 2043 1866
rect 2095 1870 2099 1871
rect 2095 1865 2099 1866
rect 2103 1870 2107 1871
rect 2103 1865 2107 1866
rect 2183 1870 2187 1871
rect 2183 1865 2187 1866
rect 2583 1870 2587 1871
rect 2583 1865 2587 1866
rect 2030 1855 2036 1856
rect 1998 1850 2004 1851
rect 2006 1853 2012 1854
rect 1918 1848 1924 1849
rect 1934 1826 1940 1827
rect 1934 1822 1935 1826
rect 1939 1822 1940 1826
rect 1934 1821 1940 1822
rect 1910 1819 1916 1820
rect 1910 1815 1911 1819
rect 1915 1815 1916 1819
rect 1936 1815 1938 1821
rect 2000 1820 2002 1850
rect 2006 1849 2007 1853
rect 2011 1849 2012 1853
rect 2030 1851 2031 1855
rect 2035 1851 2036 1855
rect 2096 1854 2098 1865
rect 2174 1855 2180 1856
rect 2030 1850 2036 1851
rect 2094 1853 2100 1854
rect 2006 1848 2012 1849
rect 2094 1849 2095 1853
rect 2099 1849 2100 1853
rect 2174 1851 2175 1855
rect 2179 1851 2180 1855
rect 2184 1854 2186 1865
rect 2206 1855 2212 1856
rect 2174 1850 2180 1851
rect 2182 1853 2188 1854
rect 2094 1848 2100 1849
rect 2022 1826 2028 1827
rect 2022 1822 2023 1826
rect 2027 1822 2028 1826
rect 2022 1821 2028 1822
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2110 1821 2116 1822
rect 1998 1819 2004 1820
rect 1998 1815 1999 1819
rect 2003 1815 2004 1819
rect 2024 1815 2026 1821
rect 2082 1819 2088 1820
rect 2082 1815 2083 1819
rect 2087 1815 2088 1819
rect 2112 1815 2114 1821
rect 2176 1820 2178 1850
rect 2182 1849 2183 1853
rect 2187 1849 2188 1853
rect 2206 1851 2207 1855
rect 2211 1851 2212 1855
rect 2584 1853 2586 1865
rect 2206 1850 2212 1851
rect 2582 1852 2588 1853
rect 2182 1848 2188 1849
rect 2208 1829 2210 1850
rect 2582 1848 2583 1852
rect 2587 1848 2588 1852
rect 2582 1847 2588 1848
rect 2582 1835 2588 1836
rect 2582 1831 2583 1835
rect 2587 1831 2588 1835
rect 2582 1830 2588 1831
rect 2207 1828 2211 1829
rect 2198 1826 2204 1827
rect 2198 1822 2199 1826
rect 2203 1822 2204 1826
rect 2207 1823 2211 1824
rect 2198 1821 2204 1822
rect 2174 1819 2180 1820
rect 2174 1815 2175 1819
rect 2179 1815 2180 1819
rect 2200 1815 2202 1821
rect 2584 1815 2586 1830
rect 1826 1814 1832 1815
rect 1839 1814 1843 1815
rect 1759 1809 1763 1810
rect 1839 1809 1843 1810
rect 1847 1814 1851 1815
rect 1910 1814 1916 1815
rect 1935 1814 1939 1815
rect 1847 1809 1851 1810
rect 1935 1809 1939 1810
rect 1951 1814 1955 1815
rect 1998 1814 2004 1815
rect 2023 1814 2027 1815
rect 1951 1809 1955 1810
rect 2023 1809 2027 1810
rect 2063 1814 2067 1815
rect 2082 1814 2088 1815
rect 2111 1814 2115 1815
rect 2174 1814 2180 1815
rect 2183 1814 2187 1815
rect 2063 1809 2067 1810
rect 1714 1807 1720 1808
rect 1714 1803 1715 1807
rect 1719 1803 1720 1807
rect 1736 1803 1738 1809
rect 1840 1803 1842 1809
rect 1926 1807 1932 1808
rect 1926 1803 1927 1807
rect 1931 1803 1932 1807
rect 1952 1803 1954 1809
rect 1970 1807 1976 1808
rect 1970 1803 1971 1807
rect 1975 1803 1976 1807
rect 2064 1803 2066 1809
rect 1714 1802 1720 1803
rect 1734 1802 1740 1803
rect 1734 1798 1735 1802
rect 1739 1798 1740 1802
rect 1734 1797 1740 1798
rect 1838 1802 1844 1803
rect 1926 1802 1932 1803
rect 1950 1802 1956 1803
rect 1970 1802 1976 1803
rect 2062 1802 2068 1803
rect 1838 1798 1839 1802
rect 1843 1798 1844 1802
rect 1838 1797 1844 1798
rect 1928 1784 1930 1802
rect 1950 1798 1951 1802
rect 1955 1798 1956 1802
rect 1950 1797 1956 1798
rect 1926 1783 1932 1784
rect 1926 1779 1927 1783
rect 1931 1779 1932 1783
rect 1926 1778 1932 1779
rect 1718 1775 1724 1776
rect 1606 1770 1612 1771
rect 1642 1771 1648 1772
rect 1530 1766 1536 1767
rect 1608 1759 1610 1770
rect 1642 1767 1643 1771
rect 1647 1767 1648 1771
rect 1718 1771 1719 1775
rect 1723 1771 1724 1775
rect 1718 1770 1724 1771
rect 1822 1775 1828 1776
rect 1822 1771 1823 1775
rect 1827 1771 1828 1775
rect 1934 1775 1940 1776
rect 1822 1770 1828 1771
rect 1918 1771 1924 1772
rect 1642 1766 1648 1767
rect 1720 1759 1722 1770
rect 1824 1759 1826 1770
rect 1918 1767 1919 1771
rect 1923 1767 1924 1771
rect 1934 1771 1935 1775
rect 1939 1771 1940 1775
rect 1972 1772 1974 1802
rect 2062 1798 2063 1802
rect 2067 1798 2068 1802
rect 2062 1797 2068 1798
rect 2046 1775 2052 1776
rect 1934 1770 1940 1771
rect 1970 1771 1976 1772
rect 1918 1766 1924 1767
rect 1439 1758 1443 1759
rect 1439 1753 1443 1754
rect 1495 1758 1499 1759
rect 1495 1753 1499 1754
rect 1519 1758 1523 1759
rect 1519 1753 1523 1754
rect 1607 1758 1611 1759
rect 1607 1753 1611 1754
rect 1615 1758 1619 1759
rect 1615 1753 1619 1754
rect 1719 1758 1723 1759
rect 1719 1753 1723 1754
rect 1823 1758 1827 1759
rect 1823 1753 1827 1754
rect 1406 1747 1412 1748
rect 1406 1743 1407 1747
rect 1411 1743 1412 1747
rect 1406 1742 1412 1743
rect 1440 1742 1442 1753
rect 1520 1742 1522 1753
rect 1616 1742 1618 1753
rect 1720 1742 1722 1753
rect 1774 1747 1780 1748
rect 1774 1743 1775 1747
rect 1779 1743 1780 1747
rect 1774 1742 1780 1743
rect 1824 1742 1826 1753
rect 1438 1741 1444 1742
rect 1366 1740 1372 1741
rect 919 1738 923 1739
rect 919 1733 923 1734
rect 935 1738 939 1739
rect 935 1733 939 1734
rect 1015 1738 1019 1739
rect 1015 1733 1019 1734
rect 1103 1738 1107 1739
rect 1103 1733 1107 1734
rect 1111 1738 1115 1739
rect 1111 1733 1115 1734
rect 1207 1738 1211 1739
rect 1207 1733 1211 1734
rect 1327 1738 1331 1739
rect 1366 1736 1367 1740
rect 1371 1736 1372 1740
rect 1438 1737 1439 1741
rect 1443 1737 1444 1741
rect 1438 1736 1444 1737
rect 1518 1741 1524 1742
rect 1518 1737 1519 1741
rect 1523 1737 1524 1741
rect 1518 1736 1524 1737
rect 1614 1741 1620 1742
rect 1614 1737 1615 1741
rect 1619 1737 1620 1741
rect 1614 1736 1620 1737
rect 1718 1741 1724 1742
rect 1718 1737 1719 1741
rect 1723 1737 1724 1741
rect 1718 1736 1724 1737
rect 1366 1735 1372 1736
rect 1327 1733 1331 1734
rect 862 1731 868 1732
rect 862 1727 863 1731
rect 867 1727 868 1731
rect 862 1726 868 1727
rect 920 1722 922 1733
rect 1016 1722 1018 1733
rect 1102 1723 1108 1724
rect 582 1718 588 1719
rect 638 1721 644 1722
rect 550 1716 556 1717
rect 566 1694 572 1695
rect 566 1690 567 1694
rect 571 1690 572 1694
rect 566 1689 572 1690
rect 542 1687 548 1688
rect 542 1683 543 1687
rect 547 1683 548 1687
rect 542 1682 548 1683
rect 568 1679 570 1689
rect 584 1680 586 1718
rect 638 1717 639 1721
rect 643 1717 644 1721
rect 638 1716 644 1717
rect 726 1721 732 1722
rect 726 1717 727 1721
rect 731 1717 732 1721
rect 726 1716 732 1717
rect 822 1721 828 1722
rect 822 1717 823 1721
rect 827 1717 828 1721
rect 822 1716 828 1717
rect 918 1721 924 1722
rect 918 1717 919 1721
rect 923 1717 924 1721
rect 918 1716 924 1717
rect 1014 1721 1020 1722
rect 1014 1717 1015 1721
rect 1019 1717 1020 1721
rect 1102 1719 1103 1723
rect 1107 1719 1108 1723
rect 1112 1722 1114 1733
rect 1198 1723 1204 1724
rect 1102 1718 1108 1719
rect 1110 1721 1116 1722
rect 1014 1716 1020 1717
rect 654 1694 660 1695
rect 654 1690 655 1694
rect 659 1690 660 1694
rect 654 1689 660 1690
rect 742 1694 748 1695
rect 742 1690 743 1694
rect 747 1690 748 1694
rect 742 1689 748 1690
rect 838 1694 844 1695
rect 838 1690 839 1694
rect 843 1690 844 1694
rect 838 1689 844 1690
rect 934 1694 940 1695
rect 934 1690 935 1694
rect 939 1690 940 1694
rect 934 1689 940 1690
rect 1030 1694 1036 1695
rect 1030 1690 1031 1694
rect 1035 1690 1036 1694
rect 1030 1689 1036 1690
rect 582 1679 588 1680
rect 656 1679 658 1689
rect 744 1679 746 1689
rect 818 1687 824 1688
rect 818 1683 819 1687
rect 823 1683 824 1687
rect 818 1682 824 1683
rect 111 1678 115 1679
rect 111 1673 115 1674
rect 367 1678 371 1679
rect 367 1673 371 1674
rect 399 1678 403 1679
rect 399 1673 403 1674
rect 423 1678 427 1679
rect 423 1673 427 1674
rect 455 1678 459 1679
rect 455 1673 459 1674
rect 487 1678 491 1679
rect 487 1673 491 1674
rect 511 1678 515 1679
rect 511 1673 515 1674
rect 567 1678 571 1679
rect 567 1673 571 1674
rect 575 1678 579 1679
rect 582 1675 583 1679
rect 587 1675 588 1679
rect 582 1674 588 1675
rect 647 1678 651 1679
rect 575 1673 579 1674
rect 647 1673 651 1674
rect 655 1678 659 1679
rect 655 1673 659 1674
rect 727 1678 731 1679
rect 727 1673 731 1674
rect 743 1678 747 1679
rect 743 1673 747 1674
rect 807 1678 811 1679
rect 807 1673 811 1674
rect 112 1658 114 1673
rect 400 1667 402 1673
rect 456 1667 458 1673
rect 470 1671 476 1672
rect 470 1667 471 1671
rect 475 1667 476 1671
rect 512 1667 514 1673
rect 530 1671 536 1672
rect 530 1667 531 1671
rect 535 1667 536 1671
rect 576 1667 578 1673
rect 594 1671 600 1672
rect 594 1667 595 1671
rect 599 1667 600 1671
rect 648 1667 650 1673
rect 666 1671 672 1672
rect 666 1667 667 1671
rect 671 1667 672 1671
rect 728 1667 730 1673
rect 766 1671 772 1672
rect 766 1667 767 1671
rect 771 1667 772 1671
rect 808 1667 810 1673
rect 398 1666 404 1667
rect 398 1662 399 1666
rect 403 1662 404 1666
rect 398 1661 404 1662
rect 454 1666 460 1667
rect 470 1666 476 1667
rect 510 1666 516 1667
rect 530 1666 536 1667
rect 574 1666 580 1667
rect 594 1666 600 1667
rect 646 1666 652 1667
rect 666 1666 672 1667
rect 726 1666 732 1667
rect 766 1666 772 1667
rect 806 1666 812 1667
rect 454 1662 455 1666
rect 459 1662 460 1666
rect 454 1661 460 1662
rect 110 1657 116 1658
rect 110 1653 111 1657
rect 115 1653 116 1657
rect 110 1652 116 1653
rect 110 1640 116 1641
rect 110 1636 111 1640
rect 115 1636 116 1640
rect 110 1635 116 1636
rect 382 1639 388 1640
rect 382 1635 383 1639
rect 387 1635 388 1639
rect 112 1607 114 1635
rect 382 1634 388 1635
rect 438 1639 444 1640
rect 438 1635 439 1639
rect 443 1635 444 1639
rect 472 1636 474 1666
rect 510 1662 511 1666
rect 515 1662 516 1666
rect 510 1661 516 1662
rect 494 1639 500 1640
rect 438 1634 444 1635
rect 470 1635 476 1636
rect 384 1607 386 1634
rect 440 1607 442 1634
rect 470 1631 471 1635
rect 475 1631 476 1635
rect 494 1635 495 1639
rect 499 1635 500 1639
rect 532 1636 534 1666
rect 574 1662 575 1666
rect 579 1662 580 1666
rect 574 1661 580 1662
rect 558 1639 564 1640
rect 494 1634 500 1635
rect 530 1635 536 1636
rect 470 1630 476 1631
rect 496 1607 498 1634
rect 530 1631 531 1635
rect 535 1631 536 1635
rect 558 1635 559 1639
rect 563 1635 564 1639
rect 596 1636 598 1666
rect 646 1662 647 1666
rect 651 1662 652 1666
rect 646 1661 652 1662
rect 630 1639 636 1640
rect 558 1634 564 1635
rect 594 1635 600 1636
rect 530 1630 536 1631
rect 560 1607 562 1634
rect 594 1631 595 1635
rect 599 1631 600 1635
rect 630 1635 631 1639
rect 635 1635 636 1639
rect 668 1636 670 1666
rect 726 1662 727 1666
rect 731 1662 732 1666
rect 726 1661 732 1662
rect 768 1640 770 1666
rect 806 1662 807 1666
rect 811 1662 812 1666
rect 806 1661 812 1662
rect 710 1639 716 1640
rect 630 1634 636 1635
rect 666 1635 672 1636
rect 594 1630 600 1631
rect 632 1607 634 1634
rect 666 1631 667 1635
rect 671 1631 672 1635
rect 710 1635 711 1639
rect 715 1635 716 1639
rect 710 1634 716 1635
rect 766 1639 772 1640
rect 766 1635 767 1639
rect 771 1635 772 1639
rect 766 1634 772 1635
rect 790 1639 796 1640
rect 790 1635 791 1639
rect 795 1635 796 1639
rect 820 1636 822 1682
rect 840 1679 842 1689
rect 936 1679 938 1689
rect 982 1687 988 1688
rect 982 1683 983 1687
rect 987 1683 988 1687
rect 982 1682 988 1683
rect 839 1678 843 1679
rect 839 1673 843 1674
rect 887 1678 891 1679
rect 887 1673 891 1674
rect 935 1678 939 1679
rect 935 1673 939 1674
rect 967 1678 971 1679
rect 967 1673 971 1674
rect 854 1671 860 1672
rect 854 1667 855 1671
rect 859 1667 860 1671
rect 888 1667 890 1673
rect 968 1667 970 1673
rect 854 1666 860 1667
rect 886 1666 892 1667
rect 790 1634 796 1635
rect 818 1635 824 1636
rect 666 1630 672 1631
rect 712 1607 714 1634
rect 792 1607 794 1634
rect 818 1631 819 1635
rect 823 1631 824 1635
rect 818 1630 824 1631
rect 111 1606 115 1607
rect 111 1601 115 1602
rect 287 1606 291 1607
rect 287 1601 291 1602
rect 367 1606 371 1607
rect 367 1601 371 1602
rect 383 1606 387 1607
rect 383 1601 387 1602
rect 439 1606 443 1607
rect 439 1601 443 1602
rect 455 1606 459 1607
rect 455 1601 459 1602
rect 495 1606 499 1607
rect 495 1601 499 1602
rect 551 1606 555 1607
rect 551 1601 555 1602
rect 559 1606 563 1607
rect 559 1601 563 1602
rect 631 1606 635 1607
rect 631 1601 635 1602
rect 647 1606 651 1607
rect 647 1601 651 1602
rect 711 1606 715 1607
rect 711 1601 715 1602
rect 735 1606 739 1607
rect 735 1601 739 1602
rect 791 1606 795 1607
rect 791 1601 795 1602
rect 823 1606 827 1607
rect 823 1601 827 1602
rect 112 1589 114 1601
rect 288 1590 290 1601
rect 358 1591 364 1592
rect 286 1589 292 1590
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 286 1585 287 1589
rect 291 1585 292 1589
rect 358 1587 359 1591
rect 363 1587 364 1591
rect 368 1590 370 1601
rect 446 1591 452 1592
rect 358 1586 364 1587
rect 366 1589 372 1590
rect 286 1584 292 1585
rect 110 1583 116 1584
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 110 1566 116 1567
rect 112 1551 114 1566
rect 302 1562 308 1563
rect 302 1558 303 1562
rect 307 1558 308 1562
rect 302 1557 308 1558
rect 294 1555 300 1556
rect 294 1551 295 1555
rect 299 1551 300 1555
rect 304 1551 306 1557
rect 360 1556 362 1586
rect 366 1585 367 1589
rect 371 1585 372 1589
rect 446 1587 447 1591
rect 451 1587 452 1591
rect 456 1590 458 1601
rect 534 1591 540 1592
rect 446 1586 452 1587
rect 454 1589 460 1590
rect 366 1584 372 1585
rect 382 1562 388 1563
rect 382 1558 383 1562
rect 387 1558 388 1562
rect 382 1557 388 1558
rect 358 1555 364 1556
rect 358 1551 359 1555
rect 363 1551 364 1555
rect 384 1551 386 1557
rect 448 1556 450 1586
rect 454 1585 455 1589
rect 459 1585 460 1589
rect 534 1587 535 1591
rect 539 1587 540 1591
rect 552 1590 554 1601
rect 638 1591 644 1592
rect 534 1586 540 1587
rect 550 1589 556 1590
rect 454 1584 460 1585
rect 470 1562 476 1563
rect 470 1558 471 1562
rect 475 1558 476 1562
rect 470 1557 476 1558
rect 446 1555 452 1556
rect 414 1551 420 1552
rect 111 1550 115 1551
rect 111 1545 115 1546
rect 279 1550 283 1551
rect 294 1550 300 1551
rect 303 1550 307 1551
rect 279 1545 283 1546
rect 112 1530 114 1545
rect 254 1543 260 1544
rect 254 1539 255 1543
rect 259 1539 260 1543
rect 280 1539 282 1545
rect 254 1538 260 1539
rect 278 1538 284 1539
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 256 1520 258 1538
rect 278 1534 279 1538
rect 283 1534 284 1538
rect 278 1533 284 1534
rect 254 1519 260 1520
rect 254 1515 255 1519
rect 259 1515 260 1519
rect 254 1514 260 1515
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 262 1511 268 1512
rect 262 1507 263 1511
rect 267 1507 268 1511
rect 296 1508 298 1550
rect 303 1545 307 1546
rect 335 1550 339 1551
rect 358 1550 364 1551
rect 383 1550 387 1551
rect 335 1545 339 1546
rect 383 1545 387 1546
rect 399 1550 403 1551
rect 414 1547 415 1551
rect 419 1547 420 1551
rect 446 1551 447 1555
rect 451 1551 452 1555
rect 472 1551 474 1557
rect 536 1556 538 1586
rect 550 1585 551 1589
rect 555 1585 556 1589
rect 638 1587 639 1591
rect 643 1587 644 1591
rect 648 1590 650 1601
rect 670 1591 676 1592
rect 638 1586 644 1587
rect 646 1589 652 1590
rect 550 1584 556 1585
rect 566 1562 572 1563
rect 566 1558 567 1562
rect 571 1558 572 1562
rect 566 1557 572 1558
rect 534 1555 540 1556
rect 534 1551 535 1555
rect 539 1551 540 1555
rect 568 1551 570 1557
rect 640 1556 642 1586
rect 646 1585 647 1589
rect 651 1585 652 1589
rect 670 1587 671 1591
rect 675 1587 676 1591
rect 736 1590 738 1601
rect 814 1591 820 1592
rect 670 1586 676 1587
rect 734 1589 740 1590
rect 646 1584 652 1585
rect 662 1562 668 1563
rect 662 1558 663 1562
rect 667 1558 668 1562
rect 662 1557 668 1558
rect 638 1555 644 1556
rect 638 1551 639 1555
rect 643 1551 644 1555
rect 664 1551 666 1557
rect 672 1552 674 1586
rect 734 1585 735 1589
rect 739 1585 740 1589
rect 814 1587 815 1591
rect 819 1587 820 1591
rect 824 1590 826 1601
rect 856 1592 858 1666
rect 886 1662 887 1666
rect 891 1662 892 1666
rect 886 1661 892 1662
rect 966 1666 972 1667
rect 966 1662 967 1666
rect 971 1662 972 1666
rect 966 1661 972 1662
rect 870 1639 876 1640
rect 870 1635 871 1639
rect 875 1635 876 1639
rect 870 1634 876 1635
rect 950 1639 956 1640
rect 950 1635 951 1639
rect 955 1635 956 1639
rect 984 1636 986 1682
rect 1032 1679 1034 1689
rect 1104 1688 1106 1718
rect 1110 1717 1111 1721
rect 1115 1717 1116 1721
rect 1198 1719 1199 1723
rect 1203 1719 1204 1723
rect 1208 1722 1210 1733
rect 1230 1723 1236 1724
rect 1198 1718 1204 1719
rect 1206 1721 1212 1722
rect 1110 1716 1116 1717
rect 1126 1694 1132 1695
rect 1126 1690 1127 1694
rect 1131 1690 1132 1694
rect 1126 1689 1132 1690
rect 1102 1687 1108 1688
rect 1102 1683 1103 1687
rect 1107 1683 1108 1687
rect 1102 1682 1108 1683
rect 1128 1679 1130 1689
rect 1200 1688 1202 1718
rect 1206 1717 1207 1721
rect 1211 1717 1212 1721
rect 1230 1719 1231 1723
rect 1235 1719 1236 1723
rect 1328 1721 1330 1733
rect 1366 1723 1372 1724
rect 1230 1718 1236 1719
rect 1326 1720 1332 1721
rect 1206 1716 1212 1717
rect 1222 1694 1228 1695
rect 1222 1690 1223 1694
rect 1227 1690 1228 1694
rect 1222 1689 1228 1690
rect 1198 1687 1204 1688
rect 1198 1683 1199 1687
rect 1203 1683 1204 1687
rect 1198 1682 1204 1683
rect 1224 1679 1226 1689
rect 1031 1678 1035 1679
rect 1031 1673 1035 1674
rect 1047 1678 1051 1679
rect 1047 1673 1051 1674
rect 1127 1678 1131 1679
rect 1127 1673 1131 1674
rect 1135 1678 1139 1679
rect 1135 1673 1139 1674
rect 1223 1678 1227 1679
rect 1232 1676 1234 1718
rect 1326 1716 1327 1720
rect 1331 1716 1332 1720
rect 1366 1719 1367 1723
rect 1371 1719 1372 1723
rect 1366 1718 1372 1719
rect 1326 1715 1332 1716
rect 1326 1703 1332 1704
rect 1326 1699 1327 1703
rect 1331 1699 1332 1703
rect 1326 1698 1332 1699
rect 1328 1679 1330 1698
rect 1368 1691 1370 1718
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1534 1714 1540 1715
rect 1534 1710 1535 1714
rect 1539 1710 1540 1714
rect 1534 1709 1540 1710
rect 1630 1714 1636 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 1734 1714 1740 1715
rect 1734 1710 1735 1714
rect 1739 1710 1740 1714
rect 1734 1709 1740 1710
rect 1456 1691 1458 1709
rect 1536 1691 1538 1709
rect 1632 1691 1634 1709
rect 1722 1707 1728 1708
rect 1722 1703 1723 1707
rect 1727 1703 1728 1707
rect 1722 1702 1728 1703
rect 1367 1690 1371 1691
rect 1367 1685 1371 1686
rect 1455 1690 1459 1691
rect 1455 1685 1459 1686
rect 1535 1690 1539 1691
rect 1535 1685 1539 1686
rect 1559 1690 1563 1691
rect 1559 1685 1563 1686
rect 1631 1690 1635 1691
rect 1631 1685 1635 1686
rect 1711 1690 1715 1691
rect 1711 1685 1715 1686
rect 1287 1678 1291 1679
rect 1223 1673 1227 1674
rect 1230 1675 1236 1676
rect 1022 1671 1028 1672
rect 1022 1667 1023 1671
rect 1027 1667 1028 1671
rect 1048 1667 1050 1673
rect 1066 1671 1072 1672
rect 1066 1667 1067 1671
rect 1071 1667 1072 1671
rect 1136 1667 1138 1673
rect 1224 1667 1226 1673
rect 1230 1671 1231 1675
rect 1235 1671 1236 1675
rect 1287 1673 1291 1674
rect 1327 1678 1331 1679
rect 1327 1673 1331 1674
rect 1230 1670 1236 1671
rect 1242 1671 1248 1672
rect 1242 1667 1243 1671
rect 1247 1667 1248 1671
rect 1288 1667 1290 1673
rect 1022 1666 1028 1667
rect 1046 1666 1052 1667
rect 1066 1666 1072 1667
rect 1134 1666 1140 1667
rect 1024 1648 1026 1666
rect 1046 1662 1047 1666
rect 1051 1662 1052 1666
rect 1046 1661 1052 1662
rect 1022 1647 1028 1648
rect 1022 1643 1023 1647
rect 1027 1643 1028 1647
rect 1022 1642 1028 1643
rect 1030 1639 1036 1640
rect 950 1634 956 1635
rect 982 1635 988 1636
rect 872 1607 874 1634
rect 952 1607 954 1634
rect 982 1631 983 1635
rect 987 1631 988 1635
rect 1030 1635 1031 1639
rect 1035 1635 1036 1639
rect 1068 1636 1070 1666
rect 1134 1662 1135 1666
rect 1139 1662 1140 1666
rect 1134 1661 1140 1662
rect 1222 1666 1228 1667
rect 1242 1666 1248 1667
rect 1286 1666 1292 1667
rect 1222 1662 1223 1666
rect 1227 1662 1228 1666
rect 1222 1661 1228 1662
rect 1118 1639 1124 1640
rect 1030 1634 1036 1635
rect 1066 1635 1072 1636
rect 982 1630 988 1631
rect 1032 1607 1034 1634
rect 1066 1631 1067 1635
rect 1071 1631 1072 1635
rect 1118 1635 1119 1639
rect 1123 1635 1124 1639
rect 1206 1639 1212 1640
rect 1118 1634 1124 1635
rect 1142 1635 1148 1636
rect 1066 1630 1072 1631
rect 1120 1607 1122 1634
rect 1142 1631 1143 1635
rect 1147 1631 1148 1635
rect 1206 1635 1207 1639
rect 1211 1635 1212 1639
rect 1244 1636 1246 1666
rect 1286 1662 1287 1666
rect 1291 1662 1292 1666
rect 1286 1661 1292 1662
rect 1328 1658 1330 1673
rect 1368 1670 1370 1685
rect 1550 1683 1556 1684
rect 1550 1679 1551 1683
rect 1555 1679 1556 1683
rect 1560 1679 1562 1685
rect 1578 1683 1584 1684
rect 1578 1679 1579 1683
rect 1583 1679 1584 1683
rect 1632 1679 1634 1685
rect 1650 1683 1656 1684
rect 1650 1679 1651 1683
rect 1655 1679 1656 1683
rect 1712 1679 1714 1685
rect 1550 1678 1556 1679
rect 1558 1678 1564 1679
rect 1578 1678 1584 1679
rect 1630 1678 1636 1679
rect 1650 1678 1656 1679
rect 1710 1678 1716 1679
rect 1366 1669 1372 1670
rect 1366 1665 1367 1669
rect 1371 1665 1372 1669
rect 1366 1664 1372 1665
rect 1326 1657 1332 1658
rect 1326 1653 1327 1657
rect 1331 1653 1332 1657
rect 1326 1652 1332 1653
rect 1366 1652 1372 1653
rect 1366 1648 1367 1652
rect 1371 1648 1372 1652
rect 1366 1647 1372 1648
rect 1542 1651 1548 1652
rect 1542 1647 1543 1651
rect 1547 1647 1548 1651
rect 1326 1640 1332 1641
rect 1270 1639 1276 1640
rect 1206 1634 1212 1635
rect 1242 1635 1248 1636
rect 1142 1630 1148 1631
rect 871 1606 875 1607
rect 871 1601 875 1602
rect 903 1606 907 1607
rect 903 1601 907 1602
rect 951 1606 955 1607
rect 951 1601 955 1602
rect 983 1606 987 1607
rect 983 1601 987 1602
rect 1031 1606 1035 1607
rect 1031 1601 1035 1602
rect 1063 1606 1067 1607
rect 1063 1601 1067 1602
rect 1119 1606 1123 1607
rect 1119 1601 1123 1602
rect 854 1591 860 1592
rect 814 1586 820 1587
rect 822 1589 828 1590
rect 734 1584 740 1585
rect 750 1562 756 1563
rect 750 1558 751 1562
rect 755 1558 756 1562
rect 750 1557 756 1558
rect 706 1555 712 1556
rect 670 1551 676 1552
rect 706 1551 707 1555
rect 711 1551 712 1555
rect 752 1551 754 1557
rect 816 1556 818 1586
rect 822 1585 823 1589
rect 827 1585 828 1589
rect 854 1587 855 1591
rect 859 1587 860 1591
rect 904 1590 906 1601
rect 910 1599 916 1600
rect 910 1595 911 1599
rect 915 1595 916 1599
rect 910 1594 916 1595
rect 854 1586 860 1587
rect 902 1589 908 1590
rect 822 1584 828 1585
rect 902 1585 903 1589
rect 907 1585 908 1589
rect 902 1584 908 1585
rect 838 1562 844 1563
rect 838 1558 839 1562
rect 843 1558 844 1562
rect 838 1557 844 1558
rect 814 1555 820 1556
rect 814 1551 815 1555
rect 819 1551 820 1555
rect 840 1551 842 1557
rect 912 1556 914 1594
rect 984 1590 986 1601
rect 1030 1591 1036 1592
rect 982 1589 988 1590
rect 982 1585 983 1589
rect 987 1585 988 1589
rect 1030 1587 1031 1591
rect 1035 1587 1036 1591
rect 1064 1590 1066 1601
rect 1030 1586 1036 1587
rect 1062 1589 1068 1590
rect 982 1584 988 1585
rect 918 1562 924 1563
rect 918 1558 919 1562
rect 923 1558 924 1562
rect 918 1557 924 1558
rect 998 1562 1004 1563
rect 998 1558 999 1562
rect 1003 1558 1004 1562
rect 998 1557 1004 1558
rect 910 1555 916 1556
rect 910 1551 911 1555
rect 915 1551 916 1555
rect 920 1551 922 1557
rect 1000 1551 1002 1557
rect 446 1550 452 1551
rect 471 1550 475 1551
rect 534 1550 540 1551
rect 543 1550 547 1551
rect 414 1546 420 1547
rect 399 1545 403 1546
rect 336 1539 338 1545
rect 390 1543 396 1544
rect 390 1539 391 1543
rect 395 1539 396 1543
rect 400 1539 402 1545
rect 334 1538 340 1539
rect 390 1538 396 1539
rect 398 1538 404 1539
rect 334 1534 335 1538
rect 339 1534 340 1538
rect 334 1533 340 1534
rect 318 1511 324 1512
rect 112 1491 114 1507
rect 262 1506 268 1507
rect 294 1507 300 1508
rect 264 1491 266 1506
rect 294 1503 295 1507
rect 299 1503 300 1507
rect 318 1507 319 1511
rect 323 1507 324 1511
rect 318 1506 324 1507
rect 382 1511 388 1512
rect 382 1507 383 1511
rect 387 1507 388 1511
rect 382 1506 388 1507
rect 294 1502 300 1503
rect 320 1491 322 1506
rect 384 1491 386 1506
rect 111 1490 115 1491
rect 111 1485 115 1486
rect 199 1490 203 1491
rect 199 1485 203 1486
rect 263 1490 267 1491
rect 263 1485 267 1486
rect 287 1490 291 1491
rect 287 1485 291 1486
rect 319 1490 323 1491
rect 319 1485 323 1486
rect 383 1490 387 1491
rect 383 1485 387 1486
rect 112 1473 114 1485
rect 200 1474 202 1485
rect 278 1475 284 1476
rect 198 1473 204 1474
rect 110 1472 116 1473
rect 110 1468 111 1472
rect 115 1468 116 1472
rect 198 1469 199 1473
rect 203 1469 204 1473
rect 278 1471 279 1475
rect 283 1471 284 1475
rect 288 1474 290 1485
rect 374 1475 380 1476
rect 278 1470 284 1471
rect 286 1473 292 1474
rect 198 1468 204 1469
rect 110 1467 116 1468
rect 110 1455 116 1456
rect 110 1451 111 1455
rect 115 1451 116 1455
rect 110 1450 116 1451
rect 112 1431 114 1450
rect 214 1446 220 1447
rect 214 1442 215 1446
rect 219 1442 220 1446
rect 214 1441 220 1442
rect 174 1439 180 1440
rect 174 1435 175 1439
rect 179 1435 180 1439
rect 174 1434 180 1435
rect 111 1430 115 1431
rect 111 1425 115 1426
rect 159 1430 163 1431
rect 159 1425 163 1426
rect 112 1410 114 1425
rect 134 1423 140 1424
rect 134 1419 135 1423
rect 139 1419 140 1423
rect 160 1419 162 1425
rect 134 1418 140 1419
rect 158 1418 164 1419
rect 110 1409 116 1410
rect 110 1405 111 1409
rect 115 1405 116 1409
rect 110 1404 116 1405
rect 136 1400 138 1418
rect 158 1414 159 1418
rect 163 1414 164 1418
rect 158 1413 164 1414
rect 134 1399 140 1400
rect 134 1395 135 1399
rect 139 1395 140 1399
rect 134 1394 140 1395
rect 110 1392 116 1393
rect 110 1388 111 1392
rect 115 1388 116 1392
rect 110 1387 116 1388
rect 142 1391 148 1392
rect 142 1387 143 1391
rect 147 1387 148 1391
rect 176 1388 178 1434
rect 216 1431 218 1441
rect 280 1440 282 1470
rect 286 1469 287 1473
rect 291 1469 292 1473
rect 374 1471 375 1475
rect 379 1471 380 1475
rect 384 1474 386 1485
rect 392 1480 394 1538
rect 398 1534 399 1538
rect 403 1534 404 1538
rect 398 1533 404 1534
rect 416 1508 418 1546
rect 471 1545 475 1546
rect 543 1545 547 1546
rect 567 1550 571 1551
rect 567 1545 571 1546
rect 615 1550 619 1551
rect 638 1550 644 1551
rect 663 1550 667 1551
rect 615 1545 619 1546
rect 670 1547 671 1551
rect 675 1547 676 1551
rect 670 1546 676 1547
rect 687 1550 691 1551
rect 706 1550 712 1551
rect 751 1550 755 1551
rect 663 1545 667 1546
rect 687 1545 691 1546
rect 446 1543 452 1544
rect 446 1539 447 1543
rect 451 1539 452 1543
rect 472 1539 474 1545
rect 490 1543 496 1544
rect 490 1539 491 1543
rect 495 1539 496 1543
rect 544 1539 546 1545
rect 616 1539 618 1545
rect 678 1543 684 1544
rect 678 1539 679 1543
rect 683 1539 684 1543
rect 688 1539 690 1545
rect 446 1538 452 1539
rect 470 1538 476 1539
rect 490 1538 496 1539
rect 542 1538 548 1539
rect 448 1520 450 1538
rect 470 1534 471 1538
rect 475 1534 476 1538
rect 470 1533 476 1534
rect 446 1519 452 1520
rect 446 1515 447 1519
rect 451 1515 452 1519
rect 446 1514 452 1515
rect 454 1511 460 1512
rect 414 1507 420 1508
rect 414 1503 415 1507
rect 419 1503 420 1507
rect 454 1507 455 1511
rect 459 1507 460 1511
rect 492 1508 494 1538
rect 542 1534 543 1538
rect 547 1534 548 1538
rect 542 1533 548 1534
rect 614 1538 620 1539
rect 678 1538 684 1539
rect 686 1538 692 1539
rect 614 1534 615 1538
rect 619 1534 620 1538
rect 614 1533 620 1534
rect 526 1511 532 1512
rect 454 1506 460 1507
rect 490 1507 496 1508
rect 414 1502 420 1503
rect 456 1491 458 1506
rect 490 1503 491 1507
rect 495 1503 496 1507
rect 526 1507 527 1511
rect 531 1507 532 1511
rect 598 1511 604 1512
rect 526 1506 532 1507
rect 574 1507 580 1508
rect 490 1502 496 1503
rect 528 1491 530 1506
rect 574 1503 575 1507
rect 579 1503 580 1507
rect 598 1507 599 1511
rect 603 1507 604 1511
rect 598 1506 604 1507
rect 670 1511 676 1512
rect 670 1507 671 1511
rect 675 1507 676 1511
rect 670 1506 676 1507
rect 574 1502 580 1503
rect 455 1490 459 1491
rect 455 1485 459 1486
rect 487 1490 491 1491
rect 487 1485 491 1486
rect 527 1490 531 1491
rect 527 1485 531 1486
rect 390 1479 396 1480
rect 390 1475 391 1479
rect 395 1475 396 1479
rect 390 1474 396 1475
rect 488 1474 490 1485
rect 510 1475 516 1476
rect 374 1470 380 1471
rect 382 1473 388 1474
rect 286 1468 292 1469
rect 302 1446 308 1447
rect 302 1442 303 1446
rect 307 1442 308 1446
rect 302 1441 308 1442
rect 278 1439 284 1440
rect 278 1435 279 1439
rect 283 1435 284 1439
rect 278 1434 284 1435
rect 304 1431 306 1441
rect 376 1440 378 1470
rect 382 1469 383 1473
rect 387 1469 388 1473
rect 382 1468 388 1469
rect 486 1473 492 1474
rect 486 1469 487 1473
rect 491 1469 492 1473
rect 510 1471 511 1475
rect 515 1471 516 1475
rect 510 1470 516 1471
rect 486 1468 492 1469
rect 398 1446 404 1447
rect 398 1442 399 1446
rect 403 1442 404 1446
rect 398 1441 404 1442
rect 502 1446 508 1447
rect 502 1442 503 1446
rect 507 1442 508 1446
rect 502 1441 508 1442
rect 374 1439 380 1440
rect 374 1435 375 1439
rect 379 1435 380 1439
rect 374 1434 380 1435
rect 358 1431 364 1432
rect 400 1431 402 1441
rect 504 1431 506 1441
rect 512 1432 514 1470
rect 576 1440 578 1502
rect 600 1491 602 1506
rect 672 1491 674 1506
rect 680 1500 682 1538
rect 686 1534 687 1538
rect 691 1534 692 1538
rect 686 1533 692 1534
rect 708 1508 710 1550
rect 751 1545 755 1546
rect 759 1550 763 1551
rect 814 1550 820 1551
rect 831 1550 835 1551
rect 759 1545 763 1546
rect 831 1545 835 1546
rect 839 1550 843 1551
rect 839 1545 843 1546
rect 903 1550 907 1551
rect 910 1550 916 1551
rect 919 1550 923 1551
rect 903 1545 907 1546
rect 919 1545 923 1546
rect 975 1550 979 1551
rect 975 1545 979 1546
rect 999 1550 1003 1551
rect 999 1545 1003 1546
rect 734 1543 740 1544
rect 734 1539 735 1543
rect 739 1539 740 1543
rect 760 1539 762 1545
rect 806 1543 812 1544
rect 806 1539 807 1543
rect 811 1539 812 1543
rect 832 1539 834 1545
rect 878 1543 884 1544
rect 878 1539 879 1543
rect 883 1539 884 1543
rect 904 1539 906 1545
rect 966 1543 972 1544
rect 966 1539 967 1543
rect 971 1539 972 1543
rect 976 1539 978 1545
rect 1032 1544 1034 1586
rect 1062 1585 1063 1589
rect 1067 1585 1068 1589
rect 1062 1584 1068 1585
rect 1078 1562 1084 1563
rect 1078 1558 1079 1562
rect 1083 1558 1084 1562
rect 1078 1557 1084 1558
rect 1080 1551 1082 1557
rect 1144 1556 1146 1630
rect 1208 1607 1210 1634
rect 1242 1631 1243 1635
rect 1247 1631 1248 1635
rect 1270 1635 1271 1639
rect 1275 1635 1276 1639
rect 1326 1636 1327 1640
rect 1331 1636 1332 1640
rect 1326 1635 1332 1636
rect 1270 1634 1276 1635
rect 1242 1630 1248 1631
rect 1272 1607 1274 1634
rect 1328 1607 1330 1635
rect 1368 1623 1370 1647
rect 1542 1646 1548 1647
rect 1544 1623 1546 1646
rect 1367 1622 1371 1623
rect 1367 1617 1371 1618
rect 1543 1622 1547 1623
rect 1543 1617 1547 1618
rect 1151 1606 1155 1607
rect 1151 1601 1155 1602
rect 1207 1606 1211 1607
rect 1207 1601 1211 1602
rect 1271 1606 1275 1607
rect 1271 1601 1275 1602
rect 1327 1606 1331 1607
rect 1368 1605 1370 1617
rect 1552 1612 1554 1678
rect 1558 1674 1559 1678
rect 1563 1674 1564 1678
rect 1558 1673 1564 1674
rect 1580 1648 1582 1678
rect 1630 1674 1631 1678
rect 1635 1674 1636 1678
rect 1630 1673 1636 1674
rect 1614 1651 1620 1652
rect 1578 1647 1584 1648
rect 1578 1643 1579 1647
rect 1583 1643 1584 1647
rect 1614 1647 1615 1651
rect 1619 1647 1620 1651
rect 1652 1648 1654 1678
rect 1710 1674 1711 1678
rect 1715 1674 1716 1678
rect 1710 1673 1716 1674
rect 1694 1651 1700 1652
rect 1614 1646 1620 1647
rect 1650 1647 1656 1648
rect 1578 1642 1584 1643
rect 1616 1623 1618 1646
rect 1650 1643 1651 1647
rect 1655 1643 1656 1647
rect 1694 1647 1695 1651
rect 1699 1647 1700 1651
rect 1724 1648 1726 1702
rect 1736 1691 1738 1709
rect 1735 1690 1739 1691
rect 1735 1685 1739 1686
rect 1776 1684 1778 1742
rect 1822 1741 1828 1742
rect 1822 1737 1823 1741
rect 1827 1737 1828 1741
rect 1822 1736 1828 1737
rect 1838 1714 1844 1715
rect 1838 1710 1839 1714
rect 1843 1710 1844 1714
rect 1838 1709 1844 1710
rect 1840 1691 1842 1709
rect 1920 1708 1922 1766
rect 1936 1759 1938 1770
rect 1970 1767 1971 1771
rect 1975 1767 1976 1771
rect 2046 1771 2047 1775
rect 2051 1771 2052 1775
rect 2084 1772 2086 1814
rect 2111 1809 2115 1810
rect 2183 1809 2187 1810
rect 2199 1814 2203 1815
rect 2199 1809 2203 1810
rect 2303 1814 2307 1815
rect 2303 1809 2307 1810
rect 2431 1814 2435 1815
rect 2431 1809 2435 1810
rect 2543 1814 2547 1815
rect 2543 1809 2547 1810
rect 2583 1814 2587 1815
rect 2583 1809 2587 1810
rect 2154 1807 2160 1808
rect 2154 1803 2155 1807
rect 2159 1803 2160 1807
rect 2184 1803 2186 1809
rect 2234 1807 2240 1808
rect 2234 1803 2235 1807
rect 2239 1803 2240 1807
rect 2304 1803 2306 1809
rect 2322 1807 2328 1808
rect 2322 1803 2323 1807
rect 2327 1803 2328 1807
rect 2432 1803 2434 1809
rect 2534 1807 2540 1808
rect 2534 1803 2535 1807
rect 2539 1803 2540 1807
rect 2544 1803 2546 1809
rect 2154 1802 2160 1803
rect 2182 1802 2188 1803
rect 2234 1802 2240 1803
rect 2302 1802 2308 1803
rect 2322 1802 2328 1803
rect 2430 1802 2436 1803
rect 2534 1802 2540 1803
rect 2542 1802 2548 1803
rect 2046 1770 2052 1771
rect 2082 1771 2088 1772
rect 1970 1766 1976 1767
rect 2048 1759 2050 1770
rect 2082 1767 2083 1771
rect 2087 1767 2088 1771
rect 2082 1766 2088 1767
rect 1927 1758 1931 1759
rect 1927 1753 1931 1754
rect 1935 1758 1939 1759
rect 1935 1753 1939 1754
rect 2023 1758 2027 1759
rect 2023 1753 2027 1754
rect 2047 1758 2051 1759
rect 2047 1753 2051 1754
rect 2119 1758 2123 1759
rect 2119 1753 2123 1754
rect 1928 1742 1930 1753
rect 2024 1742 2026 1753
rect 2110 1743 2116 1744
rect 1926 1741 1932 1742
rect 1926 1737 1927 1741
rect 1931 1737 1932 1741
rect 1926 1736 1932 1737
rect 2022 1741 2028 1742
rect 2022 1737 2023 1741
rect 2027 1737 2028 1741
rect 2110 1739 2111 1743
rect 2115 1739 2116 1743
rect 2120 1742 2122 1753
rect 2156 1744 2158 1802
rect 2182 1798 2183 1802
rect 2187 1798 2188 1802
rect 2182 1797 2188 1798
rect 2166 1775 2172 1776
rect 2166 1771 2167 1775
rect 2171 1771 2172 1775
rect 2236 1772 2238 1802
rect 2302 1798 2303 1802
rect 2307 1798 2308 1802
rect 2302 1797 2308 1798
rect 2286 1775 2292 1776
rect 2166 1770 2172 1771
rect 2234 1771 2240 1772
rect 2168 1759 2170 1770
rect 2234 1767 2235 1771
rect 2239 1767 2240 1771
rect 2286 1771 2287 1775
rect 2291 1771 2292 1775
rect 2324 1772 2326 1802
rect 2430 1798 2431 1802
rect 2435 1798 2436 1802
rect 2430 1797 2436 1798
rect 2414 1775 2420 1776
rect 2286 1770 2292 1771
rect 2322 1771 2328 1772
rect 2234 1766 2240 1767
rect 2288 1759 2290 1770
rect 2322 1767 2323 1771
rect 2327 1767 2328 1771
rect 2414 1771 2415 1775
rect 2419 1771 2420 1775
rect 2414 1770 2420 1771
rect 2526 1775 2532 1776
rect 2526 1771 2527 1775
rect 2531 1771 2532 1775
rect 2526 1770 2532 1771
rect 2322 1766 2328 1767
rect 2416 1759 2418 1770
rect 2470 1767 2476 1768
rect 2470 1763 2471 1767
rect 2475 1763 2476 1767
rect 2470 1762 2476 1763
rect 2167 1758 2171 1759
rect 2167 1753 2171 1754
rect 2207 1758 2211 1759
rect 2207 1753 2211 1754
rect 2287 1758 2291 1759
rect 2287 1753 2291 1754
rect 2375 1758 2379 1759
rect 2375 1753 2379 1754
rect 2415 1758 2419 1759
rect 2415 1753 2419 1754
rect 2463 1758 2467 1759
rect 2463 1753 2467 1754
rect 2154 1743 2160 1744
rect 2110 1738 2116 1739
rect 2118 1741 2124 1742
rect 2022 1736 2028 1737
rect 2019 1716 2023 1717
rect 1942 1714 1948 1715
rect 1942 1710 1943 1714
rect 1947 1710 1948 1714
rect 2019 1711 2023 1712
rect 2038 1714 2044 1715
rect 1942 1709 1948 1710
rect 1918 1707 1924 1708
rect 1918 1703 1919 1707
rect 1923 1703 1924 1707
rect 1918 1702 1924 1703
rect 1944 1691 1946 1709
rect 2020 1708 2022 1711
rect 2038 1710 2039 1714
rect 2043 1710 2044 1714
rect 2038 1709 2044 1710
rect 2018 1707 2024 1708
rect 2018 1703 2019 1707
rect 2023 1703 2024 1707
rect 2018 1702 2024 1703
rect 2040 1691 2042 1709
rect 2112 1708 2114 1738
rect 2118 1737 2119 1741
rect 2123 1737 2124 1741
rect 2154 1739 2155 1743
rect 2159 1739 2160 1743
rect 2208 1742 2210 1753
rect 2278 1743 2284 1744
rect 2154 1738 2160 1739
rect 2206 1741 2212 1742
rect 2118 1736 2124 1737
rect 2206 1737 2207 1741
rect 2211 1737 2212 1741
rect 2278 1739 2279 1743
rect 2283 1739 2284 1743
rect 2288 1742 2290 1753
rect 2366 1743 2372 1744
rect 2278 1738 2284 1739
rect 2286 1741 2292 1742
rect 2206 1736 2212 1737
rect 2134 1714 2140 1715
rect 2134 1710 2135 1714
rect 2139 1710 2140 1714
rect 2134 1709 2140 1710
rect 2222 1714 2228 1715
rect 2222 1710 2223 1714
rect 2227 1710 2228 1714
rect 2222 1709 2228 1710
rect 2110 1707 2116 1708
rect 2110 1703 2111 1707
rect 2115 1703 2116 1707
rect 2110 1702 2116 1703
rect 2136 1691 2138 1709
rect 2224 1691 2226 1709
rect 2280 1708 2282 1738
rect 2286 1737 2287 1741
rect 2291 1737 2292 1741
rect 2366 1739 2367 1743
rect 2371 1739 2372 1743
rect 2376 1742 2378 1753
rect 2398 1743 2404 1744
rect 2366 1738 2372 1739
rect 2374 1741 2380 1742
rect 2286 1736 2292 1737
rect 2302 1714 2308 1715
rect 2302 1710 2303 1714
rect 2307 1710 2308 1714
rect 2302 1709 2308 1710
rect 2230 1707 2236 1708
rect 2230 1703 2231 1707
rect 2235 1703 2236 1707
rect 2230 1702 2236 1703
rect 2278 1707 2284 1708
rect 2278 1703 2279 1707
rect 2283 1703 2284 1707
rect 2278 1702 2284 1703
rect 1799 1690 1803 1691
rect 1799 1685 1803 1686
rect 1839 1690 1843 1691
rect 1839 1685 1843 1686
rect 1887 1690 1891 1691
rect 1887 1685 1891 1686
rect 1943 1690 1947 1691
rect 1943 1685 1947 1686
rect 1975 1690 1979 1691
rect 1975 1685 1979 1686
rect 2039 1690 2043 1691
rect 2039 1685 2043 1686
rect 2063 1690 2067 1691
rect 2063 1685 2067 1686
rect 2135 1690 2139 1691
rect 2135 1685 2139 1686
rect 2143 1690 2147 1691
rect 2143 1685 2147 1686
rect 2215 1690 2219 1691
rect 2215 1685 2219 1686
rect 2223 1690 2227 1691
rect 2223 1685 2227 1686
rect 1774 1683 1780 1684
rect 1774 1679 1775 1683
rect 1779 1679 1780 1683
rect 1800 1679 1802 1685
rect 1818 1683 1824 1684
rect 1818 1679 1819 1683
rect 1823 1679 1824 1683
rect 1888 1679 1890 1685
rect 1902 1683 1908 1684
rect 1902 1679 1903 1683
rect 1907 1679 1908 1683
rect 1976 1679 1978 1685
rect 2064 1679 2066 1685
rect 2082 1683 2088 1684
rect 2082 1679 2083 1683
rect 2087 1679 2088 1683
rect 2144 1679 2146 1685
rect 2162 1683 2168 1684
rect 2162 1679 2163 1683
rect 2167 1679 2168 1683
rect 2216 1679 2218 1685
rect 1774 1678 1780 1679
rect 1798 1678 1804 1679
rect 1818 1678 1824 1679
rect 1886 1678 1892 1679
rect 1902 1678 1908 1679
rect 1974 1678 1980 1679
rect 1798 1674 1799 1678
rect 1803 1674 1804 1678
rect 1798 1673 1804 1674
rect 1782 1651 1788 1652
rect 1694 1646 1700 1647
rect 1722 1647 1728 1648
rect 1650 1642 1656 1643
rect 1696 1623 1698 1646
rect 1722 1643 1723 1647
rect 1727 1643 1728 1647
rect 1782 1647 1783 1651
rect 1787 1647 1788 1651
rect 1820 1648 1822 1678
rect 1886 1674 1887 1678
rect 1891 1674 1892 1678
rect 1886 1673 1892 1674
rect 1870 1651 1876 1652
rect 1782 1646 1788 1647
rect 1818 1647 1824 1648
rect 1722 1642 1728 1643
rect 1784 1623 1786 1646
rect 1818 1643 1819 1647
rect 1823 1643 1824 1647
rect 1870 1647 1871 1651
rect 1875 1647 1876 1651
rect 1904 1648 1906 1678
rect 1974 1674 1975 1678
rect 1979 1674 1980 1678
rect 1974 1673 1980 1674
rect 2062 1678 2068 1679
rect 2082 1678 2088 1679
rect 2142 1678 2148 1679
rect 2162 1678 2168 1679
rect 2214 1678 2220 1679
rect 2062 1674 2063 1678
rect 2067 1674 2068 1678
rect 2062 1673 2068 1674
rect 1958 1651 1964 1652
rect 1870 1646 1876 1647
rect 1902 1647 1908 1648
rect 1818 1642 1824 1643
rect 1872 1623 1874 1646
rect 1902 1643 1903 1647
rect 1907 1643 1908 1647
rect 1958 1647 1959 1651
rect 1963 1647 1964 1651
rect 2046 1651 2052 1652
rect 1958 1646 1964 1647
rect 1982 1647 1988 1648
rect 1902 1642 1908 1643
rect 1960 1623 1962 1646
rect 1982 1643 1983 1647
rect 1987 1643 1988 1647
rect 2046 1647 2047 1651
rect 2051 1647 2052 1651
rect 2084 1648 2086 1678
rect 2142 1674 2143 1678
rect 2147 1674 2148 1678
rect 2142 1673 2148 1674
rect 2126 1651 2132 1652
rect 2046 1646 2052 1647
rect 2082 1647 2088 1648
rect 1982 1642 1988 1643
rect 1575 1622 1579 1623
rect 1575 1617 1579 1618
rect 1615 1622 1619 1623
rect 1615 1617 1619 1618
rect 1631 1622 1635 1623
rect 1631 1617 1635 1618
rect 1687 1622 1691 1623
rect 1687 1617 1691 1618
rect 1695 1622 1699 1623
rect 1695 1617 1699 1618
rect 1751 1622 1755 1623
rect 1751 1617 1755 1618
rect 1783 1622 1787 1623
rect 1783 1617 1787 1618
rect 1831 1622 1835 1623
rect 1831 1617 1835 1618
rect 1871 1622 1875 1623
rect 1871 1617 1875 1618
rect 1919 1622 1923 1623
rect 1919 1617 1923 1618
rect 1959 1622 1963 1623
rect 1959 1617 1963 1618
rect 1550 1611 1556 1612
rect 1550 1607 1551 1611
rect 1555 1607 1556 1611
rect 1550 1606 1556 1607
rect 1576 1606 1578 1617
rect 1632 1606 1634 1617
rect 1688 1606 1690 1617
rect 1752 1606 1754 1617
rect 1832 1606 1834 1617
rect 1920 1606 1922 1617
rect 1574 1605 1580 1606
rect 1327 1601 1331 1602
rect 1366 1604 1372 1605
rect 1152 1590 1154 1601
rect 1150 1589 1156 1590
rect 1328 1589 1330 1601
rect 1366 1600 1367 1604
rect 1371 1600 1372 1604
rect 1574 1601 1575 1605
rect 1579 1601 1580 1605
rect 1574 1600 1580 1601
rect 1630 1605 1636 1606
rect 1630 1601 1631 1605
rect 1635 1601 1636 1605
rect 1630 1600 1636 1601
rect 1686 1605 1692 1606
rect 1686 1601 1687 1605
rect 1691 1601 1692 1605
rect 1686 1600 1692 1601
rect 1750 1605 1756 1606
rect 1750 1601 1751 1605
rect 1755 1601 1756 1605
rect 1750 1600 1756 1601
rect 1830 1605 1836 1606
rect 1830 1601 1831 1605
rect 1835 1601 1836 1605
rect 1830 1600 1836 1601
rect 1918 1605 1924 1606
rect 1918 1601 1919 1605
rect 1923 1601 1924 1605
rect 1918 1600 1924 1601
rect 1366 1599 1372 1600
rect 1150 1585 1151 1589
rect 1155 1585 1156 1589
rect 1150 1584 1156 1585
rect 1326 1588 1332 1589
rect 1326 1584 1327 1588
rect 1331 1584 1332 1588
rect 1326 1583 1332 1584
rect 1366 1587 1372 1588
rect 1366 1583 1367 1587
rect 1371 1583 1372 1587
rect 1366 1582 1372 1583
rect 1326 1571 1332 1572
rect 1326 1567 1327 1571
rect 1331 1567 1332 1571
rect 1326 1566 1332 1567
rect 1166 1562 1172 1563
rect 1166 1558 1167 1562
rect 1171 1558 1172 1562
rect 1166 1557 1172 1558
rect 1142 1555 1148 1556
rect 1142 1551 1143 1555
rect 1147 1551 1148 1555
rect 1168 1551 1170 1557
rect 1328 1551 1330 1566
rect 1368 1563 1370 1582
rect 1590 1578 1596 1579
rect 1590 1574 1591 1578
rect 1595 1574 1596 1578
rect 1590 1573 1596 1574
rect 1646 1578 1652 1579
rect 1646 1574 1647 1578
rect 1651 1574 1652 1578
rect 1646 1573 1652 1574
rect 1702 1578 1708 1579
rect 1702 1574 1703 1578
rect 1707 1574 1708 1578
rect 1702 1573 1708 1574
rect 1766 1578 1772 1579
rect 1766 1574 1767 1578
rect 1771 1574 1772 1578
rect 1766 1573 1772 1574
rect 1846 1578 1852 1579
rect 1846 1574 1847 1578
rect 1851 1574 1852 1578
rect 1846 1573 1852 1574
rect 1934 1578 1940 1579
rect 1934 1574 1935 1578
rect 1939 1574 1940 1578
rect 1934 1573 1940 1574
rect 1592 1563 1594 1573
rect 1648 1563 1650 1573
rect 1704 1563 1706 1573
rect 1768 1563 1770 1573
rect 1848 1563 1850 1573
rect 1902 1571 1908 1572
rect 1902 1567 1903 1571
rect 1907 1567 1908 1571
rect 1902 1566 1908 1567
rect 1367 1562 1371 1563
rect 1367 1557 1371 1558
rect 1591 1562 1595 1563
rect 1591 1557 1595 1558
rect 1647 1562 1651 1563
rect 1647 1557 1651 1558
rect 1679 1562 1683 1563
rect 1679 1557 1683 1558
rect 1703 1562 1707 1563
rect 1703 1557 1707 1558
rect 1735 1562 1739 1563
rect 1735 1557 1739 1558
rect 1767 1562 1771 1563
rect 1767 1557 1771 1558
rect 1791 1562 1795 1563
rect 1791 1557 1795 1558
rect 1847 1562 1851 1563
rect 1847 1557 1851 1558
rect 1855 1562 1859 1563
rect 1855 1557 1859 1558
rect 1055 1550 1059 1551
rect 1055 1545 1059 1546
rect 1079 1550 1083 1551
rect 1142 1550 1148 1551
rect 1167 1550 1171 1551
rect 1079 1545 1083 1546
rect 1167 1545 1171 1546
rect 1327 1550 1331 1551
rect 1327 1545 1331 1546
rect 1030 1543 1036 1544
rect 1030 1539 1031 1543
rect 1035 1539 1036 1543
rect 1056 1539 1058 1545
rect 734 1538 740 1539
rect 758 1538 764 1539
rect 806 1538 812 1539
rect 830 1538 836 1539
rect 878 1538 884 1539
rect 902 1538 908 1539
rect 966 1538 972 1539
rect 974 1538 980 1539
rect 1030 1538 1036 1539
rect 1054 1538 1060 1539
rect 736 1520 738 1538
rect 758 1534 759 1538
rect 763 1534 764 1538
rect 758 1533 764 1534
rect 734 1519 740 1520
rect 734 1515 735 1519
rect 739 1515 740 1519
rect 734 1514 740 1515
rect 742 1511 748 1512
rect 706 1507 712 1508
rect 706 1503 707 1507
rect 711 1503 712 1507
rect 742 1507 743 1511
rect 747 1507 748 1511
rect 742 1506 748 1507
rect 706 1502 712 1503
rect 678 1499 684 1500
rect 678 1495 679 1499
rect 683 1495 684 1499
rect 678 1494 684 1495
rect 744 1491 746 1506
rect 583 1490 587 1491
rect 583 1485 587 1486
rect 599 1490 603 1491
rect 599 1485 603 1486
rect 671 1490 675 1491
rect 671 1485 675 1486
rect 679 1490 683 1491
rect 679 1485 683 1486
rect 743 1490 747 1491
rect 743 1485 747 1486
rect 775 1490 779 1491
rect 775 1485 779 1486
rect 584 1474 586 1485
rect 680 1474 682 1485
rect 766 1475 772 1476
rect 582 1473 588 1474
rect 582 1469 583 1473
rect 587 1469 588 1473
rect 582 1468 588 1469
rect 678 1473 684 1474
rect 678 1469 679 1473
rect 683 1469 684 1473
rect 766 1471 767 1475
rect 771 1471 772 1475
rect 776 1474 778 1485
rect 808 1476 810 1538
rect 830 1534 831 1538
rect 835 1534 836 1538
rect 830 1533 836 1534
rect 880 1520 882 1538
rect 902 1534 903 1538
rect 907 1534 908 1538
rect 902 1533 908 1534
rect 878 1519 884 1520
rect 878 1515 879 1519
rect 883 1515 884 1519
rect 878 1514 884 1515
rect 814 1511 820 1512
rect 814 1507 815 1511
rect 819 1507 820 1511
rect 814 1506 820 1507
rect 886 1511 892 1512
rect 886 1507 887 1511
rect 891 1507 892 1511
rect 958 1511 964 1512
rect 886 1506 892 1507
rect 910 1507 916 1508
rect 816 1491 818 1506
rect 888 1491 890 1506
rect 910 1503 911 1507
rect 915 1503 916 1507
rect 958 1507 959 1511
rect 963 1507 964 1511
rect 958 1506 964 1507
rect 910 1502 916 1503
rect 815 1490 819 1491
rect 815 1485 819 1486
rect 863 1490 867 1491
rect 863 1485 867 1486
rect 887 1490 891 1491
rect 887 1485 891 1486
rect 806 1475 812 1476
rect 766 1470 772 1471
rect 774 1473 780 1474
rect 678 1468 684 1469
rect 598 1446 604 1447
rect 598 1442 599 1446
rect 603 1442 604 1446
rect 598 1441 604 1442
rect 694 1446 700 1447
rect 694 1442 695 1446
rect 699 1442 700 1446
rect 694 1441 700 1442
rect 574 1439 580 1440
rect 574 1435 575 1439
rect 579 1435 580 1439
rect 574 1434 580 1435
rect 510 1431 516 1432
rect 600 1431 602 1441
rect 696 1431 698 1441
rect 768 1440 770 1470
rect 774 1469 775 1473
rect 779 1469 780 1473
rect 806 1471 807 1475
rect 811 1471 812 1475
rect 864 1474 866 1485
rect 806 1470 812 1471
rect 862 1473 868 1474
rect 774 1468 780 1469
rect 862 1469 863 1473
rect 867 1469 868 1473
rect 862 1468 868 1469
rect 790 1446 796 1447
rect 790 1442 791 1446
rect 795 1442 796 1446
rect 790 1441 796 1442
rect 878 1446 884 1447
rect 878 1442 879 1446
rect 883 1442 884 1446
rect 878 1441 884 1442
rect 758 1439 764 1440
rect 758 1435 759 1439
rect 763 1435 764 1439
rect 758 1434 764 1435
rect 766 1439 772 1440
rect 766 1435 767 1439
rect 771 1435 772 1439
rect 766 1434 772 1435
rect 215 1430 219 1431
rect 215 1425 219 1426
rect 247 1430 251 1431
rect 247 1425 251 1426
rect 303 1430 307 1431
rect 303 1425 307 1426
rect 343 1430 347 1431
rect 358 1427 359 1431
rect 363 1427 364 1431
rect 358 1426 364 1427
rect 399 1430 403 1431
rect 343 1425 347 1426
rect 248 1419 250 1425
rect 334 1423 340 1424
rect 334 1419 335 1423
rect 339 1419 340 1423
rect 344 1419 346 1425
rect 246 1418 252 1419
rect 334 1418 340 1419
rect 342 1418 348 1419
rect 246 1414 247 1418
rect 251 1414 252 1418
rect 246 1413 252 1414
rect 230 1391 236 1392
rect 112 1375 114 1387
rect 142 1386 148 1387
rect 174 1387 180 1388
rect 144 1375 146 1386
rect 174 1383 175 1387
rect 179 1383 180 1387
rect 230 1387 231 1391
rect 235 1387 236 1391
rect 230 1386 236 1387
rect 326 1391 332 1392
rect 326 1387 327 1391
rect 331 1387 332 1391
rect 326 1386 332 1387
rect 174 1382 180 1383
rect 232 1375 234 1386
rect 328 1375 330 1386
rect 111 1374 115 1375
rect 111 1369 115 1370
rect 143 1374 147 1375
rect 143 1369 147 1370
rect 207 1374 211 1375
rect 207 1369 211 1370
rect 231 1374 235 1375
rect 231 1369 235 1370
rect 295 1374 299 1375
rect 295 1369 299 1370
rect 327 1374 331 1375
rect 327 1369 331 1370
rect 112 1357 114 1369
rect 144 1358 146 1369
rect 198 1359 204 1360
rect 142 1357 148 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 142 1353 143 1357
rect 147 1353 148 1357
rect 198 1355 199 1359
rect 203 1355 204 1359
rect 208 1358 210 1369
rect 286 1359 292 1360
rect 198 1354 204 1355
rect 206 1357 212 1358
rect 142 1352 148 1353
rect 110 1351 116 1352
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 110 1334 116 1335
rect 112 1319 114 1334
rect 158 1330 164 1331
rect 158 1326 159 1330
rect 163 1326 164 1330
rect 158 1325 164 1326
rect 160 1319 162 1325
rect 200 1324 202 1354
rect 206 1353 207 1357
rect 211 1353 212 1357
rect 286 1355 287 1359
rect 291 1355 292 1359
rect 296 1358 298 1369
rect 336 1368 338 1418
rect 342 1414 343 1418
rect 347 1414 348 1418
rect 342 1413 348 1414
rect 360 1388 362 1426
rect 399 1425 403 1426
rect 447 1430 451 1431
rect 447 1425 451 1426
rect 503 1430 507 1431
rect 510 1427 511 1431
rect 515 1427 516 1431
rect 510 1426 516 1427
rect 551 1430 555 1431
rect 503 1425 507 1426
rect 551 1425 555 1426
rect 599 1430 603 1431
rect 599 1425 603 1426
rect 663 1430 667 1431
rect 663 1425 667 1426
rect 695 1430 699 1431
rect 695 1425 699 1426
rect 448 1419 450 1425
rect 466 1423 472 1424
rect 466 1419 467 1423
rect 471 1419 472 1423
rect 552 1419 554 1425
rect 570 1423 576 1424
rect 570 1419 571 1423
rect 575 1419 576 1423
rect 664 1419 666 1425
rect 742 1423 748 1424
rect 742 1419 743 1423
rect 747 1419 748 1423
rect 446 1418 452 1419
rect 466 1418 472 1419
rect 550 1418 556 1419
rect 570 1418 576 1419
rect 662 1418 668 1419
rect 742 1418 748 1419
rect 446 1414 447 1418
rect 451 1414 452 1418
rect 446 1413 452 1414
rect 430 1391 436 1392
rect 358 1387 364 1388
rect 358 1383 359 1387
rect 363 1383 364 1387
rect 430 1387 431 1391
rect 435 1387 436 1391
rect 468 1388 470 1418
rect 550 1414 551 1418
rect 555 1414 556 1418
rect 550 1413 556 1414
rect 534 1391 540 1392
rect 430 1386 436 1387
rect 466 1387 472 1388
rect 358 1382 364 1383
rect 432 1375 434 1386
rect 466 1383 467 1387
rect 471 1383 472 1387
rect 534 1387 535 1391
rect 539 1387 540 1391
rect 572 1388 574 1418
rect 662 1414 663 1418
rect 667 1414 668 1418
rect 662 1413 668 1414
rect 744 1400 746 1418
rect 742 1399 748 1400
rect 742 1395 743 1399
rect 747 1395 748 1399
rect 742 1394 748 1395
rect 646 1391 652 1392
rect 534 1386 540 1387
rect 570 1387 576 1388
rect 466 1382 472 1383
rect 536 1375 538 1386
rect 570 1383 571 1387
rect 575 1383 576 1387
rect 646 1387 647 1391
rect 651 1387 652 1391
rect 750 1391 756 1392
rect 646 1386 652 1387
rect 670 1387 676 1388
rect 570 1382 576 1383
rect 648 1375 650 1386
rect 670 1383 671 1387
rect 675 1383 676 1387
rect 750 1387 751 1391
rect 755 1387 756 1391
rect 750 1386 756 1387
rect 670 1382 676 1383
rect 399 1374 403 1375
rect 399 1369 403 1370
rect 431 1374 435 1375
rect 431 1369 435 1370
rect 511 1374 515 1375
rect 511 1369 515 1370
rect 535 1374 539 1375
rect 535 1369 539 1370
rect 623 1374 627 1375
rect 623 1369 627 1370
rect 647 1374 651 1375
rect 647 1369 651 1370
rect 334 1367 340 1368
rect 334 1363 335 1367
rect 339 1363 340 1367
rect 334 1362 340 1363
rect 390 1359 396 1360
rect 286 1354 292 1355
rect 294 1357 300 1358
rect 206 1352 212 1353
rect 222 1330 228 1331
rect 222 1326 223 1330
rect 227 1326 228 1330
rect 222 1325 228 1326
rect 174 1323 180 1324
rect 174 1319 175 1323
rect 179 1319 180 1323
rect 111 1318 115 1319
rect 111 1313 115 1314
rect 159 1318 163 1319
rect 174 1318 180 1319
rect 198 1323 204 1324
rect 198 1319 199 1323
rect 203 1319 204 1323
rect 224 1319 226 1325
rect 288 1324 290 1354
rect 294 1353 295 1357
rect 299 1353 300 1357
rect 390 1355 391 1359
rect 395 1355 396 1359
rect 400 1358 402 1369
rect 474 1363 480 1364
rect 474 1359 475 1363
rect 479 1359 480 1363
rect 474 1358 480 1359
rect 512 1358 514 1369
rect 624 1358 626 1369
rect 390 1354 396 1355
rect 398 1357 404 1358
rect 294 1352 300 1353
rect 310 1330 316 1331
rect 310 1326 311 1330
rect 315 1326 316 1330
rect 310 1325 316 1326
rect 286 1323 292 1324
rect 286 1319 287 1323
rect 291 1319 292 1323
rect 312 1319 314 1325
rect 392 1324 394 1354
rect 398 1353 399 1357
rect 403 1353 404 1357
rect 398 1352 404 1353
rect 414 1330 420 1331
rect 414 1326 415 1330
rect 419 1326 420 1330
rect 414 1325 420 1326
rect 390 1323 396 1324
rect 342 1319 348 1320
rect 198 1318 204 1319
rect 223 1318 227 1319
rect 159 1313 163 1314
rect 112 1298 114 1313
rect 134 1311 140 1312
rect 134 1307 135 1311
rect 139 1307 140 1311
rect 160 1307 162 1313
rect 134 1306 140 1307
rect 158 1306 164 1307
rect 110 1297 116 1298
rect 110 1293 111 1297
rect 115 1293 116 1297
rect 110 1292 116 1293
rect 136 1288 138 1306
rect 158 1302 159 1306
rect 163 1302 164 1306
rect 158 1301 164 1302
rect 134 1287 140 1288
rect 134 1283 135 1287
rect 139 1283 140 1287
rect 134 1282 140 1283
rect 110 1280 116 1281
rect 110 1276 111 1280
rect 115 1276 116 1280
rect 110 1275 116 1276
rect 142 1279 148 1280
rect 142 1275 143 1279
rect 147 1275 148 1279
rect 176 1276 178 1318
rect 223 1313 227 1314
rect 231 1318 235 1319
rect 286 1318 292 1319
rect 311 1318 315 1319
rect 231 1313 235 1314
rect 311 1313 315 1314
rect 327 1318 331 1319
rect 342 1315 343 1319
rect 347 1315 348 1319
rect 390 1319 391 1323
rect 395 1319 396 1323
rect 416 1319 418 1325
rect 390 1318 396 1319
rect 415 1318 419 1319
rect 342 1314 348 1315
rect 327 1313 331 1314
rect 232 1307 234 1313
rect 302 1311 308 1312
rect 302 1307 303 1311
rect 307 1307 308 1311
rect 328 1307 330 1313
rect 230 1306 236 1307
rect 302 1306 308 1307
rect 326 1306 332 1307
rect 230 1302 231 1306
rect 235 1302 236 1306
rect 230 1301 236 1302
rect 214 1279 220 1280
rect 112 1251 114 1275
rect 142 1274 148 1275
rect 174 1275 180 1276
rect 144 1251 146 1274
rect 174 1271 175 1275
rect 179 1271 180 1275
rect 214 1275 215 1279
rect 219 1275 220 1279
rect 214 1274 220 1275
rect 174 1270 180 1271
rect 216 1251 218 1274
rect 111 1250 115 1251
rect 111 1245 115 1246
rect 143 1250 147 1251
rect 143 1245 147 1246
rect 199 1250 203 1251
rect 199 1245 203 1246
rect 215 1250 219 1251
rect 215 1245 219 1246
rect 279 1250 283 1251
rect 279 1245 283 1246
rect 112 1233 114 1245
rect 144 1234 146 1245
rect 150 1243 156 1244
rect 150 1239 151 1243
rect 155 1239 156 1243
rect 150 1238 156 1239
rect 142 1233 148 1234
rect 110 1232 116 1233
rect 110 1228 111 1232
rect 115 1228 116 1232
rect 142 1229 143 1233
rect 147 1229 148 1233
rect 142 1228 148 1229
rect 110 1227 116 1228
rect 110 1215 116 1216
rect 110 1211 111 1215
rect 115 1211 116 1215
rect 110 1210 116 1211
rect 112 1191 114 1210
rect 152 1200 154 1238
rect 190 1235 196 1236
rect 190 1231 191 1235
rect 195 1231 196 1235
rect 200 1234 202 1245
rect 270 1235 276 1236
rect 190 1230 196 1231
rect 198 1233 204 1234
rect 158 1206 164 1207
rect 158 1202 159 1206
rect 163 1202 164 1206
rect 158 1201 164 1202
rect 150 1199 156 1200
rect 150 1195 151 1199
rect 155 1195 156 1199
rect 150 1194 156 1195
rect 160 1191 162 1201
rect 192 1200 194 1230
rect 198 1229 199 1233
rect 203 1229 204 1233
rect 270 1231 271 1235
rect 275 1231 276 1235
rect 280 1234 282 1245
rect 304 1236 306 1306
rect 326 1302 327 1306
rect 331 1302 332 1306
rect 326 1301 332 1302
rect 310 1279 316 1280
rect 310 1275 311 1279
rect 315 1275 316 1279
rect 344 1276 346 1314
rect 415 1313 419 1314
rect 431 1318 435 1319
rect 476 1316 478 1358
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 622 1357 628 1358
rect 622 1353 623 1357
rect 627 1353 628 1357
rect 622 1352 628 1353
rect 526 1330 532 1331
rect 526 1326 527 1330
rect 531 1326 532 1330
rect 526 1325 532 1326
rect 638 1330 644 1331
rect 638 1326 639 1330
rect 643 1326 644 1330
rect 638 1325 644 1326
rect 528 1319 530 1325
rect 640 1319 642 1325
rect 672 1324 674 1382
rect 752 1375 754 1386
rect 760 1384 762 1434
rect 792 1431 794 1441
rect 880 1431 882 1441
rect 912 1440 914 1502
rect 960 1491 962 1506
rect 968 1500 970 1538
rect 974 1534 975 1538
rect 979 1534 980 1538
rect 974 1533 980 1534
rect 1054 1534 1055 1538
rect 1059 1534 1060 1538
rect 1054 1533 1060 1534
rect 1328 1530 1330 1545
rect 1368 1542 1370 1557
rect 1670 1555 1676 1556
rect 1670 1551 1671 1555
rect 1675 1551 1676 1555
rect 1680 1551 1682 1557
rect 1736 1551 1738 1557
rect 1754 1555 1760 1556
rect 1754 1551 1755 1555
rect 1759 1551 1760 1555
rect 1792 1551 1794 1557
rect 1810 1555 1816 1556
rect 1810 1551 1811 1555
rect 1815 1551 1816 1555
rect 1856 1551 1858 1557
rect 1874 1555 1880 1556
rect 1874 1551 1875 1555
rect 1879 1551 1880 1555
rect 1670 1550 1676 1551
rect 1678 1550 1684 1551
rect 1366 1541 1372 1542
rect 1366 1537 1367 1541
rect 1371 1537 1372 1541
rect 1366 1536 1372 1537
rect 1326 1529 1332 1530
rect 1326 1525 1327 1529
rect 1331 1525 1332 1529
rect 1326 1524 1332 1525
rect 1366 1524 1372 1525
rect 1366 1520 1367 1524
rect 1371 1520 1372 1524
rect 1366 1519 1372 1520
rect 1662 1523 1668 1524
rect 1662 1519 1663 1523
rect 1667 1519 1668 1523
rect 1326 1512 1332 1513
rect 1038 1511 1044 1512
rect 1038 1507 1039 1511
rect 1043 1507 1044 1511
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1326 1507 1332 1508
rect 1038 1506 1044 1507
rect 966 1499 972 1500
rect 966 1495 967 1499
rect 971 1495 972 1499
rect 966 1494 972 1495
rect 1040 1491 1042 1506
rect 1328 1491 1330 1507
rect 1368 1499 1370 1519
rect 1662 1518 1668 1519
rect 1664 1499 1666 1518
rect 1367 1498 1371 1499
rect 1367 1493 1371 1494
rect 1519 1498 1523 1499
rect 1519 1493 1523 1494
rect 1575 1498 1579 1499
rect 1575 1493 1579 1494
rect 1647 1498 1651 1499
rect 1647 1493 1651 1494
rect 1663 1498 1667 1499
rect 1663 1493 1667 1494
rect 951 1490 955 1491
rect 951 1485 955 1486
rect 959 1490 963 1491
rect 959 1485 963 1486
rect 1039 1490 1043 1491
rect 1039 1485 1043 1486
rect 1135 1490 1139 1491
rect 1135 1485 1139 1486
rect 1327 1490 1331 1491
rect 1327 1485 1331 1486
rect 942 1475 948 1476
rect 942 1471 943 1475
rect 947 1471 948 1475
rect 952 1474 954 1485
rect 1030 1475 1036 1476
rect 942 1470 948 1471
rect 950 1473 956 1474
rect 944 1440 946 1470
rect 950 1469 951 1473
rect 955 1469 956 1473
rect 1030 1471 1031 1475
rect 1035 1471 1036 1475
rect 1040 1474 1042 1485
rect 1126 1475 1132 1476
rect 1030 1470 1036 1471
rect 1038 1473 1044 1474
rect 950 1468 956 1469
rect 966 1446 972 1447
rect 966 1442 967 1446
rect 971 1442 972 1446
rect 966 1441 972 1442
rect 910 1439 916 1440
rect 910 1435 911 1439
rect 915 1435 916 1439
rect 910 1434 916 1435
rect 942 1439 948 1440
rect 942 1435 943 1439
rect 947 1435 948 1439
rect 942 1434 948 1435
rect 968 1431 970 1441
rect 1032 1440 1034 1470
rect 1038 1469 1039 1473
rect 1043 1469 1044 1473
rect 1126 1471 1127 1475
rect 1131 1471 1132 1475
rect 1136 1474 1138 1485
rect 1190 1475 1196 1476
rect 1126 1470 1132 1471
rect 1134 1473 1140 1474
rect 1038 1468 1044 1469
rect 1054 1446 1060 1447
rect 1054 1442 1055 1446
rect 1059 1442 1060 1446
rect 1054 1441 1060 1442
rect 1030 1439 1036 1440
rect 1030 1435 1031 1439
rect 1035 1435 1036 1439
rect 1030 1434 1036 1435
rect 1056 1431 1058 1441
rect 1128 1440 1130 1470
rect 1134 1469 1135 1473
rect 1139 1469 1140 1473
rect 1190 1471 1191 1475
rect 1195 1471 1196 1475
rect 1328 1473 1330 1485
rect 1368 1481 1370 1493
rect 1520 1482 1522 1493
rect 1566 1483 1572 1484
rect 1518 1481 1524 1482
rect 1366 1480 1372 1481
rect 1366 1476 1367 1480
rect 1371 1476 1372 1480
rect 1518 1477 1519 1481
rect 1523 1477 1524 1481
rect 1566 1479 1567 1483
rect 1571 1479 1572 1483
rect 1576 1482 1578 1493
rect 1638 1483 1644 1484
rect 1566 1478 1572 1479
rect 1574 1481 1580 1482
rect 1518 1476 1524 1477
rect 1366 1475 1372 1476
rect 1190 1470 1196 1471
rect 1326 1472 1332 1473
rect 1134 1468 1140 1469
rect 1150 1446 1156 1447
rect 1150 1442 1151 1446
rect 1155 1442 1156 1446
rect 1150 1441 1156 1442
rect 1126 1439 1132 1440
rect 1126 1435 1127 1439
rect 1131 1435 1132 1439
rect 1126 1434 1132 1435
rect 1118 1431 1124 1432
rect 1152 1431 1154 1441
rect 767 1430 771 1431
rect 767 1425 771 1426
rect 791 1430 795 1431
rect 791 1425 795 1426
rect 879 1430 883 1431
rect 879 1425 883 1426
rect 967 1430 971 1431
rect 967 1425 971 1426
rect 991 1430 995 1431
rect 991 1425 995 1426
rect 1055 1430 1059 1431
rect 1055 1425 1059 1426
rect 1103 1430 1107 1431
rect 1118 1427 1119 1431
rect 1123 1427 1124 1431
rect 1118 1426 1124 1427
rect 1151 1430 1155 1431
rect 1103 1425 1107 1426
rect 768 1419 770 1425
rect 870 1423 876 1424
rect 870 1419 871 1423
rect 875 1419 876 1423
rect 880 1419 882 1425
rect 992 1419 994 1425
rect 1078 1423 1084 1424
rect 1078 1419 1079 1423
rect 1083 1419 1084 1423
rect 1104 1419 1106 1425
rect 766 1418 772 1419
rect 870 1418 876 1419
rect 878 1418 884 1419
rect 766 1414 767 1418
rect 771 1414 772 1418
rect 766 1413 772 1414
rect 862 1391 868 1392
rect 862 1387 863 1391
rect 867 1387 868 1391
rect 862 1386 868 1387
rect 758 1383 764 1384
rect 758 1379 759 1383
rect 763 1379 764 1383
rect 758 1378 764 1379
rect 864 1375 866 1386
rect 735 1374 739 1375
rect 735 1369 739 1370
rect 751 1374 755 1375
rect 751 1369 755 1370
rect 847 1374 851 1375
rect 847 1369 851 1370
rect 863 1374 867 1375
rect 863 1369 867 1370
rect 736 1358 738 1369
rect 838 1359 844 1360
rect 734 1357 740 1358
rect 734 1353 735 1357
rect 739 1353 740 1357
rect 838 1355 839 1359
rect 843 1355 844 1359
rect 848 1358 850 1369
rect 872 1360 874 1418
rect 878 1414 879 1418
rect 883 1414 884 1418
rect 878 1413 884 1414
rect 990 1418 996 1419
rect 1078 1418 1084 1419
rect 1102 1418 1108 1419
rect 990 1414 991 1418
rect 995 1414 996 1418
rect 990 1413 996 1414
rect 1080 1400 1082 1418
rect 1102 1414 1103 1418
rect 1107 1414 1108 1418
rect 1102 1413 1108 1414
rect 1078 1399 1084 1400
rect 1078 1395 1079 1399
rect 1083 1395 1084 1399
rect 1078 1394 1084 1395
rect 974 1391 980 1392
rect 974 1387 975 1391
rect 979 1387 980 1391
rect 1086 1391 1092 1392
rect 974 1386 980 1387
rect 998 1387 1004 1388
rect 976 1375 978 1386
rect 998 1383 999 1387
rect 1003 1383 1004 1387
rect 1086 1387 1087 1391
rect 1091 1387 1092 1391
rect 1120 1388 1122 1426
rect 1151 1425 1155 1426
rect 1192 1424 1194 1470
rect 1326 1468 1327 1472
rect 1331 1468 1332 1472
rect 1326 1467 1332 1468
rect 1366 1463 1372 1464
rect 1366 1459 1367 1463
rect 1371 1459 1372 1463
rect 1366 1458 1372 1459
rect 1326 1455 1332 1456
rect 1326 1451 1327 1455
rect 1331 1451 1332 1455
rect 1326 1450 1332 1451
rect 1328 1431 1330 1450
rect 1368 1435 1370 1458
rect 1534 1454 1540 1455
rect 1534 1450 1535 1454
rect 1539 1450 1540 1454
rect 1534 1449 1540 1450
rect 1536 1435 1538 1449
rect 1568 1448 1570 1478
rect 1574 1477 1575 1481
rect 1579 1477 1580 1481
rect 1638 1479 1639 1483
rect 1643 1479 1644 1483
rect 1648 1482 1650 1493
rect 1672 1492 1674 1550
rect 1678 1546 1679 1550
rect 1683 1546 1684 1550
rect 1678 1545 1684 1546
rect 1734 1550 1740 1551
rect 1754 1550 1760 1551
rect 1790 1550 1796 1551
rect 1810 1550 1816 1551
rect 1854 1550 1860 1551
rect 1874 1550 1880 1551
rect 1734 1546 1735 1550
rect 1739 1546 1740 1550
rect 1734 1545 1740 1546
rect 1718 1523 1724 1524
rect 1718 1519 1719 1523
rect 1723 1519 1724 1523
rect 1756 1520 1758 1550
rect 1790 1546 1791 1550
rect 1795 1546 1796 1550
rect 1790 1545 1796 1546
rect 1774 1523 1780 1524
rect 1718 1518 1724 1519
rect 1754 1519 1760 1520
rect 1720 1499 1722 1518
rect 1754 1515 1755 1519
rect 1759 1515 1760 1519
rect 1774 1519 1775 1523
rect 1779 1519 1780 1523
rect 1812 1520 1814 1550
rect 1854 1546 1855 1550
rect 1859 1546 1860 1550
rect 1854 1545 1860 1546
rect 1838 1523 1844 1524
rect 1774 1518 1780 1519
rect 1810 1519 1816 1520
rect 1754 1514 1760 1515
rect 1776 1499 1778 1518
rect 1810 1515 1811 1519
rect 1815 1515 1816 1519
rect 1838 1519 1839 1523
rect 1843 1519 1844 1523
rect 1876 1520 1878 1550
rect 1904 1532 1906 1566
rect 1936 1563 1938 1573
rect 1984 1572 1986 1642
rect 2048 1623 2050 1646
rect 2082 1643 2083 1647
rect 2087 1643 2088 1647
rect 2126 1647 2127 1651
rect 2131 1647 2132 1651
rect 2164 1648 2166 1678
rect 2214 1674 2215 1678
rect 2219 1674 2220 1678
rect 2214 1673 2220 1674
rect 2198 1651 2204 1652
rect 2126 1646 2132 1647
rect 2162 1647 2168 1648
rect 2082 1642 2088 1643
rect 2128 1623 2130 1646
rect 2162 1643 2163 1647
rect 2167 1643 2168 1647
rect 2198 1647 2199 1651
rect 2203 1647 2204 1651
rect 2232 1648 2234 1702
rect 2294 1691 2300 1692
rect 2304 1691 2306 1709
rect 2368 1708 2370 1738
rect 2374 1737 2375 1741
rect 2379 1737 2380 1741
rect 2398 1739 2399 1743
rect 2403 1739 2404 1743
rect 2464 1742 2466 1753
rect 2398 1738 2404 1739
rect 2462 1741 2468 1742
rect 2374 1736 2380 1737
rect 2400 1717 2402 1738
rect 2462 1737 2463 1741
rect 2467 1737 2468 1741
rect 2462 1736 2468 1737
rect 2399 1716 2403 1717
rect 2390 1714 2396 1715
rect 2390 1710 2391 1714
rect 2395 1710 2396 1714
rect 2399 1711 2403 1712
rect 2390 1709 2396 1710
rect 2366 1707 2372 1708
rect 2366 1703 2367 1707
rect 2371 1703 2372 1707
rect 2366 1702 2372 1703
rect 2392 1691 2394 1709
rect 2472 1708 2474 1762
rect 2528 1759 2530 1770
rect 2527 1758 2531 1759
rect 2527 1753 2531 1754
rect 2494 1743 2500 1744
rect 2494 1739 2495 1743
rect 2499 1739 2500 1743
rect 2528 1742 2530 1753
rect 2536 1748 2538 1802
rect 2542 1798 2543 1802
rect 2547 1798 2548 1802
rect 2542 1797 2548 1798
rect 2584 1794 2586 1809
rect 2582 1793 2588 1794
rect 2582 1789 2583 1793
rect 2587 1789 2588 1793
rect 2582 1788 2588 1789
rect 2582 1776 2588 1777
rect 2582 1772 2583 1776
rect 2587 1772 2588 1776
rect 2582 1771 2588 1772
rect 2584 1759 2586 1771
rect 2583 1758 2587 1759
rect 2583 1753 2587 1754
rect 2534 1747 2540 1748
rect 2534 1743 2535 1747
rect 2539 1743 2540 1747
rect 2534 1742 2540 1743
rect 2494 1738 2500 1739
rect 2526 1741 2532 1742
rect 2584 1741 2586 1753
rect 2478 1714 2484 1715
rect 2478 1710 2479 1714
rect 2483 1710 2484 1714
rect 2478 1709 2484 1710
rect 2470 1707 2476 1708
rect 2470 1703 2471 1707
rect 2475 1703 2476 1707
rect 2470 1702 2476 1703
rect 2434 1691 2440 1692
rect 2480 1691 2482 1709
rect 2287 1690 2291 1691
rect 2294 1687 2295 1691
rect 2299 1687 2300 1691
rect 2294 1686 2300 1687
rect 2303 1690 2307 1691
rect 2287 1685 2291 1686
rect 2262 1683 2268 1684
rect 2262 1679 2263 1683
rect 2267 1679 2268 1683
rect 2288 1679 2290 1685
rect 2262 1678 2268 1679
rect 2286 1678 2292 1679
rect 2264 1660 2266 1678
rect 2286 1674 2287 1678
rect 2291 1674 2292 1678
rect 2286 1673 2292 1674
rect 2262 1659 2268 1660
rect 2262 1655 2263 1659
rect 2267 1655 2268 1659
rect 2262 1654 2268 1655
rect 2270 1651 2276 1652
rect 2198 1646 2204 1647
rect 2230 1647 2236 1648
rect 2162 1642 2168 1643
rect 2200 1623 2202 1646
rect 2230 1643 2231 1647
rect 2235 1643 2236 1647
rect 2270 1647 2271 1651
rect 2275 1647 2276 1651
rect 2296 1648 2298 1686
rect 2303 1685 2307 1686
rect 2351 1690 2355 1691
rect 2351 1685 2355 1686
rect 2391 1690 2395 1691
rect 2391 1685 2395 1686
rect 2423 1690 2427 1691
rect 2434 1687 2435 1691
rect 2439 1687 2440 1691
rect 2434 1686 2440 1687
rect 2479 1690 2483 1691
rect 2423 1685 2427 1686
rect 2352 1679 2354 1685
rect 2398 1683 2404 1684
rect 2398 1679 2399 1683
rect 2403 1679 2404 1683
rect 2424 1679 2426 1685
rect 2350 1678 2356 1679
rect 2398 1678 2404 1679
rect 2422 1678 2428 1679
rect 2350 1674 2351 1678
rect 2355 1674 2356 1678
rect 2350 1673 2356 1674
rect 2400 1660 2402 1678
rect 2422 1674 2423 1678
rect 2427 1674 2428 1678
rect 2422 1673 2428 1674
rect 2398 1659 2404 1660
rect 2398 1655 2399 1659
rect 2403 1655 2404 1659
rect 2398 1654 2404 1655
rect 2334 1651 2340 1652
rect 2270 1646 2276 1647
rect 2294 1647 2300 1648
rect 2230 1642 2236 1643
rect 2272 1623 2274 1646
rect 2294 1643 2295 1647
rect 2299 1643 2300 1647
rect 2334 1647 2335 1651
rect 2339 1647 2340 1651
rect 2334 1646 2340 1647
rect 2406 1651 2412 1652
rect 2406 1647 2407 1651
rect 2411 1647 2412 1651
rect 2436 1648 2438 1686
rect 2479 1685 2483 1686
rect 2487 1690 2491 1691
rect 2496 1688 2498 1738
rect 2526 1737 2527 1741
rect 2531 1737 2532 1741
rect 2526 1736 2532 1737
rect 2582 1740 2588 1741
rect 2582 1736 2583 1740
rect 2587 1736 2588 1740
rect 2582 1735 2588 1736
rect 2582 1723 2588 1724
rect 2582 1719 2583 1723
rect 2587 1719 2588 1723
rect 2582 1718 2588 1719
rect 2542 1714 2548 1715
rect 2542 1710 2543 1714
rect 2547 1710 2548 1714
rect 2542 1709 2548 1710
rect 2544 1691 2546 1709
rect 2558 1707 2564 1708
rect 2558 1703 2559 1707
rect 2563 1703 2564 1707
rect 2558 1702 2564 1703
rect 2543 1690 2547 1691
rect 2487 1685 2491 1686
rect 2494 1687 2500 1688
rect 2488 1679 2490 1685
rect 2494 1683 2495 1687
rect 2499 1683 2500 1687
rect 2543 1685 2547 1686
rect 2494 1682 2500 1683
rect 2534 1683 2540 1684
rect 2534 1679 2535 1683
rect 2539 1679 2540 1683
rect 2544 1679 2546 1685
rect 2486 1678 2492 1679
rect 2534 1678 2540 1679
rect 2542 1678 2548 1679
rect 2486 1674 2487 1678
rect 2491 1674 2492 1678
rect 2486 1673 2492 1674
rect 2470 1651 2476 1652
rect 2406 1646 2412 1647
rect 2434 1647 2440 1648
rect 2294 1642 2300 1643
rect 2336 1623 2338 1646
rect 2408 1623 2410 1646
rect 2434 1643 2435 1647
rect 2439 1643 2440 1647
rect 2470 1647 2471 1651
rect 2475 1647 2476 1651
rect 2470 1646 2476 1647
rect 2526 1651 2532 1652
rect 2526 1647 2527 1651
rect 2531 1647 2532 1651
rect 2526 1646 2532 1647
rect 2434 1642 2440 1643
rect 2472 1623 2474 1646
rect 2528 1623 2530 1646
rect 2007 1622 2011 1623
rect 2007 1617 2011 1618
rect 2047 1622 2051 1623
rect 2047 1617 2051 1618
rect 2103 1622 2107 1623
rect 2103 1617 2107 1618
rect 2127 1622 2131 1623
rect 2127 1617 2131 1618
rect 2199 1622 2203 1623
rect 2199 1617 2203 1618
rect 2207 1622 2211 1623
rect 2207 1617 2211 1618
rect 2271 1622 2275 1623
rect 2271 1617 2275 1618
rect 2319 1622 2323 1623
rect 2319 1617 2323 1618
rect 2335 1622 2339 1623
rect 2335 1617 2339 1618
rect 2407 1622 2411 1623
rect 2407 1617 2411 1618
rect 2431 1622 2435 1623
rect 2431 1617 2435 1618
rect 2471 1622 2475 1623
rect 2471 1617 2475 1618
rect 2527 1622 2531 1623
rect 2527 1617 2531 1618
rect 1998 1607 2004 1608
rect 1998 1603 1999 1607
rect 2003 1603 2004 1607
rect 2008 1606 2010 1617
rect 2094 1607 2100 1608
rect 1998 1602 2004 1603
rect 2006 1605 2012 1606
rect 2000 1572 2002 1602
rect 2006 1601 2007 1605
rect 2011 1601 2012 1605
rect 2094 1603 2095 1607
rect 2099 1603 2100 1607
rect 2104 1606 2106 1617
rect 2126 1607 2132 1608
rect 2094 1602 2100 1603
rect 2102 1605 2108 1606
rect 2006 1600 2012 1601
rect 2022 1578 2028 1579
rect 2022 1574 2023 1578
rect 2027 1574 2028 1578
rect 2022 1573 2028 1574
rect 1982 1571 1988 1572
rect 1982 1567 1983 1571
rect 1987 1567 1988 1571
rect 1982 1566 1988 1567
rect 1998 1571 2004 1572
rect 1998 1567 1999 1571
rect 2003 1567 2004 1571
rect 1998 1566 2004 1567
rect 2024 1563 2026 1573
rect 2096 1572 2098 1602
rect 2102 1601 2103 1605
rect 2107 1601 2108 1605
rect 2126 1603 2127 1607
rect 2131 1603 2132 1607
rect 2208 1606 2210 1617
rect 2310 1607 2316 1608
rect 2126 1602 2132 1603
rect 2206 1605 2212 1606
rect 2102 1600 2108 1601
rect 2118 1578 2124 1579
rect 2118 1574 2119 1578
rect 2123 1574 2124 1578
rect 2118 1573 2124 1574
rect 2094 1571 2100 1572
rect 2094 1567 2095 1571
rect 2099 1567 2100 1571
rect 2094 1566 2100 1567
rect 2120 1563 2122 1573
rect 1927 1562 1931 1563
rect 1927 1557 1931 1558
rect 1935 1562 1939 1563
rect 1935 1557 1939 1558
rect 2007 1562 2011 1563
rect 2007 1557 2011 1558
rect 2023 1562 2027 1563
rect 2023 1557 2027 1558
rect 2087 1562 2091 1563
rect 2087 1557 2091 1558
rect 2119 1562 2123 1563
rect 2128 1560 2130 1602
rect 2206 1601 2207 1605
rect 2211 1601 2212 1605
rect 2310 1603 2311 1607
rect 2315 1603 2316 1607
rect 2320 1606 2322 1617
rect 2422 1607 2428 1608
rect 2310 1602 2316 1603
rect 2318 1605 2324 1606
rect 2206 1600 2212 1601
rect 2222 1578 2228 1579
rect 2222 1574 2223 1578
rect 2227 1574 2228 1578
rect 2222 1573 2228 1574
rect 2224 1563 2226 1573
rect 2312 1572 2314 1602
rect 2318 1601 2319 1605
rect 2323 1601 2324 1605
rect 2422 1603 2423 1607
rect 2427 1603 2428 1607
rect 2432 1606 2434 1617
rect 2462 1607 2468 1608
rect 2422 1602 2428 1603
rect 2430 1605 2436 1606
rect 2318 1600 2324 1601
rect 2334 1578 2340 1579
rect 2334 1574 2335 1578
rect 2339 1574 2340 1578
rect 2334 1573 2340 1574
rect 2310 1571 2316 1572
rect 2310 1567 2311 1571
rect 2315 1567 2316 1571
rect 2310 1566 2316 1567
rect 2336 1563 2338 1573
rect 2424 1572 2426 1602
rect 2430 1601 2431 1605
rect 2435 1601 2436 1605
rect 2462 1603 2463 1607
rect 2467 1603 2468 1607
rect 2528 1606 2530 1617
rect 2536 1612 2538 1678
rect 2542 1674 2543 1678
rect 2547 1674 2548 1678
rect 2542 1673 2548 1674
rect 2560 1648 2562 1702
rect 2584 1691 2586 1718
rect 2583 1690 2587 1691
rect 2583 1685 2587 1686
rect 2584 1670 2586 1685
rect 2582 1669 2588 1670
rect 2582 1665 2583 1669
rect 2587 1665 2588 1669
rect 2582 1664 2588 1665
rect 2582 1652 2588 1653
rect 2582 1648 2583 1652
rect 2587 1648 2588 1652
rect 2558 1647 2564 1648
rect 2582 1647 2588 1648
rect 2558 1643 2559 1647
rect 2563 1643 2564 1647
rect 2558 1642 2564 1643
rect 2584 1623 2586 1647
rect 2583 1622 2587 1623
rect 2583 1617 2587 1618
rect 2534 1611 2540 1612
rect 2534 1607 2535 1611
rect 2539 1607 2540 1611
rect 2534 1606 2540 1607
rect 2462 1602 2468 1603
rect 2526 1605 2532 1606
rect 2584 1605 2586 1617
rect 2430 1600 2436 1601
rect 2446 1578 2452 1579
rect 2446 1574 2447 1578
rect 2451 1574 2452 1578
rect 2446 1573 2452 1574
rect 2422 1571 2428 1572
rect 2422 1567 2423 1571
rect 2427 1567 2428 1571
rect 2422 1566 2428 1567
rect 2342 1563 2348 1564
rect 2448 1563 2450 1573
rect 2167 1562 2171 1563
rect 2119 1557 2123 1558
rect 2126 1559 2132 1560
rect 1928 1551 1930 1557
rect 1946 1555 1952 1556
rect 1946 1551 1947 1555
rect 1951 1551 1952 1555
rect 2008 1551 2010 1557
rect 2088 1551 2090 1557
rect 2126 1555 2127 1559
rect 2131 1555 2132 1559
rect 2167 1557 2171 1558
rect 2223 1562 2227 1563
rect 2223 1557 2227 1558
rect 2247 1562 2251 1563
rect 2247 1557 2251 1558
rect 2327 1562 2331 1563
rect 2327 1557 2331 1558
rect 2335 1562 2339 1563
rect 2342 1559 2343 1563
rect 2347 1559 2348 1563
rect 2342 1558 2348 1559
rect 2407 1562 2411 1563
rect 2335 1557 2339 1558
rect 2126 1554 2132 1555
rect 2142 1555 2148 1556
rect 2142 1551 2143 1555
rect 2147 1551 2148 1555
rect 2168 1551 2170 1557
rect 2248 1551 2250 1557
rect 2266 1555 2272 1556
rect 2266 1551 2267 1555
rect 2271 1551 2272 1555
rect 2328 1551 2330 1557
rect 1926 1550 1932 1551
rect 1946 1550 1952 1551
rect 2006 1550 2012 1551
rect 1926 1546 1927 1550
rect 1931 1546 1932 1550
rect 1926 1545 1932 1546
rect 1902 1531 1908 1532
rect 1902 1527 1903 1531
rect 1907 1527 1908 1531
rect 1902 1526 1908 1527
rect 1910 1523 1916 1524
rect 1838 1518 1844 1519
rect 1874 1519 1880 1520
rect 1810 1514 1816 1515
rect 1840 1499 1842 1518
rect 1874 1515 1875 1519
rect 1879 1515 1880 1519
rect 1910 1519 1911 1523
rect 1915 1519 1916 1523
rect 1948 1520 1950 1550
rect 2006 1546 2007 1550
rect 2011 1546 2012 1550
rect 2006 1545 2012 1546
rect 2086 1550 2092 1551
rect 2142 1550 2148 1551
rect 2166 1550 2172 1551
rect 2086 1546 2087 1550
rect 2091 1546 2092 1550
rect 2086 1545 2092 1546
rect 2144 1532 2146 1550
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2246 1550 2252 1551
rect 2266 1550 2272 1551
rect 2326 1550 2332 1551
rect 2246 1546 2247 1550
rect 2251 1546 2252 1550
rect 2246 1545 2252 1546
rect 2142 1531 2148 1532
rect 2142 1527 2143 1531
rect 2147 1527 2148 1531
rect 2142 1526 2148 1527
rect 1990 1523 1996 1524
rect 1910 1518 1916 1519
rect 1946 1519 1952 1520
rect 1874 1514 1880 1515
rect 1912 1499 1914 1518
rect 1946 1515 1947 1519
rect 1951 1515 1952 1519
rect 1990 1519 1991 1523
rect 1995 1519 1996 1523
rect 1990 1518 1996 1519
rect 2070 1523 2076 1524
rect 2070 1519 2071 1523
rect 2075 1519 2076 1523
rect 2070 1518 2076 1519
rect 2150 1523 2156 1524
rect 2150 1519 2151 1523
rect 2155 1519 2156 1523
rect 2150 1518 2156 1519
rect 2230 1523 2236 1524
rect 2230 1519 2231 1523
rect 2235 1519 2236 1523
rect 2230 1518 2236 1519
rect 1946 1514 1952 1515
rect 1992 1499 1994 1518
rect 2034 1515 2040 1516
rect 2034 1511 2035 1515
rect 2039 1511 2040 1515
rect 2034 1510 2040 1511
rect 1719 1498 1723 1499
rect 1719 1493 1723 1494
rect 1727 1498 1731 1499
rect 1727 1493 1731 1494
rect 1775 1498 1779 1499
rect 1775 1493 1779 1494
rect 1807 1498 1811 1499
rect 1807 1493 1811 1494
rect 1839 1498 1843 1499
rect 1839 1493 1843 1494
rect 1895 1498 1899 1499
rect 1895 1493 1899 1494
rect 1911 1498 1915 1499
rect 1911 1493 1915 1494
rect 1983 1498 1987 1499
rect 1983 1493 1987 1494
rect 1991 1498 1995 1499
rect 1991 1493 1995 1494
rect 1670 1491 1676 1492
rect 1670 1487 1671 1491
rect 1675 1487 1676 1491
rect 1670 1486 1676 1487
rect 1718 1483 1724 1484
rect 1638 1478 1644 1479
rect 1646 1481 1652 1482
rect 1574 1476 1580 1477
rect 1590 1454 1596 1455
rect 1590 1450 1591 1454
rect 1595 1450 1596 1454
rect 1590 1449 1596 1450
rect 1566 1447 1572 1448
rect 1566 1443 1567 1447
rect 1571 1443 1572 1447
rect 1566 1442 1572 1443
rect 1592 1435 1594 1449
rect 1640 1448 1642 1478
rect 1646 1477 1647 1481
rect 1651 1477 1652 1481
rect 1718 1479 1719 1483
rect 1723 1479 1724 1483
rect 1728 1482 1730 1493
rect 1798 1483 1804 1484
rect 1718 1478 1724 1479
rect 1726 1481 1732 1482
rect 1646 1476 1652 1477
rect 1662 1454 1668 1455
rect 1662 1450 1663 1454
rect 1667 1450 1668 1454
rect 1662 1449 1668 1450
rect 1638 1447 1644 1448
rect 1638 1443 1639 1447
rect 1643 1443 1644 1447
rect 1638 1442 1644 1443
rect 1664 1435 1666 1449
rect 1720 1448 1722 1478
rect 1726 1477 1727 1481
rect 1731 1477 1732 1481
rect 1798 1479 1799 1483
rect 1803 1479 1804 1483
rect 1808 1482 1810 1493
rect 1886 1483 1892 1484
rect 1798 1478 1804 1479
rect 1806 1481 1812 1482
rect 1726 1476 1732 1477
rect 1742 1454 1748 1455
rect 1742 1450 1743 1454
rect 1747 1450 1748 1454
rect 1742 1449 1748 1450
rect 1718 1447 1724 1448
rect 1718 1443 1719 1447
rect 1723 1443 1724 1447
rect 1718 1442 1724 1443
rect 1744 1435 1746 1449
rect 1800 1448 1802 1478
rect 1806 1477 1807 1481
rect 1811 1477 1812 1481
rect 1886 1479 1887 1483
rect 1891 1479 1892 1483
rect 1896 1482 1898 1493
rect 1984 1482 1986 1493
rect 2006 1483 2012 1484
rect 1886 1478 1892 1479
rect 1894 1481 1900 1482
rect 1806 1476 1812 1477
rect 1822 1454 1828 1455
rect 1822 1450 1823 1454
rect 1827 1450 1828 1454
rect 1822 1449 1828 1450
rect 1798 1447 1804 1448
rect 1798 1443 1799 1447
rect 1803 1443 1804 1447
rect 1798 1442 1804 1443
rect 1824 1435 1826 1449
rect 1888 1448 1890 1478
rect 1894 1477 1895 1481
rect 1899 1477 1900 1481
rect 1894 1476 1900 1477
rect 1982 1481 1988 1482
rect 1982 1477 1983 1481
rect 1987 1477 1988 1481
rect 2006 1479 2007 1483
rect 2011 1479 2012 1483
rect 2006 1478 2012 1479
rect 1982 1476 1988 1477
rect 1910 1454 1916 1455
rect 1910 1450 1911 1454
rect 1915 1450 1916 1454
rect 1910 1449 1916 1450
rect 1998 1454 2004 1455
rect 1998 1450 1999 1454
rect 2003 1450 2004 1454
rect 1998 1449 2004 1450
rect 1886 1447 1892 1448
rect 1886 1443 1887 1447
rect 1891 1443 1892 1447
rect 1886 1442 1892 1443
rect 1838 1439 1844 1440
rect 1838 1435 1839 1439
rect 1843 1435 1844 1439
rect 1912 1435 1914 1449
rect 2000 1435 2002 1449
rect 2008 1436 2010 1478
rect 2036 1448 2038 1510
rect 2072 1499 2074 1518
rect 2152 1499 2154 1518
rect 2232 1499 2234 1518
rect 2071 1498 2075 1499
rect 2071 1493 2075 1494
rect 2151 1498 2155 1499
rect 2151 1493 2155 1494
rect 2231 1498 2235 1499
rect 2231 1493 2235 1494
rect 2072 1482 2074 1493
rect 2142 1483 2148 1484
rect 2070 1481 2076 1482
rect 2070 1477 2071 1481
rect 2075 1477 2076 1481
rect 2142 1479 2143 1483
rect 2147 1479 2148 1483
rect 2152 1482 2154 1493
rect 2222 1483 2228 1484
rect 2142 1478 2148 1479
rect 2150 1481 2156 1482
rect 2070 1476 2076 1477
rect 2086 1454 2092 1455
rect 2086 1450 2087 1454
rect 2091 1450 2092 1454
rect 2086 1449 2092 1450
rect 2034 1447 2040 1448
rect 2034 1443 2035 1447
rect 2039 1443 2040 1447
rect 2034 1442 2040 1443
rect 2042 1447 2048 1448
rect 2042 1443 2043 1447
rect 2047 1443 2048 1447
rect 2042 1442 2048 1443
rect 2006 1435 2012 1436
rect 1367 1434 1371 1435
rect 1215 1430 1219 1431
rect 1215 1425 1219 1426
rect 1327 1430 1331 1431
rect 1367 1429 1371 1430
rect 1415 1434 1419 1435
rect 1415 1429 1419 1430
rect 1471 1434 1475 1435
rect 1471 1429 1475 1430
rect 1535 1434 1539 1435
rect 1535 1429 1539 1430
rect 1591 1434 1595 1435
rect 1591 1429 1595 1430
rect 1623 1434 1627 1435
rect 1623 1429 1627 1430
rect 1663 1434 1667 1435
rect 1663 1429 1667 1430
rect 1719 1434 1723 1435
rect 1719 1429 1723 1430
rect 1743 1434 1747 1435
rect 1743 1429 1747 1430
rect 1823 1434 1827 1435
rect 1838 1434 1844 1435
rect 1911 1434 1915 1435
rect 1823 1429 1827 1430
rect 1327 1425 1331 1426
rect 1190 1423 1196 1424
rect 1190 1419 1191 1423
rect 1195 1419 1196 1423
rect 1216 1419 1218 1425
rect 1190 1418 1196 1419
rect 1214 1418 1220 1419
rect 1214 1414 1215 1418
rect 1219 1414 1220 1418
rect 1214 1413 1220 1414
rect 1328 1410 1330 1425
rect 1368 1414 1370 1429
rect 1406 1427 1412 1428
rect 1406 1423 1407 1427
rect 1411 1423 1412 1427
rect 1416 1423 1418 1429
rect 1434 1427 1440 1428
rect 1434 1423 1435 1427
rect 1439 1423 1440 1427
rect 1472 1423 1474 1429
rect 1502 1427 1508 1428
rect 1502 1423 1503 1427
rect 1507 1423 1508 1427
rect 1536 1423 1538 1429
rect 1554 1427 1560 1428
rect 1554 1423 1555 1427
rect 1559 1423 1560 1427
rect 1624 1423 1626 1429
rect 1642 1427 1648 1428
rect 1642 1423 1643 1427
rect 1647 1423 1648 1427
rect 1720 1423 1722 1429
rect 1824 1423 1826 1429
rect 1406 1422 1412 1423
rect 1414 1422 1420 1423
rect 1434 1422 1440 1423
rect 1470 1422 1476 1423
rect 1502 1422 1508 1423
rect 1534 1422 1540 1423
rect 1554 1422 1560 1423
rect 1622 1422 1628 1423
rect 1642 1422 1648 1423
rect 1718 1422 1724 1423
rect 1366 1413 1372 1414
rect 1326 1409 1332 1410
rect 1326 1405 1327 1409
rect 1331 1405 1332 1409
rect 1366 1409 1367 1413
rect 1371 1409 1372 1413
rect 1366 1408 1372 1409
rect 1326 1404 1332 1405
rect 1366 1396 1372 1397
rect 1326 1392 1332 1393
rect 1198 1391 1204 1392
rect 1086 1386 1092 1387
rect 1118 1387 1124 1388
rect 998 1382 1004 1383
rect 959 1374 963 1375
rect 959 1369 963 1370
rect 975 1374 979 1375
rect 975 1369 979 1370
rect 870 1359 876 1360
rect 838 1354 844 1355
rect 846 1357 852 1358
rect 734 1352 740 1353
rect 750 1330 756 1331
rect 750 1326 751 1330
rect 755 1326 756 1330
rect 750 1325 756 1326
rect 670 1323 676 1324
rect 670 1319 671 1323
rect 675 1319 676 1323
rect 742 1323 748 1324
rect 742 1319 743 1323
rect 747 1319 748 1323
rect 752 1319 754 1325
rect 840 1324 842 1354
rect 846 1353 847 1357
rect 851 1353 852 1357
rect 870 1355 871 1359
rect 875 1355 876 1359
rect 960 1358 962 1369
rect 870 1354 876 1355
rect 958 1357 964 1358
rect 846 1352 852 1353
rect 958 1353 959 1357
rect 963 1353 964 1357
rect 958 1352 964 1353
rect 891 1332 895 1333
rect 862 1330 868 1331
rect 862 1326 863 1330
rect 867 1326 868 1330
rect 891 1327 895 1328
rect 974 1330 980 1331
rect 862 1325 868 1326
rect 838 1323 844 1324
rect 838 1319 839 1323
rect 843 1319 844 1323
rect 864 1319 866 1325
rect 527 1318 531 1319
rect 431 1313 435 1314
rect 474 1315 480 1316
rect 432 1307 434 1313
rect 474 1311 475 1315
rect 479 1311 480 1315
rect 527 1313 531 1314
rect 535 1318 539 1319
rect 535 1313 539 1314
rect 631 1318 635 1319
rect 631 1313 635 1314
rect 639 1318 643 1319
rect 670 1318 676 1319
rect 727 1318 731 1319
rect 742 1318 748 1319
rect 751 1318 755 1319
rect 639 1313 643 1314
rect 727 1313 731 1314
rect 474 1310 480 1311
rect 482 1311 488 1312
rect 482 1307 483 1311
rect 487 1307 488 1311
rect 536 1307 538 1313
rect 606 1311 612 1312
rect 606 1307 607 1311
rect 611 1307 612 1311
rect 632 1307 634 1313
rect 650 1311 656 1312
rect 650 1307 651 1311
rect 655 1307 656 1311
rect 728 1307 730 1313
rect 430 1306 436 1307
rect 482 1306 488 1307
rect 534 1306 540 1307
rect 606 1306 612 1307
rect 630 1306 636 1307
rect 650 1306 656 1307
rect 726 1306 732 1307
rect 430 1302 431 1306
rect 435 1302 436 1306
rect 430 1301 436 1302
rect 414 1279 420 1280
rect 310 1274 316 1275
rect 342 1275 348 1276
rect 312 1251 314 1274
rect 342 1271 343 1275
rect 347 1271 348 1275
rect 414 1275 415 1279
rect 419 1275 420 1279
rect 484 1276 486 1306
rect 534 1302 535 1306
rect 539 1302 540 1306
rect 534 1301 540 1302
rect 608 1288 610 1306
rect 630 1302 631 1306
rect 635 1302 636 1306
rect 630 1301 636 1302
rect 606 1287 612 1288
rect 606 1283 607 1287
rect 611 1283 612 1287
rect 606 1282 612 1283
rect 518 1279 524 1280
rect 414 1274 420 1275
rect 482 1275 488 1276
rect 342 1270 348 1271
rect 416 1251 418 1274
rect 482 1271 483 1275
rect 487 1271 488 1275
rect 518 1275 519 1279
rect 523 1275 524 1279
rect 614 1279 620 1280
rect 518 1274 524 1275
rect 542 1275 548 1276
rect 482 1270 488 1271
rect 520 1251 522 1274
rect 542 1271 543 1275
rect 547 1271 548 1275
rect 614 1275 615 1279
rect 619 1275 620 1279
rect 652 1276 654 1306
rect 726 1302 727 1306
rect 731 1302 732 1306
rect 726 1301 732 1302
rect 710 1279 716 1280
rect 614 1274 620 1275
rect 650 1275 656 1276
rect 542 1270 548 1271
rect 311 1250 315 1251
rect 311 1245 315 1246
rect 359 1250 363 1251
rect 359 1245 363 1246
rect 415 1250 419 1251
rect 415 1245 419 1246
rect 439 1250 443 1251
rect 439 1245 443 1246
rect 519 1250 523 1251
rect 519 1245 523 1246
rect 302 1235 308 1236
rect 270 1230 276 1231
rect 278 1233 284 1234
rect 198 1228 204 1229
rect 214 1206 220 1207
rect 214 1202 215 1206
rect 219 1202 220 1206
rect 214 1201 220 1202
rect 190 1199 196 1200
rect 190 1195 191 1199
rect 195 1195 196 1199
rect 190 1194 196 1195
rect 216 1191 218 1201
rect 272 1200 274 1230
rect 278 1229 279 1233
rect 283 1229 284 1233
rect 302 1231 303 1235
rect 307 1231 308 1235
rect 360 1234 362 1245
rect 440 1234 442 1245
rect 494 1239 500 1240
rect 486 1235 492 1236
rect 302 1230 308 1231
rect 358 1233 364 1234
rect 278 1228 284 1229
rect 358 1229 359 1233
rect 363 1229 364 1233
rect 358 1228 364 1229
rect 438 1233 444 1234
rect 438 1229 439 1233
rect 443 1229 444 1233
rect 486 1231 487 1235
rect 491 1231 492 1235
rect 494 1235 495 1239
rect 499 1235 500 1239
rect 494 1234 500 1235
rect 520 1234 522 1245
rect 486 1230 492 1231
rect 438 1228 444 1229
rect 294 1206 300 1207
rect 294 1202 295 1206
rect 299 1202 300 1206
rect 294 1201 300 1202
rect 374 1206 380 1207
rect 374 1202 375 1206
rect 379 1202 380 1206
rect 374 1201 380 1202
rect 454 1206 460 1207
rect 454 1202 455 1206
rect 459 1202 460 1206
rect 454 1201 460 1202
rect 270 1199 276 1200
rect 270 1195 271 1199
rect 275 1195 276 1199
rect 270 1194 276 1195
rect 296 1191 298 1201
rect 346 1199 352 1200
rect 346 1195 347 1199
rect 351 1195 352 1199
rect 346 1194 352 1195
rect 111 1190 115 1191
rect 111 1185 115 1186
rect 159 1190 163 1191
rect 159 1185 163 1186
rect 215 1190 219 1191
rect 215 1185 219 1186
rect 239 1190 243 1191
rect 239 1185 243 1186
rect 295 1190 299 1191
rect 295 1185 299 1186
rect 327 1190 331 1191
rect 327 1185 331 1186
rect 112 1170 114 1185
rect 134 1183 140 1184
rect 134 1179 135 1183
rect 139 1179 140 1183
rect 160 1179 162 1185
rect 240 1179 242 1185
rect 258 1183 264 1184
rect 258 1179 259 1183
rect 263 1179 264 1183
rect 328 1179 330 1185
rect 134 1178 140 1179
rect 158 1178 164 1179
rect 110 1169 116 1170
rect 110 1165 111 1169
rect 115 1165 116 1169
rect 110 1164 116 1165
rect 136 1160 138 1178
rect 158 1174 159 1178
rect 163 1174 164 1178
rect 158 1173 164 1174
rect 238 1178 244 1179
rect 258 1178 264 1179
rect 326 1178 332 1179
rect 238 1174 239 1178
rect 243 1174 244 1178
rect 238 1173 244 1174
rect 134 1159 140 1160
rect 134 1155 135 1159
rect 139 1155 140 1159
rect 134 1154 140 1155
rect 110 1152 116 1153
rect 110 1148 111 1152
rect 115 1148 116 1152
rect 110 1147 116 1148
rect 142 1151 148 1152
rect 142 1147 143 1151
rect 147 1147 148 1151
rect 112 1127 114 1147
rect 142 1146 148 1147
rect 222 1151 228 1152
rect 222 1147 223 1151
rect 227 1147 228 1151
rect 260 1148 262 1178
rect 326 1174 327 1178
rect 331 1174 332 1178
rect 326 1173 332 1174
rect 310 1151 316 1152
rect 222 1146 228 1147
rect 258 1147 264 1148
rect 144 1127 146 1146
rect 224 1127 226 1146
rect 258 1143 259 1147
rect 263 1143 264 1147
rect 310 1147 311 1151
rect 315 1147 316 1151
rect 348 1148 350 1194
rect 376 1191 378 1201
rect 456 1191 458 1201
rect 375 1190 379 1191
rect 375 1185 379 1186
rect 423 1190 427 1191
rect 423 1185 427 1186
rect 455 1190 459 1191
rect 455 1185 459 1186
rect 354 1183 360 1184
rect 354 1179 355 1183
rect 359 1179 360 1183
rect 424 1179 426 1185
rect 488 1184 490 1230
rect 496 1200 498 1234
rect 518 1233 524 1234
rect 518 1229 519 1233
rect 523 1229 524 1233
rect 518 1228 524 1229
rect 534 1206 540 1207
rect 534 1202 535 1206
rect 539 1202 540 1206
rect 534 1201 540 1202
rect 494 1199 500 1200
rect 494 1195 495 1199
rect 499 1195 500 1199
rect 494 1194 500 1195
rect 536 1191 538 1201
rect 544 1200 546 1270
rect 616 1251 618 1274
rect 650 1271 651 1275
rect 655 1271 656 1275
rect 710 1275 711 1279
rect 715 1275 716 1279
rect 744 1276 746 1318
rect 751 1313 755 1314
rect 823 1318 827 1319
rect 838 1318 844 1319
rect 863 1318 867 1319
rect 823 1313 827 1314
rect 863 1313 867 1314
rect 778 1311 784 1312
rect 778 1307 779 1311
rect 783 1307 784 1311
rect 824 1307 826 1313
rect 892 1312 894 1327
rect 974 1326 975 1330
rect 979 1326 980 1330
rect 974 1325 980 1326
rect 976 1319 978 1325
rect 1000 1324 1002 1382
rect 1088 1375 1090 1386
rect 1118 1383 1119 1387
rect 1123 1383 1124 1387
rect 1198 1387 1199 1391
rect 1203 1387 1204 1391
rect 1326 1388 1327 1392
rect 1331 1388 1332 1392
rect 1366 1392 1367 1396
rect 1371 1392 1372 1396
rect 1366 1391 1372 1392
rect 1398 1395 1404 1396
rect 1398 1391 1399 1395
rect 1403 1391 1404 1395
rect 1326 1387 1332 1388
rect 1198 1386 1204 1387
rect 1118 1382 1124 1383
rect 1200 1375 1202 1386
rect 1328 1375 1330 1387
rect 1071 1374 1075 1375
rect 1071 1369 1075 1370
rect 1087 1374 1091 1375
rect 1087 1369 1091 1370
rect 1183 1374 1187 1375
rect 1183 1369 1187 1370
rect 1199 1374 1203 1375
rect 1199 1369 1203 1370
rect 1271 1374 1275 1375
rect 1271 1369 1275 1370
rect 1327 1374 1331 1375
rect 1368 1371 1370 1391
rect 1398 1390 1404 1391
rect 1400 1371 1402 1390
rect 1327 1369 1331 1370
rect 1367 1370 1371 1371
rect 1062 1359 1068 1360
rect 1062 1355 1063 1359
rect 1067 1355 1068 1359
rect 1072 1358 1074 1369
rect 1174 1359 1180 1360
rect 1062 1354 1068 1355
rect 1070 1357 1076 1358
rect 1064 1324 1066 1354
rect 1070 1353 1071 1357
rect 1075 1353 1076 1357
rect 1174 1355 1175 1359
rect 1179 1355 1180 1359
rect 1184 1358 1186 1369
rect 1262 1359 1268 1360
rect 1174 1354 1180 1355
rect 1182 1357 1188 1358
rect 1070 1352 1076 1353
rect 1086 1330 1092 1331
rect 1086 1326 1087 1330
rect 1091 1326 1092 1330
rect 1086 1325 1092 1326
rect 998 1323 1004 1324
rect 998 1319 999 1323
rect 1003 1319 1004 1323
rect 911 1318 915 1319
rect 911 1313 915 1314
rect 975 1318 979 1319
rect 975 1313 979 1314
rect 991 1318 995 1319
rect 998 1318 1004 1319
rect 1062 1323 1068 1324
rect 1062 1319 1063 1323
rect 1067 1319 1068 1323
rect 1088 1319 1090 1325
rect 1176 1324 1178 1354
rect 1182 1353 1183 1357
rect 1187 1353 1188 1357
rect 1262 1355 1263 1359
rect 1267 1355 1268 1359
rect 1272 1358 1274 1369
rect 1294 1359 1300 1360
rect 1262 1354 1268 1355
rect 1270 1357 1276 1358
rect 1182 1352 1188 1353
rect 1198 1330 1204 1331
rect 1198 1326 1199 1330
rect 1203 1326 1204 1330
rect 1198 1325 1204 1326
rect 1174 1323 1180 1324
rect 1174 1319 1175 1323
rect 1179 1319 1180 1323
rect 1200 1319 1202 1325
rect 1264 1324 1266 1354
rect 1270 1353 1271 1357
rect 1275 1353 1276 1357
rect 1294 1355 1295 1359
rect 1299 1355 1300 1359
rect 1328 1357 1330 1369
rect 1367 1365 1371 1366
rect 1399 1370 1403 1371
rect 1399 1365 1403 1366
rect 1294 1354 1300 1355
rect 1326 1356 1332 1357
rect 1270 1352 1276 1353
rect 1296 1333 1298 1354
rect 1326 1352 1327 1356
rect 1331 1352 1332 1356
rect 1368 1353 1370 1365
rect 1400 1354 1402 1365
rect 1408 1357 1410 1422
rect 1414 1418 1415 1422
rect 1419 1418 1420 1422
rect 1414 1417 1420 1418
rect 1436 1392 1438 1422
rect 1470 1418 1471 1422
rect 1475 1418 1476 1422
rect 1470 1417 1476 1418
rect 1454 1395 1460 1396
rect 1434 1391 1440 1392
rect 1434 1387 1435 1391
rect 1439 1387 1440 1391
rect 1454 1391 1455 1395
rect 1459 1391 1460 1395
rect 1504 1392 1506 1422
rect 1534 1418 1535 1422
rect 1539 1418 1540 1422
rect 1534 1417 1540 1418
rect 1518 1395 1524 1396
rect 1454 1390 1460 1391
rect 1502 1391 1508 1392
rect 1434 1386 1440 1387
rect 1456 1371 1458 1390
rect 1502 1387 1503 1391
rect 1507 1387 1508 1391
rect 1518 1391 1519 1395
rect 1523 1391 1524 1395
rect 1556 1392 1558 1422
rect 1622 1418 1623 1422
rect 1627 1418 1628 1422
rect 1622 1417 1628 1418
rect 1606 1395 1612 1396
rect 1518 1390 1524 1391
rect 1554 1391 1560 1392
rect 1502 1386 1508 1387
rect 1520 1371 1522 1390
rect 1554 1387 1555 1391
rect 1559 1387 1560 1391
rect 1606 1391 1607 1395
rect 1611 1391 1612 1395
rect 1644 1392 1646 1422
rect 1718 1418 1719 1422
rect 1723 1418 1724 1422
rect 1718 1417 1724 1418
rect 1822 1422 1828 1423
rect 1822 1418 1823 1422
rect 1827 1418 1828 1422
rect 1822 1417 1828 1418
rect 1702 1395 1708 1396
rect 1606 1390 1612 1391
rect 1642 1391 1648 1392
rect 1554 1386 1560 1387
rect 1608 1371 1610 1390
rect 1642 1387 1643 1391
rect 1647 1387 1648 1391
rect 1702 1391 1703 1395
rect 1707 1391 1708 1395
rect 1702 1390 1708 1391
rect 1806 1395 1812 1396
rect 1806 1391 1807 1395
rect 1811 1391 1812 1395
rect 1840 1392 1842 1434
rect 1911 1429 1915 1430
rect 1927 1434 1931 1435
rect 1927 1429 1931 1430
rect 1999 1434 2003 1435
rect 2006 1431 2007 1435
rect 2011 1431 2012 1435
rect 2006 1430 2012 1431
rect 2023 1434 2027 1435
rect 1999 1429 2003 1430
rect 2023 1429 2027 1430
rect 1928 1423 1930 1429
rect 2024 1423 2026 1429
rect 1926 1422 1932 1423
rect 1926 1418 1927 1422
rect 1931 1418 1932 1422
rect 1926 1417 1932 1418
rect 2022 1422 2028 1423
rect 2022 1418 2023 1422
rect 2027 1418 2028 1422
rect 2022 1417 2028 1418
rect 1910 1395 1916 1396
rect 1806 1390 1812 1391
rect 1838 1391 1844 1392
rect 1642 1386 1648 1387
rect 1704 1371 1706 1390
rect 1808 1371 1810 1390
rect 1838 1387 1839 1391
rect 1843 1387 1844 1391
rect 1910 1391 1911 1395
rect 1915 1391 1916 1395
rect 2006 1395 2012 1396
rect 1910 1390 1916 1391
rect 1934 1391 1940 1392
rect 1838 1386 1844 1387
rect 1912 1371 1914 1390
rect 1934 1387 1935 1391
rect 1939 1387 1940 1391
rect 2006 1391 2007 1395
rect 2011 1391 2012 1395
rect 2044 1392 2046 1442
rect 2088 1435 2090 1449
rect 2144 1448 2146 1478
rect 2150 1477 2151 1481
rect 2155 1477 2156 1481
rect 2222 1479 2223 1483
rect 2227 1479 2228 1483
rect 2232 1482 2234 1493
rect 2268 1484 2270 1550
rect 2326 1546 2327 1550
rect 2331 1546 2332 1550
rect 2326 1545 2332 1546
rect 2310 1523 2316 1524
rect 2310 1519 2311 1523
rect 2315 1519 2316 1523
rect 2344 1520 2346 1558
rect 2407 1557 2411 1558
rect 2447 1562 2451 1563
rect 2447 1557 2451 1558
rect 2382 1555 2388 1556
rect 2382 1551 2383 1555
rect 2387 1551 2388 1555
rect 2408 1551 2410 1557
rect 2464 1556 2466 1602
rect 2526 1601 2527 1605
rect 2531 1601 2532 1605
rect 2526 1600 2532 1601
rect 2582 1604 2588 1605
rect 2582 1600 2583 1604
rect 2587 1600 2588 1604
rect 2582 1599 2588 1600
rect 2582 1587 2588 1588
rect 2582 1583 2583 1587
rect 2587 1583 2588 1587
rect 2582 1582 2588 1583
rect 2542 1578 2548 1579
rect 2542 1574 2543 1578
rect 2547 1574 2548 1578
rect 2542 1573 2548 1574
rect 2544 1563 2546 1573
rect 2558 1571 2564 1572
rect 2558 1567 2559 1571
rect 2563 1567 2564 1571
rect 2558 1566 2564 1567
rect 2487 1562 2491 1563
rect 2487 1557 2491 1558
rect 2543 1562 2547 1563
rect 2543 1557 2547 1558
rect 2462 1555 2468 1556
rect 2462 1551 2463 1555
rect 2467 1551 2468 1555
rect 2488 1551 2490 1557
rect 2534 1555 2540 1556
rect 2534 1551 2535 1555
rect 2539 1551 2540 1555
rect 2544 1551 2546 1557
rect 2382 1550 2388 1551
rect 2406 1550 2412 1551
rect 2462 1550 2468 1551
rect 2486 1550 2492 1551
rect 2534 1550 2540 1551
rect 2542 1550 2548 1551
rect 2384 1532 2386 1550
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2486 1546 2487 1550
rect 2491 1546 2492 1550
rect 2486 1545 2492 1546
rect 2382 1531 2388 1532
rect 2382 1527 2383 1531
rect 2387 1527 2388 1531
rect 2382 1526 2388 1527
rect 2390 1523 2396 1524
rect 2310 1518 2316 1519
rect 2342 1519 2348 1520
rect 2312 1499 2314 1518
rect 2342 1515 2343 1519
rect 2347 1515 2348 1519
rect 2390 1519 2391 1523
rect 2395 1519 2396 1523
rect 2470 1523 2476 1524
rect 2390 1518 2396 1519
rect 2414 1519 2420 1520
rect 2342 1514 2348 1515
rect 2392 1499 2394 1518
rect 2414 1515 2415 1519
rect 2419 1515 2420 1519
rect 2470 1519 2471 1523
rect 2475 1519 2476 1523
rect 2470 1518 2476 1519
rect 2526 1523 2532 1524
rect 2526 1519 2527 1523
rect 2531 1519 2532 1523
rect 2526 1518 2532 1519
rect 2414 1514 2420 1515
rect 2311 1498 2315 1499
rect 2311 1493 2315 1494
rect 2391 1498 2395 1499
rect 2391 1493 2395 1494
rect 2282 1487 2288 1488
rect 2266 1483 2272 1484
rect 2222 1478 2228 1479
rect 2230 1481 2236 1482
rect 2150 1476 2156 1477
rect 2166 1454 2172 1455
rect 2166 1450 2167 1454
rect 2171 1450 2172 1454
rect 2166 1449 2172 1450
rect 2142 1447 2148 1448
rect 2142 1443 2143 1447
rect 2147 1443 2148 1447
rect 2142 1442 2148 1443
rect 2134 1435 2140 1436
rect 2168 1435 2170 1449
rect 2224 1448 2226 1478
rect 2230 1477 2231 1481
rect 2235 1477 2236 1481
rect 2266 1479 2267 1483
rect 2271 1479 2272 1483
rect 2282 1483 2283 1487
rect 2287 1483 2288 1487
rect 2282 1482 2288 1483
rect 2312 1482 2314 1493
rect 2354 1487 2360 1488
rect 2354 1483 2355 1487
rect 2359 1483 2360 1487
rect 2354 1482 2360 1483
rect 2392 1482 2394 1493
rect 2266 1478 2272 1479
rect 2230 1476 2236 1477
rect 2246 1454 2252 1455
rect 2246 1450 2247 1454
rect 2251 1450 2252 1454
rect 2246 1449 2252 1450
rect 2222 1447 2228 1448
rect 2222 1443 2223 1447
rect 2227 1443 2228 1447
rect 2222 1442 2228 1443
rect 2248 1435 2250 1449
rect 2087 1434 2091 1435
rect 2087 1429 2091 1430
rect 2119 1434 2123 1435
rect 2134 1431 2135 1435
rect 2139 1431 2140 1435
rect 2134 1430 2140 1431
rect 2167 1434 2171 1435
rect 2119 1429 2123 1430
rect 2094 1427 2100 1428
rect 2094 1423 2095 1427
rect 2099 1423 2100 1427
rect 2120 1423 2122 1429
rect 2094 1422 2100 1423
rect 2118 1422 2124 1423
rect 2096 1404 2098 1422
rect 2118 1418 2119 1422
rect 2123 1418 2124 1422
rect 2118 1417 2124 1418
rect 2094 1403 2100 1404
rect 2094 1399 2095 1403
rect 2099 1399 2100 1403
rect 2094 1398 2100 1399
rect 2102 1395 2108 1396
rect 2006 1390 2012 1391
rect 2042 1391 2048 1392
rect 1934 1386 1940 1387
rect 1455 1370 1459 1371
rect 1455 1365 1459 1366
rect 1519 1370 1523 1371
rect 1519 1365 1523 1366
rect 1543 1370 1547 1371
rect 1543 1365 1547 1366
rect 1607 1370 1611 1371
rect 1607 1365 1611 1366
rect 1631 1370 1635 1371
rect 1631 1365 1635 1366
rect 1703 1370 1707 1371
rect 1703 1365 1707 1366
rect 1719 1370 1723 1371
rect 1719 1365 1723 1366
rect 1807 1370 1811 1371
rect 1807 1365 1811 1366
rect 1887 1370 1891 1371
rect 1887 1365 1891 1366
rect 1911 1370 1915 1371
rect 1911 1365 1915 1366
rect 1407 1356 1411 1357
rect 1398 1353 1404 1354
rect 1326 1351 1332 1352
rect 1366 1352 1372 1353
rect 1366 1348 1367 1352
rect 1371 1348 1372 1352
rect 1398 1349 1399 1353
rect 1403 1349 1404 1353
rect 1407 1351 1411 1352
rect 1446 1355 1452 1356
rect 1446 1351 1447 1355
rect 1451 1351 1452 1355
rect 1456 1354 1458 1365
rect 1534 1355 1540 1356
rect 1446 1350 1452 1351
rect 1454 1353 1460 1354
rect 1398 1348 1404 1349
rect 1366 1347 1372 1348
rect 1326 1339 1332 1340
rect 1326 1335 1327 1339
rect 1331 1335 1332 1339
rect 1326 1334 1332 1335
rect 1366 1335 1372 1336
rect 1295 1332 1299 1333
rect 1286 1330 1292 1331
rect 1286 1326 1287 1330
rect 1291 1326 1292 1330
rect 1295 1327 1299 1328
rect 1286 1325 1292 1326
rect 1262 1323 1268 1324
rect 1262 1319 1263 1323
rect 1267 1319 1268 1323
rect 1288 1319 1290 1325
rect 1306 1319 1312 1320
rect 1328 1319 1330 1334
rect 1366 1331 1367 1335
rect 1371 1331 1372 1335
rect 1366 1330 1372 1331
rect 1062 1318 1068 1319
rect 1071 1318 1075 1319
rect 991 1313 995 1314
rect 1071 1313 1075 1314
rect 1087 1318 1091 1319
rect 1087 1313 1091 1314
rect 1151 1318 1155 1319
rect 1174 1318 1180 1319
rect 1199 1318 1203 1319
rect 1151 1313 1155 1314
rect 1199 1313 1203 1314
rect 1231 1318 1235 1319
rect 1262 1318 1268 1319
rect 1287 1318 1291 1319
rect 1231 1313 1235 1314
rect 1306 1315 1307 1319
rect 1311 1315 1312 1319
rect 1306 1314 1312 1315
rect 1327 1318 1331 1319
rect 1287 1313 1291 1314
rect 890 1311 896 1312
rect 890 1307 891 1311
rect 895 1307 896 1311
rect 912 1307 914 1313
rect 930 1311 936 1312
rect 930 1307 931 1311
rect 935 1307 936 1311
rect 992 1307 994 1313
rect 1010 1311 1016 1312
rect 1010 1307 1011 1311
rect 1015 1307 1016 1311
rect 1072 1307 1074 1313
rect 1110 1311 1116 1312
rect 1110 1307 1111 1311
rect 1115 1307 1116 1311
rect 1152 1307 1154 1313
rect 1170 1311 1176 1312
rect 1170 1307 1171 1311
rect 1175 1307 1176 1311
rect 1232 1307 1234 1313
rect 1250 1311 1256 1312
rect 1250 1307 1251 1311
rect 1255 1307 1256 1311
rect 1288 1307 1290 1313
rect 778 1306 784 1307
rect 822 1306 828 1307
rect 890 1306 896 1307
rect 910 1306 916 1307
rect 930 1306 936 1307
rect 990 1306 996 1307
rect 1010 1306 1016 1307
rect 1070 1306 1076 1307
rect 1110 1306 1116 1307
rect 1150 1306 1156 1307
rect 1170 1306 1176 1307
rect 1230 1306 1236 1307
rect 1250 1306 1256 1307
rect 1286 1306 1292 1307
rect 710 1274 716 1275
rect 742 1275 748 1276
rect 650 1270 656 1271
rect 712 1251 714 1274
rect 742 1271 743 1275
rect 747 1271 748 1275
rect 742 1270 748 1271
rect 599 1250 603 1251
rect 599 1245 603 1246
rect 615 1250 619 1251
rect 615 1245 619 1246
rect 671 1250 675 1251
rect 671 1245 675 1246
rect 711 1250 715 1251
rect 711 1245 715 1246
rect 743 1250 747 1251
rect 743 1245 747 1246
rect 600 1234 602 1245
rect 662 1235 668 1236
rect 598 1233 604 1234
rect 598 1229 599 1233
rect 603 1229 604 1233
rect 662 1231 663 1235
rect 667 1231 668 1235
rect 672 1234 674 1245
rect 734 1235 740 1236
rect 662 1230 668 1231
rect 670 1233 676 1234
rect 598 1228 604 1229
rect 614 1206 620 1207
rect 614 1202 615 1206
rect 619 1202 620 1206
rect 614 1201 620 1202
rect 542 1199 548 1200
rect 542 1195 543 1199
rect 547 1195 548 1199
rect 542 1194 548 1195
rect 616 1191 618 1201
rect 664 1200 666 1230
rect 670 1229 671 1233
rect 675 1229 676 1233
rect 734 1231 735 1235
rect 739 1231 740 1235
rect 744 1234 746 1245
rect 780 1236 782 1306
rect 822 1302 823 1306
rect 827 1302 828 1306
rect 822 1301 828 1302
rect 910 1302 911 1306
rect 915 1302 916 1306
rect 910 1301 916 1302
rect 806 1279 812 1280
rect 806 1275 807 1279
rect 811 1275 812 1279
rect 806 1274 812 1275
rect 894 1279 900 1280
rect 894 1275 895 1279
rect 899 1275 900 1279
rect 932 1276 934 1306
rect 990 1302 991 1306
rect 995 1302 996 1306
rect 990 1301 996 1302
rect 974 1279 980 1280
rect 894 1274 900 1275
rect 930 1275 936 1276
rect 808 1251 810 1274
rect 896 1251 898 1274
rect 930 1271 931 1275
rect 935 1271 936 1275
rect 974 1275 975 1279
rect 979 1275 980 1279
rect 1012 1276 1014 1306
rect 1070 1302 1071 1306
rect 1075 1302 1076 1306
rect 1070 1301 1076 1302
rect 1112 1280 1114 1306
rect 1150 1302 1151 1306
rect 1155 1302 1156 1306
rect 1150 1301 1156 1302
rect 1054 1279 1060 1280
rect 974 1274 980 1275
rect 1010 1275 1016 1276
rect 930 1270 936 1271
rect 976 1251 978 1274
rect 1010 1271 1011 1275
rect 1015 1271 1016 1275
rect 1054 1275 1055 1279
rect 1059 1275 1060 1279
rect 1054 1274 1060 1275
rect 1110 1279 1116 1280
rect 1110 1275 1111 1279
rect 1115 1275 1116 1279
rect 1110 1274 1116 1275
rect 1134 1279 1140 1280
rect 1134 1275 1135 1279
rect 1139 1275 1140 1279
rect 1172 1276 1174 1306
rect 1230 1302 1231 1306
rect 1235 1302 1236 1306
rect 1230 1301 1236 1302
rect 1214 1279 1220 1280
rect 1134 1274 1140 1275
rect 1170 1275 1176 1276
rect 1010 1270 1016 1271
rect 1056 1251 1058 1274
rect 1136 1251 1138 1274
rect 1170 1271 1171 1275
rect 1175 1271 1176 1275
rect 1214 1275 1215 1279
rect 1219 1275 1220 1279
rect 1252 1276 1254 1306
rect 1286 1302 1287 1306
rect 1291 1302 1292 1306
rect 1286 1301 1292 1302
rect 1270 1279 1276 1280
rect 1214 1274 1220 1275
rect 1250 1275 1256 1276
rect 1170 1270 1176 1271
rect 1216 1251 1218 1274
rect 1250 1271 1251 1275
rect 1255 1271 1256 1275
rect 1270 1275 1271 1279
rect 1275 1275 1276 1279
rect 1308 1276 1310 1314
rect 1327 1313 1331 1314
rect 1328 1298 1330 1313
rect 1368 1311 1370 1330
rect 1414 1326 1420 1327
rect 1414 1322 1415 1326
rect 1419 1322 1420 1326
rect 1414 1321 1420 1322
rect 1416 1311 1418 1321
rect 1448 1320 1450 1350
rect 1454 1349 1455 1353
rect 1459 1349 1460 1353
rect 1534 1351 1535 1355
rect 1539 1351 1540 1355
rect 1544 1354 1546 1365
rect 1622 1355 1628 1356
rect 1534 1350 1540 1351
rect 1542 1353 1548 1354
rect 1454 1348 1460 1349
rect 1470 1326 1476 1327
rect 1470 1322 1471 1326
rect 1475 1322 1476 1326
rect 1470 1321 1476 1322
rect 1446 1319 1452 1320
rect 1446 1315 1447 1319
rect 1451 1315 1452 1319
rect 1446 1314 1452 1315
rect 1472 1311 1474 1321
rect 1536 1320 1538 1350
rect 1542 1349 1543 1353
rect 1547 1349 1548 1353
rect 1622 1351 1623 1355
rect 1627 1351 1628 1355
rect 1632 1354 1634 1365
rect 1710 1355 1716 1356
rect 1622 1350 1628 1351
rect 1630 1353 1636 1354
rect 1542 1348 1548 1349
rect 1558 1326 1564 1327
rect 1558 1322 1559 1326
rect 1563 1322 1564 1326
rect 1558 1321 1564 1322
rect 1534 1319 1540 1320
rect 1534 1315 1535 1319
rect 1539 1315 1540 1319
rect 1534 1314 1540 1315
rect 1560 1311 1562 1321
rect 1624 1320 1626 1350
rect 1630 1349 1631 1353
rect 1635 1349 1636 1353
rect 1710 1351 1711 1355
rect 1715 1351 1716 1355
rect 1720 1354 1722 1365
rect 1751 1356 1755 1357
rect 1710 1350 1716 1351
rect 1718 1353 1724 1354
rect 1630 1348 1636 1349
rect 1646 1326 1652 1327
rect 1646 1322 1647 1326
rect 1651 1322 1652 1326
rect 1646 1321 1652 1322
rect 1622 1319 1628 1320
rect 1622 1315 1623 1319
rect 1627 1315 1628 1319
rect 1622 1314 1628 1315
rect 1648 1311 1650 1321
rect 1712 1320 1714 1350
rect 1718 1349 1719 1353
rect 1723 1349 1724 1353
rect 1750 1351 1751 1356
rect 1755 1351 1756 1356
rect 1808 1354 1810 1365
rect 1838 1355 1844 1356
rect 1750 1350 1756 1351
rect 1806 1353 1812 1354
rect 1718 1348 1724 1349
rect 1806 1349 1807 1353
rect 1811 1349 1812 1353
rect 1838 1351 1839 1355
rect 1843 1351 1844 1355
rect 1888 1354 1890 1365
rect 1838 1350 1844 1351
rect 1886 1353 1892 1354
rect 1806 1348 1812 1349
rect 1734 1326 1740 1327
rect 1734 1322 1735 1326
rect 1739 1322 1740 1326
rect 1734 1321 1740 1322
rect 1822 1326 1828 1327
rect 1822 1322 1823 1326
rect 1827 1322 1828 1326
rect 1822 1321 1828 1322
rect 1710 1319 1716 1320
rect 1710 1315 1711 1319
rect 1715 1315 1716 1319
rect 1710 1314 1716 1315
rect 1736 1311 1738 1321
rect 1824 1311 1826 1321
rect 1367 1310 1371 1311
rect 1367 1305 1371 1306
rect 1415 1310 1419 1311
rect 1415 1305 1419 1306
rect 1471 1310 1475 1311
rect 1471 1305 1475 1306
rect 1559 1310 1563 1311
rect 1559 1305 1563 1306
rect 1647 1310 1651 1311
rect 1647 1305 1651 1306
rect 1671 1310 1675 1311
rect 1671 1305 1675 1306
rect 1735 1310 1739 1311
rect 1735 1305 1739 1306
rect 1767 1310 1771 1311
rect 1823 1310 1827 1311
rect 1767 1305 1771 1306
rect 1790 1307 1796 1308
rect 1326 1297 1332 1298
rect 1326 1293 1327 1297
rect 1331 1293 1332 1297
rect 1326 1292 1332 1293
rect 1368 1290 1370 1305
rect 1672 1299 1674 1305
rect 1768 1299 1770 1305
rect 1790 1303 1791 1307
rect 1795 1303 1796 1307
rect 1823 1305 1827 1306
rect 1840 1304 1842 1350
rect 1886 1349 1887 1353
rect 1891 1349 1892 1353
rect 1886 1348 1892 1349
rect 1902 1326 1908 1327
rect 1902 1322 1903 1326
rect 1907 1322 1908 1326
rect 1902 1321 1908 1322
rect 1904 1311 1906 1321
rect 1936 1320 1938 1386
rect 2008 1371 2010 1390
rect 2042 1387 2043 1391
rect 2047 1387 2048 1391
rect 2102 1391 2103 1395
rect 2107 1391 2108 1395
rect 2136 1392 2138 1430
rect 2167 1429 2171 1430
rect 2215 1434 2219 1435
rect 2247 1434 2251 1435
rect 2215 1429 2219 1430
rect 2238 1431 2244 1432
rect 2216 1423 2218 1429
rect 2238 1427 2239 1431
rect 2243 1427 2244 1431
rect 2247 1429 2251 1430
rect 2284 1428 2286 1482
rect 2310 1481 2316 1482
rect 2310 1477 2311 1481
rect 2315 1477 2316 1481
rect 2310 1476 2316 1477
rect 2326 1454 2332 1455
rect 2326 1450 2327 1454
rect 2331 1450 2332 1454
rect 2326 1449 2332 1450
rect 2328 1435 2330 1449
rect 2356 1448 2358 1482
rect 2390 1481 2396 1482
rect 2390 1477 2391 1481
rect 2395 1477 2396 1481
rect 2390 1476 2396 1477
rect 2406 1454 2412 1455
rect 2406 1450 2407 1454
rect 2411 1450 2412 1454
rect 2406 1449 2412 1450
rect 2354 1447 2360 1448
rect 2354 1443 2355 1447
rect 2359 1443 2360 1447
rect 2354 1442 2360 1443
rect 2408 1435 2410 1449
rect 2416 1448 2418 1514
rect 2472 1499 2474 1518
rect 2528 1499 2530 1518
rect 2471 1498 2475 1499
rect 2471 1493 2475 1494
rect 2527 1498 2531 1499
rect 2527 1493 2531 1494
rect 2472 1482 2474 1493
rect 2518 1483 2524 1484
rect 2470 1481 2476 1482
rect 2470 1477 2471 1481
rect 2475 1477 2476 1481
rect 2518 1479 2519 1483
rect 2523 1479 2524 1483
rect 2528 1482 2530 1493
rect 2536 1488 2538 1550
rect 2542 1546 2543 1550
rect 2547 1546 2548 1550
rect 2542 1545 2548 1546
rect 2560 1520 2562 1566
rect 2584 1563 2586 1582
rect 2583 1562 2587 1563
rect 2583 1557 2587 1558
rect 2584 1542 2586 1557
rect 2582 1541 2588 1542
rect 2582 1537 2583 1541
rect 2587 1537 2588 1541
rect 2582 1536 2588 1537
rect 2582 1524 2588 1525
rect 2582 1520 2583 1524
rect 2587 1520 2588 1524
rect 2558 1519 2564 1520
rect 2582 1519 2588 1520
rect 2558 1515 2559 1519
rect 2563 1515 2564 1519
rect 2558 1514 2564 1515
rect 2584 1499 2586 1519
rect 2583 1498 2587 1499
rect 2583 1493 2587 1494
rect 2534 1487 2540 1488
rect 2534 1483 2535 1487
rect 2539 1483 2540 1487
rect 2534 1482 2540 1483
rect 2518 1478 2524 1479
rect 2526 1481 2532 1482
rect 2584 1481 2586 1493
rect 2470 1476 2476 1477
rect 2486 1454 2492 1455
rect 2486 1450 2487 1454
rect 2491 1450 2492 1454
rect 2486 1449 2492 1450
rect 2414 1447 2420 1448
rect 2414 1443 2415 1447
rect 2419 1443 2420 1447
rect 2414 1442 2420 1443
rect 2488 1435 2490 1449
rect 2520 1448 2522 1478
rect 2526 1477 2527 1481
rect 2531 1477 2532 1481
rect 2526 1476 2532 1477
rect 2582 1480 2588 1481
rect 2582 1476 2583 1480
rect 2587 1476 2588 1480
rect 2582 1475 2588 1476
rect 2582 1463 2588 1464
rect 2582 1459 2583 1463
rect 2587 1459 2588 1463
rect 2582 1458 2588 1459
rect 2542 1454 2548 1455
rect 2542 1450 2543 1454
rect 2547 1450 2548 1454
rect 2542 1449 2548 1450
rect 2518 1447 2524 1448
rect 2518 1443 2519 1447
rect 2523 1443 2524 1447
rect 2518 1442 2524 1443
rect 2544 1435 2546 1449
rect 2558 1439 2564 1440
rect 2558 1435 2559 1439
rect 2563 1435 2564 1439
rect 2584 1435 2586 1458
rect 2303 1434 2307 1435
rect 2303 1429 2307 1430
rect 2327 1434 2331 1435
rect 2327 1429 2331 1430
rect 2391 1434 2395 1435
rect 2391 1429 2395 1430
rect 2407 1434 2411 1435
rect 2407 1429 2411 1430
rect 2479 1434 2483 1435
rect 2479 1429 2483 1430
rect 2487 1434 2491 1435
rect 2487 1429 2491 1430
rect 2543 1434 2547 1435
rect 2558 1434 2564 1435
rect 2583 1434 2587 1435
rect 2543 1429 2547 1430
rect 2238 1426 2244 1427
rect 2282 1427 2288 1428
rect 2214 1422 2220 1423
rect 2214 1418 2215 1422
rect 2219 1418 2220 1422
rect 2214 1417 2220 1418
rect 2198 1395 2204 1396
rect 2102 1390 2108 1391
rect 2134 1391 2140 1392
rect 2042 1386 2048 1387
rect 2104 1371 2106 1390
rect 2134 1387 2135 1391
rect 2139 1387 2140 1391
rect 2198 1391 2199 1395
rect 2203 1391 2204 1395
rect 2198 1390 2204 1391
rect 2134 1386 2140 1387
rect 2200 1371 2202 1390
rect 1967 1370 1971 1371
rect 1967 1365 1971 1366
rect 2007 1370 2011 1371
rect 2007 1365 2011 1366
rect 2047 1370 2051 1371
rect 2047 1365 2051 1366
rect 2103 1370 2107 1371
rect 2103 1365 2107 1366
rect 2127 1370 2131 1371
rect 2127 1365 2131 1366
rect 2199 1370 2203 1371
rect 2199 1365 2203 1366
rect 2207 1370 2211 1371
rect 2207 1365 2211 1366
rect 1968 1354 1970 1365
rect 2038 1355 2044 1356
rect 1966 1353 1972 1354
rect 1966 1349 1967 1353
rect 1971 1349 1972 1353
rect 2038 1351 2039 1355
rect 2043 1351 2044 1355
rect 2048 1354 2050 1365
rect 2118 1355 2124 1356
rect 2038 1350 2044 1351
rect 2046 1353 2052 1354
rect 1966 1348 1972 1349
rect 1982 1326 1988 1327
rect 1982 1322 1983 1326
rect 1987 1322 1988 1326
rect 1982 1321 1988 1322
rect 1934 1319 1940 1320
rect 1934 1315 1935 1319
rect 1939 1315 1940 1319
rect 1934 1314 1940 1315
rect 1974 1319 1980 1320
rect 1974 1315 1975 1319
rect 1979 1315 1980 1319
rect 1974 1314 1980 1315
rect 1863 1310 1867 1311
rect 1863 1305 1867 1306
rect 1903 1310 1907 1311
rect 1903 1305 1907 1306
rect 1959 1310 1963 1311
rect 1959 1305 1963 1306
rect 1790 1302 1796 1303
rect 1838 1303 1844 1304
rect 1670 1298 1676 1299
rect 1670 1294 1671 1298
rect 1675 1294 1676 1298
rect 1670 1293 1676 1294
rect 1766 1298 1772 1299
rect 1766 1294 1767 1298
rect 1771 1294 1772 1298
rect 1766 1293 1772 1294
rect 1366 1289 1372 1290
rect 1366 1285 1367 1289
rect 1371 1285 1372 1289
rect 1366 1284 1372 1285
rect 1326 1280 1332 1281
rect 1326 1276 1327 1280
rect 1331 1276 1332 1280
rect 1270 1274 1276 1275
rect 1306 1275 1312 1276
rect 1326 1275 1332 1276
rect 1250 1270 1256 1271
rect 1272 1251 1274 1274
rect 1306 1271 1307 1275
rect 1311 1271 1312 1275
rect 1306 1270 1312 1271
rect 1328 1251 1330 1275
rect 1366 1272 1372 1273
rect 1366 1268 1367 1272
rect 1371 1268 1372 1272
rect 1366 1267 1372 1268
rect 1654 1271 1660 1272
rect 1654 1267 1655 1271
rect 1659 1267 1660 1271
rect 1368 1255 1370 1267
rect 1654 1266 1660 1267
rect 1750 1271 1756 1272
rect 1750 1267 1751 1271
rect 1755 1267 1756 1271
rect 1750 1266 1756 1267
rect 1656 1255 1658 1266
rect 1662 1263 1668 1264
rect 1662 1259 1663 1263
rect 1667 1259 1668 1263
rect 1662 1258 1668 1259
rect 1367 1254 1371 1255
rect 807 1250 811 1251
rect 807 1245 811 1246
rect 815 1250 819 1251
rect 815 1245 819 1246
rect 895 1250 899 1251
rect 895 1245 899 1246
rect 975 1250 979 1251
rect 975 1245 979 1246
rect 1055 1250 1059 1251
rect 1055 1245 1059 1246
rect 1135 1250 1139 1251
rect 1135 1245 1139 1246
rect 1215 1250 1219 1251
rect 1215 1245 1219 1246
rect 1271 1250 1275 1251
rect 1271 1245 1275 1246
rect 1327 1250 1331 1251
rect 1367 1249 1371 1250
rect 1495 1254 1499 1255
rect 1495 1249 1499 1250
rect 1559 1254 1563 1255
rect 1559 1249 1563 1250
rect 1623 1254 1627 1255
rect 1623 1249 1627 1250
rect 1655 1254 1659 1255
rect 1655 1249 1659 1250
rect 1327 1245 1331 1246
rect 778 1235 784 1236
rect 734 1230 740 1231
rect 742 1233 748 1234
rect 670 1228 676 1229
rect 686 1206 692 1207
rect 686 1202 687 1206
rect 691 1202 692 1206
rect 686 1201 692 1202
rect 662 1199 668 1200
rect 662 1195 663 1199
rect 667 1195 668 1199
rect 662 1194 668 1195
rect 688 1191 690 1201
rect 736 1200 738 1230
rect 742 1229 743 1233
rect 747 1229 748 1233
rect 778 1231 779 1235
rect 783 1231 784 1235
rect 816 1234 818 1245
rect 822 1243 828 1244
rect 822 1239 823 1243
rect 827 1239 828 1243
rect 822 1238 828 1239
rect 778 1230 784 1231
rect 814 1233 820 1234
rect 742 1228 748 1229
rect 814 1229 815 1233
rect 819 1229 820 1233
rect 814 1228 820 1229
rect 758 1206 764 1207
rect 758 1202 759 1206
rect 763 1202 764 1206
rect 758 1201 764 1202
rect 734 1199 740 1200
rect 734 1195 735 1199
rect 739 1195 740 1199
rect 734 1194 740 1195
rect 760 1191 762 1201
rect 824 1200 826 1238
rect 846 1235 852 1236
rect 846 1231 847 1235
rect 851 1231 852 1235
rect 896 1234 898 1245
rect 846 1230 852 1231
rect 894 1233 900 1234
rect 1328 1233 1330 1245
rect 1368 1237 1370 1249
rect 1496 1238 1498 1249
rect 1518 1247 1524 1248
rect 1518 1243 1519 1247
rect 1523 1243 1524 1247
rect 1518 1242 1524 1243
rect 1494 1237 1500 1238
rect 1366 1236 1372 1237
rect 830 1206 836 1207
rect 830 1202 831 1206
rect 835 1202 836 1206
rect 830 1201 836 1202
rect 822 1199 828 1200
rect 822 1195 823 1199
rect 827 1195 828 1199
rect 822 1194 828 1195
rect 832 1191 834 1201
rect 848 1192 850 1230
rect 894 1229 895 1233
rect 899 1229 900 1233
rect 894 1228 900 1229
rect 1326 1232 1332 1233
rect 1326 1228 1327 1232
rect 1331 1228 1332 1232
rect 1366 1232 1367 1236
rect 1371 1232 1372 1236
rect 1494 1233 1495 1237
rect 1499 1233 1500 1237
rect 1494 1232 1500 1233
rect 1366 1231 1372 1232
rect 1326 1227 1332 1228
rect 1366 1219 1372 1220
rect 1326 1215 1332 1216
rect 1326 1211 1327 1215
rect 1331 1211 1332 1215
rect 1366 1215 1367 1219
rect 1371 1215 1372 1219
rect 1366 1214 1372 1215
rect 1326 1210 1332 1211
rect 910 1206 916 1207
rect 910 1202 911 1206
rect 915 1202 916 1206
rect 910 1201 916 1202
rect 858 1199 864 1200
rect 858 1195 859 1199
rect 863 1195 864 1199
rect 858 1194 864 1195
rect 846 1191 852 1192
rect 511 1190 515 1191
rect 511 1185 515 1186
rect 535 1190 539 1191
rect 535 1185 539 1186
rect 599 1190 603 1191
rect 599 1185 603 1186
rect 615 1190 619 1191
rect 615 1185 619 1186
rect 687 1190 691 1191
rect 687 1185 691 1186
rect 759 1190 763 1191
rect 759 1185 763 1186
rect 767 1190 771 1191
rect 767 1185 771 1186
rect 831 1190 835 1191
rect 831 1185 835 1186
rect 839 1190 843 1191
rect 846 1187 847 1191
rect 851 1187 852 1191
rect 846 1186 852 1187
rect 839 1185 843 1186
rect 486 1183 492 1184
rect 486 1179 487 1183
rect 491 1179 492 1183
rect 512 1179 514 1185
rect 600 1179 602 1185
rect 678 1183 684 1184
rect 678 1179 679 1183
rect 683 1179 684 1183
rect 688 1179 690 1185
rect 706 1183 712 1184
rect 706 1179 707 1183
rect 711 1179 712 1183
rect 768 1179 770 1185
rect 786 1183 792 1184
rect 786 1179 787 1183
rect 791 1179 792 1183
rect 840 1179 842 1185
rect 354 1178 360 1179
rect 422 1178 428 1179
rect 486 1178 492 1179
rect 510 1178 516 1179
rect 310 1146 316 1147
rect 346 1147 352 1148
rect 258 1142 264 1143
rect 312 1127 314 1146
rect 346 1143 347 1147
rect 351 1143 352 1147
rect 346 1142 352 1143
rect 111 1126 115 1127
rect 111 1121 115 1122
rect 143 1126 147 1127
rect 143 1121 147 1122
rect 223 1126 227 1127
rect 223 1121 227 1122
rect 311 1126 315 1127
rect 311 1121 315 1122
rect 319 1126 323 1127
rect 319 1121 323 1122
rect 112 1109 114 1121
rect 224 1110 226 1121
rect 310 1111 316 1112
rect 222 1109 228 1110
rect 110 1108 116 1109
rect 110 1104 111 1108
rect 115 1104 116 1108
rect 222 1105 223 1109
rect 227 1105 228 1109
rect 310 1107 311 1111
rect 315 1107 316 1111
rect 320 1110 322 1121
rect 356 1112 358 1178
rect 422 1174 423 1178
rect 427 1174 428 1178
rect 422 1173 428 1174
rect 510 1174 511 1178
rect 515 1174 516 1178
rect 510 1173 516 1174
rect 598 1178 604 1179
rect 678 1178 684 1179
rect 686 1178 692 1179
rect 706 1178 712 1179
rect 766 1178 772 1179
rect 786 1178 792 1179
rect 838 1178 844 1179
rect 598 1174 599 1178
rect 603 1174 604 1178
rect 598 1173 604 1174
rect 406 1151 412 1152
rect 406 1147 407 1151
rect 411 1147 412 1151
rect 406 1146 412 1147
rect 494 1151 500 1152
rect 494 1147 495 1151
rect 499 1147 500 1151
rect 494 1146 500 1147
rect 582 1151 588 1152
rect 582 1147 583 1151
rect 587 1147 588 1151
rect 670 1151 676 1152
rect 582 1146 588 1147
rect 618 1147 624 1148
rect 408 1127 410 1146
rect 496 1127 498 1146
rect 584 1127 586 1146
rect 618 1143 619 1147
rect 623 1143 624 1147
rect 670 1147 671 1151
rect 675 1147 676 1151
rect 670 1146 676 1147
rect 618 1142 624 1143
rect 407 1126 411 1127
rect 407 1121 411 1122
rect 423 1126 427 1127
rect 423 1121 427 1122
rect 495 1126 499 1127
rect 495 1121 499 1122
rect 527 1126 531 1127
rect 527 1121 531 1122
rect 583 1126 587 1127
rect 583 1121 587 1122
rect 354 1111 360 1112
rect 310 1106 316 1107
rect 318 1109 324 1110
rect 222 1104 228 1105
rect 110 1103 116 1104
rect 110 1091 116 1092
rect 110 1087 111 1091
rect 115 1087 116 1091
rect 110 1086 116 1087
rect 112 1067 114 1086
rect 219 1084 223 1085
rect 219 1079 223 1080
rect 238 1082 244 1083
rect 220 1076 222 1079
rect 238 1078 239 1082
rect 243 1078 244 1082
rect 238 1077 244 1078
rect 218 1075 224 1076
rect 218 1071 219 1075
rect 223 1071 224 1075
rect 218 1070 224 1071
rect 240 1067 242 1077
rect 312 1076 314 1106
rect 318 1105 319 1109
rect 323 1105 324 1109
rect 354 1107 355 1111
rect 359 1107 360 1111
rect 424 1110 426 1121
rect 518 1111 524 1112
rect 354 1106 360 1107
rect 422 1109 428 1110
rect 318 1104 324 1105
rect 422 1105 423 1109
rect 427 1105 428 1109
rect 518 1107 519 1111
rect 523 1107 524 1111
rect 528 1110 530 1121
rect 550 1111 556 1112
rect 518 1106 524 1107
rect 526 1109 532 1110
rect 422 1104 428 1105
rect 334 1082 340 1083
rect 334 1078 335 1082
rect 339 1078 340 1082
rect 334 1077 340 1078
rect 438 1082 444 1083
rect 438 1078 439 1082
rect 443 1078 444 1082
rect 438 1077 444 1078
rect 310 1075 316 1076
rect 310 1071 311 1075
rect 315 1071 316 1075
rect 310 1070 316 1071
rect 336 1067 338 1077
rect 440 1067 442 1077
rect 520 1076 522 1106
rect 526 1105 527 1109
rect 531 1105 532 1109
rect 550 1107 551 1111
rect 555 1107 556 1111
rect 550 1106 556 1107
rect 526 1104 532 1105
rect 552 1085 554 1106
rect 551 1084 555 1085
rect 542 1082 548 1083
rect 542 1078 543 1082
rect 547 1078 548 1082
rect 551 1079 555 1080
rect 542 1077 548 1078
rect 454 1075 460 1076
rect 454 1071 455 1075
rect 459 1071 460 1075
rect 454 1070 460 1071
rect 518 1075 524 1076
rect 518 1071 519 1075
rect 523 1071 524 1075
rect 518 1070 524 1071
rect 111 1066 115 1067
rect 111 1061 115 1062
rect 239 1066 243 1067
rect 239 1061 243 1062
rect 311 1066 315 1067
rect 311 1061 315 1062
rect 335 1066 339 1067
rect 335 1061 339 1062
rect 367 1066 371 1067
rect 367 1061 371 1062
rect 439 1066 443 1067
rect 439 1061 443 1062
rect 112 1046 114 1061
rect 312 1055 314 1061
rect 368 1055 370 1061
rect 386 1059 392 1060
rect 386 1055 387 1059
rect 391 1055 392 1059
rect 440 1055 442 1061
rect 310 1054 316 1055
rect 310 1050 311 1054
rect 315 1050 316 1054
rect 310 1049 316 1050
rect 366 1054 372 1055
rect 386 1054 392 1055
rect 438 1054 444 1055
rect 366 1050 367 1054
rect 371 1050 372 1054
rect 366 1049 372 1050
rect 110 1045 116 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 110 1023 116 1024
rect 294 1027 300 1028
rect 294 1023 295 1027
rect 299 1023 300 1027
rect 112 1007 114 1023
rect 294 1022 300 1023
rect 350 1027 356 1028
rect 350 1023 351 1027
rect 355 1023 356 1027
rect 388 1024 390 1054
rect 438 1050 439 1054
rect 443 1050 444 1054
rect 438 1049 444 1050
rect 422 1027 428 1028
rect 350 1022 356 1023
rect 386 1023 392 1024
rect 296 1007 298 1022
rect 352 1007 354 1022
rect 386 1019 387 1023
rect 391 1019 392 1023
rect 422 1023 423 1027
rect 427 1023 428 1027
rect 456 1024 458 1070
rect 534 1067 540 1068
rect 544 1067 546 1077
rect 620 1076 622 1142
rect 672 1127 674 1146
rect 680 1140 682 1178
rect 686 1174 687 1178
rect 691 1174 692 1178
rect 686 1173 692 1174
rect 708 1148 710 1178
rect 766 1174 767 1178
rect 771 1174 772 1178
rect 766 1173 772 1174
rect 750 1151 756 1152
rect 706 1147 712 1148
rect 706 1143 707 1147
rect 711 1143 712 1147
rect 750 1147 751 1151
rect 755 1147 756 1151
rect 788 1148 790 1178
rect 838 1174 839 1178
rect 843 1174 844 1178
rect 838 1173 844 1174
rect 822 1151 828 1152
rect 750 1146 756 1147
rect 786 1147 792 1148
rect 706 1142 712 1143
rect 678 1139 684 1140
rect 678 1135 679 1139
rect 683 1135 684 1139
rect 678 1134 684 1135
rect 752 1127 754 1146
rect 786 1143 787 1147
rect 791 1143 792 1147
rect 822 1147 823 1151
rect 827 1147 828 1151
rect 860 1148 862 1194
rect 912 1191 914 1201
rect 1328 1191 1330 1210
rect 1368 1191 1370 1214
rect 1510 1210 1516 1211
rect 1510 1206 1511 1210
rect 1515 1206 1516 1210
rect 1510 1205 1516 1206
rect 1512 1191 1514 1205
rect 1520 1204 1522 1242
rect 1550 1239 1556 1240
rect 1550 1235 1551 1239
rect 1555 1235 1556 1239
rect 1560 1238 1562 1249
rect 1586 1239 1592 1240
rect 1550 1234 1556 1235
rect 1558 1237 1564 1238
rect 1552 1204 1554 1234
rect 1558 1233 1559 1237
rect 1563 1233 1564 1237
rect 1586 1235 1587 1239
rect 1591 1235 1592 1239
rect 1624 1238 1626 1249
rect 1586 1234 1592 1235
rect 1622 1237 1628 1238
rect 1558 1232 1564 1233
rect 1574 1210 1580 1211
rect 1574 1206 1575 1210
rect 1579 1206 1580 1210
rect 1574 1205 1580 1206
rect 1518 1203 1524 1204
rect 1518 1199 1519 1203
rect 1523 1199 1524 1203
rect 1518 1198 1524 1199
rect 1550 1203 1556 1204
rect 1550 1199 1551 1203
rect 1555 1199 1556 1203
rect 1550 1198 1556 1199
rect 1576 1191 1578 1205
rect 911 1190 915 1191
rect 911 1185 915 1186
rect 983 1190 987 1191
rect 983 1185 987 1186
rect 1063 1190 1067 1191
rect 1063 1185 1067 1186
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1415 1190 1419 1191
rect 1415 1185 1419 1186
rect 1503 1190 1507 1191
rect 1503 1185 1507 1186
rect 1511 1190 1515 1191
rect 1511 1185 1515 1186
rect 1575 1190 1579 1191
rect 1588 1188 1590 1234
rect 1622 1233 1623 1237
rect 1627 1233 1628 1237
rect 1622 1232 1628 1233
rect 1638 1210 1644 1211
rect 1638 1206 1639 1210
rect 1643 1206 1644 1210
rect 1638 1205 1644 1206
rect 1640 1191 1642 1205
rect 1664 1204 1666 1258
rect 1752 1255 1754 1266
rect 1687 1254 1691 1255
rect 1687 1249 1691 1250
rect 1751 1254 1755 1255
rect 1751 1249 1755 1250
rect 1759 1254 1763 1255
rect 1759 1249 1763 1250
rect 1688 1238 1690 1249
rect 1694 1247 1700 1248
rect 1694 1243 1695 1247
rect 1699 1243 1700 1247
rect 1694 1242 1700 1243
rect 1686 1237 1692 1238
rect 1686 1233 1687 1237
rect 1691 1233 1692 1237
rect 1686 1232 1692 1233
rect 1696 1204 1698 1242
rect 1750 1239 1756 1240
rect 1750 1235 1751 1239
rect 1755 1235 1756 1239
rect 1760 1238 1762 1249
rect 1792 1240 1794 1302
rect 1838 1299 1839 1303
rect 1843 1299 1844 1303
rect 1864 1299 1866 1305
rect 1960 1299 1962 1305
rect 1838 1298 1844 1299
rect 1862 1298 1868 1299
rect 1862 1294 1863 1298
rect 1867 1294 1868 1298
rect 1862 1293 1868 1294
rect 1958 1298 1964 1299
rect 1958 1294 1959 1298
rect 1963 1294 1964 1298
rect 1958 1293 1964 1294
rect 1846 1271 1852 1272
rect 1846 1267 1847 1271
rect 1851 1267 1852 1271
rect 1942 1271 1948 1272
rect 1846 1266 1852 1267
rect 1934 1267 1940 1268
rect 1848 1255 1850 1266
rect 1934 1263 1935 1267
rect 1939 1263 1940 1267
rect 1942 1267 1943 1271
rect 1947 1267 1948 1271
rect 1976 1268 1978 1314
rect 1984 1311 1986 1321
rect 2040 1320 2042 1350
rect 2046 1349 2047 1353
rect 2051 1349 2052 1353
rect 2118 1351 2119 1355
rect 2123 1351 2124 1355
rect 2128 1354 2130 1365
rect 2198 1355 2204 1356
rect 2118 1350 2124 1351
rect 2126 1353 2132 1354
rect 2046 1348 2052 1349
rect 2062 1326 2068 1327
rect 2062 1322 2063 1326
rect 2067 1322 2068 1326
rect 2062 1321 2068 1322
rect 2038 1319 2044 1320
rect 2038 1315 2039 1319
rect 2043 1315 2044 1319
rect 2038 1314 2044 1315
rect 2054 1311 2060 1312
rect 2064 1311 2066 1321
rect 2120 1320 2122 1350
rect 2126 1349 2127 1353
rect 2131 1349 2132 1353
rect 2198 1351 2199 1355
rect 2203 1351 2204 1355
rect 2208 1354 2210 1365
rect 2240 1356 2242 1426
rect 2282 1423 2283 1427
rect 2287 1423 2288 1427
rect 2304 1423 2306 1429
rect 2392 1423 2394 1429
rect 2480 1423 2482 1429
rect 2506 1427 2512 1428
rect 2506 1423 2507 1427
rect 2511 1423 2512 1427
rect 2544 1423 2546 1429
rect 2282 1422 2288 1423
rect 2302 1422 2308 1423
rect 2302 1418 2303 1422
rect 2307 1418 2308 1422
rect 2302 1417 2308 1418
rect 2390 1422 2396 1423
rect 2390 1418 2391 1422
rect 2395 1418 2396 1422
rect 2390 1417 2396 1418
rect 2478 1422 2484 1423
rect 2506 1422 2512 1423
rect 2542 1422 2548 1423
rect 2478 1418 2479 1422
rect 2483 1418 2484 1422
rect 2478 1417 2484 1418
rect 2286 1395 2292 1396
rect 2286 1391 2287 1395
rect 2291 1391 2292 1395
rect 2286 1390 2292 1391
rect 2374 1395 2380 1396
rect 2374 1391 2375 1395
rect 2379 1391 2380 1395
rect 2374 1390 2380 1391
rect 2462 1395 2468 1396
rect 2462 1391 2463 1395
rect 2467 1391 2468 1395
rect 2508 1392 2510 1422
rect 2542 1418 2543 1422
rect 2547 1418 2548 1422
rect 2542 1417 2548 1418
rect 2526 1395 2532 1396
rect 2462 1390 2468 1391
rect 2506 1391 2512 1392
rect 2288 1371 2290 1390
rect 2376 1371 2378 1390
rect 2464 1371 2466 1390
rect 2506 1387 2507 1391
rect 2511 1387 2512 1391
rect 2526 1391 2527 1395
rect 2531 1391 2532 1395
rect 2560 1392 2562 1434
rect 2583 1429 2587 1430
rect 2584 1414 2586 1429
rect 2582 1413 2588 1414
rect 2582 1409 2583 1413
rect 2587 1409 2588 1413
rect 2582 1408 2588 1409
rect 2582 1396 2588 1397
rect 2582 1392 2583 1396
rect 2587 1392 2588 1396
rect 2526 1390 2532 1391
rect 2558 1391 2564 1392
rect 2582 1391 2588 1392
rect 2506 1386 2512 1387
rect 2528 1371 2530 1390
rect 2558 1387 2559 1391
rect 2563 1387 2564 1391
rect 2558 1386 2564 1387
rect 2584 1371 2586 1391
rect 2287 1370 2291 1371
rect 2287 1365 2291 1366
rect 2375 1370 2379 1371
rect 2375 1365 2379 1366
rect 2463 1370 2467 1371
rect 2463 1365 2467 1366
rect 2527 1370 2531 1371
rect 2527 1365 2531 1366
rect 2583 1370 2587 1371
rect 2583 1365 2587 1366
rect 2238 1355 2244 1356
rect 2198 1350 2204 1351
rect 2206 1353 2212 1354
rect 2126 1348 2132 1349
rect 2142 1326 2148 1327
rect 2142 1322 2143 1326
rect 2147 1322 2148 1326
rect 2142 1321 2148 1322
rect 2118 1319 2124 1320
rect 2118 1315 2119 1319
rect 2123 1315 2124 1319
rect 2118 1314 2124 1315
rect 2144 1311 2146 1321
rect 2200 1320 2202 1350
rect 2206 1349 2207 1353
rect 2211 1349 2212 1353
rect 2238 1351 2239 1355
rect 2243 1351 2244 1355
rect 2584 1353 2586 1365
rect 2238 1350 2244 1351
rect 2582 1352 2588 1353
rect 2206 1348 2212 1349
rect 2582 1348 2583 1352
rect 2587 1348 2588 1352
rect 2582 1347 2588 1348
rect 2582 1335 2588 1336
rect 2582 1331 2583 1335
rect 2587 1331 2588 1335
rect 2582 1330 2588 1331
rect 2222 1326 2228 1327
rect 2222 1322 2223 1326
rect 2227 1322 2228 1326
rect 2222 1321 2228 1322
rect 2198 1319 2204 1320
rect 2198 1315 2199 1319
rect 2203 1315 2204 1319
rect 2198 1314 2204 1315
rect 2224 1311 2226 1321
rect 2246 1311 2252 1312
rect 2584 1311 2586 1330
rect 1983 1310 1987 1311
rect 1983 1305 1987 1306
rect 2047 1310 2051 1311
rect 2054 1307 2055 1311
rect 2059 1307 2060 1311
rect 2054 1306 2060 1307
rect 2063 1310 2067 1311
rect 2047 1305 2051 1306
rect 2022 1303 2028 1304
rect 2022 1299 2023 1303
rect 2027 1299 2028 1303
rect 2048 1299 2050 1305
rect 2022 1298 2028 1299
rect 2046 1298 2052 1299
rect 2024 1280 2026 1298
rect 2046 1294 2047 1298
rect 2051 1294 2052 1298
rect 2046 1293 2052 1294
rect 2022 1279 2028 1280
rect 2022 1275 2023 1279
rect 2027 1275 2028 1279
rect 2022 1274 2028 1275
rect 2030 1271 2036 1272
rect 1942 1266 1948 1267
rect 1974 1267 1980 1268
rect 1934 1262 1940 1263
rect 1823 1254 1827 1255
rect 1823 1249 1827 1250
rect 1847 1254 1851 1255
rect 1847 1249 1851 1250
rect 1887 1254 1891 1255
rect 1887 1249 1891 1250
rect 1790 1239 1796 1240
rect 1750 1234 1756 1235
rect 1758 1237 1764 1238
rect 1702 1210 1708 1211
rect 1702 1206 1703 1210
rect 1707 1206 1708 1210
rect 1702 1205 1708 1206
rect 1662 1203 1668 1204
rect 1662 1199 1663 1203
rect 1667 1199 1668 1203
rect 1662 1198 1668 1199
rect 1694 1203 1700 1204
rect 1694 1199 1695 1203
rect 1699 1199 1700 1203
rect 1694 1198 1700 1199
rect 1704 1191 1706 1205
rect 1752 1204 1754 1234
rect 1758 1233 1759 1237
rect 1763 1233 1764 1237
rect 1790 1235 1791 1239
rect 1795 1235 1796 1239
rect 1824 1238 1826 1249
rect 1888 1238 1890 1249
rect 1790 1234 1796 1235
rect 1822 1237 1828 1238
rect 1758 1232 1764 1233
rect 1822 1233 1823 1237
rect 1827 1233 1828 1237
rect 1822 1232 1828 1233
rect 1886 1237 1892 1238
rect 1886 1233 1887 1237
rect 1891 1233 1892 1237
rect 1886 1232 1892 1233
rect 1774 1210 1780 1211
rect 1774 1206 1775 1210
rect 1779 1206 1780 1210
rect 1774 1205 1780 1206
rect 1838 1210 1844 1211
rect 1838 1206 1839 1210
rect 1843 1206 1844 1210
rect 1838 1205 1844 1206
rect 1902 1210 1908 1211
rect 1902 1206 1903 1210
rect 1907 1206 1908 1210
rect 1902 1205 1908 1206
rect 1750 1203 1756 1204
rect 1750 1199 1751 1203
rect 1755 1199 1756 1203
rect 1750 1198 1756 1199
rect 1776 1191 1778 1205
rect 1840 1191 1842 1205
rect 1904 1191 1906 1205
rect 1936 1204 1938 1262
rect 1944 1255 1946 1266
rect 1974 1263 1975 1267
rect 1979 1263 1980 1267
rect 2030 1267 2031 1271
rect 2035 1267 2036 1271
rect 2056 1268 2058 1306
rect 2063 1305 2067 1306
rect 2135 1310 2139 1311
rect 2135 1305 2139 1306
rect 2143 1310 2147 1311
rect 2143 1305 2147 1306
rect 2223 1310 2227 1311
rect 2223 1305 2227 1306
rect 2231 1310 2235 1311
rect 2246 1307 2247 1311
rect 2251 1307 2252 1311
rect 2246 1306 2252 1307
rect 2583 1310 2587 1311
rect 2231 1305 2235 1306
rect 2136 1299 2138 1305
rect 2186 1303 2192 1304
rect 2186 1299 2187 1303
rect 2191 1299 2192 1303
rect 2232 1299 2234 1305
rect 2134 1298 2140 1299
rect 2186 1298 2192 1299
rect 2230 1298 2236 1299
rect 2134 1294 2135 1298
rect 2139 1294 2140 1298
rect 2134 1293 2140 1294
rect 2118 1271 2124 1272
rect 2030 1266 2036 1267
rect 2054 1267 2060 1268
rect 1974 1262 1980 1263
rect 2032 1255 2034 1266
rect 2054 1263 2055 1267
rect 2059 1263 2060 1267
rect 2118 1267 2119 1271
rect 2123 1267 2124 1271
rect 2118 1266 2124 1267
rect 2054 1262 2060 1263
rect 2120 1255 2122 1266
rect 1943 1254 1947 1255
rect 1943 1249 1947 1250
rect 1951 1254 1955 1255
rect 1951 1249 1955 1250
rect 2015 1254 2019 1255
rect 2015 1249 2019 1250
rect 2031 1254 2035 1255
rect 2031 1249 2035 1250
rect 2079 1254 2083 1255
rect 2079 1249 2083 1250
rect 2119 1254 2123 1255
rect 2119 1249 2123 1250
rect 2151 1254 2155 1255
rect 2151 1249 2155 1250
rect 1952 1238 1954 1249
rect 2006 1239 2012 1240
rect 1950 1237 1956 1238
rect 1950 1233 1951 1237
rect 1955 1233 1956 1237
rect 2006 1235 2007 1239
rect 2011 1235 2012 1239
rect 2016 1238 2018 1249
rect 2038 1239 2044 1240
rect 2006 1234 2012 1235
rect 2014 1237 2020 1238
rect 1950 1232 1956 1233
rect 1966 1210 1972 1211
rect 1966 1206 1967 1210
rect 1971 1206 1972 1210
rect 1966 1205 1972 1206
rect 1926 1203 1932 1204
rect 1926 1199 1927 1203
rect 1931 1199 1932 1203
rect 1926 1198 1932 1199
rect 1934 1203 1940 1204
rect 1934 1199 1935 1203
rect 1939 1199 1940 1203
rect 1934 1198 1940 1199
rect 1599 1190 1603 1191
rect 1575 1185 1579 1186
rect 1586 1187 1592 1188
rect 886 1183 892 1184
rect 886 1179 887 1183
rect 891 1179 892 1183
rect 912 1179 914 1185
rect 984 1179 986 1185
rect 1002 1183 1008 1184
rect 1002 1179 1003 1183
rect 1007 1179 1008 1183
rect 1064 1179 1066 1185
rect 886 1178 892 1179
rect 910 1178 916 1179
rect 888 1160 890 1178
rect 910 1174 911 1178
rect 915 1174 916 1178
rect 910 1173 916 1174
rect 982 1178 988 1179
rect 1002 1178 1008 1179
rect 1062 1178 1068 1179
rect 982 1174 983 1178
rect 987 1174 988 1178
rect 982 1173 988 1174
rect 886 1159 892 1160
rect 886 1155 887 1159
rect 891 1155 892 1159
rect 886 1154 892 1155
rect 894 1151 900 1152
rect 822 1146 828 1147
rect 858 1147 864 1148
rect 786 1142 792 1143
rect 824 1127 826 1146
rect 858 1143 859 1147
rect 863 1143 864 1147
rect 894 1147 895 1151
rect 899 1147 900 1151
rect 894 1146 900 1147
rect 966 1151 972 1152
rect 966 1147 967 1151
rect 971 1147 972 1151
rect 1004 1148 1006 1178
rect 1062 1174 1063 1178
rect 1067 1174 1068 1178
rect 1062 1173 1068 1174
rect 1328 1170 1330 1185
rect 1368 1170 1370 1185
rect 1390 1183 1396 1184
rect 1390 1179 1391 1183
rect 1395 1179 1396 1183
rect 1416 1179 1418 1185
rect 1494 1183 1500 1184
rect 1494 1179 1495 1183
rect 1499 1179 1500 1183
rect 1504 1179 1506 1185
rect 1586 1183 1587 1187
rect 1591 1183 1592 1187
rect 1599 1185 1603 1186
rect 1639 1190 1643 1191
rect 1639 1185 1643 1186
rect 1703 1190 1707 1191
rect 1703 1185 1707 1186
rect 1775 1190 1779 1191
rect 1775 1185 1779 1186
rect 1807 1190 1811 1191
rect 1807 1185 1811 1186
rect 1839 1190 1843 1191
rect 1839 1185 1843 1186
rect 1903 1190 1907 1191
rect 1903 1185 1907 1186
rect 1911 1190 1915 1191
rect 1911 1185 1915 1186
rect 1586 1182 1592 1183
rect 1600 1179 1602 1185
rect 1618 1183 1624 1184
rect 1618 1179 1619 1183
rect 1623 1179 1624 1183
rect 1704 1179 1706 1185
rect 1722 1183 1728 1184
rect 1722 1179 1723 1183
rect 1727 1179 1728 1183
rect 1808 1179 1810 1185
rect 1826 1183 1832 1184
rect 1826 1179 1827 1183
rect 1831 1179 1832 1183
rect 1912 1179 1914 1185
rect 1390 1178 1396 1179
rect 1414 1178 1420 1179
rect 1494 1178 1500 1179
rect 1502 1178 1508 1179
rect 1326 1169 1332 1170
rect 1326 1165 1327 1169
rect 1331 1165 1332 1169
rect 1326 1164 1332 1165
rect 1366 1169 1372 1170
rect 1366 1165 1367 1169
rect 1371 1165 1372 1169
rect 1366 1164 1372 1165
rect 1392 1160 1394 1178
rect 1414 1174 1415 1178
rect 1419 1174 1420 1178
rect 1414 1173 1420 1174
rect 1390 1159 1396 1160
rect 1390 1155 1391 1159
rect 1395 1155 1396 1159
rect 1390 1154 1396 1155
rect 1326 1152 1332 1153
rect 1046 1151 1052 1152
rect 966 1146 972 1147
rect 1002 1147 1008 1148
rect 858 1142 864 1143
rect 896 1127 898 1146
rect 968 1127 970 1146
rect 1002 1143 1003 1147
rect 1007 1143 1008 1147
rect 1046 1147 1047 1151
rect 1051 1147 1052 1151
rect 1326 1148 1327 1152
rect 1331 1148 1332 1152
rect 1326 1147 1332 1148
rect 1366 1152 1372 1153
rect 1366 1148 1367 1152
rect 1371 1148 1372 1152
rect 1366 1147 1372 1148
rect 1398 1151 1404 1152
rect 1398 1147 1399 1151
rect 1403 1147 1404 1151
rect 1486 1151 1492 1152
rect 1046 1146 1052 1147
rect 1002 1142 1008 1143
rect 1048 1127 1050 1146
rect 1328 1127 1330 1147
rect 1368 1131 1370 1147
rect 1398 1146 1404 1147
rect 1422 1147 1428 1148
rect 1400 1131 1402 1146
rect 1422 1143 1423 1147
rect 1427 1143 1428 1147
rect 1486 1147 1487 1151
rect 1491 1147 1492 1151
rect 1486 1146 1492 1147
rect 1422 1142 1428 1143
rect 1367 1130 1371 1131
rect 631 1126 635 1127
rect 631 1121 635 1122
rect 671 1126 675 1127
rect 671 1121 675 1122
rect 727 1126 731 1127
rect 727 1121 731 1122
rect 751 1126 755 1127
rect 751 1121 755 1122
rect 823 1126 827 1127
rect 823 1121 827 1122
rect 895 1126 899 1127
rect 895 1121 899 1122
rect 911 1126 915 1127
rect 911 1121 915 1122
rect 967 1126 971 1127
rect 967 1121 971 1122
rect 991 1126 995 1127
rect 991 1121 995 1122
rect 1047 1126 1051 1127
rect 1047 1121 1051 1122
rect 1079 1126 1083 1127
rect 1079 1121 1083 1122
rect 1167 1126 1171 1127
rect 1167 1121 1171 1122
rect 1327 1126 1331 1127
rect 1367 1125 1371 1126
rect 1399 1130 1403 1131
rect 1399 1125 1403 1126
rect 1327 1121 1331 1122
rect 632 1110 634 1121
rect 678 1111 684 1112
rect 630 1109 636 1110
rect 630 1105 631 1109
rect 635 1105 636 1109
rect 678 1107 679 1111
rect 683 1107 684 1111
rect 728 1110 730 1121
rect 814 1111 820 1112
rect 678 1106 684 1107
rect 726 1109 732 1110
rect 630 1104 636 1105
rect 646 1082 652 1083
rect 646 1078 647 1082
rect 651 1078 652 1082
rect 646 1077 652 1078
rect 618 1075 624 1076
rect 618 1071 619 1075
rect 623 1071 624 1075
rect 618 1070 624 1071
rect 648 1067 650 1077
rect 519 1066 523 1067
rect 534 1063 535 1067
rect 539 1063 540 1067
rect 534 1062 540 1063
rect 543 1066 547 1067
rect 519 1061 523 1062
rect 494 1059 500 1060
rect 494 1055 495 1059
rect 499 1055 500 1059
rect 520 1055 522 1061
rect 494 1054 500 1055
rect 518 1054 524 1055
rect 496 1036 498 1054
rect 518 1050 519 1054
rect 523 1050 524 1054
rect 518 1049 524 1050
rect 494 1035 500 1036
rect 494 1031 495 1035
rect 499 1031 500 1035
rect 494 1030 500 1031
rect 502 1027 508 1028
rect 422 1022 428 1023
rect 454 1023 460 1024
rect 386 1018 392 1019
rect 424 1007 426 1022
rect 454 1019 455 1023
rect 459 1019 460 1023
rect 502 1023 503 1027
rect 507 1023 508 1027
rect 536 1024 538 1062
rect 543 1061 547 1062
rect 607 1066 611 1067
rect 607 1061 611 1062
rect 647 1066 651 1067
rect 647 1061 651 1062
rect 562 1059 568 1060
rect 562 1055 563 1059
rect 567 1055 568 1059
rect 608 1055 610 1061
rect 680 1060 682 1106
rect 726 1105 727 1109
rect 731 1105 732 1109
rect 814 1107 815 1111
rect 819 1107 820 1111
rect 824 1110 826 1121
rect 902 1111 908 1112
rect 814 1106 820 1107
rect 822 1109 828 1110
rect 726 1104 732 1105
rect 742 1082 748 1083
rect 742 1078 743 1082
rect 747 1078 748 1082
rect 742 1077 748 1078
rect 744 1067 746 1077
rect 816 1076 818 1106
rect 822 1105 823 1109
rect 827 1105 828 1109
rect 902 1107 903 1111
rect 907 1107 908 1111
rect 912 1110 914 1121
rect 992 1110 994 1121
rect 1014 1119 1020 1120
rect 1014 1115 1015 1119
rect 1019 1115 1020 1119
rect 1014 1114 1020 1115
rect 902 1106 908 1107
rect 910 1109 916 1110
rect 822 1104 828 1105
rect 838 1082 844 1083
rect 838 1078 839 1082
rect 843 1078 844 1082
rect 838 1077 844 1078
rect 814 1075 820 1076
rect 814 1071 815 1075
rect 819 1071 820 1075
rect 814 1070 820 1071
rect 840 1067 842 1077
rect 904 1076 906 1106
rect 910 1105 911 1109
rect 915 1105 916 1109
rect 910 1104 916 1105
rect 990 1109 996 1110
rect 990 1105 991 1109
rect 995 1105 996 1109
rect 990 1104 996 1105
rect 926 1082 932 1083
rect 926 1078 927 1082
rect 931 1078 932 1082
rect 926 1077 932 1078
rect 1006 1082 1012 1083
rect 1006 1078 1007 1082
rect 1011 1078 1012 1082
rect 1006 1077 1012 1078
rect 902 1075 908 1076
rect 902 1071 903 1075
rect 907 1071 908 1075
rect 902 1070 908 1071
rect 928 1067 930 1077
rect 1008 1067 1010 1077
rect 1016 1076 1018 1114
rect 1022 1111 1028 1112
rect 1022 1107 1023 1111
rect 1027 1107 1028 1111
rect 1080 1110 1082 1121
rect 1158 1111 1164 1112
rect 1022 1106 1028 1107
rect 1078 1109 1084 1110
rect 1014 1075 1020 1076
rect 1014 1071 1015 1075
rect 1019 1071 1020 1075
rect 1014 1070 1020 1071
rect 1024 1068 1026 1106
rect 1078 1105 1079 1109
rect 1083 1105 1084 1109
rect 1158 1107 1159 1111
rect 1163 1107 1164 1111
rect 1168 1110 1170 1121
rect 1158 1106 1164 1107
rect 1166 1109 1172 1110
rect 1328 1109 1330 1121
rect 1368 1113 1370 1125
rect 1400 1114 1402 1125
rect 1398 1113 1404 1114
rect 1366 1112 1372 1113
rect 1078 1104 1084 1105
rect 1094 1082 1100 1083
rect 1094 1078 1095 1082
rect 1099 1078 1100 1082
rect 1094 1077 1100 1078
rect 1070 1075 1076 1076
rect 1070 1071 1071 1075
rect 1075 1071 1076 1075
rect 1070 1070 1076 1071
rect 1022 1067 1028 1068
rect 703 1066 707 1067
rect 703 1061 707 1062
rect 743 1066 747 1067
rect 743 1061 747 1062
rect 799 1066 803 1067
rect 799 1061 803 1062
rect 839 1066 843 1067
rect 839 1061 843 1062
rect 887 1066 891 1067
rect 887 1061 891 1062
rect 927 1066 931 1067
rect 927 1061 931 1062
rect 975 1066 979 1067
rect 975 1061 979 1062
rect 1007 1066 1011 1067
rect 1022 1063 1023 1067
rect 1027 1063 1028 1067
rect 1022 1062 1028 1063
rect 1055 1066 1059 1067
rect 1007 1061 1011 1062
rect 1055 1061 1059 1062
rect 678 1059 684 1060
rect 678 1055 679 1059
rect 683 1055 684 1059
rect 704 1055 706 1061
rect 722 1059 728 1060
rect 722 1055 723 1059
rect 727 1055 728 1059
rect 800 1055 802 1061
rect 878 1059 884 1060
rect 878 1055 879 1059
rect 883 1055 884 1059
rect 888 1055 890 1061
rect 906 1059 912 1060
rect 906 1055 907 1059
rect 911 1055 912 1059
rect 976 1055 978 1061
rect 994 1059 1000 1060
rect 994 1055 995 1059
rect 999 1055 1000 1059
rect 1056 1055 1058 1061
rect 1062 1059 1068 1060
rect 1062 1055 1063 1059
rect 1067 1055 1068 1059
rect 562 1054 568 1055
rect 606 1054 612 1055
rect 678 1054 684 1055
rect 702 1054 708 1055
rect 722 1054 728 1055
rect 798 1054 804 1055
rect 878 1054 884 1055
rect 886 1054 892 1055
rect 906 1054 912 1055
rect 974 1054 980 1055
rect 994 1054 1000 1055
rect 1054 1054 1060 1055
rect 1062 1054 1068 1055
rect 502 1022 508 1023
rect 534 1023 540 1024
rect 454 1018 460 1019
rect 504 1007 506 1022
rect 534 1019 535 1023
rect 539 1019 540 1023
rect 534 1018 540 1019
rect 111 1006 115 1007
rect 111 1001 115 1002
rect 295 1006 299 1007
rect 295 1001 299 1002
rect 351 1006 355 1007
rect 351 1001 355 1002
rect 415 1006 419 1007
rect 415 1001 419 1002
rect 423 1006 427 1007
rect 423 1001 427 1002
rect 471 1006 475 1007
rect 471 1001 475 1002
rect 503 1006 507 1007
rect 503 1001 507 1002
rect 527 1006 531 1007
rect 527 1001 531 1002
rect 112 989 114 1001
rect 416 990 418 1001
rect 438 999 444 1000
rect 438 995 439 999
rect 443 995 444 999
rect 438 994 444 995
rect 414 989 420 990
rect 110 988 116 989
rect 110 984 111 988
rect 115 984 116 988
rect 414 985 415 989
rect 419 985 420 989
rect 414 984 420 985
rect 110 983 116 984
rect 110 971 116 972
rect 110 967 111 971
rect 115 967 116 971
rect 110 966 116 967
rect 112 947 114 966
rect 430 962 436 963
rect 430 958 431 962
rect 435 958 436 962
rect 430 957 436 958
rect 432 947 434 957
rect 440 956 442 994
rect 462 991 468 992
rect 462 987 463 991
rect 467 987 468 991
rect 472 990 474 1001
rect 518 991 524 992
rect 462 986 468 987
rect 470 989 476 990
rect 464 956 466 986
rect 470 985 471 989
rect 475 985 476 989
rect 518 987 519 991
rect 523 987 524 991
rect 528 990 530 1001
rect 564 992 566 1054
rect 606 1050 607 1054
rect 611 1050 612 1054
rect 606 1049 612 1050
rect 702 1050 703 1054
rect 707 1050 708 1054
rect 702 1049 708 1050
rect 590 1027 596 1028
rect 590 1023 591 1027
rect 595 1023 596 1027
rect 590 1022 596 1023
rect 686 1027 692 1028
rect 686 1023 687 1027
rect 691 1023 692 1027
rect 724 1024 726 1054
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 880 1029 882 1054
rect 886 1050 887 1054
rect 891 1050 892 1054
rect 886 1049 892 1050
rect 879 1028 883 1029
rect 782 1027 788 1028
rect 686 1022 692 1023
rect 722 1023 728 1024
rect 592 1007 594 1022
rect 688 1007 690 1022
rect 722 1019 723 1023
rect 727 1019 728 1023
rect 782 1023 783 1027
rect 787 1023 788 1027
rect 782 1022 788 1023
rect 870 1027 876 1028
rect 870 1023 871 1027
rect 875 1023 876 1027
rect 908 1024 910 1054
rect 974 1050 975 1054
rect 979 1050 980 1054
rect 974 1049 980 1050
rect 958 1027 964 1028
rect 879 1023 883 1024
rect 906 1023 912 1024
rect 870 1022 876 1023
rect 722 1018 728 1019
rect 754 1019 760 1020
rect 754 1015 755 1019
rect 759 1015 760 1019
rect 754 1014 760 1015
rect 591 1006 595 1007
rect 591 1001 595 1002
rect 655 1006 659 1007
rect 655 1001 659 1002
rect 687 1006 691 1007
rect 687 1001 691 1002
rect 719 1006 723 1007
rect 719 1001 723 1002
rect 562 991 568 992
rect 518 986 524 987
rect 526 989 532 990
rect 470 984 476 985
rect 486 962 492 963
rect 486 958 487 962
rect 491 958 492 962
rect 486 957 492 958
rect 438 955 444 956
rect 438 951 439 955
rect 443 951 444 955
rect 438 950 444 951
rect 462 955 468 956
rect 462 951 463 955
rect 467 951 468 955
rect 462 950 468 951
rect 488 947 490 957
rect 520 956 522 986
rect 526 985 527 989
rect 531 985 532 989
rect 562 987 563 991
rect 567 987 568 991
rect 592 990 594 1001
rect 638 995 644 996
rect 638 991 639 995
rect 643 991 644 995
rect 638 990 644 991
rect 656 990 658 1001
rect 720 990 722 1001
rect 746 991 752 992
rect 562 986 568 987
rect 590 989 596 990
rect 526 984 532 985
rect 590 985 591 989
rect 595 985 596 989
rect 590 984 596 985
rect 542 962 548 963
rect 542 958 543 962
rect 547 958 548 962
rect 542 957 548 958
rect 606 962 612 963
rect 606 958 607 962
rect 611 958 612 962
rect 606 957 612 958
rect 518 955 524 956
rect 518 951 519 955
rect 523 951 524 955
rect 518 950 524 951
rect 544 947 546 957
rect 608 947 610 957
rect 640 956 642 990
rect 654 989 660 990
rect 654 985 655 989
rect 659 985 660 989
rect 654 984 660 985
rect 718 989 724 990
rect 718 985 719 989
rect 723 985 724 989
rect 746 987 747 991
rect 751 987 752 991
rect 746 986 752 987
rect 718 984 724 985
rect 670 962 676 963
rect 670 958 671 962
rect 675 958 676 962
rect 670 957 676 958
rect 734 962 740 963
rect 734 958 735 962
rect 739 958 740 962
rect 734 957 740 958
rect 638 955 644 956
rect 638 951 639 955
rect 643 951 644 955
rect 638 950 644 951
rect 662 955 668 956
rect 662 951 663 955
rect 667 951 668 955
rect 662 950 668 951
rect 111 946 115 947
rect 111 941 115 942
rect 423 946 427 947
rect 423 941 427 942
rect 431 946 435 947
rect 431 941 435 942
rect 479 946 483 947
rect 479 941 483 942
rect 487 946 491 947
rect 487 941 491 942
rect 535 946 539 947
rect 535 941 539 942
rect 543 946 547 947
rect 543 941 547 942
rect 591 946 595 947
rect 591 941 595 942
rect 607 946 611 947
rect 607 941 611 942
rect 647 946 651 947
rect 647 941 651 942
rect 112 926 114 941
rect 414 939 420 940
rect 414 935 415 939
rect 419 935 420 939
rect 424 935 426 941
rect 442 939 448 940
rect 442 935 443 939
rect 447 935 448 939
rect 480 935 482 941
rect 498 939 504 940
rect 498 935 499 939
rect 503 935 504 939
rect 536 935 538 941
rect 554 939 560 940
rect 554 935 555 939
rect 559 935 560 939
rect 592 935 594 941
rect 648 935 650 941
rect 414 934 420 935
rect 422 934 428 935
rect 442 934 448 935
rect 478 934 484 935
rect 498 934 504 935
rect 534 934 540 935
rect 554 934 560 935
rect 590 934 596 935
rect 110 925 116 926
rect 110 921 111 925
rect 115 921 116 925
rect 110 920 116 921
rect 110 908 116 909
rect 110 904 111 908
rect 115 904 116 908
rect 110 903 116 904
rect 406 907 412 908
rect 406 903 407 907
rect 411 903 412 907
rect 112 891 114 903
rect 406 902 412 903
rect 408 891 410 902
rect 111 890 115 891
rect 111 885 115 886
rect 279 890 283 891
rect 279 885 283 886
rect 335 890 339 891
rect 335 885 339 886
rect 391 890 395 891
rect 391 885 395 886
rect 407 890 411 891
rect 407 885 411 886
rect 112 873 114 885
rect 280 874 282 885
rect 326 875 332 876
rect 278 873 284 874
rect 110 872 116 873
rect 110 868 111 872
rect 115 868 116 872
rect 278 869 279 873
rect 283 869 284 873
rect 326 871 327 875
rect 331 871 332 875
rect 336 874 338 885
rect 382 875 388 876
rect 326 870 332 871
rect 334 873 340 874
rect 278 868 284 869
rect 110 867 116 868
rect 110 855 116 856
rect 110 851 111 855
rect 115 851 116 855
rect 110 850 116 851
rect 112 827 114 850
rect 294 846 300 847
rect 294 842 295 846
rect 299 842 300 846
rect 294 841 300 842
rect 296 827 298 841
rect 328 840 330 870
rect 334 869 335 873
rect 339 869 340 873
rect 382 871 383 875
rect 387 871 388 875
rect 392 874 394 885
rect 416 884 418 934
rect 422 930 423 934
rect 427 930 428 934
rect 422 929 428 930
rect 444 904 446 934
rect 478 930 479 934
rect 483 930 484 934
rect 478 929 484 930
rect 462 907 468 908
rect 442 903 448 904
rect 442 899 443 903
rect 447 899 448 903
rect 462 903 463 907
rect 467 903 468 907
rect 500 904 502 934
rect 534 930 535 934
rect 539 930 540 934
rect 534 929 540 930
rect 518 907 524 908
rect 462 902 468 903
rect 498 903 504 904
rect 442 898 448 899
rect 464 891 466 902
rect 498 899 499 903
rect 503 899 504 903
rect 518 903 519 907
rect 523 903 524 907
rect 556 904 558 934
rect 590 930 591 934
rect 595 930 596 934
rect 590 929 596 930
rect 646 934 652 935
rect 646 930 647 934
rect 651 930 652 934
rect 646 929 652 930
rect 574 907 580 908
rect 518 902 524 903
rect 554 903 560 904
rect 498 898 504 899
rect 520 891 522 902
rect 554 899 555 903
rect 559 899 560 903
rect 574 903 575 907
rect 579 903 580 907
rect 574 902 580 903
rect 630 907 636 908
rect 630 903 631 907
rect 635 903 636 907
rect 664 904 666 950
rect 672 947 674 957
rect 736 947 738 957
rect 671 946 675 947
rect 671 941 675 942
rect 703 946 707 947
rect 703 941 707 942
rect 735 946 739 947
rect 748 944 750 986
rect 756 956 758 1014
rect 784 1007 786 1022
rect 872 1007 874 1022
rect 906 1019 907 1023
rect 911 1019 912 1023
rect 958 1023 959 1027
rect 963 1023 964 1027
rect 996 1024 998 1054
rect 1054 1050 1055 1054
rect 1059 1050 1060 1054
rect 1054 1049 1060 1050
rect 1038 1027 1044 1028
rect 958 1022 964 1023
rect 994 1023 1000 1024
rect 906 1018 912 1019
rect 946 1011 952 1012
rect 946 1007 947 1011
rect 951 1007 952 1011
rect 960 1007 962 1022
rect 994 1019 995 1023
rect 999 1019 1000 1023
rect 1038 1023 1039 1027
rect 1043 1023 1044 1027
rect 1038 1022 1044 1023
rect 994 1018 1000 1019
rect 1040 1007 1042 1022
rect 1064 1012 1066 1054
rect 1072 1024 1074 1070
rect 1096 1067 1098 1077
rect 1160 1076 1162 1106
rect 1166 1105 1167 1109
rect 1171 1105 1172 1109
rect 1166 1104 1172 1105
rect 1326 1108 1332 1109
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1366 1108 1367 1112
rect 1371 1108 1372 1112
rect 1398 1109 1399 1113
rect 1403 1109 1404 1113
rect 1398 1108 1404 1109
rect 1366 1107 1372 1108
rect 1326 1103 1332 1104
rect 1366 1095 1372 1096
rect 1326 1091 1332 1092
rect 1326 1087 1327 1091
rect 1331 1087 1332 1091
rect 1366 1091 1367 1095
rect 1371 1091 1372 1095
rect 1366 1090 1372 1091
rect 1326 1086 1332 1087
rect 1182 1082 1188 1083
rect 1182 1078 1183 1082
rect 1187 1078 1188 1082
rect 1182 1077 1188 1078
rect 1158 1075 1164 1076
rect 1158 1071 1159 1075
rect 1163 1071 1164 1075
rect 1158 1070 1164 1071
rect 1184 1067 1186 1077
rect 1328 1067 1330 1086
rect 1368 1071 1370 1090
rect 1414 1086 1420 1087
rect 1414 1082 1415 1086
rect 1419 1082 1420 1086
rect 1414 1081 1420 1082
rect 1416 1071 1418 1081
rect 1424 1080 1426 1142
rect 1488 1131 1490 1146
rect 1496 1140 1498 1178
rect 1502 1174 1503 1178
rect 1507 1174 1508 1178
rect 1502 1173 1508 1174
rect 1598 1178 1604 1179
rect 1618 1178 1624 1179
rect 1702 1178 1708 1179
rect 1722 1178 1728 1179
rect 1806 1178 1812 1179
rect 1826 1178 1832 1179
rect 1910 1178 1916 1179
rect 1598 1174 1599 1178
rect 1603 1174 1604 1178
rect 1598 1173 1604 1174
rect 1582 1151 1588 1152
rect 1582 1147 1583 1151
rect 1587 1147 1588 1151
rect 1582 1146 1588 1147
rect 1494 1139 1500 1140
rect 1494 1135 1495 1139
rect 1499 1135 1500 1139
rect 1494 1134 1500 1135
rect 1584 1131 1586 1146
rect 1479 1130 1483 1131
rect 1479 1125 1483 1126
rect 1487 1130 1491 1131
rect 1487 1125 1491 1126
rect 1583 1130 1587 1131
rect 1583 1125 1587 1126
rect 1470 1115 1476 1116
rect 1470 1111 1471 1115
rect 1475 1111 1476 1115
rect 1480 1114 1482 1125
rect 1502 1115 1508 1116
rect 1470 1110 1476 1111
rect 1478 1113 1484 1114
rect 1472 1080 1474 1110
rect 1478 1109 1479 1113
rect 1483 1109 1484 1113
rect 1502 1111 1503 1115
rect 1507 1111 1508 1115
rect 1584 1114 1586 1125
rect 1620 1116 1622 1178
rect 1702 1174 1703 1178
rect 1707 1174 1708 1178
rect 1702 1173 1708 1174
rect 1686 1151 1692 1152
rect 1686 1147 1687 1151
rect 1691 1147 1692 1151
rect 1724 1148 1726 1178
rect 1806 1174 1807 1178
rect 1811 1174 1812 1178
rect 1806 1173 1812 1174
rect 1790 1151 1796 1152
rect 1686 1146 1692 1147
rect 1722 1147 1728 1148
rect 1688 1131 1690 1146
rect 1722 1143 1723 1147
rect 1727 1143 1728 1147
rect 1790 1147 1791 1151
rect 1795 1147 1796 1151
rect 1828 1148 1830 1178
rect 1910 1174 1911 1178
rect 1915 1174 1916 1178
rect 1910 1173 1916 1174
rect 1894 1151 1900 1152
rect 1790 1146 1796 1147
rect 1826 1147 1832 1148
rect 1722 1142 1728 1143
rect 1792 1131 1794 1146
rect 1826 1143 1827 1147
rect 1831 1143 1832 1147
rect 1894 1147 1895 1151
rect 1899 1147 1900 1151
rect 1928 1148 1930 1198
rect 1968 1191 1970 1205
rect 2008 1204 2010 1234
rect 2014 1233 2015 1237
rect 2019 1233 2020 1237
rect 2038 1235 2039 1239
rect 2043 1235 2044 1239
rect 2080 1238 2082 1249
rect 2086 1247 2092 1248
rect 2086 1243 2087 1247
rect 2091 1243 2092 1247
rect 2086 1242 2092 1243
rect 2038 1234 2044 1235
rect 2078 1237 2084 1238
rect 2014 1232 2020 1233
rect 2030 1210 2036 1211
rect 2030 1206 2031 1210
rect 2035 1206 2036 1210
rect 2030 1205 2036 1206
rect 2006 1203 2012 1204
rect 2006 1199 2007 1203
rect 2011 1199 2012 1203
rect 2006 1198 2012 1199
rect 2032 1191 2034 1205
rect 1967 1190 1971 1191
rect 1967 1185 1971 1186
rect 2015 1190 2019 1191
rect 2015 1185 2019 1186
rect 2031 1190 2035 1191
rect 2040 1188 2042 1234
rect 2078 1233 2079 1237
rect 2083 1233 2084 1237
rect 2078 1232 2084 1233
rect 2088 1204 2090 1242
rect 2138 1239 2144 1240
rect 2138 1235 2139 1239
rect 2143 1235 2144 1239
rect 2152 1238 2154 1249
rect 2188 1240 2190 1298
rect 2230 1294 2231 1298
rect 2235 1294 2236 1298
rect 2230 1293 2236 1294
rect 2214 1271 2220 1272
rect 2214 1267 2215 1271
rect 2219 1267 2220 1271
rect 2248 1268 2250 1306
rect 2583 1305 2587 1306
rect 2584 1290 2586 1305
rect 2582 1289 2588 1290
rect 2582 1285 2583 1289
rect 2587 1285 2588 1289
rect 2582 1284 2588 1285
rect 2582 1272 2588 1273
rect 2582 1268 2583 1272
rect 2587 1268 2588 1272
rect 2214 1266 2220 1267
rect 2246 1267 2252 1268
rect 2582 1267 2588 1268
rect 2216 1255 2218 1266
rect 2246 1263 2247 1267
rect 2251 1263 2252 1267
rect 2246 1262 2252 1263
rect 2584 1255 2586 1267
rect 2215 1254 2219 1255
rect 2215 1249 2219 1250
rect 2223 1254 2227 1255
rect 2223 1249 2227 1250
rect 2295 1254 2299 1255
rect 2295 1249 2299 1250
rect 2583 1254 2587 1255
rect 2583 1249 2587 1250
rect 2186 1239 2192 1240
rect 2138 1234 2144 1235
rect 2150 1237 2156 1238
rect 2094 1210 2100 1211
rect 2094 1206 2095 1210
rect 2099 1206 2100 1210
rect 2094 1205 2100 1206
rect 2086 1203 2092 1204
rect 2086 1199 2087 1203
rect 2091 1199 2092 1203
rect 2086 1198 2092 1199
rect 2096 1191 2098 1205
rect 2140 1204 2142 1234
rect 2150 1233 2151 1237
rect 2155 1233 2156 1237
rect 2186 1235 2187 1239
rect 2191 1235 2192 1239
rect 2224 1238 2226 1249
rect 2286 1239 2292 1240
rect 2186 1234 2192 1235
rect 2222 1237 2228 1238
rect 2150 1232 2156 1233
rect 2222 1233 2223 1237
rect 2227 1233 2228 1237
rect 2286 1235 2287 1239
rect 2291 1235 2292 1239
rect 2296 1238 2298 1249
rect 2286 1234 2292 1235
rect 2294 1237 2300 1238
rect 2584 1237 2586 1249
rect 2222 1232 2228 1233
rect 2166 1210 2172 1211
rect 2166 1206 2167 1210
rect 2171 1206 2172 1210
rect 2166 1205 2172 1206
rect 2238 1210 2244 1211
rect 2238 1206 2239 1210
rect 2243 1206 2244 1210
rect 2238 1205 2244 1206
rect 2138 1203 2144 1204
rect 2138 1199 2139 1203
rect 2143 1199 2144 1203
rect 2138 1198 2144 1199
rect 2168 1191 2170 1205
rect 2218 1203 2224 1204
rect 2218 1199 2219 1203
rect 2223 1199 2224 1203
rect 2218 1198 2224 1199
rect 2095 1190 2099 1191
rect 2031 1185 2035 1186
rect 2038 1187 2044 1188
rect 2016 1179 2018 1185
rect 2038 1183 2039 1187
rect 2043 1183 2044 1187
rect 2095 1185 2099 1186
rect 2111 1190 2115 1191
rect 2111 1185 2115 1186
rect 2167 1190 2171 1191
rect 2167 1185 2171 1186
rect 2207 1190 2211 1191
rect 2207 1185 2211 1186
rect 2038 1182 2044 1183
rect 2086 1183 2092 1184
rect 2086 1179 2087 1183
rect 2091 1179 2092 1183
rect 2112 1179 2114 1185
rect 2130 1183 2136 1184
rect 2130 1179 2131 1183
rect 2135 1179 2136 1183
rect 2208 1179 2210 1185
rect 2014 1178 2020 1179
rect 2086 1178 2092 1179
rect 2110 1178 2116 1179
rect 2130 1178 2136 1179
rect 2206 1178 2212 1179
rect 2014 1174 2015 1178
rect 2019 1174 2020 1178
rect 2014 1173 2020 1174
rect 2088 1160 2090 1178
rect 2110 1174 2111 1178
rect 2115 1174 2116 1178
rect 2110 1173 2116 1174
rect 2086 1159 2092 1160
rect 2086 1155 2087 1159
rect 2091 1155 2092 1159
rect 2086 1154 2092 1155
rect 1998 1151 2004 1152
rect 1894 1146 1900 1147
rect 1926 1147 1932 1148
rect 1826 1142 1832 1143
rect 1896 1131 1898 1146
rect 1926 1143 1927 1147
rect 1931 1143 1932 1147
rect 1998 1147 1999 1151
rect 2003 1147 2004 1151
rect 1998 1146 2004 1147
rect 2094 1151 2100 1152
rect 2094 1147 2095 1151
rect 2099 1147 2100 1151
rect 2132 1148 2134 1178
rect 2206 1174 2207 1178
rect 2211 1174 2212 1178
rect 2206 1173 2212 1174
rect 2190 1151 2196 1152
rect 2094 1146 2100 1147
rect 2130 1147 2136 1148
rect 1926 1142 1932 1143
rect 2000 1131 2002 1146
rect 2096 1131 2098 1146
rect 2130 1143 2131 1147
rect 2135 1143 2136 1147
rect 2190 1147 2191 1151
rect 2195 1147 2196 1151
rect 2220 1148 2222 1198
rect 2240 1191 2242 1205
rect 2288 1204 2290 1234
rect 2294 1233 2295 1237
rect 2299 1233 2300 1237
rect 2294 1232 2300 1233
rect 2582 1236 2588 1237
rect 2582 1232 2583 1236
rect 2587 1232 2588 1236
rect 2582 1231 2588 1232
rect 2582 1219 2588 1220
rect 2582 1215 2583 1219
rect 2587 1215 2588 1219
rect 2582 1214 2588 1215
rect 2310 1210 2316 1211
rect 2310 1206 2311 1210
rect 2315 1206 2316 1210
rect 2310 1205 2316 1206
rect 2286 1203 2292 1204
rect 2286 1199 2287 1203
rect 2291 1199 2292 1203
rect 2286 1198 2292 1199
rect 2312 1191 2314 1205
rect 2584 1191 2586 1214
rect 2239 1190 2243 1191
rect 2239 1185 2243 1186
rect 2303 1190 2307 1191
rect 2303 1185 2307 1186
rect 2311 1190 2315 1191
rect 2311 1185 2315 1186
rect 2399 1190 2403 1191
rect 2399 1185 2403 1186
rect 2583 1190 2587 1191
rect 2583 1185 2587 1186
rect 2294 1183 2300 1184
rect 2294 1179 2295 1183
rect 2299 1179 2300 1183
rect 2304 1179 2306 1185
rect 2322 1183 2328 1184
rect 2322 1179 2323 1183
rect 2327 1179 2328 1183
rect 2400 1179 2402 1185
rect 2294 1178 2300 1179
rect 2302 1178 2308 1179
rect 2322 1178 2328 1179
rect 2398 1178 2404 1179
rect 2286 1151 2292 1152
rect 2190 1146 2196 1147
rect 2218 1147 2224 1148
rect 2130 1142 2136 1143
rect 2192 1131 2194 1146
rect 2218 1143 2219 1147
rect 2223 1143 2224 1147
rect 2286 1147 2287 1151
rect 2291 1147 2292 1151
rect 2286 1146 2292 1147
rect 2218 1142 2224 1143
rect 2288 1131 2290 1146
rect 1687 1130 1691 1131
rect 1687 1125 1691 1126
rect 1791 1130 1795 1131
rect 1791 1125 1795 1126
rect 1887 1130 1891 1131
rect 1887 1125 1891 1126
rect 1895 1130 1899 1131
rect 1895 1125 1899 1126
rect 1975 1130 1979 1131
rect 1975 1125 1979 1126
rect 1999 1130 2003 1131
rect 1999 1125 2003 1126
rect 2063 1130 2067 1131
rect 2063 1125 2067 1126
rect 2095 1130 2099 1131
rect 2095 1125 2099 1126
rect 2143 1130 2147 1131
rect 2143 1125 2147 1126
rect 2191 1130 2195 1131
rect 2191 1125 2195 1126
rect 2215 1130 2219 1131
rect 2215 1125 2219 1126
rect 2279 1130 2283 1131
rect 2279 1125 2283 1126
rect 2287 1130 2291 1131
rect 2287 1125 2291 1126
rect 1626 1119 1632 1120
rect 1618 1115 1624 1116
rect 1502 1110 1508 1111
rect 1582 1113 1588 1114
rect 1478 1108 1484 1109
rect 1494 1086 1500 1087
rect 1494 1082 1495 1086
rect 1499 1082 1500 1086
rect 1494 1081 1500 1082
rect 1422 1079 1428 1080
rect 1422 1075 1423 1079
rect 1427 1075 1428 1079
rect 1422 1074 1428 1075
rect 1470 1079 1476 1080
rect 1470 1075 1471 1079
rect 1475 1075 1476 1079
rect 1470 1074 1476 1075
rect 1496 1071 1498 1081
rect 1367 1070 1371 1071
rect 1095 1066 1099 1067
rect 1095 1061 1099 1062
rect 1135 1066 1139 1067
rect 1135 1061 1139 1062
rect 1183 1066 1187 1067
rect 1183 1061 1187 1062
rect 1223 1066 1227 1067
rect 1223 1061 1227 1062
rect 1287 1066 1291 1067
rect 1287 1061 1291 1062
rect 1327 1066 1331 1067
rect 1367 1065 1371 1066
rect 1415 1070 1419 1071
rect 1415 1065 1419 1066
rect 1471 1070 1475 1071
rect 1471 1065 1475 1066
rect 1495 1070 1499 1071
rect 1504 1068 1506 1110
rect 1582 1109 1583 1113
rect 1587 1109 1588 1113
rect 1618 1111 1619 1115
rect 1623 1111 1624 1115
rect 1626 1115 1627 1119
rect 1631 1115 1632 1119
rect 1626 1114 1632 1115
rect 1688 1114 1690 1125
rect 1792 1114 1794 1125
rect 1888 1114 1890 1125
rect 1966 1115 1972 1116
rect 1618 1110 1624 1111
rect 1582 1108 1588 1109
rect 1598 1086 1604 1087
rect 1598 1082 1599 1086
rect 1603 1082 1604 1086
rect 1598 1081 1604 1082
rect 1600 1071 1602 1081
rect 1628 1080 1630 1114
rect 1686 1113 1692 1114
rect 1686 1109 1687 1113
rect 1691 1109 1692 1113
rect 1686 1108 1692 1109
rect 1790 1113 1796 1114
rect 1790 1109 1791 1113
rect 1795 1109 1796 1113
rect 1790 1108 1796 1109
rect 1886 1113 1892 1114
rect 1886 1109 1887 1113
rect 1891 1109 1892 1113
rect 1966 1111 1967 1115
rect 1971 1111 1972 1115
rect 1976 1114 1978 1125
rect 2038 1115 2044 1116
rect 1966 1110 1972 1111
rect 1974 1113 1980 1114
rect 1886 1108 1892 1109
rect 1702 1086 1708 1087
rect 1702 1082 1703 1086
rect 1707 1082 1708 1086
rect 1702 1081 1708 1082
rect 1806 1086 1812 1087
rect 1806 1082 1807 1086
rect 1811 1082 1812 1086
rect 1806 1081 1812 1082
rect 1902 1086 1908 1087
rect 1902 1082 1903 1086
rect 1907 1082 1908 1086
rect 1902 1081 1908 1082
rect 1626 1079 1632 1080
rect 1626 1075 1627 1079
rect 1631 1075 1632 1079
rect 1626 1074 1632 1075
rect 1704 1071 1706 1081
rect 1808 1071 1810 1081
rect 1854 1079 1860 1080
rect 1854 1075 1855 1079
rect 1859 1075 1860 1079
rect 1854 1074 1860 1075
rect 1535 1070 1539 1071
rect 1495 1065 1499 1066
rect 1502 1067 1508 1068
rect 1327 1061 1331 1062
rect 1136 1055 1138 1061
rect 1154 1059 1160 1060
rect 1154 1055 1155 1059
rect 1159 1055 1160 1059
rect 1224 1055 1226 1061
rect 1288 1055 1290 1061
rect 1134 1054 1140 1055
rect 1154 1054 1160 1055
rect 1222 1054 1228 1055
rect 1134 1050 1135 1054
rect 1139 1050 1140 1054
rect 1134 1049 1140 1050
rect 1118 1027 1124 1028
rect 1070 1023 1076 1024
rect 1070 1019 1071 1023
rect 1075 1019 1076 1023
rect 1118 1023 1119 1027
rect 1123 1023 1124 1027
rect 1156 1024 1158 1054
rect 1222 1050 1223 1054
rect 1227 1050 1228 1054
rect 1222 1049 1228 1050
rect 1286 1054 1292 1055
rect 1286 1050 1287 1054
rect 1291 1050 1292 1054
rect 1286 1049 1292 1050
rect 1328 1046 1330 1061
rect 1368 1050 1370 1065
rect 1416 1059 1418 1065
rect 1472 1059 1474 1065
rect 1502 1063 1503 1067
rect 1507 1063 1508 1067
rect 1535 1065 1539 1066
rect 1599 1070 1603 1071
rect 1599 1065 1603 1066
rect 1623 1070 1627 1071
rect 1623 1065 1627 1066
rect 1703 1070 1707 1071
rect 1703 1065 1707 1066
rect 1727 1070 1731 1071
rect 1727 1065 1731 1066
rect 1807 1070 1811 1071
rect 1807 1065 1811 1066
rect 1839 1070 1843 1071
rect 1839 1065 1843 1066
rect 1502 1062 1508 1063
rect 1526 1063 1532 1064
rect 1526 1059 1527 1063
rect 1531 1059 1532 1063
rect 1536 1059 1538 1065
rect 1554 1063 1560 1064
rect 1554 1059 1555 1063
rect 1559 1059 1560 1063
rect 1624 1059 1626 1065
rect 1642 1063 1648 1064
rect 1642 1059 1643 1063
rect 1647 1059 1648 1063
rect 1728 1059 1730 1065
rect 1746 1063 1752 1064
rect 1746 1059 1747 1063
rect 1751 1059 1752 1063
rect 1840 1059 1842 1065
rect 1414 1058 1420 1059
rect 1414 1054 1415 1058
rect 1419 1054 1420 1058
rect 1414 1053 1420 1054
rect 1470 1058 1476 1059
rect 1526 1058 1532 1059
rect 1534 1058 1540 1059
rect 1554 1058 1560 1059
rect 1622 1058 1628 1059
rect 1642 1058 1648 1059
rect 1726 1058 1732 1059
rect 1746 1058 1752 1059
rect 1838 1058 1844 1059
rect 1470 1054 1471 1058
rect 1475 1054 1476 1058
rect 1470 1053 1476 1054
rect 1366 1049 1372 1050
rect 1326 1045 1332 1046
rect 1326 1041 1327 1045
rect 1331 1041 1332 1045
rect 1366 1045 1367 1049
rect 1371 1045 1372 1049
rect 1366 1044 1372 1045
rect 1326 1040 1332 1041
rect 1366 1032 1372 1033
rect 1235 1028 1239 1029
rect 1326 1028 1332 1029
rect 1206 1027 1212 1028
rect 1118 1022 1124 1023
rect 1154 1023 1160 1024
rect 1070 1018 1076 1019
rect 1062 1011 1068 1012
rect 1062 1007 1063 1011
rect 1067 1007 1068 1011
rect 1120 1007 1122 1022
rect 1154 1019 1155 1023
rect 1159 1019 1160 1023
rect 1206 1023 1207 1027
rect 1211 1023 1212 1027
rect 1270 1027 1276 1028
rect 1206 1022 1212 1023
rect 1234 1023 1240 1024
rect 1154 1018 1160 1019
rect 1208 1007 1210 1022
rect 1234 1019 1235 1023
rect 1239 1019 1240 1023
rect 1270 1023 1271 1027
rect 1275 1023 1276 1027
rect 1326 1024 1327 1028
rect 1331 1024 1332 1028
rect 1366 1028 1367 1032
rect 1371 1028 1372 1032
rect 1366 1027 1372 1028
rect 1398 1031 1404 1032
rect 1398 1027 1399 1031
rect 1403 1027 1404 1031
rect 1270 1022 1276 1023
rect 1294 1023 1300 1024
rect 1326 1023 1332 1024
rect 1234 1018 1240 1019
rect 1272 1007 1274 1022
rect 1294 1019 1295 1023
rect 1299 1019 1300 1023
rect 1294 1018 1300 1019
rect 783 1006 787 1007
rect 783 1001 787 1002
rect 847 1006 851 1007
rect 847 1001 851 1002
rect 871 1006 875 1007
rect 871 1001 875 1002
rect 911 1006 915 1007
rect 946 1006 952 1007
rect 959 1006 963 1007
rect 911 1001 915 1002
rect 784 990 786 1001
rect 806 999 812 1000
rect 806 995 807 999
rect 811 995 812 999
rect 806 994 812 995
rect 782 989 788 990
rect 782 985 783 989
rect 787 985 788 989
rect 782 984 788 985
rect 798 962 804 963
rect 798 958 799 962
rect 803 958 804 962
rect 798 957 804 958
rect 754 955 760 956
rect 754 951 755 955
rect 759 951 760 955
rect 754 950 760 951
rect 800 947 802 957
rect 808 956 810 994
rect 838 991 844 992
rect 838 987 839 991
rect 843 987 844 991
rect 848 990 850 1001
rect 902 991 908 992
rect 838 986 844 987
rect 846 989 852 990
rect 840 956 842 986
rect 846 985 847 989
rect 851 985 852 989
rect 902 987 903 991
rect 907 987 908 991
rect 912 990 914 1001
rect 948 992 950 1006
rect 959 1001 963 1002
rect 975 1006 979 1007
rect 975 1001 979 1002
rect 1039 1006 1043 1007
rect 1062 1006 1068 1007
rect 1103 1006 1107 1007
rect 1039 1001 1043 1002
rect 1103 1001 1107 1002
rect 1119 1006 1123 1007
rect 1119 1001 1123 1002
rect 1159 1006 1163 1007
rect 1159 1001 1163 1002
rect 1207 1006 1211 1007
rect 1207 1001 1211 1002
rect 1215 1006 1219 1007
rect 1215 1001 1219 1002
rect 1271 1006 1275 1007
rect 1271 1001 1275 1002
rect 946 991 952 992
rect 902 986 908 987
rect 910 989 916 990
rect 846 984 852 985
rect 862 962 868 963
rect 862 958 863 962
rect 867 958 868 962
rect 862 957 868 958
rect 806 955 812 956
rect 806 951 807 955
rect 811 951 812 955
rect 806 950 812 951
rect 838 955 844 956
rect 838 951 839 955
rect 843 951 844 955
rect 838 950 844 951
rect 864 947 866 957
rect 904 956 906 986
rect 910 985 911 989
rect 915 985 916 989
rect 946 987 947 991
rect 951 987 952 991
rect 976 990 978 1001
rect 1040 990 1042 1001
rect 1104 990 1106 1001
rect 1160 990 1162 1001
rect 1216 990 1218 1001
rect 1272 990 1274 1001
rect 946 986 952 987
rect 974 989 980 990
rect 910 984 916 985
rect 974 985 975 989
rect 979 985 980 989
rect 974 984 980 985
rect 1038 989 1044 990
rect 1038 985 1039 989
rect 1043 985 1044 989
rect 1038 984 1044 985
rect 1102 989 1108 990
rect 1102 985 1103 989
rect 1107 985 1108 989
rect 1102 984 1108 985
rect 1158 989 1164 990
rect 1158 985 1159 989
rect 1163 985 1164 989
rect 1158 984 1164 985
rect 1214 989 1220 990
rect 1214 985 1215 989
rect 1219 985 1220 989
rect 1214 984 1220 985
rect 1270 989 1276 990
rect 1270 985 1271 989
rect 1275 985 1276 989
rect 1270 984 1276 985
rect 926 962 932 963
rect 926 958 927 962
rect 931 958 932 962
rect 926 957 932 958
rect 990 962 996 963
rect 990 958 991 962
rect 995 958 996 962
rect 990 957 996 958
rect 1054 962 1060 963
rect 1054 958 1055 962
rect 1059 958 1060 962
rect 1054 957 1060 958
rect 1118 962 1124 963
rect 1118 958 1119 962
rect 1123 958 1124 962
rect 1118 957 1124 958
rect 1174 962 1180 963
rect 1174 958 1175 962
rect 1179 958 1180 962
rect 1174 957 1180 958
rect 1230 962 1236 963
rect 1230 958 1231 962
rect 1235 958 1236 962
rect 1230 957 1236 958
rect 1286 962 1292 963
rect 1286 958 1287 962
rect 1291 958 1292 962
rect 1286 957 1292 958
rect 902 955 908 956
rect 902 951 903 955
rect 907 951 908 955
rect 902 950 908 951
rect 928 947 930 957
rect 992 947 994 957
rect 1056 947 1058 957
rect 1120 947 1122 957
rect 1176 947 1178 957
rect 1232 947 1234 957
rect 1288 947 1290 957
rect 1296 956 1298 1018
rect 1328 1007 1330 1023
rect 1327 1006 1331 1007
rect 1327 1001 1331 1002
rect 1328 989 1330 1001
rect 1368 999 1370 1027
rect 1398 1026 1404 1027
rect 1454 1031 1460 1032
rect 1454 1027 1455 1031
rect 1459 1027 1460 1031
rect 1454 1026 1460 1027
rect 1518 1031 1524 1032
rect 1518 1027 1519 1031
rect 1523 1027 1524 1031
rect 1518 1026 1524 1027
rect 1400 999 1402 1026
rect 1456 999 1458 1026
rect 1520 999 1522 1026
rect 1367 998 1371 999
rect 1367 993 1371 994
rect 1399 998 1403 999
rect 1399 993 1403 994
rect 1455 998 1459 999
rect 1455 993 1459 994
rect 1511 998 1515 999
rect 1511 993 1515 994
rect 1519 998 1523 999
rect 1519 993 1523 994
rect 1326 988 1332 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1368 981 1370 993
rect 1400 982 1402 993
rect 1446 983 1452 984
rect 1398 981 1404 982
rect 1366 980 1372 981
rect 1366 976 1367 980
rect 1371 976 1372 980
rect 1398 977 1399 981
rect 1403 977 1404 981
rect 1446 979 1447 983
rect 1451 979 1452 983
rect 1456 982 1458 993
rect 1502 983 1508 984
rect 1446 978 1452 979
rect 1454 981 1460 982
rect 1398 976 1404 977
rect 1366 975 1372 976
rect 1326 971 1332 972
rect 1326 967 1327 971
rect 1331 967 1332 971
rect 1326 966 1332 967
rect 1294 955 1300 956
rect 1294 951 1295 955
rect 1299 951 1300 955
rect 1294 950 1300 951
rect 1328 947 1330 966
rect 1366 963 1372 964
rect 1366 959 1367 963
rect 1371 959 1372 963
rect 1366 958 1372 959
rect 759 946 763 947
rect 735 941 739 942
rect 746 943 752 944
rect 678 939 684 940
rect 678 935 679 939
rect 683 935 684 939
rect 704 935 706 941
rect 746 939 747 943
rect 751 939 752 943
rect 759 941 763 942
rect 799 946 803 947
rect 799 941 803 942
rect 815 946 819 947
rect 815 941 819 942
rect 863 946 867 947
rect 863 941 867 942
rect 927 946 931 947
rect 927 941 931 942
rect 991 946 995 947
rect 991 941 995 942
rect 1055 946 1059 947
rect 1055 941 1059 942
rect 1119 946 1123 947
rect 1119 941 1123 942
rect 1175 946 1179 947
rect 1175 941 1179 942
rect 1231 946 1235 947
rect 1231 941 1235 942
rect 1287 946 1291 947
rect 1287 941 1291 942
rect 1327 946 1331 947
rect 1327 941 1331 942
rect 746 938 752 939
rect 760 935 762 941
rect 778 939 784 940
rect 778 935 779 939
rect 783 935 784 939
rect 816 935 818 941
rect 678 934 684 935
rect 702 934 708 935
rect 680 916 682 934
rect 702 930 703 934
rect 707 930 708 934
rect 702 929 708 930
rect 758 934 764 935
rect 778 934 784 935
rect 814 934 820 935
rect 758 930 759 934
rect 763 930 764 934
rect 758 929 764 930
rect 678 915 684 916
rect 678 911 679 915
rect 683 911 684 915
rect 678 910 684 911
rect 686 907 692 908
rect 630 902 636 903
rect 662 903 668 904
rect 554 898 560 899
rect 576 891 578 902
rect 632 891 634 902
rect 662 899 663 903
rect 667 899 668 903
rect 686 903 687 907
rect 691 903 692 907
rect 686 902 692 903
rect 742 907 748 908
rect 742 903 743 907
rect 747 903 748 907
rect 780 904 782 934
rect 814 930 815 934
rect 819 930 820 934
rect 814 929 820 930
rect 1328 926 1330 941
rect 1368 935 1370 958
rect 1414 954 1420 955
rect 1414 950 1415 954
rect 1419 950 1420 954
rect 1414 949 1420 950
rect 1416 935 1418 949
rect 1448 948 1450 978
rect 1454 977 1455 981
rect 1459 977 1460 981
rect 1502 979 1503 983
rect 1507 979 1508 983
rect 1512 982 1514 993
rect 1528 992 1530 1058
rect 1534 1054 1535 1058
rect 1539 1054 1540 1058
rect 1534 1053 1540 1054
rect 1556 1028 1558 1058
rect 1622 1054 1623 1058
rect 1627 1054 1628 1058
rect 1622 1053 1628 1054
rect 1606 1031 1612 1032
rect 1554 1027 1560 1028
rect 1554 1023 1555 1027
rect 1559 1023 1560 1027
rect 1606 1027 1607 1031
rect 1611 1027 1612 1031
rect 1644 1028 1646 1058
rect 1726 1054 1727 1058
rect 1731 1054 1732 1058
rect 1726 1053 1732 1054
rect 1710 1031 1716 1032
rect 1606 1026 1612 1027
rect 1642 1027 1648 1028
rect 1554 1022 1560 1023
rect 1608 999 1610 1026
rect 1642 1023 1643 1027
rect 1647 1023 1648 1027
rect 1710 1027 1711 1031
rect 1715 1027 1716 1031
rect 1748 1028 1750 1058
rect 1838 1054 1839 1058
rect 1843 1054 1844 1058
rect 1838 1053 1844 1054
rect 1822 1031 1828 1032
rect 1710 1026 1716 1027
rect 1746 1027 1752 1028
rect 1642 1022 1648 1023
rect 1712 999 1714 1026
rect 1746 1023 1747 1027
rect 1751 1023 1752 1027
rect 1822 1027 1823 1031
rect 1827 1027 1828 1031
rect 1856 1028 1858 1074
rect 1904 1071 1906 1081
rect 1968 1080 1970 1110
rect 1974 1109 1975 1113
rect 1979 1109 1980 1113
rect 2038 1111 2039 1115
rect 2043 1111 2044 1115
rect 2064 1114 2066 1125
rect 2134 1115 2140 1116
rect 2038 1110 2044 1111
rect 2062 1113 2068 1114
rect 1974 1108 1980 1109
rect 1990 1086 1996 1087
rect 1990 1082 1991 1086
rect 1995 1082 1996 1086
rect 1990 1081 1996 1082
rect 1966 1079 1972 1080
rect 1966 1075 1967 1079
rect 1971 1075 1972 1079
rect 1966 1074 1972 1075
rect 1992 1071 1994 1081
rect 1903 1070 1907 1071
rect 1903 1065 1907 1066
rect 1951 1070 1955 1071
rect 1951 1065 1955 1066
rect 1991 1070 1995 1071
rect 1991 1065 1995 1066
rect 1926 1063 1932 1064
rect 1926 1059 1927 1063
rect 1931 1059 1932 1063
rect 1952 1059 1954 1065
rect 2040 1064 2042 1110
rect 2062 1109 2063 1113
rect 2067 1109 2068 1113
rect 2134 1111 2135 1115
rect 2139 1111 2140 1115
rect 2144 1114 2146 1125
rect 2206 1115 2212 1116
rect 2134 1110 2140 1111
rect 2142 1113 2148 1114
rect 2062 1108 2068 1109
rect 2078 1086 2084 1087
rect 2078 1082 2079 1086
rect 2083 1082 2084 1086
rect 2078 1081 2084 1082
rect 2080 1071 2082 1081
rect 2136 1080 2138 1110
rect 2142 1109 2143 1113
rect 2147 1109 2148 1113
rect 2206 1111 2207 1115
rect 2211 1111 2212 1115
rect 2216 1114 2218 1125
rect 2270 1115 2276 1116
rect 2206 1110 2212 1111
rect 2214 1113 2220 1114
rect 2142 1108 2148 1109
rect 2158 1086 2164 1087
rect 2158 1082 2159 1086
rect 2163 1082 2164 1086
rect 2158 1081 2164 1082
rect 2126 1079 2132 1080
rect 2126 1075 2127 1079
rect 2131 1075 2132 1079
rect 2126 1074 2132 1075
rect 2134 1079 2140 1080
rect 2134 1075 2135 1079
rect 2139 1075 2140 1079
rect 2134 1074 2140 1075
rect 2063 1070 2067 1071
rect 2063 1065 2067 1066
rect 2079 1070 2083 1071
rect 2079 1065 2083 1066
rect 2038 1063 2044 1064
rect 2038 1059 2039 1063
rect 2043 1059 2044 1063
rect 2064 1059 2066 1065
rect 1926 1058 1932 1059
rect 1950 1058 1956 1059
rect 2038 1058 2044 1059
rect 2062 1058 2068 1059
rect 1928 1040 1930 1058
rect 1950 1054 1951 1058
rect 1955 1054 1956 1058
rect 1950 1053 1956 1054
rect 2062 1054 2063 1058
rect 2067 1054 2068 1058
rect 2062 1053 2068 1054
rect 1926 1039 1932 1040
rect 1926 1035 1927 1039
rect 1931 1035 1932 1039
rect 1926 1034 1932 1035
rect 1934 1031 1940 1032
rect 1822 1026 1828 1027
rect 1854 1027 1860 1028
rect 1746 1022 1752 1023
rect 1824 999 1826 1026
rect 1854 1023 1855 1027
rect 1859 1023 1860 1027
rect 1934 1027 1935 1031
rect 1939 1027 1940 1031
rect 1934 1026 1940 1027
rect 2046 1031 2052 1032
rect 2046 1027 2047 1031
rect 2051 1027 2052 1031
rect 2046 1026 2052 1027
rect 1854 1022 1860 1023
rect 1936 999 1938 1026
rect 2048 999 2050 1026
rect 2128 1024 2130 1074
rect 2160 1071 2162 1081
rect 2208 1080 2210 1110
rect 2214 1109 2215 1113
rect 2219 1109 2220 1113
rect 2270 1111 2271 1115
rect 2275 1111 2276 1115
rect 2280 1114 2282 1125
rect 2296 1120 2298 1178
rect 2302 1174 2303 1178
rect 2307 1174 2308 1178
rect 2302 1173 2308 1174
rect 2324 1148 2326 1178
rect 2398 1174 2399 1178
rect 2403 1174 2404 1178
rect 2398 1173 2404 1174
rect 2584 1170 2586 1185
rect 2582 1169 2588 1170
rect 2582 1165 2583 1169
rect 2587 1165 2588 1169
rect 2582 1164 2588 1165
rect 2582 1152 2588 1153
rect 2382 1151 2388 1152
rect 2322 1147 2328 1148
rect 2322 1143 2323 1147
rect 2327 1143 2328 1147
rect 2382 1147 2383 1151
rect 2387 1147 2388 1151
rect 2582 1148 2583 1152
rect 2587 1148 2588 1152
rect 2582 1147 2588 1148
rect 2382 1146 2388 1147
rect 2322 1142 2328 1143
rect 2384 1131 2386 1146
rect 2584 1131 2586 1147
rect 2343 1130 2347 1131
rect 2343 1125 2347 1126
rect 2383 1130 2387 1131
rect 2383 1125 2387 1126
rect 2407 1130 2411 1131
rect 2407 1125 2411 1126
rect 2471 1130 2475 1131
rect 2471 1125 2475 1126
rect 2527 1130 2531 1131
rect 2527 1125 2531 1126
rect 2583 1130 2587 1131
rect 2583 1125 2587 1126
rect 2294 1119 2300 1120
rect 2294 1115 2295 1119
rect 2299 1115 2300 1119
rect 2294 1114 2300 1115
rect 2344 1114 2346 1125
rect 2374 1115 2380 1116
rect 2270 1110 2276 1111
rect 2278 1113 2284 1114
rect 2214 1108 2220 1109
rect 2230 1086 2236 1087
rect 2230 1082 2231 1086
rect 2235 1082 2236 1086
rect 2230 1081 2236 1082
rect 2206 1079 2212 1080
rect 2206 1075 2207 1079
rect 2211 1075 2212 1079
rect 2206 1074 2212 1075
rect 2232 1071 2234 1081
rect 2272 1080 2274 1110
rect 2278 1109 2279 1113
rect 2283 1109 2284 1113
rect 2278 1108 2284 1109
rect 2342 1113 2348 1114
rect 2342 1109 2343 1113
rect 2347 1109 2348 1113
rect 2374 1111 2375 1115
rect 2379 1111 2380 1115
rect 2408 1114 2410 1125
rect 2438 1123 2444 1124
rect 2438 1119 2439 1123
rect 2443 1119 2444 1123
rect 2438 1118 2444 1119
rect 2374 1110 2380 1111
rect 2406 1113 2412 1114
rect 2342 1108 2348 1109
rect 2294 1086 2300 1087
rect 2294 1082 2295 1086
rect 2299 1082 2300 1086
rect 2294 1081 2300 1082
rect 2358 1086 2364 1087
rect 2358 1082 2359 1086
rect 2363 1082 2364 1086
rect 2358 1081 2364 1082
rect 2270 1079 2276 1080
rect 2270 1075 2271 1079
rect 2275 1075 2276 1079
rect 2270 1074 2276 1075
rect 2286 1071 2292 1072
rect 2296 1071 2298 1081
rect 2360 1071 2362 1081
rect 2159 1070 2163 1071
rect 2159 1065 2163 1066
rect 2167 1070 2171 1071
rect 2167 1065 2171 1066
rect 2231 1070 2235 1071
rect 2231 1065 2235 1066
rect 2271 1070 2275 1071
rect 2286 1067 2287 1071
rect 2291 1067 2292 1071
rect 2286 1066 2292 1067
rect 2295 1070 2299 1071
rect 2271 1065 2275 1066
rect 2168 1059 2170 1065
rect 2246 1063 2252 1064
rect 2246 1059 2247 1063
rect 2251 1059 2252 1063
rect 2272 1059 2274 1065
rect 2166 1058 2172 1059
rect 2246 1058 2252 1059
rect 2270 1058 2276 1059
rect 2166 1054 2167 1058
rect 2171 1054 2172 1058
rect 2166 1053 2172 1054
rect 2248 1040 2250 1058
rect 2270 1054 2271 1058
rect 2275 1054 2276 1058
rect 2270 1053 2276 1054
rect 2246 1039 2252 1040
rect 2246 1035 2247 1039
rect 2251 1035 2252 1039
rect 2246 1034 2252 1035
rect 2150 1031 2156 1032
rect 2150 1027 2151 1031
rect 2155 1027 2156 1031
rect 2150 1026 2156 1027
rect 2254 1031 2260 1032
rect 2254 1027 2255 1031
rect 2259 1027 2260 1031
rect 2288 1028 2290 1066
rect 2295 1065 2299 1066
rect 2359 1070 2363 1071
rect 2359 1065 2363 1066
rect 2367 1070 2371 1071
rect 2376 1068 2378 1110
rect 2406 1109 2407 1113
rect 2411 1109 2412 1113
rect 2406 1108 2412 1109
rect 2422 1086 2428 1087
rect 2422 1082 2423 1086
rect 2427 1082 2428 1086
rect 2422 1081 2428 1082
rect 2424 1071 2426 1081
rect 2440 1080 2442 1118
rect 2472 1114 2474 1125
rect 2518 1115 2524 1116
rect 2470 1113 2476 1114
rect 2470 1109 2471 1113
rect 2475 1109 2476 1113
rect 2518 1111 2519 1115
rect 2523 1111 2524 1115
rect 2528 1114 2530 1125
rect 2518 1110 2524 1111
rect 2526 1113 2532 1114
rect 2584 1113 2586 1125
rect 2470 1108 2476 1109
rect 2486 1086 2492 1087
rect 2486 1082 2487 1086
rect 2491 1082 2492 1086
rect 2486 1081 2492 1082
rect 2438 1079 2444 1080
rect 2438 1075 2439 1079
rect 2443 1075 2444 1079
rect 2438 1074 2444 1075
rect 2478 1079 2484 1080
rect 2478 1075 2479 1079
rect 2483 1075 2484 1079
rect 2478 1074 2484 1075
rect 2423 1070 2427 1071
rect 2367 1065 2371 1066
rect 2374 1067 2380 1068
rect 2368 1059 2370 1065
rect 2374 1063 2375 1067
rect 2379 1063 2380 1067
rect 2423 1065 2427 1066
rect 2463 1070 2467 1071
rect 2463 1065 2467 1066
rect 2374 1062 2380 1063
rect 2438 1063 2444 1064
rect 2438 1059 2439 1063
rect 2443 1059 2444 1063
rect 2464 1059 2466 1065
rect 2366 1058 2372 1059
rect 2438 1058 2444 1059
rect 2462 1058 2468 1059
rect 2366 1054 2367 1058
rect 2371 1054 2372 1058
rect 2366 1053 2372 1054
rect 2440 1040 2442 1058
rect 2462 1054 2463 1058
rect 2467 1054 2468 1058
rect 2462 1053 2468 1054
rect 2438 1039 2444 1040
rect 2438 1035 2439 1039
rect 2443 1035 2444 1039
rect 2438 1034 2444 1035
rect 2350 1031 2356 1032
rect 2254 1026 2260 1027
rect 2286 1027 2292 1028
rect 2126 1023 2132 1024
rect 2126 1019 2127 1023
rect 2131 1019 2132 1023
rect 2126 1018 2132 1019
rect 2152 999 2154 1026
rect 2256 999 2258 1026
rect 2286 1023 2287 1027
rect 2291 1023 2292 1027
rect 2350 1027 2351 1031
rect 2355 1027 2356 1031
rect 2350 1026 2356 1027
rect 2446 1031 2452 1032
rect 2446 1027 2447 1031
rect 2451 1027 2452 1031
rect 2480 1028 2482 1074
rect 2488 1071 2490 1081
rect 2520 1080 2522 1110
rect 2526 1109 2527 1113
rect 2531 1109 2532 1113
rect 2526 1108 2532 1109
rect 2582 1112 2588 1113
rect 2582 1108 2583 1112
rect 2587 1108 2588 1112
rect 2582 1107 2588 1108
rect 2582 1095 2588 1096
rect 2582 1091 2583 1095
rect 2587 1091 2588 1095
rect 2582 1090 2588 1091
rect 2542 1086 2548 1087
rect 2542 1082 2543 1086
rect 2547 1082 2548 1086
rect 2542 1081 2548 1082
rect 2518 1079 2524 1080
rect 2518 1075 2519 1079
rect 2523 1075 2524 1079
rect 2518 1074 2524 1075
rect 2544 1071 2546 1081
rect 2584 1071 2586 1090
rect 2487 1070 2491 1071
rect 2487 1065 2491 1066
rect 2543 1070 2547 1071
rect 2543 1065 2547 1066
rect 2583 1070 2587 1071
rect 2583 1065 2587 1066
rect 2534 1063 2540 1064
rect 2534 1059 2535 1063
rect 2539 1059 2540 1063
rect 2544 1059 2546 1065
rect 2534 1058 2540 1059
rect 2542 1058 2548 1059
rect 2526 1031 2532 1032
rect 2446 1026 2452 1027
rect 2478 1027 2484 1028
rect 2286 1022 2292 1023
rect 2352 999 2354 1026
rect 2448 999 2450 1026
rect 2478 1023 2479 1027
rect 2483 1023 2484 1027
rect 2526 1027 2527 1031
rect 2531 1027 2532 1031
rect 2526 1026 2532 1027
rect 2478 1022 2484 1023
rect 2528 999 2530 1026
rect 1567 998 1571 999
rect 1567 993 1571 994
rect 1607 998 1611 999
rect 1607 993 1611 994
rect 1639 998 1643 999
rect 1639 993 1643 994
rect 1711 998 1715 999
rect 1711 993 1715 994
rect 1719 998 1723 999
rect 1719 993 1723 994
rect 1807 998 1811 999
rect 1807 993 1811 994
rect 1823 998 1827 999
rect 1823 993 1827 994
rect 1903 998 1907 999
rect 1903 993 1907 994
rect 1935 998 1939 999
rect 1935 993 1939 994
rect 2015 998 2019 999
rect 2015 993 2019 994
rect 2047 998 2051 999
rect 2047 993 2051 994
rect 2143 998 2147 999
rect 2143 993 2147 994
rect 2151 998 2155 999
rect 2151 993 2155 994
rect 2255 998 2259 999
rect 2255 993 2259 994
rect 2271 998 2275 999
rect 2271 993 2275 994
rect 2351 998 2355 999
rect 2351 993 2355 994
rect 2407 998 2411 999
rect 2407 993 2411 994
rect 2447 998 2451 999
rect 2447 993 2451 994
rect 2527 998 2531 999
rect 2527 993 2531 994
rect 1526 991 1532 992
rect 1526 987 1527 991
rect 1531 987 1532 991
rect 1526 986 1532 987
rect 1558 983 1564 984
rect 1502 978 1508 979
rect 1510 981 1516 982
rect 1454 976 1460 977
rect 1470 954 1476 955
rect 1470 950 1471 954
rect 1475 950 1476 954
rect 1470 949 1476 950
rect 1430 947 1436 948
rect 1430 943 1431 947
rect 1435 943 1436 947
rect 1430 942 1436 943
rect 1446 947 1452 948
rect 1446 943 1447 947
rect 1451 943 1452 947
rect 1446 942 1452 943
rect 1367 934 1371 935
rect 1367 929 1371 930
rect 1415 934 1419 935
rect 1415 929 1419 930
rect 1326 925 1332 926
rect 1326 921 1327 925
rect 1331 921 1332 925
rect 1326 920 1332 921
rect 1368 914 1370 929
rect 1416 923 1418 929
rect 1414 922 1420 923
rect 1414 918 1415 922
rect 1419 918 1420 922
rect 1414 917 1420 918
rect 1366 913 1372 914
rect 1366 909 1367 913
rect 1371 909 1372 913
rect 1326 908 1332 909
rect 1366 908 1372 909
rect 798 907 804 908
rect 742 902 748 903
rect 778 903 784 904
rect 662 898 668 899
rect 688 891 690 902
rect 694 899 700 900
rect 694 895 695 899
rect 699 895 700 899
rect 694 894 700 895
rect 455 890 459 891
rect 455 885 459 886
rect 463 890 467 891
rect 463 885 467 886
rect 519 890 523 891
rect 519 885 523 886
rect 575 890 579 891
rect 575 885 579 886
rect 583 890 587 891
rect 583 885 587 886
rect 631 890 635 891
rect 631 885 635 886
rect 647 890 651 891
rect 647 885 651 886
rect 687 890 691 891
rect 687 885 691 886
rect 414 883 420 884
rect 414 879 415 883
rect 419 879 420 883
rect 414 878 420 879
rect 446 875 452 876
rect 382 870 388 871
rect 390 873 396 874
rect 334 868 340 869
rect 350 846 356 847
rect 350 842 351 846
rect 355 842 356 846
rect 350 841 356 842
rect 326 839 332 840
rect 326 835 327 839
rect 331 835 332 839
rect 326 834 332 835
rect 352 827 354 841
rect 384 840 386 870
rect 390 869 391 873
rect 395 869 396 873
rect 446 871 447 875
rect 451 871 452 875
rect 456 874 458 885
rect 510 875 516 876
rect 446 870 452 871
rect 454 873 460 874
rect 390 868 396 869
rect 406 846 412 847
rect 406 842 407 846
rect 411 842 412 846
rect 406 841 412 842
rect 382 839 388 840
rect 382 835 383 839
rect 387 835 388 839
rect 382 834 388 835
rect 408 827 410 841
rect 448 840 450 870
rect 454 869 455 873
rect 459 869 460 873
rect 510 871 511 875
rect 515 871 516 875
rect 520 874 522 885
rect 574 875 580 876
rect 510 870 516 871
rect 518 873 524 874
rect 454 868 460 869
rect 470 846 476 847
rect 470 842 471 846
rect 475 842 476 846
rect 470 841 476 842
rect 446 839 452 840
rect 446 835 447 839
rect 451 835 452 839
rect 446 834 452 835
rect 472 827 474 841
rect 512 840 514 870
rect 518 869 519 873
rect 523 869 524 873
rect 574 871 575 875
rect 579 871 580 875
rect 584 874 586 885
rect 648 874 650 885
rect 574 870 580 871
rect 582 873 588 874
rect 518 868 524 869
rect 534 846 540 847
rect 534 842 535 846
rect 539 842 540 846
rect 534 841 540 842
rect 510 839 516 840
rect 510 835 511 839
rect 515 835 516 839
rect 510 834 516 835
rect 536 827 538 841
rect 576 840 578 870
rect 582 869 583 873
rect 587 869 588 873
rect 582 868 588 869
rect 646 873 652 874
rect 646 869 647 873
rect 651 869 652 873
rect 646 868 652 869
rect 598 846 604 847
rect 598 842 599 846
rect 603 842 604 846
rect 598 841 604 842
rect 662 846 668 847
rect 662 842 663 846
rect 667 842 668 846
rect 662 841 668 842
rect 574 839 580 840
rect 574 835 575 839
rect 579 835 580 839
rect 574 834 580 835
rect 590 831 596 832
rect 590 827 591 831
rect 595 827 596 831
rect 600 827 602 841
rect 664 827 666 841
rect 696 840 698 894
rect 744 891 746 902
rect 778 899 779 903
rect 783 899 784 903
rect 798 903 799 907
rect 803 903 804 907
rect 1326 904 1327 908
rect 1331 904 1332 908
rect 1326 903 1332 904
rect 798 902 804 903
rect 778 898 784 899
rect 800 891 802 902
rect 1328 891 1330 903
rect 1366 896 1372 897
rect 1366 892 1367 896
rect 1371 892 1372 896
rect 1366 891 1372 892
rect 1398 895 1404 896
rect 1398 891 1399 895
rect 1403 891 1404 895
rect 1432 892 1434 942
rect 1472 935 1474 949
rect 1504 948 1506 978
rect 1510 977 1511 981
rect 1515 977 1516 981
rect 1558 979 1559 983
rect 1563 979 1564 983
rect 1568 982 1570 993
rect 1630 983 1636 984
rect 1558 978 1564 979
rect 1566 981 1572 982
rect 1510 976 1516 977
rect 1526 954 1532 955
rect 1526 950 1527 954
rect 1531 950 1532 954
rect 1526 949 1532 950
rect 1502 947 1508 948
rect 1502 943 1503 947
rect 1507 943 1508 947
rect 1502 942 1508 943
rect 1486 935 1492 936
rect 1528 935 1530 949
rect 1560 948 1562 978
rect 1566 977 1567 981
rect 1571 977 1572 981
rect 1630 979 1631 983
rect 1635 979 1636 983
rect 1640 982 1642 993
rect 1710 983 1716 984
rect 1630 978 1636 979
rect 1638 981 1644 982
rect 1566 976 1572 977
rect 1582 954 1588 955
rect 1582 950 1583 954
rect 1587 950 1588 954
rect 1582 949 1588 950
rect 1558 947 1564 948
rect 1558 943 1559 947
rect 1563 943 1564 947
rect 1558 942 1564 943
rect 1584 935 1586 949
rect 1632 948 1634 978
rect 1638 977 1639 981
rect 1643 977 1644 981
rect 1710 979 1711 983
rect 1715 979 1716 983
rect 1720 982 1722 993
rect 1808 982 1810 993
rect 1894 983 1900 984
rect 1710 978 1716 979
rect 1718 981 1724 982
rect 1638 976 1644 977
rect 1654 954 1660 955
rect 1654 950 1655 954
rect 1659 950 1660 954
rect 1654 949 1660 950
rect 1630 947 1636 948
rect 1630 943 1631 947
rect 1635 943 1636 947
rect 1630 942 1636 943
rect 1630 935 1636 936
rect 1656 935 1658 949
rect 1712 948 1714 978
rect 1718 977 1719 981
rect 1723 977 1724 981
rect 1718 976 1724 977
rect 1806 981 1812 982
rect 1806 977 1807 981
rect 1811 977 1812 981
rect 1894 979 1895 983
rect 1899 979 1900 983
rect 1904 982 1906 993
rect 2006 983 2012 984
rect 1894 978 1900 979
rect 1902 981 1908 982
rect 1806 976 1812 977
rect 1734 954 1740 955
rect 1734 950 1735 954
rect 1739 950 1740 954
rect 1734 949 1740 950
rect 1822 954 1828 955
rect 1822 950 1823 954
rect 1827 950 1828 954
rect 1822 949 1828 950
rect 1710 947 1716 948
rect 1710 943 1711 947
rect 1715 943 1716 947
rect 1710 942 1716 943
rect 1736 935 1738 949
rect 1824 935 1826 949
rect 1896 948 1898 978
rect 1902 977 1903 981
rect 1907 977 1908 981
rect 2006 979 2007 983
rect 2011 979 2012 983
rect 2016 982 2018 993
rect 2134 983 2140 984
rect 2006 978 2012 979
rect 2014 981 2020 982
rect 1902 976 1908 977
rect 1918 954 1924 955
rect 1918 950 1919 954
rect 1923 950 1924 954
rect 1918 949 1924 950
rect 1894 947 1900 948
rect 1894 943 1895 947
rect 1899 943 1900 947
rect 1894 942 1900 943
rect 1920 935 1922 949
rect 2008 948 2010 978
rect 2014 977 2015 981
rect 2019 977 2020 981
rect 2134 979 2135 983
rect 2139 979 2140 983
rect 2144 982 2146 993
rect 2262 983 2268 984
rect 2134 978 2140 979
rect 2142 981 2148 982
rect 2014 976 2020 977
rect 2030 954 2036 955
rect 2030 950 2031 954
rect 2035 950 2036 954
rect 2030 949 2036 950
rect 2006 947 2012 948
rect 2006 943 2007 947
rect 2011 943 2012 947
rect 2006 942 2012 943
rect 2032 935 2034 949
rect 2136 948 2138 978
rect 2142 977 2143 981
rect 2147 977 2148 981
rect 2262 979 2263 983
rect 2267 979 2268 983
rect 2272 982 2274 993
rect 2294 983 2300 984
rect 2262 978 2268 979
rect 2270 981 2276 982
rect 2142 976 2148 977
rect 2158 954 2164 955
rect 2158 950 2159 954
rect 2163 950 2164 954
rect 2158 949 2164 950
rect 2134 947 2140 948
rect 2134 943 2135 947
rect 2139 943 2140 947
rect 2134 942 2140 943
rect 2078 935 2084 936
rect 2160 935 2162 949
rect 2264 948 2266 978
rect 2270 977 2271 981
rect 2275 977 2276 981
rect 2294 979 2295 983
rect 2299 979 2300 983
rect 2408 982 2410 993
rect 2518 983 2524 984
rect 2294 978 2300 979
rect 2406 981 2412 982
rect 2270 976 2276 977
rect 2286 954 2292 955
rect 2286 950 2287 954
rect 2291 950 2292 954
rect 2286 949 2292 950
rect 2262 947 2268 948
rect 2262 943 2263 947
rect 2267 943 2268 947
rect 2262 942 2268 943
rect 2288 935 2290 949
rect 2296 936 2298 978
rect 2406 977 2407 981
rect 2411 977 2412 981
rect 2518 979 2519 983
rect 2523 979 2524 983
rect 2528 982 2530 993
rect 2536 988 2538 1058
rect 2542 1054 2543 1058
rect 2547 1054 2548 1058
rect 2542 1053 2548 1054
rect 2584 1050 2586 1065
rect 2582 1049 2588 1050
rect 2582 1045 2583 1049
rect 2587 1045 2588 1049
rect 2582 1044 2588 1045
rect 2582 1032 2588 1033
rect 2582 1028 2583 1032
rect 2587 1028 2588 1032
rect 2582 1027 2588 1028
rect 2584 999 2586 1027
rect 2583 998 2587 999
rect 2583 993 2587 994
rect 2534 987 2540 988
rect 2534 983 2535 987
rect 2539 983 2540 987
rect 2534 982 2540 983
rect 2518 978 2524 979
rect 2526 981 2532 982
rect 2584 981 2586 993
rect 2406 976 2412 977
rect 2422 954 2428 955
rect 2422 950 2423 954
rect 2427 950 2428 954
rect 2422 949 2428 950
rect 2330 947 2336 948
rect 2330 943 2331 947
rect 2335 943 2336 947
rect 2330 942 2336 943
rect 2294 935 2300 936
rect 1471 934 1475 935
rect 1486 931 1487 935
rect 1491 931 1492 935
rect 1486 930 1492 931
rect 1527 934 1531 935
rect 1471 929 1475 930
rect 1446 927 1452 928
rect 1446 923 1447 927
rect 1451 923 1452 927
rect 1472 923 1474 929
rect 1446 922 1452 923
rect 1470 922 1476 923
rect 1448 904 1450 922
rect 1470 918 1471 922
rect 1475 918 1476 922
rect 1470 917 1476 918
rect 1446 903 1452 904
rect 1446 899 1447 903
rect 1451 899 1452 903
rect 1446 898 1452 899
rect 1454 895 1460 896
rect 711 890 715 891
rect 711 885 715 886
rect 743 890 747 891
rect 743 885 747 886
rect 775 890 779 891
rect 775 885 779 886
rect 799 890 803 891
rect 799 885 803 886
rect 847 890 851 891
rect 847 885 851 886
rect 919 890 923 891
rect 919 885 923 886
rect 1327 890 1331 891
rect 1327 885 1331 886
rect 702 875 708 876
rect 702 871 703 875
rect 707 871 708 875
rect 712 874 714 885
rect 766 875 772 876
rect 702 870 708 871
rect 710 873 716 874
rect 704 840 706 870
rect 710 869 711 873
rect 715 869 716 873
rect 766 871 767 875
rect 771 871 772 875
rect 776 874 778 885
rect 838 875 844 876
rect 766 870 772 871
rect 774 873 780 874
rect 710 868 716 869
rect 726 846 732 847
rect 726 842 727 846
rect 731 842 732 846
rect 726 841 732 842
rect 694 839 700 840
rect 694 835 695 839
rect 699 835 700 839
rect 694 834 700 835
rect 702 839 708 840
rect 702 835 703 839
rect 707 835 708 839
rect 702 834 708 835
rect 728 827 730 841
rect 768 840 770 870
rect 774 869 775 873
rect 779 869 780 873
rect 838 871 839 875
rect 843 871 844 875
rect 848 874 850 885
rect 910 875 916 876
rect 838 870 844 871
rect 846 873 852 874
rect 774 868 780 869
rect 790 846 796 847
rect 790 842 791 846
rect 795 842 796 846
rect 790 841 796 842
rect 766 839 772 840
rect 766 835 767 839
rect 771 835 772 839
rect 766 834 772 835
rect 792 827 794 841
rect 840 840 842 870
rect 846 869 847 873
rect 851 869 852 873
rect 910 871 911 875
rect 915 871 916 875
rect 920 874 922 885
rect 942 875 948 876
rect 910 870 916 871
rect 918 873 924 874
rect 846 868 852 869
rect 862 846 868 847
rect 862 842 863 846
rect 867 842 868 846
rect 862 841 868 842
rect 838 839 844 840
rect 838 835 839 839
rect 843 835 844 839
rect 838 834 844 835
rect 864 827 866 841
rect 912 840 914 870
rect 918 869 919 873
rect 923 869 924 873
rect 942 871 943 875
rect 947 871 948 875
rect 1328 873 1330 885
rect 1368 879 1370 891
rect 1398 890 1404 891
rect 1430 891 1436 892
rect 1400 879 1402 890
rect 1430 887 1431 891
rect 1435 887 1436 891
rect 1454 891 1455 895
rect 1459 891 1460 895
rect 1488 892 1490 930
rect 1527 929 1531 930
rect 1583 934 1587 935
rect 1583 929 1587 930
rect 1615 934 1619 935
rect 1630 931 1631 935
rect 1635 931 1636 935
rect 1630 930 1636 931
rect 1655 934 1659 935
rect 1615 929 1619 930
rect 1528 923 1530 929
rect 1590 927 1596 928
rect 1590 923 1591 927
rect 1595 923 1596 927
rect 1616 923 1618 929
rect 1526 922 1532 923
rect 1590 922 1596 923
rect 1614 922 1620 923
rect 1526 918 1527 922
rect 1531 918 1532 922
rect 1526 917 1532 918
rect 1592 904 1594 922
rect 1614 918 1615 922
rect 1619 918 1620 922
rect 1614 917 1620 918
rect 1590 903 1596 904
rect 1590 899 1591 903
rect 1595 899 1596 903
rect 1590 898 1596 899
rect 1510 895 1516 896
rect 1454 890 1460 891
rect 1486 891 1492 892
rect 1430 886 1436 887
rect 1456 879 1458 890
rect 1486 887 1487 891
rect 1491 887 1492 891
rect 1510 891 1511 895
rect 1515 891 1516 895
rect 1510 890 1516 891
rect 1598 895 1604 896
rect 1598 891 1599 895
rect 1603 891 1604 895
rect 1632 892 1634 930
rect 1655 929 1659 930
rect 1711 934 1715 935
rect 1711 929 1715 930
rect 1735 934 1739 935
rect 1735 929 1739 930
rect 1823 934 1827 935
rect 1823 929 1827 930
rect 1919 934 1923 935
rect 1919 929 1923 930
rect 1943 934 1947 935
rect 1943 929 1947 930
rect 2031 934 2035 935
rect 2031 929 2035 930
rect 2063 934 2067 935
rect 2078 931 2079 935
rect 2083 931 2084 935
rect 2078 930 2084 931
rect 2159 934 2163 935
rect 2063 929 2067 930
rect 1712 923 1714 929
rect 1824 923 1826 929
rect 1944 923 1946 929
rect 2038 927 2044 928
rect 2038 923 2039 927
rect 2043 923 2044 927
rect 2064 923 2066 929
rect 1710 922 1716 923
rect 1710 918 1711 922
rect 1715 918 1716 922
rect 1710 917 1716 918
rect 1822 922 1828 923
rect 1822 918 1823 922
rect 1827 918 1828 922
rect 1822 917 1828 918
rect 1942 922 1948 923
rect 2038 922 2044 923
rect 2062 922 2068 923
rect 1942 918 1943 922
rect 1947 918 1948 922
rect 1942 917 1948 918
rect 2040 904 2042 922
rect 2062 918 2063 922
rect 2067 918 2068 922
rect 2062 917 2068 918
rect 2038 903 2044 904
rect 2038 899 2039 903
rect 2043 899 2044 903
rect 2038 898 2044 899
rect 1694 895 1700 896
rect 1598 890 1604 891
rect 1630 891 1636 892
rect 1486 886 1492 887
rect 1512 879 1514 890
rect 1600 879 1602 890
rect 1630 887 1631 891
rect 1635 887 1636 891
rect 1694 891 1695 895
rect 1699 891 1700 895
rect 1694 890 1700 891
rect 1806 895 1812 896
rect 1806 891 1807 895
rect 1811 891 1812 895
rect 1806 890 1812 891
rect 1926 895 1932 896
rect 1926 891 1927 895
rect 1931 891 1932 895
rect 2046 895 2052 896
rect 1926 890 1932 891
rect 1950 891 1956 892
rect 1630 886 1636 887
rect 1696 879 1698 890
rect 1808 879 1810 890
rect 1928 879 1930 890
rect 1950 887 1951 891
rect 1955 887 1956 891
rect 2046 891 2047 895
rect 2051 891 2052 895
rect 2080 892 2082 930
rect 2159 929 2163 930
rect 2183 934 2187 935
rect 2183 929 2187 930
rect 2287 934 2291 935
rect 2294 931 2295 935
rect 2299 931 2300 935
rect 2294 930 2300 931
rect 2311 934 2315 935
rect 2287 929 2291 930
rect 2311 929 2315 930
rect 2184 923 2186 929
rect 2312 923 2314 929
rect 2182 922 2188 923
rect 2182 918 2183 922
rect 2187 918 2188 922
rect 2182 917 2188 918
rect 2310 922 2316 923
rect 2310 918 2311 922
rect 2315 918 2316 922
rect 2310 917 2316 918
rect 2166 895 2172 896
rect 2046 890 2052 891
rect 2078 891 2084 892
rect 1950 886 1956 887
rect 1367 878 1371 879
rect 1367 873 1371 874
rect 1399 878 1403 879
rect 1399 873 1403 874
rect 1455 878 1459 879
rect 1455 873 1459 874
rect 1471 878 1475 879
rect 1471 873 1475 874
rect 1511 878 1515 879
rect 1511 873 1515 874
rect 1551 878 1555 879
rect 1551 873 1555 874
rect 1599 878 1603 879
rect 1599 873 1603 874
rect 1639 878 1643 879
rect 1639 873 1643 874
rect 1695 878 1699 879
rect 1695 873 1699 874
rect 1727 878 1731 879
rect 1727 873 1731 874
rect 1807 878 1811 879
rect 1807 873 1811 874
rect 1815 878 1819 879
rect 1815 873 1819 874
rect 1903 878 1907 879
rect 1903 873 1907 874
rect 1927 878 1931 879
rect 1927 873 1931 874
rect 942 870 948 871
rect 1326 872 1332 873
rect 918 868 924 869
rect 934 846 940 847
rect 934 842 935 846
rect 939 842 940 846
rect 934 841 940 842
rect 910 839 916 840
rect 910 835 911 839
rect 915 835 916 839
rect 910 834 916 835
rect 936 827 938 841
rect 944 828 946 870
rect 1326 868 1327 872
rect 1331 868 1332 872
rect 1326 867 1332 868
rect 1368 861 1370 873
rect 1472 862 1474 873
rect 1542 863 1548 864
rect 1470 861 1476 862
rect 1366 860 1372 861
rect 1366 856 1367 860
rect 1371 856 1372 860
rect 1470 857 1471 861
rect 1475 857 1476 861
rect 1542 859 1543 863
rect 1547 859 1548 863
rect 1552 862 1554 873
rect 1630 863 1636 864
rect 1542 858 1548 859
rect 1550 861 1556 862
rect 1470 856 1476 857
rect 1326 855 1332 856
rect 1366 855 1372 856
rect 1326 851 1327 855
rect 1331 851 1332 855
rect 1326 850 1332 851
rect 942 827 948 828
rect 1328 827 1330 850
rect 1366 843 1372 844
rect 1366 839 1367 843
rect 1371 839 1372 843
rect 1366 838 1372 839
rect 111 826 115 827
rect 111 821 115 822
rect 167 826 171 827
rect 167 821 171 822
rect 231 826 235 827
rect 231 821 235 822
rect 295 826 299 827
rect 295 821 299 822
rect 311 826 315 827
rect 311 821 315 822
rect 351 826 355 827
rect 351 821 355 822
rect 399 826 403 827
rect 399 821 403 822
rect 407 826 411 827
rect 407 821 411 822
rect 471 826 475 827
rect 471 821 475 822
rect 487 826 491 827
rect 487 821 491 822
rect 535 826 539 827
rect 535 821 539 822
rect 583 826 587 827
rect 590 826 596 827
rect 599 826 603 827
rect 583 821 587 822
rect 112 806 114 821
rect 158 819 164 820
rect 158 815 159 819
rect 163 815 164 819
rect 168 815 170 821
rect 186 819 192 820
rect 186 815 187 819
rect 191 815 192 819
rect 232 815 234 821
rect 250 819 256 820
rect 250 815 251 819
rect 255 815 256 819
rect 312 815 314 821
rect 330 819 336 820
rect 330 815 331 819
rect 335 815 336 819
rect 400 815 402 821
rect 418 819 424 820
rect 418 815 419 819
rect 423 815 424 819
rect 488 815 490 821
rect 506 819 512 820
rect 506 815 507 819
rect 511 815 512 819
rect 584 815 586 821
rect 158 814 164 815
rect 166 814 172 815
rect 186 814 192 815
rect 230 814 236 815
rect 250 814 256 815
rect 310 814 316 815
rect 330 814 336 815
rect 398 814 404 815
rect 418 814 424 815
rect 486 814 492 815
rect 506 814 512 815
rect 582 814 588 815
rect 110 805 116 806
rect 110 801 111 805
rect 115 801 116 805
rect 110 800 116 801
rect 110 788 116 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 150 787 156 788
rect 150 783 151 787
rect 155 783 156 787
rect 112 763 114 783
rect 150 782 156 783
rect 152 763 154 782
rect 111 762 115 763
rect 111 757 115 758
rect 143 762 147 763
rect 143 757 147 758
rect 151 762 155 763
rect 151 757 155 758
rect 112 745 114 757
rect 144 746 146 757
rect 160 756 162 814
rect 166 810 167 814
rect 171 810 172 814
rect 166 809 172 810
rect 188 784 190 814
rect 230 810 231 814
rect 235 810 236 814
rect 230 809 236 810
rect 214 787 220 788
rect 186 783 192 784
rect 186 779 187 783
rect 191 779 192 783
rect 214 783 215 787
rect 219 783 220 787
rect 252 784 254 814
rect 310 810 311 814
rect 315 810 316 814
rect 310 809 316 810
rect 294 787 300 788
rect 214 782 220 783
rect 250 783 256 784
rect 186 778 192 779
rect 216 763 218 782
rect 250 779 251 783
rect 255 779 256 783
rect 294 783 295 787
rect 299 783 300 787
rect 332 784 334 814
rect 398 810 399 814
rect 403 810 404 814
rect 398 809 404 810
rect 382 787 388 788
rect 294 782 300 783
rect 330 783 336 784
rect 250 778 256 779
rect 296 763 298 782
rect 330 779 331 783
rect 335 779 336 783
rect 382 783 383 787
rect 387 783 388 787
rect 420 784 422 814
rect 486 810 487 814
rect 491 810 492 814
rect 486 809 492 810
rect 470 787 476 788
rect 382 782 388 783
rect 418 783 424 784
rect 330 778 336 779
rect 384 763 386 782
rect 418 779 419 783
rect 423 779 424 783
rect 470 783 471 787
rect 475 783 476 787
rect 508 784 510 814
rect 582 810 583 814
rect 587 810 588 814
rect 582 809 588 810
rect 566 787 572 788
rect 470 782 476 783
rect 506 783 512 784
rect 418 778 424 779
rect 472 763 474 782
rect 506 779 507 783
rect 511 779 512 783
rect 566 783 567 787
rect 571 783 572 787
rect 592 784 594 826
rect 599 821 603 822
rect 663 826 667 827
rect 663 821 667 822
rect 671 826 675 827
rect 671 821 675 822
rect 727 826 731 827
rect 727 821 731 822
rect 759 826 763 827
rect 759 821 763 822
rect 791 826 795 827
rect 791 821 795 822
rect 839 826 843 827
rect 839 821 843 822
rect 863 826 867 827
rect 863 821 867 822
rect 919 826 923 827
rect 919 821 923 822
rect 935 826 939 827
rect 942 823 943 827
rect 947 823 948 827
rect 942 822 948 823
rect 1007 826 1011 827
rect 935 821 939 822
rect 1007 821 1011 822
rect 1095 826 1099 827
rect 1095 821 1099 822
rect 1327 826 1331 827
rect 1327 821 1331 822
rect 672 815 674 821
rect 690 819 696 820
rect 690 815 691 819
rect 695 815 696 819
rect 760 815 762 821
rect 778 819 784 820
rect 778 815 779 819
rect 783 815 784 819
rect 840 815 842 821
rect 920 815 922 821
rect 1008 815 1010 821
rect 1026 819 1032 820
rect 1026 815 1027 819
rect 1031 815 1032 819
rect 1096 815 1098 821
rect 670 814 676 815
rect 690 814 696 815
rect 758 814 764 815
rect 778 814 784 815
rect 838 814 844 815
rect 670 810 671 814
rect 675 810 676 814
rect 670 809 676 810
rect 654 787 660 788
rect 566 782 572 783
rect 590 783 596 784
rect 506 778 512 779
rect 568 763 570 782
rect 590 779 591 783
rect 595 779 596 783
rect 654 783 655 787
rect 659 783 660 787
rect 692 784 694 814
rect 758 810 759 814
rect 763 810 764 814
rect 758 809 764 810
rect 742 787 748 788
rect 654 782 660 783
rect 690 783 696 784
rect 590 778 596 779
rect 656 763 658 782
rect 690 779 691 783
rect 695 779 696 783
rect 742 783 743 787
rect 747 783 748 787
rect 780 784 782 814
rect 838 810 839 814
rect 843 810 844 814
rect 838 809 844 810
rect 918 814 924 815
rect 918 810 919 814
rect 923 810 924 814
rect 918 809 924 810
rect 1006 814 1012 815
rect 1026 814 1032 815
rect 1094 814 1100 815
rect 1006 810 1007 814
rect 1011 810 1012 814
rect 1006 809 1012 810
rect 822 787 828 788
rect 742 782 748 783
rect 778 783 784 784
rect 690 778 696 779
rect 744 763 746 782
rect 778 779 779 783
rect 783 779 784 783
rect 822 783 823 787
rect 827 783 828 787
rect 822 782 828 783
rect 902 787 908 788
rect 902 783 903 787
rect 907 783 908 787
rect 902 782 908 783
rect 990 787 996 788
rect 990 783 991 787
rect 995 783 996 787
rect 1028 784 1030 814
rect 1094 810 1095 814
rect 1099 810 1100 814
rect 1094 809 1100 810
rect 1328 806 1330 821
rect 1368 815 1370 838
rect 1486 834 1492 835
rect 1486 830 1487 834
rect 1491 830 1492 834
rect 1486 829 1492 830
rect 1488 815 1490 829
rect 1544 828 1546 858
rect 1550 857 1551 861
rect 1555 857 1556 861
rect 1630 859 1631 863
rect 1635 859 1636 863
rect 1640 862 1642 873
rect 1728 862 1730 873
rect 1750 871 1756 872
rect 1750 867 1751 871
rect 1755 867 1756 871
rect 1750 866 1756 867
rect 1630 858 1636 859
rect 1638 861 1644 862
rect 1550 856 1556 857
rect 1566 834 1572 835
rect 1566 830 1567 834
rect 1571 830 1572 834
rect 1566 829 1572 830
rect 1542 827 1548 828
rect 1542 823 1543 827
rect 1547 823 1548 827
rect 1542 822 1548 823
rect 1568 815 1570 829
rect 1632 828 1634 858
rect 1638 857 1639 861
rect 1643 857 1644 861
rect 1638 856 1644 857
rect 1726 861 1732 862
rect 1726 857 1727 861
rect 1731 857 1732 861
rect 1726 856 1732 857
rect 1654 834 1660 835
rect 1654 830 1655 834
rect 1659 830 1660 834
rect 1654 829 1660 830
rect 1742 834 1748 835
rect 1742 830 1743 834
rect 1747 830 1748 834
rect 1742 829 1748 830
rect 1630 827 1636 828
rect 1630 823 1631 827
rect 1635 823 1636 827
rect 1630 822 1636 823
rect 1656 815 1658 829
rect 1744 815 1746 829
rect 1752 828 1754 866
rect 1758 863 1764 864
rect 1758 859 1759 863
rect 1763 859 1764 863
rect 1816 862 1818 873
rect 1904 862 1906 873
rect 1758 858 1764 859
rect 1814 861 1820 862
rect 1750 827 1756 828
rect 1750 823 1751 827
rect 1755 823 1756 827
rect 1760 824 1762 858
rect 1814 857 1815 861
rect 1819 857 1820 861
rect 1814 856 1820 857
rect 1902 861 1908 862
rect 1902 857 1903 861
rect 1907 857 1908 861
rect 1902 856 1908 857
rect 1830 834 1836 835
rect 1830 830 1831 834
rect 1835 830 1836 834
rect 1830 829 1836 830
rect 1918 834 1924 835
rect 1918 830 1919 834
rect 1923 830 1924 834
rect 1918 829 1924 830
rect 1770 827 1776 828
rect 1750 822 1756 823
rect 1758 823 1764 824
rect 1758 819 1759 823
rect 1763 819 1764 823
rect 1770 823 1771 827
rect 1775 823 1776 827
rect 1770 822 1776 823
rect 1758 818 1764 819
rect 1367 814 1371 815
rect 1367 809 1371 810
rect 1487 814 1491 815
rect 1487 809 1491 810
rect 1567 814 1571 815
rect 1567 809 1571 810
rect 1631 814 1635 815
rect 1631 809 1635 810
rect 1655 814 1659 815
rect 1655 809 1659 810
rect 1687 814 1691 815
rect 1687 809 1691 810
rect 1743 814 1747 815
rect 1743 809 1747 810
rect 1751 814 1755 815
rect 1751 809 1755 810
rect 1326 805 1332 806
rect 1326 801 1327 805
rect 1331 801 1332 805
rect 1326 800 1332 801
rect 1368 794 1370 809
rect 1632 803 1634 809
rect 1688 803 1690 809
rect 1706 807 1712 808
rect 1706 803 1707 807
rect 1711 803 1712 807
rect 1752 803 1754 809
rect 1630 802 1636 803
rect 1630 798 1631 802
rect 1635 798 1636 802
rect 1630 797 1636 798
rect 1686 802 1692 803
rect 1706 802 1712 803
rect 1750 802 1756 803
rect 1686 798 1687 802
rect 1691 798 1692 802
rect 1686 797 1692 798
rect 1366 793 1372 794
rect 1366 789 1367 793
rect 1371 789 1372 793
rect 1326 788 1332 789
rect 1366 788 1372 789
rect 1078 787 1084 788
rect 990 782 996 783
rect 1026 783 1032 784
rect 778 778 784 779
rect 824 763 826 782
rect 904 763 906 782
rect 992 763 994 782
rect 1026 779 1027 783
rect 1031 779 1032 783
rect 1078 783 1079 787
rect 1083 783 1084 787
rect 1326 784 1327 788
rect 1331 784 1332 788
rect 1078 782 1084 783
rect 1102 783 1108 784
rect 1326 783 1332 784
rect 1026 778 1032 779
rect 1080 763 1082 782
rect 1102 779 1103 783
rect 1107 779 1108 783
rect 1102 778 1108 779
rect 199 762 203 763
rect 199 757 203 758
rect 215 762 219 763
rect 215 757 219 758
rect 279 762 283 763
rect 279 757 283 758
rect 295 762 299 763
rect 295 757 299 758
rect 383 762 387 763
rect 383 757 387 758
rect 471 762 475 763
rect 471 757 475 758
rect 487 762 491 763
rect 487 757 491 758
rect 567 762 571 763
rect 567 757 571 758
rect 599 762 603 763
rect 599 757 603 758
rect 655 762 659 763
rect 655 757 659 758
rect 703 762 707 763
rect 703 757 707 758
rect 743 762 747 763
rect 743 757 747 758
rect 807 762 811 763
rect 807 757 811 758
rect 823 762 827 763
rect 823 757 827 758
rect 903 762 907 763
rect 903 757 907 758
rect 991 762 995 763
rect 991 757 995 758
rect 1079 762 1083 763
rect 1079 757 1083 758
rect 158 755 164 756
rect 158 751 159 755
rect 163 751 164 755
rect 158 750 164 751
rect 190 747 196 748
rect 142 745 148 746
rect 110 744 116 745
rect 110 740 111 744
rect 115 740 116 744
rect 142 741 143 745
rect 147 741 148 745
rect 190 743 191 747
rect 195 743 196 747
rect 200 746 202 757
rect 270 747 276 748
rect 190 742 196 743
rect 198 745 204 746
rect 142 740 148 741
rect 110 739 116 740
rect 110 727 116 728
rect 110 723 111 727
rect 115 723 116 727
rect 110 722 116 723
rect 112 703 114 722
rect 158 718 164 719
rect 158 714 159 718
rect 163 714 164 718
rect 158 713 164 714
rect 160 703 162 713
rect 192 712 194 742
rect 198 741 199 745
rect 203 741 204 745
rect 270 743 271 747
rect 275 743 276 747
rect 280 746 282 757
rect 374 747 380 748
rect 270 742 276 743
rect 278 745 284 746
rect 198 740 204 741
rect 214 718 220 719
rect 214 714 215 718
rect 219 714 220 718
rect 214 713 220 714
rect 190 711 196 712
rect 190 707 191 711
rect 195 707 196 711
rect 190 706 196 707
rect 216 703 218 713
rect 272 712 274 742
rect 278 741 279 745
rect 283 741 284 745
rect 374 743 375 747
rect 379 743 380 747
rect 384 746 386 757
rect 478 747 484 748
rect 374 742 380 743
rect 382 745 388 746
rect 278 740 284 741
rect 294 718 300 719
rect 294 714 295 718
rect 299 714 300 718
rect 294 713 300 714
rect 270 711 276 712
rect 270 707 271 711
rect 275 707 276 711
rect 270 706 276 707
rect 296 703 298 713
rect 376 712 378 742
rect 382 741 383 745
rect 387 741 388 745
rect 478 743 479 747
rect 483 743 484 747
rect 488 746 490 757
rect 590 747 596 748
rect 478 742 484 743
rect 486 745 492 746
rect 382 740 388 741
rect 398 718 404 719
rect 398 714 399 718
rect 403 714 404 718
rect 398 713 404 714
rect 374 711 380 712
rect 374 707 375 711
rect 379 707 380 711
rect 374 706 380 707
rect 366 703 372 704
rect 400 703 402 713
rect 480 712 482 742
rect 486 741 487 745
rect 491 741 492 745
rect 590 743 591 747
rect 595 743 596 747
rect 600 746 602 757
rect 704 746 706 757
rect 798 747 804 748
rect 590 742 596 743
rect 598 745 604 746
rect 486 740 492 741
rect 502 718 508 719
rect 502 714 503 718
rect 507 714 508 718
rect 502 713 508 714
rect 478 711 484 712
rect 478 707 479 711
rect 483 707 484 711
rect 478 706 484 707
rect 504 703 506 713
rect 592 712 594 742
rect 598 741 599 745
rect 603 741 604 745
rect 598 740 604 741
rect 702 745 708 746
rect 702 741 703 745
rect 707 741 708 745
rect 798 743 799 747
rect 803 743 804 747
rect 808 746 810 757
rect 894 747 900 748
rect 798 742 804 743
rect 806 745 812 746
rect 702 740 708 741
rect 614 718 620 719
rect 614 714 615 718
rect 619 714 620 718
rect 718 718 724 719
rect 614 713 620 714
rect 699 716 703 717
rect 590 711 596 712
rect 590 707 591 711
rect 595 707 596 711
rect 590 706 596 707
rect 616 703 618 713
rect 718 714 719 718
rect 723 714 724 718
rect 718 713 724 714
rect 698 711 704 712
rect 698 707 699 711
rect 703 707 704 711
rect 698 706 704 707
rect 720 703 722 713
rect 800 712 802 742
rect 806 741 807 745
rect 811 741 812 745
rect 894 743 895 747
rect 899 743 900 747
rect 904 746 906 757
rect 982 747 988 748
rect 894 742 900 743
rect 902 745 908 746
rect 806 740 812 741
rect 822 718 828 719
rect 822 714 823 718
rect 827 714 828 718
rect 822 713 828 714
rect 798 711 804 712
rect 798 707 799 711
rect 803 707 804 711
rect 798 706 804 707
rect 726 703 732 704
rect 824 703 826 713
rect 896 712 898 742
rect 902 741 903 745
rect 907 741 908 745
rect 982 743 983 747
rect 987 743 988 747
rect 992 746 994 757
rect 1070 747 1076 748
rect 982 742 988 743
rect 990 745 996 746
rect 902 740 908 741
rect 918 718 924 719
rect 918 714 919 718
rect 923 714 924 718
rect 918 713 924 714
rect 894 711 900 712
rect 894 707 895 711
rect 899 707 900 711
rect 894 706 900 707
rect 886 703 892 704
rect 920 703 922 713
rect 984 712 986 742
rect 990 741 991 745
rect 995 741 996 745
rect 1070 743 1071 747
rect 1075 743 1076 747
rect 1080 746 1082 757
rect 1070 742 1076 743
rect 1078 745 1084 746
rect 990 740 996 741
rect 1006 718 1012 719
rect 1006 714 1007 718
rect 1011 714 1012 718
rect 1006 713 1012 714
rect 982 711 988 712
rect 982 707 983 711
rect 987 707 988 711
rect 982 706 988 707
rect 1008 703 1010 713
rect 1072 712 1074 742
rect 1078 741 1079 745
rect 1083 741 1084 745
rect 1078 740 1084 741
rect 1094 718 1100 719
rect 1094 714 1095 718
rect 1099 714 1100 718
rect 1104 717 1106 778
rect 1328 763 1330 783
rect 1366 776 1372 777
rect 1366 772 1367 776
rect 1371 772 1372 776
rect 1366 771 1372 772
rect 1614 775 1620 776
rect 1614 771 1615 775
rect 1619 771 1620 775
rect 1175 762 1179 763
rect 1175 757 1179 758
rect 1327 762 1331 763
rect 1327 757 1331 758
rect 1166 747 1172 748
rect 1166 743 1167 747
rect 1171 743 1172 747
rect 1176 746 1178 757
rect 1198 747 1204 748
rect 1166 742 1172 743
rect 1174 745 1180 746
rect 1094 713 1100 714
rect 1103 716 1107 717
rect 1070 711 1076 712
rect 1070 707 1071 711
rect 1075 707 1076 711
rect 1070 706 1076 707
rect 1096 703 1098 713
rect 1168 712 1170 742
rect 1174 741 1175 745
rect 1179 741 1180 745
rect 1198 743 1199 747
rect 1203 743 1204 747
rect 1328 745 1330 757
rect 1368 755 1370 771
rect 1614 770 1620 771
rect 1670 775 1676 776
rect 1670 771 1671 775
rect 1675 771 1676 775
rect 1708 772 1710 802
rect 1750 798 1751 802
rect 1755 798 1756 802
rect 1750 797 1756 798
rect 1734 775 1740 776
rect 1670 770 1676 771
rect 1706 771 1712 772
rect 1616 755 1618 770
rect 1672 755 1674 770
rect 1706 767 1707 771
rect 1711 767 1712 771
rect 1734 771 1735 775
rect 1739 771 1740 775
rect 1772 772 1774 822
rect 1832 815 1834 829
rect 1838 815 1844 816
rect 1920 815 1922 829
rect 1952 828 1954 886
rect 2048 879 2050 890
rect 2078 887 2079 891
rect 2083 887 2084 891
rect 2166 891 2167 895
rect 2171 891 2172 895
rect 2166 890 2172 891
rect 2294 895 2300 896
rect 2294 891 2295 895
rect 2299 891 2300 895
rect 2332 892 2334 942
rect 2424 935 2426 949
rect 2520 948 2522 978
rect 2526 977 2527 981
rect 2531 977 2532 981
rect 2526 976 2532 977
rect 2582 980 2588 981
rect 2582 976 2583 980
rect 2587 976 2588 980
rect 2582 975 2588 976
rect 2582 963 2588 964
rect 2582 959 2583 963
rect 2587 959 2588 963
rect 2582 958 2588 959
rect 2542 954 2548 955
rect 2542 950 2543 954
rect 2547 950 2548 954
rect 2542 949 2548 950
rect 2518 947 2524 948
rect 2518 943 2519 947
rect 2523 943 2524 947
rect 2518 942 2524 943
rect 2454 935 2460 936
rect 2544 935 2546 949
rect 2584 935 2586 958
rect 2423 934 2427 935
rect 2423 929 2427 930
rect 2439 934 2443 935
rect 2454 931 2455 935
rect 2459 931 2460 935
rect 2454 930 2460 931
rect 2543 934 2547 935
rect 2439 929 2443 930
rect 2414 927 2420 928
rect 2414 923 2415 927
rect 2419 923 2420 927
rect 2440 923 2442 929
rect 2414 922 2420 923
rect 2438 922 2444 923
rect 2416 904 2418 922
rect 2438 918 2439 922
rect 2443 918 2444 922
rect 2438 917 2444 918
rect 2414 903 2420 904
rect 2414 899 2415 903
rect 2419 899 2420 903
rect 2414 898 2420 899
rect 2422 895 2428 896
rect 2294 890 2300 891
rect 2330 891 2336 892
rect 2078 886 2084 887
rect 2168 879 2170 890
rect 2296 879 2298 890
rect 2330 887 2331 891
rect 2335 887 2336 891
rect 2422 891 2423 895
rect 2427 891 2428 895
rect 2456 892 2458 930
rect 2543 929 2547 930
rect 2583 934 2587 935
rect 2583 929 2587 930
rect 2534 927 2540 928
rect 2534 923 2535 927
rect 2539 923 2540 927
rect 2544 923 2546 929
rect 2534 922 2540 923
rect 2542 922 2548 923
rect 2526 895 2532 896
rect 2422 890 2428 891
rect 2454 891 2460 892
rect 2330 886 2336 887
rect 2424 879 2426 890
rect 2454 887 2455 891
rect 2459 887 2460 891
rect 2526 891 2527 895
rect 2531 891 2532 895
rect 2526 890 2532 891
rect 2454 886 2460 887
rect 2528 879 2530 890
rect 1991 878 1995 879
rect 1991 873 1995 874
rect 2047 878 2051 879
rect 2047 873 2051 874
rect 2071 878 2075 879
rect 2071 873 2075 874
rect 2143 878 2147 879
rect 2143 873 2147 874
rect 2167 878 2171 879
rect 2167 873 2171 874
rect 2215 878 2219 879
rect 2215 873 2219 874
rect 2279 878 2283 879
rect 2279 873 2283 874
rect 2295 878 2299 879
rect 2295 873 2299 874
rect 2343 878 2347 879
rect 2343 873 2347 874
rect 2407 878 2411 879
rect 2407 873 2411 874
rect 2423 878 2427 879
rect 2423 873 2427 874
rect 2471 878 2475 879
rect 2471 873 2475 874
rect 2527 878 2531 879
rect 2527 873 2531 874
rect 1982 863 1988 864
rect 1982 859 1983 863
rect 1987 859 1988 863
rect 1992 862 1994 873
rect 2046 863 2052 864
rect 1982 858 1988 859
rect 1990 861 1996 862
rect 1984 828 1986 858
rect 1990 857 1991 861
rect 1995 857 1996 861
rect 2046 859 2047 863
rect 2051 859 2052 863
rect 2072 862 2074 873
rect 2134 863 2140 864
rect 2046 858 2052 859
rect 2070 861 2076 862
rect 1990 856 1996 857
rect 2006 834 2012 835
rect 2006 830 2007 834
rect 2011 830 2012 834
rect 2006 829 2012 830
rect 1950 827 1956 828
rect 1950 823 1951 827
rect 1955 823 1956 827
rect 1950 822 1956 823
rect 1982 827 1988 828
rect 1982 823 1983 827
rect 1987 823 1988 827
rect 1982 822 1988 823
rect 1998 815 2004 816
rect 2008 815 2010 829
rect 1823 814 1827 815
rect 1823 809 1827 810
rect 1831 814 1835 815
rect 1838 811 1839 815
rect 1843 811 1844 815
rect 1838 810 1844 811
rect 1903 814 1907 815
rect 1831 809 1835 810
rect 1798 807 1804 808
rect 1798 803 1799 807
rect 1803 803 1804 807
rect 1824 803 1826 809
rect 1798 802 1804 803
rect 1822 802 1828 803
rect 1800 784 1802 802
rect 1822 798 1823 802
rect 1827 798 1828 802
rect 1822 797 1828 798
rect 1798 783 1804 784
rect 1798 779 1799 783
rect 1803 779 1804 783
rect 1798 778 1804 779
rect 1806 775 1812 776
rect 1734 770 1740 771
rect 1770 771 1776 772
rect 1706 766 1712 767
rect 1736 755 1738 770
rect 1770 767 1771 771
rect 1775 767 1776 771
rect 1806 771 1807 775
rect 1811 771 1812 775
rect 1840 772 1842 810
rect 1903 809 1907 810
rect 1919 814 1923 815
rect 1919 809 1923 810
rect 1991 814 1995 815
rect 1998 811 1999 815
rect 2003 811 2004 815
rect 1998 810 2004 811
rect 2007 814 2011 815
rect 1991 809 1995 810
rect 1904 803 1906 809
rect 1992 803 1994 809
rect 1902 802 1908 803
rect 1902 798 1903 802
rect 1907 798 1908 802
rect 1902 797 1908 798
rect 1990 802 1996 803
rect 1990 798 1991 802
rect 1995 798 1996 802
rect 1990 797 1996 798
rect 1886 775 1892 776
rect 1806 770 1812 771
rect 1838 771 1844 772
rect 1770 766 1776 767
rect 1808 755 1810 770
rect 1838 767 1839 771
rect 1843 767 1844 771
rect 1886 771 1887 775
rect 1891 771 1892 775
rect 1886 770 1892 771
rect 1974 775 1980 776
rect 1974 771 1975 775
rect 1979 771 1980 775
rect 2000 772 2002 810
rect 2007 809 2011 810
rect 2048 808 2050 858
rect 2070 857 2071 861
rect 2075 857 2076 861
rect 2134 859 2135 863
rect 2139 859 2140 863
rect 2144 862 2146 873
rect 2206 863 2212 864
rect 2134 858 2140 859
rect 2142 861 2148 862
rect 2070 856 2076 857
rect 2086 834 2092 835
rect 2086 830 2087 834
rect 2091 830 2092 834
rect 2086 829 2092 830
rect 2088 815 2090 829
rect 2136 828 2138 858
rect 2142 857 2143 861
rect 2147 857 2148 861
rect 2206 859 2207 863
rect 2211 859 2212 863
rect 2216 862 2218 873
rect 2270 863 2276 864
rect 2206 858 2212 859
rect 2214 861 2220 862
rect 2142 856 2148 857
rect 2158 834 2164 835
rect 2158 830 2159 834
rect 2163 830 2164 834
rect 2158 829 2164 830
rect 2126 827 2132 828
rect 2126 823 2127 827
rect 2131 823 2132 827
rect 2126 822 2132 823
rect 2134 827 2140 828
rect 2134 823 2135 827
rect 2139 823 2140 827
rect 2134 822 2140 823
rect 2071 814 2075 815
rect 2071 809 2075 810
rect 2087 814 2091 815
rect 2087 809 2091 810
rect 2046 807 2052 808
rect 2046 803 2047 807
rect 2051 803 2052 807
rect 2072 803 2074 809
rect 2046 802 2052 803
rect 2070 802 2076 803
rect 2070 798 2071 802
rect 2075 798 2076 802
rect 2070 797 2076 798
rect 2128 781 2130 822
rect 2160 815 2162 829
rect 2208 828 2210 858
rect 2214 857 2215 861
rect 2219 857 2220 861
rect 2270 859 2271 863
rect 2275 859 2276 863
rect 2280 862 2282 873
rect 2334 863 2340 864
rect 2270 858 2276 859
rect 2278 861 2284 862
rect 2214 856 2220 857
rect 2230 834 2236 835
rect 2230 830 2231 834
rect 2235 830 2236 834
rect 2230 829 2236 830
rect 2206 827 2212 828
rect 2206 823 2207 827
rect 2211 823 2212 827
rect 2206 822 2212 823
rect 2232 815 2234 829
rect 2272 828 2274 858
rect 2278 857 2279 861
rect 2283 857 2284 861
rect 2334 859 2335 863
rect 2339 859 2340 863
rect 2344 862 2346 873
rect 2398 863 2404 864
rect 2334 858 2340 859
rect 2342 861 2348 862
rect 2278 856 2284 857
rect 2294 834 2300 835
rect 2294 830 2295 834
rect 2299 830 2300 834
rect 2294 829 2300 830
rect 2270 827 2276 828
rect 2270 823 2271 827
rect 2275 823 2276 827
rect 2270 822 2276 823
rect 2296 815 2298 829
rect 2336 828 2338 858
rect 2342 857 2343 861
rect 2347 857 2348 861
rect 2398 859 2399 863
rect 2403 859 2404 863
rect 2408 862 2410 873
rect 2462 863 2468 864
rect 2398 858 2404 859
rect 2406 861 2412 862
rect 2342 856 2348 857
rect 2358 834 2364 835
rect 2358 830 2359 834
rect 2363 830 2364 834
rect 2358 829 2364 830
rect 2334 827 2340 828
rect 2334 823 2335 827
rect 2339 823 2340 827
rect 2334 822 2340 823
rect 2360 815 2362 829
rect 2400 828 2402 858
rect 2406 857 2407 861
rect 2411 857 2412 861
rect 2462 859 2463 863
rect 2467 859 2468 863
rect 2472 862 2474 873
rect 2518 863 2524 864
rect 2462 858 2468 859
rect 2470 861 2476 862
rect 2406 856 2412 857
rect 2422 834 2428 835
rect 2422 830 2423 834
rect 2427 830 2428 834
rect 2422 829 2428 830
rect 2398 827 2404 828
rect 2398 823 2399 827
rect 2403 823 2404 827
rect 2398 822 2404 823
rect 2424 815 2426 829
rect 2464 828 2466 858
rect 2470 857 2471 861
rect 2475 857 2476 861
rect 2518 859 2519 863
rect 2523 859 2524 863
rect 2528 862 2530 873
rect 2536 868 2538 922
rect 2542 918 2543 922
rect 2547 918 2548 922
rect 2542 917 2548 918
rect 2584 914 2586 929
rect 2582 913 2588 914
rect 2582 909 2583 913
rect 2587 909 2588 913
rect 2582 908 2588 909
rect 2582 896 2588 897
rect 2582 892 2583 896
rect 2587 892 2588 896
rect 2582 891 2588 892
rect 2584 879 2586 891
rect 2583 878 2587 879
rect 2583 873 2587 874
rect 2534 867 2540 868
rect 2534 863 2535 867
rect 2539 863 2540 867
rect 2534 862 2540 863
rect 2518 858 2524 859
rect 2526 861 2532 862
rect 2584 861 2586 873
rect 2470 856 2476 857
rect 2486 834 2492 835
rect 2486 830 2487 834
rect 2491 830 2492 834
rect 2486 829 2492 830
rect 2462 827 2468 828
rect 2462 823 2463 827
rect 2467 823 2468 827
rect 2462 822 2468 823
rect 2488 815 2490 829
rect 2520 828 2522 858
rect 2526 857 2527 861
rect 2531 857 2532 861
rect 2526 856 2532 857
rect 2582 860 2588 861
rect 2582 856 2583 860
rect 2587 856 2588 860
rect 2582 855 2588 856
rect 2582 843 2588 844
rect 2582 839 2583 843
rect 2587 839 2588 843
rect 2582 838 2588 839
rect 2542 834 2548 835
rect 2542 830 2543 834
rect 2547 830 2548 834
rect 2542 829 2548 830
rect 2518 827 2524 828
rect 2518 823 2519 827
rect 2523 823 2524 827
rect 2518 822 2524 823
rect 2544 815 2546 829
rect 2584 815 2586 838
rect 2159 814 2163 815
rect 2159 809 2163 810
rect 2231 814 2235 815
rect 2231 809 2235 810
rect 2247 814 2251 815
rect 2247 809 2251 810
rect 2295 814 2299 815
rect 2295 809 2299 810
rect 2335 814 2339 815
rect 2335 809 2339 810
rect 2359 814 2363 815
rect 2359 809 2363 810
rect 2423 814 2427 815
rect 2423 809 2427 810
rect 2487 814 2491 815
rect 2487 809 2491 810
rect 2543 814 2547 815
rect 2543 809 2547 810
rect 2583 814 2587 815
rect 2583 809 2587 810
rect 2150 807 2156 808
rect 2150 803 2151 807
rect 2155 803 2156 807
rect 2160 803 2162 809
rect 2178 807 2184 808
rect 2178 803 2179 807
rect 2183 803 2184 807
rect 2248 803 2250 809
rect 2266 807 2272 808
rect 2266 803 2267 807
rect 2271 803 2272 807
rect 2336 803 2338 809
rect 2424 803 2426 809
rect 2150 802 2156 803
rect 2158 802 2164 803
rect 2178 802 2184 803
rect 2246 802 2252 803
rect 2266 802 2272 803
rect 2334 802 2340 803
rect 2127 780 2131 781
rect 2054 775 2060 776
rect 2127 775 2131 776
rect 2142 775 2148 776
rect 1974 770 1980 771
rect 1998 771 2004 772
rect 1838 766 1844 767
rect 1888 755 1890 770
rect 1976 755 1978 770
rect 1998 767 1999 771
rect 2003 767 2004 771
rect 2054 771 2055 775
rect 2059 771 2060 775
rect 2054 770 2060 771
rect 2086 771 2092 772
rect 1998 766 2004 767
rect 2056 755 2058 770
rect 2086 767 2087 771
rect 2091 767 2092 771
rect 2142 771 2143 775
rect 2147 771 2148 775
rect 2142 770 2148 771
rect 2086 766 2092 767
rect 1367 754 1371 755
rect 1367 749 1371 750
rect 1567 754 1571 755
rect 1567 749 1571 750
rect 1615 754 1619 755
rect 1615 749 1619 750
rect 1623 754 1627 755
rect 1623 749 1627 750
rect 1671 754 1675 755
rect 1671 749 1675 750
rect 1687 754 1691 755
rect 1687 749 1691 750
rect 1735 754 1739 755
rect 1735 749 1739 750
rect 1759 754 1763 755
rect 1759 749 1763 750
rect 1807 754 1811 755
rect 1807 749 1811 750
rect 1839 754 1843 755
rect 1839 749 1843 750
rect 1887 754 1891 755
rect 1887 749 1891 750
rect 1919 754 1923 755
rect 1919 749 1923 750
rect 1975 754 1979 755
rect 1975 749 1979 750
rect 1999 754 2003 755
rect 1999 749 2003 750
rect 2055 754 2059 755
rect 2055 749 2059 750
rect 2079 754 2083 755
rect 2079 749 2083 750
rect 1198 742 1204 743
rect 1326 744 1332 745
rect 1174 740 1180 741
rect 1190 718 1196 719
rect 1190 714 1191 718
rect 1195 714 1196 718
rect 1190 713 1196 714
rect 1103 711 1107 712
rect 1166 711 1172 712
rect 1166 707 1167 711
rect 1171 707 1172 711
rect 1166 706 1172 707
rect 1192 703 1194 713
rect 111 702 115 703
rect 111 697 115 698
rect 159 702 163 703
rect 159 697 163 698
rect 215 702 219 703
rect 215 697 219 698
rect 279 702 283 703
rect 279 697 283 698
rect 295 702 299 703
rect 295 697 299 698
rect 359 702 363 703
rect 366 699 367 703
rect 371 699 372 703
rect 366 698 372 699
rect 399 702 403 703
rect 359 697 363 698
rect 112 682 114 697
rect 134 695 140 696
rect 134 691 135 695
rect 139 691 140 695
rect 160 691 162 697
rect 178 695 184 696
rect 178 691 179 695
rect 183 691 184 695
rect 216 691 218 697
rect 242 695 248 696
rect 242 691 243 695
rect 247 691 248 695
rect 280 691 282 697
rect 360 691 362 697
rect 134 690 140 691
rect 158 690 164 691
rect 178 690 184 691
rect 214 690 220 691
rect 242 690 248 691
rect 278 690 284 691
rect 110 681 116 682
rect 110 677 111 681
rect 115 677 116 681
rect 110 676 116 677
rect 136 672 138 690
rect 158 686 159 690
rect 163 686 164 690
rect 158 685 164 686
rect 134 671 140 672
rect 134 667 135 671
rect 139 667 140 671
rect 134 666 140 667
rect 110 664 116 665
rect 110 660 111 664
rect 115 660 116 664
rect 110 659 116 660
rect 142 663 148 664
rect 142 659 143 663
rect 147 659 148 663
rect 180 660 182 690
rect 214 686 215 690
rect 219 686 220 690
rect 214 685 220 686
rect 198 663 204 664
rect 112 639 114 659
rect 142 658 148 659
rect 178 659 184 660
rect 144 639 146 658
rect 178 655 179 659
rect 183 655 184 659
rect 198 659 199 663
rect 203 659 204 663
rect 244 660 246 690
rect 278 686 279 690
rect 283 686 284 690
rect 278 685 284 686
rect 358 690 364 691
rect 358 686 359 690
rect 363 686 364 690
rect 358 685 364 686
rect 262 663 268 664
rect 198 658 204 659
rect 242 659 248 660
rect 178 654 184 655
rect 200 639 202 658
rect 242 655 243 659
rect 247 655 248 659
rect 262 659 263 663
rect 267 659 268 663
rect 262 658 268 659
rect 342 663 348 664
rect 342 659 343 663
rect 347 659 348 663
rect 368 660 370 698
rect 399 697 403 698
rect 447 702 451 703
rect 447 697 451 698
rect 503 702 507 703
rect 503 697 507 698
rect 535 702 539 703
rect 535 697 539 698
rect 615 702 619 703
rect 615 697 619 698
rect 623 702 627 703
rect 623 697 627 698
rect 711 702 715 703
rect 711 697 715 698
rect 719 702 723 703
rect 726 699 727 703
rect 731 699 732 703
rect 726 698 732 699
rect 791 702 795 703
rect 719 697 723 698
rect 374 695 380 696
rect 374 691 375 695
rect 379 691 380 695
rect 448 691 450 697
rect 466 695 472 696
rect 466 691 467 695
rect 471 691 472 695
rect 536 691 538 697
rect 624 691 626 697
rect 686 695 692 696
rect 686 691 687 695
rect 691 691 692 695
rect 712 691 714 697
rect 374 690 380 691
rect 446 690 452 691
rect 466 690 472 691
rect 534 690 540 691
rect 342 658 348 659
rect 366 659 372 660
rect 242 654 248 655
rect 264 639 266 658
rect 344 639 346 658
rect 366 655 367 659
rect 371 655 372 659
rect 366 654 372 655
rect 376 640 378 690
rect 446 686 447 690
rect 451 686 452 690
rect 446 685 452 686
rect 430 663 436 664
rect 430 659 431 663
rect 435 659 436 663
rect 468 660 470 690
rect 534 686 535 690
rect 539 686 540 690
rect 534 685 540 686
rect 622 690 628 691
rect 686 690 692 691
rect 710 690 716 691
rect 622 686 623 690
rect 627 686 628 690
rect 622 685 628 686
rect 688 672 690 690
rect 710 686 711 690
rect 715 686 716 690
rect 710 685 716 686
rect 686 671 692 672
rect 686 667 687 671
rect 691 667 692 671
rect 686 666 692 667
rect 518 663 524 664
rect 430 658 436 659
rect 466 659 472 660
rect 374 639 380 640
rect 432 639 434 658
rect 466 655 467 659
rect 471 655 472 659
rect 518 659 519 663
rect 523 659 524 663
rect 518 658 524 659
rect 606 663 612 664
rect 606 659 607 663
rect 611 659 612 663
rect 694 663 700 664
rect 606 658 612 659
rect 630 659 636 660
rect 466 654 472 655
rect 520 639 522 658
rect 608 639 610 658
rect 630 655 631 659
rect 635 655 636 659
rect 694 659 695 663
rect 699 659 700 663
rect 728 660 730 698
rect 791 697 795 698
rect 823 702 827 703
rect 823 697 827 698
rect 871 702 875 703
rect 886 699 887 703
rect 891 699 892 703
rect 886 698 892 699
rect 919 702 923 703
rect 871 697 875 698
rect 792 691 794 697
rect 846 695 852 696
rect 846 691 847 695
rect 851 691 852 695
rect 872 691 874 697
rect 790 690 796 691
rect 846 690 852 691
rect 870 690 876 691
rect 790 686 791 690
rect 795 686 796 690
rect 790 685 796 686
rect 848 672 850 690
rect 870 686 871 690
rect 875 686 876 690
rect 870 685 876 686
rect 846 671 852 672
rect 846 667 847 671
rect 851 667 852 671
rect 846 666 852 667
rect 774 663 780 664
rect 694 658 700 659
rect 726 659 732 660
rect 630 654 636 655
rect 111 638 115 639
rect 111 633 115 634
rect 143 638 147 639
rect 143 633 147 634
rect 199 638 203 639
rect 199 633 203 634
rect 255 638 259 639
rect 255 633 259 634
rect 263 638 267 639
rect 263 633 267 634
rect 311 638 315 639
rect 311 633 315 634
rect 343 638 347 639
rect 374 635 375 639
rect 379 635 380 639
rect 374 634 380 635
rect 391 638 395 639
rect 343 633 347 634
rect 391 633 395 634
rect 431 638 435 639
rect 431 633 435 634
rect 479 638 483 639
rect 479 633 483 634
rect 519 638 523 639
rect 519 633 523 634
rect 575 638 579 639
rect 575 633 579 634
rect 607 638 611 639
rect 607 633 611 634
rect 112 621 114 633
rect 144 622 146 633
rect 190 623 196 624
rect 142 621 148 622
rect 110 620 116 621
rect 110 616 111 620
rect 115 616 116 620
rect 142 617 143 621
rect 147 617 148 621
rect 190 619 191 623
rect 195 619 196 623
rect 200 622 202 633
rect 246 623 252 624
rect 190 618 196 619
rect 198 621 204 622
rect 142 616 148 617
rect 110 615 116 616
rect 110 603 116 604
rect 110 599 111 603
rect 115 599 116 603
rect 110 598 116 599
rect 112 579 114 598
rect 158 594 164 595
rect 158 590 159 594
rect 163 590 164 594
rect 158 589 164 590
rect 160 579 162 589
rect 192 588 194 618
rect 198 617 199 621
rect 203 617 204 621
rect 246 619 247 623
rect 251 619 252 623
rect 256 622 258 633
rect 312 622 314 633
rect 334 631 340 632
rect 334 627 335 631
rect 339 627 340 631
rect 334 626 340 627
rect 246 618 252 619
rect 254 621 260 622
rect 198 616 204 617
rect 214 594 220 595
rect 214 590 215 594
rect 219 590 220 594
rect 214 589 220 590
rect 190 587 196 588
rect 190 583 191 587
rect 195 583 196 587
rect 190 582 196 583
rect 216 579 218 589
rect 248 588 250 618
rect 254 617 255 621
rect 259 617 260 621
rect 254 616 260 617
rect 310 621 316 622
rect 310 617 311 621
rect 315 617 316 621
rect 310 616 316 617
rect 270 594 276 595
rect 270 590 271 594
rect 275 590 276 594
rect 270 589 276 590
rect 326 594 332 595
rect 326 590 327 594
rect 331 590 332 594
rect 326 589 332 590
rect 246 587 252 588
rect 246 583 247 587
rect 251 583 252 587
rect 246 582 252 583
rect 272 579 274 589
rect 328 579 330 589
rect 336 588 338 626
rect 342 623 348 624
rect 342 619 343 623
rect 347 619 348 623
rect 392 622 394 633
rect 470 623 476 624
rect 342 618 348 619
rect 390 621 396 622
rect 334 587 340 588
rect 334 583 335 587
rect 339 583 340 587
rect 334 582 340 583
rect 344 580 346 618
rect 390 617 391 621
rect 395 617 396 621
rect 470 619 471 623
rect 475 619 476 623
rect 480 622 482 633
rect 576 622 578 633
rect 470 618 476 619
rect 478 621 484 622
rect 390 616 396 617
rect 406 594 412 595
rect 406 590 407 594
rect 411 590 412 594
rect 406 589 412 590
rect 354 587 360 588
rect 354 583 355 587
rect 359 583 360 587
rect 354 582 360 583
rect 342 579 348 580
rect 111 578 115 579
rect 111 573 115 574
rect 159 578 163 579
rect 159 573 163 574
rect 199 578 203 579
rect 199 573 203 574
rect 215 578 219 579
rect 215 573 219 574
rect 263 578 267 579
rect 263 573 267 574
rect 271 578 275 579
rect 271 573 275 574
rect 327 578 331 579
rect 327 573 331 574
rect 335 578 339 579
rect 342 575 343 579
rect 347 575 348 579
rect 342 574 348 575
rect 335 573 339 574
rect 112 558 114 573
rect 190 571 196 572
rect 190 567 191 571
rect 195 567 196 571
rect 200 567 202 573
rect 264 567 266 573
rect 336 567 338 573
rect 190 566 196 567
rect 198 566 204 567
rect 110 557 116 558
rect 110 553 111 557
rect 115 553 116 557
rect 110 552 116 553
rect 110 540 116 541
rect 110 536 111 540
rect 115 536 116 540
rect 110 535 116 536
rect 182 539 188 540
rect 182 535 183 539
rect 187 535 188 539
rect 112 515 114 535
rect 182 534 188 535
rect 184 515 186 534
rect 192 528 194 566
rect 198 562 199 566
rect 203 562 204 566
rect 198 561 204 562
rect 262 566 268 567
rect 262 562 263 566
rect 267 562 268 566
rect 262 561 268 562
rect 334 566 340 567
rect 334 562 335 566
rect 339 562 340 566
rect 334 561 340 562
rect 246 539 252 540
rect 246 535 247 539
rect 251 535 252 539
rect 246 534 252 535
rect 318 539 324 540
rect 318 535 319 539
rect 323 535 324 539
rect 356 536 358 582
rect 408 579 410 589
rect 472 588 474 618
rect 478 617 479 621
rect 483 617 484 621
rect 478 616 484 617
rect 574 621 580 622
rect 574 617 575 621
rect 579 617 580 621
rect 574 616 580 617
rect 494 594 500 595
rect 494 590 495 594
rect 499 590 500 594
rect 494 589 500 590
rect 590 594 596 595
rect 590 590 591 594
rect 595 590 596 594
rect 590 589 596 590
rect 470 587 476 588
rect 470 583 471 587
rect 475 583 476 587
rect 470 582 476 583
rect 496 579 498 589
rect 592 579 594 589
rect 632 588 634 654
rect 696 639 698 658
rect 726 655 727 659
rect 731 655 732 659
rect 774 659 775 663
rect 779 659 780 663
rect 774 658 780 659
rect 854 663 860 664
rect 854 659 855 663
rect 859 659 860 663
rect 888 660 890 698
rect 919 697 923 698
rect 951 702 955 703
rect 951 697 955 698
rect 1007 702 1011 703
rect 1007 697 1011 698
rect 1039 702 1043 703
rect 1039 697 1043 698
rect 1095 702 1099 703
rect 1095 697 1099 698
rect 1191 702 1195 703
rect 1200 700 1202 742
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 1326 739 1332 740
rect 1368 737 1370 749
rect 1568 738 1570 749
rect 1614 739 1620 740
rect 1566 737 1572 738
rect 1366 736 1372 737
rect 1366 732 1367 736
rect 1371 732 1372 736
rect 1566 733 1567 737
rect 1571 733 1572 737
rect 1614 735 1615 739
rect 1619 735 1620 739
rect 1624 738 1626 749
rect 1678 739 1684 740
rect 1614 734 1620 735
rect 1622 737 1628 738
rect 1566 732 1572 733
rect 1366 731 1372 732
rect 1326 727 1332 728
rect 1326 723 1327 727
rect 1331 723 1332 727
rect 1326 722 1332 723
rect 1328 703 1330 722
rect 1366 719 1372 720
rect 1366 715 1367 719
rect 1371 715 1372 719
rect 1366 714 1372 715
rect 1327 702 1331 703
rect 1191 697 1195 698
rect 1198 699 1204 700
rect 942 695 948 696
rect 942 691 943 695
rect 947 691 948 695
rect 952 691 954 697
rect 1040 691 1042 697
rect 1198 695 1199 699
rect 1203 695 1204 699
rect 1327 697 1331 698
rect 1198 694 1204 695
rect 942 690 948 691
rect 950 690 956 691
rect 934 663 940 664
rect 854 658 860 659
rect 886 659 892 660
rect 726 654 732 655
rect 776 639 778 658
rect 856 639 858 658
rect 886 655 887 659
rect 891 655 892 659
rect 934 659 935 663
rect 939 659 940 663
rect 934 658 940 659
rect 886 654 892 655
rect 936 639 938 658
rect 944 652 946 690
rect 950 686 951 690
rect 955 686 956 690
rect 950 685 956 686
rect 1038 690 1044 691
rect 1038 686 1039 690
rect 1043 686 1044 690
rect 1038 685 1044 686
rect 1328 682 1330 697
rect 1368 695 1370 714
rect 1582 710 1588 711
rect 1582 706 1583 710
rect 1587 706 1588 710
rect 1582 705 1588 706
rect 1584 695 1586 705
rect 1616 704 1618 734
rect 1622 733 1623 737
rect 1627 733 1628 737
rect 1678 735 1679 739
rect 1683 735 1684 739
rect 1688 738 1690 749
rect 1750 739 1756 740
rect 1678 734 1684 735
rect 1686 737 1692 738
rect 1622 732 1628 733
rect 1638 710 1644 711
rect 1638 706 1639 710
rect 1643 706 1644 710
rect 1638 705 1644 706
rect 1614 703 1620 704
rect 1614 699 1615 703
rect 1619 699 1620 703
rect 1614 698 1620 699
rect 1640 695 1642 705
rect 1680 704 1682 734
rect 1686 733 1687 737
rect 1691 733 1692 737
rect 1750 735 1751 739
rect 1755 735 1756 739
rect 1760 738 1762 749
rect 1830 739 1836 740
rect 1750 734 1756 735
rect 1758 737 1764 738
rect 1686 732 1692 733
rect 1702 710 1708 711
rect 1702 706 1703 710
rect 1707 706 1708 710
rect 1702 705 1708 706
rect 1678 703 1684 704
rect 1678 699 1679 703
rect 1683 699 1684 703
rect 1678 698 1684 699
rect 1704 695 1706 705
rect 1752 704 1754 734
rect 1758 733 1759 737
rect 1763 733 1764 737
rect 1830 735 1831 739
rect 1835 735 1836 739
rect 1840 738 1842 749
rect 1910 739 1916 740
rect 1830 734 1836 735
rect 1838 737 1844 738
rect 1758 732 1764 733
rect 1774 710 1780 711
rect 1774 706 1775 710
rect 1779 706 1780 710
rect 1774 705 1780 706
rect 1750 703 1756 704
rect 1750 699 1751 703
rect 1755 699 1756 703
rect 1750 698 1756 699
rect 1776 695 1778 705
rect 1832 704 1834 734
rect 1838 733 1839 737
rect 1843 733 1844 737
rect 1910 735 1911 739
rect 1915 735 1916 739
rect 1920 738 1922 749
rect 2000 738 2002 749
rect 2054 743 2060 744
rect 2030 739 2036 740
rect 1910 734 1916 735
rect 1918 737 1924 738
rect 1838 732 1844 733
rect 1854 710 1860 711
rect 1854 706 1855 710
rect 1859 706 1860 710
rect 1854 705 1860 706
rect 1830 703 1836 704
rect 1830 699 1831 703
rect 1835 699 1836 703
rect 1830 698 1836 699
rect 1838 695 1844 696
rect 1856 695 1858 705
rect 1912 704 1914 734
rect 1918 733 1919 737
rect 1923 733 1924 737
rect 1918 732 1924 733
rect 1998 737 2004 738
rect 1998 733 1999 737
rect 2003 733 2004 737
rect 2030 735 2031 739
rect 2035 735 2036 739
rect 2054 739 2055 743
rect 2059 739 2060 743
rect 2054 738 2060 739
rect 2080 738 2082 749
rect 2030 734 2036 735
rect 1998 732 2004 733
rect 1934 710 1940 711
rect 1934 706 1935 710
rect 1939 706 1940 710
rect 1934 705 1940 706
rect 2014 710 2020 711
rect 2014 706 2015 710
rect 2019 706 2020 710
rect 2014 705 2020 706
rect 1910 703 1916 704
rect 1910 699 1911 703
rect 1915 699 1916 703
rect 1910 698 1916 699
rect 1936 695 1938 705
rect 2016 695 2018 705
rect 2032 696 2034 734
rect 2056 704 2058 738
rect 2078 737 2084 738
rect 2078 733 2079 737
rect 2083 733 2084 737
rect 2078 732 2084 733
rect 2088 704 2090 766
rect 2144 755 2146 770
rect 2143 754 2147 755
rect 2143 749 2147 750
rect 2152 748 2154 802
rect 2158 798 2159 802
rect 2163 798 2164 802
rect 2158 797 2164 798
rect 2180 772 2182 802
rect 2246 798 2247 802
rect 2251 798 2252 802
rect 2246 797 2252 798
rect 2230 775 2236 776
rect 2178 771 2184 772
rect 2178 767 2179 771
rect 2183 767 2184 771
rect 2230 771 2231 775
rect 2235 771 2236 775
rect 2268 772 2270 802
rect 2334 798 2335 802
rect 2339 798 2340 802
rect 2334 797 2340 798
rect 2422 802 2428 803
rect 2422 798 2423 802
rect 2427 798 2428 802
rect 2422 797 2428 798
rect 2584 794 2586 809
rect 2582 793 2588 794
rect 2582 789 2583 793
rect 2587 789 2588 793
rect 2582 788 2588 789
rect 2439 780 2443 781
rect 2318 775 2324 776
rect 2230 770 2236 771
rect 2266 771 2272 772
rect 2178 766 2184 767
rect 2232 755 2234 770
rect 2266 767 2267 771
rect 2271 767 2272 771
rect 2318 771 2319 775
rect 2323 771 2324 775
rect 2318 770 2324 771
rect 2406 775 2412 776
rect 2439 775 2443 776
rect 2582 776 2588 777
rect 2406 771 2407 775
rect 2411 771 2412 775
rect 2440 772 2442 775
rect 2582 772 2583 776
rect 2587 772 2588 776
rect 2406 770 2412 771
rect 2438 771 2444 772
rect 2582 771 2588 772
rect 2266 766 2272 767
rect 2320 755 2322 770
rect 2408 755 2410 770
rect 2438 767 2439 771
rect 2443 767 2444 771
rect 2438 766 2444 767
rect 2584 755 2586 771
rect 2159 754 2163 755
rect 2159 749 2163 750
rect 2231 754 2235 755
rect 2231 749 2235 750
rect 2247 754 2251 755
rect 2247 749 2251 750
rect 2319 754 2323 755
rect 2319 749 2323 750
rect 2335 754 2339 755
rect 2335 749 2339 750
rect 2407 754 2411 755
rect 2407 749 2411 750
rect 2583 754 2587 755
rect 2583 749 2587 750
rect 2150 747 2156 748
rect 2150 743 2151 747
rect 2155 743 2156 747
rect 2150 742 2156 743
rect 2160 738 2162 749
rect 2238 739 2244 740
rect 2158 737 2164 738
rect 2158 733 2159 737
rect 2163 733 2164 737
rect 2238 735 2239 739
rect 2243 735 2244 739
rect 2248 738 2250 749
rect 2326 739 2332 740
rect 2238 734 2244 735
rect 2246 737 2252 738
rect 2158 732 2164 733
rect 2094 710 2100 711
rect 2094 706 2095 710
rect 2099 706 2100 710
rect 2094 705 2100 706
rect 2174 710 2180 711
rect 2174 706 2175 710
rect 2179 706 2180 710
rect 2174 705 2180 706
rect 2054 703 2060 704
rect 2054 699 2055 703
rect 2059 699 2060 703
rect 2054 698 2060 699
rect 2086 703 2092 704
rect 2086 699 2087 703
rect 2091 699 2092 703
rect 2086 698 2092 699
rect 2030 695 2036 696
rect 2096 695 2098 705
rect 2138 703 2144 704
rect 2138 699 2139 703
rect 2143 699 2144 703
rect 2138 698 2144 699
rect 1367 694 1371 695
rect 1367 689 1371 690
rect 1415 694 1419 695
rect 1415 689 1419 690
rect 1511 694 1515 695
rect 1511 689 1515 690
rect 1583 694 1587 695
rect 1583 689 1587 690
rect 1615 694 1619 695
rect 1615 689 1619 690
rect 1639 694 1643 695
rect 1639 689 1643 690
rect 1703 694 1707 695
rect 1703 689 1707 690
rect 1719 694 1723 695
rect 1719 689 1723 690
rect 1775 694 1779 695
rect 1775 689 1779 690
rect 1823 694 1827 695
rect 1838 691 1839 695
rect 1843 691 1844 695
rect 1838 690 1844 691
rect 1855 694 1859 695
rect 1823 689 1827 690
rect 1326 681 1332 682
rect 1326 677 1327 681
rect 1331 677 1332 681
rect 1326 676 1332 677
rect 1368 674 1370 689
rect 1406 687 1412 688
rect 1406 683 1407 687
rect 1411 683 1412 687
rect 1416 683 1418 689
rect 1434 687 1440 688
rect 1434 683 1435 687
rect 1439 683 1440 687
rect 1512 683 1514 689
rect 1616 683 1618 689
rect 1720 683 1722 689
rect 1738 687 1744 688
rect 1738 683 1739 687
rect 1743 683 1744 687
rect 1824 683 1826 689
rect 1406 682 1412 683
rect 1414 682 1420 683
rect 1434 682 1440 683
rect 1510 682 1516 683
rect 1366 673 1372 674
rect 1366 669 1367 673
rect 1371 669 1372 673
rect 1366 668 1372 669
rect 1326 664 1332 665
rect 1022 663 1028 664
rect 1022 659 1023 663
rect 1027 659 1028 663
rect 1326 660 1327 664
rect 1331 660 1332 664
rect 1326 659 1332 660
rect 1022 658 1028 659
rect 942 651 948 652
rect 942 647 943 651
rect 947 647 948 651
rect 942 646 948 647
rect 1024 639 1026 658
rect 1328 639 1330 659
rect 1366 656 1372 657
rect 1366 652 1367 656
rect 1371 652 1372 656
rect 1366 651 1372 652
rect 1398 655 1404 656
rect 1398 651 1399 655
rect 1403 651 1404 655
rect 1368 639 1370 651
rect 1398 650 1404 651
rect 1400 639 1402 650
rect 679 638 683 639
rect 679 633 683 634
rect 695 638 699 639
rect 695 633 699 634
rect 775 638 779 639
rect 775 633 779 634
rect 783 638 787 639
rect 783 633 787 634
rect 855 638 859 639
rect 855 633 859 634
rect 887 638 891 639
rect 887 633 891 634
rect 935 638 939 639
rect 935 633 939 634
rect 991 638 995 639
rect 991 633 995 634
rect 1023 638 1027 639
rect 1023 633 1027 634
rect 1087 638 1091 639
rect 1087 633 1091 634
rect 1191 638 1195 639
rect 1191 633 1195 634
rect 1271 638 1275 639
rect 1271 633 1275 634
rect 1327 638 1331 639
rect 1327 633 1331 634
rect 1367 638 1371 639
rect 1367 633 1371 634
rect 1399 638 1403 639
rect 1399 633 1403 634
rect 670 623 676 624
rect 670 619 671 623
rect 675 619 676 623
rect 680 622 682 633
rect 774 623 780 624
rect 670 618 676 619
rect 678 621 684 622
rect 672 588 674 618
rect 678 617 679 621
rect 683 617 684 621
rect 774 619 775 623
rect 779 619 780 623
rect 784 622 786 633
rect 878 623 884 624
rect 774 618 780 619
rect 782 621 788 622
rect 678 616 684 617
rect 694 594 700 595
rect 694 590 695 594
rect 699 590 700 594
rect 694 589 700 590
rect 630 587 636 588
rect 630 583 631 587
rect 635 583 636 587
rect 630 582 636 583
rect 670 587 676 588
rect 670 583 671 587
rect 675 583 676 587
rect 670 582 676 583
rect 696 579 698 589
rect 776 588 778 618
rect 782 617 783 621
rect 787 617 788 621
rect 878 619 879 623
rect 883 619 884 623
rect 888 622 890 633
rect 918 623 924 624
rect 878 618 884 619
rect 886 621 892 622
rect 782 616 788 617
rect 798 594 804 595
rect 798 590 799 594
rect 803 590 804 594
rect 798 589 804 590
rect 774 587 780 588
rect 774 583 775 587
rect 779 583 780 587
rect 774 582 780 583
rect 800 579 802 589
rect 880 588 882 618
rect 886 617 887 621
rect 891 617 892 621
rect 918 619 919 623
rect 923 619 924 623
rect 992 622 994 633
rect 1078 623 1084 624
rect 918 618 924 619
rect 990 621 996 622
rect 886 616 892 617
rect 902 594 908 595
rect 902 590 903 594
rect 907 590 908 594
rect 902 589 908 590
rect 878 587 884 588
rect 878 583 879 587
rect 883 583 884 587
rect 878 582 884 583
rect 846 579 852 580
rect 904 579 906 589
rect 407 578 411 579
rect 407 573 411 574
rect 415 578 419 579
rect 415 573 419 574
rect 495 578 499 579
rect 495 573 499 574
rect 511 578 515 579
rect 511 573 515 574
rect 591 578 595 579
rect 591 573 595 574
rect 615 578 619 579
rect 615 573 619 574
rect 695 578 699 579
rect 695 573 699 574
rect 719 578 723 579
rect 719 573 723 574
rect 799 578 803 579
rect 799 573 803 574
rect 831 578 835 579
rect 846 575 847 579
rect 851 575 852 579
rect 846 574 852 575
rect 903 578 907 579
rect 831 573 835 574
rect 390 571 396 572
rect 390 567 391 571
rect 395 567 396 571
rect 416 567 418 573
rect 512 567 514 573
rect 530 571 536 572
rect 530 567 531 571
rect 535 567 536 571
rect 616 567 618 573
rect 720 567 722 573
rect 806 571 812 572
rect 806 567 807 571
rect 811 567 812 571
rect 832 567 834 573
rect 390 566 396 567
rect 414 566 420 567
rect 392 548 394 566
rect 414 562 415 566
rect 419 562 420 566
rect 414 561 420 562
rect 510 566 516 567
rect 530 566 536 567
rect 614 566 620 567
rect 510 562 511 566
rect 515 562 516 566
rect 510 561 516 562
rect 390 547 396 548
rect 390 543 391 547
rect 395 543 396 547
rect 390 542 396 543
rect 398 539 404 540
rect 318 534 324 535
rect 354 535 360 536
rect 190 527 196 528
rect 190 523 191 527
rect 195 523 196 527
rect 190 522 196 523
rect 248 515 250 534
rect 320 515 322 534
rect 354 531 355 535
rect 359 531 360 535
rect 398 535 399 539
rect 403 535 404 539
rect 398 534 404 535
rect 494 539 500 540
rect 494 535 495 539
rect 499 535 500 539
rect 532 536 534 566
rect 614 562 615 566
rect 619 562 620 566
rect 614 561 620 562
rect 718 566 724 567
rect 806 566 812 567
rect 830 566 836 567
rect 718 562 719 566
rect 723 562 724 566
rect 718 561 724 562
rect 808 548 810 566
rect 830 562 831 566
rect 835 562 836 566
rect 830 561 836 562
rect 806 547 812 548
rect 806 543 807 547
rect 811 543 812 547
rect 806 542 812 543
rect 598 539 604 540
rect 494 534 500 535
rect 530 535 536 536
rect 354 530 360 531
rect 400 515 402 534
rect 496 515 498 534
rect 530 531 531 535
rect 535 531 536 535
rect 598 535 599 539
rect 603 535 604 539
rect 598 534 604 535
rect 702 539 708 540
rect 702 535 703 539
rect 707 535 708 539
rect 814 539 820 540
rect 702 534 708 535
rect 726 535 732 536
rect 530 530 536 531
rect 600 515 602 534
rect 704 515 706 534
rect 726 531 727 535
rect 731 531 732 535
rect 814 535 815 539
rect 819 535 820 539
rect 848 536 850 574
rect 903 573 907 574
rect 920 572 922 618
rect 990 617 991 621
rect 995 617 996 621
rect 1078 619 1079 623
rect 1083 619 1084 623
rect 1088 622 1090 633
rect 1182 623 1188 624
rect 1078 618 1084 619
rect 1086 621 1092 622
rect 990 616 996 617
rect 1006 594 1012 595
rect 1006 590 1007 594
rect 1011 590 1012 594
rect 1006 589 1012 590
rect 1008 579 1010 589
rect 1080 588 1082 618
rect 1086 617 1087 621
rect 1091 617 1092 621
rect 1182 619 1183 623
rect 1187 619 1188 623
rect 1192 622 1194 633
rect 1262 623 1268 624
rect 1182 618 1188 619
rect 1190 621 1196 622
rect 1086 616 1092 617
rect 1102 594 1108 595
rect 1102 590 1103 594
rect 1107 590 1108 594
rect 1102 589 1108 590
rect 1070 587 1076 588
rect 1070 583 1071 587
rect 1075 583 1076 587
rect 1070 582 1076 583
rect 1078 587 1084 588
rect 1078 583 1079 587
rect 1083 583 1084 587
rect 1078 582 1084 583
rect 943 578 947 579
rect 943 573 947 574
rect 1007 578 1011 579
rect 1007 573 1011 574
rect 1063 578 1067 579
rect 1063 573 1067 574
rect 918 571 924 572
rect 918 567 919 571
rect 923 567 924 571
rect 944 567 946 573
rect 1064 567 1066 573
rect 918 566 924 567
rect 942 566 948 567
rect 942 562 943 566
rect 947 562 948 566
rect 942 561 948 562
rect 1062 566 1068 567
rect 1062 562 1063 566
rect 1067 562 1068 566
rect 1062 561 1068 562
rect 926 539 932 540
rect 814 534 820 535
rect 846 535 852 536
rect 726 530 732 531
rect 111 514 115 515
rect 111 509 115 510
rect 183 514 187 515
rect 183 509 187 510
rect 247 514 251 515
rect 247 509 251 510
rect 303 514 307 515
rect 303 509 307 510
rect 319 514 323 515
rect 319 509 323 510
rect 359 514 363 515
rect 359 509 363 510
rect 399 514 403 515
rect 399 509 403 510
rect 423 514 427 515
rect 423 509 427 510
rect 495 514 499 515
rect 495 509 499 510
rect 575 514 579 515
rect 575 509 579 510
rect 599 514 603 515
rect 599 509 603 510
rect 647 514 651 515
rect 647 509 651 510
rect 703 514 707 515
rect 703 509 707 510
rect 719 514 723 515
rect 719 509 723 510
rect 112 497 114 509
rect 304 498 306 509
rect 350 499 356 500
rect 302 497 308 498
rect 110 496 116 497
rect 110 492 111 496
rect 115 492 116 496
rect 302 493 303 497
rect 307 493 308 497
rect 350 495 351 499
rect 355 495 356 499
rect 360 498 362 509
rect 414 499 420 500
rect 350 494 356 495
rect 358 497 364 498
rect 302 492 308 493
rect 110 491 116 492
rect 110 479 116 480
rect 110 475 111 479
rect 115 475 116 479
rect 110 474 116 475
rect 112 455 114 474
rect 318 470 324 471
rect 318 466 319 470
rect 323 466 324 470
rect 318 465 324 466
rect 320 455 322 465
rect 352 464 354 494
rect 358 493 359 497
rect 363 493 364 497
rect 414 495 415 499
rect 419 495 420 499
rect 424 498 426 509
rect 496 498 498 509
rect 518 507 524 508
rect 518 503 519 507
rect 523 503 524 507
rect 518 502 524 503
rect 414 494 420 495
rect 422 497 428 498
rect 358 492 364 493
rect 374 470 380 471
rect 374 466 375 470
rect 379 466 380 470
rect 374 465 380 466
rect 350 463 356 464
rect 350 459 351 463
rect 355 459 356 463
rect 350 458 356 459
rect 376 455 378 465
rect 416 464 418 494
rect 422 493 423 497
rect 427 493 428 497
rect 422 492 428 493
rect 494 497 500 498
rect 494 493 495 497
rect 499 493 500 497
rect 494 492 500 493
rect 438 470 444 471
rect 438 466 439 470
rect 443 466 444 470
rect 438 465 444 466
rect 510 470 516 471
rect 510 466 511 470
rect 515 466 516 470
rect 510 465 516 466
rect 414 463 420 464
rect 414 459 415 463
rect 419 459 420 463
rect 414 458 420 459
rect 440 455 442 465
rect 512 455 514 465
rect 520 464 522 502
rect 526 499 532 500
rect 526 495 527 499
rect 531 495 532 499
rect 576 498 578 509
rect 638 499 644 500
rect 526 494 532 495
rect 574 497 580 498
rect 518 463 524 464
rect 518 459 519 463
rect 523 459 524 463
rect 518 458 524 459
rect 528 456 530 494
rect 574 493 575 497
rect 579 493 580 497
rect 638 495 639 499
rect 643 495 644 499
rect 648 498 650 509
rect 720 498 722 509
rect 638 494 644 495
rect 646 497 652 498
rect 574 492 580 493
rect 590 470 596 471
rect 590 466 591 470
rect 595 466 596 470
rect 590 465 596 466
rect 582 463 588 464
rect 582 459 583 463
rect 587 459 588 463
rect 582 458 588 459
rect 526 455 532 456
rect 111 454 115 455
rect 111 449 115 450
rect 319 454 323 455
rect 319 449 323 450
rect 375 454 379 455
rect 375 449 379 450
rect 439 454 443 455
rect 439 449 443 450
rect 455 454 459 455
rect 455 449 459 450
rect 511 454 515 455
rect 526 451 527 455
rect 531 451 532 455
rect 526 450 532 451
rect 575 454 579 455
rect 511 449 515 450
rect 575 449 579 450
rect 112 434 114 449
rect 430 447 436 448
rect 430 443 431 447
rect 435 443 436 447
rect 456 443 458 449
rect 470 447 476 448
rect 470 443 471 447
rect 475 443 476 447
rect 512 443 514 449
rect 530 447 536 448
rect 530 443 531 447
rect 535 443 536 447
rect 576 443 578 449
rect 430 442 436 443
rect 454 442 460 443
rect 470 442 476 443
rect 510 442 516 443
rect 530 442 536 443
rect 574 442 580 443
rect 110 433 116 434
rect 110 429 111 433
rect 115 429 116 433
rect 110 428 116 429
rect 432 424 434 442
rect 454 438 455 442
rect 459 438 460 442
rect 454 437 460 438
rect 430 423 436 424
rect 430 419 431 423
rect 435 419 436 423
rect 430 418 436 419
rect 110 416 116 417
rect 110 412 111 416
rect 115 412 116 416
rect 110 411 116 412
rect 438 415 444 416
rect 438 411 439 415
rect 443 411 444 415
rect 472 412 474 442
rect 510 438 511 442
rect 515 438 516 442
rect 510 437 516 438
rect 494 415 500 416
rect 112 395 114 411
rect 438 410 444 411
rect 470 411 476 412
rect 440 395 442 410
rect 470 407 471 411
rect 475 407 476 411
rect 494 411 495 415
rect 499 411 500 415
rect 532 412 534 442
rect 574 438 575 442
rect 579 438 580 442
rect 574 437 580 438
rect 558 415 564 416
rect 494 410 500 411
rect 530 411 536 412
rect 470 406 476 407
rect 496 395 498 410
rect 530 407 531 411
rect 535 407 536 411
rect 558 411 559 415
rect 563 411 564 415
rect 584 412 586 458
rect 592 455 594 465
rect 640 464 642 494
rect 646 493 647 497
rect 651 493 652 497
rect 646 492 652 493
rect 718 497 724 498
rect 718 493 719 497
rect 723 493 724 497
rect 718 492 724 493
rect 662 470 668 471
rect 662 466 663 470
rect 667 466 668 470
rect 662 465 668 466
rect 638 463 644 464
rect 638 459 639 463
rect 643 459 644 463
rect 638 458 644 459
rect 664 455 666 465
rect 728 464 730 530
rect 816 515 818 534
rect 846 531 847 535
rect 851 531 852 535
rect 926 535 927 539
rect 931 535 932 539
rect 926 534 932 535
rect 1046 539 1052 540
rect 1046 535 1047 539
rect 1051 535 1052 539
rect 1072 536 1074 582
rect 1104 579 1106 589
rect 1184 588 1186 618
rect 1190 617 1191 621
rect 1195 617 1196 621
rect 1262 619 1263 623
rect 1267 619 1268 623
rect 1272 622 1274 633
rect 1262 618 1268 619
rect 1270 621 1276 622
rect 1328 621 1330 633
rect 1368 621 1370 633
rect 1400 622 1402 633
rect 1408 629 1410 682
rect 1414 678 1415 682
rect 1419 678 1420 682
rect 1414 677 1420 678
rect 1436 652 1438 682
rect 1510 678 1511 682
rect 1515 678 1516 682
rect 1510 677 1516 678
rect 1614 682 1620 683
rect 1614 678 1615 682
rect 1619 678 1620 682
rect 1614 677 1620 678
rect 1718 682 1724 683
rect 1738 682 1744 683
rect 1822 682 1828 683
rect 1718 678 1719 682
rect 1723 678 1724 682
rect 1718 677 1724 678
rect 1494 655 1500 656
rect 1434 651 1440 652
rect 1434 647 1435 651
rect 1439 647 1440 651
rect 1494 651 1495 655
rect 1499 651 1500 655
rect 1494 650 1500 651
rect 1598 655 1604 656
rect 1598 651 1599 655
rect 1603 651 1604 655
rect 1598 650 1604 651
rect 1702 655 1708 656
rect 1702 651 1703 655
rect 1707 651 1708 655
rect 1740 652 1742 682
rect 1822 678 1823 682
rect 1827 678 1828 682
rect 1822 677 1828 678
rect 1806 655 1812 656
rect 1702 650 1708 651
rect 1738 651 1744 652
rect 1434 646 1440 647
rect 1496 639 1498 650
rect 1600 639 1602 650
rect 1704 639 1706 650
rect 1738 647 1739 651
rect 1743 647 1744 651
rect 1806 651 1807 655
rect 1811 651 1812 655
rect 1840 652 1842 690
rect 1855 689 1859 690
rect 1927 694 1931 695
rect 1927 689 1931 690
rect 1935 694 1939 695
rect 1935 689 1939 690
rect 2015 694 2019 695
rect 2015 689 2019 690
rect 2023 694 2027 695
rect 2030 691 2031 695
rect 2035 691 2036 695
rect 2030 690 2036 691
rect 2095 694 2099 695
rect 2023 689 2027 690
rect 2095 689 2099 690
rect 2119 694 2123 695
rect 2119 689 2123 690
rect 1928 683 1930 689
rect 1946 687 1952 688
rect 1946 683 1947 687
rect 1951 683 1952 687
rect 2024 683 2026 689
rect 2120 683 2122 689
rect 1926 682 1932 683
rect 1946 682 1952 683
rect 2022 682 2028 683
rect 1926 678 1927 682
rect 1931 678 1932 682
rect 1926 677 1932 678
rect 1910 655 1916 656
rect 1806 650 1812 651
rect 1838 651 1844 652
rect 1738 646 1744 647
rect 1808 639 1810 650
rect 1838 647 1839 651
rect 1843 647 1844 651
rect 1910 651 1911 655
rect 1915 651 1916 655
rect 1948 652 1950 682
rect 2022 678 2023 682
rect 2027 678 2028 682
rect 2022 677 2028 678
rect 2118 682 2124 683
rect 2118 678 2119 682
rect 2123 678 2124 682
rect 2118 677 2124 678
rect 2006 655 2012 656
rect 1910 650 1916 651
rect 1946 651 1952 652
rect 1838 646 1844 647
rect 1912 639 1914 650
rect 1946 647 1947 651
rect 1951 647 1952 651
rect 2006 651 2007 655
rect 2011 651 2012 655
rect 2102 655 2108 656
rect 2006 650 2012 651
rect 2030 651 2036 652
rect 1946 646 1952 647
rect 2008 639 2010 650
rect 2030 647 2031 651
rect 2035 647 2036 651
rect 2102 651 2103 655
rect 2107 651 2108 655
rect 2140 652 2142 698
rect 2176 695 2178 705
rect 2240 704 2242 734
rect 2246 733 2247 737
rect 2251 733 2252 737
rect 2326 735 2327 739
rect 2331 735 2332 739
rect 2336 738 2338 749
rect 2326 734 2332 735
rect 2334 737 2340 738
rect 2584 737 2586 749
rect 2246 732 2252 733
rect 2262 710 2268 711
rect 2262 706 2263 710
rect 2267 706 2268 710
rect 2262 705 2268 706
rect 2238 703 2244 704
rect 2238 699 2239 703
rect 2243 699 2244 703
rect 2238 698 2244 699
rect 2222 695 2228 696
rect 2264 695 2266 705
rect 2328 704 2330 734
rect 2334 733 2335 737
rect 2339 733 2340 737
rect 2334 732 2340 733
rect 2582 736 2588 737
rect 2582 732 2583 736
rect 2587 732 2588 736
rect 2582 731 2588 732
rect 2582 719 2588 720
rect 2582 715 2583 719
rect 2587 715 2588 719
rect 2582 714 2588 715
rect 2350 710 2356 711
rect 2350 706 2351 710
rect 2355 706 2356 710
rect 2350 705 2356 706
rect 2326 703 2332 704
rect 2326 699 2327 703
rect 2331 699 2332 703
rect 2326 698 2332 699
rect 2352 695 2354 705
rect 2584 695 2586 714
rect 2175 694 2179 695
rect 2175 689 2179 690
rect 2207 694 2211 695
rect 2222 691 2223 695
rect 2227 691 2228 695
rect 2222 690 2228 691
rect 2263 694 2267 695
rect 2207 689 2211 690
rect 2182 687 2188 688
rect 2182 683 2183 687
rect 2187 683 2188 687
rect 2208 683 2210 689
rect 2182 682 2188 683
rect 2206 682 2212 683
rect 2184 664 2186 682
rect 2206 678 2207 682
rect 2211 678 2212 682
rect 2206 677 2212 678
rect 2182 663 2188 664
rect 2182 659 2183 663
rect 2187 659 2188 663
rect 2182 658 2188 659
rect 2190 655 2196 656
rect 2102 650 2108 651
rect 2138 651 2144 652
rect 2030 646 2036 647
rect 1495 638 1499 639
rect 1495 633 1499 634
rect 1511 638 1515 639
rect 1511 633 1515 634
rect 1599 638 1603 639
rect 1647 638 1651 639
rect 1599 633 1603 634
rect 1638 635 1644 636
rect 1407 628 1411 629
rect 1407 623 1411 624
rect 1422 623 1428 624
rect 1398 621 1404 622
rect 1190 616 1196 617
rect 1206 594 1212 595
rect 1206 590 1207 594
rect 1211 590 1212 594
rect 1206 589 1212 590
rect 1182 587 1188 588
rect 1182 583 1183 587
rect 1187 583 1188 587
rect 1182 582 1188 583
rect 1198 579 1204 580
rect 1208 579 1210 589
rect 1264 588 1266 618
rect 1270 617 1271 621
rect 1275 617 1276 621
rect 1270 616 1276 617
rect 1326 620 1332 621
rect 1326 616 1327 620
rect 1331 616 1332 620
rect 1326 615 1332 616
rect 1366 620 1372 621
rect 1366 616 1367 620
rect 1371 616 1372 620
rect 1398 617 1399 621
rect 1403 617 1404 621
rect 1422 619 1423 623
rect 1427 619 1428 623
rect 1512 622 1514 633
rect 1638 631 1639 635
rect 1643 631 1644 635
rect 1647 633 1651 634
rect 1703 638 1707 639
rect 1703 633 1707 634
rect 1783 638 1787 639
rect 1783 633 1787 634
rect 1807 638 1811 639
rect 1807 633 1811 634
rect 1911 638 1915 639
rect 1911 633 1915 634
rect 2007 638 2011 639
rect 2007 633 2011 634
rect 1638 630 1644 631
rect 1422 618 1428 619
rect 1510 621 1516 622
rect 1398 616 1404 617
rect 1366 615 1372 616
rect 1326 603 1332 604
rect 1326 599 1327 603
rect 1331 599 1332 603
rect 1326 598 1332 599
rect 1366 603 1372 604
rect 1366 599 1367 603
rect 1371 599 1372 603
rect 1366 598 1372 599
rect 1286 594 1292 595
rect 1286 590 1287 594
rect 1291 590 1292 594
rect 1286 589 1292 590
rect 1262 587 1268 588
rect 1262 583 1263 587
rect 1267 583 1268 587
rect 1262 582 1268 583
rect 1288 579 1290 589
rect 1328 579 1330 598
rect 1103 578 1107 579
rect 1103 573 1107 574
rect 1183 578 1187 579
rect 1198 575 1199 579
rect 1203 575 1204 579
rect 1198 574 1204 575
rect 1207 578 1211 579
rect 1183 573 1187 574
rect 1158 571 1164 572
rect 1158 567 1159 571
rect 1163 567 1164 571
rect 1184 567 1186 573
rect 1158 566 1164 567
rect 1182 566 1188 567
rect 1160 548 1162 566
rect 1182 562 1183 566
rect 1187 562 1188 566
rect 1182 561 1188 562
rect 1158 547 1164 548
rect 1158 543 1159 547
rect 1163 543 1164 547
rect 1158 542 1164 543
rect 1166 539 1172 540
rect 1046 534 1052 535
rect 1070 535 1076 536
rect 846 530 852 531
rect 928 515 930 534
rect 1048 515 1050 534
rect 1070 531 1071 535
rect 1075 531 1076 535
rect 1166 535 1167 539
rect 1171 535 1172 539
rect 1200 536 1202 574
rect 1207 573 1211 574
rect 1287 578 1291 579
rect 1287 573 1291 574
rect 1327 578 1331 579
rect 1368 575 1370 598
rect 1414 594 1420 595
rect 1414 590 1415 594
rect 1419 590 1420 594
rect 1414 589 1420 590
rect 1416 575 1418 589
rect 1424 576 1426 618
rect 1510 617 1511 621
rect 1515 617 1516 621
rect 1510 616 1516 617
rect 1526 594 1532 595
rect 1526 590 1527 594
rect 1531 590 1532 594
rect 1526 589 1532 590
rect 1490 587 1496 588
rect 1490 583 1491 587
rect 1495 583 1496 587
rect 1490 582 1496 583
rect 1422 575 1428 576
rect 1327 573 1331 574
rect 1367 574 1371 575
rect 1288 567 1290 573
rect 1286 566 1292 567
rect 1286 562 1287 566
rect 1291 562 1292 566
rect 1286 561 1292 562
rect 1328 558 1330 573
rect 1367 569 1371 570
rect 1415 574 1419 575
rect 1422 571 1423 575
rect 1427 571 1428 575
rect 1422 570 1428 571
rect 1471 574 1475 575
rect 1415 569 1419 570
rect 1471 569 1475 570
rect 1326 557 1332 558
rect 1326 553 1327 557
rect 1331 553 1332 557
rect 1368 554 1370 569
rect 1390 567 1396 568
rect 1390 563 1391 567
rect 1395 563 1396 567
rect 1416 563 1418 569
rect 1434 567 1440 568
rect 1434 563 1435 567
rect 1439 563 1440 567
rect 1472 563 1474 569
rect 1390 562 1396 563
rect 1414 562 1420 563
rect 1434 562 1440 563
rect 1470 562 1476 563
rect 1326 552 1332 553
rect 1366 553 1372 554
rect 1366 549 1367 553
rect 1371 549 1372 553
rect 1366 548 1372 549
rect 1392 544 1394 562
rect 1414 558 1415 562
rect 1419 558 1420 562
rect 1414 557 1420 558
rect 1390 543 1396 544
rect 1326 540 1332 541
rect 1270 539 1276 540
rect 1166 534 1172 535
rect 1198 535 1204 536
rect 1070 530 1076 531
rect 1168 515 1170 534
rect 1198 531 1199 535
rect 1203 531 1204 535
rect 1270 535 1271 539
rect 1275 535 1276 539
rect 1326 536 1327 540
rect 1331 536 1332 540
rect 1390 539 1391 543
rect 1395 539 1396 543
rect 1390 538 1396 539
rect 1326 535 1332 536
rect 1366 536 1372 537
rect 1270 534 1276 535
rect 1198 530 1204 531
rect 1272 515 1274 534
rect 1328 515 1330 535
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1398 535 1404 536
rect 1398 531 1399 535
rect 1403 531 1404 535
rect 1436 532 1438 562
rect 1470 558 1471 562
rect 1475 558 1476 562
rect 1470 557 1476 558
rect 1454 535 1460 536
rect 1368 519 1370 531
rect 1398 530 1404 531
rect 1434 531 1440 532
rect 1400 519 1402 530
rect 1434 527 1435 531
rect 1439 527 1440 531
rect 1454 531 1455 535
rect 1459 531 1460 535
rect 1492 532 1494 582
rect 1528 575 1530 589
rect 1640 588 1642 630
rect 1648 622 1650 633
rect 1774 623 1780 624
rect 1646 621 1652 622
rect 1646 617 1647 621
rect 1651 617 1652 621
rect 1774 619 1775 623
rect 1779 619 1780 623
rect 1784 622 1786 633
rect 1815 628 1819 629
rect 1814 623 1820 624
rect 1774 618 1780 619
rect 1782 621 1788 622
rect 1646 616 1652 617
rect 1662 594 1668 595
rect 1662 590 1663 594
rect 1667 590 1668 594
rect 1662 589 1668 590
rect 1638 587 1644 588
rect 1638 583 1639 587
rect 1643 583 1644 587
rect 1638 582 1644 583
rect 1654 575 1660 576
rect 1664 575 1666 589
rect 1776 588 1778 618
rect 1782 617 1783 621
rect 1787 617 1788 621
rect 1814 619 1815 623
rect 1819 619 1820 623
rect 1912 622 1914 633
rect 1938 623 1944 624
rect 1814 618 1820 619
rect 1910 621 1916 622
rect 1782 616 1788 617
rect 1910 617 1911 621
rect 1915 617 1916 621
rect 1938 619 1939 623
rect 1943 619 1944 623
rect 1938 618 1944 619
rect 1910 616 1916 617
rect 1798 594 1804 595
rect 1798 590 1799 594
rect 1803 590 1804 594
rect 1798 589 1804 590
rect 1926 594 1932 595
rect 1926 590 1927 594
rect 1931 590 1932 594
rect 1926 589 1932 590
rect 1774 587 1780 588
rect 1774 583 1775 587
rect 1779 583 1780 587
rect 1774 582 1780 583
rect 1800 575 1802 589
rect 1928 575 1930 589
rect 1527 574 1531 575
rect 1527 569 1531 570
rect 1551 574 1555 575
rect 1551 569 1555 570
rect 1647 574 1651 575
rect 1654 571 1655 575
rect 1659 571 1660 575
rect 1654 570 1660 571
rect 1663 574 1667 575
rect 1647 569 1651 570
rect 1552 563 1554 569
rect 1622 567 1628 568
rect 1622 563 1623 567
rect 1627 563 1628 567
rect 1648 563 1650 569
rect 1550 562 1556 563
rect 1622 562 1628 563
rect 1646 562 1652 563
rect 1550 558 1551 562
rect 1555 558 1556 562
rect 1550 557 1556 558
rect 1624 544 1626 562
rect 1646 558 1647 562
rect 1651 558 1652 562
rect 1646 557 1652 558
rect 1622 543 1628 544
rect 1622 539 1623 543
rect 1627 539 1628 543
rect 1622 538 1628 539
rect 1534 535 1540 536
rect 1454 530 1460 531
rect 1490 531 1496 532
rect 1434 526 1440 527
rect 1456 519 1458 530
rect 1490 527 1491 531
rect 1495 527 1496 531
rect 1534 531 1535 535
rect 1539 531 1540 535
rect 1534 530 1540 531
rect 1630 535 1636 536
rect 1630 531 1631 535
rect 1635 531 1636 535
rect 1656 532 1658 570
rect 1663 569 1667 570
rect 1751 574 1755 575
rect 1751 569 1755 570
rect 1799 574 1803 575
rect 1799 569 1803 570
rect 1855 574 1859 575
rect 1855 569 1859 570
rect 1927 574 1931 575
rect 1927 569 1931 570
rect 1718 567 1724 568
rect 1718 563 1719 567
rect 1723 563 1724 567
rect 1752 563 1754 569
rect 1770 567 1776 568
rect 1770 563 1771 567
rect 1775 563 1776 567
rect 1856 563 1858 569
rect 1940 568 1942 618
rect 2032 588 2034 646
rect 2104 639 2106 650
rect 2138 647 2139 651
rect 2143 647 2144 651
rect 2190 651 2191 655
rect 2195 651 2196 655
rect 2224 652 2226 690
rect 2263 689 2267 690
rect 2295 694 2299 695
rect 2295 689 2299 690
rect 2351 694 2355 695
rect 2351 689 2355 690
rect 2391 694 2395 695
rect 2583 694 2587 695
rect 2391 689 2395 690
rect 2438 691 2444 692
rect 2286 687 2292 688
rect 2286 683 2287 687
rect 2291 683 2292 687
rect 2296 683 2298 689
rect 2392 683 2394 689
rect 2438 687 2439 691
rect 2443 687 2444 691
rect 2583 689 2587 690
rect 2438 686 2444 687
rect 2286 682 2292 683
rect 2294 682 2300 683
rect 2278 655 2284 656
rect 2190 650 2196 651
rect 2222 651 2228 652
rect 2138 646 2144 647
rect 2192 639 2194 650
rect 2222 647 2223 651
rect 2227 647 2228 651
rect 2278 651 2279 655
rect 2283 651 2284 655
rect 2278 650 2284 651
rect 2222 646 2228 647
rect 2280 639 2282 650
rect 2288 644 2290 682
rect 2294 678 2295 682
rect 2299 678 2300 682
rect 2294 677 2300 678
rect 2390 682 2396 683
rect 2390 678 2391 682
rect 2395 678 2396 682
rect 2390 677 2396 678
rect 2374 655 2380 656
rect 2374 651 2375 655
rect 2379 651 2380 655
rect 2374 650 2380 651
rect 2286 643 2292 644
rect 2286 639 2287 643
rect 2291 639 2292 643
rect 2376 639 2378 650
rect 2039 638 2043 639
rect 2039 633 2043 634
rect 2103 638 2107 639
rect 2103 633 2107 634
rect 2159 638 2163 639
rect 2159 633 2163 634
rect 2191 638 2195 639
rect 2191 633 2195 634
rect 2279 638 2283 639
rect 2286 638 2292 639
rect 2375 638 2379 639
rect 2279 633 2283 634
rect 2375 633 2379 634
rect 2407 638 2411 639
rect 2407 633 2411 634
rect 2040 622 2042 633
rect 2160 622 2162 633
rect 2270 623 2276 624
rect 2038 621 2044 622
rect 2038 617 2039 621
rect 2043 617 2044 621
rect 2038 616 2044 617
rect 2158 621 2164 622
rect 2158 617 2159 621
rect 2163 617 2164 621
rect 2270 619 2271 623
rect 2275 619 2276 623
rect 2280 622 2282 633
rect 2398 623 2404 624
rect 2270 618 2276 619
rect 2278 621 2284 622
rect 2158 616 2164 617
rect 2054 594 2060 595
rect 2054 590 2055 594
rect 2059 590 2060 594
rect 2054 589 2060 590
rect 2174 594 2180 595
rect 2174 590 2175 594
rect 2179 590 2180 594
rect 2174 589 2180 590
rect 2030 587 2036 588
rect 2030 583 2031 587
rect 2035 583 2036 587
rect 2030 582 2036 583
rect 2056 575 2058 589
rect 2176 575 2178 589
rect 2272 588 2274 618
rect 2278 617 2279 621
rect 2283 617 2284 621
rect 2398 619 2399 623
rect 2403 619 2404 623
rect 2408 622 2410 633
rect 2440 624 2442 686
rect 2584 674 2586 689
rect 2582 673 2588 674
rect 2582 669 2583 673
rect 2587 669 2588 673
rect 2582 668 2588 669
rect 2582 656 2588 657
rect 2582 652 2583 656
rect 2587 652 2588 656
rect 2582 651 2588 652
rect 2584 639 2586 651
rect 2583 638 2587 639
rect 2583 633 2587 634
rect 2438 623 2444 624
rect 2398 618 2404 619
rect 2406 621 2412 622
rect 2278 616 2284 617
rect 2294 594 2300 595
rect 2294 590 2295 594
rect 2299 590 2300 594
rect 2294 589 2300 590
rect 2254 587 2260 588
rect 2254 583 2255 587
rect 2259 583 2260 587
rect 2254 582 2260 583
rect 2270 587 2276 588
rect 2270 583 2271 587
rect 2275 583 2276 587
rect 2270 582 2276 583
rect 1959 574 1963 575
rect 1959 569 1963 570
rect 2055 574 2059 575
rect 2055 569 2059 570
rect 2151 574 2155 575
rect 2151 569 2155 570
rect 2175 574 2179 575
rect 2175 569 2179 570
rect 2239 574 2243 575
rect 2239 569 2243 570
rect 1938 567 1944 568
rect 1938 563 1939 567
rect 1943 563 1944 567
rect 1960 563 1962 569
rect 2056 563 2058 569
rect 2074 567 2080 568
rect 2074 563 2075 567
rect 2079 563 2080 567
rect 2152 563 2154 569
rect 2214 567 2220 568
rect 2214 563 2215 567
rect 2219 563 2220 567
rect 2240 563 2242 569
rect 1718 562 1724 563
rect 1750 562 1756 563
rect 1770 562 1776 563
rect 1854 562 1860 563
rect 1938 562 1944 563
rect 1958 562 1964 563
rect 1630 530 1636 531
rect 1654 531 1660 532
rect 1490 526 1496 527
rect 1536 519 1538 530
rect 1632 519 1634 530
rect 1654 527 1655 531
rect 1659 527 1660 531
rect 1654 526 1660 527
rect 1367 518 1371 519
rect 791 514 795 515
rect 791 509 795 510
rect 815 514 819 515
rect 815 509 819 510
rect 863 514 867 515
rect 863 509 867 510
rect 927 514 931 515
rect 927 509 931 510
rect 935 514 939 515
rect 935 509 939 510
rect 1007 514 1011 515
rect 1007 509 1011 510
rect 1047 514 1051 515
rect 1047 509 1051 510
rect 1087 514 1091 515
rect 1087 509 1091 510
rect 1167 514 1171 515
rect 1167 509 1171 510
rect 1271 514 1275 515
rect 1271 509 1275 510
rect 1327 514 1331 515
rect 1367 513 1371 514
rect 1399 518 1403 519
rect 1399 513 1403 514
rect 1455 518 1459 519
rect 1455 513 1459 514
rect 1535 518 1539 519
rect 1535 513 1539 514
rect 1599 518 1603 519
rect 1599 513 1603 514
rect 1631 518 1635 519
rect 1631 513 1635 514
rect 1671 518 1675 519
rect 1671 513 1675 514
rect 1327 509 1331 510
rect 774 499 780 500
rect 774 495 775 499
rect 779 495 780 499
rect 792 498 794 509
rect 854 499 860 500
rect 774 494 780 495
rect 790 497 796 498
rect 734 470 740 471
rect 734 466 735 470
rect 739 466 740 470
rect 734 465 740 466
rect 726 463 732 464
rect 726 459 727 463
rect 731 459 732 463
rect 726 458 732 459
rect 736 455 738 465
rect 776 464 778 494
rect 790 493 791 497
rect 795 493 796 497
rect 854 495 855 499
rect 859 495 860 499
rect 864 498 866 509
rect 926 499 932 500
rect 854 494 860 495
rect 862 497 868 498
rect 790 492 796 493
rect 806 470 812 471
rect 806 466 807 470
rect 811 466 812 470
rect 806 465 812 466
rect 774 463 780 464
rect 774 459 775 463
rect 779 459 780 463
rect 774 458 780 459
rect 742 455 748 456
rect 808 455 810 465
rect 856 464 858 494
rect 862 493 863 497
rect 867 493 868 497
rect 926 495 927 499
rect 931 495 932 499
rect 936 498 938 509
rect 998 499 1004 500
rect 926 494 932 495
rect 934 497 940 498
rect 862 492 868 493
rect 878 470 884 471
rect 878 466 879 470
rect 883 466 884 470
rect 878 465 884 466
rect 854 463 860 464
rect 854 459 855 463
rect 859 459 860 463
rect 854 458 860 459
rect 880 455 882 465
rect 928 464 930 494
rect 934 493 935 497
rect 939 493 940 497
rect 998 495 999 499
rect 1003 495 1004 499
rect 1008 498 1010 509
rect 1078 499 1084 500
rect 998 494 1004 495
rect 1006 497 1012 498
rect 934 492 940 493
rect 950 470 956 471
rect 950 466 951 470
rect 955 466 956 470
rect 950 465 956 466
rect 926 463 932 464
rect 926 459 927 463
rect 931 459 932 463
rect 926 458 932 459
rect 952 455 954 465
rect 1000 464 1002 494
rect 1006 493 1007 497
rect 1011 493 1012 497
rect 1078 495 1079 499
rect 1083 495 1084 499
rect 1088 498 1090 509
rect 1110 499 1116 500
rect 1078 494 1084 495
rect 1086 497 1092 498
rect 1006 492 1012 493
rect 1022 470 1028 471
rect 1022 466 1023 470
rect 1027 466 1028 470
rect 1022 465 1028 466
rect 998 463 1004 464
rect 998 459 999 463
rect 1003 459 1004 463
rect 998 458 1004 459
rect 1024 455 1026 465
rect 1080 464 1082 494
rect 1086 493 1087 497
rect 1091 493 1092 497
rect 1110 495 1111 499
rect 1115 495 1116 499
rect 1328 497 1330 509
rect 1368 501 1370 513
rect 1536 502 1538 513
rect 1542 511 1548 512
rect 1542 507 1543 511
rect 1547 507 1548 511
rect 1542 506 1548 507
rect 1534 501 1540 502
rect 1366 500 1372 501
rect 1110 494 1116 495
rect 1326 496 1332 497
rect 1086 492 1092 493
rect 1102 470 1108 471
rect 1102 466 1103 470
rect 1107 466 1108 470
rect 1102 465 1108 466
rect 1078 463 1084 464
rect 1078 459 1079 463
rect 1083 459 1084 463
rect 1078 458 1084 459
rect 1104 455 1106 465
rect 1112 456 1114 494
rect 1326 492 1327 496
rect 1331 492 1332 496
rect 1366 496 1367 500
rect 1371 496 1372 500
rect 1534 497 1535 501
rect 1539 497 1540 501
rect 1534 496 1540 497
rect 1366 495 1372 496
rect 1326 491 1332 492
rect 1366 483 1372 484
rect 1326 479 1332 480
rect 1326 475 1327 479
rect 1331 475 1332 479
rect 1366 479 1367 483
rect 1371 479 1372 483
rect 1366 478 1372 479
rect 1326 474 1332 475
rect 1110 455 1116 456
rect 1328 455 1330 474
rect 1368 455 1370 478
rect 1544 468 1546 506
rect 1590 503 1596 504
rect 1590 499 1591 503
rect 1595 499 1596 503
rect 1600 502 1602 513
rect 1662 503 1668 504
rect 1590 498 1596 499
rect 1598 501 1604 502
rect 1550 474 1556 475
rect 1550 470 1551 474
rect 1555 470 1556 474
rect 1550 469 1556 470
rect 1542 467 1548 468
rect 1542 463 1543 467
rect 1547 463 1548 467
rect 1542 462 1548 463
rect 1552 455 1554 469
rect 1592 468 1594 498
rect 1598 497 1599 501
rect 1603 497 1604 501
rect 1662 499 1663 503
rect 1667 499 1668 503
rect 1672 502 1674 513
rect 1720 504 1722 562
rect 1750 558 1751 562
rect 1755 558 1756 562
rect 1750 557 1756 558
rect 1734 535 1740 536
rect 1734 531 1735 535
rect 1739 531 1740 535
rect 1772 532 1774 562
rect 1854 558 1855 562
rect 1859 558 1860 562
rect 1854 557 1860 558
rect 1958 558 1959 562
rect 1963 558 1964 562
rect 1958 557 1964 558
rect 2054 562 2060 563
rect 2074 562 2080 563
rect 2150 562 2156 563
rect 2214 562 2220 563
rect 2238 562 2244 563
rect 2054 558 2055 562
rect 2059 558 2060 562
rect 2054 557 2060 558
rect 1838 535 1844 536
rect 1734 530 1740 531
rect 1770 531 1776 532
rect 1736 519 1738 530
rect 1770 527 1771 531
rect 1775 527 1776 531
rect 1838 531 1839 535
rect 1843 531 1844 535
rect 1838 530 1844 531
rect 1942 535 1948 536
rect 1942 531 1943 535
rect 1947 531 1948 535
rect 1942 530 1948 531
rect 2038 535 2044 536
rect 2038 531 2039 535
rect 2043 531 2044 535
rect 2076 532 2078 562
rect 2150 558 2151 562
rect 2155 558 2156 562
rect 2150 557 2156 558
rect 2216 544 2218 562
rect 2238 558 2239 562
rect 2243 558 2244 562
rect 2238 557 2244 558
rect 2214 543 2220 544
rect 2214 539 2215 543
rect 2219 539 2220 543
rect 2214 538 2220 539
rect 2134 535 2140 536
rect 2038 530 2044 531
rect 2074 531 2080 532
rect 1770 526 1776 527
rect 1840 519 1842 530
rect 1944 519 1946 530
rect 2022 523 2028 524
rect 2022 519 2023 523
rect 2027 519 2028 523
rect 2040 519 2042 530
rect 2074 527 2075 531
rect 2079 527 2080 531
rect 2134 531 2135 535
rect 2139 531 2140 535
rect 2134 530 2140 531
rect 2222 535 2228 536
rect 2222 531 2223 535
rect 2227 531 2228 535
rect 2256 532 2258 582
rect 2296 575 2298 589
rect 2400 588 2402 618
rect 2406 617 2407 621
rect 2411 617 2412 621
rect 2438 619 2439 623
rect 2443 619 2444 623
rect 2584 621 2586 633
rect 2438 618 2444 619
rect 2582 620 2588 621
rect 2406 616 2412 617
rect 2582 616 2583 620
rect 2587 616 2588 620
rect 2582 615 2588 616
rect 2582 603 2588 604
rect 2582 599 2583 603
rect 2587 599 2588 603
rect 2582 598 2588 599
rect 2422 594 2428 595
rect 2422 590 2423 594
rect 2427 590 2428 594
rect 2422 589 2428 590
rect 2398 587 2404 588
rect 2398 583 2399 587
rect 2403 583 2404 587
rect 2398 582 2404 583
rect 2414 575 2420 576
rect 2424 575 2426 589
rect 2584 575 2586 598
rect 2295 574 2299 575
rect 2295 569 2299 570
rect 2319 574 2323 575
rect 2319 569 2323 570
rect 2399 574 2403 575
rect 2414 571 2415 575
rect 2419 571 2420 575
rect 2414 570 2420 571
rect 2423 574 2427 575
rect 2399 569 2403 570
rect 2320 563 2322 569
rect 2374 567 2380 568
rect 2374 563 2375 567
rect 2379 563 2380 567
rect 2400 563 2402 569
rect 2318 562 2324 563
rect 2374 562 2380 563
rect 2398 562 2404 563
rect 2318 558 2319 562
rect 2323 558 2324 562
rect 2318 557 2324 558
rect 2376 544 2378 562
rect 2398 558 2399 562
rect 2403 558 2404 562
rect 2398 557 2404 558
rect 2374 543 2380 544
rect 2374 539 2375 543
rect 2379 539 2380 543
rect 2374 538 2380 539
rect 2302 535 2308 536
rect 2222 530 2228 531
rect 2254 531 2260 532
rect 2074 526 2080 527
rect 2136 519 2138 530
rect 2224 519 2226 530
rect 2254 527 2255 531
rect 2259 527 2260 531
rect 2302 531 2303 535
rect 2307 531 2308 535
rect 2302 530 2308 531
rect 2382 535 2388 536
rect 2382 531 2383 535
rect 2387 531 2388 535
rect 2416 532 2418 570
rect 2423 569 2427 570
rect 2479 574 2483 575
rect 2479 569 2483 570
rect 2543 574 2547 575
rect 2543 569 2547 570
rect 2583 574 2587 575
rect 2583 569 2587 570
rect 2434 567 2440 568
rect 2434 563 2435 567
rect 2439 563 2440 567
rect 2480 563 2482 569
rect 2498 567 2504 568
rect 2498 563 2499 567
rect 2503 563 2504 567
rect 2544 563 2546 569
rect 2434 562 2440 563
rect 2478 562 2484 563
rect 2498 562 2504 563
rect 2542 562 2548 563
rect 2382 530 2388 531
rect 2414 531 2420 532
rect 2254 526 2260 527
rect 2304 519 2306 530
rect 2384 519 2386 530
rect 2414 527 2415 531
rect 2419 527 2420 531
rect 2414 526 2420 527
rect 1735 518 1739 519
rect 1735 513 1739 514
rect 1751 518 1755 519
rect 1751 513 1755 514
rect 1839 518 1843 519
rect 1839 513 1843 514
rect 1927 518 1931 519
rect 1927 513 1931 514
rect 1943 518 1947 519
rect 1943 513 1947 514
rect 2015 518 2019 519
rect 2022 518 2028 519
rect 2039 518 2043 519
rect 2015 513 2019 514
rect 1718 503 1724 504
rect 1662 498 1668 499
rect 1670 501 1676 502
rect 1598 496 1604 497
rect 1614 474 1620 475
rect 1614 470 1615 474
rect 1619 470 1620 474
rect 1614 469 1620 470
rect 1590 467 1596 468
rect 1590 463 1591 467
rect 1595 463 1596 467
rect 1590 462 1596 463
rect 1616 455 1618 469
rect 1664 468 1666 498
rect 1670 497 1671 501
rect 1675 497 1676 501
rect 1718 499 1719 503
rect 1723 499 1724 503
rect 1752 502 1754 513
rect 1830 503 1836 504
rect 1718 498 1724 499
rect 1750 501 1756 502
rect 1670 496 1676 497
rect 1750 497 1751 501
rect 1755 497 1756 501
rect 1830 499 1831 503
rect 1835 499 1836 503
rect 1840 502 1842 513
rect 1918 503 1924 504
rect 1830 498 1836 499
rect 1838 501 1844 502
rect 1750 496 1756 497
rect 1686 474 1692 475
rect 1686 470 1687 474
rect 1691 470 1692 474
rect 1686 469 1692 470
rect 1766 474 1772 475
rect 1766 470 1767 474
rect 1771 470 1772 474
rect 1766 469 1772 470
rect 1662 467 1668 468
rect 1662 463 1663 467
rect 1667 463 1668 467
rect 1662 462 1668 463
rect 1688 455 1690 469
rect 1768 455 1770 469
rect 1832 468 1834 498
rect 1838 497 1839 501
rect 1843 497 1844 501
rect 1918 499 1919 503
rect 1923 499 1924 503
rect 1928 502 1930 513
rect 2016 502 2018 513
rect 1918 498 1924 499
rect 1926 501 1932 502
rect 1838 496 1844 497
rect 1854 474 1860 475
rect 1854 470 1855 474
rect 1859 470 1860 474
rect 1854 469 1860 470
rect 1774 467 1780 468
rect 1774 463 1775 467
rect 1779 463 1780 467
rect 1774 462 1780 463
rect 1830 467 1836 468
rect 1830 463 1831 467
rect 1835 463 1836 467
rect 1830 462 1836 463
rect 591 454 595 455
rect 591 449 595 450
rect 647 454 651 455
rect 647 449 651 450
rect 663 454 667 455
rect 663 449 667 450
rect 727 454 731 455
rect 727 449 731 450
rect 735 454 739 455
rect 742 451 743 455
rect 747 451 748 455
rect 742 450 748 451
rect 799 454 803 455
rect 735 449 739 450
rect 648 443 650 449
rect 702 447 708 448
rect 702 443 703 447
rect 707 443 708 447
rect 728 443 730 449
rect 646 442 652 443
rect 702 442 708 443
rect 726 442 732 443
rect 646 438 647 442
rect 651 438 652 442
rect 646 437 652 438
rect 704 424 706 442
rect 726 438 727 442
rect 731 438 732 442
rect 726 437 732 438
rect 702 423 708 424
rect 702 419 703 423
rect 707 419 708 423
rect 702 418 708 419
rect 630 415 636 416
rect 558 410 564 411
rect 582 411 588 412
rect 530 406 536 407
rect 560 395 562 410
rect 582 407 583 411
rect 587 407 588 411
rect 630 411 631 415
rect 635 411 636 415
rect 630 410 636 411
rect 710 415 716 416
rect 710 411 711 415
rect 715 411 716 415
rect 744 412 746 450
rect 799 449 803 450
rect 807 454 811 455
rect 807 449 811 450
rect 871 454 875 455
rect 871 449 875 450
rect 879 454 883 455
rect 879 449 883 450
rect 943 454 947 455
rect 943 449 947 450
rect 951 454 955 455
rect 951 449 955 450
rect 1015 454 1019 455
rect 1015 449 1019 450
rect 1023 454 1027 455
rect 1023 449 1027 450
rect 1087 454 1091 455
rect 1087 449 1091 450
rect 1103 454 1107 455
rect 1110 451 1111 455
rect 1115 451 1116 455
rect 1110 450 1116 451
rect 1159 454 1163 455
rect 1103 449 1107 450
rect 1159 449 1163 450
rect 1239 454 1243 455
rect 1239 449 1243 450
rect 1327 454 1331 455
rect 1327 449 1331 450
rect 1367 454 1371 455
rect 1367 449 1371 450
rect 1551 454 1555 455
rect 1551 449 1555 450
rect 1615 454 1619 455
rect 1615 449 1619 450
rect 1647 454 1651 455
rect 1647 449 1651 450
rect 1687 454 1691 455
rect 1687 449 1691 450
rect 1703 454 1707 455
rect 1703 449 1707 450
rect 1759 454 1763 455
rect 1759 449 1763 450
rect 1767 454 1771 455
rect 1767 449 1771 450
rect 790 447 796 448
rect 790 443 791 447
rect 795 443 796 447
rect 800 443 802 449
rect 872 443 874 449
rect 890 447 896 448
rect 890 443 891 447
rect 895 443 896 447
rect 944 443 946 449
rect 962 447 968 448
rect 962 443 963 447
rect 967 443 968 447
rect 1016 443 1018 449
rect 1034 447 1040 448
rect 1034 443 1035 447
rect 1039 443 1040 447
rect 1088 443 1090 449
rect 1122 447 1128 448
rect 1122 443 1123 447
rect 1127 443 1128 447
rect 1160 443 1162 449
rect 1178 447 1184 448
rect 1178 443 1179 447
rect 1183 443 1184 447
rect 1240 443 1242 449
rect 790 442 796 443
rect 798 442 804 443
rect 782 415 788 416
rect 710 410 716 411
rect 742 411 748 412
rect 582 406 588 407
rect 632 395 634 410
rect 712 395 714 410
rect 742 407 743 411
rect 747 407 748 411
rect 782 411 783 415
rect 787 411 788 415
rect 782 410 788 411
rect 742 406 748 407
rect 784 395 786 410
rect 111 394 115 395
rect 111 389 115 390
rect 415 394 419 395
rect 415 389 419 390
rect 439 394 443 395
rect 439 389 443 390
rect 471 394 475 395
rect 471 389 475 390
rect 495 394 499 395
rect 495 389 499 390
rect 535 394 539 395
rect 535 389 539 390
rect 559 394 563 395
rect 559 389 563 390
rect 607 394 611 395
rect 607 389 611 390
rect 631 394 635 395
rect 631 389 635 390
rect 687 394 691 395
rect 687 389 691 390
rect 711 394 715 395
rect 711 389 715 390
rect 767 394 771 395
rect 767 389 771 390
rect 783 394 787 395
rect 783 389 787 390
rect 112 377 114 389
rect 416 378 418 389
rect 462 379 468 380
rect 414 377 420 378
rect 110 376 116 377
rect 110 372 111 376
rect 115 372 116 376
rect 414 373 415 377
rect 419 373 420 377
rect 462 375 463 379
rect 467 375 468 379
rect 472 378 474 389
rect 526 379 532 380
rect 462 374 468 375
rect 470 377 476 378
rect 414 372 420 373
rect 110 371 116 372
rect 110 359 116 360
rect 110 355 111 359
rect 115 355 116 359
rect 110 354 116 355
rect 112 335 114 354
rect 430 350 436 351
rect 430 346 431 350
rect 435 346 436 350
rect 430 345 436 346
rect 432 335 434 345
rect 464 344 466 374
rect 470 373 471 377
rect 475 373 476 377
rect 526 375 527 379
rect 531 375 532 379
rect 536 378 538 389
rect 598 379 604 380
rect 526 374 532 375
rect 534 377 540 378
rect 470 372 476 373
rect 486 350 492 351
rect 486 346 487 350
rect 491 346 492 350
rect 486 345 492 346
rect 454 343 460 344
rect 454 339 455 343
rect 459 339 460 343
rect 454 338 460 339
rect 462 343 468 344
rect 462 339 463 343
rect 467 339 468 343
rect 462 338 468 339
rect 111 334 115 335
rect 111 329 115 330
rect 431 334 435 335
rect 431 329 435 330
rect 112 314 114 329
rect 438 327 444 328
rect 438 323 439 327
rect 443 323 444 327
rect 438 322 444 323
rect 110 313 116 314
rect 110 309 111 313
rect 115 309 116 313
rect 110 308 116 309
rect 440 304 442 322
rect 438 303 444 304
rect 438 299 439 303
rect 443 299 444 303
rect 438 298 444 299
rect 110 296 116 297
rect 110 292 111 296
rect 115 292 116 296
rect 110 291 116 292
rect 446 295 452 296
rect 446 291 447 295
rect 451 291 452 295
rect 112 275 114 291
rect 446 290 452 291
rect 448 275 450 290
rect 456 288 458 338
rect 488 335 490 345
rect 528 344 530 374
rect 534 373 535 377
rect 539 373 540 377
rect 598 375 599 379
rect 603 375 604 379
rect 608 378 610 389
rect 678 379 684 380
rect 598 374 604 375
rect 606 377 612 378
rect 534 372 540 373
rect 550 350 556 351
rect 550 346 551 350
rect 555 346 556 350
rect 550 345 556 346
rect 526 343 532 344
rect 526 339 527 343
rect 531 339 532 343
rect 526 338 532 339
rect 552 335 554 345
rect 600 344 602 374
rect 606 373 607 377
rect 611 373 612 377
rect 678 375 679 379
rect 683 375 684 379
rect 688 378 690 389
rect 710 379 716 380
rect 678 374 684 375
rect 686 377 692 378
rect 606 372 612 373
rect 622 350 628 351
rect 622 346 623 350
rect 627 346 628 350
rect 622 345 628 346
rect 598 343 604 344
rect 598 339 599 343
rect 603 339 604 343
rect 598 338 604 339
rect 624 335 626 345
rect 680 344 682 374
rect 686 373 687 377
rect 691 373 692 377
rect 710 375 711 379
rect 715 375 716 379
rect 768 378 770 389
rect 792 380 794 442
rect 798 438 799 442
rect 803 438 804 442
rect 798 437 804 438
rect 870 442 876 443
rect 890 442 896 443
rect 942 442 948 443
rect 962 442 968 443
rect 1014 442 1020 443
rect 1034 442 1040 443
rect 1086 442 1092 443
rect 1122 442 1128 443
rect 1158 442 1164 443
rect 1178 442 1184 443
rect 1238 442 1244 443
rect 870 438 871 442
rect 875 438 876 442
rect 870 437 876 438
rect 854 415 860 416
rect 854 411 855 415
rect 859 411 860 415
rect 892 412 894 442
rect 942 438 943 442
rect 947 438 948 442
rect 942 437 948 438
rect 926 415 932 416
rect 854 410 860 411
rect 890 411 896 412
rect 856 395 858 410
rect 890 407 891 411
rect 895 407 896 411
rect 926 411 927 415
rect 931 411 932 415
rect 964 412 966 442
rect 1014 438 1015 442
rect 1019 438 1020 442
rect 1014 437 1020 438
rect 998 415 1004 416
rect 926 410 932 411
rect 962 411 968 412
rect 890 406 896 407
rect 928 395 930 410
rect 962 407 963 411
rect 967 407 968 411
rect 998 411 999 415
rect 1003 411 1004 415
rect 1036 412 1038 442
rect 1086 438 1087 442
rect 1091 438 1092 442
rect 1086 437 1092 438
rect 1124 416 1126 442
rect 1158 438 1159 442
rect 1163 438 1164 442
rect 1158 437 1164 438
rect 1070 415 1076 416
rect 998 410 1004 411
rect 1034 411 1040 412
rect 962 406 968 407
rect 1000 395 1002 410
rect 1034 407 1035 411
rect 1039 407 1040 411
rect 1070 411 1071 415
rect 1075 411 1076 415
rect 1070 410 1076 411
rect 1122 415 1128 416
rect 1122 411 1123 415
rect 1127 411 1128 415
rect 1122 410 1128 411
rect 1142 415 1148 416
rect 1142 411 1143 415
rect 1147 411 1148 415
rect 1180 412 1182 442
rect 1238 438 1239 442
rect 1243 438 1244 442
rect 1238 437 1244 438
rect 1328 434 1330 449
rect 1368 434 1370 449
rect 1622 447 1628 448
rect 1622 443 1623 447
rect 1627 443 1628 447
rect 1648 443 1650 449
rect 1666 447 1672 448
rect 1666 443 1667 447
rect 1671 443 1672 447
rect 1704 443 1706 449
rect 1722 447 1728 448
rect 1722 443 1723 447
rect 1727 443 1728 447
rect 1760 443 1762 449
rect 1622 442 1628 443
rect 1646 442 1652 443
rect 1666 442 1672 443
rect 1702 442 1708 443
rect 1722 442 1728 443
rect 1758 442 1764 443
rect 1326 433 1332 434
rect 1326 429 1327 433
rect 1331 429 1332 433
rect 1326 428 1332 429
rect 1366 433 1372 434
rect 1366 429 1367 433
rect 1371 429 1372 433
rect 1366 428 1372 429
rect 1624 424 1626 442
rect 1646 438 1647 442
rect 1651 438 1652 442
rect 1646 437 1652 438
rect 1622 423 1628 424
rect 1622 419 1623 423
rect 1627 419 1628 423
rect 1622 418 1628 419
rect 1326 416 1332 417
rect 1222 415 1228 416
rect 1142 410 1148 411
rect 1178 411 1184 412
rect 1034 406 1040 407
rect 1072 395 1074 410
rect 1144 395 1146 410
rect 1178 407 1179 411
rect 1183 407 1184 411
rect 1222 411 1223 415
rect 1227 411 1228 415
rect 1326 412 1327 416
rect 1331 412 1332 416
rect 1222 410 1228 411
rect 1254 411 1260 412
rect 1326 411 1332 412
rect 1366 416 1372 417
rect 1366 412 1367 416
rect 1371 412 1372 416
rect 1366 411 1372 412
rect 1630 415 1636 416
rect 1630 411 1631 415
rect 1635 411 1636 415
rect 1668 412 1670 442
rect 1702 438 1703 442
rect 1707 438 1708 442
rect 1702 437 1708 438
rect 1686 415 1692 416
rect 1178 406 1184 407
rect 1224 395 1226 410
rect 1254 407 1255 411
rect 1259 407 1260 411
rect 1254 406 1260 407
rect 847 394 851 395
rect 847 389 851 390
rect 855 394 859 395
rect 855 389 859 390
rect 927 394 931 395
rect 927 389 931 390
rect 999 394 1003 395
rect 999 389 1003 390
rect 1007 394 1011 395
rect 1007 389 1011 390
rect 1071 394 1075 395
rect 1071 389 1075 390
rect 1087 394 1091 395
rect 1087 389 1091 390
rect 1143 394 1147 395
rect 1143 389 1147 390
rect 1175 394 1179 395
rect 1175 389 1179 390
rect 1223 394 1227 395
rect 1223 389 1227 390
rect 790 379 796 380
rect 710 374 716 375
rect 766 377 772 378
rect 686 372 692 373
rect 702 350 708 351
rect 702 346 703 350
rect 707 346 708 350
rect 702 345 708 346
rect 678 343 684 344
rect 678 339 679 343
rect 683 339 684 343
rect 678 338 684 339
rect 704 335 706 345
rect 712 336 714 374
rect 766 373 767 377
rect 771 373 772 377
rect 790 375 791 379
rect 795 375 796 379
rect 848 378 850 389
rect 928 378 930 389
rect 934 387 940 388
rect 934 383 935 387
rect 939 383 940 387
rect 934 382 940 383
rect 790 374 796 375
rect 846 377 852 378
rect 766 372 772 373
rect 846 373 847 377
rect 851 373 852 377
rect 846 372 852 373
rect 926 377 932 378
rect 926 373 927 377
rect 931 373 932 377
rect 926 372 932 373
rect 782 350 788 351
rect 782 346 783 350
rect 787 346 788 350
rect 782 345 788 346
rect 862 350 868 351
rect 862 346 863 350
rect 867 346 868 350
rect 862 345 868 346
rect 710 335 716 336
rect 784 335 786 345
rect 854 343 860 344
rect 854 339 855 343
rect 859 339 860 343
rect 854 338 860 339
rect 463 334 467 335
rect 463 329 467 330
rect 487 334 491 335
rect 487 329 491 330
rect 519 334 523 335
rect 519 329 523 330
rect 551 334 555 335
rect 551 329 555 330
rect 575 334 579 335
rect 575 329 579 330
rect 623 334 627 335
rect 623 329 627 330
rect 631 334 635 335
rect 631 329 635 330
rect 695 334 699 335
rect 695 329 699 330
rect 703 334 707 335
rect 710 331 711 335
rect 715 331 716 335
rect 710 330 716 331
rect 767 334 771 335
rect 703 329 707 330
rect 767 329 771 330
rect 783 334 787 335
rect 783 329 787 330
rect 847 334 851 335
rect 847 329 851 330
rect 464 323 466 329
rect 510 327 516 328
rect 510 323 511 327
rect 515 323 516 327
rect 520 323 522 329
rect 576 323 578 329
rect 594 327 600 328
rect 594 323 595 327
rect 599 323 600 327
rect 632 323 634 329
rect 650 327 656 328
rect 650 323 651 327
rect 655 323 656 327
rect 696 323 698 329
rect 768 323 770 329
rect 848 323 850 329
rect 462 322 468 323
rect 510 322 516 323
rect 518 322 524 323
rect 462 318 463 322
rect 467 318 468 322
rect 462 317 468 318
rect 502 295 508 296
rect 502 291 503 295
rect 507 291 508 295
rect 502 290 508 291
rect 454 287 460 288
rect 454 283 455 287
rect 459 283 460 287
rect 454 282 460 283
rect 504 275 506 290
rect 111 274 115 275
rect 111 269 115 270
rect 287 274 291 275
rect 287 269 291 270
rect 359 274 363 275
rect 359 269 363 270
rect 439 274 443 275
rect 439 269 443 270
rect 447 274 451 275
rect 447 269 451 270
rect 503 274 507 275
rect 503 269 507 270
rect 112 257 114 269
rect 288 258 290 269
rect 342 259 348 260
rect 286 257 292 258
rect 110 256 116 257
rect 110 252 111 256
rect 115 252 116 256
rect 286 253 287 257
rect 291 253 292 257
rect 342 255 343 259
rect 347 255 348 259
rect 360 258 362 269
rect 430 259 436 260
rect 342 254 348 255
rect 358 257 364 258
rect 286 252 292 253
rect 110 251 116 252
rect 110 239 116 240
rect 110 235 111 239
rect 115 235 116 239
rect 110 234 116 235
rect 112 219 114 234
rect 302 230 308 231
rect 302 226 303 230
rect 307 226 308 230
rect 302 225 308 226
rect 304 219 306 225
rect 344 224 346 254
rect 358 253 359 257
rect 363 253 364 257
rect 430 255 431 259
rect 435 255 436 259
rect 440 258 442 269
rect 512 268 514 322
rect 518 318 519 322
rect 523 318 524 322
rect 518 317 524 318
rect 574 322 580 323
rect 594 322 600 323
rect 630 322 636 323
rect 650 322 656 323
rect 694 322 700 323
rect 574 318 575 322
rect 579 318 580 322
rect 574 317 580 318
rect 558 295 564 296
rect 558 291 559 295
rect 563 291 564 295
rect 596 292 598 322
rect 630 318 631 322
rect 635 318 636 322
rect 630 317 636 318
rect 614 295 620 296
rect 558 290 564 291
rect 594 291 600 292
rect 560 275 562 290
rect 594 287 595 291
rect 599 287 600 291
rect 614 291 615 295
rect 619 291 620 295
rect 652 292 654 322
rect 694 318 695 322
rect 699 318 700 322
rect 694 317 700 318
rect 766 322 772 323
rect 766 318 767 322
rect 771 318 772 322
rect 766 317 772 318
rect 846 322 852 323
rect 846 318 847 322
rect 851 318 852 322
rect 846 317 852 318
rect 678 295 684 296
rect 614 290 620 291
rect 650 291 656 292
rect 594 286 600 287
rect 616 275 618 290
rect 650 287 651 291
rect 655 287 656 291
rect 678 291 679 295
rect 683 291 684 295
rect 750 295 756 296
rect 678 290 684 291
rect 710 291 716 292
rect 650 286 656 287
rect 680 275 682 290
rect 710 287 711 291
rect 715 287 716 291
rect 750 291 751 295
rect 755 291 756 295
rect 750 290 756 291
rect 830 295 836 296
rect 830 291 831 295
rect 835 291 836 295
rect 856 292 858 338
rect 864 335 866 345
rect 936 344 938 382
rect 998 379 1004 380
rect 998 375 999 379
rect 1003 375 1004 379
rect 1008 378 1010 389
rect 1078 379 1084 380
rect 998 374 1004 375
rect 1006 377 1012 378
rect 942 350 948 351
rect 942 346 943 350
rect 947 346 948 350
rect 942 345 948 346
rect 934 343 940 344
rect 934 339 935 343
rect 939 339 940 343
rect 934 338 940 339
rect 934 335 940 336
rect 944 335 946 345
rect 1000 344 1002 374
rect 1006 373 1007 377
rect 1011 373 1012 377
rect 1078 375 1079 379
rect 1083 375 1084 379
rect 1088 378 1090 389
rect 1176 378 1178 389
rect 1078 374 1084 375
rect 1086 377 1092 378
rect 1006 372 1012 373
rect 1022 350 1028 351
rect 1022 346 1023 350
rect 1027 346 1028 350
rect 1022 345 1028 346
rect 998 343 1004 344
rect 998 339 999 343
rect 1003 339 1004 343
rect 998 338 1004 339
rect 1024 335 1026 345
rect 863 334 867 335
rect 863 329 867 330
rect 927 334 931 335
rect 934 331 935 335
rect 939 331 940 335
rect 934 330 940 331
rect 943 334 947 335
rect 927 329 931 330
rect 902 327 908 328
rect 902 323 903 327
rect 907 323 908 327
rect 928 323 930 329
rect 902 322 908 323
rect 926 322 932 323
rect 904 304 906 322
rect 926 318 927 322
rect 931 318 932 322
rect 926 317 932 318
rect 902 303 908 304
rect 902 299 903 303
rect 907 299 908 303
rect 902 298 908 299
rect 910 295 916 296
rect 830 290 836 291
rect 854 291 860 292
rect 710 286 716 287
rect 527 274 531 275
rect 527 269 531 270
rect 559 274 563 275
rect 559 269 563 270
rect 615 274 619 275
rect 615 269 619 270
rect 623 274 627 275
rect 623 269 627 270
rect 679 274 683 275
rect 679 269 683 270
rect 510 267 516 268
rect 510 263 511 267
rect 515 263 516 267
rect 510 262 516 263
rect 518 259 524 260
rect 430 254 436 255
rect 438 257 444 258
rect 358 252 364 253
rect 374 230 380 231
rect 374 226 375 230
rect 379 226 380 230
rect 374 225 380 226
rect 334 223 340 224
rect 334 219 335 223
rect 339 219 340 223
rect 111 218 115 219
rect 111 213 115 214
rect 199 218 203 219
rect 199 213 203 214
rect 271 218 275 219
rect 271 213 275 214
rect 303 218 307 219
rect 334 218 340 219
rect 342 223 348 224
rect 342 219 343 223
rect 347 219 348 223
rect 376 219 378 225
rect 432 224 434 254
rect 438 253 439 257
rect 443 253 444 257
rect 518 255 519 259
rect 523 255 524 259
rect 528 258 530 269
rect 614 259 620 260
rect 518 254 524 255
rect 526 257 532 258
rect 438 252 444 253
rect 454 230 460 231
rect 454 226 455 230
rect 459 226 460 230
rect 454 225 460 226
rect 430 223 436 224
rect 430 219 431 223
rect 435 219 436 223
rect 456 219 458 225
rect 520 224 522 254
rect 526 253 527 257
rect 531 253 532 257
rect 614 255 615 259
rect 619 255 620 259
rect 624 258 626 269
rect 614 254 620 255
rect 622 257 628 258
rect 526 252 532 253
rect 542 230 548 231
rect 542 226 543 230
rect 547 226 548 230
rect 542 225 548 226
rect 518 223 524 224
rect 518 219 519 223
rect 523 219 524 223
rect 544 219 546 225
rect 616 224 618 254
rect 622 253 623 257
rect 627 253 628 257
rect 622 252 628 253
rect 638 230 644 231
rect 638 226 639 230
rect 643 226 644 230
rect 638 225 644 226
rect 614 223 620 224
rect 614 219 615 223
rect 619 219 620 223
rect 640 219 642 225
rect 712 224 714 286
rect 752 275 754 290
rect 832 275 834 290
rect 854 287 855 291
rect 859 287 860 291
rect 910 291 911 295
rect 915 291 916 295
rect 936 292 938 330
rect 943 329 947 330
rect 1015 334 1019 335
rect 1015 329 1019 330
rect 1023 334 1027 335
rect 1023 329 1027 330
rect 962 327 968 328
rect 962 323 963 327
rect 967 323 968 327
rect 1016 323 1018 329
rect 1080 328 1082 374
rect 1086 373 1087 377
rect 1091 373 1092 377
rect 1086 372 1092 373
rect 1174 377 1180 378
rect 1174 373 1175 377
rect 1179 373 1180 377
rect 1174 372 1180 373
rect 1102 350 1108 351
rect 1102 346 1103 350
rect 1107 346 1108 350
rect 1102 345 1108 346
rect 1190 350 1196 351
rect 1190 346 1191 350
rect 1195 346 1196 350
rect 1190 345 1196 346
rect 1104 335 1106 345
rect 1192 335 1194 345
rect 1256 344 1258 406
rect 1328 395 1330 411
rect 1368 399 1370 411
rect 1630 410 1636 411
rect 1666 411 1672 412
rect 1632 399 1634 410
rect 1666 407 1667 411
rect 1671 407 1672 411
rect 1686 411 1687 415
rect 1691 411 1692 415
rect 1724 412 1726 442
rect 1758 438 1759 442
rect 1763 438 1764 442
rect 1758 437 1764 438
rect 1742 415 1748 416
rect 1686 410 1692 411
rect 1722 411 1728 412
rect 1666 406 1672 407
rect 1688 399 1690 410
rect 1722 407 1723 411
rect 1727 407 1728 411
rect 1742 411 1743 415
rect 1747 411 1748 415
rect 1776 412 1778 462
rect 1856 455 1858 469
rect 1920 468 1922 498
rect 1926 497 1927 501
rect 1931 497 1932 501
rect 1926 496 1932 497
rect 2014 501 2020 502
rect 2014 497 2015 501
rect 2019 497 2020 501
rect 2014 496 2020 497
rect 1942 474 1948 475
rect 1942 470 1943 474
rect 1947 470 1948 474
rect 1942 469 1948 470
rect 1918 467 1924 468
rect 1918 463 1919 467
rect 1923 463 1924 467
rect 1918 462 1924 463
rect 1886 455 1892 456
rect 1944 455 1946 469
rect 2024 468 2026 518
rect 2039 513 2043 514
rect 2095 518 2099 519
rect 2095 513 2099 514
rect 2135 518 2139 519
rect 2135 513 2139 514
rect 2175 518 2179 519
rect 2175 513 2179 514
rect 2223 518 2227 519
rect 2223 513 2227 514
rect 2255 518 2259 519
rect 2255 513 2259 514
rect 2303 518 2307 519
rect 2303 513 2307 514
rect 2327 518 2331 519
rect 2327 513 2331 514
rect 2383 518 2387 519
rect 2383 513 2387 514
rect 2399 518 2403 519
rect 2399 513 2403 514
rect 2086 503 2092 504
rect 2086 499 2087 503
rect 2091 499 2092 503
rect 2096 502 2098 513
rect 2166 503 2172 504
rect 2086 498 2092 499
rect 2094 501 2100 502
rect 2030 474 2036 475
rect 2030 470 2031 474
rect 2035 470 2036 474
rect 2030 469 2036 470
rect 2022 467 2028 468
rect 2022 463 2023 467
rect 2027 463 2028 467
rect 2022 462 2028 463
rect 2032 455 2034 469
rect 2088 468 2090 498
rect 2094 497 2095 501
rect 2099 497 2100 501
rect 2166 499 2167 503
rect 2171 499 2172 503
rect 2176 502 2178 513
rect 2198 503 2204 504
rect 2166 498 2172 499
rect 2174 501 2180 502
rect 2094 496 2100 497
rect 2110 474 2116 475
rect 2110 470 2111 474
rect 2115 470 2116 474
rect 2110 469 2116 470
rect 2086 467 2092 468
rect 2086 463 2087 467
rect 2091 463 2092 467
rect 2086 462 2092 463
rect 2112 455 2114 469
rect 2168 468 2170 498
rect 2174 497 2175 501
rect 2179 497 2180 501
rect 2198 499 2199 503
rect 2203 499 2204 503
rect 2256 502 2258 513
rect 2318 503 2324 504
rect 2198 498 2204 499
rect 2254 501 2260 502
rect 2174 496 2180 497
rect 2190 474 2196 475
rect 2190 470 2191 474
rect 2195 470 2196 474
rect 2190 469 2196 470
rect 2166 467 2172 468
rect 2166 463 2167 467
rect 2171 463 2172 467
rect 2166 462 2172 463
rect 2192 455 2194 469
rect 1815 454 1819 455
rect 1815 449 1819 450
rect 1855 454 1859 455
rect 1855 449 1859 450
rect 1871 454 1875 455
rect 1886 451 1887 455
rect 1891 451 1892 455
rect 1886 450 1892 451
rect 1927 454 1931 455
rect 1871 449 1875 450
rect 1816 443 1818 449
rect 1846 447 1852 448
rect 1846 443 1847 447
rect 1851 443 1852 447
rect 1872 443 1874 449
rect 1814 442 1820 443
rect 1846 442 1852 443
rect 1870 442 1876 443
rect 1814 438 1815 442
rect 1819 438 1820 442
rect 1814 437 1820 438
rect 1848 424 1850 442
rect 1870 438 1871 442
rect 1875 438 1876 442
rect 1870 437 1876 438
rect 1846 423 1852 424
rect 1846 419 1847 423
rect 1851 419 1852 423
rect 1846 418 1852 419
rect 1798 415 1804 416
rect 1742 410 1748 411
rect 1774 411 1780 412
rect 1722 406 1728 407
rect 1744 399 1746 410
rect 1774 407 1775 411
rect 1779 407 1780 411
rect 1798 411 1799 415
rect 1803 411 1804 415
rect 1798 410 1804 411
rect 1854 415 1860 416
rect 1854 411 1855 415
rect 1859 411 1860 415
rect 1888 412 1890 450
rect 1927 449 1931 450
rect 1943 454 1947 455
rect 1943 449 1947 450
rect 1999 454 2003 455
rect 1999 449 2003 450
rect 2031 454 2035 455
rect 2031 449 2035 450
rect 2087 454 2091 455
rect 2087 449 2091 450
rect 2111 454 2115 455
rect 2111 449 2115 450
rect 2191 454 2195 455
rect 2200 452 2202 498
rect 2254 497 2255 501
rect 2259 497 2260 501
rect 2318 499 2319 503
rect 2323 499 2324 503
rect 2328 502 2330 513
rect 2390 503 2396 504
rect 2318 498 2324 499
rect 2326 501 2332 502
rect 2254 496 2260 497
rect 2270 474 2276 475
rect 2270 470 2271 474
rect 2275 470 2276 474
rect 2270 469 2276 470
rect 2272 455 2274 469
rect 2320 468 2322 498
rect 2326 497 2327 501
rect 2331 497 2332 501
rect 2390 499 2391 503
rect 2395 499 2396 503
rect 2400 502 2402 513
rect 2436 504 2438 562
rect 2478 558 2479 562
rect 2483 558 2484 562
rect 2478 557 2484 558
rect 2462 535 2468 536
rect 2462 531 2463 535
rect 2467 531 2468 535
rect 2500 532 2502 562
rect 2542 558 2543 562
rect 2547 558 2548 562
rect 2542 557 2548 558
rect 2584 554 2586 569
rect 2582 553 2588 554
rect 2582 549 2583 553
rect 2587 549 2588 553
rect 2582 548 2588 549
rect 2582 536 2588 537
rect 2526 535 2532 536
rect 2462 530 2468 531
rect 2498 531 2504 532
rect 2464 519 2466 530
rect 2498 527 2499 531
rect 2503 527 2504 531
rect 2526 531 2527 535
rect 2531 531 2532 535
rect 2582 532 2583 536
rect 2587 532 2588 536
rect 2582 531 2588 532
rect 2526 530 2532 531
rect 2498 526 2504 527
rect 2528 519 2530 530
rect 2584 519 2586 531
rect 2463 518 2467 519
rect 2463 513 2467 514
rect 2471 518 2475 519
rect 2471 513 2475 514
rect 2527 518 2531 519
rect 2527 513 2531 514
rect 2583 518 2587 519
rect 2583 513 2587 514
rect 2434 503 2440 504
rect 2390 498 2396 499
rect 2398 501 2404 502
rect 2326 496 2332 497
rect 2342 474 2348 475
rect 2342 470 2343 474
rect 2347 470 2348 474
rect 2342 469 2348 470
rect 2318 467 2324 468
rect 2318 463 2319 467
rect 2323 463 2324 467
rect 2318 462 2324 463
rect 2344 455 2346 469
rect 2392 468 2394 498
rect 2398 497 2399 501
rect 2403 497 2404 501
rect 2434 499 2435 503
rect 2439 499 2440 503
rect 2472 502 2474 513
rect 2494 503 2500 504
rect 2434 498 2440 499
rect 2470 501 2476 502
rect 2398 496 2404 497
rect 2470 497 2471 501
rect 2475 497 2476 501
rect 2494 499 2495 503
rect 2499 499 2500 503
rect 2528 502 2530 513
rect 2494 498 2500 499
rect 2526 501 2532 502
rect 2584 501 2586 513
rect 2470 496 2476 497
rect 2414 474 2420 475
rect 2414 470 2415 474
rect 2419 470 2420 474
rect 2414 469 2420 470
rect 2486 474 2492 475
rect 2486 470 2487 474
rect 2491 470 2492 474
rect 2486 469 2492 470
rect 2390 467 2396 468
rect 2390 463 2391 467
rect 2395 463 2396 467
rect 2390 462 2396 463
rect 2416 455 2418 469
rect 2488 455 2490 469
rect 2496 460 2498 498
rect 2526 497 2527 501
rect 2531 497 2532 501
rect 2526 496 2532 497
rect 2582 500 2588 501
rect 2582 496 2583 500
rect 2587 496 2588 500
rect 2582 495 2588 496
rect 2582 483 2588 484
rect 2582 479 2583 483
rect 2587 479 2588 483
rect 2582 478 2588 479
rect 2542 474 2548 475
rect 2542 470 2543 474
rect 2547 470 2548 474
rect 2542 469 2548 470
rect 2494 459 2500 460
rect 2494 455 2495 459
rect 2499 455 2500 459
rect 2544 455 2546 469
rect 2558 467 2564 468
rect 2558 463 2559 467
rect 2563 463 2564 467
rect 2558 462 2564 463
rect 2271 454 2275 455
rect 2191 449 2195 450
rect 2198 451 2204 452
rect 1918 447 1924 448
rect 1918 443 1919 447
rect 1923 443 1924 447
rect 1928 443 1930 449
rect 1974 447 1980 448
rect 1974 443 1975 447
rect 1979 443 1980 447
rect 2000 443 2002 449
rect 2078 447 2084 448
rect 2078 443 2079 447
rect 2083 443 2084 447
rect 2088 443 2090 449
rect 2192 443 2194 449
rect 2198 447 2199 451
rect 2203 447 2204 451
rect 2271 449 2275 450
rect 2311 454 2315 455
rect 2311 449 2315 450
rect 2343 454 2347 455
rect 2343 449 2347 450
rect 2415 454 2419 455
rect 2415 449 2419 450
rect 2439 454 2443 455
rect 2439 449 2443 450
rect 2487 454 2491 455
rect 2494 454 2500 455
rect 2543 454 2547 455
rect 2487 449 2491 450
rect 2543 449 2547 450
rect 2198 446 2204 447
rect 2210 447 2216 448
rect 2210 443 2211 447
rect 2215 443 2216 447
rect 2312 443 2314 449
rect 2330 447 2336 448
rect 2330 443 2331 447
rect 2335 443 2336 447
rect 2440 443 2442 449
rect 2534 447 2540 448
rect 2534 443 2535 447
rect 2539 443 2540 447
rect 2544 443 2546 449
rect 1918 442 1924 443
rect 1926 442 1932 443
rect 1974 442 1980 443
rect 1998 442 2004 443
rect 2078 442 2084 443
rect 2086 442 2092 443
rect 1910 415 1916 416
rect 1854 410 1860 411
rect 1886 411 1892 412
rect 1774 406 1780 407
rect 1800 399 1802 410
rect 1856 399 1858 410
rect 1886 407 1887 411
rect 1891 407 1892 411
rect 1910 411 1911 415
rect 1915 411 1916 415
rect 1910 410 1916 411
rect 1886 406 1892 407
rect 1912 399 1914 410
rect 1367 398 1371 399
rect 1263 394 1267 395
rect 1263 389 1267 390
rect 1327 394 1331 395
rect 1367 393 1371 394
rect 1631 398 1635 399
rect 1631 393 1635 394
rect 1655 398 1659 399
rect 1655 393 1659 394
rect 1687 398 1691 399
rect 1687 393 1691 394
rect 1711 398 1715 399
rect 1711 393 1715 394
rect 1743 398 1747 399
rect 1743 393 1747 394
rect 1767 398 1771 399
rect 1767 393 1771 394
rect 1799 398 1803 399
rect 1799 393 1803 394
rect 1823 398 1827 399
rect 1823 393 1827 394
rect 1855 398 1859 399
rect 1855 393 1859 394
rect 1879 398 1883 399
rect 1879 393 1883 394
rect 1911 398 1915 399
rect 1911 393 1915 394
rect 1327 389 1331 390
rect 1264 378 1266 389
rect 1262 377 1268 378
rect 1328 377 1330 389
rect 1368 381 1370 393
rect 1656 382 1658 393
rect 1702 383 1708 384
rect 1654 381 1660 382
rect 1366 380 1372 381
rect 1262 373 1263 377
rect 1267 373 1268 377
rect 1262 372 1268 373
rect 1326 376 1332 377
rect 1326 372 1327 376
rect 1331 372 1332 376
rect 1366 376 1367 380
rect 1371 376 1372 380
rect 1654 377 1655 381
rect 1659 377 1660 381
rect 1702 379 1703 383
rect 1707 379 1708 383
rect 1712 382 1714 393
rect 1758 383 1764 384
rect 1702 378 1708 379
rect 1710 381 1716 382
rect 1654 376 1660 377
rect 1366 375 1372 376
rect 1326 371 1332 372
rect 1366 363 1372 364
rect 1326 359 1332 360
rect 1326 355 1327 359
rect 1331 355 1332 359
rect 1366 359 1367 363
rect 1371 359 1372 363
rect 1366 358 1372 359
rect 1326 354 1332 355
rect 1278 350 1284 351
rect 1278 346 1279 350
rect 1283 346 1284 350
rect 1278 345 1284 346
rect 1254 343 1260 344
rect 1254 339 1255 343
rect 1259 339 1260 343
rect 1254 338 1260 339
rect 1280 335 1282 345
rect 1328 335 1330 354
rect 1368 335 1370 358
rect 1670 354 1676 355
rect 1670 350 1671 354
rect 1675 350 1676 354
rect 1670 349 1676 350
rect 1672 335 1674 349
rect 1704 348 1706 378
rect 1710 377 1711 381
rect 1715 377 1716 381
rect 1758 379 1759 383
rect 1763 379 1764 383
rect 1768 382 1770 393
rect 1814 383 1820 384
rect 1758 378 1764 379
rect 1766 381 1772 382
rect 1710 376 1716 377
rect 1726 354 1732 355
rect 1726 350 1727 354
rect 1731 350 1732 354
rect 1726 349 1732 350
rect 1702 347 1708 348
rect 1702 343 1703 347
rect 1707 343 1708 347
rect 1702 342 1708 343
rect 1728 335 1730 349
rect 1760 348 1762 378
rect 1766 377 1767 381
rect 1771 377 1772 381
rect 1814 379 1815 383
rect 1819 379 1820 383
rect 1824 382 1826 393
rect 1870 383 1876 384
rect 1814 378 1820 379
rect 1822 381 1828 382
rect 1766 376 1772 377
rect 1782 354 1788 355
rect 1782 350 1783 354
rect 1787 350 1788 354
rect 1782 349 1788 350
rect 1758 347 1764 348
rect 1758 343 1759 347
rect 1763 343 1764 347
rect 1758 342 1764 343
rect 1784 335 1786 349
rect 1816 348 1818 378
rect 1822 377 1823 381
rect 1827 377 1828 381
rect 1870 379 1871 383
rect 1875 379 1876 383
rect 1880 382 1882 393
rect 1920 392 1922 442
rect 1926 438 1927 442
rect 1931 438 1932 442
rect 1926 437 1932 438
rect 1976 424 1978 442
rect 1998 438 1999 442
rect 2003 438 2004 442
rect 1998 437 2004 438
rect 1974 423 1980 424
rect 1974 419 1975 423
rect 1979 419 1980 423
rect 2080 421 2082 442
rect 2086 438 2087 442
rect 2091 438 2092 442
rect 2086 437 2092 438
rect 2190 442 2196 443
rect 2210 442 2216 443
rect 2310 442 2316 443
rect 2330 442 2336 443
rect 2438 442 2444 443
rect 2534 442 2540 443
rect 2542 442 2548 443
rect 2190 438 2191 442
rect 2195 438 2196 442
rect 2190 437 2196 438
rect 1974 418 1980 419
rect 2079 420 2083 421
rect 1982 415 1988 416
rect 1982 411 1983 415
rect 1987 411 1988 415
rect 2070 415 2076 416
rect 2079 415 2083 416
rect 2174 415 2180 416
rect 1982 410 1988 411
rect 2018 411 2024 412
rect 1984 399 1986 410
rect 2018 407 2019 411
rect 2023 407 2024 411
rect 2070 411 2071 415
rect 2075 411 2076 415
rect 2070 410 2076 411
rect 2174 411 2175 415
rect 2179 411 2180 415
rect 2212 412 2214 442
rect 2310 438 2311 442
rect 2315 438 2316 442
rect 2310 437 2316 438
rect 2294 415 2300 416
rect 2174 410 2180 411
rect 2210 411 2216 412
rect 2018 406 2024 407
rect 1951 398 1955 399
rect 1951 393 1955 394
rect 1983 398 1987 399
rect 1983 393 1987 394
rect 1918 391 1924 392
rect 1918 387 1919 391
rect 1923 387 1924 391
rect 1918 386 1924 387
rect 1942 383 1948 384
rect 1870 378 1876 379
rect 1878 381 1884 382
rect 1822 376 1828 377
rect 1838 354 1844 355
rect 1838 350 1839 354
rect 1843 350 1844 354
rect 1838 349 1844 350
rect 1814 347 1820 348
rect 1814 343 1815 347
rect 1819 343 1820 347
rect 1814 342 1820 343
rect 1840 335 1842 349
rect 1872 348 1874 378
rect 1878 377 1879 381
rect 1883 377 1884 381
rect 1942 379 1943 383
rect 1947 379 1948 383
rect 1952 382 1954 393
rect 1942 378 1948 379
rect 1950 381 1956 382
rect 1878 376 1884 377
rect 1894 354 1900 355
rect 1894 350 1895 354
rect 1899 350 1900 354
rect 1894 349 1900 350
rect 1870 347 1876 348
rect 1870 343 1871 347
rect 1875 343 1876 347
rect 1870 342 1876 343
rect 1896 335 1898 349
rect 1944 348 1946 378
rect 1950 377 1951 381
rect 1955 377 1956 381
rect 1950 376 1956 377
rect 1966 354 1972 355
rect 1966 350 1967 354
rect 1971 350 1972 354
rect 1966 349 1972 350
rect 1942 347 1948 348
rect 1942 343 1943 347
rect 1947 343 1948 347
rect 1942 342 1948 343
rect 1968 335 1970 349
rect 2020 348 2022 406
rect 2072 399 2074 410
rect 2176 399 2178 410
rect 2210 407 2211 411
rect 2215 407 2216 411
rect 2294 411 2295 415
rect 2299 411 2300 415
rect 2332 412 2334 442
rect 2438 438 2439 442
rect 2443 438 2444 442
rect 2438 437 2444 438
rect 2455 420 2459 421
rect 2422 415 2428 416
rect 2455 415 2459 416
rect 2526 415 2532 416
rect 2294 410 2300 411
rect 2330 411 2336 412
rect 2210 406 2216 407
rect 2296 399 2298 410
rect 2330 407 2331 411
rect 2335 407 2336 411
rect 2422 411 2423 415
rect 2427 411 2428 415
rect 2456 412 2458 415
rect 2422 410 2428 411
rect 2454 411 2460 412
rect 2330 406 2336 407
rect 2424 399 2426 410
rect 2454 407 2455 411
rect 2459 407 2460 411
rect 2526 411 2527 415
rect 2531 411 2532 415
rect 2526 410 2532 411
rect 2454 406 2460 407
rect 2528 399 2530 410
rect 2039 398 2043 399
rect 2039 393 2043 394
rect 2071 398 2075 399
rect 2071 393 2075 394
rect 2151 398 2155 399
rect 2151 393 2155 394
rect 2175 398 2179 399
rect 2175 393 2179 394
rect 2279 398 2283 399
rect 2279 393 2283 394
rect 2295 398 2299 399
rect 2295 393 2299 394
rect 2415 398 2419 399
rect 2415 393 2419 394
rect 2423 398 2427 399
rect 2423 393 2427 394
rect 2527 398 2531 399
rect 2527 393 2531 394
rect 2040 382 2042 393
rect 2142 383 2148 384
rect 2038 381 2044 382
rect 2038 377 2039 381
rect 2043 377 2044 381
rect 2142 379 2143 383
rect 2147 379 2148 383
rect 2152 382 2154 393
rect 2270 383 2276 384
rect 2142 378 2148 379
rect 2150 381 2156 382
rect 2038 376 2044 377
rect 2123 356 2127 357
rect 2054 354 2060 355
rect 2054 350 2055 354
rect 2059 350 2060 354
rect 2123 351 2127 352
rect 2054 349 2060 350
rect 2018 347 2024 348
rect 2018 343 2019 347
rect 2023 343 2024 347
rect 2018 342 2024 343
rect 1982 339 1988 340
rect 1982 335 1983 339
rect 1987 335 1988 339
rect 2056 335 2058 349
rect 1103 334 1107 335
rect 1103 329 1107 330
rect 1111 334 1115 335
rect 1111 329 1115 330
rect 1191 334 1195 335
rect 1191 329 1195 330
rect 1215 334 1219 335
rect 1215 329 1219 330
rect 1279 334 1283 335
rect 1279 329 1283 330
rect 1327 334 1331 335
rect 1327 329 1331 330
rect 1367 334 1371 335
rect 1367 329 1371 330
rect 1631 334 1635 335
rect 1631 329 1635 330
rect 1671 334 1675 335
rect 1671 329 1675 330
rect 1687 334 1691 335
rect 1687 329 1691 330
rect 1727 334 1731 335
rect 1727 329 1731 330
rect 1743 334 1747 335
rect 1743 329 1747 330
rect 1783 334 1787 335
rect 1783 329 1787 330
rect 1807 334 1811 335
rect 1807 329 1811 330
rect 1839 334 1843 335
rect 1839 329 1843 330
rect 1887 334 1891 335
rect 1887 329 1891 330
rect 1895 334 1899 335
rect 1895 329 1899 330
rect 1967 334 1971 335
rect 1982 334 1988 335
rect 2055 334 2059 335
rect 1967 329 1971 330
rect 1078 327 1084 328
rect 1078 323 1079 327
rect 1083 323 1084 327
rect 1112 323 1114 329
rect 1130 327 1136 328
rect 1130 323 1131 327
rect 1135 323 1136 327
rect 1216 323 1218 329
rect 962 322 968 323
rect 1014 322 1020 323
rect 1078 322 1084 323
rect 1110 322 1116 323
rect 1130 322 1136 323
rect 1214 322 1220 323
rect 910 290 916 291
rect 934 291 940 292
rect 854 286 860 287
rect 912 275 914 290
rect 934 287 935 291
rect 939 287 940 291
rect 934 286 940 287
rect 719 274 723 275
rect 719 269 723 270
rect 751 274 755 275
rect 751 269 755 270
rect 823 274 827 275
rect 823 269 827 270
rect 831 274 835 275
rect 831 269 835 270
rect 911 274 915 275
rect 911 269 915 270
rect 927 274 931 275
rect 927 269 931 270
rect 720 258 722 269
rect 766 259 772 260
rect 718 257 724 258
rect 718 253 719 257
rect 723 253 724 257
rect 766 255 767 259
rect 771 255 772 259
rect 824 258 826 269
rect 846 267 852 268
rect 846 263 847 267
rect 851 263 852 267
rect 846 262 852 263
rect 766 254 772 255
rect 822 257 828 258
rect 718 252 724 253
rect 734 230 740 231
rect 734 226 735 230
rect 739 226 740 230
rect 734 225 740 226
rect 710 223 716 224
rect 710 219 711 223
rect 715 219 716 223
rect 736 219 738 225
rect 342 218 348 219
rect 359 218 363 219
rect 303 213 307 214
rect 112 198 114 213
rect 190 211 196 212
rect 190 207 191 211
rect 195 207 196 211
rect 200 207 202 213
rect 218 211 224 212
rect 218 207 219 211
rect 223 207 224 211
rect 272 207 274 213
rect 290 211 296 212
rect 290 207 291 211
rect 295 207 296 211
rect 190 206 196 207
rect 198 206 204 207
rect 218 206 224 207
rect 270 206 276 207
rect 290 206 296 207
rect 110 197 116 198
rect 110 193 111 197
rect 115 193 116 197
rect 110 192 116 193
rect 110 180 116 181
rect 110 176 111 180
rect 115 176 116 180
rect 110 175 116 176
rect 182 179 188 180
rect 182 175 183 179
rect 187 175 188 179
rect 112 139 114 175
rect 182 174 188 175
rect 184 139 186 174
rect 192 165 194 206
rect 198 202 199 206
rect 203 202 204 206
rect 198 201 204 202
rect 220 176 222 206
rect 270 202 271 206
rect 275 202 276 206
rect 270 201 276 202
rect 254 179 260 180
rect 218 175 224 176
rect 218 171 219 175
rect 223 171 224 175
rect 254 175 255 179
rect 259 175 260 179
rect 292 176 294 206
rect 336 188 338 218
rect 359 213 363 214
rect 375 218 379 219
rect 430 218 436 219
rect 455 218 459 219
rect 375 213 379 214
rect 455 213 459 214
rect 463 218 467 219
rect 518 218 524 219
rect 543 218 547 219
rect 463 213 467 214
rect 543 213 547 214
rect 567 218 571 219
rect 614 218 620 219
rect 639 218 643 219
rect 567 213 571 214
rect 639 213 643 214
rect 679 218 683 219
rect 710 218 716 219
rect 735 218 739 219
rect 679 213 683 214
rect 735 213 739 214
rect 360 207 362 213
rect 464 207 466 213
rect 482 211 488 212
rect 482 207 483 211
rect 487 207 488 211
rect 568 207 570 213
rect 654 211 660 212
rect 654 207 655 211
rect 659 207 660 211
rect 680 207 682 213
rect 768 212 770 254
rect 822 253 823 257
rect 827 253 828 257
rect 822 252 828 253
rect 838 230 844 231
rect 838 226 839 230
rect 843 226 844 230
rect 838 225 844 226
rect 840 219 842 225
rect 848 224 850 262
rect 918 259 924 260
rect 918 255 919 259
rect 923 255 924 259
rect 928 258 930 269
rect 964 260 966 322
rect 1014 318 1015 322
rect 1019 318 1020 322
rect 1014 317 1020 318
rect 1110 318 1111 322
rect 1115 318 1116 322
rect 1110 317 1116 318
rect 998 295 1004 296
rect 998 291 999 295
rect 1003 291 1004 295
rect 998 290 1004 291
rect 1094 295 1100 296
rect 1094 291 1095 295
rect 1099 291 1100 295
rect 1132 292 1134 322
rect 1214 318 1215 322
rect 1219 318 1220 322
rect 1214 317 1220 318
rect 1328 314 1330 329
rect 1368 314 1370 329
rect 1622 327 1628 328
rect 1622 323 1623 327
rect 1627 323 1628 327
rect 1632 323 1634 329
rect 1650 327 1656 328
rect 1650 323 1651 327
rect 1655 323 1656 327
rect 1688 323 1690 329
rect 1706 327 1712 328
rect 1706 323 1707 327
rect 1711 323 1712 327
rect 1744 323 1746 329
rect 1762 327 1768 328
rect 1762 323 1763 327
rect 1767 323 1768 327
rect 1808 323 1810 329
rect 1826 327 1832 328
rect 1826 323 1827 327
rect 1831 323 1832 327
rect 1888 323 1890 329
rect 1906 327 1912 328
rect 1906 323 1907 327
rect 1911 323 1912 327
rect 1968 323 1970 329
rect 1622 322 1628 323
rect 1630 322 1636 323
rect 1650 322 1656 323
rect 1686 322 1692 323
rect 1706 322 1712 323
rect 1742 322 1748 323
rect 1762 322 1768 323
rect 1806 322 1812 323
rect 1826 322 1832 323
rect 1886 322 1892 323
rect 1906 322 1912 323
rect 1966 322 1972 323
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1326 308 1332 309
rect 1366 313 1372 314
rect 1366 309 1367 313
rect 1371 309 1372 313
rect 1366 308 1372 309
rect 1326 296 1332 297
rect 1198 295 1204 296
rect 1094 290 1100 291
rect 1130 291 1136 292
rect 1000 275 1002 290
rect 1096 275 1098 290
rect 1130 287 1131 291
rect 1135 287 1136 291
rect 1198 291 1199 295
rect 1203 291 1204 295
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1198 290 1204 291
rect 1222 291 1228 292
rect 1326 291 1332 292
rect 1366 296 1372 297
rect 1366 292 1367 296
rect 1371 292 1372 296
rect 1366 291 1372 292
rect 1614 295 1620 296
rect 1614 291 1615 295
rect 1619 291 1620 295
rect 1130 286 1136 287
rect 1200 275 1202 290
rect 1222 287 1223 291
rect 1227 287 1228 291
rect 1222 286 1228 287
rect 999 274 1003 275
rect 999 269 1003 270
rect 1031 274 1035 275
rect 1031 269 1035 270
rect 1095 274 1099 275
rect 1095 269 1099 270
rect 1143 274 1147 275
rect 1143 269 1147 270
rect 1199 274 1203 275
rect 1199 269 1203 270
rect 962 259 968 260
rect 918 254 924 255
rect 926 257 932 258
rect 920 224 922 254
rect 926 253 927 257
rect 931 253 932 257
rect 962 255 963 259
rect 967 255 968 259
rect 1032 258 1034 269
rect 1144 258 1146 269
rect 962 254 968 255
rect 1030 257 1036 258
rect 926 252 932 253
rect 1030 253 1031 257
rect 1035 253 1036 257
rect 1030 252 1036 253
rect 1142 257 1148 258
rect 1142 253 1143 257
rect 1147 253 1148 257
rect 1142 252 1148 253
rect 942 230 948 231
rect 942 226 943 230
rect 947 226 948 230
rect 942 225 948 226
rect 1046 230 1052 231
rect 1046 226 1047 230
rect 1051 226 1052 230
rect 1046 225 1052 226
rect 1158 230 1164 231
rect 1158 226 1159 230
rect 1163 226 1164 230
rect 1158 225 1164 226
rect 846 223 852 224
rect 846 219 847 223
rect 851 219 852 223
rect 918 223 924 224
rect 918 219 919 223
rect 923 219 924 223
rect 944 219 946 225
rect 1038 223 1044 224
rect 1038 219 1039 223
rect 1043 219 1044 223
rect 1048 219 1050 225
rect 1160 219 1162 225
rect 1224 224 1226 286
rect 1328 275 1330 291
rect 1368 279 1370 291
rect 1614 290 1620 291
rect 1616 279 1618 290
rect 1367 278 1371 279
rect 1255 274 1259 275
rect 1255 269 1259 270
rect 1327 274 1331 275
rect 1367 273 1371 274
rect 1535 278 1539 279
rect 1535 273 1539 274
rect 1607 278 1611 279
rect 1607 273 1611 274
rect 1615 278 1619 279
rect 1615 273 1619 274
rect 1327 269 1331 270
rect 1246 259 1252 260
rect 1246 255 1247 259
rect 1251 255 1252 259
rect 1256 258 1258 269
rect 1278 259 1284 260
rect 1246 254 1252 255
rect 1254 257 1260 258
rect 1248 224 1250 254
rect 1254 253 1255 257
rect 1259 253 1260 257
rect 1278 255 1279 259
rect 1283 255 1284 259
rect 1328 257 1330 269
rect 1368 261 1370 273
rect 1536 262 1538 273
rect 1598 263 1604 264
rect 1534 261 1540 262
rect 1366 260 1372 261
rect 1278 254 1284 255
rect 1326 256 1332 257
rect 1254 252 1260 253
rect 1270 230 1276 231
rect 1270 226 1271 230
rect 1275 226 1276 230
rect 1270 225 1276 226
rect 1222 223 1228 224
rect 1222 219 1223 223
rect 1227 219 1228 223
rect 791 218 795 219
rect 791 213 795 214
rect 839 218 843 219
rect 846 218 852 219
rect 911 218 915 219
rect 918 218 924 219
rect 943 218 947 219
rect 839 213 843 214
rect 911 213 915 214
rect 943 213 947 214
rect 1031 218 1035 219
rect 1038 218 1044 219
rect 1047 218 1051 219
rect 1031 213 1035 214
rect 766 211 772 212
rect 766 207 767 211
rect 771 207 772 211
rect 792 207 794 213
rect 886 211 892 212
rect 886 207 887 211
rect 891 207 892 211
rect 912 207 914 213
rect 930 211 936 212
rect 930 207 931 211
rect 935 207 936 211
rect 1032 207 1034 213
rect 358 206 364 207
rect 358 202 359 206
rect 363 202 364 206
rect 358 201 364 202
rect 462 206 468 207
rect 482 206 488 207
rect 566 206 572 207
rect 654 206 660 207
rect 678 206 684 207
rect 766 206 772 207
rect 790 206 796 207
rect 886 206 892 207
rect 910 206 916 207
rect 930 206 936 207
rect 1030 206 1036 207
rect 462 202 463 206
rect 467 202 468 206
rect 462 201 468 202
rect 334 187 340 188
rect 334 183 335 187
rect 339 183 340 187
rect 334 182 340 183
rect 342 179 348 180
rect 254 174 260 175
rect 290 175 296 176
rect 218 170 224 171
rect 191 164 195 165
rect 191 159 195 160
rect 256 139 258 174
rect 290 171 291 175
rect 295 171 296 175
rect 342 175 343 179
rect 347 175 348 179
rect 342 174 348 175
rect 446 179 452 180
rect 446 175 447 179
rect 451 175 452 179
rect 484 176 486 206
rect 566 202 567 206
rect 571 202 572 206
rect 566 201 572 202
rect 656 188 658 206
rect 678 202 679 206
rect 683 202 684 206
rect 678 201 684 202
rect 790 202 791 206
rect 795 202 796 206
rect 790 201 796 202
rect 888 188 890 206
rect 910 202 911 206
rect 915 202 916 206
rect 910 201 916 202
rect 654 187 660 188
rect 654 183 655 187
rect 659 183 660 187
rect 654 182 660 183
rect 886 187 892 188
rect 886 183 887 187
rect 891 183 892 187
rect 886 182 892 183
rect 550 179 556 180
rect 446 174 452 175
rect 482 175 488 176
rect 290 170 296 171
rect 344 139 346 174
rect 448 139 450 174
rect 482 171 483 175
rect 487 171 488 175
rect 550 175 551 179
rect 555 175 556 179
rect 550 174 556 175
rect 662 179 668 180
rect 662 175 663 179
rect 667 175 668 179
rect 774 179 780 180
rect 662 174 668 175
rect 686 175 692 176
rect 482 170 488 171
rect 552 139 554 174
rect 623 164 627 165
rect 623 159 627 160
rect 111 138 115 139
rect 111 133 115 134
rect 143 138 147 139
rect 143 133 147 134
rect 183 138 187 139
rect 183 133 187 134
rect 199 138 203 139
rect 199 133 203 134
rect 255 138 259 139
rect 255 133 259 134
rect 311 138 315 139
rect 311 133 315 134
rect 343 138 347 139
rect 343 133 347 134
rect 367 138 371 139
rect 367 133 371 134
rect 423 138 427 139
rect 423 133 427 134
rect 447 138 451 139
rect 447 133 451 134
rect 479 138 483 139
rect 479 133 483 134
rect 535 138 539 139
rect 535 133 539 134
rect 551 138 555 139
rect 551 133 555 134
rect 591 138 595 139
rect 591 133 595 134
rect 112 121 114 133
rect 144 122 146 133
rect 190 123 196 124
rect 142 121 148 122
rect 110 120 116 121
rect 110 116 111 120
rect 115 116 116 120
rect 142 117 143 121
rect 147 117 148 121
rect 190 119 191 123
rect 195 119 196 123
rect 200 122 202 133
rect 246 123 252 124
rect 190 118 196 119
rect 198 121 204 122
rect 142 116 148 117
rect 110 115 116 116
rect 110 103 116 104
rect 110 99 111 103
rect 115 99 116 103
rect 110 98 116 99
rect 112 83 114 98
rect 158 94 164 95
rect 158 90 159 94
rect 163 90 164 94
rect 158 89 164 90
rect 160 83 162 89
rect 192 88 194 118
rect 198 117 199 121
rect 203 117 204 121
rect 246 119 247 123
rect 251 119 252 123
rect 256 122 258 133
rect 302 123 308 124
rect 246 118 252 119
rect 254 121 260 122
rect 198 116 204 117
rect 214 94 220 95
rect 214 90 215 94
rect 219 90 220 94
rect 214 89 220 90
rect 190 87 196 88
rect 190 83 191 87
rect 195 83 196 87
rect 216 83 218 89
rect 248 88 250 118
rect 254 117 255 121
rect 259 117 260 121
rect 302 119 303 123
rect 307 119 308 123
rect 312 122 314 133
rect 358 123 364 124
rect 302 118 308 119
rect 310 121 316 122
rect 254 116 260 117
rect 270 94 276 95
rect 270 90 271 94
rect 275 90 276 94
rect 270 89 276 90
rect 246 87 252 88
rect 246 83 247 87
rect 251 83 252 87
rect 272 83 274 89
rect 304 88 306 118
rect 310 117 311 121
rect 315 117 316 121
rect 358 119 359 123
rect 363 119 364 123
rect 368 122 370 133
rect 414 123 420 124
rect 358 118 364 119
rect 366 121 372 122
rect 310 116 316 117
rect 326 94 332 95
rect 326 90 327 94
rect 331 90 332 94
rect 326 89 332 90
rect 302 87 308 88
rect 302 83 303 87
rect 307 83 308 87
rect 328 83 330 89
rect 360 88 362 118
rect 366 117 367 121
rect 371 117 372 121
rect 414 119 415 123
rect 419 119 420 123
rect 424 122 426 133
rect 470 123 476 124
rect 414 118 420 119
rect 422 121 428 122
rect 366 116 372 117
rect 382 94 388 95
rect 382 90 383 94
rect 387 90 388 94
rect 382 89 388 90
rect 358 87 364 88
rect 358 83 359 87
rect 363 83 364 87
rect 384 83 386 89
rect 416 88 418 118
rect 422 117 423 121
rect 427 117 428 121
rect 470 119 471 123
rect 475 119 476 123
rect 480 122 482 133
rect 526 123 532 124
rect 470 118 476 119
rect 478 121 484 122
rect 422 116 428 117
rect 438 94 444 95
rect 438 90 439 94
rect 443 90 444 94
rect 438 89 444 90
rect 414 87 420 88
rect 414 83 415 87
rect 419 83 420 87
rect 440 83 442 89
rect 472 88 474 118
rect 478 117 479 121
rect 483 117 484 121
rect 526 119 527 123
rect 531 119 532 123
rect 536 122 538 133
rect 582 123 588 124
rect 526 118 532 119
rect 534 121 540 122
rect 478 116 484 117
rect 494 94 500 95
rect 494 90 495 94
rect 499 90 500 94
rect 494 89 500 90
rect 470 87 476 88
rect 470 83 471 87
rect 475 83 476 87
rect 496 83 498 89
rect 528 88 530 118
rect 534 117 535 121
rect 539 117 540 121
rect 582 119 583 123
rect 587 119 588 123
rect 592 122 594 133
rect 624 124 626 159
rect 664 139 666 174
rect 686 171 687 175
rect 691 171 692 175
rect 774 175 775 179
rect 779 175 780 179
rect 774 174 780 175
rect 894 179 900 180
rect 894 175 895 179
rect 899 175 900 179
rect 932 176 934 206
rect 1030 202 1031 206
rect 1035 202 1036 206
rect 1030 201 1036 202
rect 1014 179 1020 180
rect 894 174 900 175
rect 930 175 936 176
rect 686 170 692 171
rect 647 138 651 139
rect 647 133 651 134
rect 663 138 667 139
rect 663 133 667 134
rect 622 123 628 124
rect 582 118 588 119
rect 590 121 596 122
rect 534 116 540 117
rect 550 94 556 95
rect 550 90 551 94
rect 555 90 556 94
rect 550 89 556 90
rect 526 87 532 88
rect 526 83 527 87
rect 531 83 532 87
rect 552 83 554 89
rect 584 88 586 118
rect 590 117 591 121
rect 595 117 596 121
rect 622 119 623 123
rect 627 119 628 123
rect 648 122 650 133
rect 622 118 628 119
rect 646 121 652 122
rect 590 116 596 117
rect 646 117 647 121
rect 651 117 652 121
rect 646 116 652 117
rect 606 94 612 95
rect 606 90 607 94
rect 611 90 612 94
rect 606 89 612 90
rect 662 94 668 95
rect 662 90 663 94
rect 667 90 668 94
rect 662 89 668 90
rect 582 87 588 88
rect 582 83 583 87
rect 587 83 588 87
rect 608 83 610 89
rect 664 83 666 89
rect 688 88 690 170
rect 776 139 778 174
rect 896 139 898 174
rect 930 171 931 175
rect 935 171 936 175
rect 1014 175 1015 179
rect 1019 175 1020 179
rect 1040 176 1042 218
rect 1047 213 1051 214
rect 1151 218 1155 219
rect 1151 213 1155 214
rect 1159 218 1163 219
rect 1222 218 1228 219
rect 1246 223 1252 224
rect 1246 219 1247 223
rect 1251 219 1252 223
rect 1272 219 1274 225
rect 1246 218 1252 219
rect 1271 218 1275 219
rect 1159 213 1163 214
rect 1280 216 1282 254
rect 1326 252 1327 256
rect 1331 252 1332 256
rect 1366 256 1367 260
rect 1371 256 1372 260
rect 1534 257 1535 261
rect 1539 257 1540 261
rect 1598 259 1599 263
rect 1603 259 1604 263
rect 1608 262 1610 273
rect 1624 272 1626 322
rect 1630 318 1631 322
rect 1635 318 1636 322
rect 1630 317 1636 318
rect 1652 292 1654 322
rect 1686 318 1687 322
rect 1691 318 1692 322
rect 1686 317 1692 318
rect 1670 295 1676 296
rect 1650 291 1656 292
rect 1650 287 1651 291
rect 1655 287 1656 291
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1708 292 1710 322
rect 1742 318 1743 322
rect 1747 318 1748 322
rect 1742 317 1748 318
rect 1726 295 1732 296
rect 1670 290 1676 291
rect 1706 291 1712 292
rect 1650 286 1656 287
rect 1672 279 1674 290
rect 1706 287 1707 291
rect 1711 287 1712 291
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1764 292 1766 322
rect 1806 318 1807 322
rect 1811 318 1812 322
rect 1806 317 1812 318
rect 1790 295 1796 296
rect 1726 290 1732 291
rect 1762 291 1768 292
rect 1706 286 1712 287
rect 1728 279 1730 290
rect 1762 287 1763 291
rect 1767 287 1768 291
rect 1790 291 1791 295
rect 1795 291 1796 295
rect 1828 292 1830 322
rect 1886 318 1887 322
rect 1891 318 1892 322
rect 1886 317 1892 318
rect 1870 295 1876 296
rect 1790 290 1796 291
rect 1826 291 1832 292
rect 1762 286 1768 287
rect 1792 279 1794 290
rect 1826 287 1827 291
rect 1831 287 1832 291
rect 1870 291 1871 295
rect 1875 291 1876 295
rect 1908 292 1910 322
rect 1966 318 1967 322
rect 1971 318 1972 322
rect 1966 317 1972 318
rect 1950 295 1956 296
rect 1870 290 1876 291
rect 1906 291 1912 292
rect 1826 286 1832 287
rect 1872 279 1874 290
rect 1906 287 1907 291
rect 1911 287 1912 291
rect 1950 291 1951 295
rect 1955 291 1956 295
rect 1984 292 1986 334
rect 2055 329 2059 330
rect 2030 327 2036 328
rect 2030 323 2031 327
rect 2035 323 2036 327
rect 2056 323 2058 329
rect 2124 328 2126 351
rect 2144 348 2146 378
rect 2150 377 2151 381
rect 2155 377 2156 381
rect 2270 379 2271 383
rect 2275 379 2276 383
rect 2280 382 2282 393
rect 2406 383 2412 384
rect 2270 378 2276 379
rect 2278 381 2284 382
rect 2150 376 2156 377
rect 2166 354 2172 355
rect 2166 350 2167 354
rect 2171 350 2172 354
rect 2166 349 2172 350
rect 2142 347 2148 348
rect 2142 343 2143 347
rect 2147 343 2148 347
rect 2142 342 2148 343
rect 2168 335 2170 349
rect 2272 348 2274 378
rect 2278 377 2279 381
rect 2283 377 2284 381
rect 2406 379 2407 383
rect 2411 379 2412 383
rect 2416 382 2418 393
rect 2438 383 2444 384
rect 2406 378 2412 379
rect 2414 381 2420 382
rect 2278 376 2284 377
rect 2294 354 2300 355
rect 2294 350 2295 354
rect 2299 350 2300 354
rect 2294 349 2300 350
rect 2270 347 2276 348
rect 2270 343 2271 347
rect 2275 343 2276 347
rect 2270 342 2276 343
rect 2296 335 2298 349
rect 2408 348 2410 378
rect 2414 377 2415 381
rect 2419 377 2420 381
rect 2438 379 2439 383
rect 2443 379 2444 383
rect 2528 382 2530 393
rect 2536 388 2538 442
rect 2542 438 2543 442
rect 2547 438 2548 442
rect 2542 437 2548 438
rect 2560 412 2562 462
rect 2584 455 2586 478
rect 2583 454 2587 455
rect 2583 449 2587 450
rect 2584 434 2586 449
rect 2582 433 2588 434
rect 2582 429 2583 433
rect 2587 429 2588 433
rect 2582 428 2588 429
rect 2582 416 2588 417
rect 2582 412 2583 416
rect 2587 412 2588 416
rect 2558 411 2564 412
rect 2582 411 2588 412
rect 2558 407 2559 411
rect 2563 407 2564 411
rect 2558 406 2564 407
rect 2584 399 2586 411
rect 2583 398 2587 399
rect 2583 393 2587 394
rect 2534 387 2540 388
rect 2534 383 2535 387
rect 2539 383 2540 387
rect 2534 382 2540 383
rect 2438 378 2444 379
rect 2526 381 2532 382
rect 2584 381 2586 393
rect 2414 376 2420 377
rect 2440 357 2442 378
rect 2526 377 2527 381
rect 2531 377 2532 381
rect 2526 376 2532 377
rect 2582 380 2588 381
rect 2582 376 2583 380
rect 2587 376 2588 380
rect 2582 375 2588 376
rect 2582 363 2588 364
rect 2582 359 2583 363
rect 2587 359 2588 363
rect 2582 358 2588 359
rect 2439 356 2443 357
rect 2430 354 2436 355
rect 2430 350 2431 354
rect 2435 350 2436 354
rect 2439 351 2443 352
rect 2542 354 2548 355
rect 2430 349 2436 350
rect 2542 350 2543 354
rect 2547 350 2548 354
rect 2542 349 2548 350
rect 2406 347 2412 348
rect 2406 343 2407 347
rect 2411 343 2412 347
rect 2406 342 2412 343
rect 2432 335 2434 349
rect 2544 335 2546 349
rect 2558 347 2564 348
rect 2558 343 2559 347
rect 2563 343 2564 347
rect 2558 342 2564 343
rect 2143 334 2147 335
rect 2143 329 2147 330
rect 2167 334 2171 335
rect 2167 329 2171 330
rect 2231 334 2235 335
rect 2231 329 2235 330
rect 2295 334 2299 335
rect 2295 329 2299 330
rect 2311 334 2315 335
rect 2311 329 2315 330
rect 2391 334 2395 335
rect 2391 329 2395 330
rect 2431 334 2435 335
rect 2431 329 2435 330
rect 2479 334 2483 335
rect 2479 329 2483 330
rect 2543 334 2547 335
rect 2543 329 2547 330
rect 2122 327 2128 328
rect 2122 323 2123 327
rect 2127 323 2128 327
rect 2144 323 2146 329
rect 2222 327 2228 328
rect 2222 323 2223 327
rect 2227 323 2228 327
rect 2232 323 2234 329
rect 2250 327 2256 328
rect 2250 323 2251 327
rect 2255 323 2256 327
rect 2312 323 2314 329
rect 2330 327 2336 328
rect 2330 323 2331 327
rect 2335 323 2336 327
rect 2392 323 2394 329
rect 2454 327 2460 328
rect 2454 323 2455 327
rect 2459 323 2460 327
rect 2480 323 2482 329
rect 2498 327 2504 328
rect 2498 323 2499 327
rect 2503 323 2504 327
rect 2544 323 2546 329
rect 2030 322 2036 323
rect 2054 322 2060 323
rect 2122 322 2128 323
rect 2142 322 2148 323
rect 2222 322 2228 323
rect 2230 322 2236 323
rect 2250 322 2256 323
rect 2310 322 2316 323
rect 2330 322 2336 323
rect 2390 322 2396 323
rect 2454 322 2460 323
rect 2478 322 2484 323
rect 2498 322 2504 323
rect 2542 322 2548 323
rect 2032 304 2034 322
rect 2054 318 2055 322
rect 2059 318 2060 322
rect 2054 317 2060 318
rect 2142 318 2143 322
rect 2147 318 2148 322
rect 2142 317 2148 318
rect 2030 303 2036 304
rect 2030 299 2031 303
rect 2035 299 2036 303
rect 2030 298 2036 299
rect 2038 295 2044 296
rect 1950 290 1956 291
rect 1982 291 1988 292
rect 1906 286 1912 287
rect 1952 279 1954 290
rect 1982 287 1983 291
rect 1987 287 1988 291
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2126 295 2132 296
rect 2126 291 2127 295
rect 2131 291 2132 295
rect 2126 290 2132 291
rect 2214 295 2220 296
rect 2214 291 2215 295
rect 2219 291 2220 295
rect 2214 290 2220 291
rect 1982 286 1988 287
rect 2040 279 2042 290
rect 2128 279 2130 290
rect 2216 279 2218 290
rect 1671 278 1675 279
rect 1671 273 1675 274
rect 1687 278 1691 279
rect 1687 273 1691 274
rect 1727 278 1731 279
rect 1727 273 1731 274
rect 1775 278 1779 279
rect 1775 273 1779 274
rect 1791 278 1795 279
rect 1791 273 1795 274
rect 1863 278 1867 279
rect 1863 273 1867 274
rect 1871 278 1875 279
rect 1871 273 1875 274
rect 1951 278 1955 279
rect 1951 273 1955 274
rect 2039 278 2043 279
rect 2039 273 2043 274
rect 2119 278 2123 279
rect 2119 273 2123 274
rect 2127 278 2131 279
rect 2127 273 2131 274
rect 2199 278 2203 279
rect 2199 273 2203 274
rect 2215 278 2219 279
rect 2215 273 2219 274
rect 1622 271 1628 272
rect 1622 267 1623 271
rect 1627 267 1628 271
rect 1622 266 1628 267
rect 1678 263 1684 264
rect 1598 258 1604 259
rect 1606 261 1612 262
rect 1534 256 1540 257
rect 1366 255 1372 256
rect 1326 251 1332 252
rect 1366 243 1372 244
rect 1326 239 1332 240
rect 1326 235 1327 239
rect 1331 235 1332 239
rect 1366 239 1367 243
rect 1371 239 1372 243
rect 1366 238 1372 239
rect 1326 234 1332 235
rect 1328 219 1330 234
rect 1368 223 1370 238
rect 1550 234 1556 235
rect 1550 230 1551 234
rect 1555 230 1556 234
rect 1550 229 1556 230
rect 1552 223 1554 229
rect 1600 228 1602 258
rect 1606 257 1607 261
rect 1611 257 1612 261
rect 1678 259 1679 263
rect 1683 259 1684 263
rect 1688 262 1690 273
rect 1766 263 1772 264
rect 1678 258 1684 259
rect 1686 261 1692 262
rect 1606 256 1612 257
rect 1622 234 1628 235
rect 1622 230 1623 234
rect 1627 230 1628 234
rect 1622 229 1628 230
rect 1590 227 1596 228
rect 1590 223 1591 227
rect 1595 223 1596 227
rect 1367 222 1371 223
rect 1327 218 1331 219
rect 1271 213 1275 214
rect 1278 215 1284 216
rect 1114 211 1120 212
rect 1114 207 1115 211
rect 1119 207 1120 211
rect 1152 207 1154 213
rect 1272 207 1274 213
rect 1278 211 1279 215
rect 1283 211 1284 215
rect 1367 217 1371 218
rect 1415 222 1419 223
rect 1415 217 1419 218
rect 1479 222 1483 223
rect 1479 217 1483 218
rect 1551 222 1555 223
rect 1551 217 1555 218
rect 1559 222 1563 223
rect 1590 222 1596 223
rect 1598 227 1604 228
rect 1598 223 1599 227
rect 1603 223 1604 227
rect 1624 223 1626 229
rect 1680 228 1682 258
rect 1686 257 1687 261
rect 1691 257 1692 261
rect 1766 259 1767 263
rect 1771 259 1772 263
rect 1776 262 1778 273
rect 1846 263 1852 264
rect 1766 258 1772 259
rect 1774 261 1780 262
rect 1686 256 1692 257
rect 1702 234 1708 235
rect 1702 230 1703 234
rect 1707 230 1708 234
rect 1702 229 1708 230
rect 1678 227 1684 228
rect 1678 223 1679 227
rect 1683 223 1684 227
rect 1704 223 1706 229
rect 1768 228 1770 258
rect 1774 257 1775 261
rect 1779 257 1780 261
rect 1846 259 1847 263
rect 1851 259 1852 263
rect 1864 262 1866 273
rect 1952 262 1954 273
rect 2030 263 2036 264
rect 1846 258 1852 259
rect 1862 261 1868 262
rect 1774 256 1780 257
rect 1790 234 1796 235
rect 1790 230 1791 234
rect 1795 230 1796 234
rect 1790 229 1796 230
rect 1766 227 1772 228
rect 1766 223 1767 227
rect 1771 223 1772 227
rect 1792 223 1794 229
rect 1848 228 1850 258
rect 1862 257 1863 261
rect 1867 257 1868 261
rect 1862 256 1868 257
rect 1950 261 1956 262
rect 1950 257 1951 261
rect 1955 257 1956 261
rect 2030 259 2031 263
rect 2035 259 2036 263
rect 2040 262 2042 273
rect 2070 263 2076 264
rect 2030 258 2036 259
rect 2038 261 2044 262
rect 1950 256 1956 257
rect 1878 234 1884 235
rect 1878 230 1879 234
rect 1883 230 1884 234
rect 1878 229 1884 230
rect 1966 234 1972 235
rect 1966 230 1967 234
rect 1971 230 1972 234
rect 1966 229 1972 230
rect 1846 227 1852 228
rect 1846 223 1847 227
rect 1851 223 1852 227
rect 1880 223 1882 229
rect 1968 223 1970 229
rect 2032 228 2034 258
rect 2038 257 2039 261
rect 2043 257 2044 261
rect 2070 259 2071 263
rect 2075 259 2076 263
rect 2120 262 2122 273
rect 2190 263 2196 264
rect 2070 258 2076 259
rect 2118 261 2124 262
rect 2038 256 2044 257
rect 2054 234 2060 235
rect 2054 230 2055 234
rect 2059 230 2060 234
rect 2054 229 2060 230
rect 2030 227 2036 228
rect 2030 223 2031 227
rect 2035 223 2036 227
rect 2056 223 2058 229
rect 1598 222 1604 223
rect 1623 222 1627 223
rect 1559 217 1563 218
rect 1327 213 1331 214
rect 1278 210 1284 211
rect 1114 206 1120 207
rect 1150 206 1156 207
rect 1014 174 1020 175
rect 1038 175 1044 176
rect 930 170 936 171
rect 1016 139 1018 174
rect 1038 171 1039 175
rect 1043 171 1044 175
rect 1038 170 1044 171
rect 703 138 707 139
rect 703 133 707 134
rect 759 138 763 139
rect 759 133 763 134
rect 775 138 779 139
rect 775 133 779 134
rect 823 138 827 139
rect 823 133 827 134
rect 887 138 891 139
rect 887 133 891 134
rect 895 138 899 139
rect 895 133 899 134
rect 951 138 955 139
rect 951 133 955 134
rect 1015 138 1019 139
rect 1015 133 1019 134
rect 1079 138 1083 139
rect 1079 133 1083 134
rect 694 123 700 124
rect 694 119 695 123
rect 699 119 700 123
rect 704 122 706 133
rect 750 123 756 124
rect 694 118 700 119
rect 702 121 708 122
rect 696 88 698 118
rect 702 117 703 121
rect 707 117 708 121
rect 750 119 751 123
rect 755 119 756 123
rect 760 122 762 133
rect 814 123 820 124
rect 750 118 756 119
rect 758 121 764 122
rect 702 116 708 117
rect 718 94 724 95
rect 718 90 719 94
rect 723 90 724 94
rect 718 89 724 90
rect 686 87 692 88
rect 686 83 687 87
rect 691 83 692 87
rect 111 82 115 83
rect 111 77 115 78
rect 159 82 163 83
rect 190 82 196 83
rect 215 82 219 83
rect 246 82 252 83
rect 271 82 275 83
rect 302 82 308 83
rect 327 82 331 83
rect 358 82 364 83
rect 383 82 387 83
rect 414 82 420 83
rect 439 82 443 83
rect 470 82 476 83
rect 495 82 499 83
rect 526 82 532 83
rect 551 82 555 83
rect 582 82 588 83
rect 607 82 611 83
rect 159 77 163 78
rect 215 77 219 78
rect 271 77 275 78
rect 327 77 331 78
rect 383 77 387 78
rect 439 77 443 78
rect 495 77 499 78
rect 551 77 555 78
rect 607 77 611 78
rect 663 82 667 83
rect 686 82 692 83
rect 694 87 700 88
rect 694 83 695 87
rect 699 83 700 87
rect 720 83 722 89
rect 752 88 754 118
rect 758 117 759 121
rect 763 117 764 121
rect 814 119 815 123
rect 819 119 820 123
rect 824 122 826 133
rect 878 123 884 124
rect 814 118 820 119
rect 822 121 828 122
rect 758 116 764 117
rect 774 94 780 95
rect 774 90 775 94
rect 779 90 780 94
rect 774 89 780 90
rect 750 87 756 88
rect 750 83 751 87
rect 755 83 756 87
rect 776 83 778 89
rect 816 88 818 118
rect 822 117 823 121
rect 827 117 828 121
rect 878 119 879 123
rect 883 119 884 123
rect 888 122 890 133
rect 942 123 948 124
rect 878 118 884 119
rect 886 121 892 122
rect 822 116 828 117
rect 838 94 844 95
rect 838 90 839 94
rect 843 90 844 94
rect 838 89 844 90
rect 814 87 820 88
rect 814 83 815 87
rect 819 83 820 87
rect 840 83 842 89
rect 880 88 882 118
rect 886 117 887 121
rect 891 117 892 121
rect 942 119 943 123
rect 947 119 948 123
rect 952 122 954 133
rect 1006 123 1012 124
rect 942 118 948 119
rect 950 121 956 122
rect 886 116 892 117
rect 902 94 908 95
rect 902 90 903 94
rect 907 90 908 94
rect 902 89 908 90
rect 878 87 884 88
rect 878 83 879 87
rect 883 83 884 87
rect 904 83 906 89
rect 944 88 946 118
rect 950 117 951 121
rect 955 117 956 121
rect 1006 119 1007 123
rect 1011 119 1012 123
rect 1016 122 1018 133
rect 1070 123 1076 124
rect 1006 118 1012 119
rect 1014 121 1020 122
rect 950 116 956 117
rect 966 94 972 95
rect 966 90 967 94
rect 971 90 972 94
rect 966 89 972 90
rect 942 87 948 88
rect 942 83 943 87
rect 947 83 948 87
rect 968 83 970 89
rect 1008 88 1010 118
rect 1014 117 1015 121
rect 1019 117 1020 121
rect 1070 119 1071 123
rect 1075 119 1076 123
rect 1080 122 1082 133
rect 1116 124 1118 206
rect 1150 202 1151 206
rect 1155 202 1156 206
rect 1150 201 1156 202
rect 1270 206 1276 207
rect 1270 202 1271 206
rect 1275 202 1276 206
rect 1270 201 1276 202
rect 1328 198 1330 213
rect 1368 202 1370 217
rect 1406 215 1412 216
rect 1406 211 1407 215
rect 1411 211 1412 215
rect 1416 211 1418 217
rect 1434 215 1440 216
rect 1434 211 1435 215
rect 1439 211 1440 215
rect 1480 211 1482 217
rect 1498 215 1504 216
rect 1498 211 1499 215
rect 1503 211 1504 215
rect 1560 211 1562 217
rect 1578 215 1584 216
rect 1578 211 1579 215
rect 1583 211 1584 215
rect 1406 210 1412 211
rect 1414 210 1420 211
rect 1434 210 1440 211
rect 1478 210 1484 211
rect 1498 210 1504 211
rect 1558 210 1564 211
rect 1578 210 1584 211
rect 1366 201 1372 202
rect 1326 197 1332 198
rect 1326 193 1327 197
rect 1331 193 1332 197
rect 1366 197 1367 201
rect 1371 197 1372 201
rect 1366 196 1372 197
rect 1326 192 1332 193
rect 1366 184 1372 185
rect 1326 180 1332 181
rect 1134 179 1140 180
rect 1134 175 1135 179
rect 1139 175 1140 179
rect 1134 174 1140 175
rect 1254 179 1260 180
rect 1254 175 1255 179
rect 1259 175 1260 179
rect 1326 176 1327 180
rect 1331 176 1332 180
rect 1366 180 1367 184
rect 1371 180 1372 184
rect 1366 179 1372 180
rect 1398 183 1404 184
rect 1398 179 1399 183
rect 1403 179 1404 183
rect 1326 175 1332 176
rect 1254 174 1260 175
rect 1136 139 1138 174
rect 1198 171 1204 172
rect 1198 167 1199 171
rect 1203 167 1204 171
rect 1198 166 1204 167
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1151 138 1155 139
rect 1151 133 1155 134
rect 1114 123 1120 124
rect 1070 118 1076 119
rect 1078 121 1084 122
rect 1014 116 1020 117
rect 1030 94 1036 95
rect 1030 90 1031 94
rect 1035 90 1036 94
rect 1030 89 1036 90
rect 1006 87 1012 88
rect 1006 83 1007 87
rect 1011 83 1012 87
rect 1032 83 1034 89
rect 1072 88 1074 118
rect 1078 117 1079 121
rect 1083 117 1084 121
rect 1114 119 1115 123
rect 1119 119 1120 123
rect 1152 122 1154 133
rect 1114 118 1120 119
rect 1150 121 1156 122
rect 1078 116 1084 117
rect 1150 117 1151 121
rect 1155 117 1156 121
rect 1150 116 1156 117
rect 1094 94 1100 95
rect 1094 90 1095 94
rect 1099 90 1100 94
rect 1094 89 1100 90
rect 1166 94 1172 95
rect 1166 90 1167 94
rect 1171 90 1172 94
rect 1166 89 1172 90
rect 1070 87 1076 88
rect 1070 83 1071 87
rect 1075 83 1076 87
rect 1096 83 1098 89
rect 1168 83 1170 89
rect 1200 88 1202 166
rect 1256 139 1258 174
rect 1328 139 1330 175
rect 1368 151 1370 179
rect 1398 178 1404 179
rect 1400 151 1402 178
rect 1367 150 1371 151
rect 1367 145 1371 146
rect 1399 150 1403 151
rect 1399 145 1403 146
rect 1215 138 1219 139
rect 1215 133 1219 134
rect 1255 138 1259 139
rect 1255 133 1259 134
rect 1271 138 1275 139
rect 1271 133 1275 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1368 133 1370 145
rect 1400 134 1402 145
rect 1408 141 1410 210
rect 1414 206 1415 210
rect 1419 206 1420 210
rect 1414 205 1420 206
rect 1436 180 1438 210
rect 1478 206 1479 210
rect 1483 206 1484 210
rect 1478 205 1484 206
rect 1462 183 1468 184
rect 1434 179 1440 180
rect 1434 175 1435 179
rect 1439 175 1440 179
rect 1462 179 1463 183
rect 1467 179 1468 183
rect 1500 180 1502 210
rect 1558 206 1559 210
rect 1563 206 1564 210
rect 1558 205 1564 206
rect 1542 183 1548 184
rect 1462 178 1468 179
rect 1498 179 1504 180
rect 1434 174 1440 175
rect 1464 151 1466 178
rect 1498 175 1499 179
rect 1503 175 1504 179
rect 1542 179 1543 183
rect 1547 179 1548 183
rect 1580 180 1582 210
rect 1592 189 1594 222
rect 1623 217 1627 218
rect 1655 222 1659 223
rect 1678 222 1684 223
rect 1703 222 1707 223
rect 1655 217 1659 218
rect 1703 217 1707 218
rect 1751 222 1755 223
rect 1766 222 1772 223
rect 1791 222 1795 223
rect 1846 222 1852 223
rect 1855 222 1859 223
rect 1751 217 1755 218
rect 1791 217 1795 218
rect 1855 217 1859 218
rect 1879 222 1883 223
rect 1879 217 1883 218
rect 1959 222 1963 223
rect 1959 217 1963 218
rect 1967 222 1971 223
rect 2030 222 2036 223
rect 2055 222 2059 223
rect 1967 217 1971 218
rect 2055 217 2059 218
rect 2063 222 2067 223
rect 2072 220 2074 258
rect 2118 257 2119 261
rect 2123 257 2124 261
rect 2190 259 2191 263
rect 2195 259 2196 263
rect 2200 262 2202 273
rect 2224 272 2226 322
rect 2230 318 2231 322
rect 2235 318 2236 322
rect 2230 317 2236 318
rect 2252 292 2254 322
rect 2310 318 2311 322
rect 2315 318 2316 322
rect 2310 317 2316 318
rect 2294 295 2300 296
rect 2250 291 2256 292
rect 2250 287 2251 291
rect 2255 287 2256 291
rect 2294 291 2295 295
rect 2299 291 2300 295
rect 2332 292 2334 322
rect 2390 318 2391 322
rect 2395 318 2396 322
rect 2390 317 2396 318
rect 2374 295 2380 296
rect 2294 290 2300 291
rect 2330 291 2336 292
rect 2250 286 2256 287
rect 2296 279 2298 290
rect 2330 287 2331 291
rect 2335 287 2336 291
rect 2374 291 2375 295
rect 2379 291 2380 295
rect 2374 290 2380 291
rect 2398 291 2404 292
rect 2330 286 2336 287
rect 2376 279 2378 290
rect 2398 287 2399 291
rect 2403 287 2404 291
rect 2398 286 2404 287
rect 2271 278 2275 279
rect 2271 273 2275 274
rect 2295 278 2299 279
rect 2295 273 2299 274
rect 2335 278 2339 279
rect 2335 273 2339 274
rect 2375 278 2379 279
rect 2375 273 2379 274
rect 2222 271 2228 272
rect 2222 267 2223 271
rect 2227 267 2228 271
rect 2222 266 2228 267
rect 2254 263 2260 264
rect 2190 258 2196 259
rect 2198 261 2204 262
rect 2118 256 2124 257
rect 2134 234 2140 235
rect 2134 230 2135 234
rect 2139 230 2140 234
rect 2134 229 2140 230
rect 2136 223 2138 229
rect 2192 228 2194 258
rect 2198 257 2199 261
rect 2203 257 2204 261
rect 2254 259 2255 263
rect 2259 259 2260 263
rect 2272 262 2274 273
rect 2326 263 2332 264
rect 2254 258 2260 259
rect 2270 261 2276 262
rect 2198 256 2204 257
rect 2214 234 2220 235
rect 2214 230 2215 234
rect 2219 230 2220 234
rect 2214 229 2220 230
rect 2182 227 2188 228
rect 2182 223 2183 227
rect 2187 223 2188 227
rect 2135 222 2139 223
rect 2063 217 2067 218
rect 2070 219 2076 220
rect 1656 211 1658 217
rect 1674 215 1680 216
rect 1674 211 1675 215
rect 1679 211 1680 215
rect 1752 211 1754 217
rect 1770 215 1776 216
rect 1770 211 1771 215
rect 1775 211 1776 215
rect 1856 211 1858 217
rect 1934 215 1940 216
rect 1934 211 1935 215
rect 1939 211 1940 215
rect 1960 211 1962 217
rect 2064 211 2066 217
rect 2070 215 2071 219
rect 2075 215 2076 219
rect 2135 217 2139 218
rect 2167 222 2171 223
rect 2182 222 2188 223
rect 2190 227 2196 228
rect 2190 223 2191 227
rect 2195 223 2196 227
rect 2216 223 2218 229
rect 2256 228 2258 258
rect 2270 257 2271 261
rect 2275 257 2276 261
rect 2326 259 2327 263
rect 2331 259 2332 263
rect 2336 262 2338 273
rect 2326 258 2332 259
rect 2334 261 2340 262
rect 2270 256 2276 257
rect 2286 234 2292 235
rect 2286 230 2287 234
rect 2291 230 2292 234
rect 2286 229 2292 230
rect 2254 227 2260 228
rect 2254 223 2255 227
rect 2259 223 2260 227
rect 2288 223 2290 229
rect 2328 228 2330 258
rect 2334 257 2335 261
rect 2339 257 2340 261
rect 2334 256 2340 257
rect 2350 234 2356 235
rect 2350 230 2351 234
rect 2355 230 2356 234
rect 2350 229 2356 230
rect 2326 227 2332 228
rect 2326 223 2327 227
rect 2331 223 2332 227
rect 2352 223 2354 229
rect 2400 228 2402 286
rect 2407 278 2411 279
rect 2407 273 2411 274
rect 2408 262 2410 273
rect 2456 272 2458 322
rect 2478 318 2479 322
rect 2483 318 2484 322
rect 2478 317 2484 318
rect 2462 295 2468 296
rect 2462 291 2463 295
rect 2467 291 2468 295
rect 2500 292 2502 322
rect 2542 318 2543 322
rect 2547 318 2548 322
rect 2542 317 2548 318
rect 2526 295 2532 296
rect 2462 290 2468 291
rect 2498 291 2504 292
rect 2464 279 2466 290
rect 2498 287 2499 291
rect 2503 287 2504 291
rect 2526 291 2527 295
rect 2531 291 2532 295
rect 2560 292 2562 342
rect 2584 335 2586 358
rect 2583 334 2587 335
rect 2583 329 2587 330
rect 2584 314 2586 329
rect 2582 313 2588 314
rect 2582 309 2583 313
rect 2587 309 2588 313
rect 2582 308 2588 309
rect 2582 296 2588 297
rect 2582 292 2583 296
rect 2587 292 2588 296
rect 2526 290 2532 291
rect 2558 291 2564 292
rect 2582 291 2588 292
rect 2498 286 2504 287
rect 2528 279 2530 290
rect 2558 287 2559 291
rect 2563 287 2564 291
rect 2558 286 2564 287
rect 2584 279 2586 291
rect 2463 278 2467 279
rect 2463 273 2467 274
rect 2471 278 2475 279
rect 2471 273 2475 274
rect 2527 278 2531 279
rect 2527 273 2531 274
rect 2583 278 2587 279
rect 2583 273 2587 274
rect 2454 271 2460 272
rect 2454 267 2455 271
rect 2459 267 2460 271
rect 2454 266 2460 267
rect 2472 262 2474 273
rect 2494 263 2500 264
rect 2406 261 2412 262
rect 2406 257 2407 261
rect 2411 257 2412 261
rect 2406 256 2412 257
rect 2470 261 2476 262
rect 2470 257 2471 261
rect 2475 257 2476 261
rect 2494 259 2495 263
rect 2499 259 2500 263
rect 2528 262 2530 273
rect 2494 258 2500 259
rect 2526 261 2532 262
rect 2584 261 2586 273
rect 2470 256 2476 257
rect 2422 234 2428 235
rect 2422 230 2423 234
rect 2427 230 2428 234
rect 2422 229 2428 230
rect 2486 234 2492 235
rect 2486 230 2487 234
rect 2491 230 2492 234
rect 2486 229 2492 230
rect 2398 227 2404 228
rect 2398 223 2399 227
rect 2403 223 2404 227
rect 2424 223 2426 229
rect 2488 223 2490 229
rect 2496 224 2498 258
rect 2526 257 2527 261
rect 2531 257 2532 261
rect 2526 256 2532 257
rect 2582 260 2588 261
rect 2582 256 2583 260
rect 2587 256 2588 260
rect 2582 255 2588 256
rect 2582 243 2588 244
rect 2582 239 2583 243
rect 2587 239 2588 243
rect 2582 238 2588 239
rect 2542 234 2548 235
rect 2542 230 2543 234
rect 2547 230 2548 234
rect 2542 229 2548 230
rect 2494 223 2500 224
rect 2544 223 2546 229
rect 2558 227 2564 228
rect 2558 223 2559 227
rect 2563 223 2564 227
rect 2584 223 2586 238
rect 2190 222 2196 223
rect 2215 222 2219 223
rect 2254 222 2260 223
rect 2263 222 2267 223
rect 2167 217 2171 218
rect 2070 214 2076 215
rect 2158 215 2164 216
rect 2158 211 2159 215
rect 2163 211 2164 215
rect 2168 211 2170 217
rect 1654 210 1660 211
rect 1674 210 1680 211
rect 1750 210 1756 211
rect 1770 210 1776 211
rect 1854 210 1860 211
rect 1934 210 1940 211
rect 1958 210 1964 211
rect 1654 206 1655 210
rect 1659 206 1660 210
rect 1654 205 1660 206
rect 1591 188 1595 189
rect 1591 183 1595 184
rect 1638 183 1644 184
rect 1542 178 1548 179
rect 1578 179 1584 180
rect 1498 174 1504 175
rect 1544 151 1546 178
rect 1578 175 1579 179
rect 1583 175 1584 179
rect 1638 179 1639 183
rect 1643 179 1644 183
rect 1676 180 1678 210
rect 1750 206 1751 210
rect 1755 206 1756 210
rect 1750 205 1756 206
rect 1734 183 1740 184
rect 1638 178 1644 179
rect 1674 179 1680 180
rect 1578 174 1584 175
rect 1640 151 1642 178
rect 1674 175 1675 179
rect 1679 175 1680 179
rect 1734 179 1735 183
rect 1739 179 1740 183
rect 1772 180 1774 210
rect 1854 206 1855 210
rect 1859 206 1860 210
rect 1854 205 1860 206
rect 1936 192 1938 210
rect 1958 206 1959 210
rect 1963 206 1964 210
rect 1958 205 1964 206
rect 2062 210 2068 211
rect 2158 210 2164 211
rect 2166 210 2172 211
rect 2062 206 2063 210
rect 2067 206 2068 210
rect 2062 205 2068 206
rect 1934 191 1940 192
rect 1871 188 1875 189
rect 1934 187 1935 191
rect 1939 187 1940 191
rect 1934 186 1940 187
rect 1838 183 1844 184
rect 1871 183 1875 184
rect 1942 183 1948 184
rect 1734 178 1740 179
rect 1770 179 1776 180
rect 1674 174 1680 175
rect 1736 151 1738 178
rect 1770 175 1771 179
rect 1775 175 1776 179
rect 1838 179 1839 183
rect 1843 179 1844 183
rect 1872 180 1874 183
rect 1838 178 1844 179
rect 1870 179 1876 180
rect 1770 174 1776 175
rect 1840 151 1842 178
rect 1870 175 1871 179
rect 1875 175 1876 179
rect 1942 179 1943 183
rect 1947 179 1948 183
rect 1942 178 1948 179
rect 2046 183 2052 184
rect 2046 179 2047 183
rect 2051 179 2052 183
rect 2046 178 2052 179
rect 2150 183 2156 184
rect 2150 179 2151 183
rect 2155 179 2156 183
rect 2150 178 2156 179
rect 1870 174 1876 175
rect 1894 175 1900 176
rect 1894 171 1895 175
rect 1899 171 1900 175
rect 1894 170 1900 171
rect 1455 150 1459 151
rect 1455 145 1459 146
rect 1463 150 1467 151
rect 1463 145 1467 146
rect 1511 150 1515 151
rect 1511 145 1515 146
rect 1543 150 1547 151
rect 1543 145 1547 146
rect 1567 150 1571 151
rect 1567 145 1571 146
rect 1631 150 1635 151
rect 1631 145 1635 146
rect 1639 150 1643 151
rect 1639 145 1643 146
rect 1711 150 1715 151
rect 1711 145 1715 146
rect 1735 150 1739 151
rect 1735 145 1739 146
rect 1791 150 1795 151
rect 1791 145 1795 146
rect 1839 150 1843 151
rect 1839 145 1843 146
rect 1871 150 1875 151
rect 1871 145 1875 146
rect 1407 140 1411 141
rect 1407 135 1411 136
rect 1446 135 1452 136
rect 1398 133 1404 134
rect 1206 123 1212 124
rect 1206 119 1207 123
rect 1211 119 1212 123
rect 1216 122 1218 133
rect 1262 123 1268 124
rect 1206 118 1212 119
rect 1214 121 1220 122
rect 1208 88 1210 118
rect 1214 117 1215 121
rect 1219 117 1220 121
rect 1262 119 1263 123
rect 1267 119 1268 123
rect 1272 122 1274 133
rect 1262 118 1268 119
rect 1270 121 1276 122
rect 1328 121 1330 133
rect 1366 132 1372 133
rect 1366 128 1367 132
rect 1371 128 1372 132
rect 1398 129 1399 133
rect 1403 129 1404 133
rect 1446 131 1447 135
rect 1451 131 1452 135
rect 1456 134 1458 145
rect 1502 135 1508 136
rect 1446 130 1452 131
rect 1454 133 1460 134
rect 1398 128 1404 129
rect 1366 127 1372 128
rect 1214 116 1220 117
rect 1230 94 1236 95
rect 1230 90 1231 94
rect 1235 90 1236 94
rect 1230 89 1236 90
rect 1198 87 1204 88
rect 1198 83 1199 87
rect 1203 83 1204 87
rect 694 82 700 83
rect 719 82 723 83
rect 750 82 756 83
rect 775 82 779 83
rect 814 82 820 83
rect 839 82 843 83
rect 878 82 884 83
rect 903 82 907 83
rect 942 82 948 83
rect 967 82 971 83
rect 1006 82 1012 83
rect 1031 82 1035 83
rect 1070 82 1076 83
rect 1095 82 1099 83
rect 663 77 667 78
rect 719 77 723 78
rect 775 77 779 78
rect 839 77 843 78
rect 903 77 907 78
rect 967 77 971 78
rect 1031 77 1035 78
rect 1095 77 1099 78
rect 1167 82 1171 83
rect 1198 82 1204 83
rect 1206 87 1212 88
rect 1206 83 1207 87
rect 1211 83 1212 87
rect 1232 83 1234 89
rect 1264 88 1266 118
rect 1270 117 1271 121
rect 1275 117 1276 121
rect 1270 116 1276 117
rect 1326 120 1332 121
rect 1326 116 1327 120
rect 1331 116 1332 120
rect 1326 115 1332 116
rect 1366 115 1372 116
rect 1366 111 1367 115
rect 1371 111 1372 115
rect 1366 110 1372 111
rect 1326 103 1332 104
rect 1326 99 1327 103
rect 1331 99 1332 103
rect 1326 98 1332 99
rect 1286 94 1292 95
rect 1286 90 1287 94
rect 1291 90 1292 94
rect 1286 89 1292 90
rect 1262 87 1268 88
rect 1262 83 1263 87
rect 1267 83 1268 87
rect 1288 83 1290 89
rect 1328 83 1330 98
rect 1368 95 1370 110
rect 1414 106 1420 107
rect 1414 102 1415 106
rect 1419 102 1420 106
rect 1414 101 1420 102
rect 1416 95 1418 101
rect 1448 100 1450 130
rect 1454 129 1455 133
rect 1459 129 1460 133
rect 1502 131 1503 135
rect 1507 131 1508 135
rect 1512 134 1514 145
rect 1558 135 1564 136
rect 1502 130 1508 131
rect 1510 133 1516 134
rect 1454 128 1460 129
rect 1470 106 1476 107
rect 1470 102 1471 106
rect 1475 102 1476 106
rect 1470 101 1476 102
rect 1446 99 1452 100
rect 1446 95 1447 99
rect 1451 95 1452 99
rect 1472 95 1474 101
rect 1504 100 1506 130
rect 1510 129 1511 133
rect 1515 129 1516 133
rect 1558 131 1559 135
rect 1563 131 1564 135
rect 1568 134 1570 145
rect 1622 135 1628 136
rect 1558 130 1564 131
rect 1566 133 1572 134
rect 1510 128 1516 129
rect 1526 106 1532 107
rect 1526 102 1527 106
rect 1531 102 1532 106
rect 1526 101 1532 102
rect 1502 99 1508 100
rect 1502 95 1503 99
rect 1507 95 1508 99
rect 1528 95 1530 101
rect 1560 100 1562 130
rect 1566 129 1567 133
rect 1571 129 1572 133
rect 1622 131 1623 135
rect 1627 131 1628 135
rect 1632 134 1634 145
rect 1702 135 1708 136
rect 1622 130 1628 131
rect 1630 133 1636 134
rect 1566 128 1572 129
rect 1582 106 1588 107
rect 1582 102 1583 106
rect 1587 102 1588 106
rect 1582 101 1588 102
rect 1558 99 1564 100
rect 1558 95 1559 99
rect 1563 95 1564 99
rect 1584 95 1586 101
rect 1624 100 1626 130
rect 1630 129 1631 133
rect 1635 129 1636 133
rect 1702 131 1703 135
rect 1707 131 1708 135
rect 1712 134 1714 145
rect 1782 135 1788 136
rect 1702 130 1708 131
rect 1710 133 1716 134
rect 1630 128 1636 129
rect 1646 106 1652 107
rect 1646 102 1647 106
rect 1651 102 1652 106
rect 1646 101 1652 102
rect 1622 99 1628 100
rect 1622 95 1623 99
rect 1627 95 1628 99
rect 1648 95 1650 101
rect 1704 100 1706 130
rect 1710 129 1711 133
rect 1715 129 1716 133
rect 1782 131 1783 135
rect 1787 131 1788 135
rect 1792 134 1794 145
rect 1823 140 1827 141
rect 1822 135 1828 136
rect 1782 130 1788 131
rect 1790 133 1796 134
rect 1710 128 1716 129
rect 1726 106 1732 107
rect 1726 102 1727 106
rect 1731 102 1732 106
rect 1726 101 1732 102
rect 1702 99 1708 100
rect 1702 95 1703 99
rect 1707 95 1708 99
rect 1728 95 1730 101
rect 1784 100 1786 130
rect 1790 129 1791 133
rect 1795 129 1796 133
rect 1822 131 1823 135
rect 1827 131 1828 135
rect 1872 134 1874 145
rect 1822 130 1828 131
rect 1870 133 1876 134
rect 1790 128 1796 129
rect 1870 129 1871 133
rect 1875 129 1876 133
rect 1870 128 1876 129
rect 1806 106 1812 107
rect 1806 102 1807 106
rect 1811 102 1812 106
rect 1806 101 1812 102
rect 1886 106 1892 107
rect 1886 102 1887 106
rect 1891 102 1892 106
rect 1886 101 1892 102
rect 1782 99 1788 100
rect 1782 95 1783 99
rect 1787 95 1788 99
rect 1808 95 1810 101
rect 1888 95 1890 101
rect 1896 100 1898 170
rect 1944 151 1946 178
rect 2048 151 2050 178
rect 2152 151 2154 178
rect 2160 172 2162 210
rect 2166 206 2167 210
rect 2171 206 2172 210
rect 2166 205 2172 206
rect 2184 180 2186 222
rect 2215 217 2219 218
rect 2263 217 2267 218
rect 2287 222 2291 223
rect 2326 222 2332 223
rect 2351 222 2355 223
rect 2287 217 2291 218
rect 2351 217 2355 218
rect 2359 222 2363 223
rect 2398 222 2404 223
rect 2423 222 2427 223
rect 2359 217 2363 218
rect 2423 217 2427 218
rect 2463 222 2467 223
rect 2463 217 2467 218
rect 2487 222 2491 223
rect 2494 219 2495 223
rect 2499 219 2500 223
rect 2494 218 2500 219
rect 2543 222 2547 223
rect 2558 222 2564 223
rect 2583 222 2587 223
rect 2487 217 2491 218
rect 2543 217 2547 218
rect 2238 215 2244 216
rect 2238 211 2239 215
rect 2243 211 2244 215
rect 2264 211 2266 217
rect 2334 215 2340 216
rect 2334 211 2335 215
rect 2339 211 2340 215
rect 2360 211 2362 217
rect 2464 211 2466 217
rect 2544 211 2546 217
rect 2238 210 2244 211
rect 2262 210 2268 211
rect 2334 210 2340 211
rect 2358 210 2364 211
rect 2240 192 2242 210
rect 2262 206 2263 210
rect 2267 206 2268 210
rect 2262 205 2268 206
rect 2238 191 2244 192
rect 2238 187 2239 191
rect 2243 187 2244 191
rect 2238 186 2244 187
rect 2246 183 2252 184
rect 2182 179 2188 180
rect 2182 175 2183 179
rect 2187 175 2188 179
rect 2246 179 2247 183
rect 2251 179 2252 183
rect 2246 178 2252 179
rect 2182 174 2188 175
rect 2158 171 2164 172
rect 2158 167 2159 171
rect 2163 167 2164 171
rect 2158 166 2164 167
rect 2248 151 2250 178
rect 1943 150 1947 151
rect 1943 145 1947 146
rect 2015 150 2019 151
rect 2015 145 2019 146
rect 2047 150 2051 151
rect 2047 145 2051 146
rect 2079 150 2083 151
rect 2079 145 2083 146
rect 2143 150 2147 151
rect 2143 145 2147 146
rect 2151 150 2155 151
rect 2151 145 2155 146
rect 2207 150 2211 151
rect 2207 145 2211 146
rect 2247 150 2251 151
rect 2247 145 2251 146
rect 2271 150 2275 151
rect 2271 145 2275 146
rect 1934 135 1940 136
rect 1934 131 1935 135
rect 1939 131 1940 135
rect 1944 134 1946 145
rect 2006 135 2012 136
rect 1934 130 1940 131
rect 1942 133 1948 134
rect 1936 100 1938 130
rect 1942 129 1943 133
rect 1947 129 1948 133
rect 2006 131 2007 135
rect 2011 131 2012 135
rect 2016 134 2018 145
rect 2070 135 2076 136
rect 2006 130 2012 131
rect 2014 133 2020 134
rect 1942 128 1948 129
rect 1958 106 1964 107
rect 1958 102 1959 106
rect 1963 102 1964 106
rect 1958 101 1964 102
rect 1894 99 1900 100
rect 1894 95 1895 99
rect 1899 95 1900 99
rect 1367 94 1371 95
rect 1367 89 1371 90
rect 1415 94 1419 95
rect 1446 94 1452 95
rect 1471 94 1475 95
rect 1502 94 1508 95
rect 1527 94 1531 95
rect 1558 94 1564 95
rect 1583 94 1587 95
rect 1622 94 1628 95
rect 1647 94 1651 95
rect 1702 94 1708 95
rect 1727 94 1731 95
rect 1782 94 1788 95
rect 1807 94 1811 95
rect 1415 89 1419 90
rect 1471 89 1475 90
rect 1527 89 1531 90
rect 1583 89 1587 90
rect 1647 89 1651 90
rect 1727 89 1731 90
rect 1807 89 1811 90
rect 1887 94 1891 95
rect 1894 94 1900 95
rect 1934 99 1940 100
rect 1934 95 1935 99
rect 1939 95 1940 99
rect 1960 95 1962 101
rect 2008 100 2010 130
rect 2014 129 2015 133
rect 2019 129 2020 133
rect 2070 131 2071 135
rect 2075 131 2076 135
rect 2080 134 2082 145
rect 2134 135 2140 136
rect 2070 130 2076 131
rect 2078 133 2084 134
rect 2014 128 2020 129
rect 2030 106 2036 107
rect 2030 102 2031 106
rect 2035 102 2036 106
rect 2030 101 2036 102
rect 2006 99 2012 100
rect 2006 95 2007 99
rect 2011 95 2012 99
rect 2032 95 2034 101
rect 2072 100 2074 130
rect 2078 129 2079 133
rect 2083 129 2084 133
rect 2134 131 2135 135
rect 2139 131 2140 135
rect 2144 134 2146 145
rect 2198 135 2204 136
rect 2134 130 2140 131
rect 2142 133 2148 134
rect 2078 128 2084 129
rect 2094 106 2100 107
rect 2094 102 2095 106
rect 2099 102 2100 106
rect 2094 101 2100 102
rect 2070 99 2076 100
rect 2070 95 2071 99
rect 2075 95 2076 99
rect 2096 95 2098 101
rect 2136 100 2138 130
rect 2142 129 2143 133
rect 2147 129 2148 133
rect 2198 131 2199 135
rect 2203 131 2204 135
rect 2208 134 2210 145
rect 2262 135 2268 136
rect 2198 130 2204 131
rect 2206 133 2212 134
rect 2142 128 2148 129
rect 2158 106 2164 107
rect 2158 102 2159 106
rect 2163 102 2164 106
rect 2158 101 2164 102
rect 2134 99 2140 100
rect 2134 95 2135 99
rect 2139 95 2140 99
rect 2160 95 2162 101
rect 2200 100 2202 130
rect 2206 129 2207 133
rect 2211 129 2212 133
rect 2262 131 2263 135
rect 2267 131 2268 135
rect 2272 134 2274 145
rect 2336 144 2338 210
rect 2358 206 2359 210
rect 2363 206 2364 210
rect 2358 205 2364 206
rect 2462 210 2468 211
rect 2462 206 2463 210
rect 2467 206 2468 210
rect 2462 205 2468 206
rect 2542 210 2548 211
rect 2542 206 2543 210
rect 2547 206 2548 210
rect 2542 205 2548 206
rect 2342 183 2348 184
rect 2342 179 2343 183
rect 2347 179 2348 183
rect 2342 178 2348 179
rect 2446 183 2452 184
rect 2446 179 2447 183
rect 2451 179 2452 183
rect 2446 178 2452 179
rect 2526 183 2532 184
rect 2526 179 2527 183
rect 2531 179 2532 183
rect 2560 180 2562 222
rect 2583 217 2587 218
rect 2584 202 2586 217
rect 2582 201 2588 202
rect 2582 197 2583 201
rect 2587 197 2588 201
rect 2582 196 2588 197
rect 2582 184 2588 185
rect 2582 180 2583 184
rect 2587 180 2588 184
rect 2526 178 2532 179
rect 2558 179 2564 180
rect 2582 179 2588 180
rect 2344 151 2346 178
rect 2448 151 2450 178
rect 2528 151 2530 178
rect 2558 175 2559 179
rect 2563 175 2564 179
rect 2558 174 2564 175
rect 2584 151 2586 179
rect 2343 150 2347 151
rect 2343 145 2347 146
rect 2415 150 2419 151
rect 2415 145 2419 146
rect 2447 150 2451 151
rect 2447 145 2451 146
rect 2527 150 2531 151
rect 2527 145 2531 146
rect 2583 150 2587 151
rect 2583 145 2587 146
rect 2334 143 2340 144
rect 2334 139 2335 143
rect 2339 139 2340 143
rect 2334 138 2340 139
rect 2334 135 2340 136
rect 2262 130 2268 131
rect 2270 133 2276 134
rect 2206 128 2212 129
rect 2222 106 2228 107
rect 2222 102 2223 106
rect 2227 102 2228 106
rect 2222 101 2228 102
rect 2198 99 2204 100
rect 2198 95 2199 99
rect 2203 95 2204 99
rect 2224 95 2226 101
rect 2264 100 2266 130
rect 2270 129 2271 133
rect 2275 129 2276 133
rect 2334 131 2335 135
rect 2339 131 2340 135
rect 2344 134 2346 145
rect 2406 135 2412 136
rect 2334 130 2340 131
rect 2342 133 2348 134
rect 2270 128 2276 129
rect 2286 106 2292 107
rect 2286 102 2287 106
rect 2291 102 2292 106
rect 2286 101 2292 102
rect 2262 99 2268 100
rect 2262 95 2263 99
rect 2267 95 2268 99
rect 2288 95 2290 101
rect 2336 100 2338 130
rect 2342 129 2343 133
rect 2347 129 2348 133
rect 2406 131 2407 135
rect 2411 131 2412 135
rect 2416 134 2418 145
rect 2406 130 2412 131
rect 2414 133 2420 134
rect 2584 133 2586 145
rect 2342 128 2348 129
rect 2358 106 2364 107
rect 2358 102 2359 106
rect 2363 102 2364 106
rect 2358 101 2364 102
rect 2334 99 2340 100
rect 2334 95 2335 99
rect 2339 95 2340 99
rect 2360 95 2362 101
rect 2408 100 2410 130
rect 2414 129 2415 133
rect 2419 129 2420 133
rect 2414 128 2420 129
rect 2582 132 2588 133
rect 2582 128 2583 132
rect 2587 128 2588 132
rect 2582 127 2588 128
rect 2582 115 2588 116
rect 2582 111 2583 115
rect 2587 111 2588 115
rect 2582 110 2588 111
rect 2430 106 2436 107
rect 2430 102 2431 106
rect 2435 102 2436 106
rect 2430 101 2436 102
rect 2406 99 2412 100
rect 2406 95 2407 99
rect 2411 95 2412 99
rect 2432 95 2434 101
rect 2584 95 2586 110
rect 1934 94 1940 95
rect 1959 94 1963 95
rect 2006 94 2012 95
rect 2031 94 2035 95
rect 2070 94 2076 95
rect 2095 94 2099 95
rect 2134 94 2140 95
rect 2159 94 2163 95
rect 2198 94 2204 95
rect 2223 94 2227 95
rect 2262 94 2268 95
rect 2287 94 2291 95
rect 2334 94 2340 95
rect 2359 94 2363 95
rect 2406 94 2412 95
rect 2431 94 2435 95
rect 1887 89 1891 90
rect 1959 89 1963 90
rect 2031 89 2035 90
rect 2095 89 2099 90
rect 2159 89 2163 90
rect 2223 89 2227 90
rect 2287 89 2291 90
rect 2359 89 2363 90
rect 2431 89 2435 90
rect 2583 94 2587 95
rect 2583 89 2587 90
rect 1206 82 1212 83
rect 1231 82 1235 83
rect 1262 82 1268 83
rect 1287 82 1291 83
rect 1167 77 1171 78
rect 1231 77 1235 78
rect 1287 77 1291 78
rect 1327 82 1331 83
rect 1327 77 1331 78
<< m4c >>
rect 111 2638 115 2642
rect 551 2638 555 2642
rect 607 2638 611 2642
rect 663 2638 667 2642
rect 719 2638 723 2642
rect 775 2638 779 2642
rect 111 2582 115 2586
rect 215 2582 219 2586
rect 271 2582 275 2586
rect 327 2582 331 2586
rect 383 2582 387 2586
rect 439 2582 443 2586
rect 495 2582 499 2586
rect 535 2582 539 2586
rect 551 2582 555 2586
rect 111 2522 115 2526
rect 231 2522 235 2526
rect 287 2522 291 2526
rect 343 2522 347 2526
rect 1327 2638 1331 2642
rect 591 2582 595 2586
rect 607 2582 611 2586
rect 647 2582 651 2586
rect 663 2582 667 2586
rect 703 2582 707 2586
rect 719 2582 723 2586
rect 1367 2634 1371 2638
rect 1551 2634 1555 2638
rect 1607 2634 1611 2638
rect 1663 2634 1667 2638
rect 759 2582 763 2586
rect 775 2582 779 2586
rect 831 2582 835 2586
rect 887 2582 891 2586
rect 943 2582 947 2586
rect 999 2582 1003 2586
rect 1055 2582 1059 2586
rect 1111 2582 1115 2586
rect 1327 2582 1331 2586
rect 1719 2634 1723 2638
rect 1775 2634 1779 2638
rect 1367 2578 1371 2582
rect 1439 2578 1443 2582
rect 367 2522 371 2526
rect 399 2522 403 2526
rect 423 2522 427 2526
rect 455 2522 459 2526
rect 487 2522 491 2526
rect 511 2522 515 2526
rect 551 2522 555 2526
rect 567 2522 571 2526
rect 615 2522 619 2526
rect 623 2522 627 2526
rect 679 2522 683 2526
rect 735 2522 739 2526
rect 743 2522 747 2526
rect 791 2522 795 2526
rect 807 2522 811 2526
rect 847 2522 851 2526
rect 871 2522 875 2526
rect 903 2522 907 2526
rect 943 2522 947 2526
rect 959 2522 963 2526
rect 1015 2522 1019 2526
rect 1071 2522 1075 2526
rect 111 2462 115 2466
rect 271 2462 275 2466
rect 335 2462 339 2466
rect 351 2462 355 2466
rect 399 2462 403 2466
rect 407 2462 411 2466
rect 471 2462 475 2466
rect 535 2462 539 2466
rect 551 2462 555 2466
rect 599 2462 603 2466
rect 111 2402 115 2406
rect 247 2402 251 2406
rect 287 2402 291 2406
rect 335 2402 339 2406
rect 351 2402 355 2406
rect 415 2402 419 2406
rect 1127 2522 1131 2526
rect 1327 2522 1331 2526
rect 1831 2634 1835 2638
rect 1887 2634 1891 2638
rect 1943 2634 1947 2638
rect 1999 2634 2003 2638
rect 2055 2634 2059 2638
rect 2111 2634 2115 2638
rect 2167 2634 2171 2638
rect 2583 2634 2587 2638
rect 1535 2578 1539 2582
rect 1543 2578 1547 2582
rect 1591 2578 1595 2582
rect 1647 2578 1651 2582
rect 1655 2578 1659 2582
rect 1703 2578 1707 2582
rect 1759 2578 1763 2582
rect 1767 2578 1771 2582
rect 1815 2578 1819 2582
rect 1871 2578 1875 2582
rect 1879 2578 1883 2582
rect 1927 2578 1931 2582
rect 1983 2578 1987 2582
rect 1991 2578 1995 2582
rect 1543 2528 1547 2532
rect 1367 2514 1371 2518
rect 1455 2514 1459 2518
rect 2039 2578 2043 2582
rect 2095 2578 2099 2582
rect 2111 2578 2115 2582
rect 2151 2578 2155 2582
rect 2231 2578 2235 2582
rect 2351 2578 2355 2582
rect 2583 2578 2587 2582
rect 1903 2528 1907 2532
rect 1551 2514 1555 2518
rect 1559 2514 1563 2518
rect 1631 2514 1635 2518
rect 1671 2514 1675 2518
rect 1719 2514 1723 2518
rect 1783 2514 1787 2518
rect 1807 2514 1811 2518
rect 1895 2514 1899 2518
rect 1903 2514 1907 2518
rect 1999 2514 2003 2518
rect 2007 2514 2011 2518
rect 2095 2514 2099 2518
rect 2127 2514 2131 2518
rect 2191 2514 2195 2518
rect 2247 2514 2251 2518
rect 2295 2514 2299 2518
rect 631 2462 635 2466
rect 663 2462 667 2466
rect 711 2462 715 2466
rect 727 2462 731 2466
rect 783 2462 787 2466
rect 791 2462 795 2466
rect 855 2462 859 2466
rect 863 2462 867 2466
rect 927 2462 931 2466
rect 943 2462 947 2466
rect 999 2462 1003 2466
rect 1023 2462 1027 2466
rect 1327 2462 1331 2466
rect 1367 2458 1371 2462
rect 1535 2458 1539 2462
rect 1615 2458 1619 2462
rect 1647 2458 1651 2462
rect 431 2402 435 2406
rect 487 2402 491 2406
rect 527 2402 531 2406
rect 567 2402 571 2406
rect 631 2402 635 2406
rect 647 2402 651 2406
rect 727 2402 731 2406
rect 799 2402 803 2406
rect 823 2402 827 2406
rect 879 2402 883 2406
rect 919 2402 923 2406
rect 239 2368 243 2372
rect 111 2346 115 2350
rect 159 2346 163 2350
rect 231 2346 235 2350
rect 263 2346 267 2350
rect 319 2346 323 2350
rect 111 2286 115 2290
rect 159 2286 163 2290
rect 175 2286 179 2290
rect 247 2286 251 2290
rect 279 2286 283 2290
rect 647 2368 651 2372
rect 959 2402 963 2406
rect 1015 2402 1019 2406
rect 1039 2402 1043 2406
rect 1111 2402 1115 2406
rect 1327 2402 1331 2406
rect 1703 2458 1707 2462
rect 1767 2458 1771 2462
rect 1791 2458 1795 2462
rect 1839 2458 1843 2462
rect 1887 2458 1891 2462
rect 1911 2458 1915 2462
rect 2367 2514 2371 2518
rect 2399 2514 2403 2518
rect 2583 2514 2587 2518
rect 1983 2458 1987 2462
rect 1991 2458 1995 2462
rect 2079 2458 2083 2462
rect 2167 2458 2171 2462
rect 2175 2458 2179 2462
rect 1367 2398 1371 2402
rect 1455 2398 1459 2402
rect 1559 2398 1563 2402
rect 1663 2398 1667 2402
rect 1719 2398 1723 2402
rect 1759 2398 1763 2402
rect 1783 2398 1787 2402
rect 1855 2398 1859 2402
rect 1927 2398 1931 2402
rect 1943 2398 1947 2402
rect 375 2346 379 2350
rect 415 2346 419 2350
rect 487 2346 491 2350
rect 511 2346 515 2350
rect 599 2346 603 2350
rect 615 2346 619 2350
rect 711 2346 715 2350
rect 807 2346 811 2350
rect 815 2346 819 2350
rect 903 2346 907 2350
rect 911 2346 915 2350
rect 999 2346 1003 2350
rect 1007 2346 1011 2350
rect 1095 2346 1099 2350
rect 1103 2346 1107 2350
rect 1199 2346 1203 2350
rect 1327 2346 1331 2350
rect 375 2286 379 2290
rect 391 2286 395 2290
rect 503 2286 507 2290
rect 511 2286 515 2290
rect 615 2286 619 2290
rect 639 2286 643 2290
rect 727 2286 731 2290
rect 111 2222 115 2226
rect 143 2222 147 2226
rect 139 2184 143 2188
rect 111 2162 115 2166
rect 767 2286 771 2290
rect 831 2286 835 2290
rect 887 2286 891 2290
rect 927 2286 931 2290
rect 999 2286 1003 2290
rect 1367 2342 1371 2346
rect 1399 2342 1403 2346
rect 1439 2342 1443 2346
rect 1455 2342 1459 2346
rect 1511 2342 1515 2346
rect 1023 2286 1027 2290
rect 1103 2286 1107 2290
rect 1119 2286 1123 2290
rect 1207 2286 1211 2290
rect 1215 2286 1219 2290
rect 1287 2286 1291 2290
rect 231 2222 235 2226
rect 359 2222 363 2226
rect 495 2222 499 2226
rect 623 2222 627 2226
rect 751 2222 755 2226
rect 871 2222 875 2226
rect 983 2222 987 2226
rect 1087 2222 1091 2226
rect 1191 2222 1195 2226
rect 647 2184 651 2188
rect 159 2162 163 2166
rect 215 2162 219 2166
rect 247 2162 251 2166
rect 311 2162 315 2166
rect 375 2162 379 2166
rect 423 2162 427 2166
rect 511 2162 515 2166
rect 543 2162 547 2166
rect 639 2162 643 2166
rect 663 2162 667 2166
rect 767 2162 771 2166
rect 775 2162 779 2166
rect 111 2098 115 2102
rect 143 2098 147 2102
rect 199 2098 203 2102
rect 263 2098 267 2102
rect 295 2098 299 2102
rect 327 2098 331 2102
rect 399 2098 403 2102
rect 407 2098 411 2102
rect 479 2098 483 2102
rect 527 2098 531 2102
rect 567 2098 571 2102
rect 647 2098 651 2102
rect 655 2098 659 2102
rect 259 2072 263 2076
rect 735 2098 739 2102
rect 1327 2286 1331 2290
rect 2007 2398 2011 2402
rect 2039 2398 2043 2402
rect 2095 2398 2099 2402
rect 1543 2342 1547 2346
rect 1567 2342 1571 2346
rect 1639 2342 1643 2346
rect 1647 2342 1651 2346
rect 1727 2342 1731 2346
rect 1743 2342 1747 2346
rect 1823 2342 1827 2346
rect 1839 2342 1843 2346
rect 1367 2278 1371 2282
rect 1415 2278 1419 2282
rect 1471 2278 1475 2282
rect 1495 2278 1499 2282
rect 1527 2278 1531 2282
rect 1583 2278 1587 2282
rect 1615 2278 1619 2282
rect 1655 2278 1659 2282
rect 1735 2278 1739 2282
rect 1743 2278 1747 2282
rect 1271 2222 1275 2226
rect 1327 2222 1331 2226
rect 1367 2210 1371 2214
rect 1399 2210 1403 2214
rect 1455 2210 1459 2214
rect 1479 2210 1483 2214
rect 1535 2210 1539 2214
rect 1599 2210 1603 2214
rect 1631 2210 1635 2214
rect 879 2162 883 2166
rect 887 2162 891 2166
rect 975 2162 979 2166
rect 999 2162 1003 2166
rect 1071 2162 1075 2166
rect 1103 2162 1107 2166
rect 1167 2162 1171 2166
rect 1207 2162 1211 2166
rect 1271 2162 1275 2166
rect 1287 2162 1291 2166
rect 1327 2162 1331 2166
rect 855 2128 859 2132
rect 2135 2398 2139 2402
rect 2183 2398 2187 2402
rect 2263 2458 2267 2462
rect 2279 2458 2283 2462
rect 2359 2458 2363 2462
rect 2383 2458 2387 2462
rect 2455 2458 2459 2462
rect 2527 2458 2531 2462
rect 2583 2458 2587 2462
rect 2231 2398 2235 2402
rect 2279 2398 2283 2402
rect 2335 2398 2339 2402
rect 2375 2398 2379 2402
rect 1927 2342 1931 2346
rect 1943 2342 1947 2346
rect 2023 2342 2027 2346
rect 2079 2342 2083 2346
rect 2119 2342 2123 2346
rect 2215 2342 2219 2346
rect 2223 2342 2227 2346
rect 2319 2342 2323 2346
rect 2383 2342 2387 2346
rect 1839 2278 1843 2282
rect 1855 2278 1859 2282
rect 1959 2278 1963 2282
rect 1967 2278 1971 2282
rect 2071 2278 2075 2282
rect 2095 2278 2099 2282
rect 2167 2278 2171 2282
rect 2239 2278 2243 2282
rect 2255 2278 2259 2282
rect 2335 2278 2339 2282
rect 2399 2278 2403 2282
rect 2407 2278 2411 2282
rect 1719 2210 1723 2214
rect 1743 2210 1747 2214
rect 1839 2210 1843 2214
rect 1863 2210 1867 2214
rect 1951 2210 1955 2214
rect 1983 2210 1987 2214
rect 2055 2210 2059 2214
rect 2095 2210 2099 2214
rect 2151 2210 2155 2214
rect 2207 2210 2211 2214
rect 2239 2210 2243 2214
rect 2311 2210 2315 2214
rect 2319 2210 2323 2214
rect 1367 2154 1371 2158
rect 1471 2154 1475 2158
rect 1535 2154 1539 2158
rect 1551 2154 1555 2158
rect 1631 2154 1635 2158
rect 1647 2154 1651 2158
rect 1735 2154 1739 2158
rect 1759 2154 1763 2158
rect 1839 2154 1843 2158
rect 1879 2154 1883 2158
rect 1951 2154 1955 2158
rect 1999 2154 2003 2158
rect 2447 2398 2451 2402
rect 2471 2398 2475 2402
rect 2543 2398 2547 2402
rect 2431 2342 2435 2346
rect 2527 2342 2531 2346
rect 2583 2398 2587 2402
rect 2583 2342 2587 2346
rect 2487 2278 2491 2282
rect 2543 2278 2547 2282
rect 2583 2278 2587 2282
rect 2391 2210 2395 2214
rect 2423 2210 2427 2214
rect 2471 2210 2475 2214
rect 2527 2210 2531 2214
rect 2583 2210 2587 2214
rect 1287 2128 1291 2132
rect 2055 2154 2059 2158
rect 759 2098 763 2102
rect 815 2098 819 2102
rect 863 2098 867 2102
rect 887 2098 891 2102
rect 959 2098 963 2102
rect 967 2098 971 2102
rect 1047 2098 1051 2102
rect 1055 2098 1059 2102
rect 1127 2098 1131 2102
rect 1151 2098 1155 2102
rect 1255 2098 1259 2102
rect 1327 2098 1331 2102
rect 1367 2098 1371 2102
rect 1431 2098 1435 2102
rect 1519 2098 1523 2102
rect 1535 2098 1539 2102
rect 1615 2098 1619 2102
rect 1647 2098 1651 2102
rect 671 2072 675 2076
rect 1719 2098 1723 2102
rect 1759 2098 1763 2102
rect 1823 2098 1827 2102
rect 1367 2042 1371 2046
rect 1415 2042 1419 2046
rect 111 2034 115 2038
rect 279 2034 283 2038
rect 343 2034 347 2038
rect 415 2034 419 2038
rect 471 2034 475 2038
rect 495 2034 499 2038
rect 527 2034 531 2038
rect 583 2034 587 2038
rect 639 2034 643 2038
rect 671 2034 675 2038
rect 695 2034 699 2038
rect 751 2034 755 2038
rect 807 2034 811 2038
rect 831 2034 835 2038
rect 863 2034 867 2038
rect 903 2034 907 2038
rect 919 2034 923 2038
rect 975 2034 979 2038
rect 983 2034 987 2038
rect 1031 2034 1035 2038
rect 111 1974 115 1978
rect 335 1974 339 1978
rect 391 1974 395 1978
rect 399 1974 403 1978
rect 447 1974 451 1978
rect 455 1974 459 1978
rect 503 1974 507 1978
rect 511 1974 515 1978
rect 567 1974 571 1978
rect 111 1918 115 1922
rect 159 1918 163 1922
rect 231 1918 235 1922
rect 327 1918 331 1922
rect 351 1918 355 1922
rect 407 1918 411 1922
rect 431 1918 435 1922
rect 463 1918 467 1922
rect 743 1992 747 1996
rect 1063 2034 1067 2038
rect 1143 2034 1147 2038
rect 1327 2034 1331 2038
rect 1447 2042 1451 2046
rect 1503 2042 1507 2046
rect 1551 2042 1555 2046
rect 1607 2042 1611 2046
rect 1663 2042 1667 2046
rect 1711 2042 1715 2046
rect 1775 2042 1779 2046
rect 2111 2154 2115 2158
rect 2159 2154 2163 2158
rect 2223 2154 2227 2158
rect 2263 2154 2267 2158
rect 2327 2154 2331 2158
rect 2359 2154 2363 2158
rect 2439 2154 2443 2158
rect 2463 2154 2467 2158
rect 2543 2154 2547 2158
rect 1863 2098 1867 2102
rect 1935 2098 1939 2102
rect 1967 2098 1971 2102
rect 2039 2098 2043 2102
rect 2071 2098 2075 2102
rect 2143 2098 2147 2102
rect 2175 2098 2179 2102
rect 2247 2098 2251 2102
rect 2271 2098 2275 2102
rect 1807 2042 1811 2046
rect 1879 2042 1883 2046
rect 1903 2042 1907 2046
rect 1983 2042 1987 2046
rect 2343 2098 2347 2102
rect 2359 2098 2363 2102
rect 2447 2098 2451 2102
rect 2455 2098 2459 2102
rect 2007 2042 2011 2046
rect 1175 1992 1179 1996
rect 623 1974 627 1978
rect 647 1974 651 1978
rect 679 1974 683 1978
rect 735 1974 739 1978
rect 743 1974 747 1978
rect 791 1974 795 1978
rect 847 1974 851 1978
rect 863 1974 867 1978
rect 903 1974 907 1978
rect 959 1974 963 1978
rect 999 1974 1003 1978
rect 1015 1974 1019 1978
rect 1143 1974 1147 1978
rect 519 1918 523 1922
rect 543 1918 547 1922
rect 583 1918 587 1922
rect 655 1918 659 1922
rect 1367 1986 1371 1990
rect 1399 1986 1403 1990
rect 1479 1986 1483 1990
rect 1487 1986 1491 1990
rect 1271 1974 1275 1978
rect 1327 1974 1331 1978
rect 1583 1986 1587 1990
rect 1591 1986 1595 1990
rect 1679 1986 1683 1990
rect 1695 1986 1699 1990
rect 1367 1926 1371 1930
rect 1415 1926 1419 1930
rect 1495 1926 1499 1930
rect 1599 1926 1603 1930
rect 1695 1926 1699 1930
rect 1767 1986 1771 1990
rect 1791 1986 1795 1990
rect 1847 1986 1851 1990
rect 1887 1986 1891 1990
rect 2087 2042 2091 2046
rect 2111 2042 2115 2046
rect 2191 2042 2195 2046
rect 2215 2042 2219 2046
rect 2287 2042 2291 2046
rect 2327 2042 2331 2046
rect 2375 2042 2379 2046
rect 2527 2098 2531 2102
rect 2583 2154 2587 2158
rect 2583 2098 2587 2102
rect 2447 2042 2451 2046
rect 2471 2042 2475 2046
rect 2543 2042 2547 2046
rect 2583 2042 2587 2046
rect 1927 1986 1931 1990
rect 1991 1986 1995 1990
rect 2007 1986 2011 1990
rect 2087 1986 2091 1990
rect 2095 1986 2099 1990
rect 2199 1986 2203 1990
rect 2311 1986 2315 1990
rect 2431 1986 2435 1990
rect 2527 1986 2531 1990
rect 2583 1986 2587 1990
rect 663 1918 667 1922
rect 111 1854 115 1858
rect 143 1854 147 1858
rect 759 1918 763 1922
rect 767 1918 771 1922
rect 879 1918 883 1922
rect 983 1918 987 1922
rect 1015 1918 1019 1922
rect 1087 1918 1091 1922
rect 1159 1918 1163 1922
rect 1199 1918 1203 1922
rect 199 1854 203 1858
rect 215 1854 219 1858
rect 263 1854 267 1858
rect 311 1854 315 1858
rect 351 1854 355 1858
rect 415 1854 419 1858
rect 439 1854 443 1858
rect 527 1854 531 1858
rect 535 1854 539 1858
rect 623 1854 627 1858
rect 639 1854 643 1858
rect 711 1854 715 1858
rect 751 1854 755 1858
rect 791 1854 795 1858
rect 863 1854 867 1858
rect 871 1854 875 1858
rect 951 1854 955 1858
rect 967 1854 971 1858
rect 111 1794 115 1798
rect 159 1794 163 1798
rect 215 1794 219 1798
rect 231 1794 235 1798
rect 279 1794 283 1798
rect 295 1794 299 1798
rect 367 1794 371 1798
rect 447 1794 451 1798
rect 455 1794 459 1798
rect 535 1794 539 1798
rect 551 1794 555 1798
rect 623 1794 627 1798
rect 111 1734 115 1738
rect 215 1734 219 1738
rect 279 1734 283 1738
rect 351 1734 355 1738
rect 1287 1918 1291 1922
rect 1327 1918 1331 1922
rect 1719 1926 1723 1930
rect 1775 1926 1779 1930
rect 1783 1926 1787 1930
rect 1831 1926 1835 1930
rect 1863 1926 1867 1930
rect 1887 1926 1891 1930
rect 1943 1926 1947 1930
rect 1999 1926 2003 1930
rect 1367 1866 1371 1870
rect 1399 1866 1403 1870
rect 1463 1866 1467 1870
rect 1559 1866 1563 1870
rect 1655 1866 1659 1870
rect 1703 1866 1707 1870
rect 1743 1866 1747 1870
rect 1759 1866 1763 1870
rect 1039 1854 1043 1858
rect 1071 1854 1075 1858
rect 1183 1854 1187 1858
rect 1271 1854 1275 1858
rect 1327 1854 1331 1858
rect 639 1794 643 1798
rect 711 1794 715 1798
rect 727 1794 731 1798
rect 791 1794 795 1798
rect 807 1794 811 1798
rect 871 1794 875 1798
rect 887 1794 891 1798
rect 951 1794 955 1798
rect 407 1734 411 1738
rect 431 1734 435 1738
rect 471 1734 475 1738
rect 519 1734 523 1738
rect 551 1734 555 1738
rect 607 1734 611 1738
rect 639 1734 643 1738
rect 695 1734 699 1738
rect 727 1734 731 1738
rect 775 1734 779 1738
rect 823 1734 827 1738
rect 855 1734 859 1738
rect 1367 1810 1371 1814
rect 1415 1810 1419 1814
rect 1479 1810 1483 1814
rect 1511 1810 1515 1814
rect 1575 1810 1579 1814
rect 1623 1810 1627 1814
rect 967 1794 971 1798
rect 1031 1794 1035 1798
rect 1055 1794 1059 1798
rect 1119 1794 1123 1798
rect 1327 1794 1331 1798
rect 1367 1754 1371 1758
rect 1399 1754 1403 1758
rect 1671 1810 1675 1814
rect 2023 1926 2027 1930
rect 2055 1926 2059 1930
rect 2103 1926 2107 1930
rect 2119 1926 2123 1930
rect 2583 1926 2587 1930
rect 1815 1866 1819 1870
rect 1831 1866 1835 1870
rect 1871 1866 1875 1870
rect 1919 1866 1923 1870
rect 1927 1866 1931 1870
rect 1983 1866 1987 1870
rect 2007 1866 2011 1870
rect 1827 1824 1831 1828
rect 1735 1810 1739 1814
rect 2039 1866 2043 1870
rect 2095 1866 2099 1870
rect 2103 1866 2107 1870
rect 2183 1866 2187 1870
rect 2583 1866 2587 1870
rect 2207 1824 2211 1828
rect 1759 1810 1763 1814
rect 1839 1810 1843 1814
rect 1847 1810 1851 1814
rect 1935 1810 1939 1814
rect 1951 1810 1955 1814
rect 2023 1810 2027 1814
rect 2063 1810 2067 1814
rect 1439 1754 1443 1758
rect 1495 1754 1499 1758
rect 1519 1754 1523 1758
rect 1607 1754 1611 1758
rect 1615 1754 1619 1758
rect 1719 1754 1723 1758
rect 1823 1754 1827 1758
rect 919 1734 923 1738
rect 935 1734 939 1738
rect 1015 1734 1019 1738
rect 1103 1734 1107 1738
rect 1111 1734 1115 1738
rect 1207 1734 1211 1738
rect 1327 1734 1331 1738
rect 111 1674 115 1678
rect 367 1674 371 1678
rect 399 1674 403 1678
rect 423 1674 427 1678
rect 455 1674 459 1678
rect 487 1674 491 1678
rect 511 1674 515 1678
rect 567 1674 571 1678
rect 575 1674 579 1678
rect 647 1674 651 1678
rect 655 1674 659 1678
rect 727 1674 731 1678
rect 743 1674 747 1678
rect 807 1674 811 1678
rect 839 1674 843 1678
rect 887 1674 891 1678
rect 935 1674 939 1678
rect 967 1674 971 1678
rect 111 1602 115 1606
rect 287 1602 291 1606
rect 367 1602 371 1606
rect 383 1602 387 1606
rect 439 1602 443 1606
rect 455 1602 459 1606
rect 495 1602 499 1606
rect 551 1602 555 1606
rect 559 1602 563 1606
rect 631 1602 635 1606
rect 647 1602 651 1606
rect 711 1602 715 1606
rect 735 1602 739 1606
rect 791 1602 795 1606
rect 823 1602 827 1606
rect 111 1546 115 1550
rect 279 1546 283 1550
rect 303 1546 307 1550
rect 335 1546 339 1550
rect 383 1546 387 1550
rect 399 1546 403 1550
rect 1031 1674 1035 1678
rect 1047 1674 1051 1678
rect 1127 1674 1131 1678
rect 1135 1674 1139 1678
rect 1223 1674 1227 1678
rect 1367 1686 1371 1690
rect 1455 1686 1459 1690
rect 1535 1686 1539 1690
rect 1559 1686 1563 1690
rect 1631 1686 1635 1690
rect 1711 1686 1715 1690
rect 1287 1674 1291 1678
rect 1327 1674 1331 1678
rect 871 1602 875 1606
rect 903 1602 907 1606
rect 951 1602 955 1606
rect 983 1602 987 1606
rect 1031 1602 1035 1606
rect 1063 1602 1067 1606
rect 1119 1602 1123 1606
rect 471 1546 475 1550
rect 111 1486 115 1490
rect 199 1486 203 1490
rect 263 1486 267 1490
rect 287 1486 291 1490
rect 319 1486 323 1490
rect 383 1486 387 1490
rect 111 1426 115 1430
rect 159 1426 163 1430
rect 543 1546 547 1550
rect 567 1546 571 1550
rect 615 1546 619 1550
rect 663 1546 667 1550
rect 687 1546 691 1550
rect 455 1486 459 1490
rect 487 1486 491 1490
rect 527 1486 531 1490
rect 751 1546 755 1550
rect 759 1546 763 1550
rect 831 1546 835 1550
rect 839 1546 843 1550
rect 903 1546 907 1550
rect 919 1546 923 1550
rect 975 1546 979 1550
rect 999 1546 1003 1550
rect 1367 1618 1371 1622
rect 1543 1618 1547 1622
rect 1151 1602 1155 1606
rect 1207 1602 1211 1606
rect 1271 1602 1275 1606
rect 1327 1602 1331 1606
rect 1735 1686 1739 1690
rect 2111 1810 2115 1814
rect 2183 1810 2187 1814
rect 2199 1810 2203 1814
rect 2303 1810 2307 1814
rect 2431 1810 2435 1814
rect 2543 1810 2547 1814
rect 2583 1810 2587 1814
rect 1927 1754 1931 1758
rect 1935 1754 1939 1758
rect 2023 1754 2027 1758
rect 2047 1754 2051 1758
rect 2119 1754 2123 1758
rect 2167 1754 2171 1758
rect 2207 1754 2211 1758
rect 2287 1754 2291 1758
rect 2375 1754 2379 1758
rect 2415 1754 2419 1758
rect 2463 1754 2467 1758
rect 2019 1712 2023 1716
rect 1799 1686 1803 1690
rect 1839 1686 1843 1690
rect 1887 1686 1891 1690
rect 1943 1686 1947 1690
rect 1975 1686 1979 1690
rect 2039 1686 2043 1690
rect 2063 1686 2067 1690
rect 2135 1686 2139 1690
rect 2143 1686 2147 1690
rect 2215 1686 2219 1690
rect 2223 1686 2227 1690
rect 1575 1618 1579 1622
rect 1615 1618 1619 1622
rect 1631 1618 1635 1622
rect 1687 1618 1691 1622
rect 1695 1618 1699 1622
rect 1751 1618 1755 1622
rect 1783 1618 1787 1622
rect 1831 1618 1835 1622
rect 1871 1618 1875 1622
rect 1919 1618 1923 1622
rect 1959 1618 1963 1622
rect 1367 1558 1371 1562
rect 1591 1558 1595 1562
rect 1647 1558 1651 1562
rect 1679 1558 1683 1562
rect 1703 1558 1707 1562
rect 1735 1558 1739 1562
rect 1767 1558 1771 1562
rect 1791 1558 1795 1562
rect 1847 1558 1851 1562
rect 1855 1558 1859 1562
rect 1055 1546 1059 1550
rect 1079 1546 1083 1550
rect 1167 1546 1171 1550
rect 1327 1546 1331 1550
rect 583 1486 587 1490
rect 599 1486 603 1490
rect 671 1486 675 1490
rect 679 1486 683 1490
rect 743 1486 747 1490
rect 775 1486 779 1490
rect 815 1486 819 1490
rect 863 1486 867 1490
rect 887 1486 891 1490
rect 215 1426 219 1430
rect 247 1426 251 1430
rect 303 1426 307 1430
rect 343 1426 347 1430
rect 399 1426 403 1430
rect 111 1370 115 1374
rect 143 1370 147 1374
rect 207 1370 211 1374
rect 231 1370 235 1374
rect 295 1370 299 1374
rect 327 1370 331 1374
rect 447 1426 451 1430
rect 503 1426 507 1430
rect 551 1426 555 1430
rect 599 1426 603 1430
rect 663 1426 667 1430
rect 695 1426 699 1430
rect 399 1370 403 1374
rect 431 1370 435 1374
rect 511 1370 515 1374
rect 535 1370 539 1374
rect 623 1370 627 1374
rect 647 1370 651 1374
rect 111 1314 115 1318
rect 159 1314 163 1318
rect 223 1314 227 1318
rect 231 1314 235 1318
rect 311 1314 315 1318
rect 327 1314 331 1318
rect 415 1314 419 1318
rect 111 1246 115 1250
rect 143 1246 147 1250
rect 199 1246 203 1250
rect 215 1246 219 1250
rect 279 1246 283 1250
rect 431 1314 435 1318
rect 1367 1494 1371 1498
rect 1519 1494 1523 1498
rect 1575 1494 1579 1498
rect 1647 1494 1651 1498
rect 1663 1494 1667 1498
rect 951 1486 955 1490
rect 959 1486 963 1490
rect 1039 1486 1043 1490
rect 1135 1486 1139 1490
rect 1327 1486 1331 1490
rect 767 1426 771 1430
rect 791 1426 795 1430
rect 879 1426 883 1430
rect 967 1426 971 1430
rect 991 1426 995 1430
rect 1055 1426 1059 1430
rect 1103 1426 1107 1430
rect 1151 1426 1155 1430
rect 735 1370 739 1374
rect 751 1370 755 1374
rect 847 1370 851 1374
rect 863 1370 867 1374
rect 2399 1712 2403 1716
rect 2527 1754 2531 1758
rect 2583 1754 2587 1758
rect 2287 1686 2291 1690
rect 2303 1686 2307 1690
rect 2351 1686 2355 1690
rect 2391 1686 2395 1690
rect 2423 1686 2427 1690
rect 2479 1686 2483 1690
rect 2487 1686 2491 1690
rect 2543 1686 2547 1690
rect 2007 1618 2011 1622
rect 2047 1618 2051 1622
rect 2103 1618 2107 1622
rect 2127 1618 2131 1622
rect 2199 1618 2203 1622
rect 2207 1618 2211 1622
rect 2271 1618 2275 1622
rect 2319 1618 2323 1622
rect 2335 1618 2339 1622
rect 2407 1618 2411 1622
rect 2431 1618 2435 1622
rect 2471 1618 2475 1622
rect 2527 1618 2531 1622
rect 1927 1558 1931 1562
rect 1935 1558 1939 1562
rect 2007 1558 2011 1562
rect 2023 1558 2027 1562
rect 2087 1558 2091 1562
rect 2119 1558 2123 1562
rect 2583 1686 2587 1690
rect 2583 1618 2587 1622
rect 2167 1558 2171 1562
rect 2223 1558 2227 1562
rect 2247 1558 2251 1562
rect 2327 1558 2331 1562
rect 2335 1558 2339 1562
rect 2407 1558 2411 1562
rect 1719 1494 1723 1498
rect 1727 1494 1731 1498
rect 1775 1494 1779 1498
rect 1807 1494 1811 1498
rect 1839 1494 1843 1498
rect 1895 1494 1899 1498
rect 1911 1494 1915 1498
rect 1983 1494 1987 1498
rect 1991 1494 1995 1498
rect 2071 1494 2075 1498
rect 2151 1494 2155 1498
rect 2231 1494 2235 1498
rect 1215 1426 1219 1430
rect 1327 1426 1331 1430
rect 1367 1430 1371 1434
rect 1415 1430 1419 1434
rect 1471 1430 1475 1434
rect 1535 1430 1539 1434
rect 1591 1430 1595 1434
rect 1623 1430 1627 1434
rect 1663 1430 1667 1434
rect 1719 1430 1723 1434
rect 1743 1430 1747 1434
rect 1823 1430 1827 1434
rect 959 1370 963 1374
rect 975 1370 979 1374
rect 891 1328 895 1332
rect 527 1314 531 1318
rect 535 1314 539 1318
rect 631 1314 635 1318
rect 639 1314 643 1318
rect 727 1314 731 1318
rect 311 1246 315 1250
rect 359 1246 363 1250
rect 415 1246 419 1250
rect 439 1246 443 1250
rect 519 1246 523 1250
rect 111 1186 115 1190
rect 159 1186 163 1190
rect 215 1186 219 1190
rect 239 1186 243 1190
rect 295 1186 299 1190
rect 327 1186 331 1190
rect 375 1186 379 1190
rect 423 1186 427 1190
rect 455 1186 459 1190
rect 751 1314 755 1318
rect 823 1314 827 1318
rect 863 1314 867 1318
rect 1071 1370 1075 1374
rect 1087 1370 1091 1374
rect 1183 1370 1187 1374
rect 1199 1370 1203 1374
rect 1271 1370 1275 1374
rect 1327 1370 1331 1374
rect 911 1314 915 1318
rect 975 1314 979 1318
rect 1367 1366 1371 1370
rect 1399 1366 1403 1370
rect 1911 1430 1915 1434
rect 1927 1430 1931 1434
rect 1999 1430 2003 1434
rect 2023 1430 2027 1434
rect 2447 1558 2451 1562
rect 2487 1558 2491 1562
rect 2543 1558 2547 1562
rect 2311 1494 2315 1498
rect 2391 1494 2395 1498
rect 2087 1430 2091 1434
rect 2119 1430 2123 1434
rect 2167 1430 2171 1434
rect 1455 1366 1459 1370
rect 1519 1366 1523 1370
rect 1543 1366 1547 1370
rect 1607 1366 1611 1370
rect 1631 1366 1635 1370
rect 1703 1366 1707 1370
rect 1719 1366 1723 1370
rect 1807 1366 1811 1370
rect 1887 1366 1891 1370
rect 1911 1366 1915 1370
rect 1407 1352 1411 1356
rect 1295 1328 1299 1332
rect 991 1314 995 1318
rect 1071 1314 1075 1318
rect 1087 1314 1091 1318
rect 1151 1314 1155 1318
rect 1199 1314 1203 1318
rect 1231 1314 1235 1318
rect 1287 1314 1291 1318
rect 1327 1314 1331 1318
rect 599 1246 603 1250
rect 615 1246 619 1250
rect 671 1246 675 1250
rect 711 1246 715 1250
rect 743 1246 747 1250
rect 1751 1355 1755 1356
rect 1751 1352 1755 1355
rect 1367 1306 1371 1310
rect 1415 1306 1419 1310
rect 1471 1306 1475 1310
rect 1559 1306 1563 1310
rect 1647 1306 1651 1310
rect 1671 1306 1675 1310
rect 1735 1306 1739 1310
rect 1767 1306 1771 1310
rect 1823 1306 1827 1310
rect 2215 1430 2219 1434
rect 2247 1430 2251 1434
rect 2471 1494 2475 1498
rect 2527 1494 2531 1498
rect 2583 1558 2587 1562
rect 2583 1494 2587 1498
rect 2303 1430 2307 1434
rect 2327 1430 2331 1434
rect 2391 1430 2395 1434
rect 2407 1430 2411 1434
rect 2479 1430 2483 1434
rect 2487 1430 2491 1434
rect 2543 1430 2547 1434
rect 1967 1366 1971 1370
rect 2007 1366 2011 1370
rect 2047 1366 2051 1370
rect 2103 1366 2107 1370
rect 2127 1366 2131 1370
rect 2199 1366 2203 1370
rect 2207 1366 2211 1370
rect 1863 1306 1867 1310
rect 1903 1306 1907 1310
rect 1959 1306 1963 1310
rect 807 1246 811 1250
rect 815 1246 819 1250
rect 895 1246 899 1250
rect 975 1246 979 1250
rect 1055 1246 1059 1250
rect 1135 1246 1139 1250
rect 1215 1246 1219 1250
rect 1271 1246 1275 1250
rect 1327 1246 1331 1250
rect 1367 1250 1371 1254
rect 1495 1250 1499 1254
rect 1559 1250 1563 1254
rect 1623 1250 1627 1254
rect 1655 1250 1659 1254
rect 511 1186 515 1190
rect 535 1186 539 1190
rect 599 1186 603 1190
rect 615 1186 619 1190
rect 687 1186 691 1190
rect 759 1186 763 1190
rect 767 1186 771 1190
rect 831 1186 835 1190
rect 839 1186 843 1190
rect 111 1122 115 1126
rect 143 1122 147 1126
rect 223 1122 227 1126
rect 311 1122 315 1126
rect 319 1122 323 1126
rect 407 1122 411 1126
rect 423 1122 427 1126
rect 495 1122 499 1126
rect 527 1122 531 1126
rect 583 1122 587 1126
rect 219 1080 223 1084
rect 551 1080 555 1084
rect 111 1062 115 1066
rect 239 1062 243 1066
rect 311 1062 315 1066
rect 335 1062 339 1066
rect 367 1062 371 1066
rect 439 1062 443 1066
rect 911 1186 915 1190
rect 983 1186 987 1190
rect 1063 1186 1067 1190
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1415 1186 1419 1190
rect 1503 1186 1507 1190
rect 1511 1186 1515 1190
rect 1575 1186 1579 1190
rect 1687 1250 1691 1254
rect 1751 1250 1755 1254
rect 1759 1250 1763 1254
rect 2583 1430 2587 1434
rect 2287 1366 2291 1370
rect 2375 1366 2379 1370
rect 2463 1366 2467 1370
rect 2527 1366 2531 1370
rect 2583 1366 2587 1370
rect 1983 1306 1987 1310
rect 2047 1306 2051 1310
rect 2063 1306 2067 1310
rect 1823 1250 1827 1254
rect 1847 1250 1851 1254
rect 1887 1250 1891 1254
rect 2135 1306 2139 1310
rect 2143 1306 2147 1310
rect 2223 1306 2227 1310
rect 2231 1306 2235 1310
rect 2583 1306 2587 1310
rect 1943 1250 1947 1254
rect 1951 1250 1955 1254
rect 2015 1250 2019 1254
rect 2031 1250 2035 1254
rect 2079 1250 2083 1254
rect 2119 1250 2123 1254
rect 2151 1250 2155 1254
rect 1599 1186 1603 1190
rect 1639 1186 1643 1190
rect 1703 1186 1707 1190
rect 1775 1186 1779 1190
rect 1807 1186 1811 1190
rect 1839 1186 1843 1190
rect 1903 1186 1907 1190
rect 1911 1186 1915 1190
rect 631 1122 635 1126
rect 671 1122 675 1126
rect 727 1122 731 1126
rect 751 1122 755 1126
rect 823 1122 827 1126
rect 895 1122 899 1126
rect 911 1122 915 1126
rect 967 1122 971 1126
rect 991 1122 995 1126
rect 1047 1122 1051 1126
rect 1079 1122 1083 1126
rect 1167 1122 1171 1126
rect 1327 1122 1331 1126
rect 1367 1126 1371 1130
rect 1399 1126 1403 1130
rect 519 1062 523 1066
rect 543 1062 547 1066
rect 607 1062 611 1066
rect 647 1062 651 1066
rect 703 1062 707 1066
rect 743 1062 747 1066
rect 799 1062 803 1066
rect 839 1062 843 1066
rect 887 1062 891 1066
rect 927 1062 931 1066
rect 975 1062 979 1066
rect 1007 1062 1011 1066
rect 1055 1062 1059 1066
rect 111 1002 115 1006
rect 295 1002 299 1006
rect 351 1002 355 1006
rect 415 1002 419 1006
rect 423 1002 427 1006
rect 471 1002 475 1006
rect 503 1002 507 1006
rect 527 1002 531 1006
rect 879 1024 883 1028
rect 591 1002 595 1006
rect 655 1002 659 1006
rect 687 1002 691 1006
rect 719 1002 723 1006
rect 111 942 115 946
rect 423 942 427 946
rect 431 942 435 946
rect 479 942 483 946
rect 487 942 491 946
rect 535 942 539 946
rect 543 942 547 946
rect 591 942 595 946
rect 607 942 611 946
rect 647 942 651 946
rect 111 886 115 890
rect 279 886 283 890
rect 335 886 339 890
rect 391 886 395 890
rect 407 886 411 890
rect 671 942 675 946
rect 703 942 707 946
rect 735 942 739 946
rect 1479 1126 1483 1130
rect 1487 1126 1491 1130
rect 1583 1126 1587 1130
rect 1967 1186 1971 1190
rect 2015 1186 2019 1190
rect 2031 1186 2035 1190
rect 2215 1250 2219 1254
rect 2223 1250 2227 1254
rect 2295 1250 2299 1254
rect 2583 1250 2587 1254
rect 2095 1186 2099 1190
rect 2111 1186 2115 1190
rect 2167 1186 2171 1190
rect 2207 1186 2211 1190
rect 2239 1186 2243 1190
rect 2303 1186 2307 1190
rect 2311 1186 2315 1190
rect 2399 1186 2403 1190
rect 2583 1186 2587 1190
rect 1687 1126 1691 1130
rect 1791 1126 1795 1130
rect 1887 1126 1891 1130
rect 1895 1126 1899 1130
rect 1975 1126 1979 1130
rect 1999 1126 2003 1130
rect 2063 1126 2067 1130
rect 2095 1126 2099 1130
rect 2143 1126 2147 1130
rect 2191 1126 2195 1130
rect 2215 1126 2219 1130
rect 2279 1126 2283 1130
rect 2287 1126 2291 1130
rect 1095 1062 1099 1066
rect 1135 1062 1139 1066
rect 1183 1062 1187 1066
rect 1223 1062 1227 1066
rect 1287 1062 1291 1066
rect 1327 1062 1331 1066
rect 1367 1066 1371 1070
rect 1415 1066 1419 1070
rect 1471 1066 1475 1070
rect 1495 1066 1499 1070
rect 1535 1066 1539 1070
rect 1599 1066 1603 1070
rect 1623 1066 1627 1070
rect 1703 1066 1707 1070
rect 1727 1066 1731 1070
rect 1807 1066 1811 1070
rect 1839 1066 1843 1070
rect 1235 1024 1239 1028
rect 783 1002 787 1006
rect 847 1002 851 1006
rect 871 1002 875 1006
rect 911 1002 915 1006
rect 959 1002 963 1006
rect 975 1002 979 1006
rect 1039 1002 1043 1006
rect 1103 1002 1107 1006
rect 1119 1002 1123 1006
rect 1159 1002 1163 1006
rect 1207 1002 1211 1006
rect 1215 1002 1219 1006
rect 1271 1002 1275 1006
rect 1327 1002 1331 1006
rect 1367 994 1371 998
rect 1399 994 1403 998
rect 1455 994 1459 998
rect 1511 994 1515 998
rect 1519 994 1523 998
rect 759 942 763 946
rect 799 942 803 946
rect 815 942 819 946
rect 863 942 867 946
rect 927 942 931 946
rect 991 942 995 946
rect 1055 942 1059 946
rect 1119 942 1123 946
rect 1175 942 1179 946
rect 1231 942 1235 946
rect 1287 942 1291 946
rect 1327 942 1331 946
rect 1903 1066 1907 1070
rect 1951 1066 1955 1070
rect 1991 1066 1995 1070
rect 2063 1066 2067 1070
rect 2079 1066 2083 1070
rect 2343 1126 2347 1130
rect 2383 1126 2387 1130
rect 2407 1126 2411 1130
rect 2471 1126 2475 1130
rect 2527 1126 2531 1130
rect 2583 1126 2587 1130
rect 2159 1066 2163 1070
rect 2167 1066 2171 1070
rect 2231 1066 2235 1070
rect 2271 1066 2275 1070
rect 2295 1066 2299 1070
rect 2359 1066 2363 1070
rect 2367 1066 2371 1070
rect 2423 1066 2427 1070
rect 2463 1066 2467 1070
rect 2487 1066 2491 1070
rect 2543 1066 2547 1070
rect 2583 1066 2587 1070
rect 1567 994 1571 998
rect 1607 994 1611 998
rect 1639 994 1643 998
rect 1711 994 1715 998
rect 1719 994 1723 998
rect 1807 994 1811 998
rect 1823 994 1827 998
rect 1903 994 1907 998
rect 1935 994 1939 998
rect 2015 994 2019 998
rect 2047 994 2051 998
rect 2143 994 2147 998
rect 2151 994 2155 998
rect 2255 994 2259 998
rect 2271 994 2275 998
rect 2351 994 2355 998
rect 2407 994 2411 998
rect 2447 994 2451 998
rect 2527 994 2531 998
rect 1367 930 1371 934
rect 1415 930 1419 934
rect 455 886 459 890
rect 463 886 467 890
rect 519 886 523 890
rect 575 886 579 890
rect 583 886 587 890
rect 631 886 635 890
rect 647 886 651 890
rect 687 886 691 890
rect 2583 994 2587 998
rect 1471 930 1475 934
rect 1527 930 1531 934
rect 711 886 715 890
rect 743 886 747 890
rect 775 886 779 890
rect 799 886 803 890
rect 847 886 851 890
rect 919 886 923 890
rect 1327 886 1331 890
rect 1583 930 1587 934
rect 1615 930 1619 934
rect 1655 930 1659 934
rect 1711 930 1715 934
rect 1735 930 1739 934
rect 1823 930 1827 934
rect 1919 930 1923 934
rect 1943 930 1947 934
rect 2031 930 2035 934
rect 2063 930 2067 934
rect 2159 930 2163 934
rect 2183 930 2187 934
rect 2287 930 2291 934
rect 2311 930 2315 934
rect 1367 874 1371 878
rect 1399 874 1403 878
rect 1455 874 1459 878
rect 1471 874 1475 878
rect 1511 874 1515 878
rect 1551 874 1555 878
rect 1599 874 1603 878
rect 1639 874 1643 878
rect 1695 874 1699 878
rect 1727 874 1731 878
rect 1807 874 1811 878
rect 1815 874 1819 878
rect 1903 874 1907 878
rect 1927 874 1931 878
rect 111 822 115 826
rect 167 822 171 826
rect 231 822 235 826
rect 295 822 299 826
rect 311 822 315 826
rect 351 822 355 826
rect 399 822 403 826
rect 407 822 411 826
rect 471 822 475 826
rect 487 822 491 826
rect 535 822 539 826
rect 583 822 587 826
rect 111 758 115 762
rect 143 758 147 762
rect 151 758 155 762
rect 599 822 603 826
rect 663 822 667 826
rect 671 822 675 826
rect 727 822 731 826
rect 759 822 763 826
rect 791 822 795 826
rect 839 822 843 826
rect 863 822 867 826
rect 919 822 923 826
rect 935 822 939 826
rect 1007 822 1011 826
rect 1095 822 1099 826
rect 1327 822 1331 826
rect 1367 810 1371 814
rect 1487 810 1491 814
rect 1567 810 1571 814
rect 1631 810 1635 814
rect 1655 810 1659 814
rect 1687 810 1691 814
rect 1743 810 1747 814
rect 1751 810 1755 814
rect 199 758 203 762
rect 215 758 219 762
rect 279 758 283 762
rect 295 758 299 762
rect 383 758 387 762
rect 471 758 475 762
rect 487 758 491 762
rect 567 758 571 762
rect 599 758 603 762
rect 655 758 659 762
rect 703 758 707 762
rect 743 758 747 762
rect 807 758 811 762
rect 823 758 827 762
rect 903 758 907 762
rect 991 758 995 762
rect 1079 758 1083 762
rect 699 712 703 716
rect 1175 758 1179 762
rect 1327 758 1331 762
rect 1103 712 1107 716
rect 2423 930 2427 934
rect 2439 930 2443 934
rect 2543 930 2547 934
rect 2583 930 2587 934
rect 1991 874 1995 878
rect 2047 874 2051 878
rect 2071 874 2075 878
rect 2143 874 2147 878
rect 2167 874 2171 878
rect 2215 874 2219 878
rect 2279 874 2283 878
rect 2295 874 2299 878
rect 2343 874 2347 878
rect 2407 874 2411 878
rect 2423 874 2427 878
rect 2471 874 2475 878
rect 2527 874 2531 878
rect 1823 810 1827 814
rect 1831 810 1835 814
rect 1903 810 1907 814
rect 1919 810 1923 814
rect 1991 810 1995 814
rect 2007 810 2011 814
rect 2071 810 2075 814
rect 2087 810 2091 814
rect 2583 874 2587 878
rect 2159 810 2163 814
rect 2231 810 2235 814
rect 2247 810 2251 814
rect 2295 810 2299 814
rect 2335 810 2339 814
rect 2359 810 2363 814
rect 2423 810 2427 814
rect 2487 810 2491 814
rect 2543 810 2547 814
rect 2583 810 2587 814
rect 2127 776 2131 780
rect 1367 750 1371 754
rect 1567 750 1571 754
rect 1615 750 1619 754
rect 1623 750 1627 754
rect 1671 750 1675 754
rect 1687 750 1691 754
rect 1735 750 1739 754
rect 1759 750 1763 754
rect 1807 750 1811 754
rect 1839 750 1843 754
rect 1887 750 1891 754
rect 1919 750 1923 754
rect 1975 750 1979 754
rect 1999 750 2003 754
rect 2055 750 2059 754
rect 2079 750 2083 754
rect 111 698 115 702
rect 159 698 163 702
rect 215 698 219 702
rect 279 698 283 702
rect 295 698 299 702
rect 359 698 363 702
rect 399 698 403 702
rect 447 698 451 702
rect 503 698 507 702
rect 535 698 539 702
rect 615 698 619 702
rect 623 698 627 702
rect 711 698 715 702
rect 719 698 723 702
rect 791 698 795 702
rect 823 698 827 702
rect 871 698 875 702
rect 919 698 923 702
rect 111 634 115 638
rect 143 634 147 638
rect 199 634 203 638
rect 255 634 259 638
rect 263 634 267 638
rect 311 634 315 638
rect 343 634 347 638
rect 391 634 395 638
rect 431 634 435 638
rect 479 634 483 638
rect 519 634 523 638
rect 575 634 579 638
rect 607 634 611 638
rect 111 574 115 578
rect 159 574 163 578
rect 199 574 203 578
rect 215 574 219 578
rect 263 574 267 578
rect 271 574 275 578
rect 327 574 331 578
rect 335 574 339 578
rect 951 698 955 702
rect 1007 698 1011 702
rect 1039 698 1043 702
rect 1095 698 1099 702
rect 1191 698 1195 702
rect 1327 698 1331 702
rect 2143 750 2147 754
rect 2439 776 2443 780
rect 2159 750 2163 754
rect 2231 750 2235 754
rect 2247 750 2251 754
rect 2319 750 2323 754
rect 2335 750 2339 754
rect 2407 750 2411 754
rect 2583 750 2587 754
rect 1367 690 1371 694
rect 1415 690 1419 694
rect 1511 690 1515 694
rect 1583 690 1587 694
rect 1615 690 1619 694
rect 1639 690 1643 694
rect 1703 690 1707 694
rect 1719 690 1723 694
rect 1775 690 1779 694
rect 1823 690 1827 694
rect 1855 690 1859 694
rect 679 634 683 638
rect 695 634 699 638
rect 775 634 779 638
rect 783 634 787 638
rect 855 634 859 638
rect 887 634 891 638
rect 935 634 939 638
rect 991 634 995 638
rect 1023 634 1027 638
rect 1087 634 1091 638
rect 1191 634 1195 638
rect 1271 634 1275 638
rect 1327 634 1331 638
rect 1367 634 1371 638
rect 1399 634 1403 638
rect 407 574 411 578
rect 415 574 419 578
rect 495 574 499 578
rect 511 574 515 578
rect 591 574 595 578
rect 615 574 619 578
rect 695 574 699 578
rect 719 574 723 578
rect 799 574 803 578
rect 831 574 835 578
rect 903 574 907 578
rect 943 574 947 578
rect 1007 574 1011 578
rect 1063 574 1067 578
rect 111 510 115 514
rect 183 510 187 514
rect 247 510 251 514
rect 303 510 307 514
rect 319 510 323 514
rect 359 510 363 514
rect 399 510 403 514
rect 423 510 427 514
rect 495 510 499 514
rect 575 510 579 514
rect 599 510 603 514
rect 647 510 651 514
rect 703 510 707 514
rect 719 510 723 514
rect 111 450 115 454
rect 319 450 323 454
rect 375 450 379 454
rect 439 450 443 454
rect 455 450 459 454
rect 511 450 515 454
rect 575 450 579 454
rect 1927 690 1931 694
rect 1935 690 1939 694
rect 2015 690 2019 694
rect 2023 690 2027 694
rect 2095 690 2099 694
rect 2119 690 2123 694
rect 2175 690 2179 694
rect 2207 690 2211 694
rect 2263 690 2267 694
rect 1495 634 1499 638
rect 1511 634 1515 638
rect 1599 634 1603 638
rect 1407 624 1411 628
rect 1647 634 1651 638
rect 1703 634 1707 638
rect 1783 634 1787 638
rect 1807 634 1811 638
rect 1911 634 1915 638
rect 2007 634 2011 638
rect 1103 574 1107 578
rect 1183 574 1187 578
rect 1207 574 1211 578
rect 1287 574 1291 578
rect 1327 574 1331 578
rect 1367 570 1371 574
rect 1415 570 1419 574
rect 1471 570 1475 574
rect 1815 624 1819 628
rect 1527 570 1531 574
rect 1551 570 1555 574
rect 1647 570 1651 574
rect 1663 570 1667 574
rect 1751 570 1755 574
rect 1799 570 1803 574
rect 1855 570 1859 574
rect 1927 570 1931 574
rect 2295 690 2299 694
rect 2351 690 2355 694
rect 2391 690 2395 694
rect 2583 690 2587 694
rect 2039 634 2043 638
rect 2103 634 2107 638
rect 2159 634 2163 638
rect 2191 634 2195 638
rect 2279 634 2283 638
rect 2375 634 2379 638
rect 2407 634 2411 638
rect 2583 634 2587 638
rect 1959 570 1963 574
rect 2055 570 2059 574
rect 2151 570 2155 574
rect 2175 570 2179 574
rect 2239 570 2243 574
rect 791 510 795 514
rect 815 510 819 514
rect 863 510 867 514
rect 927 510 931 514
rect 935 510 939 514
rect 1007 510 1011 514
rect 1047 510 1051 514
rect 1087 510 1091 514
rect 1167 510 1171 514
rect 1271 510 1275 514
rect 1327 510 1331 514
rect 1367 514 1371 518
rect 1399 514 1403 518
rect 1455 514 1459 518
rect 1535 514 1539 518
rect 1599 514 1603 518
rect 1631 514 1635 518
rect 1671 514 1675 518
rect 2295 570 2299 574
rect 2319 570 2323 574
rect 2399 570 2403 574
rect 2423 570 2427 574
rect 2479 570 2483 574
rect 2543 570 2547 574
rect 2583 570 2587 574
rect 1735 514 1739 518
rect 1751 514 1755 518
rect 1839 514 1843 518
rect 1927 514 1931 518
rect 1943 514 1947 518
rect 2015 514 2019 518
rect 591 450 595 454
rect 647 450 651 454
rect 663 450 667 454
rect 727 450 731 454
rect 735 450 739 454
rect 799 450 803 454
rect 807 450 811 454
rect 871 450 875 454
rect 879 450 883 454
rect 943 450 947 454
rect 951 450 955 454
rect 1015 450 1019 454
rect 1023 450 1027 454
rect 1087 450 1091 454
rect 1103 450 1107 454
rect 1159 450 1163 454
rect 1239 450 1243 454
rect 1327 450 1331 454
rect 1367 450 1371 454
rect 1551 450 1555 454
rect 1615 450 1619 454
rect 1647 450 1651 454
rect 1687 450 1691 454
rect 1703 450 1707 454
rect 1759 450 1763 454
rect 1767 450 1771 454
rect 111 390 115 394
rect 415 390 419 394
rect 439 390 443 394
rect 471 390 475 394
rect 495 390 499 394
rect 535 390 539 394
rect 559 390 563 394
rect 607 390 611 394
rect 631 390 635 394
rect 687 390 691 394
rect 711 390 715 394
rect 767 390 771 394
rect 783 390 787 394
rect 111 330 115 334
rect 431 330 435 334
rect 847 390 851 394
rect 855 390 859 394
rect 927 390 931 394
rect 999 390 1003 394
rect 1007 390 1011 394
rect 1071 390 1075 394
rect 1087 390 1091 394
rect 1143 390 1147 394
rect 1175 390 1179 394
rect 1223 390 1227 394
rect 463 330 467 334
rect 487 330 491 334
rect 519 330 523 334
rect 551 330 555 334
rect 575 330 579 334
rect 623 330 627 334
rect 631 330 635 334
rect 695 330 699 334
rect 703 330 707 334
rect 767 330 771 334
rect 783 330 787 334
rect 847 330 851 334
rect 111 270 115 274
rect 287 270 291 274
rect 359 270 363 274
rect 439 270 443 274
rect 447 270 451 274
rect 503 270 507 274
rect 863 330 867 334
rect 927 330 931 334
rect 943 330 947 334
rect 527 270 531 274
rect 559 270 563 274
rect 615 270 619 274
rect 623 270 627 274
rect 679 270 683 274
rect 111 214 115 218
rect 199 214 203 218
rect 271 214 275 218
rect 1015 330 1019 334
rect 1023 330 1027 334
rect 2039 514 2043 518
rect 2095 514 2099 518
rect 2135 514 2139 518
rect 2175 514 2179 518
rect 2223 514 2227 518
rect 2255 514 2259 518
rect 2303 514 2307 518
rect 2327 514 2331 518
rect 2383 514 2387 518
rect 2399 514 2403 518
rect 1815 450 1819 454
rect 1855 450 1859 454
rect 1871 450 1875 454
rect 1927 450 1931 454
rect 1943 450 1947 454
rect 1999 450 2003 454
rect 2031 450 2035 454
rect 2087 450 2091 454
rect 2111 450 2115 454
rect 2191 450 2195 454
rect 2463 514 2467 518
rect 2471 514 2475 518
rect 2527 514 2531 518
rect 2583 514 2587 518
rect 2271 450 2275 454
rect 2311 450 2315 454
rect 2343 450 2347 454
rect 2415 450 2419 454
rect 2439 450 2443 454
rect 2487 450 2491 454
rect 2543 450 2547 454
rect 1263 390 1267 394
rect 1327 390 1331 394
rect 1367 394 1371 398
rect 1631 394 1635 398
rect 1655 394 1659 398
rect 1687 394 1691 398
rect 1711 394 1715 398
rect 1743 394 1747 398
rect 1767 394 1771 398
rect 1799 394 1803 398
rect 1823 394 1827 398
rect 1855 394 1859 398
rect 1879 394 1883 398
rect 1911 394 1915 398
rect 2079 416 2083 420
rect 1951 394 1955 398
rect 1983 394 1987 398
rect 2455 416 2459 420
rect 2039 394 2043 398
rect 2071 394 2075 398
rect 2151 394 2155 398
rect 2175 394 2179 398
rect 2279 394 2283 398
rect 2295 394 2299 398
rect 2415 394 2419 398
rect 2423 394 2427 398
rect 2527 394 2531 398
rect 2123 352 2127 356
rect 1103 330 1107 334
rect 1111 330 1115 334
rect 1191 330 1195 334
rect 1215 330 1219 334
rect 1279 330 1283 334
rect 1327 330 1331 334
rect 1367 330 1371 334
rect 1631 330 1635 334
rect 1671 330 1675 334
rect 1687 330 1691 334
rect 1727 330 1731 334
rect 1743 330 1747 334
rect 1783 330 1787 334
rect 1807 330 1811 334
rect 1839 330 1843 334
rect 1887 330 1891 334
rect 1895 330 1899 334
rect 1967 330 1971 334
rect 719 270 723 274
rect 751 270 755 274
rect 823 270 827 274
rect 831 270 835 274
rect 911 270 915 274
rect 927 270 931 274
rect 303 214 307 218
rect 359 214 363 218
rect 375 214 379 218
rect 455 214 459 218
rect 463 214 467 218
rect 543 214 547 218
rect 567 214 571 218
rect 639 214 643 218
rect 679 214 683 218
rect 735 214 739 218
rect 999 270 1003 274
rect 1031 270 1035 274
rect 1095 270 1099 274
rect 1143 270 1147 274
rect 1199 270 1203 274
rect 1255 270 1259 274
rect 1327 270 1331 274
rect 1367 274 1371 278
rect 1535 274 1539 278
rect 1607 274 1611 278
rect 1615 274 1619 278
rect 791 214 795 218
rect 839 214 843 218
rect 911 214 915 218
rect 943 214 947 218
rect 1031 214 1035 218
rect 191 160 195 164
rect 623 160 627 164
rect 111 134 115 138
rect 143 134 147 138
rect 183 134 187 138
rect 199 134 203 138
rect 255 134 259 138
rect 311 134 315 138
rect 343 134 347 138
rect 367 134 371 138
rect 423 134 427 138
rect 447 134 451 138
rect 479 134 483 138
rect 535 134 539 138
rect 551 134 555 138
rect 591 134 595 138
rect 647 134 651 138
rect 663 134 667 138
rect 1047 214 1051 218
rect 1151 214 1155 218
rect 1159 214 1163 218
rect 1271 214 1275 218
rect 2055 330 2059 334
rect 2583 450 2587 454
rect 2583 394 2587 398
rect 2439 352 2443 356
rect 2143 330 2147 334
rect 2167 330 2171 334
rect 2231 330 2235 334
rect 2295 330 2299 334
rect 2311 330 2315 334
rect 2391 330 2395 334
rect 2431 330 2435 334
rect 2479 330 2483 334
rect 2543 330 2547 334
rect 1671 274 1675 278
rect 1687 274 1691 278
rect 1727 274 1731 278
rect 1775 274 1779 278
rect 1791 274 1795 278
rect 1863 274 1867 278
rect 1871 274 1875 278
rect 1951 274 1955 278
rect 2039 274 2043 278
rect 2119 274 2123 278
rect 2127 274 2131 278
rect 2199 274 2203 278
rect 2215 274 2219 278
rect 1327 214 1331 218
rect 1367 218 1371 222
rect 1415 218 1419 222
rect 1479 218 1483 222
rect 1551 218 1555 222
rect 1559 218 1563 222
rect 703 134 707 138
rect 759 134 763 138
rect 775 134 779 138
rect 823 134 827 138
rect 887 134 891 138
rect 895 134 899 138
rect 951 134 955 138
rect 1015 134 1019 138
rect 1079 134 1083 138
rect 111 78 115 82
rect 159 78 163 82
rect 215 78 219 82
rect 271 78 275 82
rect 327 78 331 82
rect 383 78 387 82
rect 439 78 443 82
rect 495 78 499 82
rect 551 78 555 82
rect 607 78 611 82
rect 1135 134 1139 138
rect 1151 134 1155 138
rect 1367 146 1371 150
rect 1399 146 1403 150
rect 1215 134 1219 138
rect 1255 134 1259 138
rect 1271 134 1275 138
rect 1327 134 1331 138
rect 1623 218 1627 222
rect 1655 218 1659 222
rect 1703 218 1707 222
rect 1751 218 1755 222
rect 1791 218 1795 222
rect 1855 218 1859 222
rect 1879 218 1883 222
rect 1959 218 1963 222
rect 1967 218 1971 222
rect 2055 218 2059 222
rect 2063 218 2067 222
rect 2271 274 2275 278
rect 2295 274 2299 278
rect 2335 274 2339 278
rect 2375 274 2379 278
rect 2135 218 2139 222
rect 2407 274 2411 278
rect 2583 330 2587 334
rect 2463 274 2467 278
rect 2471 274 2475 278
rect 2527 274 2531 278
rect 2583 274 2587 278
rect 2167 218 2171 222
rect 1591 184 1595 188
rect 1871 184 1875 188
rect 1455 146 1459 150
rect 1463 146 1467 150
rect 1511 146 1515 150
rect 1543 146 1547 150
rect 1567 146 1571 150
rect 1631 146 1635 150
rect 1639 146 1643 150
rect 1711 146 1715 150
rect 1735 146 1739 150
rect 1791 146 1795 150
rect 1839 146 1843 150
rect 1871 146 1875 150
rect 1407 136 1411 140
rect 663 78 667 82
rect 719 78 723 82
rect 775 78 779 82
rect 839 78 843 82
rect 903 78 907 82
rect 967 78 971 82
rect 1031 78 1035 82
rect 1095 78 1099 82
rect 1823 136 1827 140
rect 2215 218 2219 222
rect 2263 218 2267 222
rect 2287 218 2291 222
rect 2351 218 2355 222
rect 2359 218 2363 222
rect 2423 218 2427 222
rect 2463 218 2467 222
rect 2487 218 2491 222
rect 2543 218 2547 222
rect 1943 146 1947 150
rect 2015 146 2019 150
rect 2047 146 2051 150
rect 2079 146 2083 150
rect 2143 146 2147 150
rect 2151 146 2155 150
rect 2207 146 2211 150
rect 2247 146 2251 150
rect 2271 146 2275 150
rect 1367 90 1371 94
rect 1415 90 1419 94
rect 1471 90 1475 94
rect 1527 90 1531 94
rect 1583 90 1587 94
rect 1647 90 1651 94
rect 1727 90 1731 94
rect 1807 90 1811 94
rect 2583 218 2587 222
rect 2343 146 2347 150
rect 2415 146 2419 150
rect 2447 146 2451 150
rect 2527 146 2531 150
rect 2583 146 2587 150
rect 1887 90 1891 94
rect 1959 90 1963 94
rect 2031 90 2035 94
rect 2095 90 2099 94
rect 2159 90 2163 94
rect 2223 90 2227 94
rect 2287 90 2291 94
rect 2359 90 2363 94
rect 2431 90 2435 94
rect 2583 90 2587 94
rect 1167 78 1171 82
rect 1231 78 1235 82
rect 1287 78 1291 82
rect 1327 78 1331 82
<< m4 >>
rect 84 2637 85 2643
rect 91 2642 1339 2643
rect 91 2638 111 2642
rect 115 2638 551 2642
rect 555 2638 607 2642
rect 611 2638 663 2642
rect 667 2638 719 2642
rect 723 2638 775 2642
rect 779 2638 1327 2642
rect 1331 2638 1339 2642
rect 91 2637 1339 2638
rect 1345 2639 1346 2643
rect 1345 2638 2618 2639
rect 1345 2637 1367 2638
rect 1338 2634 1367 2637
rect 1371 2634 1551 2638
rect 1555 2634 1607 2638
rect 1611 2634 1663 2638
rect 1667 2634 1719 2638
rect 1723 2634 1775 2638
rect 1779 2634 1831 2638
rect 1835 2634 1887 2638
rect 1891 2634 1943 2638
rect 1947 2634 1999 2638
rect 2003 2634 2055 2638
rect 2059 2634 2111 2638
rect 2115 2634 2167 2638
rect 2171 2634 2583 2638
rect 2587 2634 2618 2638
rect 1338 2633 2618 2634
rect 96 2581 97 2587
rect 103 2586 1351 2587
rect 103 2582 111 2586
rect 115 2582 215 2586
rect 219 2582 271 2586
rect 275 2582 327 2586
rect 331 2582 383 2586
rect 387 2582 439 2586
rect 443 2582 495 2586
rect 499 2582 535 2586
rect 539 2582 551 2586
rect 555 2582 591 2586
rect 595 2582 607 2586
rect 611 2582 647 2586
rect 651 2582 663 2586
rect 667 2582 703 2586
rect 707 2582 719 2586
rect 723 2582 759 2586
rect 763 2582 775 2586
rect 779 2582 831 2586
rect 835 2582 887 2586
rect 891 2582 943 2586
rect 947 2582 999 2586
rect 1003 2582 1055 2586
rect 1059 2582 1111 2586
rect 1115 2582 1327 2586
rect 1331 2582 1351 2586
rect 103 2581 1351 2582
rect 1357 2583 1358 2587
rect 1357 2582 2630 2583
rect 1357 2581 1367 2582
rect 1350 2578 1367 2581
rect 1371 2578 1439 2582
rect 1443 2578 1535 2582
rect 1539 2578 1543 2582
rect 1547 2578 1591 2582
rect 1595 2578 1647 2582
rect 1651 2578 1655 2582
rect 1659 2578 1703 2582
rect 1707 2578 1759 2582
rect 1763 2578 1767 2582
rect 1771 2578 1815 2582
rect 1819 2578 1871 2582
rect 1875 2578 1879 2582
rect 1883 2578 1927 2582
rect 1931 2578 1983 2582
rect 1987 2578 1991 2582
rect 1995 2578 2039 2582
rect 2043 2578 2095 2582
rect 2099 2578 2111 2582
rect 2115 2578 2151 2582
rect 2155 2578 2231 2582
rect 2235 2578 2351 2582
rect 2355 2578 2583 2582
rect 2587 2578 2630 2582
rect 1350 2577 2630 2578
rect 1542 2532 1548 2533
rect 1902 2532 1908 2533
rect 1542 2528 1543 2532
rect 1547 2528 1903 2532
rect 1907 2528 1908 2532
rect 1542 2527 1548 2528
rect 1902 2527 1908 2528
rect 84 2521 85 2527
rect 91 2526 1339 2527
rect 91 2522 111 2526
rect 115 2522 231 2526
rect 235 2522 287 2526
rect 291 2522 343 2526
rect 347 2522 367 2526
rect 371 2522 399 2526
rect 403 2522 423 2526
rect 427 2522 455 2526
rect 459 2522 487 2526
rect 491 2522 511 2526
rect 515 2522 551 2526
rect 555 2522 567 2526
rect 571 2522 615 2526
rect 619 2522 623 2526
rect 627 2522 679 2526
rect 683 2522 735 2526
rect 739 2522 743 2526
rect 747 2522 791 2526
rect 795 2522 807 2526
rect 811 2522 847 2526
rect 851 2522 871 2526
rect 875 2522 903 2526
rect 907 2522 943 2526
rect 947 2522 959 2526
rect 963 2522 1015 2526
rect 1019 2522 1071 2526
rect 1075 2522 1127 2526
rect 1131 2522 1327 2526
rect 1331 2522 1339 2526
rect 91 2521 1339 2522
rect 1345 2521 1346 2527
rect 1338 2519 1346 2521
rect 1338 2513 1339 2519
rect 1345 2518 2611 2519
rect 1345 2514 1367 2518
rect 1371 2514 1455 2518
rect 1459 2514 1551 2518
rect 1555 2514 1559 2518
rect 1563 2514 1631 2518
rect 1635 2514 1671 2518
rect 1675 2514 1719 2518
rect 1723 2514 1783 2518
rect 1787 2514 1807 2518
rect 1811 2514 1895 2518
rect 1899 2514 1903 2518
rect 1907 2514 1999 2518
rect 2003 2514 2007 2518
rect 2011 2514 2095 2518
rect 2099 2514 2127 2518
rect 2131 2514 2191 2518
rect 2195 2514 2247 2518
rect 2251 2514 2295 2518
rect 2299 2514 2367 2518
rect 2371 2514 2399 2518
rect 2403 2514 2583 2518
rect 2587 2514 2611 2518
rect 1345 2513 2611 2514
rect 2617 2513 2618 2519
rect 96 2461 97 2467
rect 103 2466 1351 2467
rect 103 2462 111 2466
rect 115 2462 271 2466
rect 275 2462 335 2466
rect 339 2462 351 2466
rect 355 2462 399 2466
rect 403 2462 407 2466
rect 411 2462 471 2466
rect 475 2462 535 2466
rect 539 2462 551 2466
rect 555 2462 599 2466
rect 603 2462 631 2466
rect 635 2462 663 2466
rect 667 2462 711 2466
rect 715 2462 727 2466
rect 731 2462 783 2466
rect 787 2462 791 2466
rect 795 2462 855 2466
rect 859 2462 863 2466
rect 867 2462 927 2466
rect 931 2462 943 2466
rect 947 2462 999 2466
rect 1003 2462 1023 2466
rect 1027 2462 1327 2466
rect 1331 2462 1351 2466
rect 103 2461 1351 2462
rect 1357 2463 1358 2467
rect 1357 2462 2630 2463
rect 1357 2461 1367 2462
rect 1350 2458 1367 2461
rect 1371 2458 1535 2462
rect 1539 2458 1615 2462
rect 1619 2458 1647 2462
rect 1651 2458 1703 2462
rect 1707 2458 1767 2462
rect 1771 2458 1791 2462
rect 1795 2458 1839 2462
rect 1843 2458 1887 2462
rect 1891 2458 1911 2462
rect 1915 2458 1983 2462
rect 1987 2458 1991 2462
rect 1995 2458 2079 2462
rect 2083 2458 2167 2462
rect 2171 2458 2175 2462
rect 2179 2458 2263 2462
rect 2267 2458 2279 2462
rect 2283 2458 2359 2462
rect 2363 2458 2383 2462
rect 2387 2458 2455 2462
rect 2459 2458 2527 2462
rect 2531 2458 2583 2462
rect 2587 2458 2630 2462
rect 1350 2457 2630 2458
rect 84 2401 85 2407
rect 91 2406 1339 2407
rect 91 2402 111 2406
rect 115 2402 247 2406
rect 251 2402 287 2406
rect 291 2402 335 2406
rect 339 2402 351 2406
rect 355 2402 415 2406
rect 419 2402 431 2406
rect 435 2402 487 2406
rect 491 2402 527 2406
rect 531 2402 567 2406
rect 571 2402 631 2406
rect 635 2402 647 2406
rect 651 2402 727 2406
rect 731 2402 799 2406
rect 803 2402 823 2406
rect 827 2402 879 2406
rect 883 2402 919 2406
rect 923 2402 959 2406
rect 963 2402 1015 2406
rect 1019 2402 1039 2406
rect 1043 2402 1111 2406
rect 1115 2402 1327 2406
rect 1331 2402 1339 2406
rect 91 2401 1339 2402
rect 1345 2403 1346 2407
rect 1345 2402 2618 2403
rect 1345 2401 1367 2402
rect 1338 2398 1367 2401
rect 1371 2398 1455 2402
rect 1459 2398 1559 2402
rect 1563 2398 1663 2402
rect 1667 2398 1719 2402
rect 1723 2398 1759 2402
rect 1763 2398 1783 2402
rect 1787 2398 1855 2402
rect 1859 2398 1927 2402
rect 1931 2398 1943 2402
rect 1947 2398 2007 2402
rect 2011 2398 2039 2402
rect 2043 2398 2095 2402
rect 2099 2398 2135 2402
rect 2139 2398 2183 2402
rect 2187 2398 2231 2402
rect 2235 2398 2279 2402
rect 2283 2398 2335 2402
rect 2339 2398 2375 2402
rect 2379 2398 2447 2402
rect 2451 2398 2471 2402
rect 2475 2398 2543 2402
rect 2547 2398 2583 2402
rect 2587 2398 2618 2402
rect 1338 2397 2618 2398
rect 238 2372 244 2373
rect 646 2372 652 2373
rect 238 2368 239 2372
rect 243 2368 647 2372
rect 651 2368 652 2372
rect 238 2367 244 2368
rect 646 2367 652 2368
rect 96 2345 97 2351
rect 103 2350 1351 2351
rect 103 2346 111 2350
rect 115 2346 159 2350
rect 163 2346 231 2350
rect 235 2346 263 2350
rect 267 2346 319 2350
rect 323 2346 375 2350
rect 379 2346 415 2350
rect 419 2346 487 2350
rect 491 2346 511 2350
rect 515 2346 599 2350
rect 603 2346 615 2350
rect 619 2346 711 2350
rect 715 2346 807 2350
rect 811 2346 815 2350
rect 819 2346 903 2350
rect 907 2346 911 2350
rect 915 2346 999 2350
rect 1003 2346 1007 2350
rect 1011 2346 1095 2350
rect 1099 2346 1103 2350
rect 1107 2346 1199 2350
rect 1203 2346 1327 2350
rect 1331 2346 1351 2350
rect 103 2345 1351 2346
rect 1357 2347 1358 2351
rect 1357 2346 2630 2347
rect 1357 2345 1367 2346
rect 1350 2342 1367 2345
rect 1371 2342 1399 2346
rect 1403 2342 1439 2346
rect 1443 2342 1455 2346
rect 1459 2342 1511 2346
rect 1515 2342 1543 2346
rect 1547 2342 1567 2346
rect 1571 2342 1639 2346
rect 1643 2342 1647 2346
rect 1651 2342 1727 2346
rect 1731 2342 1743 2346
rect 1747 2342 1823 2346
rect 1827 2342 1839 2346
rect 1843 2342 1927 2346
rect 1931 2342 1943 2346
rect 1947 2342 2023 2346
rect 2027 2342 2079 2346
rect 2083 2342 2119 2346
rect 2123 2342 2215 2346
rect 2219 2342 2223 2346
rect 2227 2342 2319 2346
rect 2323 2342 2383 2346
rect 2387 2342 2431 2346
rect 2435 2342 2527 2346
rect 2531 2342 2583 2346
rect 2587 2342 2630 2346
rect 1350 2341 2630 2342
rect 84 2285 85 2291
rect 91 2290 1339 2291
rect 91 2286 111 2290
rect 115 2286 159 2290
rect 163 2286 175 2290
rect 179 2286 247 2290
rect 251 2286 279 2290
rect 283 2286 375 2290
rect 379 2286 391 2290
rect 395 2286 503 2290
rect 507 2286 511 2290
rect 515 2286 615 2290
rect 619 2286 639 2290
rect 643 2286 727 2290
rect 731 2286 767 2290
rect 771 2286 831 2290
rect 835 2286 887 2290
rect 891 2286 927 2290
rect 931 2286 999 2290
rect 1003 2286 1023 2290
rect 1027 2286 1103 2290
rect 1107 2286 1119 2290
rect 1123 2286 1207 2290
rect 1211 2286 1215 2290
rect 1219 2286 1287 2290
rect 1291 2286 1327 2290
rect 1331 2286 1339 2290
rect 91 2285 1339 2286
rect 1345 2285 1346 2291
rect 1338 2283 1346 2285
rect 1338 2277 1339 2283
rect 1345 2282 2611 2283
rect 1345 2278 1367 2282
rect 1371 2278 1415 2282
rect 1419 2278 1471 2282
rect 1475 2278 1495 2282
rect 1499 2278 1527 2282
rect 1531 2278 1583 2282
rect 1587 2278 1615 2282
rect 1619 2278 1655 2282
rect 1659 2278 1735 2282
rect 1739 2278 1743 2282
rect 1747 2278 1839 2282
rect 1843 2278 1855 2282
rect 1859 2278 1959 2282
rect 1963 2278 1967 2282
rect 1971 2278 2071 2282
rect 2075 2278 2095 2282
rect 2099 2278 2167 2282
rect 2171 2278 2239 2282
rect 2243 2278 2255 2282
rect 2259 2278 2335 2282
rect 2339 2278 2399 2282
rect 2403 2278 2407 2282
rect 2411 2278 2487 2282
rect 2491 2278 2543 2282
rect 2547 2278 2583 2282
rect 2587 2278 2611 2282
rect 1345 2277 2611 2278
rect 2617 2277 2618 2283
rect 96 2221 97 2227
rect 103 2226 1351 2227
rect 103 2222 111 2226
rect 115 2222 143 2226
rect 147 2222 231 2226
rect 235 2222 359 2226
rect 363 2222 495 2226
rect 499 2222 623 2226
rect 627 2222 751 2226
rect 755 2222 871 2226
rect 875 2222 983 2226
rect 987 2222 1087 2226
rect 1091 2222 1191 2226
rect 1195 2222 1271 2226
rect 1275 2222 1327 2226
rect 1331 2222 1351 2226
rect 103 2221 1351 2222
rect 1357 2221 1358 2227
rect 1350 2209 1351 2215
rect 1357 2214 2623 2215
rect 1357 2210 1367 2214
rect 1371 2210 1399 2214
rect 1403 2210 1455 2214
rect 1459 2210 1479 2214
rect 1483 2210 1535 2214
rect 1539 2210 1599 2214
rect 1603 2210 1631 2214
rect 1635 2210 1719 2214
rect 1723 2210 1743 2214
rect 1747 2210 1839 2214
rect 1843 2210 1863 2214
rect 1867 2210 1951 2214
rect 1955 2210 1983 2214
rect 1987 2210 2055 2214
rect 2059 2210 2095 2214
rect 2099 2210 2151 2214
rect 2155 2210 2207 2214
rect 2211 2210 2239 2214
rect 2243 2210 2311 2214
rect 2315 2210 2319 2214
rect 2323 2210 2391 2214
rect 2395 2210 2423 2214
rect 2427 2210 2471 2214
rect 2475 2210 2527 2214
rect 2531 2210 2583 2214
rect 2587 2210 2623 2214
rect 1357 2209 2623 2210
rect 2629 2209 2630 2215
rect 138 2188 144 2189
rect 646 2188 652 2189
rect 138 2184 139 2188
rect 143 2184 647 2188
rect 651 2184 652 2188
rect 138 2183 144 2184
rect 646 2183 652 2184
rect 84 2161 85 2167
rect 91 2166 1339 2167
rect 91 2162 111 2166
rect 115 2162 159 2166
rect 163 2162 215 2166
rect 219 2162 247 2166
rect 251 2162 311 2166
rect 315 2162 375 2166
rect 379 2162 423 2166
rect 427 2162 511 2166
rect 515 2162 543 2166
rect 547 2162 639 2166
rect 643 2162 663 2166
rect 667 2162 767 2166
rect 771 2162 775 2166
rect 779 2162 879 2166
rect 883 2162 887 2166
rect 891 2162 975 2166
rect 979 2162 999 2166
rect 1003 2162 1071 2166
rect 1075 2162 1103 2166
rect 1107 2162 1167 2166
rect 1171 2162 1207 2166
rect 1211 2162 1271 2166
rect 1275 2162 1287 2166
rect 1291 2162 1327 2166
rect 1331 2162 1339 2166
rect 91 2161 1339 2162
rect 1345 2161 1346 2167
rect 1338 2159 1346 2161
rect 1338 2153 1339 2159
rect 1345 2158 2611 2159
rect 1345 2154 1367 2158
rect 1371 2154 1471 2158
rect 1475 2154 1535 2158
rect 1539 2154 1551 2158
rect 1555 2154 1631 2158
rect 1635 2154 1647 2158
rect 1651 2154 1735 2158
rect 1739 2154 1759 2158
rect 1763 2154 1839 2158
rect 1843 2154 1879 2158
rect 1883 2154 1951 2158
rect 1955 2154 1999 2158
rect 2003 2154 2055 2158
rect 2059 2154 2111 2158
rect 2115 2154 2159 2158
rect 2163 2154 2223 2158
rect 2227 2154 2263 2158
rect 2267 2154 2327 2158
rect 2331 2154 2359 2158
rect 2363 2154 2439 2158
rect 2443 2154 2463 2158
rect 2467 2154 2543 2158
rect 2547 2154 2583 2158
rect 2587 2154 2611 2158
rect 1345 2153 2611 2154
rect 2617 2153 2618 2159
rect 854 2132 860 2133
rect 1286 2132 1292 2133
rect 854 2128 855 2132
rect 859 2128 1287 2132
rect 1291 2128 1292 2132
rect 854 2127 860 2128
rect 1286 2127 1292 2128
rect 96 2097 97 2103
rect 103 2102 1351 2103
rect 103 2098 111 2102
rect 115 2098 143 2102
rect 147 2098 199 2102
rect 203 2098 263 2102
rect 267 2098 295 2102
rect 299 2098 327 2102
rect 331 2098 399 2102
rect 403 2098 407 2102
rect 411 2098 479 2102
rect 483 2098 527 2102
rect 531 2098 567 2102
rect 571 2098 647 2102
rect 651 2098 655 2102
rect 659 2098 735 2102
rect 739 2098 759 2102
rect 763 2098 815 2102
rect 819 2098 863 2102
rect 867 2098 887 2102
rect 891 2098 959 2102
rect 963 2098 967 2102
rect 971 2098 1047 2102
rect 1051 2098 1055 2102
rect 1059 2098 1127 2102
rect 1131 2098 1151 2102
rect 1155 2098 1255 2102
rect 1259 2098 1327 2102
rect 1331 2098 1351 2102
rect 103 2097 1351 2098
rect 1357 2102 2630 2103
rect 1357 2098 1367 2102
rect 1371 2098 1431 2102
rect 1435 2098 1519 2102
rect 1523 2098 1535 2102
rect 1539 2098 1615 2102
rect 1619 2098 1647 2102
rect 1651 2098 1719 2102
rect 1723 2098 1759 2102
rect 1763 2098 1823 2102
rect 1827 2098 1863 2102
rect 1867 2098 1935 2102
rect 1939 2098 1967 2102
rect 1971 2098 2039 2102
rect 2043 2098 2071 2102
rect 2075 2098 2143 2102
rect 2147 2098 2175 2102
rect 2179 2098 2247 2102
rect 2251 2098 2271 2102
rect 2275 2098 2343 2102
rect 2347 2098 2359 2102
rect 2363 2098 2447 2102
rect 2451 2098 2455 2102
rect 2459 2098 2527 2102
rect 2531 2098 2583 2102
rect 2587 2098 2630 2102
rect 1357 2097 2630 2098
rect 258 2076 264 2077
rect 670 2076 676 2077
rect 258 2072 259 2076
rect 263 2072 671 2076
rect 675 2072 676 2076
rect 258 2071 264 2072
rect 670 2071 676 2072
rect 1338 2041 1339 2047
rect 1345 2046 2611 2047
rect 1345 2042 1367 2046
rect 1371 2042 1415 2046
rect 1419 2042 1447 2046
rect 1451 2042 1503 2046
rect 1507 2042 1551 2046
rect 1555 2042 1607 2046
rect 1611 2042 1663 2046
rect 1667 2042 1711 2046
rect 1715 2042 1775 2046
rect 1779 2042 1807 2046
rect 1811 2042 1879 2046
rect 1883 2042 1903 2046
rect 1907 2042 1983 2046
rect 1987 2042 2007 2046
rect 2011 2042 2087 2046
rect 2091 2042 2111 2046
rect 2115 2042 2191 2046
rect 2195 2042 2215 2046
rect 2219 2042 2287 2046
rect 2291 2042 2327 2046
rect 2331 2042 2375 2046
rect 2379 2042 2447 2046
rect 2451 2042 2471 2046
rect 2475 2042 2543 2046
rect 2547 2042 2583 2046
rect 2587 2042 2611 2046
rect 1345 2041 2611 2042
rect 2617 2041 2618 2047
rect 1338 2039 1346 2041
rect 84 2033 85 2039
rect 91 2038 1339 2039
rect 91 2034 111 2038
rect 115 2034 279 2038
rect 283 2034 343 2038
rect 347 2034 415 2038
rect 419 2034 471 2038
rect 475 2034 495 2038
rect 499 2034 527 2038
rect 531 2034 583 2038
rect 587 2034 639 2038
rect 643 2034 671 2038
rect 675 2034 695 2038
rect 699 2034 751 2038
rect 755 2034 807 2038
rect 811 2034 831 2038
rect 835 2034 863 2038
rect 867 2034 903 2038
rect 907 2034 919 2038
rect 923 2034 975 2038
rect 979 2034 983 2038
rect 987 2034 1031 2038
rect 1035 2034 1063 2038
rect 1067 2034 1143 2038
rect 1147 2034 1327 2038
rect 1331 2034 1339 2038
rect 91 2033 1339 2034
rect 1345 2033 1346 2039
rect 742 1996 748 1997
rect 1174 1996 1180 1997
rect 742 1992 743 1996
rect 747 1992 1175 1996
rect 1179 1992 1180 1996
rect 742 1991 748 1992
rect 1174 1991 1180 1992
rect 1350 1985 1351 1991
rect 1357 1990 2623 1991
rect 1357 1986 1367 1990
rect 1371 1986 1399 1990
rect 1403 1986 1479 1990
rect 1483 1986 1487 1990
rect 1491 1986 1583 1990
rect 1587 1986 1591 1990
rect 1595 1986 1679 1990
rect 1683 1986 1695 1990
rect 1699 1986 1767 1990
rect 1771 1986 1791 1990
rect 1795 1986 1847 1990
rect 1851 1986 1887 1990
rect 1891 1986 1927 1990
rect 1931 1986 1991 1990
rect 1995 1986 2007 1990
rect 2011 1986 2087 1990
rect 2091 1986 2095 1990
rect 2099 1986 2199 1990
rect 2203 1986 2311 1990
rect 2315 1986 2431 1990
rect 2435 1986 2527 1990
rect 2531 1986 2583 1990
rect 2587 1986 2623 1990
rect 1357 1985 2623 1986
rect 2629 1985 2630 1991
rect 96 1973 97 1979
rect 103 1978 1351 1979
rect 103 1974 111 1978
rect 115 1974 335 1978
rect 339 1974 391 1978
rect 395 1974 399 1978
rect 403 1974 447 1978
rect 451 1974 455 1978
rect 459 1974 503 1978
rect 507 1974 511 1978
rect 515 1974 567 1978
rect 571 1974 623 1978
rect 627 1974 647 1978
rect 651 1974 679 1978
rect 683 1974 735 1978
rect 739 1974 743 1978
rect 747 1974 791 1978
rect 795 1974 847 1978
rect 851 1974 863 1978
rect 867 1974 903 1978
rect 907 1974 959 1978
rect 963 1974 999 1978
rect 1003 1974 1015 1978
rect 1019 1974 1143 1978
rect 1147 1974 1271 1978
rect 1275 1974 1327 1978
rect 1331 1974 1351 1978
rect 103 1973 1351 1974
rect 1357 1973 1358 1979
rect 1338 1925 1339 1931
rect 1345 1930 2611 1931
rect 1345 1926 1367 1930
rect 1371 1926 1415 1930
rect 1419 1926 1495 1930
rect 1499 1926 1599 1930
rect 1603 1926 1695 1930
rect 1699 1926 1719 1930
rect 1723 1926 1775 1930
rect 1779 1926 1783 1930
rect 1787 1926 1831 1930
rect 1835 1926 1863 1930
rect 1867 1926 1887 1930
rect 1891 1926 1943 1930
rect 1947 1926 1999 1930
rect 2003 1926 2023 1930
rect 2027 1926 2055 1930
rect 2059 1926 2103 1930
rect 2107 1926 2119 1930
rect 2123 1926 2583 1930
rect 2587 1926 2611 1930
rect 1345 1925 2611 1926
rect 2617 1925 2618 1931
rect 1338 1923 1346 1925
rect 84 1917 85 1923
rect 91 1922 1339 1923
rect 91 1918 111 1922
rect 115 1918 159 1922
rect 163 1918 231 1922
rect 235 1918 327 1922
rect 331 1918 351 1922
rect 355 1918 407 1922
rect 411 1918 431 1922
rect 435 1918 463 1922
rect 467 1918 519 1922
rect 523 1918 543 1922
rect 547 1918 583 1922
rect 587 1918 655 1922
rect 659 1918 663 1922
rect 667 1918 759 1922
rect 763 1918 767 1922
rect 771 1918 879 1922
rect 883 1918 983 1922
rect 987 1918 1015 1922
rect 1019 1918 1087 1922
rect 1091 1918 1159 1922
rect 1163 1918 1199 1922
rect 1203 1918 1287 1922
rect 1291 1918 1327 1922
rect 1331 1918 1339 1922
rect 91 1917 1339 1918
rect 1345 1917 1346 1923
rect 1350 1865 1351 1871
rect 1357 1870 2623 1871
rect 1357 1866 1367 1870
rect 1371 1866 1399 1870
rect 1403 1866 1463 1870
rect 1467 1866 1559 1870
rect 1563 1866 1655 1870
rect 1659 1866 1703 1870
rect 1707 1866 1743 1870
rect 1747 1866 1759 1870
rect 1763 1866 1815 1870
rect 1819 1866 1831 1870
rect 1835 1866 1871 1870
rect 1875 1866 1919 1870
rect 1923 1866 1927 1870
rect 1931 1866 1983 1870
rect 1987 1866 2007 1870
rect 2011 1866 2039 1870
rect 2043 1866 2095 1870
rect 2099 1866 2103 1870
rect 2107 1866 2183 1870
rect 2187 1866 2583 1870
rect 2587 1866 2623 1870
rect 1357 1865 2623 1866
rect 2629 1865 2630 1871
rect 96 1853 97 1859
rect 103 1858 1351 1859
rect 103 1854 111 1858
rect 115 1854 143 1858
rect 147 1854 199 1858
rect 203 1854 215 1858
rect 219 1854 263 1858
rect 267 1854 311 1858
rect 315 1854 351 1858
rect 355 1854 415 1858
rect 419 1854 439 1858
rect 443 1854 527 1858
rect 531 1854 535 1858
rect 539 1854 623 1858
rect 627 1854 639 1858
rect 643 1854 711 1858
rect 715 1854 751 1858
rect 755 1854 791 1858
rect 795 1854 863 1858
rect 867 1854 871 1858
rect 875 1854 951 1858
rect 955 1854 967 1858
rect 971 1854 1039 1858
rect 1043 1854 1071 1858
rect 1075 1854 1183 1858
rect 1187 1854 1271 1858
rect 1275 1854 1327 1858
rect 1331 1854 1351 1858
rect 103 1853 1351 1854
rect 1357 1853 1358 1859
rect 1826 1828 1832 1829
rect 2206 1828 2212 1829
rect 1826 1824 1827 1828
rect 1831 1824 2207 1828
rect 2211 1824 2212 1828
rect 1826 1823 1832 1824
rect 2206 1823 2212 1824
rect 1338 1809 1339 1815
rect 1345 1814 2611 1815
rect 1345 1810 1367 1814
rect 1371 1810 1415 1814
rect 1419 1810 1479 1814
rect 1483 1810 1511 1814
rect 1515 1810 1575 1814
rect 1579 1810 1623 1814
rect 1627 1810 1671 1814
rect 1675 1810 1735 1814
rect 1739 1810 1759 1814
rect 1763 1810 1839 1814
rect 1843 1810 1847 1814
rect 1851 1810 1935 1814
rect 1939 1810 1951 1814
rect 1955 1810 2023 1814
rect 2027 1810 2063 1814
rect 2067 1810 2111 1814
rect 2115 1810 2183 1814
rect 2187 1810 2199 1814
rect 2203 1810 2303 1814
rect 2307 1810 2431 1814
rect 2435 1810 2543 1814
rect 2547 1810 2583 1814
rect 2587 1810 2611 1814
rect 1345 1809 2611 1810
rect 2617 1809 2618 1815
rect 84 1793 85 1799
rect 91 1798 1339 1799
rect 91 1794 111 1798
rect 115 1794 159 1798
rect 163 1794 215 1798
rect 219 1794 231 1798
rect 235 1794 279 1798
rect 283 1794 295 1798
rect 299 1794 367 1798
rect 371 1794 447 1798
rect 451 1794 455 1798
rect 459 1794 535 1798
rect 539 1794 551 1798
rect 555 1794 623 1798
rect 627 1794 639 1798
rect 643 1794 711 1798
rect 715 1794 727 1798
rect 731 1794 791 1798
rect 795 1794 807 1798
rect 811 1794 871 1798
rect 875 1794 887 1798
rect 891 1794 951 1798
rect 955 1794 967 1798
rect 971 1794 1031 1798
rect 1035 1794 1055 1798
rect 1059 1794 1119 1798
rect 1123 1794 1327 1798
rect 1331 1794 1339 1798
rect 91 1793 1339 1794
rect 1345 1793 1346 1799
rect 1350 1753 1351 1759
rect 1357 1758 2623 1759
rect 1357 1754 1367 1758
rect 1371 1754 1399 1758
rect 1403 1754 1439 1758
rect 1443 1754 1495 1758
rect 1499 1754 1519 1758
rect 1523 1754 1607 1758
rect 1611 1754 1615 1758
rect 1619 1754 1719 1758
rect 1723 1754 1823 1758
rect 1827 1754 1927 1758
rect 1931 1754 1935 1758
rect 1939 1754 2023 1758
rect 2027 1754 2047 1758
rect 2051 1754 2119 1758
rect 2123 1754 2167 1758
rect 2171 1754 2207 1758
rect 2211 1754 2287 1758
rect 2291 1754 2375 1758
rect 2379 1754 2415 1758
rect 2419 1754 2463 1758
rect 2467 1754 2527 1758
rect 2531 1754 2583 1758
rect 2587 1754 2623 1758
rect 1357 1753 2623 1754
rect 2629 1753 2630 1759
rect 96 1733 97 1739
rect 103 1738 1351 1739
rect 103 1734 111 1738
rect 115 1734 215 1738
rect 219 1734 279 1738
rect 283 1734 351 1738
rect 355 1734 407 1738
rect 411 1734 431 1738
rect 435 1734 471 1738
rect 475 1734 519 1738
rect 523 1734 551 1738
rect 555 1734 607 1738
rect 611 1734 639 1738
rect 643 1734 695 1738
rect 699 1734 727 1738
rect 731 1734 775 1738
rect 779 1734 823 1738
rect 827 1734 855 1738
rect 859 1734 919 1738
rect 923 1734 935 1738
rect 939 1734 1015 1738
rect 1019 1734 1103 1738
rect 1107 1734 1111 1738
rect 1115 1734 1207 1738
rect 1211 1734 1327 1738
rect 1331 1734 1351 1738
rect 103 1733 1351 1734
rect 1357 1733 1358 1739
rect 2018 1716 2024 1717
rect 2398 1716 2404 1717
rect 2018 1712 2019 1716
rect 2023 1712 2399 1716
rect 2403 1712 2404 1716
rect 2018 1711 2024 1712
rect 2398 1711 2404 1712
rect 1338 1685 1339 1691
rect 1345 1690 2611 1691
rect 1345 1686 1367 1690
rect 1371 1686 1455 1690
rect 1459 1686 1535 1690
rect 1539 1686 1559 1690
rect 1563 1686 1631 1690
rect 1635 1686 1711 1690
rect 1715 1686 1735 1690
rect 1739 1686 1799 1690
rect 1803 1686 1839 1690
rect 1843 1686 1887 1690
rect 1891 1686 1943 1690
rect 1947 1686 1975 1690
rect 1979 1686 2039 1690
rect 2043 1686 2063 1690
rect 2067 1686 2135 1690
rect 2139 1686 2143 1690
rect 2147 1686 2215 1690
rect 2219 1686 2223 1690
rect 2227 1686 2287 1690
rect 2291 1686 2303 1690
rect 2307 1686 2351 1690
rect 2355 1686 2391 1690
rect 2395 1686 2423 1690
rect 2427 1686 2479 1690
rect 2483 1686 2487 1690
rect 2491 1686 2543 1690
rect 2547 1686 2583 1690
rect 2587 1686 2611 1690
rect 1345 1685 2611 1686
rect 2617 1685 2618 1691
rect 84 1673 85 1679
rect 91 1678 1339 1679
rect 91 1674 111 1678
rect 115 1674 367 1678
rect 371 1674 399 1678
rect 403 1674 423 1678
rect 427 1674 455 1678
rect 459 1674 487 1678
rect 491 1674 511 1678
rect 515 1674 567 1678
rect 571 1674 575 1678
rect 579 1674 647 1678
rect 651 1674 655 1678
rect 659 1674 727 1678
rect 731 1674 743 1678
rect 747 1674 807 1678
rect 811 1674 839 1678
rect 843 1674 887 1678
rect 891 1674 935 1678
rect 939 1674 967 1678
rect 971 1674 1031 1678
rect 1035 1674 1047 1678
rect 1051 1674 1127 1678
rect 1131 1674 1135 1678
rect 1139 1674 1223 1678
rect 1227 1674 1287 1678
rect 1291 1674 1327 1678
rect 1331 1674 1339 1678
rect 91 1673 1339 1674
rect 1345 1673 1346 1679
rect 1350 1617 1351 1623
rect 1357 1622 2623 1623
rect 1357 1618 1367 1622
rect 1371 1618 1543 1622
rect 1547 1618 1575 1622
rect 1579 1618 1615 1622
rect 1619 1618 1631 1622
rect 1635 1618 1687 1622
rect 1691 1618 1695 1622
rect 1699 1618 1751 1622
rect 1755 1618 1783 1622
rect 1787 1618 1831 1622
rect 1835 1618 1871 1622
rect 1875 1618 1919 1622
rect 1923 1618 1959 1622
rect 1963 1618 2007 1622
rect 2011 1618 2047 1622
rect 2051 1618 2103 1622
rect 2107 1618 2127 1622
rect 2131 1618 2199 1622
rect 2203 1618 2207 1622
rect 2211 1618 2271 1622
rect 2275 1618 2319 1622
rect 2323 1618 2335 1622
rect 2339 1618 2407 1622
rect 2411 1618 2431 1622
rect 2435 1618 2471 1622
rect 2475 1618 2527 1622
rect 2531 1618 2583 1622
rect 2587 1618 2623 1622
rect 1357 1617 2623 1618
rect 2629 1617 2630 1623
rect 96 1601 97 1607
rect 103 1606 1351 1607
rect 103 1602 111 1606
rect 115 1602 287 1606
rect 291 1602 367 1606
rect 371 1602 383 1606
rect 387 1602 439 1606
rect 443 1602 455 1606
rect 459 1602 495 1606
rect 499 1602 551 1606
rect 555 1602 559 1606
rect 563 1602 631 1606
rect 635 1602 647 1606
rect 651 1602 711 1606
rect 715 1602 735 1606
rect 739 1602 791 1606
rect 795 1602 823 1606
rect 827 1602 871 1606
rect 875 1602 903 1606
rect 907 1602 951 1606
rect 955 1602 983 1606
rect 987 1602 1031 1606
rect 1035 1602 1063 1606
rect 1067 1602 1119 1606
rect 1123 1602 1151 1606
rect 1155 1602 1207 1606
rect 1211 1602 1271 1606
rect 1275 1602 1327 1606
rect 1331 1602 1351 1606
rect 103 1601 1351 1602
rect 1357 1601 1358 1607
rect 1338 1557 1339 1563
rect 1345 1562 2611 1563
rect 1345 1558 1367 1562
rect 1371 1558 1591 1562
rect 1595 1558 1647 1562
rect 1651 1558 1679 1562
rect 1683 1558 1703 1562
rect 1707 1558 1735 1562
rect 1739 1558 1767 1562
rect 1771 1558 1791 1562
rect 1795 1558 1847 1562
rect 1851 1558 1855 1562
rect 1859 1558 1927 1562
rect 1931 1558 1935 1562
rect 1939 1558 2007 1562
rect 2011 1558 2023 1562
rect 2027 1558 2087 1562
rect 2091 1558 2119 1562
rect 2123 1558 2167 1562
rect 2171 1558 2223 1562
rect 2227 1558 2247 1562
rect 2251 1558 2327 1562
rect 2331 1558 2335 1562
rect 2339 1558 2407 1562
rect 2411 1558 2447 1562
rect 2451 1558 2487 1562
rect 2491 1558 2543 1562
rect 2547 1558 2583 1562
rect 2587 1558 2611 1562
rect 1345 1557 2611 1558
rect 2617 1557 2618 1563
rect 84 1545 85 1551
rect 91 1550 1339 1551
rect 91 1546 111 1550
rect 115 1546 279 1550
rect 283 1546 303 1550
rect 307 1546 335 1550
rect 339 1546 383 1550
rect 387 1546 399 1550
rect 403 1546 471 1550
rect 475 1546 543 1550
rect 547 1546 567 1550
rect 571 1546 615 1550
rect 619 1546 663 1550
rect 667 1546 687 1550
rect 691 1546 751 1550
rect 755 1546 759 1550
rect 763 1546 831 1550
rect 835 1546 839 1550
rect 843 1546 903 1550
rect 907 1546 919 1550
rect 923 1546 975 1550
rect 979 1546 999 1550
rect 1003 1546 1055 1550
rect 1059 1546 1079 1550
rect 1083 1546 1167 1550
rect 1171 1546 1327 1550
rect 1331 1546 1339 1550
rect 91 1545 1339 1546
rect 1345 1545 1346 1551
rect 1350 1493 1351 1499
rect 1357 1498 2623 1499
rect 1357 1494 1367 1498
rect 1371 1494 1519 1498
rect 1523 1494 1575 1498
rect 1579 1494 1647 1498
rect 1651 1494 1663 1498
rect 1667 1494 1719 1498
rect 1723 1494 1727 1498
rect 1731 1494 1775 1498
rect 1779 1494 1807 1498
rect 1811 1494 1839 1498
rect 1843 1494 1895 1498
rect 1899 1494 1911 1498
rect 1915 1494 1983 1498
rect 1987 1494 1991 1498
rect 1995 1494 2071 1498
rect 2075 1494 2151 1498
rect 2155 1494 2231 1498
rect 2235 1494 2311 1498
rect 2315 1494 2391 1498
rect 2395 1494 2471 1498
rect 2475 1494 2527 1498
rect 2531 1494 2583 1498
rect 2587 1494 2623 1498
rect 1357 1493 2623 1494
rect 2629 1493 2630 1499
rect 1350 1491 1358 1493
rect 96 1485 97 1491
rect 103 1490 1351 1491
rect 103 1486 111 1490
rect 115 1486 199 1490
rect 203 1486 263 1490
rect 267 1486 287 1490
rect 291 1486 319 1490
rect 323 1486 383 1490
rect 387 1486 455 1490
rect 459 1486 487 1490
rect 491 1486 527 1490
rect 531 1486 583 1490
rect 587 1486 599 1490
rect 603 1486 671 1490
rect 675 1486 679 1490
rect 683 1486 743 1490
rect 747 1486 775 1490
rect 779 1486 815 1490
rect 819 1486 863 1490
rect 867 1486 887 1490
rect 891 1486 951 1490
rect 955 1486 959 1490
rect 963 1486 1039 1490
rect 1043 1486 1135 1490
rect 1139 1486 1327 1490
rect 1331 1486 1351 1490
rect 103 1485 1351 1486
rect 1357 1485 1358 1491
rect 1338 1434 2618 1435
rect 1338 1431 1367 1434
rect 84 1425 85 1431
rect 91 1430 1339 1431
rect 91 1426 111 1430
rect 115 1426 159 1430
rect 163 1426 215 1430
rect 219 1426 247 1430
rect 251 1426 303 1430
rect 307 1426 343 1430
rect 347 1426 399 1430
rect 403 1426 447 1430
rect 451 1426 503 1430
rect 507 1426 551 1430
rect 555 1426 599 1430
rect 603 1426 663 1430
rect 667 1426 695 1430
rect 699 1426 767 1430
rect 771 1426 791 1430
rect 795 1426 879 1430
rect 883 1426 967 1430
rect 971 1426 991 1430
rect 995 1426 1055 1430
rect 1059 1426 1103 1430
rect 1107 1426 1151 1430
rect 1155 1426 1215 1430
rect 1219 1426 1327 1430
rect 1331 1426 1339 1430
rect 91 1425 1339 1426
rect 1345 1430 1367 1431
rect 1371 1430 1415 1434
rect 1419 1430 1471 1434
rect 1475 1430 1535 1434
rect 1539 1430 1591 1434
rect 1595 1430 1623 1434
rect 1627 1430 1663 1434
rect 1667 1430 1719 1434
rect 1723 1430 1743 1434
rect 1747 1430 1823 1434
rect 1827 1430 1911 1434
rect 1915 1430 1927 1434
rect 1931 1430 1999 1434
rect 2003 1430 2023 1434
rect 2027 1430 2087 1434
rect 2091 1430 2119 1434
rect 2123 1430 2167 1434
rect 2171 1430 2215 1434
rect 2219 1430 2247 1434
rect 2251 1430 2303 1434
rect 2307 1430 2327 1434
rect 2331 1430 2391 1434
rect 2395 1430 2407 1434
rect 2411 1430 2479 1434
rect 2483 1430 2487 1434
rect 2491 1430 2543 1434
rect 2547 1430 2583 1434
rect 2587 1430 2618 1434
rect 1345 1429 2618 1430
rect 1345 1425 1346 1429
rect 96 1369 97 1375
rect 103 1374 1351 1375
rect 103 1370 111 1374
rect 115 1370 143 1374
rect 147 1370 207 1374
rect 211 1370 231 1374
rect 235 1370 295 1374
rect 299 1370 327 1374
rect 331 1370 399 1374
rect 403 1370 431 1374
rect 435 1370 511 1374
rect 515 1370 535 1374
rect 539 1370 623 1374
rect 627 1370 647 1374
rect 651 1370 735 1374
rect 739 1370 751 1374
rect 755 1370 847 1374
rect 851 1370 863 1374
rect 867 1370 959 1374
rect 963 1370 975 1374
rect 979 1370 1071 1374
rect 1075 1370 1087 1374
rect 1091 1370 1183 1374
rect 1187 1370 1199 1374
rect 1203 1370 1271 1374
rect 1275 1370 1327 1374
rect 1331 1370 1351 1374
rect 103 1369 1351 1370
rect 1357 1371 1358 1375
rect 1357 1370 2630 1371
rect 1357 1369 1367 1370
rect 1350 1366 1367 1369
rect 1371 1366 1399 1370
rect 1403 1366 1455 1370
rect 1459 1366 1519 1370
rect 1523 1366 1543 1370
rect 1547 1366 1607 1370
rect 1611 1366 1631 1370
rect 1635 1366 1703 1370
rect 1707 1366 1719 1370
rect 1723 1366 1807 1370
rect 1811 1366 1887 1370
rect 1891 1366 1911 1370
rect 1915 1366 1967 1370
rect 1971 1366 2007 1370
rect 2011 1366 2047 1370
rect 2051 1366 2103 1370
rect 2107 1366 2127 1370
rect 2131 1366 2199 1370
rect 2203 1366 2207 1370
rect 2211 1366 2287 1370
rect 2291 1366 2375 1370
rect 2379 1366 2463 1370
rect 2467 1366 2527 1370
rect 2531 1366 2583 1370
rect 2587 1366 2630 1370
rect 1350 1365 2630 1366
rect 1406 1356 1412 1357
rect 1750 1356 1756 1357
rect 1406 1352 1407 1356
rect 1411 1352 1751 1356
rect 1755 1352 1756 1356
rect 1406 1351 1412 1352
rect 1750 1351 1756 1352
rect 890 1332 896 1333
rect 1294 1332 1300 1333
rect 890 1328 891 1332
rect 895 1328 1295 1332
rect 1299 1328 1300 1332
rect 890 1327 896 1328
rect 1294 1327 1300 1328
rect 84 1313 85 1319
rect 91 1318 1339 1319
rect 91 1314 111 1318
rect 115 1314 159 1318
rect 163 1314 223 1318
rect 227 1314 231 1318
rect 235 1314 311 1318
rect 315 1314 327 1318
rect 331 1314 415 1318
rect 419 1314 431 1318
rect 435 1314 527 1318
rect 531 1314 535 1318
rect 539 1314 631 1318
rect 635 1314 639 1318
rect 643 1314 727 1318
rect 731 1314 751 1318
rect 755 1314 823 1318
rect 827 1314 863 1318
rect 867 1314 911 1318
rect 915 1314 975 1318
rect 979 1314 991 1318
rect 995 1314 1071 1318
rect 1075 1314 1087 1318
rect 1091 1314 1151 1318
rect 1155 1314 1199 1318
rect 1203 1314 1231 1318
rect 1235 1314 1287 1318
rect 1291 1314 1327 1318
rect 1331 1314 1339 1318
rect 91 1313 1339 1314
rect 1345 1313 1346 1319
rect 1338 1311 1346 1313
rect 1338 1305 1339 1311
rect 1345 1310 2611 1311
rect 1345 1306 1367 1310
rect 1371 1306 1415 1310
rect 1419 1306 1471 1310
rect 1475 1306 1559 1310
rect 1563 1306 1647 1310
rect 1651 1306 1671 1310
rect 1675 1306 1735 1310
rect 1739 1306 1767 1310
rect 1771 1306 1823 1310
rect 1827 1306 1863 1310
rect 1867 1306 1903 1310
rect 1907 1306 1959 1310
rect 1963 1306 1983 1310
rect 1987 1306 2047 1310
rect 2051 1306 2063 1310
rect 2067 1306 2135 1310
rect 2139 1306 2143 1310
rect 2147 1306 2223 1310
rect 2227 1306 2231 1310
rect 2235 1306 2583 1310
rect 2587 1306 2611 1310
rect 1345 1305 2611 1306
rect 2617 1305 2618 1311
rect 1350 1254 2630 1255
rect 1350 1251 1367 1254
rect 96 1245 97 1251
rect 103 1250 1351 1251
rect 103 1246 111 1250
rect 115 1246 143 1250
rect 147 1246 199 1250
rect 203 1246 215 1250
rect 219 1246 279 1250
rect 283 1246 311 1250
rect 315 1246 359 1250
rect 363 1246 415 1250
rect 419 1246 439 1250
rect 443 1246 519 1250
rect 523 1246 599 1250
rect 603 1246 615 1250
rect 619 1246 671 1250
rect 675 1246 711 1250
rect 715 1246 743 1250
rect 747 1246 807 1250
rect 811 1246 815 1250
rect 819 1246 895 1250
rect 899 1246 975 1250
rect 979 1246 1055 1250
rect 1059 1246 1135 1250
rect 1139 1246 1215 1250
rect 1219 1246 1271 1250
rect 1275 1246 1327 1250
rect 1331 1246 1351 1250
rect 103 1245 1351 1246
rect 1357 1250 1367 1251
rect 1371 1250 1495 1254
rect 1499 1250 1559 1254
rect 1563 1250 1623 1254
rect 1627 1250 1655 1254
rect 1659 1250 1687 1254
rect 1691 1250 1751 1254
rect 1755 1250 1759 1254
rect 1763 1250 1823 1254
rect 1827 1250 1847 1254
rect 1851 1250 1887 1254
rect 1891 1250 1943 1254
rect 1947 1250 1951 1254
rect 1955 1250 2015 1254
rect 2019 1250 2031 1254
rect 2035 1250 2079 1254
rect 2083 1250 2119 1254
rect 2123 1250 2151 1254
rect 2155 1250 2215 1254
rect 2219 1250 2223 1254
rect 2227 1250 2295 1254
rect 2299 1250 2583 1254
rect 2587 1250 2630 1254
rect 1357 1249 2630 1250
rect 1357 1245 1358 1249
rect 84 1185 85 1191
rect 91 1190 1339 1191
rect 91 1186 111 1190
rect 115 1186 159 1190
rect 163 1186 215 1190
rect 219 1186 239 1190
rect 243 1186 295 1190
rect 299 1186 327 1190
rect 331 1186 375 1190
rect 379 1186 423 1190
rect 427 1186 455 1190
rect 459 1186 511 1190
rect 515 1186 535 1190
rect 539 1186 599 1190
rect 603 1186 615 1190
rect 619 1186 687 1190
rect 691 1186 759 1190
rect 763 1186 767 1190
rect 771 1186 831 1190
rect 835 1186 839 1190
rect 843 1186 911 1190
rect 915 1186 983 1190
rect 987 1186 1063 1190
rect 1067 1186 1327 1190
rect 1331 1186 1339 1190
rect 91 1185 1339 1186
rect 1345 1190 2618 1191
rect 1345 1186 1367 1190
rect 1371 1186 1415 1190
rect 1419 1186 1503 1190
rect 1507 1186 1511 1190
rect 1515 1186 1575 1190
rect 1579 1186 1599 1190
rect 1603 1186 1639 1190
rect 1643 1186 1703 1190
rect 1707 1186 1775 1190
rect 1779 1186 1807 1190
rect 1811 1186 1839 1190
rect 1843 1186 1903 1190
rect 1907 1186 1911 1190
rect 1915 1186 1967 1190
rect 1971 1186 2015 1190
rect 2019 1186 2031 1190
rect 2035 1186 2095 1190
rect 2099 1186 2111 1190
rect 2115 1186 2167 1190
rect 2171 1186 2207 1190
rect 2211 1186 2239 1190
rect 2243 1186 2303 1190
rect 2307 1186 2311 1190
rect 2315 1186 2399 1190
rect 2403 1186 2583 1190
rect 2587 1186 2618 1190
rect 1345 1185 2618 1186
rect 1350 1130 2630 1131
rect 1350 1127 1367 1130
rect 96 1121 97 1127
rect 103 1126 1351 1127
rect 103 1122 111 1126
rect 115 1122 143 1126
rect 147 1122 223 1126
rect 227 1122 311 1126
rect 315 1122 319 1126
rect 323 1122 407 1126
rect 411 1122 423 1126
rect 427 1122 495 1126
rect 499 1122 527 1126
rect 531 1122 583 1126
rect 587 1122 631 1126
rect 635 1122 671 1126
rect 675 1122 727 1126
rect 731 1122 751 1126
rect 755 1122 823 1126
rect 827 1122 895 1126
rect 899 1122 911 1126
rect 915 1122 967 1126
rect 971 1122 991 1126
rect 995 1122 1047 1126
rect 1051 1122 1079 1126
rect 1083 1122 1167 1126
rect 1171 1122 1327 1126
rect 1331 1122 1351 1126
rect 103 1121 1351 1122
rect 1357 1126 1367 1127
rect 1371 1126 1399 1130
rect 1403 1126 1479 1130
rect 1483 1126 1487 1130
rect 1491 1126 1583 1130
rect 1587 1126 1687 1130
rect 1691 1126 1791 1130
rect 1795 1126 1887 1130
rect 1891 1126 1895 1130
rect 1899 1126 1975 1130
rect 1979 1126 1999 1130
rect 2003 1126 2063 1130
rect 2067 1126 2095 1130
rect 2099 1126 2143 1130
rect 2147 1126 2191 1130
rect 2195 1126 2215 1130
rect 2219 1126 2279 1130
rect 2283 1126 2287 1130
rect 2291 1126 2343 1130
rect 2347 1126 2383 1130
rect 2387 1126 2407 1130
rect 2411 1126 2471 1130
rect 2475 1126 2527 1130
rect 2531 1126 2583 1130
rect 2587 1126 2630 1130
rect 1357 1125 2630 1126
rect 1357 1121 1358 1125
rect 218 1084 224 1085
rect 550 1084 556 1085
rect 218 1080 219 1084
rect 223 1080 551 1084
rect 555 1080 556 1084
rect 218 1079 224 1080
rect 550 1079 556 1080
rect 1338 1070 2618 1071
rect 1338 1067 1367 1070
rect 84 1061 85 1067
rect 91 1066 1339 1067
rect 91 1062 111 1066
rect 115 1062 239 1066
rect 243 1062 311 1066
rect 315 1062 335 1066
rect 339 1062 367 1066
rect 371 1062 439 1066
rect 443 1062 519 1066
rect 523 1062 543 1066
rect 547 1062 607 1066
rect 611 1062 647 1066
rect 651 1062 703 1066
rect 707 1062 743 1066
rect 747 1062 799 1066
rect 803 1062 839 1066
rect 843 1062 887 1066
rect 891 1062 927 1066
rect 931 1062 975 1066
rect 979 1062 1007 1066
rect 1011 1062 1055 1066
rect 1059 1062 1095 1066
rect 1099 1062 1135 1066
rect 1139 1062 1183 1066
rect 1187 1062 1223 1066
rect 1227 1062 1287 1066
rect 1291 1062 1327 1066
rect 1331 1062 1339 1066
rect 91 1061 1339 1062
rect 1345 1066 1367 1067
rect 1371 1066 1415 1070
rect 1419 1066 1471 1070
rect 1475 1066 1495 1070
rect 1499 1066 1535 1070
rect 1539 1066 1599 1070
rect 1603 1066 1623 1070
rect 1627 1066 1703 1070
rect 1707 1066 1727 1070
rect 1731 1066 1807 1070
rect 1811 1066 1839 1070
rect 1843 1066 1903 1070
rect 1907 1066 1951 1070
rect 1955 1066 1991 1070
rect 1995 1066 2063 1070
rect 2067 1066 2079 1070
rect 2083 1066 2159 1070
rect 2163 1066 2167 1070
rect 2171 1066 2231 1070
rect 2235 1066 2271 1070
rect 2275 1066 2295 1070
rect 2299 1066 2359 1070
rect 2363 1066 2367 1070
rect 2371 1066 2423 1070
rect 2427 1066 2463 1070
rect 2467 1066 2487 1070
rect 2491 1066 2543 1070
rect 2547 1066 2583 1070
rect 2587 1066 2618 1070
rect 1345 1065 2618 1066
rect 1345 1061 1346 1065
rect 878 1028 884 1029
rect 1234 1028 1240 1029
rect 878 1024 879 1028
rect 883 1024 1235 1028
rect 1239 1024 1240 1028
rect 878 1023 884 1024
rect 1234 1023 1240 1024
rect 96 1001 97 1007
rect 103 1006 1351 1007
rect 103 1002 111 1006
rect 115 1002 295 1006
rect 299 1002 351 1006
rect 355 1002 415 1006
rect 419 1002 423 1006
rect 427 1002 471 1006
rect 475 1002 503 1006
rect 507 1002 527 1006
rect 531 1002 591 1006
rect 595 1002 655 1006
rect 659 1002 687 1006
rect 691 1002 719 1006
rect 723 1002 783 1006
rect 787 1002 847 1006
rect 851 1002 871 1006
rect 875 1002 911 1006
rect 915 1002 959 1006
rect 963 1002 975 1006
rect 979 1002 1039 1006
rect 1043 1002 1103 1006
rect 1107 1002 1119 1006
rect 1123 1002 1159 1006
rect 1163 1002 1207 1006
rect 1211 1002 1215 1006
rect 1219 1002 1271 1006
rect 1275 1002 1327 1006
rect 1331 1002 1351 1006
rect 103 1001 1351 1002
rect 1357 1001 1358 1007
rect 1350 999 1358 1001
rect 1350 993 1351 999
rect 1357 998 2623 999
rect 1357 994 1367 998
rect 1371 994 1399 998
rect 1403 994 1455 998
rect 1459 994 1511 998
rect 1515 994 1519 998
rect 1523 994 1567 998
rect 1571 994 1607 998
rect 1611 994 1639 998
rect 1643 994 1711 998
rect 1715 994 1719 998
rect 1723 994 1807 998
rect 1811 994 1823 998
rect 1827 994 1903 998
rect 1907 994 1935 998
rect 1939 994 2015 998
rect 2019 994 2047 998
rect 2051 994 2143 998
rect 2147 994 2151 998
rect 2155 994 2255 998
rect 2259 994 2271 998
rect 2275 994 2351 998
rect 2355 994 2407 998
rect 2411 994 2447 998
rect 2451 994 2527 998
rect 2531 994 2583 998
rect 2587 994 2623 998
rect 1357 993 2623 994
rect 2629 993 2630 999
rect 84 941 85 947
rect 91 946 1339 947
rect 91 942 111 946
rect 115 942 423 946
rect 427 942 431 946
rect 435 942 479 946
rect 483 942 487 946
rect 491 942 535 946
rect 539 942 543 946
rect 547 942 591 946
rect 595 942 607 946
rect 611 942 647 946
rect 651 942 671 946
rect 675 942 703 946
rect 707 942 735 946
rect 739 942 759 946
rect 763 942 799 946
rect 803 942 815 946
rect 819 942 863 946
rect 867 942 927 946
rect 931 942 991 946
rect 995 942 1055 946
rect 1059 942 1119 946
rect 1123 942 1175 946
rect 1179 942 1231 946
rect 1235 942 1287 946
rect 1291 942 1327 946
rect 1331 942 1339 946
rect 91 941 1339 942
rect 1345 941 1346 947
rect 1338 929 1339 935
rect 1345 934 2611 935
rect 1345 930 1367 934
rect 1371 930 1415 934
rect 1419 930 1471 934
rect 1475 930 1527 934
rect 1531 930 1583 934
rect 1587 930 1615 934
rect 1619 930 1655 934
rect 1659 930 1711 934
rect 1715 930 1735 934
rect 1739 930 1823 934
rect 1827 930 1919 934
rect 1923 930 1943 934
rect 1947 930 2031 934
rect 2035 930 2063 934
rect 2067 930 2159 934
rect 2163 930 2183 934
rect 2187 930 2287 934
rect 2291 930 2311 934
rect 2315 930 2423 934
rect 2427 930 2439 934
rect 2443 930 2543 934
rect 2547 930 2583 934
rect 2587 930 2611 934
rect 1345 929 2611 930
rect 2617 929 2618 935
rect 96 885 97 891
rect 103 890 1351 891
rect 103 886 111 890
rect 115 886 279 890
rect 283 886 335 890
rect 339 886 391 890
rect 395 886 407 890
rect 411 886 455 890
rect 459 886 463 890
rect 467 886 519 890
rect 523 886 575 890
rect 579 886 583 890
rect 587 886 631 890
rect 635 886 647 890
rect 651 886 687 890
rect 691 886 711 890
rect 715 886 743 890
rect 747 886 775 890
rect 779 886 799 890
rect 803 886 847 890
rect 851 886 919 890
rect 923 886 1327 890
rect 1331 886 1351 890
rect 103 885 1351 886
rect 1357 885 1358 891
rect 1350 873 1351 879
rect 1357 878 2623 879
rect 1357 874 1367 878
rect 1371 874 1399 878
rect 1403 874 1455 878
rect 1459 874 1471 878
rect 1475 874 1511 878
rect 1515 874 1551 878
rect 1555 874 1599 878
rect 1603 874 1639 878
rect 1643 874 1695 878
rect 1699 874 1727 878
rect 1731 874 1807 878
rect 1811 874 1815 878
rect 1819 874 1903 878
rect 1907 874 1927 878
rect 1931 874 1991 878
rect 1995 874 2047 878
rect 2051 874 2071 878
rect 2075 874 2143 878
rect 2147 874 2167 878
rect 2171 874 2215 878
rect 2219 874 2279 878
rect 2283 874 2295 878
rect 2299 874 2343 878
rect 2347 874 2407 878
rect 2411 874 2423 878
rect 2427 874 2471 878
rect 2475 874 2527 878
rect 2531 874 2583 878
rect 2587 874 2623 878
rect 1357 873 2623 874
rect 2629 873 2630 879
rect 84 821 85 827
rect 91 826 1339 827
rect 91 822 111 826
rect 115 822 167 826
rect 171 822 231 826
rect 235 822 295 826
rect 299 822 311 826
rect 315 822 351 826
rect 355 822 399 826
rect 403 822 407 826
rect 411 822 471 826
rect 475 822 487 826
rect 491 822 535 826
rect 539 822 583 826
rect 587 822 599 826
rect 603 822 663 826
rect 667 822 671 826
rect 675 822 727 826
rect 731 822 759 826
rect 763 822 791 826
rect 795 822 839 826
rect 843 822 863 826
rect 867 822 919 826
rect 923 822 935 826
rect 939 822 1007 826
rect 1011 822 1095 826
rect 1099 822 1327 826
rect 1331 822 1339 826
rect 91 821 1339 822
rect 1345 821 1346 827
rect 1338 809 1339 815
rect 1345 814 2611 815
rect 1345 810 1367 814
rect 1371 810 1487 814
rect 1491 810 1567 814
rect 1571 810 1631 814
rect 1635 810 1655 814
rect 1659 810 1687 814
rect 1691 810 1743 814
rect 1747 810 1751 814
rect 1755 810 1823 814
rect 1827 810 1831 814
rect 1835 810 1903 814
rect 1907 810 1919 814
rect 1923 810 1991 814
rect 1995 810 2007 814
rect 2011 810 2071 814
rect 2075 810 2087 814
rect 2091 810 2159 814
rect 2163 810 2231 814
rect 2235 810 2247 814
rect 2251 810 2295 814
rect 2299 810 2335 814
rect 2339 810 2359 814
rect 2363 810 2423 814
rect 2427 810 2487 814
rect 2491 810 2543 814
rect 2547 810 2583 814
rect 2587 810 2611 814
rect 1345 809 2611 810
rect 2617 809 2618 815
rect 2126 780 2132 781
rect 2438 780 2444 781
rect 2126 776 2127 780
rect 2131 776 2439 780
rect 2443 776 2444 780
rect 2126 775 2132 776
rect 2438 775 2444 776
rect 96 757 97 763
rect 103 762 1351 763
rect 103 758 111 762
rect 115 758 143 762
rect 147 758 151 762
rect 155 758 199 762
rect 203 758 215 762
rect 219 758 279 762
rect 283 758 295 762
rect 299 758 383 762
rect 387 758 471 762
rect 475 758 487 762
rect 491 758 567 762
rect 571 758 599 762
rect 603 758 655 762
rect 659 758 703 762
rect 707 758 743 762
rect 747 758 807 762
rect 811 758 823 762
rect 827 758 903 762
rect 907 758 991 762
rect 995 758 1079 762
rect 1083 758 1175 762
rect 1179 758 1327 762
rect 1331 758 1351 762
rect 103 757 1351 758
rect 1357 757 1358 763
rect 1350 755 1358 757
rect 1350 749 1351 755
rect 1357 754 2623 755
rect 1357 750 1367 754
rect 1371 750 1567 754
rect 1571 750 1615 754
rect 1619 750 1623 754
rect 1627 750 1671 754
rect 1675 750 1687 754
rect 1691 750 1735 754
rect 1739 750 1759 754
rect 1763 750 1807 754
rect 1811 750 1839 754
rect 1843 750 1887 754
rect 1891 750 1919 754
rect 1923 750 1975 754
rect 1979 750 1999 754
rect 2003 750 2055 754
rect 2059 750 2079 754
rect 2083 750 2143 754
rect 2147 750 2159 754
rect 2163 750 2231 754
rect 2235 750 2247 754
rect 2251 750 2319 754
rect 2323 750 2335 754
rect 2339 750 2407 754
rect 2411 750 2583 754
rect 2587 750 2623 754
rect 1357 749 2623 750
rect 2629 749 2630 755
rect 698 716 704 717
rect 1102 716 1108 717
rect 698 712 699 716
rect 703 712 1103 716
rect 1107 712 1108 716
rect 698 711 704 712
rect 1102 711 1108 712
rect 84 697 85 703
rect 91 702 1339 703
rect 91 698 111 702
rect 115 698 159 702
rect 163 698 215 702
rect 219 698 279 702
rect 283 698 295 702
rect 299 698 359 702
rect 363 698 399 702
rect 403 698 447 702
rect 451 698 503 702
rect 507 698 535 702
rect 539 698 615 702
rect 619 698 623 702
rect 627 698 711 702
rect 715 698 719 702
rect 723 698 791 702
rect 795 698 823 702
rect 827 698 871 702
rect 875 698 919 702
rect 923 698 951 702
rect 955 698 1007 702
rect 1011 698 1039 702
rect 1043 698 1095 702
rect 1099 698 1191 702
rect 1195 698 1327 702
rect 1331 698 1339 702
rect 91 697 1339 698
rect 1345 697 1346 703
rect 1338 695 1346 697
rect 1338 689 1339 695
rect 1345 694 2611 695
rect 1345 690 1367 694
rect 1371 690 1415 694
rect 1419 690 1511 694
rect 1515 690 1583 694
rect 1587 690 1615 694
rect 1619 690 1639 694
rect 1643 690 1703 694
rect 1707 690 1719 694
rect 1723 690 1775 694
rect 1779 690 1823 694
rect 1827 690 1855 694
rect 1859 690 1927 694
rect 1931 690 1935 694
rect 1939 690 2015 694
rect 2019 690 2023 694
rect 2027 690 2095 694
rect 2099 690 2119 694
rect 2123 690 2175 694
rect 2179 690 2207 694
rect 2211 690 2263 694
rect 2267 690 2295 694
rect 2299 690 2351 694
rect 2355 690 2391 694
rect 2395 690 2583 694
rect 2587 690 2611 694
rect 1345 689 2611 690
rect 2617 689 2618 695
rect 96 633 97 639
rect 103 638 1351 639
rect 103 634 111 638
rect 115 634 143 638
rect 147 634 199 638
rect 203 634 255 638
rect 259 634 263 638
rect 267 634 311 638
rect 315 634 343 638
rect 347 634 391 638
rect 395 634 431 638
rect 435 634 479 638
rect 483 634 519 638
rect 523 634 575 638
rect 579 634 607 638
rect 611 634 679 638
rect 683 634 695 638
rect 699 634 775 638
rect 779 634 783 638
rect 787 634 855 638
rect 859 634 887 638
rect 891 634 935 638
rect 939 634 991 638
rect 995 634 1023 638
rect 1027 634 1087 638
rect 1091 634 1191 638
rect 1195 634 1271 638
rect 1275 634 1327 638
rect 1331 634 1351 638
rect 103 633 1351 634
rect 1357 638 2630 639
rect 1357 634 1367 638
rect 1371 634 1399 638
rect 1403 634 1495 638
rect 1499 634 1511 638
rect 1515 634 1599 638
rect 1603 634 1647 638
rect 1651 634 1703 638
rect 1707 634 1783 638
rect 1787 634 1807 638
rect 1811 634 1911 638
rect 1915 634 2007 638
rect 2011 634 2039 638
rect 2043 634 2103 638
rect 2107 634 2159 638
rect 2163 634 2191 638
rect 2195 634 2279 638
rect 2283 634 2375 638
rect 2379 634 2407 638
rect 2411 634 2583 638
rect 2587 634 2630 638
rect 1357 633 2630 634
rect 1406 628 1412 629
rect 1814 628 1820 629
rect 1406 624 1407 628
rect 1411 624 1815 628
rect 1819 624 1820 628
rect 1406 623 1412 624
rect 1814 623 1820 624
rect 84 573 85 579
rect 91 578 1339 579
rect 91 574 111 578
rect 115 574 159 578
rect 163 574 199 578
rect 203 574 215 578
rect 219 574 263 578
rect 267 574 271 578
rect 275 574 327 578
rect 331 574 335 578
rect 339 574 407 578
rect 411 574 415 578
rect 419 574 495 578
rect 499 574 511 578
rect 515 574 591 578
rect 595 574 615 578
rect 619 574 695 578
rect 699 574 719 578
rect 723 574 799 578
rect 803 574 831 578
rect 835 574 903 578
rect 907 574 943 578
rect 947 574 1007 578
rect 1011 574 1063 578
rect 1067 574 1103 578
rect 1107 574 1183 578
rect 1187 574 1207 578
rect 1211 574 1287 578
rect 1291 574 1327 578
rect 1331 574 1339 578
rect 91 573 1339 574
rect 1345 575 1346 579
rect 1345 574 2618 575
rect 1345 573 1367 574
rect 1338 570 1367 573
rect 1371 570 1415 574
rect 1419 570 1471 574
rect 1475 570 1527 574
rect 1531 570 1551 574
rect 1555 570 1647 574
rect 1651 570 1663 574
rect 1667 570 1751 574
rect 1755 570 1799 574
rect 1803 570 1855 574
rect 1859 570 1927 574
rect 1931 570 1959 574
rect 1963 570 2055 574
rect 2059 570 2151 574
rect 2155 570 2175 574
rect 2179 570 2239 574
rect 2243 570 2295 574
rect 2299 570 2319 574
rect 2323 570 2399 574
rect 2403 570 2423 574
rect 2427 570 2479 574
rect 2483 570 2543 574
rect 2547 570 2583 574
rect 2587 570 2618 574
rect 1338 569 2618 570
rect 1350 518 2630 519
rect 1350 515 1367 518
rect 96 509 97 515
rect 103 514 1351 515
rect 103 510 111 514
rect 115 510 183 514
rect 187 510 247 514
rect 251 510 303 514
rect 307 510 319 514
rect 323 510 359 514
rect 363 510 399 514
rect 403 510 423 514
rect 427 510 495 514
rect 499 510 575 514
rect 579 510 599 514
rect 603 510 647 514
rect 651 510 703 514
rect 707 510 719 514
rect 723 510 791 514
rect 795 510 815 514
rect 819 510 863 514
rect 867 510 927 514
rect 931 510 935 514
rect 939 510 1007 514
rect 1011 510 1047 514
rect 1051 510 1087 514
rect 1091 510 1167 514
rect 1171 510 1271 514
rect 1275 510 1327 514
rect 1331 510 1351 514
rect 103 509 1351 510
rect 1357 514 1367 515
rect 1371 514 1399 518
rect 1403 514 1455 518
rect 1459 514 1535 518
rect 1539 514 1599 518
rect 1603 514 1631 518
rect 1635 514 1671 518
rect 1675 514 1735 518
rect 1739 514 1751 518
rect 1755 514 1839 518
rect 1843 514 1927 518
rect 1931 514 1943 518
rect 1947 514 2015 518
rect 2019 514 2039 518
rect 2043 514 2095 518
rect 2099 514 2135 518
rect 2139 514 2175 518
rect 2179 514 2223 518
rect 2227 514 2255 518
rect 2259 514 2303 518
rect 2307 514 2327 518
rect 2331 514 2383 518
rect 2387 514 2399 518
rect 2403 514 2463 518
rect 2467 514 2471 518
rect 2475 514 2527 518
rect 2531 514 2583 518
rect 2587 514 2630 518
rect 1357 513 2630 514
rect 1357 509 1358 513
rect 84 449 85 455
rect 91 454 1339 455
rect 91 450 111 454
rect 115 450 319 454
rect 323 450 375 454
rect 379 450 439 454
rect 443 450 455 454
rect 459 450 511 454
rect 515 450 575 454
rect 579 450 591 454
rect 595 450 647 454
rect 651 450 663 454
rect 667 450 727 454
rect 731 450 735 454
rect 739 450 799 454
rect 803 450 807 454
rect 811 450 871 454
rect 875 450 879 454
rect 883 450 943 454
rect 947 450 951 454
rect 955 450 1015 454
rect 1019 450 1023 454
rect 1027 450 1087 454
rect 1091 450 1103 454
rect 1107 450 1159 454
rect 1163 450 1239 454
rect 1243 450 1327 454
rect 1331 450 1339 454
rect 91 449 1339 450
rect 1345 454 2618 455
rect 1345 450 1367 454
rect 1371 450 1551 454
rect 1555 450 1615 454
rect 1619 450 1647 454
rect 1651 450 1687 454
rect 1691 450 1703 454
rect 1707 450 1759 454
rect 1763 450 1767 454
rect 1771 450 1815 454
rect 1819 450 1855 454
rect 1859 450 1871 454
rect 1875 450 1927 454
rect 1931 450 1943 454
rect 1947 450 1999 454
rect 2003 450 2031 454
rect 2035 450 2087 454
rect 2091 450 2111 454
rect 2115 450 2191 454
rect 2195 450 2271 454
rect 2275 450 2311 454
rect 2315 450 2343 454
rect 2347 450 2415 454
rect 2419 450 2439 454
rect 2443 450 2487 454
rect 2491 450 2543 454
rect 2547 450 2583 454
rect 2587 450 2618 454
rect 1345 449 2618 450
rect 2078 420 2084 421
rect 2454 420 2460 421
rect 2078 416 2079 420
rect 2083 416 2455 420
rect 2459 416 2460 420
rect 2078 415 2084 416
rect 2454 415 2460 416
rect 1350 398 2630 399
rect 1350 395 1367 398
rect 96 389 97 395
rect 103 394 1351 395
rect 103 390 111 394
rect 115 390 415 394
rect 419 390 439 394
rect 443 390 471 394
rect 475 390 495 394
rect 499 390 535 394
rect 539 390 559 394
rect 563 390 607 394
rect 611 390 631 394
rect 635 390 687 394
rect 691 390 711 394
rect 715 390 767 394
rect 771 390 783 394
rect 787 390 847 394
rect 851 390 855 394
rect 859 390 927 394
rect 931 390 999 394
rect 1003 390 1007 394
rect 1011 390 1071 394
rect 1075 390 1087 394
rect 1091 390 1143 394
rect 1147 390 1175 394
rect 1179 390 1223 394
rect 1227 390 1263 394
rect 1267 390 1327 394
rect 1331 390 1351 394
rect 103 389 1351 390
rect 1357 394 1367 395
rect 1371 394 1631 398
rect 1635 394 1655 398
rect 1659 394 1687 398
rect 1691 394 1711 398
rect 1715 394 1743 398
rect 1747 394 1767 398
rect 1771 394 1799 398
rect 1803 394 1823 398
rect 1827 394 1855 398
rect 1859 394 1879 398
rect 1883 394 1911 398
rect 1915 394 1951 398
rect 1955 394 1983 398
rect 1987 394 2039 398
rect 2043 394 2071 398
rect 2075 394 2151 398
rect 2155 394 2175 398
rect 2179 394 2279 398
rect 2283 394 2295 398
rect 2299 394 2415 398
rect 2419 394 2423 398
rect 2427 394 2527 398
rect 2531 394 2583 398
rect 2587 394 2630 398
rect 1357 393 2630 394
rect 1357 389 1358 393
rect 2122 356 2128 357
rect 2438 356 2444 357
rect 2122 352 2123 356
rect 2127 352 2439 356
rect 2443 352 2444 356
rect 2122 351 2128 352
rect 2438 351 2444 352
rect 84 329 85 335
rect 91 334 1339 335
rect 91 330 111 334
rect 115 330 431 334
rect 435 330 463 334
rect 467 330 487 334
rect 491 330 519 334
rect 523 330 551 334
rect 555 330 575 334
rect 579 330 623 334
rect 627 330 631 334
rect 635 330 695 334
rect 699 330 703 334
rect 707 330 767 334
rect 771 330 783 334
rect 787 330 847 334
rect 851 330 863 334
rect 867 330 927 334
rect 931 330 943 334
rect 947 330 1015 334
rect 1019 330 1023 334
rect 1027 330 1103 334
rect 1107 330 1111 334
rect 1115 330 1191 334
rect 1195 330 1215 334
rect 1219 330 1279 334
rect 1283 330 1327 334
rect 1331 330 1339 334
rect 91 329 1339 330
rect 1345 334 2618 335
rect 1345 330 1367 334
rect 1371 330 1631 334
rect 1635 330 1671 334
rect 1675 330 1687 334
rect 1691 330 1727 334
rect 1731 330 1743 334
rect 1747 330 1783 334
rect 1787 330 1807 334
rect 1811 330 1839 334
rect 1843 330 1887 334
rect 1891 330 1895 334
rect 1899 330 1967 334
rect 1971 330 2055 334
rect 2059 330 2143 334
rect 2147 330 2167 334
rect 2171 330 2231 334
rect 2235 330 2295 334
rect 2299 330 2311 334
rect 2315 330 2391 334
rect 2395 330 2431 334
rect 2435 330 2479 334
rect 2483 330 2543 334
rect 2547 330 2583 334
rect 2587 330 2618 334
rect 1345 329 2618 330
rect 1350 278 2630 279
rect 1350 275 1367 278
rect 96 269 97 275
rect 103 274 1351 275
rect 103 270 111 274
rect 115 270 287 274
rect 291 270 359 274
rect 363 270 439 274
rect 443 270 447 274
rect 451 270 503 274
rect 507 270 527 274
rect 531 270 559 274
rect 563 270 615 274
rect 619 270 623 274
rect 627 270 679 274
rect 683 270 719 274
rect 723 270 751 274
rect 755 270 823 274
rect 827 270 831 274
rect 835 270 911 274
rect 915 270 927 274
rect 931 270 999 274
rect 1003 270 1031 274
rect 1035 270 1095 274
rect 1099 270 1143 274
rect 1147 270 1199 274
rect 1203 270 1255 274
rect 1259 270 1327 274
rect 1331 270 1351 274
rect 103 269 1351 270
rect 1357 274 1367 275
rect 1371 274 1535 278
rect 1539 274 1607 278
rect 1611 274 1615 278
rect 1619 274 1671 278
rect 1675 274 1687 278
rect 1691 274 1727 278
rect 1731 274 1775 278
rect 1779 274 1791 278
rect 1795 274 1863 278
rect 1867 274 1871 278
rect 1875 274 1951 278
rect 1955 274 2039 278
rect 2043 274 2119 278
rect 2123 274 2127 278
rect 2131 274 2199 278
rect 2203 274 2215 278
rect 2219 274 2271 278
rect 2275 274 2295 278
rect 2299 274 2335 278
rect 2339 274 2375 278
rect 2379 274 2407 278
rect 2411 274 2463 278
rect 2467 274 2471 278
rect 2475 274 2527 278
rect 2531 274 2583 278
rect 2587 274 2630 278
rect 1357 273 2630 274
rect 1357 269 1358 273
rect 1338 222 2618 223
rect 1338 219 1367 222
rect 84 213 85 219
rect 91 218 1339 219
rect 91 214 111 218
rect 115 214 199 218
rect 203 214 271 218
rect 275 214 303 218
rect 307 214 359 218
rect 363 214 375 218
rect 379 214 455 218
rect 459 214 463 218
rect 467 214 543 218
rect 547 214 567 218
rect 571 214 639 218
rect 643 214 679 218
rect 683 214 735 218
rect 739 214 791 218
rect 795 214 839 218
rect 843 214 911 218
rect 915 214 943 218
rect 947 214 1031 218
rect 1035 214 1047 218
rect 1051 214 1151 218
rect 1155 214 1159 218
rect 1163 214 1271 218
rect 1275 214 1327 218
rect 1331 214 1339 218
rect 91 213 1339 214
rect 1345 218 1367 219
rect 1371 218 1415 222
rect 1419 218 1479 222
rect 1483 218 1551 222
rect 1555 218 1559 222
rect 1563 218 1623 222
rect 1627 218 1655 222
rect 1659 218 1703 222
rect 1707 218 1751 222
rect 1755 218 1791 222
rect 1795 218 1855 222
rect 1859 218 1879 222
rect 1883 218 1959 222
rect 1963 218 1967 222
rect 1971 218 2055 222
rect 2059 218 2063 222
rect 2067 218 2135 222
rect 2139 218 2167 222
rect 2171 218 2215 222
rect 2219 218 2263 222
rect 2267 218 2287 222
rect 2291 218 2351 222
rect 2355 218 2359 222
rect 2363 218 2423 222
rect 2427 218 2463 222
rect 2467 218 2487 222
rect 2491 218 2543 222
rect 2547 218 2583 222
rect 2587 218 2618 222
rect 1345 217 2618 218
rect 1345 213 1346 217
rect 1590 188 1596 189
rect 1870 188 1876 189
rect 1590 184 1591 188
rect 1595 184 1871 188
rect 1875 184 1876 188
rect 1590 183 1596 184
rect 1870 183 1876 184
rect 190 164 196 165
rect 622 164 628 165
rect 190 160 191 164
rect 195 160 623 164
rect 627 160 628 164
rect 190 159 196 160
rect 622 159 628 160
rect 1350 145 1351 151
rect 1357 150 2623 151
rect 1357 146 1367 150
rect 1371 146 1399 150
rect 1403 146 1455 150
rect 1459 146 1463 150
rect 1467 146 1511 150
rect 1515 146 1543 150
rect 1547 146 1567 150
rect 1571 146 1631 150
rect 1635 146 1639 150
rect 1643 146 1711 150
rect 1715 146 1735 150
rect 1739 146 1791 150
rect 1795 146 1839 150
rect 1843 146 1871 150
rect 1875 146 1943 150
rect 1947 146 2015 150
rect 2019 146 2047 150
rect 2051 146 2079 150
rect 2083 146 2143 150
rect 2147 146 2151 150
rect 2155 146 2207 150
rect 2211 146 2247 150
rect 2251 146 2271 150
rect 2275 146 2343 150
rect 2347 146 2415 150
rect 2419 146 2447 150
rect 2451 146 2527 150
rect 2531 146 2583 150
rect 2587 146 2623 150
rect 1357 145 2623 146
rect 2629 145 2630 151
rect 1406 140 1412 141
rect 1822 140 1828 141
rect 96 133 97 139
rect 103 138 1351 139
rect 103 134 111 138
rect 115 134 143 138
rect 147 134 183 138
rect 187 134 199 138
rect 203 134 255 138
rect 259 134 311 138
rect 315 134 343 138
rect 347 134 367 138
rect 371 134 423 138
rect 427 134 447 138
rect 451 134 479 138
rect 483 134 535 138
rect 539 134 551 138
rect 555 134 591 138
rect 595 134 647 138
rect 651 134 663 138
rect 667 134 703 138
rect 707 134 759 138
rect 763 134 775 138
rect 779 134 823 138
rect 827 134 887 138
rect 891 134 895 138
rect 899 134 951 138
rect 955 134 1015 138
rect 1019 134 1079 138
rect 1083 134 1135 138
rect 1139 134 1151 138
rect 1155 134 1215 138
rect 1219 134 1255 138
rect 1259 134 1271 138
rect 1275 134 1327 138
rect 1331 134 1351 138
rect 103 133 1351 134
rect 1357 133 1358 139
rect 1406 136 1407 140
rect 1411 136 1823 140
rect 1827 136 1828 140
rect 1406 135 1412 136
rect 1822 135 1828 136
rect 1338 89 1339 95
rect 1345 94 2611 95
rect 1345 90 1367 94
rect 1371 90 1415 94
rect 1419 90 1471 94
rect 1475 90 1527 94
rect 1531 90 1583 94
rect 1587 90 1647 94
rect 1651 90 1727 94
rect 1731 90 1807 94
rect 1811 90 1887 94
rect 1891 90 1959 94
rect 1963 90 2031 94
rect 2035 90 2095 94
rect 2099 90 2159 94
rect 2163 90 2223 94
rect 2227 90 2287 94
rect 2291 90 2359 94
rect 2363 90 2431 94
rect 2435 90 2583 94
rect 2587 90 2611 94
rect 1345 89 2611 90
rect 2617 89 2618 95
rect 84 77 85 83
rect 91 82 1339 83
rect 91 78 111 82
rect 115 78 159 82
rect 163 78 215 82
rect 219 78 271 82
rect 275 78 327 82
rect 331 78 383 82
rect 387 78 439 82
rect 443 78 495 82
rect 499 78 551 82
rect 555 78 607 82
rect 611 78 663 82
rect 667 78 719 82
rect 723 78 775 82
rect 779 78 839 82
rect 843 78 903 82
rect 907 78 967 82
rect 971 78 1031 82
rect 1035 78 1095 82
rect 1099 78 1167 82
rect 1171 78 1231 82
rect 1235 78 1287 82
rect 1291 78 1327 82
rect 1331 78 1339 82
rect 91 77 1339 78
rect 1345 77 1346 83
<< m5c >>
rect 85 2637 91 2643
rect 1339 2637 1345 2643
rect 97 2581 103 2587
rect 1351 2581 1357 2587
rect 85 2521 91 2527
rect 1339 2521 1345 2527
rect 1339 2513 1345 2519
rect 2611 2513 2617 2519
rect 97 2461 103 2467
rect 1351 2461 1357 2467
rect 85 2401 91 2407
rect 1339 2401 1345 2407
rect 97 2345 103 2351
rect 1351 2345 1357 2351
rect 85 2285 91 2291
rect 1339 2285 1345 2291
rect 1339 2277 1345 2283
rect 2611 2277 2617 2283
rect 97 2221 103 2227
rect 1351 2221 1357 2227
rect 1351 2209 1357 2215
rect 2623 2209 2629 2215
rect 85 2161 91 2167
rect 1339 2161 1345 2167
rect 1339 2153 1345 2159
rect 2611 2153 2617 2159
rect 97 2097 103 2103
rect 1351 2097 1357 2103
rect 1339 2041 1345 2047
rect 2611 2041 2617 2047
rect 85 2033 91 2039
rect 1339 2033 1345 2039
rect 1351 1985 1357 1991
rect 2623 1985 2629 1991
rect 97 1973 103 1979
rect 1351 1973 1357 1979
rect 1339 1925 1345 1931
rect 2611 1925 2617 1931
rect 85 1917 91 1923
rect 1339 1917 1345 1923
rect 1351 1865 1357 1871
rect 2623 1865 2629 1871
rect 97 1853 103 1859
rect 1351 1853 1357 1859
rect 1339 1809 1345 1815
rect 2611 1809 2617 1815
rect 85 1793 91 1799
rect 1339 1793 1345 1799
rect 1351 1753 1357 1759
rect 2623 1753 2629 1759
rect 97 1733 103 1739
rect 1351 1733 1357 1739
rect 1339 1685 1345 1691
rect 2611 1685 2617 1691
rect 85 1673 91 1679
rect 1339 1673 1345 1679
rect 1351 1617 1357 1623
rect 2623 1617 2629 1623
rect 97 1601 103 1607
rect 1351 1601 1357 1607
rect 1339 1557 1345 1563
rect 2611 1557 2617 1563
rect 85 1545 91 1551
rect 1339 1545 1345 1551
rect 1351 1493 1357 1499
rect 2623 1493 2629 1499
rect 97 1485 103 1491
rect 1351 1485 1357 1491
rect 85 1425 91 1431
rect 1339 1425 1345 1431
rect 97 1369 103 1375
rect 1351 1369 1357 1375
rect 85 1313 91 1319
rect 1339 1313 1345 1319
rect 1339 1305 1345 1311
rect 2611 1305 2617 1311
rect 97 1245 103 1251
rect 1351 1245 1357 1251
rect 85 1185 91 1191
rect 1339 1185 1345 1191
rect 97 1121 103 1127
rect 1351 1121 1357 1127
rect 85 1061 91 1067
rect 1339 1061 1345 1067
rect 97 1001 103 1007
rect 1351 1001 1357 1007
rect 1351 993 1357 999
rect 2623 993 2629 999
rect 85 941 91 947
rect 1339 941 1345 947
rect 1339 929 1345 935
rect 2611 929 2617 935
rect 97 885 103 891
rect 1351 885 1357 891
rect 1351 873 1357 879
rect 2623 873 2629 879
rect 85 821 91 827
rect 1339 821 1345 827
rect 1339 809 1345 815
rect 2611 809 2617 815
rect 97 757 103 763
rect 1351 757 1357 763
rect 1351 749 1357 755
rect 2623 749 2629 755
rect 85 697 91 703
rect 1339 697 1345 703
rect 1339 689 1345 695
rect 2611 689 2617 695
rect 97 633 103 639
rect 1351 633 1357 639
rect 85 573 91 579
rect 1339 573 1345 579
rect 97 509 103 515
rect 1351 509 1357 515
rect 85 449 91 455
rect 1339 449 1345 455
rect 97 389 103 395
rect 1351 389 1357 395
rect 85 329 91 335
rect 1339 329 1345 335
rect 97 269 103 275
rect 1351 269 1357 275
rect 85 213 91 219
rect 1339 213 1345 219
rect 1351 145 1357 151
rect 2623 145 2629 151
rect 97 133 103 139
rect 1351 133 1357 139
rect 1339 89 1345 95
rect 2611 89 2617 95
rect 85 77 91 83
rect 1339 77 1345 83
<< m5 >>
rect 84 2643 92 2664
rect 84 2637 85 2643
rect 91 2637 92 2643
rect 84 2527 92 2637
rect 84 2521 85 2527
rect 91 2521 92 2527
rect 84 2407 92 2521
rect 84 2401 85 2407
rect 91 2401 92 2407
rect 84 2291 92 2401
rect 84 2285 85 2291
rect 91 2285 92 2291
rect 84 2167 92 2285
rect 84 2161 85 2167
rect 91 2161 92 2167
rect 84 2039 92 2161
rect 84 2033 85 2039
rect 91 2033 92 2039
rect 84 1923 92 2033
rect 84 1917 85 1923
rect 91 1917 92 1923
rect 84 1799 92 1917
rect 84 1793 85 1799
rect 91 1793 92 1799
rect 84 1679 92 1793
rect 84 1673 85 1679
rect 91 1673 92 1679
rect 84 1551 92 1673
rect 84 1545 85 1551
rect 91 1545 92 1551
rect 84 1431 92 1545
rect 84 1425 85 1431
rect 91 1425 92 1431
rect 84 1319 92 1425
rect 84 1313 85 1319
rect 91 1313 92 1319
rect 84 1191 92 1313
rect 84 1185 85 1191
rect 91 1185 92 1191
rect 84 1067 92 1185
rect 84 1061 85 1067
rect 91 1061 92 1067
rect 84 947 92 1061
rect 84 941 85 947
rect 91 941 92 947
rect 84 827 92 941
rect 84 821 85 827
rect 91 821 92 827
rect 84 703 92 821
rect 84 697 85 703
rect 91 697 92 703
rect 84 579 92 697
rect 84 573 85 579
rect 91 573 92 579
rect 84 455 92 573
rect 84 449 85 455
rect 91 449 92 455
rect 84 335 92 449
rect 84 329 85 335
rect 91 329 92 335
rect 84 219 92 329
rect 84 213 85 219
rect 91 213 92 219
rect 84 83 92 213
rect 84 77 85 83
rect 91 77 92 83
rect 84 72 92 77
rect 96 2587 104 2664
rect 96 2581 97 2587
rect 103 2581 104 2587
rect 96 2467 104 2581
rect 96 2461 97 2467
rect 103 2461 104 2467
rect 96 2351 104 2461
rect 96 2345 97 2351
rect 103 2345 104 2351
rect 96 2227 104 2345
rect 96 2221 97 2227
rect 103 2221 104 2227
rect 96 2103 104 2221
rect 96 2097 97 2103
rect 103 2097 104 2103
rect 96 1979 104 2097
rect 96 1973 97 1979
rect 103 1973 104 1979
rect 96 1859 104 1973
rect 96 1853 97 1859
rect 103 1853 104 1859
rect 96 1739 104 1853
rect 96 1733 97 1739
rect 103 1733 104 1739
rect 96 1607 104 1733
rect 96 1601 97 1607
rect 103 1601 104 1607
rect 96 1491 104 1601
rect 96 1485 97 1491
rect 103 1485 104 1491
rect 96 1375 104 1485
rect 96 1369 97 1375
rect 103 1369 104 1375
rect 96 1251 104 1369
rect 96 1245 97 1251
rect 103 1245 104 1251
rect 96 1127 104 1245
rect 96 1121 97 1127
rect 103 1121 104 1127
rect 96 1007 104 1121
rect 96 1001 97 1007
rect 103 1001 104 1007
rect 96 891 104 1001
rect 96 885 97 891
rect 103 885 104 891
rect 96 763 104 885
rect 96 757 97 763
rect 103 757 104 763
rect 96 639 104 757
rect 96 633 97 639
rect 103 633 104 639
rect 96 515 104 633
rect 96 509 97 515
rect 103 509 104 515
rect 96 395 104 509
rect 96 389 97 395
rect 103 389 104 395
rect 96 275 104 389
rect 96 269 97 275
rect 103 269 104 275
rect 96 139 104 269
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1338 2643 1346 2664
rect 1338 2637 1339 2643
rect 1345 2637 1346 2643
rect 1338 2527 1346 2637
rect 1338 2521 1339 2527
rect 1345 2521 1346 2527
rect 1338 2519 1346 2521
rect 1338 2513 1339 2519
rect 1345 2513 1346 2519
rect 1338 2407 1346 2513
rect 1338 2401 1339 2407
rect 1345 2401 1346 2407
rect 1338 2291 1346 2401
rect 1338 2285 1339 2291
rect 1345 2285 1346 2291
rect 1338 2283 1346 2285
rect 1338 2277 1339 2283
rect 1345 2277 1346 2283
rect 1338 2167 1346 2277
rect 1338 2161 1339 2167
rect 1345 2161 1346 2167
rect 1338 2159 1346 2161
rect 1338 2153 1339 2159
rect 1345 2153 1346 2159
rect 1338 2047 1346 2153
rect 1338 2041 1339 2047
rect 1345 2041 1346 2047
rect 1338 2039 1346 2041
rect 1338 2033 1339 2039
rect 1345 2033 1346 2039
rect 1338 1931 1346 2033
rect 1338 1925 1339 1931
rect 1345 1925 1346 1931
rect 1338 1923 1346 1925
rect 1338 1917 1339 1923
rect 1345 1917 1346 1923
rect 1338 1815 1346 1917
rect 1338 1809 1339 1815
rect 1345 1809 1346 1815
rect 1338 1799 1346 1809
rect 1338 1793 1339 1799
rect 1345 1793 1346 1799
rect 1338 1691 1346 1793
rect 1338 1685 1339 1691
rect 1345 1685 1346 1691
rect 1338 1679 1346 1685
rect 1338 1673 1339 1679
rect 1345 1673 1346 1679
rect 1338 1563 1346 1673
rect 1338 1557 1339 1563
rect 1345 1557 1346 1563
rect 1338 1551 1346 1557
rect 1338 1545 1339 1551
rect 1345 1545 1346 1551
rect 1338 1431 1346 1545
rect 1338 1425 1339 1431
rect 1345 1425 1346 1431
rect 1338 1319 1346 1425
rect 1338 1313 1339 1319
rect 1345 1313 1346 1319
rect 1338 1311 1346 1313
rect 1338 1305 1339 1311
rect 1345 1305 1346 1311
rect 1338 1191 1346 1305
rect 1338 1185 1339 1191
rect 1345 1185 1346 1191
rect 1338 1067 1346 1185
rect 1338 1061 1339 1067
rect 1345 1061 1346 1067
rect 1338 947 1346 1061
rect 1338 941 1339 947
rect 1345 941 1346 947
rect 1338 935 1346 941
rect 1338 929 1339 935
rect 1345 929 1346 935
rect 1338 827 1346 929
rect 1338 821 1339 827
rect 1345 821 1346 827
rect 1338 815 1346 821
rect 1338 809 1339 815
rect 1345 809 1346 815
rect 1338 703 1346 809
rect 1338 697 1339 703
rect 1345 697 1346 703
rect 1338 695 1346 697
rect 1338 689 1339 695
rect 1345 689 1346 695
rect 1338 579 1346 689
rect 1338 573 1339 579
rect 1345 573 1346 579
rect 1338 455 1346 573
rect 1338 449 1339 455
rect 1345 449 1346 455
rect 1338 335 1346 449
rect 1338 329 1339 335
rect 1345 329 1346 335
rect 1338 219 1346 329
rect 1338 213 1339 219
rect 1345 213 1346 219
rect 1338 95 1346 213
rect 1338 89 1339 95
rect 1345 89 1346 95
rect 1338 83 1346 89
rect 1338 77 1339 83
rect 1345 77 1346 83
rect 1338 72 1346 77
rect 1350 2587 1358 2664
rect 1350 2581 1351 2587
rect 1357 2581 1358 2587
rect 1350 2467 1358 2581
rect 1350 2461 1351 2467
rect 1357 2461 1358 2467
rect 1350 2351 1358 2461
rect 1350 2345 1351 2351
rect 1357 2345 1358 2351
rect 1350 2227 1358 2345
rect 1350 2221 1351 2227
rect 1357 2221 1358 2227
rect 1350 2215 1358 2221
rect 1350 2209 1351 2215
rect 1357 2209 1358 2215
rect 1350 2103 1358 2209
rect 1350 2097 1351 2103
rect 1357 2097 1358 2103
rect 1350 1991 1358 2097
rect 1350 1985 1351 1991
rect 1357 1985 1358 1991
rect 1350 1979 1358 1985
rect 1350 1973 1351 1979
rect 1357 1973 1358 1979
rect 1350 1871 1358 1973
rect 1350 1865 1351 1871
rect 1357 1865 1358 1871
rect 1350 1859 1358 1865
rect 1350 1853 1351 1859
rect 1357 1853 1358 1859
rect 1350 1759 1358 1853
rect 1350 1753 1351 1759
rect 1357 1753 1358 1759
rect 1350 1739 1358 1753
rect 1350 1733 1351 1739
rect 1357 1733 1358 1739
rect 1350 1623 1358 1733
rect 1350 1617 1351 1623
rect 1357 1617 1358 1623
rect 1350 1607 1358 1617
rect 1350 1601 1351 1607
rect 1357 1601 1358 1607
rect 1350 1499 1358 1601
rect 1350 1493 1351 1499
rect 1357 1493 1358 1499
rect 1350 1491 1358 1493
rect 1350 1485 1351 1491
rect 1357 1485 1358 1491
rect 1350 1375 1358 1485
rect 1350 1369 1351 1375
rect 1357 1369 1358 1375
rect 1350 1251 1358 1369
rect 1350 1245 1351 1251
rect 1357 1245 1358 1251
rect 1350 1127 1358 1245
rect 1350 1121 1351 1127
rect 1357 1121 1358 1127
rect 1350 1007 1358 1121
rect 1350 1001 1351 1007
rect 1357 1001 1358 1007
rect 1350 999 1358 1001
rect 1350 993 1351 999
rect 1357 993 1358 999
rect 1350 891 1358 993
rect 1350 885 1351 891
rect 1357 885 1358 891
rect 1350 879 1358 885
rect 1350 873 1351 879
rect 1357 873 1358 879
rect 1350 763 1358 873
rect 1350 757 1351 763
rect 1357 757 1358 763
rect 1350 755 1358 757
rect 1350 749 1351 755
rect 1357 749 1358 755
rect 1350 639 1358 749
rect 1350 633 1351 639
rect 1357 633 1358 639
rect 1350 515 1358 633
rect 1350 509 1351 515
rect 1357 509 1358 515
rect 1350 395 1358 509
rect 1350 389 1351 395
rect 1357 389 1358 395
rect 1350 275 1358 389
rect 1350 269 1351 275
rect 1357 269 1358 275
rect 1350 151 1358 269
rect 1350 145 1351 151
rect 1357 145 1358 151
rect 1350 139 1358 145
rect 1350 133 1351 139
rect 1357 133 1358 139
rect 1350 72 1358 133
rect 2610 2519 2618 2664
rect 2610 2513 2611 2519
rect 2617 2513 2618 2519
rect 2610 2283 2618 2513
rect 2610 2277 2611 2283
rect 2617 2277 2618 2283
rect 2610 2159 2618 2277
rect 2610 2153 2611 2159
rect 2617 2153 2618 2159
rect 2610 2047 2618 2153
rect 2610 2041 2611 2047
rect 2617 2041 2618 2047
rect 2610 1931 2618 2041
rect 2610 1925 2611 1931
rect 2617 1925 2618 1931
rect 2610 1815 2618 1925
rect 2610 1809 2611 1815
rect 2617 1809 2618 1815
rect 2610 1691 2618 1809
rect 2610 1685 2611 1691
rect 2617 1685 2618 1691
rect 2610 1563 2618 1685
rect 2610 1557 2611 1563
rect 2617 1557 2618 1563
rect 2610 1311 2618 1557
rect 2610 1305 2611 1311
rect 2617 1305 2618 1311
rect 2610 935 2618 1305
rect 2610 929 2611 935
rect 2617 929 2618 935
rect 2610 815 2618 929
rect 2610 809 2611 815
rect 2617 809 2618 815
rect 2610 695 2618 809
rect 2610 689 2611 695
rect 2617 689 2618 695
rect 2610 95 2618 689
rect 2610 89 2611 95
rect 2617 89 2618 95
rect 2610 72 2618 89
rect 2622 2215 2630 2664
rect 2622 2209 2623 2215
rect 2629 2209 2630 2215
rect 2622 1991 2630 2209
rect 2622 1985 2623 1991
rect 2629 1985 2630 1991
rect 2622 1871 2630 1985
rect 2622 1865 2623 1871
rect 2629 1865 2630 1871
rect 2622 1759 2630 1865
rect 2622 1753 2623 1759
rect 2629 1753 2630 1759
rect 2622 1623 2630 1753
rect 2622 1617 2623 1623
rect 2629 1617 2630 1623
rect 2622 1499 2630 1617
rect 2622 1493 2623 1499
rect 2629 1493 2630 1499
rect 2622 999 2630 1493
rect 2622 993 2623 999
rect 2629 993 2630 999
rect 2622 879 2630 993
rect 2622 873 2623 879
rect 2629 873 2630 879
rect 2622 755 2630 873
rect 2622 749 2623 755
rect 2629 749 2630 755
rect 2622 151 2630 749
rect 2622 145 2623 151
rect 2629 145 2630 151
rect 2622 72 2630 145
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__167
timestamp 1731220403
transform 1 0 2576 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220403
transform 1 0 1360 0 -1 2620
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220403
transform 1 0 2576 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220403
transform 1 0 1360 0 1 2540
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220403
transform 1 0 2576 0 -1 2500
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220403
transform 1 0 1360 0 -1 2500
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220403
transform 1 0 2576 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220403
transform 1 0 1360 0 1 2420
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220403
transform 1 0 2576 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220403
transform 1 0 1360 0 -1 2384
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220403
transform 1 0 2576 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220403
transform 1 0 1360 0 1 2304
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220403
transform 1 0 2576 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220403
transform 1 0 1360 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220403
transform 1 0 2576 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220403
transform 1 0 1360 0 1 2172
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220403
transform 1 0 2576 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220403
transform 1 0 1360 0 -1 2140
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220403
transform 1 0 2576 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220403
transform 1 0 1360 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220403
transform 1 0 2576 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220403
transform 1 0 1360 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220403
transform 1 0 2576 0 1 1948
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220403
transform 1 0 1360 0 1 1948
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220403
transform 1 0 2576 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220403
transform 1 0 1360 0 -1 1912
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220403
transform 1 0 2576 0 1 1828
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220403
transform 1 0 1360 0 1 1828
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220403
transform 1 0 2576 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220403
transform 1 0 1360 0 -1 1796
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220403
transform 1 0 2576 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220403
transform 1 0 1360 0 1 1716
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220403
transform 1 0 2576 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220403
transform 1 0 1360 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220403
transform 1 0 2576 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220403
transform 1 0 1360 0 1 1580
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220403
transform 1 0 2576 0 -1 1544
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220403
transform 1 0 1360 0 -1 1544
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220403
transform 1 0 2576 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220403
transform 1 0 1360 0 1 1456
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220403
transform 1 0 2576 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220403
transform 1 0 1360 0 -1 1416
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220403
transform 1 0 2576 0 1 1328
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220403
transform 1 0 1360 0 1 1328
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220403
transform 1 0 2576 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220403
transform 1 0 1360 0 -1 1292
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220403
transform 1 0 2576 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220403
transform 1 0 1360 0 1 1212
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220403
transform 1 0 2576 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220403
transform 1 0 1360 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220403
transform 1 0 2576 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220403
transform 1 0 1360 0 1 1088
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220403
transform 1 0 2576 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220403
transform 1 0 1360 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220403
transform 1 0 2576 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220403
transform 1 0 1360 0 1 956
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220403
transform 1 0 2576 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220403
transform 1 0 1360 0 -1 916
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220403
transform 1 0 2576 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220403
transform 1 0 1360 0 1 836
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220403
transform 1 0 2576 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220403
transform 1 0 1360 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220403
transform 1 0 2576 0 1 712
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220403
transform 1 0 1360 0 1 712
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220403
transform 1 0 2576 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220403
transform 1 0 1360 0 -1 676
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220403
transform 1 0 2576 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220403
transform 1 0 1360 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220403
transform 1 0 2576 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220403
transform 1 0 1360 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220403
transform 1 0 2576 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220403
transform 1 0 1360 0 1 476
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220403
transform 1 0 2576 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220403
transform 1 0 1360 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220403
transform 1 0 2576 0 1 356
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220403
transform 1 0 1360 0 1 356
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220403
transform 1 0 2576 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220403
transform 1 0 1360 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220403
transform 1 0 2576 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220403
transform 1 0 1360 0 1 236
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220403
transform 1 0 2576 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220403
transform 1 0 1360 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220403
transform 1 0 2576 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220403
transform 1 0 1360 0 1 108
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220403
transform 1 0 1320 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220403
transform 1 0 104 0 -1 2624
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220403
transform 1 0 1320 0 1 2544
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220403
transform 1 0 104 0 1 2544
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220403
transform 1 0 1320 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220403
transform 1 0 104 0 -1 2508
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220403
transform 1 0 1320 0 1 2424
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220403
transform 1 0 104 0 1 2424
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220403
transform 1 0 1320 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220403
transform 1 0 104 0 -1 2388
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220403
transform 1 0 1320 0 1 2308
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220403
transform 1 0 104 0 1 2308
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220403
transform 1 0 1320 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220403
transform 1 0 104 0 -1 2272
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220403
transform 1 0 1320 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220403
transform 1 0 104 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220403
transform 1 0 1320 0 -1 2148
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220403
transform 1 0 104 0 -1 2148
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220403
transform 1 0 1320 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220403
transform 1 0 104 0 1 2060
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220403
transform 1 0 1320 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220403
transform 1 0 104 0 -1 2020
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220403
transform 1 0 1320 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220403
transform 1 0 104 0 1 1936
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220403
transform 1 0 1320 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220403
transform 1 0 104 0 -1 1904
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220403
transform 1 0 1320 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220403
transform 1 0 104 0 1 1816
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220403
transform 1 0 1320 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220403
transform 1 0 104 0 -1 1780
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220403
transform 1 0 1320 0 1 1696
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220403
transform 1 0 104 0 1 1696
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220403
transform 1 0 1320 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220403
transform 1 0 104 0 -1 1660
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220403
transform 1 0 1320 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220403
transform 1 0 104 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220403
transform 1 0 1320 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220403
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220403
transform 1 0 1320 0 1 1448
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220403
transform 1 0 104 0 1 1448
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220403
transform 1 0 1320 0 -1 1412
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220403
transform 1 0 104 0 -1 1412
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220403
transform 1 0 1320 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220403
transform 1 0 104 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220403
transform 1 0 1320 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220403
transform 1 0 104 0 -1 1300
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220403
transform 1 0 1320 0 1 1208
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220403
transform 1 0 104 0 1 1208
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220403
transform 1 0 1320 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220403
transform 1 0 104 0 -1 1172
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220403
transform 1 0 1320 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220403
transform 1 0 104 0 1 1084
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220403
transform 1 0 1320 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220403
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220403
transform 1 0 1320 0 1 964
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220403
transform 1 0 104 0 1 964
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220403
transform 1 0 1320 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220403
transform 1 0 104 0 -1 928
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220403
transform 1 0 1320 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220403
transform 1 0 104 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220403
transform 1 0 1320 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220403
transform 1 0 104 0 -1 808
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220403
transform 1 0 1320 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220403
transform 1 0 104 0 1 720
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220403
transform 1 0 1320 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220403
transform 1 0 104 0 -1 684
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220403
transform 1 0 1320 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220403
transform 1 0 104 0 1 596
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220403
transform 1 0 1320 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220403
transform 1 0 104 0 -1 560
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220403
transform 1 0 1320 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220403
transform 1 0 104 0 1 472
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220403
transform 1 0 1320 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220403
transform 1 0 104 0 -1 436
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220403
transform 1 0 1320 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220403
transform 1 0 104 0 1 352
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220403
transform 1 0 1320 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220403
transform 1 0 104 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220403
transform 1 0 1320 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220403
transform 1 0 104 0 1 232
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220403
transform 1 0 1320 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220403
transform 1 0 104 0 -1 200
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220403
transform 1 0 1320 0 1 96
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220403
transform 1 0 104 0 1 96
box 7 3 12 24
use _0_0std_0_0cells_0_0AND2X1  tst_5999_6
timestamp 1731220403
transform 1 0 2440 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5998_6
timestamp 1731220403
transform 1 0 2512 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5997_6
timestamp 1731220403
transform 1 0 2512 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5996_6
timestamp 1731220403
transform 1 0 2512 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5995_6
timestamp 1731220403
transform 1 0 2512 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5994_6
timestamp 1731220403
transform 1 0 2456 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5993_6
timestamp 1731220403
transform 1 0 2304 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5992_6
timestamp 1731220403
transform 1 0 2224 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5991_6
timestamp 1731220403
transform 1 0 2136 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5990_6
timestamp 1731220403
transform 1 0 2040 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5989_6
timestamp 1731220403
transform 1 0 1936 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5988_6
timestamp 1731220403
transform 1 0 2368 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5987_6
timestamp 1731220403
transform 1 0 2304 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5986_6
timestamp 1731220403
transform 1 0 2200 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5985_6
timestamp 1731220403
transform 1 0 2248 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5984_6
timestamp 1731220403
transform 1 0 2160 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5983_6
timestamp 1731220403
transform 1 0 2064 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5982_6
timestamp 1731220403
transform 1 0 1968 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5981_6
timestamp 1731220403
transform 1 0 2152 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5980_6
timestamp 1731220403
transform 1 0 2064 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5979_6
timestamp 1731220403
transform 1 0 1976 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5978_6
timestamp 1731220403
transform 1 0 1912 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5977_6
timestamp 1731220403
transform 1 0 2008 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5976_6
timestamp 1731220403
transform 1 0 2104 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5975_6
timestamp 1731220403
transform 1 0 2208 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5974_6
timestamp 1731220403
transform 1 0 2064 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5973_6
timestamp 1731220403
transform 1 0 1928 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5972_6
timestamp 1731220403
transform 1 0 1808 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5971_6
timestamp 1731220403
transform 1 0 1824 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5970_6
timestamp 1731220403
transform 1 0 1728 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5969_6
timestamp 1731220403
transform 1 0 1632 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5968_6
timestamp 1731220403
transform 1 0 1528 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5967_6
timestamp 1731220403
transform 1 0 1896 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5966_6
timestamp 1731220403
transform 1 0 1824 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5965_6
timestamp 1731220403
transform 1 0 1752 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5964_6
timestamp 1731220403
transform 1 0 1688 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5963_6
timestamp 1731220403
transform 1 0 1632 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5962_6
timestamp 1731220403
transform 1 0 1872 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5961_6
timestamp 1731220403
transform 1 0 1776 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5960_6
timestamp 1731220403
transform 1 0 1688 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5959_6
timestamp 1731220403
transform 1 0 1600 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5958_6
timestamp 1731220403
transform 1 0 1520 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5957_6
timestamp 1731220403
transform 1 0 1864 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5956_6
timestamp 1731220403
transform 1 0 1752 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5955_6
timestamp 1731220403
transform 1 0 1640 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5954_6
timestamp 1731220403
transform 1 0 1528 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5953_6
timestamp 1731220403
transform 1 0 1424 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5952_6
timestamp 1731220403
transform 1 0 1520 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5951_6
timestamp 1731220403
transform 1 0 1576 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5950_6
timestamp 1731220403
transform 1 0 1632 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5949_6
timestamp 1731220403
transform 1 0 1688 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5948_6
timestamp 1731220403
transform 1 0 1744 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5947_6
timestamp 1731220403
transform 1 0 1800 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5946_6
timestamp 1731220403
transform 1 0 1856 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5945_6
timestamp 1731220403
transform 1 0 1912 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5944_6
timestamp 1731220403
transform 1 0 1968 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5943_6
timestamp 1731220403
transform 1 0 2136 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5942_6
timestamp 1731220403
transform 1 0 2080 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5941_6
timestamp 1731220403
transform 1 0 2024 0 -1 2636
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5940_6
timestamp 1731220403
transform 1 0 1976 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5939_6
timestamp 1731220403
transform 1 0 2096 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5938_6
timestamp 1731220403
transform 1 0 2216 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5937_6
timestamp 1731220403
transform 1 0 2336 0 1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5936_6
timestamp 1731220403
transform 1 0 2264 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5935_6
timestamp 1731220403
transform 1 0 2368 0 -1 2516
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5934_6
timestamp 1731220403
transform 1 0 2344 0 1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5933_6
timestamp 1731220403
transform 1 0 2416 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5932_6
timestamp 1731220403
transform 1 0 2376 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5931_6
timestamp 1731220403
transform 1 0 2408 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5930_6
timestamp 1731220403
transform 1 0 2512 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5929_6
timestamp 1731220403
transform 1 0 2512 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5928_6
timestamp 1731220403
transform 1 0 2512 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5927_6
timestamp 1731220403
transform 1 0 2512 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5926_6
timestamp 1731220403
transform 1 0 2416 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5925_6
timestamp 1731220403
transform 1 0 2344 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5924_6
timestamp 1731220403
transform 1 0 2440 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5923_6
timestamp 1731220403
transform 1 0 2432 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5922_6
timestamp 1731220403
transform 1 0 2328 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5921_6
timestamp 1731220403
transform 1 0 2296 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5920_6
timestamp 1731220403
transform 1 0 2192 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5919_6
timestamp 1731220403
transform 1 0 2080 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5918_6
timestamp 1731220403
transform 1 0 2024 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5917_6
timestamp 1731220403
transform 1 0 2128 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5916_6
timestamp 1731220403
transform 1 0 2232 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5915_6
timestamp 1731220403
transform 1 0 2256 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5914_6
timestamp 1731220403
transform 1 0 2160 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5913_6
timestamp 1731220403
transform 1 0 2056 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5912_6
timestamp 1731220403
transform 1 0 1952 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5911_6
timestamp 1731220403
transform 1 0 2296 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5910_6
timestamp 1731220403
transform 1 0 2184 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5909_6
timestamp 1731220403
transform 1 0 2080 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5908_6
timestamp 1731220403
transform 1 0 1976 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5907_6
timestamp 1731220403
transform 1 0 1872 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5906_6
timestamp 1731220403
transform 1 0 2072 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5905_6
timestamp 1731220403
transform 1 0 1992 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5904_6
timestamp 1731220403
transform 1 0 1912 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5903_6
timestamp 1731220403
transform 1 0 1832 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5902_6
timestamp 1731220403
transform 1 0 1800 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5901_6
timestamp 1731220403
transform 1 0 1856 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5900_6
timestamp 1731220403
transform 1 0 1912 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5899_6
timestamp 1731220403
transform 1 0 1968 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5898_6
timestamp 1731220403
transform 1 0 2088 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5897_6
timestamp 1731220403
transform 1 0 2024 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5896_6
timestamp 1731220403
transform 1 0 1992 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5895_6
timestamp 1731220403
transform 1 0 1904 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5894_6
timestamp 1731220403
transform 1 0 1816 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5893_6
timestamp 1731220403
transform 1 0 2168 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5892_6
timestamp 1731220403
transform 1 0 2080 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5891_6
timestamp 1731220403
transform 1 0 2032 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5890_6
timestamp 1731220403
transform 1 0 1920 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5889_6
timestamp 1731220403
transform 1 0 2400 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5888_6
timestamp 1731220403
transform 1 0 2272 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5887_6
timestamp 1731220403
transform 1 0 2152 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5886_6
timestamp 1731220403
transform 1 0 2104 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5885_6
timestamp 1731220403
transform 1 0 2008 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5884_6
timestamp 1731220403
transform 1 0 2360 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5883_6
timestamp 1731220403
transform 1 0 2272 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5882_6
timestamp 1731220403
transform 1 0 2192 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5881_6
timestamp 1731220403
transform 1 0 2184 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5880_6
timestamp 1731220403
transform 1 0 2112 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5879_6
timestamp 1731220403
transform 1 0 2032 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5878_6
timestamp 1731220403
transform 1 0 2256 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5877_6
timestamp 1731220403
transform 1 0 2320 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5876_6
timestamp 1731220403
transform 1 0 2392 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5875_6
timestamp 1731220403
transform 1 0 2456 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5874_6
timestamp 1731220403
transform 1 0 2448 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5873_6
timestamp 1731220403
transform 1 0 2512 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5872_6
timestamp 1731220403
transform 1 0 2512 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5871_6
timestamp 1731220403
transform 1 0 2512 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5870_6
timestamp 1731220403
transform 1 0 2512 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5869_6
timestamp 1731220403
transform 1 0 2512 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5868_6
timestamp 1731220403
transform 1 0 2512 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5867_6
timestamp 1731220403
transform 1 0 2456 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5866_6
timestamp 1731220403
transform 1 0 2512 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5865_6
timestamp 1731220403
transform 1 0 2448 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5864_6
timestamp 1731220403
transform 1 0 2360 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5863_6
timestamp 1731220403
transform 1 0 2272 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5862_6
timestamp 1731220403
transform 1 0 2296 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5861_6
timestamp 1731220403
transform 1 0 2376 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5860_6
timestamp 1731220403
transform 1 0 2376 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5859_6
timestamp 1731220403
transform 1 0 2456 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5858_6
timestamp 1731220403
transform 1 0 2416 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5857_6
timestamp 1731220403
transform 1 0 2304 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5856_6
timestamp 1731220403
transform 1 0 2192 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5855_6
timestamp 1731220403
transform 1 0 2136 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5854_6
timestamp 1731220403
transform 1 0 2216 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5853_6
timestamp 1731220403
transform 1 0 2296 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5852_6
timestamp 1731220403
transform 1 0 2216 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5851_6
timestamp 1731220403
transform 1 0 2136 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5850_6
timestamp 1731220403
transform 1 0 2056 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5849_6
timestamp 1731220403
transform 1 0 1992 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5848_6
timestamp 1731220403
transform 1 0 2088 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5847_6
timestamp 1731220403
transform 1 0 2184 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5846_6
timestamp 1731220403
transform 1 0 2192 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5845_6
timestamp 1731220403
transform 1 0 2112 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5844_6
timestamp 1731220403
transform 1 0 2032 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5843_6
timestamp 1731220403
transform 1 0 1952 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5842_6
timestamp 1731220403
transform 1 0 1928 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5841_6
timestamp 1731220403
transform 1 0 2016 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5840_6
timestamp 1731220403
transform 1 0 2104 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5839_6
timestamp 1731220403
transform 1 0 2200 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5838_6
timestamp 1731220403
transform 1 0 2136 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5837_6
timestamp 1731220403
transform 1 0 2064 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5836_6
timestamp 1731220403
transform 1 0 2280 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5835_6
timestamp 1731220403
transform 1 0 2208 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5834_6
timestamp 1731220403
transform 1 0 2176 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5833_6
timestamp 1731220403
transform 1 0 2080 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5832_6
timestamp 1731220403
transform 1 0 2368 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5831_6
timestamp 1731220403
transform 1 0 2272 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5830_6
timestamp 1731220403
transform 1 0 2264 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5829_6
timestamp 1731220403
transform 1 0 2200 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5828_6
timestamp 1731220403
transform 1 0 2128 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5827_6
timestamp 1731220403
transform 1 0 2048 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5826_6
timestamp 1731220403
transform 1 0 2136 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5825_6
timestamp 1731220403
transform 1 0 2240 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5824_6
timestamp 1731220403
transform 1 0 2336 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5823_6
timestamp 1731220403
transform 1 0 2328 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5822_6
timestamp 1731220403
transform 1 0 2392 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5821_6
timestamp 1731220403
transform 1 0 2512 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5820_6
timestamp 1731220403
transform 1 0 2456 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5819_6
timestamp 1731220403
transform 1 0 2432 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5818_6
timestamp 1731220403
transform 1 0 2512 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5817_6
timestamp 1731220403
transform 1 0 2512 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5816_6
timestamp 1731220403
transform 1 0 2392 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5815_6
timestamp 1731220403
transform 1 0 2280 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5814_6
timestamp 1731220403
transform 1 0 2408 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5813_6
timestamp 1731220403
transform 1 0 2512 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5812_6
timestamp 1731220403
transform 1 0 2512 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5811_6
timestamp 1731220403
transform 1 0 2456 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5810_6
timestamp 1731220403
transform 1 0 2392 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5809_6
timestamp 1731220403
transform 1 0 2328 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5808_6
timestamp 1731220403
transform 1 0 2264 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5807_6
timestamp 1731220403
transform 1 0 2200 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5806_6
timestamp 1731220403
transform 1 0 2128 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5805_6
timestamp 1731220403
transform 1 0 2056 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5804_6
timestamp 1731220403
transform 1 0 2392 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5803_6
timestamp 1731220403
transform 1 0 2304 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5802_6
timestamp 1731220403
transform 1 0 2216 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5801_6
timestamp 1731220403
transform 1 0 2128 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5800_6
timestamp 1731220403
transform 1 0 2320 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5799_6
timestamp 1731220403
transform 1 0 2232 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5798_6
timestamp 1731220403
transform 1 0 2144 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5797_6
timestamp 1731220403
transform 1 0 2088 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5796_6
timestamp 1731220403
transform 1 0 2176 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5795_6
timestamp 1731220403
transform 1 0 2264 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5794_6
timestamp 1731220403
transform 1 0 2360 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5793_6
timestamp 1731220403
transform 1 0 2392 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5792_6
timestamp 1731220403
transform 1 0 2264 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5791_6
timestamp 1731220403
transform 1 0 2144 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5790_6
timestamp 1731220403
transform 1 0 2208 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5789_6
timestamp 1731220403
transform 1 0 2288 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5788_6
timestamp 1731220403
transform 1 0 2368 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5787_6
timestamp 1731220403
transform 1 0 2512 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5786_6
timestamp 1731220403
transform 1 0 2448 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5785_6
timestamp 1731220403
transform 1 0 2384 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5784_6
timestamp 1731220403
transform 1 0 2312 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5783_6
timestamp 1731220403
transform 1 0 2240 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5782_6
timestamp 1731220403
transform 1 0 2456 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5781_6
timestamp 1731220403
transform 1 0 2512 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5780_6
timestamp 1731220403
transform 1 0 2512 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5779_6
timestamp 1731220403
transform 1 0 2512 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5778_6
timestamp 1731220403
transform 1 0 2512 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5777_6
timestamp 1731220403
transform 1 0 2448 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5776_6
timestamp 1731220403
transform 1 0 2512 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5775_6
timestamp 1731220403
transform 1 0 2512 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5774_6
timestamp 1731220403
transform 1 0 2432 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5773_6
timestamp 1731220403
transform 1 0 2456 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5772_6
timestamp 1731220403
transform 1 0 2392 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5771_6
timestamp 1731220403
transform 1 0 2360 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5770_6
timestamp 1731220403
transform 1 0 2280 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5769_6
timestamp 1731220403
transform 1 0 2200 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5768_6
timestamp 1731220403
transform 1 0 2320 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5767_6
timestamp 1731220403
transform 1 0 2256 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5766_6
timestamp 1731220403
transform 1 0 2184 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5765_6
timestamp 1731220403
transform 1 0 2104 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5764_6
timestamp 1731220403
transform 1 0 2136 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5763_6
timestamp 1731220403
transform 1 0 2232 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5762_6
timestamp 1731220403
transform 1 0 2328 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5761_6
timestamp 1731220403
transform 1 0 2400 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5760_6
timestamp 1731220403
transform 1 0 2328 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5759_6
timestamp 1731220403
transform 1 0 2256 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5758_6
timestamp 1731220403
transform 1 0 2192 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5757_6
timestamp 1731220403
transform 1 0 2128 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5756_6
timestamp 1731220403
transform 1 0 2064 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5755_6
timestamp 1731220403
transform 1 0 2000 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5754_6
timestamp 1731220403
transform 1 0 1928 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5753_6
timestamp 1731220403
transform 1 0 1856 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5752_6
timestamp 1731220403
transform 1 0 1928 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5751_6
timestamp 1731220403
transform 1 0 2032 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5750_6
timestamp 1731220403
transform 1 0 2024 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5749_6
timestamp 1731220403
transform 1 0 1936 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5748_6
timestamp 1731220403
transform 1 0 2024 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5747_6
timestamp 1731220403
transform 1 0 2112 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5746_6
timestamp 1731220403
transform 1 0 2400 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5745_6
timestamp 1731220403
transform 1 0 2264 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5744_6
timestamp 1731220403
transform 1 0 2136 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5743_6
timestamp 1731220403
transform 1 0 2024 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5742_6
timestamp 1731220403
transform 1 0 1968 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5741_6
timestamp 1731220403
transform 1 0 2056 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5740_6
timestamp 1731220403
transform 1 0 2408 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5739_6
timestamp 1731220403
transform 1 0 2280 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5738_6
timestamp 1731220403
transform 1 0 2160 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5737_6
timestamp 1731220403
transform 1 0 2160 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5736_6
timestamp 1731220403
transform 1 0 2080 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5735_6
timestamp 1731220403
transform 1 0 2000 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5734_6
timestamp 1731220403
transform 1 0 2120 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5733_6
timestamp 1731220403
transform 1 0 2024 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5732_6
timestamp 1731220403
transform 1 0 1928 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5731_6
timestamp 1731220403
transform 1 0 1896 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5730_6
timestamp 1731220403
transform 1 0 2024 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5729_6
timestamp 1731220403
transform 1 0 1992 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5728_6
timestamp 1731220403
transform 1 0 1896 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5727_6
timestamp 1731220403
transform 1 0 1984 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5726_6
timestamp 1731220403
transform 1 0 2064 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5725_6
timestamp 1731220403
transform 1 0 2040 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5724_6
timestamp 1731220403
transform 1 0 1976 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5723_6
timestamp 1731220403
transform 1 0 1888 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5722_6
timestamp 1731220403
transform 1 0 1912 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5721_6
timestamp 1731220403
transform 1 0 2032 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5720_6
timestamp 1731220403
transform 1 0 2152 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5719_6
timestamp 1731220403
transform 1 0 2256 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5718_6
timestamp 1731220403
transform 1 0 2128 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5717_6
timestamp 1731220403
transform 1 0 2000 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5716_6
timestamp 1731220403
transform 1 0 1888 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5715_6
timestamp 1731220403
transform 1 0 1792 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5714_6
timestamp 1731220403
transform 1 0 1920 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5713_6
timestamp 1731220403
transform 1 0 2032 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5712_6
timestamp 1731220403
transform 1 0 1960 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5711_6
timestamp 1731220403
transform 1 0 1872 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5710_6
timestamp 1731220403
transform 1 0 1984 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5709_6
timestamp 1731220403
transform 1 0 2000 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5708_6
timestamp 1731220403
transform 1 0 1936 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5707_6
timestamp 1731220403
transform 1 0 1832 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5706_6
timestamp 1731220403
transform 1 0 1792 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5705_6
timestamp 1731220403
transform 1 0 1872 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5704_6
timestamp 1731220403
transform 1 0 1896 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5703_6
timestamp 1731220403
transform 1 0 1968 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5702_6
timestamp 1731220403
transform 1 0 2056 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5701_6
timestamp 1731220403
transform 1 0 2088 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5700_6
timestamp 1731220403
transform 1 0 1992 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5699_6
timestamp 1731220403
transform 1 0 1904 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5698_6
timestamp 1731220403
transform 1 0 1944 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5697_6
timestamp 1731220403
transform 1 0 1856 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5696_6
timestamp 1731220403
transform 1 0 1768 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5695_6
timestamp 1731220403
transform 1 0 1808 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5694_6
timestamp 1731220403
transform 1 0 1912 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5693_6
timestamp 1731220403
transform 1 0 1808 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5692_6
timestamp 1731220403
transform 1 0 1704 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5691_6
timestamp 1731220403
transform 1 0 1728 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5690_6
timestamp 1731220403
transform 1 0 1744 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5689_6
timestamp 1731220403
transform 1 0 1688 0 -1 1928
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5688_6
timestamp 1731220403
transform 1 0 1664 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5687_6
timestamp 1731220403
transform 1 0 1568 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5686_6
timestamp 1731220403
transform 1 0 1752 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5685_6
timestamp 1731220403
transform 1 0 1680 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5684_6
timestamp 1731220403
transform 1 0 1776 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5683_6
timestamp 1731220403
transform 1 0 1744 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5682_6
timestamp 1731220403
transform 1 0 1848 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5681_6
timestamp 1731220403
transform 1 0 1808 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5680_6
timestamp 1731220403
transform 1 0 1920 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5679_6
timestamp 1731220403
transform 1 0 1968 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5678_6
timestamp 1731220403
transform 1 0 1848 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5677_6
timestamp 1731220403
transform 1 0 1728 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5676_6
timestamp 1731220403
transform 1 0 1704 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5675_6
timestamp 1731220403
transform 1 0 1824 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5674_6
timestamp 1731220403
transform 1 0 1712 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5673_6
timestamp 1731220403
transform 1 0 1624 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5672_6
timestamp 1731220403
transform 1 0 1552 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5671_6
timestamp 1731220403
transform 1 0 1424 0 -1 2400
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5670_6
timestamp 1731220403
transform 1 0 1496 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5669_6
timestamp 1731220403
transform 1 0 1440 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5668_6
timestamp 1731220403
transform 1 0 1384 0 1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5667_6
timestamp 1731220403
transform 1 0 1256 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5666_6
timestamp 1731220403
transform 1 0 1384 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5665_6
timestamp 1731220403
transform 1 0 1464 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5664_6
timestamp 1731220403
transform 1 0 1584 0 -1 2280
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5663_6
timestamp 1731220403
transform 1 0 1616 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5662_6
timestamp 1731220403
transform 1 0 1520 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5661_6
timestamp 1731220403
transform 1 0 1440 0 1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5660_6
timestamp 1731220403
transform 1 0 1504 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5659_6
timestamp 1731220403
transform 1 0 1600 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5658_6
timestamp 1731220403
transform 1 0 1704 0 -1 2156
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5657_6
timestamp 1731220403
transform 1 0 1632 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5656_6
timestamp 1731220403
transform 1 0 1520 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5655_6
timestamp 1731220403
transform 1 0 1416 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5654_6
timestamp 1731220403
transform 1 0 1384 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5653_6
timestamp 1731220403
transform 1 0 1576 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5652_6
timestamp 1731220403
transform 1 0 1472 0 -1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5651_6
timestamp 1731220403
transform 1 0 1464 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5650_6
timestamp 1731220403
transform 1 0 1384 0 1 1932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5649_6
timestamp 1731220403
transform 1 0 1256 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5648_6
timestamp 1731220403
transform 1 0 1168 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5647_6
timestamp 1731220403
transform 1 0 1056 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5646_6
timestamp 1731220403
transform 1 0 1256 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5645_6
timestamp 1731220403
transform 1 0 1384 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5644_6
timestamp 1731220403
transform 1 0 1448 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5643_6
timestamp 1731220403
transform 1 0 1544 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5642_6
timestamp 1731220403
transform 1 0 1640 0 1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5641_6
timestamp 1731220403
transform 1 0 1592 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5640_6
timestamp 1731220403
transform 1 0 1480 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5639_6
timestamp 1731220403
transform 1 0 1384 0 -1 1812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5638_6
timestamp 1731220403
transform 1 0 1424 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5637_6
timestamp 1731220403
transform 1 0 1504 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5636_6
timestamp 1731220403
transform 1 0 1600 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5635_6
timestamp 1731220403
transform 1 0 1704 0 1 1700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5634_6
timestamp 1731220403
transform 1 0 1680 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5633_6
timestamp 1731220403
transform 1 0 1600 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5632_6
timestamp 1731220403
transform 1 0 1528 0 -1 1688
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5631_6
timestamp 1731220403
transform 1 0 1560 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5630_6
timestamp 1731220403
transform 1 0 1616 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5629_6
timestamp 1731220403
transform 1 0 1672 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5628_6
timestamp 1731220403
transform 1 0 1736 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5627_6
timestamp 1731220403
transform 1 0 1816 0 1 1564
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5626_6
timestamp 1731220403
transform 1 0 1976 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5625_6
timestamp 1731220403
transform 1 0 1896 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5624_6
timestamp 1731220403
transform 1 0 1824 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5623_6
timestamp 1731220403
transform 1 0 1760 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5622_6
timestamp 1731220403
transform 1 0 1704 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5621_6
timestamp 1731220403
transform 1 0 1648 0 -1 1560
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5620_6
timestamp 1731220403
transform 1 0 1880 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5619_6
timestamp 1731220403
transform 1 0 1792 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5618_6
timestamp 1731220403
transform 1 0 1712 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5617_6
timestamp 1731220403
transform 1 0 1632 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5616_6
timestamp 1731220403
transform 1 0 1560 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5615_6
timestamp 1731220403
transform 1 0 1504 0 1 1440
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5614_6
timestamp 1731220403
transform 1 0 1792 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5613_6
timestamp 1731220403
transform 1 0 1688 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5612_6
timestamp 1731220403
transform 1 0 1592 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5611_6
timestamp 1731220403
transform 1 0 1504 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5610_6
timestamp 1731220403
transform 1 0 1440 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5609_6
timestamp 1731220403
transform 1 0 1384 0 -1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5608_6
timestamp 1731220403
transform 1 0 1704 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5607_6
timestamp 1731220403
transform 1 0 1616 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5606_6
timestamp 1731220403
transform 1 0 1528 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5605_6
timestamp 1731220403
transform 1 0 1440 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5604_6
timestamp 1731220403
transform 1 0 1384 0 1 1312
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5603_6
timestamp 1731220403
transform 1 0 1256 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5602_6
timestamp 1731220403
transform 1 0 1200 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5601_6
timestamp 1731220403
transform 1 0 1120 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5600_6
timestamp 1731220403
transform 1 0 1040 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5599_6
timestamp 1731220403
transform 1 0 960 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5598_6
timestamp 1731220403
transform 1 0 880 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5597_6
timestamp 1731220403
transform 1 0 1256 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5596_6
timestamp 1731220403
transform 1 0 1168 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5595_6
timestamp 1731220403
transform 1 0 1056 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5594_6
timestamp 1731220403
transform 1 0 944 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5593_6
timestamp 1731220403
transform 1 0 960 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5592_6
timestamp 1731220403
transform 1 0 1072 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5591_6
timestamp 1731220403
transform 1 0 1184 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5590_6
timestamp 1731220403
transform 1 0 1120 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5589_6
timestamp 1731220403
transform 1 0 1024 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5588_6
timestamp 1731220403
transform 1 0 936 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5587_6
timestamp 1731220403
transform 1 0 848 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5586_6
timestamp 1731220403
transform 1 0 872 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5585_6
timestamp 1731220403
transform 1 0 944 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5584_6
timestamp 1731220403
transform 1 0 1024 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5583_6
timestamp 1731220403
transform 1 0 968 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5582_6
timestamp 1731220403
transform 1 0 888 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5581_6
timestamp 1731220403
transform 1 0 1048 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5580_6
timestamp 1731220403
transform 1 0 1136 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5579_6
timestamp 1731220403
transform 1 0 1104 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5578_6
timestamp 1731220403
transform 1 0 1016 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5577_6
timestamp 1731220403
transform 1 0 1256 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5576_6
timestamp 1731220403
transform 1 0 1192 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5575_6
timestamp 1731220403
transform 1 0 1192 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5574_6
timestamp 1731220403
transform 1 0 1096 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5573_6
timestamp 1731220403
transform 1 0 1000 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5572_6
timestamp 1731220403
transform 1 0 1088 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5571_6
timestamp 1731220403
transform 1 0 1000 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5570_6
timestamp 1731220403
transform 1 0 856 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5569_6
timestamp 1731220403
transform 1 0 776 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5568_6
timestamp 1731220403
transform 1 0 696 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5567_6
timestamp 1731220403
transform 1 0 608 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5566_6
timestamp 1731220403
transform 1 0 592 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5565_6
timestamp 1731220403
transform 1 0 760 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5564_6
timestamp 1731220403
transform 1 0 680 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5563_6
timestamp 1731220403
transform 1 0 624 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5562_6
timestamp 1731220403
transform 1 0 712 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5561_6
timestamp 1731220403
transform 1 0 808 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5560_6
timestamp 1731220403
transform 1 0 776 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5559_6
timestamp 1731220403
transform 1 0 696 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5558_6
timestamp 1731220403
transform 1 0 616 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5557_6
timestamp 1731220403
transform 1 0 544 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5556_6
timestamp 1731220403
transform 1 0 480 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5555_6
timestamp 1731220403
transform 1 0 424 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5554_6
timestamp 1731220403
transform 1 0 368 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5553_6
timestamp 1731220403
transform 1 0 536 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5552_6
timestamp 1731220403
transform 1 0 456 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5551_6
timestamp 1731220403
transform 1 0 392 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5550_6
timestamp 1731220403
transform 1 0 336 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5549_6
timestamp 1731220403
transform 1 0 504 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5548_6
timestamp 1731220403
transform 1 0 416 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5547_6
timestamp 1731220403
transform 1 0 336 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5546_6
timestamp 1731220403
transform 1 0 264 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5545_6
timestamp 1731220403
transform 1 0 200 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5544_6
timestamp 1731220403
transform 1 0 520 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5543_6
timestamp 1731220403
transform 1 0 424 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5542_6
timestamp 1731220403
transform 1 0 336 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5541_6
timestamp 1731220403
transform 1 0 248 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5540_6
timestamp 1731220403
transform 1 0 184 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5539_6
timestamp 1731220403
transform 1 0 128 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5538_6
timestamp 1731220403
transform 1 0 128 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5537_6
timestamp 1731220403
transform 1 0 200 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5536_6
timestamp 1731220403
transform 1 0 296 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5535_6
timestamp 1731220403
transform 1 0 400 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5534_6
timestamp 1731220403
transform 1 0 512 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5533_6
timestamp 1731220403
transform 1 0 432 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5532_6
timestamp 1731220403
transform 1 0 376 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5531_6
timestamp 1731220403
transform 1 0 320 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5530_6
timestamp 1731220403
transform 1 0 488 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5529_6
timestamp 1731220403
transform 1 0 552 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5528_6
timestamp 1731220403
transform 1 0 664 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5527_6
timestamp 1731220403
transform 1 0 608 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5526_6
timestamp 1731220403
transform 1 0 552 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5525_6
timestamp 1731220403
transform 1 0 496 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5524_6
timestamp 1731220403
transform 1 0 440 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5523_6
timestamp 1731220403
transform 1 0 384 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5522_6
timestamp 1731220403
transform 1 0 640 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5521_6
timestamp 1731220403
transform 1 0 552 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5520_6
timestamp 1731220403
transform 1 0 464 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5519_6
timestamp 1731220403
transform 1 0 384 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5518_6
timestamp 1731220403
transform 1 0 312 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5517_6
timestamp 1731220403
transform 1 0 248 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5516_6
timestamp 1731220403
transform 1 0 632 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5515_6
timestamp 1731220403
transform 1 0 512 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5514_6
timestamp 1731220403
transform 1 0 392 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5513_6
timestamp 1731220403
transform 1 0 280 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5512_6
timestamp 1731220403
transform 1 0 184 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5511_6
timestamp 1731220403
transform 1 0 128 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5510_6
timestamp 1731220403
transform 1 0 608 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5509_6
timestamp 1731220403
transform 1 0 480 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5508_6
timestamp 1731220403
transform 1 0 344 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5507_6
timestamp 1731220403
transform 1 0 216 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5506_6
timestamp 1731220403
transform 1 0 128 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5505_6
timestamp 1731220403
transform 1 0 128 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5504_6
timestamp 1731220403
transform 1 0 216 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5503_6
timestamp 1731220403
transform 1 0 608 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5502_6
timestamp 1731220403
transform 1 0 480 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5501_6
timestamp 1731220403
transform 1 0 344 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5500_6
timestamp 1731220403
transform 1 0 248 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5499_6
timestamp 1731220403
transform 1 0 144 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5498_6
timestamp 1731220403
transform 1 0 584 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5497_6
timestamp 1731220403
transform 1 0 472 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5496_6
timestamp 1731220403
transform 1 0 360 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5495_6
timestamp 1731220403
transform 1 0 304 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5494_6
timestamp 1731220403
transform 1 0 216 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5493_6
timestamp 1731220403
transform 1 0 600 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5492_6
timestamp 1731220403
transform 1 0 496 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5491_6
timestamp 1731220403
transform 1 0 400 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5490_6
timestamp 1731220403
transform 1 0 384 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5489_6
timestamp 1731220403
transform 1 0 320 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5488_6
timestamp 1731220403
transform 1 0 256 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5487_6
timestamp 1731220403
transform 1 0 456 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5486_6
timestamp 1731220403
transform 1 0 536 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5485_6
timestamp 1731220403
transform 1 0 616 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5484_6
timestamp 1731220403
transform 1 0 584 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5483_6
timestamp 1731220403
transform 1 0 520 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5482_6
timestamp 1731220403
transform 1 0 456 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5481_6
timestamp 1731220403
transform 1 0 392 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5480_6
timestamp 1731220403
transform 1 0 336 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5479_6
timestamp 1731220403
transform 1 0 312 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5478_6
timestamp 1731220403
transform 1 0 256 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5477_6
timestamp 1731220403
transform 1 0 200 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5476_6
timestamp 1731220403
transform 1 0 368 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5475_6
timestamp 1731220403
transform 1 0 424 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5474_6
timestamp 1731220403
transform 1 0 480 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5473_6
timestamp 1731220403
transform 1 0 592 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5472_6
timestamp 1731220403
transform 1 0 536 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5471_6
timestamp 1731220403
transform 1 0 520 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5470_6
timestamp 1731220403
transform 1 0 576 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5469_6
timestamp 1731220403
transform 1 0 632 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5468_6
timestamp 1731220403
transform 1 0 688 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5467_6
timestamp 1731220403
transform 1 0 744 0 -1 2640
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5466_6
timestamp 1731220403
transform 1 0 704 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5465_6
timestamp 1731220403
transform 1 0 648 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5464_6
timestamp 1731220403
transform 1 0 760 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5463_6
timestamp 1731220403
transform 1 0 816 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5462_6
timestamp 1731220403
transform 1 0 872 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5461_6
timestamp 1731220403
transform 1 0 928 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5460_6
timestamp 1731220403
transform 1 0 1096 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5459_6
timestamp 1731220403
transform 1 0 1040 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5458_6
timestamp 1731220403
transform 1 0 984 0 1 2528
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5457_6
timestamp 1731220403
transform 1 0 776 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5456_6
timestamp 1731220403
transform 1 0 712 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5455_6
timestamp 1731220403
transform 1 0 648 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5454_6
timestamp 1731220403
transform 1 0 840 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5453_6
timestamp 1731220403
transform 1 0 984 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5452_6
timestamp 1731220403
transform 1 0 912 0 -1 2524
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5451_6
timestamp 1731220403
transform 1 0 848 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5450_6
timestamp 1731220403
transform 1 0 768 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5449_6
timestamp 1731220403
transform 1 0 696 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5448_6
timestamp 1731220403
transform 1 0 1008 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5447_6
timestamp 1731220403
transform 1 0 928 0 1 2408
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5446_6
timestamp 1731220403
transform 1 0 888 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5445_6
timestamp 1731220403
transform 1 0 792 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5444_6
timestamp 1731220403
transform 1 0 696 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5443_6
timestamp 1731220403
transform 1 0 1080 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5442_6
timestamp 1731220403
transform 1 0 984 0 -1 2404
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5441_6
timestamp 1731220403
transform 1 0 896 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5440_6
timestamp 1731220403
transform 1 0 800 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5439_6
timestamp 1731220403
transform 1 0 696 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5438_6
timestamp 1731220403
transform 1 0 1184 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5437_6
timestamp 1731220403
transform 1 0 1088 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5436_6
timestamp 1731220403
transform 1 0 992 0 1 2292
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5435_6
timestamp 1731220403
transform 1 0 968 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5434_6
timestamp 1731220403
transform 1 0 856 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5433_6
timestamp 1731220403
transform 1 0 736 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5432_6
timestamp 1731220403
transform 1 0 1072 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5431_6
timestamp 1731220403
transform 1 0 1176 0 -1 2288
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5430_6
timestamp 1731220403
transform 1 0 1256 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5429_6
timestamp 1731220403
transform 1 0 1176 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5428_6
timestamp 1731220403
transform 1 0 1072 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5427_6
timestamp 1731220403
transform 1 0 968 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5426_6
timestamp 1731220403
transform 1 0 856 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5425_6
timestamp 1731220403
transform 1 0 736 0 1 2168
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5424_6
timestamp 1731220403
transform 1 0 1240 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5423_6
timestamp 1731220403
transform 1 0 1136 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5422_6
timestamp 1731220403
transform 1 0 1040 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5421_6
timestamp 1731220403
transform 1 0 944 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5420_6
timestamp 1731220403
transform 1 0 848 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5419_6
timestamp 1731220403
transform 1 0 744 0 -1 2164
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5418_6
timestamp 1731220403
transform 1 0 1112 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5417_6
timestamp 1731220403
transform 1 0 1032 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5416_6
timestamp 1731220403
transform 1 0 952 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5415_6
timestamp 1731220403
transform 1 0 872 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5414_6
timestamp 1731220403
transform 1 0 800 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5413_6
timestamp 1731220403
transform 1 0 720 0 1 2044
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5412_6
timestamp 1731220403
transform 1 0 1000 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5411_6
timestamp 1731220403
transform 1 0 944 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5410_6
timestamp 1731220403
transform 1 0 888 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5409_6
timestamp 1731220403
transform 1 0 832 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5408_6
timestamp 1731220403
transform 1 0 776 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5407_6
timestamp 1731220403
transform 1 0 720 0 -1 2036
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5406_6
timestamp 1731220403
transform 1 0 1128 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5405_6
timestamp 1731220403
transform 1 0 984 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5404_6
timestamp 1731220403
transform 1 0 848 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5403_6
timestamp 1731220403
transform 1 0 728 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5402_6
timestamp 1731220403
transform 1 0 632 0 1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5401_6
timestamp 1731220403
transform 1 0 624 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5400_6
timestamp 1731220403
transform 1 0 736 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5399_6
timestamp 1731220403
transform 1 0 848 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5398_6
timestamp 1731220403
transform 1 0 952 0 -1 1920
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5397_6
timestamp 1731220403
transform 1 0 1024 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5396_6
timestamp 1731220403
transform 1 0 936 0 1 1800
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5395_6
timestamp 1731220403
transform 1 0 920 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5394_6
timestamp 1731220403
transform 1 0 840 0 -1 1796
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5393_6
timestamp 1731220403
transform 1 0 904 0 1 1680
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5392_6
timestamp 1731220403
transform 1 0 936 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5391_6
timestamp 1731220403
transform 1 0 856 0 -1 1676
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5390_6
timestamp 1731220403
transform 1 0 808 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5389_6
timestamp 1731220403
transform 1 0 720 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5388_6
timestamp 1731220403
transform 1 0 656 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5387_6
timestamp 1731220403
transform 1 0 728 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5386_6
timestamp 1731220403
transform 1 0 800 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5385_6
timestamp 1731220403
transform 1 0 760 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5384_6
timestamp 1731220403
transform 1 0 664 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5383_6
timestamp 1731220403
transform 1 0 736 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5382_6
timestamp 1731220403
transform 1 0 848 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5381_6
timestamp 1731220403
transform 1 0 832 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5380_6
timestamp 1731220403
transform 1 0 720 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5379_6
timestamp 1731220403
transform 1 0 696 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5378_6
timestamp 1731220403
transform 1 0 600 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5377_6
timestamp 1731220403
transform 1 0 792 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5376_6
timestamp 1731220403
transform 1 0 728 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5375_6
timestamp 1731220403
transform 1 0 656 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5374_6
timestamp 1731220403
transform 1 0 584 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5373_6
timestamp 1731220403
transform 1 0 800 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5372_6
timestamp 1731220403
transform 1 0 880 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5371_6
timestamp 1731220403
transform 1 0 808 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5370_6
timestamp 1731220403
transform 1 0 736 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5369_6
timestamp 1731220403
transform 1 0 656 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5368_6
timestamp 1731220403
transform 1 0 880 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5367_6
timestamp 1731220403
transform 1 0 1032 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5366_6
timestamp 1731220403
transform 1 0 952 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5365_6
timestamp 1731220403
transform 1 0 896 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5364_6
timestamp 1731220403
transform 1 0 808 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5363_6
timestamp 1731220403
transform 1 0 712 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5362_6
timestamp 1731220403
transform 1 0 976 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5361_6
timestamp 1731220403
transform 1 0 1152 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5360_6
timestamp 1731220403
transform 1 0 1064 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5359_6
timestamp 1731220403
transform 1 0 1024 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5358_6
timestamp 1731220403
transform 1 0 944 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5357_6
timestamp 1731220403
transform 1 0 856 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5356_6
timestamp 1731220403
transform 1 0 1192 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5355_6
timestamp 1731220403
transform 1 0 1104 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5354_6
timestamp 1731220403
transform 1 0 896 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5353_6
timestamp 1731220403
transform 1 0 832 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5352_6
timestamp 1731220403
transform 1 0 768 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5351_6
timestamp 1731220403
transform 1 0 960 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5350_6
timestamp 1731220403
transform 1 0 1024 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5349_6
timestamp 1731220403
transform 1 0 1088 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5348_6
timestamp 1731220403
transform 1 0 1144 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5347_6
timestamp 1731220403
transform 1 0 1200 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5346_6
timestamp 1731220403
transform 1 0 1256 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5345_6
timestamp 1731220403
transform 1 0 1256 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5344_6
timestamp 1731220403
transform 1 0 1384 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5343_6
timestamp 1731220403
transform 1 0 1440 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5342_6
timestamp 1731220403
transform 1 0 1464 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5341_6
timestamp 1731220403
transform 1 0 1384 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5340_6
timestamp 1731220403
transform 1 0 1384 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5339_6
timestamp 1731220403
transform 1 0 1472 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5338_6
timestamp 1731220403
transform 1 0 1568 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5337_6
timestamp 1731220403
transform 1 0 1544 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5336_6
timestamp 1731220403
transform 1 0 1480 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5335_6
timestamp 1731220403
transform 1 0 1608 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5334_6
timestamp 1731220403
transform 1 0 1640 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5333_6
timestamp 1731220403
transform 1 0 1736 0 -1 1308
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5332_6
timestamp 1731220403
transform 1 0 1744 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5331_6
timestamp 1731220403
transform 1 0 1672 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5330_6
timestamp 1731220403
transform 1 0 1808 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5329_6
timestamp 1731220403
transform 1 0 1872 0 1 1196
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5328_6
timestamp 1731220403
transform 1 0 1880 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5327_6
timestamp 1731220403
transform 1 0 1776 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5326_6
timestamp 1731220403
transform 1 0 1672 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5325_6
timestamp 1731220403
transform 1 0 1568 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5324_6
timestamp 1731220403
transform 1 0 1672 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5323_6
timestamp 1731220403
transform 1 0 1776 0 1 1072
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5322_6
timestamp 1731220403
transform 1 0 1808 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5321_6
timestamp 1731220403
transform 1 0 1696 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5320_6
timestamp 1731220403
transform 1 0 1592 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5319_6
timestamp 1731220403
transform 1 0 1504 0 -1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5318_6
timestamp 1731220403
transform 1 0 1704 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5317_6
timestamp 1731220403
transform 1 0 1624 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5316_6
timestamp 1731220403
transform 1 0 1552 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5315_6
timestamp 1731220403
transform 1 0 1496 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5314_6
timestamp 1731220403
transform 1 0 1440 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5313_6
timestamp 1731220403
transform 1 0 1384 0 1 940
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5312_6
timestamp 1731220403
transform 1 0 1384 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5311_6
timestamp 1731220403
transform 1 0 1440 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5310_6
timestamp 1731220403
transform 1 0 1496 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5309_6
timestamp 1731220403
transform 1 0 1584 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5308_6
timestamp 1731220403
transform 1 0 1792 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5307_6
timestamp 1731220403
transform 1 0 1680 0 -1 932
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5306_6
timestamp 1731220403
transform 1 0 1624 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5305_6
timestamp 1731220403
transform 1 0 1536 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5304_6
timestamp 1731220403
transform 1 0 1456 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5303_6
timestamp 1731220403
transform 1 0 1712 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5302_6
timestamp 1731220403
transform 1 0 1800 0 1 820
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5301_6
timestamp 1731220403
transform 1 0 1720 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5300_6
timestamp 1731220403
transform 1 0 1656 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5299_6
timestamp 1731220403
transform 1 0 1600 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5298_6
timestamp 1731220403
transform 1 0 1792 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5297_6
timestamp 1731220403
transform 1 0 1872 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5296_6
timestamp 1731220403
transform 1 0 1960 0 -1 812
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5295_6
timestamp 1731220403
transform 1 0 1904 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5294_6
timestamp 1731220403
transform 1 0 1824 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5293_6
timestamp 1731220403
transform 1 0 1744 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5292_6
timestamp 1731220403
transform 1 0 1672 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5291_6
timestamp 1731220403
transform 1 0 1608 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5290_6
timestamp 1731220403
transform 1 0 1552 0 1 696
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5289_6
timestamp 1731220403
transform 1 0 1792 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5288_6
timestamp 1731220403
transform 1 0 1688 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5287_6
timestamp 1731220403
transform 1 0 1584 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5286_6
timestamp 1731220403
transform 1 0 1480 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5285_6
timestamp 1731220403
transform 1 0 1384 0 -1 692
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5284_6
timestamp 1731220403
transform 1 0 1768 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5283_6
timestamp 1731220403
transform 1 0 1632 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5282_6
timestamp 1731220403
transform 1 0 1256 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5281_6
timestamp 1731220403
transform 1 0 1176 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5280_6
timestamp 1731220403
transform 1 0 1072 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5279_6
timestamp 1731220403
transform 1 0 976 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5278_6
timestamp 1731220403
transform 1 0 1032 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5277_6
timestamp 1731220403
transform 1 0 1152 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5276_6
timestamp 1731220403
transform 1 0 1256 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5275_6
timestamp 1731220403
transform 1 0 1384 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5274_6
timestamp 1731220403
transform 1 0 1496 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5273_6
timestamp 1731220403
transform 1 0 1440 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5272_6
timestamp 1731220403
transform 1 0 1384 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5271_6
timestamp 1731220403
transform 1 0 1520 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5270_6
timestamp 1731220403
transform 1 0 1616 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5269_6
timestamp 1731220403
transform 1 0 1824 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5268_6
timestamp 1731220403
transform 1 0 1720 0 -1 572
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5267_6
timestamp 1731220403
transform 1 0 1656 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5266_6
timestamp 1731220403
transform 1 0 1584 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5265_6
timestamp 1731220403
transform 1 0 1520 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5264_6
timestamp 1731220403
transform 1 0 1912 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5263_6
timestamp 1731220403
transform 1 0 1824 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5262_6
timestamp 1731220403
transform 1 0 1736 0 1 460
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5261_6
timestamp 1731220403
transform 1 0 1728 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5260_6
timestamp 1731220403
transform 1 0 1672 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5259_6
timestamp 1731220403
transform 1 0 1616 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5258_6
timestamp 1731220403
transform 1 0 1784 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5257_6
timestamp 1731220403
transform 1 0 1840 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5256_6
timestamp 1731220403
transform 1 0 1896 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5255_6
timestamp 1731220403
transform 1 0 1936 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5254_6
timestamp 1731220403
transform 1 0 1864 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5253_6
timestamp 1731220403
transform 1 0 1808 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5252_6
timestamp 1731220403
transform 1 0 1752 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5251_6
timestamp 1731220403
transform 1 0 1696 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5250_6
timestamp 1731220403
transform 1 0 1640 0 1 340
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5249_6
timestamp 1731220403
transform 1 0 1936 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5248_6
timestamp 1731220403
transform 1 0 1856 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5247_6
timestamp 1731220403
transform 1 0 1776 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5246_6
timestamp 1731220403
transform 1 0 1712 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5245_6
timestamp 1731220403
transform 1 0 1656 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5244_6
timestamp 1731220403
transform 1 0 1600 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5243_6
timestamp 1731220403
transform 1 0 1848 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5242_6
timestamp 1731220403
transform 1 0 1760 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5241_6
timestamp 1731220403
transform 1 0 1672 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5240_6
timestamp 1731220403
transform 1 0 1592 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5239_6
timestamp 1731220403
transform 1 0 1520 0 1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5238_6
timestamp 1731220403
transform 1 0 1824 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5237_6
timestamp 1731220403
transform 1 0 1720 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5236_6
timestamp 1731220403
transform 1 0 1624 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5235_6
timestamp 1731220403
transform 1 0 1528 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5234_6
timestamp 1731220403
transform 1 0 1448 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5233_6
timestamp 1731220403
transform 1 0 1384 0 -1 220
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5232_6
timestamp 1731220403
transform 1 0 1776 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5231_6
timestamp 1731220403
transform 1 0 1696 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5230_6
timestamp 1731220403
transform 1 0 1616 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5229_6
timestamp 1731220403
transform 1 0 1552 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5228_6
timestamp 1731220403
transform 1 0 1496 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5227_6
timestamp 1731220403
transform 1 0 1440 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5226_6
timestamp 1731220403
transform 1 0 1384 0 1 92
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5225_6
timestamp 1731220403
transform 1 0 1256 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5224_6
timestamp 1731220403
transform 1 0 1200 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5223_6
timestamp 1731220403
transform 1 0 1136 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5222_6
timestamp 1731220403
transform 1 0 1240 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5221_6
timestamp 1731220403
transform 1 0 1240 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5220_6
timestamp 1731220403
transform 1 0 1128 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5219_6
timestamp 1731220403
transform 1 0 1184 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5218_6
timestamp 1731220403
transform 1 0 1080 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5217_6
timestamp 1731220403
transform 1 0 992 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5216_6
timestamp 1731220403
transform 1 0 912 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5215_6
timestamp 1731220403
transform 1 0 1072 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5214_6
timestamp 1731220403
transform 1 0 1160 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5213_6
timestamp 1731220403
transform 1 0 1248 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5212_6
timestamp 1731220403
transform 1 0 1208 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5211_6
timestamp 1731220403
transform 1 0 1128 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5210_6
timestamp 1731220403
transform 1 0 1056 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5209_6
timestamp 1731220403
transform 1 0 984 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5208_6
timestamp 1731220403
transform 1 0 912 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5207_6
timestamp 1731220403
transform 1 0 840 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5206_6
timestamp 1731220403
transform 1 0 1072 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5205_6
timestamp 1731220403
transform 1 0 992 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5204_6
timestamp 1731220403
transform 1 0 920 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5203_6
timestamp 1731220403
transform 1 0 848 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5202_6
timestamp 1731220403
transform 1 0 776 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5201_6
timestamp 1731220403
transform 1 0 704 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5200_6
timestamp 1731220403
transform 1 0 688 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5199_6
timestamp 1731220403
transform 1 0 800 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5198_6
timestamp 1731220403
transform 1 0 912 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5197_6
timestamp 1731220403
transform 1 0 872 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5196_6
timestamp 1731220403
transform 1 0 768 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5195_6
timestamp 1731220403
transform 1 0 664 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5194_6
timestamp 1731220403
transform 1 0 560 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5193_6
timestamp 1731220403
transform 1 0 592 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5192_6
timestamp 1731220403
transform 1 0 680 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5191_6
timestamp 1731220403
transform 1 0 760 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5190_6
timestamp 1731220403
transform 1 0 840 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5189_6
timestamp 1731220403
transform 1 0 920 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5188_6
timestamp 1731220403
transform 1 0 1008 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5187_6
timestamp 1731220403
transform 1 0 1160 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5186_6
timestamp 1731220403
transform 1 0 1064 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5185_6
timestamp 1731220403
transform 1 0 976 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5184_6
timestamp 1731220403
transform 1 0 888 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5183_6
timestamp 1731220403
transform 1 0 792 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5182_6
timestamp 1731220403
transform 1 0 688 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5181_6
timestamp 1731220403
transform 1 0 1064 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5180_6
timestamp 1731220403
transform 1 0 976 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5179_6
timestamp 1731220403
transform 1 0 888 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5178_6
timestamp 1731220403
transform 1 0 808 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5177_6
timestamp 1731220403
transform 1 0 728 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5176_6
timestamp 1731220403
transform 1 0 640 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5175_6
timestamp 1731220403
transform 1 0 904 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5174_6
timestamp 1731220403
transform 1 0 832 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5173_6
timestamp 1731220403
transform 1 0 760 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5172_6
timestamp 1731220403
transform 1 0 696 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5171_6
timestamp 1731220403
transform 1 0 632 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5170_6
timestamp 1731220403
transform 1 0 672 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5169_6
timestamp 1731220403
transform 1 0 784 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5168_6
timestamp 1731220403
transform 1 0 728 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5167_6
timestamp 1731220403
transform 1 0 704 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5166_6
timestamp 1731220403
transform 1 0 768 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5165_6
timestamp 1731220403
transform 1 0 672 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5164_6
timestamp 1731220403
transform 1 0 616 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5163_6
timestamp 1731220403
transform 1 0 568 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5162_6
timestamp 1731220403
transform 1 0 480 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5161_6
timestamp 1731220403
transform 1 0 424 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5160_6
timestamp 1731220403
transform 1 0 504 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5159_6
timestamp 1731220403
transform 1 0 504 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5158_6
timestamp 1731220403
transform 1 0 400 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5157_6
timestamp 1731220403
transform 1 0 496 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5156_6
timestamp 1731220403
transform 1 0 608 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5155_6
timestamp 1731220403
transform 1 0 632 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5154_6
timestamp 1731220403
transform 1 0 520 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5153_6
timestamp 1731220403
transform 1 0 416 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5152_6
timestamp 1731220403
transform 1 0 472 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5151_6
timestamp 1731220403
transform 1 0 568 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5150_6
timestamp 1731220403
transform 1 0 512 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5149_6
timestamp 1731220403
transform 1 0 440 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5148_6
timestamp 1731220403
transform 1 0 584 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5147_6
timestamp 1731220403
transform 1 0 632 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5146_6
timestamp 1731220403
transform 1 0 536 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5145_6
timestamp 1731220403
transform 1 0 440 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5144_6
timestamp 1731220403
transform 1 0 352 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5143_6
timestamp 1731220403
transform 1 0 272 0 1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5142_6
timestamp 1731220403
transform 1 0 248 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5141_6
timestamp 1731220403
transform 1 0 304 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5140_6
timestamp 1731220403
transform 1 0 368 0 -1 1548
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5139_6
timestamp 1731220403
transform 1 0 368 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5138_6
timestamp 1731220403
transform 1 0 272 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5137_6
timestamp 1731220403
transform 1 0 184 0 1 1432
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5136_6
timestamp 1731220403
transform 1 0 128 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5135_6
timestamp 1731220403
transform 1 0 216 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5134_6
timestamp 1731220403
transform 1 0 312 0 -1 1428
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5133_6
timestamp 1731220403
transform 1 0 384 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5132_6
timestamp 1731220403
transform 1 0 280 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5131_6
timestamp 1731220403
transform 1 0 192 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5130_6
timestamp 1731220403
transform 1 0 128 0 1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5129_6
timestamp 1731220403
transform 1 0 128 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5128_6
timestamp 1731220403
transform 1 0 200 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5127_6
timestamp 1731220403
transform 1 0 296 0 -1 1316
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5126_6
timestamp 1731220403
transform 1 0 264 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5125_6
timestamp 1731220403
transform 1 0 184 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5124_6
timestamp 1731220403
transform 1 0 128 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5123_6
timestamp 1731220403
transform 1 0 344 0 1 1192
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5122_6
timestamp 1731220403
transform 1 0 296 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5121_6
timestamp 1731220403
transform 1 0 208 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5120_6
timestamp 1731220403
transform 1 0 128 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5119_6
timestamp 1731220403
transform 1 0 392 0 -1 1188
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5118_6
timestamp 1731220403
transform 1 0 304 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5117_6
timestamp 1731220403
transform 1 0 208 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5116_6
timestamp 1731220403
transform 1 0 512 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5115_6
timestamp 1731220403
transform 1 0 408 0 1 1068
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5114_6
timestamp 1731220403
transform 1 0 408 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5113_6
timestamp 1731220403
transform 1 0 336 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5112_6
timestamp 1731220403
transform 1 0 280 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5111_6
timestamp 1731220403
transform 1 0 488 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5110_6
timestamp 1731220403
transform 1 0 576 0 -1 1064
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5109_6
timestamp 1731220403
transform 1 0 512 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5108_6
timestamp 1731220403
transform 1 0 456 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5107_6
timestamp 1731220403
transform 1 0 400 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5106_6
timestamp 1731220403
transform 1 0 576 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5105_6
timestamp 1731220403
transform 1 0 640 0 1 948
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5104_6
timestamp 1731220403
transform 1 0 616 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5103_6
timestamp 1731220403
transform 1 0 560 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5102_6
timestamp 1731220403
transform 1 0 504 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5101_6
timestamp 1731220403
transform 1 0 448 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_5100_6
timestamp 1731220403
transform 1 0 392 0 -1 944
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_599_6
timestamp 1731220403
transform 1 0 568 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_598_6
timestamp 1731220403
transform 1 0 504 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_597_6
timestamp 1731220403
transform 1 0 440 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_596_6
timestamp 1731220403
transform 1 0 376 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_595_6
timestamp 1731220403
transform 1 0 320 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_594_6
timestamp 1731220403
transform 1 0 264 0 1 832
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_593_6
timestamp 1731220403
transform 1 0 552 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_592_6
timestamp 1731220403
transform 1 0 456 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_591_6
timestamp 1731220403
transform 1 0 368 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_590_6
timestamp 1731220403
transform 1 0 280 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_589_6
timestamp 1731220403
transform 1 0 200 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_588_6
timestamp 1731220403
transform 1 0 136 0 -1 824
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_587_6
timestamp 1731220403
transform 1 0 584 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_586_6
timestamp 1731220403
transform 1 0 472 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_585_6
timestamp 1731220403
transform 1 0 368 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_584_6
timestamp 1731220403
transform 1 0 264 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_583_6
timestamp 1731220403
transform 1 0 184 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_582_6
timestamp 1731220403
transform 1 0 128 0 1 704
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_581_6
timestamp 1731220403
transform 1 0 328 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_580_6
timestamp 1731220403
transform 1 0 248 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_579_6
timestamp 1731220403
transform 1 0 184 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_578_6
timestamp 1731220403
transform 1 0 128 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_577_6
timestamp 1731220403
transform 1 0 504 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_576_6
timestamp 1731220403
transform 1 0 416 0 -1 700
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_575_6
timestamp 1731220403
transform 1 0 240 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_574_6
timestamp 1731220403
transform 1 0 184 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_573_6
timestamp 1731220403
transform 1 0 128 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_572_6
timestamp 1731220403
transform 1 0 296 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_571_6
timestamp 1731220403
transform 1 0 464 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_570_6
timestamp 1731220403
transform 1 0 376 0 1 580
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_569_6
timestamp 1731220403
transform 1 0 304 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_568_6
timestamp 1731220403
transform 1 0 232 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_567_6
timestamp 1731220403
transform 1 0 168 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_566_6
timestamp 1731220403
transform 1 0 384 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_565_6
timestamp 1731220403
transform 1 0 584 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_564_6
timestamp 1731220403
transform 1 0 480 0 -1 576
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_563_6
timestamp 1731220403
transform 1 0 408 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_562_6
timestamp 1731220403
transform 1 0 344 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_561_6
timestamp 1731220403
transform 1 0 288 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_560_6
timestamp 1731220403
transform 1 0 480 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_559_6
timestamp 1731220403
transform 1 0 632 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_558_6
timestamp 1731220403
transform 1 0 560 0 1 456
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_557_6
timestamp 1731220403
transform 1 0 544 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_556_6
timestamp 1731220403
transform 1 0 480 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_555_6
timestamp 1731220403
transform 1 0 424 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_554_6
timestamp 1731220403
transform 1 0 616 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_553_6
timestamp 1731220403
transform 1 0 696 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_552_6
timestamp 1731220403
transform 1 0 768 0 -1 452
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_551_6
timestamp 1731220403
transform 1 0 752 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_550_6
timestamp 1731220403
transform 1 0 832 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_549_6
timestamp 1731220403
transform 1 0 816 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_548_6
timestamp 1731220403
transform 1 0 736 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_547_6
timestamp 1731220403
transform 1 0 896 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_546_6
timestamp 1731220403
transform 1 0 984 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_545_6
timestamp 1731220403
transform 1 0 912 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_544_6
timestamp 1731220403
transform 1 0 808 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_543_6
timestamp 1731220403
transform 1 0 1016 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_542_6
timestamp 1731220403
transform 1 0 1000 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_541_6
timestamp 1731220403
transform 1 0 880 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_540_6
timestamp 1731220403
transform 1 0 1120 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_539_6
timestamp 1731220403
transform 1 0 1064 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_538_6
timestamp 1731220403
transform 1 0 1000 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_537_6
timestamp 1731220403
transform 1 0 936 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_536_6
timestamp 1731220403
transform 1 0 872 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_535_6
timestamp 1731220403
transform 1 0 808 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_534_6
timestamp 1731220403
transform 1 0 744 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_533_6
timestamp 1731220403
transform 1 0 688 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_532_6
timestamp 1731220403
transform 1 0 632 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_531_6
timestamp 1731220403
transform 1 0 648 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_530_6
timestamp 1731220403
transform 1 0 760 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_529_6
timestamp 1731220403
transform 1 0 704 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_528_6
timestamp 1731220403
transform 1 0 664 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_527_6
timestamp 1731220403
transform 1 0 600 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_526_6
timestamp 1731220403
transform 1 0 544 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_525_6
timestamp 1731220403
transform 1 0 672 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_524_6
timestamp 1731220403
transform 1 0 592 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_523_6
timestamp 1731220403
transform 1 0 520 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_522_6
timestamp 1731220403
transform 1 0 456 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_521_6
timestamp 1731220403
transform 1 0 400 0 1 336
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_520_6
timestamp 1731220403
transform 1 0 432 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_519_6
timestamp 1731220403
transform 1 0 488 0 -1 332
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_518_6
timestamp 1731220403
transform 1 0 608 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_517_6
timestamp 1731220403
transform 1 0 512 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_516_6
timestamp 1731220403
transform 1 0 424 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_515_6
timestamp 1731220403
transform 1 0 344 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_514_6
timestamp 1731220403
transform 1 0 272 0 1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_513_6
timestamp 1731220403
transform 1 0 536 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_512_6
timestamp 1731220403
transform 1 0 432 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_511_6
timestamp 1731220403
transform 1 0 328 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_510_6
timestamp 1731220403
transform 1 0 240 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_59_6
timestamp 1731220403
transform 1 0 168 0 -1 216
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_58_6
timestamp 1731220403
transform 1 0 576 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_57_6
timestamp 1731220403
transform 1 0 520 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_56_6
timestamp 1731220403
transform 1 0 464 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_55_6
timestamp 1731220403
transform 1 0 408 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_54_6
timestamp 1731220403
transform 1 0 352 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_53_6
timestamp 1731220403
transform 1 0 296 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_52_6
timestamp 1731220403
transform 1 0 240 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_51_6
timestamp 1731220403
transform 1 0 184 0 1 80
box 8 4 52 52
use _0_0std_0_0cells_0_0AND2X1  tst_50_6
timestamp 1731220403
transform 1 0 128 0 1 80
box 8 4 52 52
<< end >>
