magic
tech sky130l
timestamp 1731220663
<< m2c >>
rect 780 2567 784 2571
rect 836 2567 840 2571
rect 892 2567 896 2571
rect 948 2567 952 2571
rect 740 2553 744 2557
rect 796 2553 800 2557
rect 852 2553 856 2557
rect 908 2553 912 2557
rect 964 2551 968 2555
rect 1404 2545 1408 2549
rect 1460 2543 1464 2547
rect 1516 2543 1520 2547
rect 1572 2543 1576 2547
rect 1628 2543 1632 2547
rect 1684 2543 1688 2547
rect 1740 2543 1744 2547
rect 1796 2543 1800 2547
rect 1852 2543 1856 2547
rect 1908 2543 1912 2547
rect 1964 2543 1968 2547
rect 2020 2543 2024 2547
rect 2076 2543 2080 2547
rect 2132 2543 2136 2547
rect 2188 2543 2192 2547
rect 1420 2529 1424 2533
rect 1476 2529 1480 2533
rect 1532 2529 1536 2533
rect 1588 2529 1592 2533
rect 1644 2529 1648 2533
rect 1700 2529 1704 2533
rect 1756 2529 1760 2533
rect 1812 2529 1816 2533
rect 1868 2529 1872 2533
rect 1924 2529 1928 2533
rect 1980 2529 1984 2533
rect 2036 2529 2040 2533
rect 2092 2529 2096 2533
rect 2148 2529 2152 2533
rect 2204 2527 2208 2531
rect 204 2499 208 2503
rect 260 2499 264 2503
rect 316 2499 320 2503
rect 380 2499 384 2503
rect 444 2499 448 2503
rect 516 2499 520 2503
rect 596 2499 600 2503
rect 676 2499 680 2503
rect 756 2499 760 2503
rect 836 2499 840 2503
rect 916 2499 920 2503
rect 996 2499 1000 2503
rect 1076 2499 1080 2503
rect 188 2483 192 2487
rect 244 2485 248 2489
rect 300 2483 304 2487
rect 364 2485 368 2489
rect 428 2485 432 2489
rect 500 2483 504 2487
rect 580 2485 584 2489
rect 660 2483 664 2487
rect 740 2483 744 2487
rect 820 2485 824 2489
rect 900 2485 904 2489
rect 980 2485 984 2489
rect 1060 2485 1064 2489
rect 188 2465 192 2469
rect 252 2463 256 2467
rect 332 2463 336 2467
rect 420 2463 424 2467
rect 508 2465 512 2469
rect 604 2463 608 2467
rect 700 2463 704 2467
rect 796 2465 800 2469
rect 1388 2467 1392 2471
rect 1460 2467 1464 2471
rect 1548 2467 1552 2471
rect 1636 2467 1640 2471
rect 1724 2467 1728 2471
rect 1812 2467 1816 2471
rect 1900 2467 1904 2471
rect 1988 2467 1992 2471
rect 2076 2467 2080 2471
rect 2164 2467 2168 2471
rect 884 2463 888 2467
rect 972 2463 976 2467
rect 1068 2463 1072 2467
rect 1164 2463 1168 2467
rect 204 2447 208 2451
rect 268 2449 272 2453
rect 348 2449 352 2453
rect 436 2447 440 2451
rect 524 2449 528 2453
rect 620 2447 624 2451
rect 716 2447 720 2451
rect 812 2449 816 2453
rect 900 2449 904 2453
rect 988 2449 992 2453
rect 1084 2449 1088 2453
rect 1372 2451 1376 2455
rect 1444 2453 1448 2457
rect 1532 2453 1536 2457
rect 1620 2453 1624 2457
rect 1708 2453 1712 2457
rect 1796 2451 1800 2455
rect 1884 2453 1888 2457
rect 1972 2453 1976 2457
rect 2060 2453 2064 2457
rect 2148 2453 2152 2457
rect 1180 2447 1184 2451
rect 1372 2423 1376 2427
rect 1444 2423 1448 2427
rect 1548 2423 1552 2427
rect 1644 2423 1648 2427
rect 1740 2423 1744 2427
rect 1828 2423 1832 2427
rect 1916 2423 1920 2427
rect 2012 2423 2016 2427
rect 2108 2423 2112 2427
rect 1388 2409 1392 2413
rect 1460 2409 1464 2413
rect 1564 2409 1568 2413
rect 1660 2407 1664 2411
rect 1756 2407 1760 2411
rect 1844 2409 1848 2413
rect 1932 2409 1936 2413
rect 2028 2409 2032 2413
rect 2124 2409 2128 2413
rect 188 2391 192 2395
rect 268 2391 272 2395
rect 356 2391 360 2395
rect 452 2391 456 2395
rect 556 2391 560 2395
rect 660 2391 664 2395
rect 764 2391 768 2395
rect 868 2391 872 2395
rect 972 2391 976 2395
rect 1076 2391 1080 2395
rect 1188 2391 1192 2395
rect 172 2375 176 2379
rect 252 2377 256 2381
rect 340 2377 344 2381
rect 436 2377 440 2381
rect 540 2375 544 2379
rect 644 2377 648 2381
rect 748 2377 752 2381
rect 852 2375 856 2379
rect 956 2377 960 2381
rect 1060 2377 1064 2381
rect 1172 2377 1176 2381
rect 180 2357 184 2361
rect 284 2355 288 2359
rect 396 2355 400 2359
rect 508 2355 512 2359
rect 628 2355 632 2359
rect 748 2355 752 2359
rect 876 2357 880 2361
rect 1004 2355 1008 2359
rect 1132 2355 1136 2359
rect 1388 2347 1392 2351
rect 1444 2347 1448 2351
rect 1532 2347 1536 2351
rect 1620 2347 1624 2351
rect 1708 2347 1712 2351
rect 1788 2347 1792 2351
rect 1868 2347 1872 2351
rect 1956 2347 1960 2351
rect 2044 2347 2048 2351
rect 2132 2347 2136 2351
rect 196 2341 200 2345
rect 300 2341 304 2345
rect 412 2341 416 2345
rect 524 2339 528 2343
rect 644 2339 648 2343
rect 764 2341 768 2345
rect 892 2341 896 2345
rect 1020 2339 1024 2343
rect 1148 2339 1152 2343
rect 1372 2333 1376 2337
rect 1428 2333 1432 2337
rect 1516 2331 1520 2335
rect 1604 2331 1608 2335
rect 1692 2333 1696 2337
rect 1772 2331 1776 2335
rect 1852 2333 1856 2337
rect 1940 2333 1944 2337
rect 2028 2333 2032 2337
rect 2116 2333 2120 2337
rect 1372 2309 1376 2313
rect 1460 2307 1464 2311
rect 1548 2307 1552 2311
rect 1644 2307 1648 2311
rect 1740 2307 1744 2311
rect 1836 2309 1840 2313
rect 1932 2307 1936 2311
rect 2020 2307 2024 2311
rect 2116 2307 2120 2311
rect 2212 2307 2216 2311
rect 1388 2293 1392 2297
rect 1476 2293 1480 2297
rect 1564 2291 1568 2295
rect 1660 2291 1664 2295
rect 1756 2293 1760 2297
rect 1852 2293 1856 2297
rect 1948 2293 1952 2297
rect 2036 2293 2040 2297
rect 2132 2293 2136 2297
rect 2228 2291 2232 2295
rect 244 2283 248 2287
rect 324 2283 328 2287
rect 412 2283 416 2287
rect 508 2283 512 2287
rect 596 2283 600 2287
rect 684 2283 688 2287
rect 772 2283 776 2287
rect 852 2283 856 2287
rect 940 2283 944 2287
rect 1028 2283 1032 2287
rect 1116 2283 1120 2287
rect 228 2267 232 2271
rect 308 2269 312 2273
rect 396 2269 400 2273
rect 492 2269 496 2273
rect 580 2267 584 2271
rect 668 2269 672 2273
rect 756 2269 760 2273
rect 836 2267 840 2271
rect 924 2269 928 2273
rect 1012 2267 1016 2271
rect 1100 2269 1104 2273
rect 268 2245 272 2249
rect 324 2243 328 2247
rect 388 2243 392 2247
rect 452 2243 456 2247
rect 508 2243 512 2247
rect 564 2243 568 2247
rect 620 2243 624 2247
rect 676 2243 680 2247
rect 732 2243 736 2247
rect 796 2243 800 2247
rect 860 2243 864 2247
rect 924 2245 928 2249
rect 988 2243 992 2247
rect 1052 2243 1056 2247
rect 1116 2243 1120 2247
rect 1492 2239 1496 2243
rect 1580 2239 1584 2243
rect 1676 2239 1680 2243
rect 1772 2239 1776 2243
rect 1876 2239 1880 2243
rect 1972 2239 1976 2243
rect 2068 2239 2072 2243
rect 2156 2239 2160 2243
rect 2252 2239 2256 2243
rect 2348 2239 2352 2243
rect 284 2229 288 2233
rect 340 2229 344 2233
rect 404 2229 408 2233
rect 468 2229 472 2233
rect 524 2227 528 2231
rect 580 2227 584 2231
rect 636 2229 640 2233
rect 692 2229 696 2233
rect 748 2229 752 2233
rect 812 2229 816 2233
rect 876 2229 880 2233
rect 940 2229 944 2233
rect 1004 2229 1008 2233
rect 1068 2229 1072 2233
rect 1132 2227 1136 2231
rect 1476 2223 1480 2227
rect 1564 2225 1568 2229
rect 1660 2225 1664 2229
rect 1756 2225 1760 2229
rect 1860 2225 1864 2229
rect 1956 2223 1960 2227
rect 2052 2225 2056 2229
rect 2140 2225 2144 2229
rect 2236 2225 2240 2229
rect 2332 2225 2336 2229
rect 1572 2199 1576 2203
rect 1628 2199 1632 2203
rect 1684 2199 1688 2203
rect 1748 2201 1752 2205
rect 1812 2199 1816 2203
rect 1876 2199 1880 2203
rect 1932 2201 1936 2205
rect 1988 2199 1992 2203
rect 2044 2199 2048 2203
rect 2100 2199 2104 2203
rect 2164 2199 2168 2203
rect 2228 2199 2232 2203
rect 2292 2199 2296 2203
rect 2348 2199 2352 2203
rect 2404 2199 2408 2203
rect 2460 2199 2464 2203
rect 1588 2183 1592 2187
rect 1644 2185 1648 2189
rect 1700 2185 1704 2189
rect 1764 2185 1768 2189
rect 1828 2185 1832 2189
rect 1892 2183 1896 2187
rect 1948 2185 1952 2189
rect 2004 2185 2008 2189
rect 2060 2185 2064 2189
rect 2116 2185 2120 2189
rect 2180 2185 2184 2189
rect 2244 2185 2248 2189
rect 2308 2185 2312 2189
rect 2364 2185 2368 2189
rect 2420 2185 2424 2189
rect 2476 2183 2480 2187
rect 372 2171 376 2175
rect 428 2171 432 2175
rect 484 2171 488 2175
rect 540 2171 544 2175
rect 596 2171 600 2175
rect 356 2155 360 2159
rect 412 2157 416 2161
rect 468 2157 472 2161
rect 524 2157 528 2161
rect 580 2157 584 2161
rect 420 2137 424 2141
rect 516 2135 520 2139
rect 612 2135 616 2139
rect 716 2135 720 2139
rect 820 2135 824 2139
rect 932 2137 936 2141
rect 1044 2135 1048 2139
rect 1156 2135 1160 2139
rect 1244 2135 1248 2139
rect 436 2121 440 2125
rect 532 2121 536 2125
rect 628 2121 632 2125
rect 732 2121 736 2125
rect 836 2119 840 2123
rect 948 2121 952 2125
rect 1060 2121 1064 2125
rect 1172 2121 1176 2125
rect 1260 2119 1264 2123
rect 1700 2119 1704 2123
rect 1756 2119 1760 2123
rect 1828 2119 1832 2123
rect 1908 2119 1912 2123
rect 2004 2119 2008 2123
rect 2116 2119 2120 2123
rect 2236 2119 2240 2123
rect 2364 2119 2368 2123
rect 2476 2119 2480 2123
rect 1684 2103 1688 2107
rect 1740 2105 1744 2109
rect 1812 2105 1816 2109
rect 1892 2103 1896 2107
rect 1988 2105 1992 2109
rect 2100 2105 2104 2109
rect 2220 2103 2224 2107
rect 2348 2103 2352 2107
rect 2460 2105 2464 2109
rect 1372 2073 1376 2077
rect 412 2067 416 2071
rect 484 2067 488 2071
rect 556 2067 560 2071
rect 636 2067 640 2071
rect 716 2067 720 2071
rect 796 2067 800 2071
rect 868 2067 872 2071
rect 940 2067 944 2071
rect 1004 2067 1008 2071
rect 1068 2067 1072 2071
rect 1140 2067 1144 2071
rect 1204 2067 1208 2071
rect 1260 2069 1264 2073
rect 1428 2071 1432 2075
rect 1508 2071 1512 2075
rect 1596 2071 1600 2075
rect 1684 2071 1688 2075
rect 1788 2073 1792 2077
rect 1900 2071 1904 2075
rect 2028 2071 2032 2075
rect 2172 2071 2176 2075
rect 2324 2071 2328 2075
rect 2460 2071 2464 2075
rect 1388 2057 1392 2061
rect 1444 2057 1448 2061
rect 1524 2057 1528 2061
rect 1612 2057 1616 2061
rect 396 2051 400 2055
rect 468 2053 472 2057
rect 540 2051 544 2055
rect 620 2053 624 2057
rect 700 2053 704 2057
rect 780 2051 784 2055
rect 852 2053 856 2057
rect 924 2053 928 2057
rect 988 2053 992 2057
rect 1052 2053 1056 2057
rect 1124 2053 1128 2057
rect 1188 2051 1192 2055
rect 1244 2053 1248 2057
rect 1700 2055 1704 2059
rect 1804 2057 1808 2061
rect 1916 2057 1920 2061
rect 2044 2057 2048 2061
rect 2188 2057 2192 2061
rect 2340 2055 2344 2059
rect 2476 2055 2480 2059
rect 300 2029 304 2033
rect 380 2027 384 2031
rect 468 2027 472 2031
rect 556 2027 560 2031
rect 644 2027 648 2031
rect 724 2027 728 2031
rect 804 2027 808 2031
rect 892 2027 896 2031
rect 980 2027 984 2031
rect 1068 2027 1072 2031
rect 316 2013 320 2017
rect 396 2011 400 2015
rect 484 2013 488 2017
rect 572 2013 576 2017
rect 660 2011 664 2015
rect 740 2013 744 2017
rect 820 2013 824 2017
rect 908 2013 912 2017
rect 996 2013 1000 2017
rect 1084 2011 1088 2015
rect 1388 2003 1392 2007
rect 1460 2003 1464 2007
rect 1556 2003 1560 2007
rect 1652 2003 1656 2007
rect 1756 2003 1760 2007
rect 1860 2003 1864 2007
rect 1972 2003 1976 2007
rect 2092 2003 2096 2007
rect 2220 2003 2224 2007
rect 2356 2003 2360 2007
rect 2476 2003 2480 2007
rect 1372 1987 1376 1991
rect 1444 1989 1448 1993
rect 1540 1989 1544 1993
rect 1636 1989 1640 1993
rect 1740 1989 1744 1993
rect 1844 1987 1848 1991
rect 1956 1989 1960 1993
rect 2076 1987 2080 1991
rect 2204 1987 2208 1991
rect 2340 1989 2344 1993
rect 2460 1987 2464 1991
rect 1460 1965 1464 1969
rect 1548 1963 1552 1967
rect 1644 1963 1648 1967
rect 1740 1963 1744 1967
rect 1844 1963 1848 1967
rect 1948 1965 1952 1969
rect 2052 1963 2056 1967
rect 2156 1963 2160 1967
rect 2260 1963 2264 1967
rect 2372 1963 2376 1967
rect 2460 1963 2464 1967
rect 172 1955 176 1959
rect 244 1955 248 1959
rect 324 1955 328 1959
rect 420 1955 424 1959
rect 524 1955 528 1959
rect 628 1955 632 1959
rect 732 1955 736 1959
rect 836 1955 840 1959
rect 940 1955 944 1959
rect 1052 1955 1056 1959
rect 1476 1949 1480 1953
rect 1564 1949 1568 1953
rect 1660 1949 1664 1953
rect 1756 1949 1760 1953
rect 1860 1947 1864 1951
rect 1964 1949 1968 1953
rect 2068 1949 2072 1953
rect 2172 1947 2176 1951
rect 2276 1949 2280 1953
rect 2388 1949 2392 1953
rect 2476 1947 2480 1951
rect 156 1939 160 1943
rect 228 1941 232 1945
rect 308 1941 312 1945
rect 404 1939 408 1943
rect 508 1941 512 1945
rect 612 1941 616 1945
rect 716 1941 720 1945
rect 820 1939 824 1943
rect 924 1939 928 1943
rect 1036 1941 1040 1945
rect 156 1911 160 1915
rect 244 1913 248 1917
rect 380 1911 384 1915
rect 532 1911 536 1915
rect 692 1911 696 1915
rect 868 1911 872 1915
rect 1044 1911 1048 1915
rect 172 1895 176 1899
rect 260 1897 264 1901
rect 396 1897 400 1901
rect 548 1897 552 1901
rect 708 1895 712 1899
rect 884 1895 888 1899
rect 1060 1897 1064 1901
rect 1564 1891 1568 1895
rect 1652 1891 1656 1895
rect 1748 1891 1752 1895
rect 1852 1891 1856 1895
rect 1956 1891 1960 1895
rect 2052 1891 2056 1895
rect 2148 1891 2152 1895
rect 2236 1891 2240 1895
rect 2324 1891 2328 1895
rect 2412 1891 2416 1895
rect 2476 1891 2480 1895
rect 1548 1875 1552 1879
rect 1636 1877 1640 1881
rect 1732 1877 1736 1881
rect 1836 1877 1840 1881
rect 1940 1877 1944 1881
rect 2036 1875 2040 1879
rect 2132 1877 2136 1881
rect 2220 1877 2224 1881
rect 2308 1877 2312 1881
rect 2396 1875 2400 1879
rect 2460 1875 2464 1879
rect 1540 1857 1544 1861
rect 1612 1855 1616 1859
rect 1692 1855 1696 1859
rect 1788 1855 1792 1859
rect 1884 1855 1888 1859
rect 1988 1855 1992 1859
rect 2084 1855 2088 1859
rect 2180 1855 2184 1859
rect 2276 1855 2280 1859
rect 2372 1855 2376 1859
rect 2460 1855 2464 1859
rect 172 1843 176 1847
rect 228 1843 232 1847
rect 300 1843 304 1847
rect 372 1843 376 1847
rect 444 1843 448 1847
rect 516 1843 520 1847
rect 588 1843 592 1847
rect 652 1843 656 1847
rect 716 1843 720 1847
rect 780 1843 784 1847
rect 852 1843 856 1847
rect 924 1843 928 1847
rect 996 1843 1000 1847
rect 1076 1843 1080 1847
rect 1556 1841 1560 1845
rect 1628 1841 1632 1845
rect 1708 1839 1712 1843
rect 1804 1839 1808 1843
rect 1900 1841 1904 1845
rect 2004 1841 2008 1845
rect 2100 1841 2104 1845
rect 2196 1841 2200 1845
rect 2292 1841 2296 1845
rect 2388 1841 2392 1845
rect 2476 1839 2480 1843
rect 156 1827 160 1831
rect 212 1827 216 1831
rect 284 1829 288 1833
rect 356 1829 360 1833
rect 428 1827 432 1831
rect 500 1829 504 1833
rect 572 1829 576 1833
rect 636 1829 640 1833
rect 700 1829 704 1833
rect 764 1829 768 1833
rect 836 1829 840 1833
rect 908 1829 912 1833
rect 980 1829 984 1833
rect 1060 1827 1064 1831
rect 156 1799 160 1803
rect 236 1799 240 1803
rect 340 1799 344 1803
rect 444 1801 448 1805
rect 540 1799 544 1803
rect 636 1799 640 1803
rect 724 1801 728 1805
rect 804 1799 808 1803
rect 884 1799 888 1803
rect 964 1799 968 1803
rect 1044 1799 1048 1803
rect 1124 1799 1128 1803
rect 172 1785 176 1789
rect 252 1785 256 1789
rect 356 1783 360 1787
rect 460 1783 464 1787
rect 556 1785 560 1789
rect 652 1783 656 1787
rect 740 1785 744 1789
rect 820 1785 824 1789
rect 900 1785 904 1789
rect 980 1783 984 1787
rect 1060 1783 1064 1787
rect 1140 1785 1144 1789
rect 1500 1783 1504 1787
rect 1596 1783 1600 1787
rect 1700 1783 1704 1787
rect 1804 1783 1808 1787
rect 1916 1783 1920 1787
rect 2020 1783 2024 1787
rect 2124 1783 2128 1787
rect 2220 1783 2224 1787
rect 2308 1783 2312 1787
rect 2404 1783 2408 1787
rect 2476 1783 2480 1787
rect 1484 1769 1488 1773
rect 1580 1767 1584 1771
rect 1684 1767 1688 1771
rect 1788 1769 1792 1773
rect 1900 1769 1904 1773
rect 2004 1767 2008 1771
rect 2108 1769 2112 1773
rect 2204 1769 2208 1773
rect 2292 1769 2296 1773
rect 2388 1769 2392 1773
rect 2460 1767 2464 1771
rect 1380 1743 1384 1747
rect 1476 1745 1480 1749
rect 1572 1743 1576 1747
rect 1676 1743 1680 1747
rect 1780 1743 1784 1747
rect 1892 1745 1896 1749
rect 2004 1743 2008 1747
rect 2116 1743 2120 1747
rect 2236 1743 2240 1747
rect 2356 1743 2360 1747
rect 2460 1743 2464 1747
rect 172 1727 176 1731
rect 276 1727 280 1731
rect 388 1727 392 1731
rect 500 1727 504 1731
rect 612 1727 616 1731
rect 716 1727 720 1731
rect 820 1727 824 1731
rect 924 1727 928 1731
rect 1028 1727 1032 1731
rect 1140 1727 1144 1731
rect 1396 1727 1400 1731
rect 1492 1729 1496 1733
rect 1588 1729 1592 1733
rect 1692 1729 1696 1733
rect 1796 1727 1800 1731
rect 1908 1729 1912 1733
rect 2020 1729 2024 1733
rect 2132 1729 2136 1733
rect 2252 1729 2256 1733
rect 2372 1727 2376 1731
rect 2476 1727 2480 1731
rect 156 1713 160 1717
rect 260 1713 264 1717
rect 372 1711 376 1715
rect 484 1713 488 1717
rect 596 1711 600 1715
rect 700 1713 704 1717
rect 804 1711 808 1715
rect 908 1713 912 1717
rect 1012 1711 1016 1715
rect 1124 1711 1128 1715
rect 196 1687 200 1691
rect 276 1687 280 1691
rect 356 1687 360 1691
rect 444 1687 448 1691
rect 540 1687 544 1691
rect 644 1687 648 1691
rect 748 1687 752 1691
rect 852 1687 856 1691
rect 956 1687 960 1691
rect 1068 1687 1072 1691
rect 1180 1687 1184 1691
rect 212 1673 216 1677
rect 292 1673 296 1677
rect 372 1671 376 1675
rect 460 1673 464 1677
rect 556 1673 560 1677
rect 660 1671 664 1675
rect 764 1673 768 1677
rect 868 1673 872 1677
rect 972 1671 976 1675
rect 1084 1673 1088 1677
rect 1388 1675 1392 1679
rect 1468 1675 1472 1679
rect 1572 1675 1576 1679
rect 1684 1675 1688 1679
rect 1796 1675 1800 1679
rect 1916 1675 1920 1679
rect 2052 1675 2056 1679
rect 2196 1675 2200 1679
rect 2348 1675 2352 1679
rect 2476 1675 2480 1679
rect 1196 1671 1200 1675
rect 1372 1659 1376 1663
rect 1452 1659 1456 1663
rect 1556 1661 1560 1665
rect 1668 1661 1672 1665
rect 1780 1659 1784 1663
rect 1900 1661 1904 1665
rect 2036 1661 2040 1665
rect 2180 1661 2184 1665
rect 2332 1661 2336 1665
rect 2460 1659 2464 1663
rect 1372 1631 1376 1635
rect 1436 1631 1440 1635
rect 1524 1631 1528 1635
rect 1604 1633 1608 1637
rect 1684 1631 1688 1635
rect 1756 1631 1760 1635
rect 1844 1631 1848 1635
rect 1940 1631 1944 1635
rect 2060 1631 2064 1635
rect 2188 1631 2192 1635
rect 2332 1631 2336 1635
rect 2460 1631 2464 1635
rect 252 1619 256 1623
rect 308 1619 312 1623
rect 372 1619 376 1623
rect 444 1619 448 1623
rect 516 1619 520 1623
rect 596 1619 600 1623
rect 684 1619 688 1623
rect 780 1619 784 1623
rect 876 1619 880 1623
rect 980 1619 984 1623
rect 1092 1619 1096 1623
rect 1212 1619 1216 1623
rect 1388 1617 1392 1621
rect 1452 1617 1456 1621
rect 1540 1615 1544 1619
rect 1620 1617 1624 1621
rect 1700 1617 1704 1621
rect 1772 1617 1776 1621
rect 1860 1617 1864 1621
rect 1956 1617 1960 1621
rect 2076 1617 2080 1621
rect 2204 1617 2208 1621
rect 2348 1615 2352 1619
rect 2476 1615 2480 1619
rect 236 1603 240 1607
rect 292 1605 296 1609
rect 356 1603 360 1607
rect 428 1605 432 1609
rect 500 1605 504 1609
rect 580 1603 584 1607
rect 668 1603 672 1607
rect 764 1605 768 1609
rect 860 1605 864 1609
rect 964 1603 968 1607
rect 1076 1605 1080 1609
rect 1196 1603 1200 1607
rect 292 1583 296 1587
rect 356 1583 360 1587
rect 428 1583 432 1587
rect 508 1583 512 1587
rect 604 1583 608 1587
rect 708 1583 712 1587
rect 820 1583 824 1587
rect 940 1583 944 1587
rect 1068 1583 1072 1587
rect 1196 1583 1200 1587
rect 308 1569 312 1573
rect 372 1569 376 1573
rect 444 1569 448 1573
rect 524 1567 528 1571
rect 620 1569 624 1573
rect 724 1567 728 1571
rect 836 1569 840 1573
rect 956 1567 960 1571
rect 1084 1569 1088 1573
rect 1212 1567 1216 1571
rect 1388 1559 1392 1563
rect 1460 1559 1464 1563
rect 1564 1559 1568 1563
rect 1684 1559 1688 1563
rect 1820 1559 1824 1563
rect 1972 1559 1976 1563
rect 2140 1559 2144 1563
rect 2316 1559 2320 1563
rect 2476 1559 2480 1563
rect 1372 1545 1376 1549
rect 1444 1543 1448 1547
rect 1548 1543 1552 1547
rect 1668 1545 1672 1549
rect 1804 1545 1808 1549
rect 1956 1545 1960 1549
rect 2124 1545 2128 1549
rect 2300 1543 2304 1547
rect 2460 1543 2464 1547
rect 1372 1523 1376 1527
rect 1444 1523 1448 1527
rect 1548 1523 1552 1527
rect 1652 1523 1656 1527
rect 1756 1523 1760 1527
rect 1860 1523 1864 1527
rect 1964 1525 1968 1529
rect 2060 1523 2064 1527
rect 2156 1525 2160 1529
rect 2252 1523 2256 1527
rect 2348 1523 2352 1527
rect 2444 1523 2448 1527
rect 508 1507 512 1511
rect 588 1507 592 1511
rect 676 1507 680 1511
rect 772 1507 776 1511
rect 876 1507 880 1511
rect 988 1507 992 1511
rect 1100 1507 1104 1511
rect 1212 1507 1216 1511
rect 1388 1509 1392 1513
rect 1460 1509 1464 1513
rect 1564 1509 1568 1513
rect 1668 1509 1672 1513
rect 1772 1509 1776 1513
rect 1876 1507 1880 1511
rect 1980 1509 1984 1513
rect 2076 1507 2080 1511
rect 2172 1509 2176 1513
rect 2268 1507 2272 1511
rect 2364 1507 2368 1511
rect 2460 1507 2464 1511
rect 492 1491 496 1495
rect 572 1493 576 1497
rect 660 1493 664 1497
rect 756 1491 760 1495
rect 860 1493 864 1497
rect 972 1491 976 1495
rect 1084 1493 1088 1497
rect 1196 1491 1200 1495
rect 380 1473 384 1477
rect 468 1471 472 1475
rect 564 1471 568 1475
rect 660 1471 664 1475
rect 756 1471 760 1475
rect 860 1473 864 1477
rect 964 1471 968 1475
rect 1068 1471 1072 1475
rect 1172 1471 1176 1475
rect 396 1457 400 1461
rect 484 1457 488 1461
rect 580 1455 584 1459
rect 676 1457 680 1461
rect 772 1455 776 1459
rect 876 1457 880 1461
rect 980 1457 984 1461
rect 1084 1457 1088 1461
rect 1188 1455 1192 1459
rect 1388 1451 1392 1455
rect 1460 1451 1464 1455
rect 1556 1451 1560 1455
rect 1652 1451 1656 1455
rect 1748 1451 1752 1455
rect 1852 1451 1856 1455
rect 1964 1451 1968 1455
rect 2084 1451 2088 1455
rect 2212 1451 2216 1455
rect 2340 1451 2344 1455
rect 2476 1451 2480 1455
rect 1372 1437 1376 1441
rect 1444 1435 1448 1439
rect 1540 1435 1544 1439
rect 1636 1437 1640 1441
rect 1732 1435 1736 1439
rect 1836 1435 1840 1439
rect 1948 1437 1952 1441
rect 2068 1437 2072 1441
rect 2196 1435 2200 1439
rect 2324 1435 2328 1439
rect 2460 1435 2464 1439
rect 1372 1411 1376 1415
rect 1428 1411 1432 1415
rect 1508 1413 1512 1417
rect 1596 1411 1600 1415
rect 1684 1411 1688 1415
rect 1780 1413 1784 1417
rect 1884 1411 1888 1415
rect 1996 1411 2000 1415
rect 2116 1411 2120 1415
rect 2236 1411 2240 1415
rect 2356 1411 2360 1415
rect 2460 1411 2464 1415
rect 268 1403 272 1407
rect 356 1403 360 1407
rect 452 1403 456 1407
rect 548 1403 552 1407
rect 652 1403 656 1407
rect 748 1403 752 1407
rect 844 1403 848 1407
rect 932 1403 936 1407
rect 1028 1403 1032 1407
rect 1124 1403 1128 1407
rect 1388 1395 1392 1399
rect 1444 1397 1448 1401
rect 1524 1397 1528 1401
rect 1612 1397 1616 1401
rect 1700 1395 1704 1399
rect 1796 1397 1800 1401
rect 1900 1397 1904 1401
rect 2012 1397 2016 1401
rect 2132 1395 2136 1399
rect 2252 1395 2256 1399
rect 2372 1397 2376 1401
rect 2476 1395 2480 1399
rect 252 1387 256 1391
rect 340 1389 344 1393
rect 436 1389 440 1393
rect 532 1389 536 1393
rect 636 1387 640 1391
rect 732 1387 736 1391
rect 828 1389 832 1393
rect 916 1389 920 1393
rect 1012 1389 1016 1393
rect 1108 1389 1112 1393
rect 156 1367 160 1371
rect 220 1367 224 1371
rect 316 1367 320 1371
rect 412 1367 416 1371
rect 516 1367 520 1371
rect 612 1369 616 1373
rect 708 1367 712 1371
rect 804 1367 808 1371
rect 900 1367 904 1371
rect 1004 1367 1008 1371
rect 172 1351 176 1355
rect 236 1353 240 1357
rect 332 1353 336 1357
rect 428 1353 432 1357
rect 532 1353 536 1357
rect 628 1353 632 1357
rect 724 1353 728 1357
rect 820 1353 824 1357
rect 916 1353 920 1357
rect 1020 1351 1024 1355
rect 1388 1339 1392 1343
rect 1444 1339 1448 1343
rect 1516 1339 1520 1343
rect 1604 1339 1608 1343
rect 1692 1339 1696 1343
rect 1788 1339 1792 1343
rect 1892 1339 1896 1343
rect 2004 1339 2008 1343
rect 2116 1339 2120 1343
rect 2236 1339 2240 1343
rect 2364 1339 2368 1343
rect 2476 1339 2480 1343
rect 1372 1323 1376 1327
rect 1428 1325 1432 1329
rect 1500 1325 1504 1329
rect 1588 1325 1592 1329
rect 1676 1325 1680 1329
rect 1772 1323 1776 1327
rect 1876 1323 1880 1327
rect 1988 1325 1992 1329
rect 2100 1325 2104 1329
rect 2220 1325 2224 1329
rect 2348 1323 2352 1327
rect 2460 1323 2464 1327
rect 172 1299 176 1303
rect 252 1299 256 1303
rect 356 1299 360 1303
rect 452 1299 456 1303
rect 548 1299 552 1303
rect 636 1299 640 1303
rect 724 1299 728 1303
rect 820 1299 824 1303
rect 916 1299 920 1303
rect 1372 1295 1376 1299
rect 1428 1295 1432 1299
rect 1524 1295 1528 1299
rect 1620 1297 1624 1301
rect 1724 1295 1728 1299
rect 1828 1295 1832 1299
rect 1924 1297 1928 1301
rect 2020 1295 2024 1299
rect 2108 1295 2112 1299
rect 2188 1295 2192 1299
rect 2260 1295 2264 1299
rect 2332 1295 2336 1299
rect 2404 1297 2408 1301
rect 2460 1295 2464 1299
rect 156 1283 160 1287
rect 236 1285 240 1289
rect 340 1285 344 1289
rect 436 1285 440 1289
rect 532 1283 536 1287
rect 620 1285 624 1289
rect 708 1285 712 1289
rect 804 1285 808 1289
rect 900 1285 904 1289
rect 1388 1281 1392 1285
rect 1444 1281 1448 1285
rect 1540 1281 1544 1285
rect 1636 1281 1640 1285
rect 1740 1279 1744 1283
rect 1844 1279 1848 1283
rect 1940 1281 1944 1285
rect 2036 1281 2040 1285
rect 2124 1281 2128 1285
rect 2204 1281 2208 1285
rect 2276 1279 2280 1283
rect 2348 1279 2352 1283
rect 2420 1281 2424 1285
rect 2476 1279 2480 1283
rect 196 1265 200 1269
rect 252 1263 256 1267
rect 308 1263 312 1267
rect 372 1263 376 1267
rect 444 1263 448 1267
rect 532 1263 536 1267
rect 644 1263 648 1267
rect 780 1263 784 1267
rect 932 1263 936 1267
rect 1100 1263 1104 1267
rect 1244 1263 1248 1267
rect 212 1249 216 1253
rect 268 1249 272 1253
rect 324 1249 328 1253
rect 388 1249 392 1253
rect 460 1249 464 1253
rect 548 1247 552 1251
rect 660 1249 664 1253
rect 796 1249 800 1253
rect 948 1249 952 1253
rect 1116 1247 1120 1251
rect 1260 1247 1264 1251
rect 1388 1211 1392 1215
rect 1484 1211 1488 1215
rect 1612 1211 1616 1215
rect 1732 1211 1736 1215
rect 1852 1211 1856 1215
rect 1964 1211 1968 1215
rect 2068 1211 2072 1215
rect 2164 1211 2168 1215
rect 2252 1211 2256 1215
rect 2332 1211 2336 1215
rect 2412 1211 2416 1215
rect 2476 1211 2480 1215
rect 388 1195 392 1199
rect 444 1195 448 1199
rect 500 1195 504 1199
rect 556 1195 560 1199
rect 612 1195 616 1199
rect 668 1195 672 1199
rect 724 1195 728 1199
rect 780 1195 784 1199
rect 836 1195 840 1199
rect 892 1195 896 1199
rect 948 1195 952 1199
rect 1372 1197 1376 1201
rect 1468 1197 1472 1201
rect 1596 1195 1600 1199
rect 1716 1197 1720 1201
rect 1836 1197 1840 1201
rect 1948 1195 1952 1199
rect 2052 1197 2056 1201
rect 2148 1197 2152 1201
rect 2236 1197 2240 1201
rect 2316 1197 2320 1201
rect 2396 1195 2400 1199
rect 2460 1195 2464 1199
rect 372 1179 376 1183
rect 428 1181 432 1185
rect 484 1181 488 1185
rect 540 1181 544 1185
rect 596 1181 600 1185
rect 652 1181 656 1185
rect 708 1179 712 1183
rect 764 1181 768 1185
rect 820 1179 824 1183
rect 876 1181 880 1185
rect 932 1179 936 1183
rect 1372 1177 1376 1181
rect 1476 1175 1480 1179
rect 1604 1175 1608 1179
rect 1740 1175 1744 1179
rect 1868 1175 1872 1179
rect 1988 1177 1992 1181
rect 2092 1175 2096 1179
rect 2196 1175 2200 1179
rect 2292 1175 2296 1179
rect 2388 1175 2392 1179
rect 2460 1175 2464 1179
rect 1388 1161 1392 1165
rect 1492 1161 1496 1165
rect 428 1157 432 1161
rect 484 1155 488 1159
rect 540 1155 544 1159
rect 596 1157 600 1161
rect 652 1155 656 1159
rect 708 1155 712 1159
rect 764 1157 768 1161
rect 1620 1159 1624 1163
rect 1756 1159 1760 1163
rect 1884 1161 1888 1165
rect 2004 1161 2008 1165
rect 2108 1159 2112 1163
rect 2212 1159 2216 1163
rect 2308 1161 2312 1165
rect 2404 1161 2408 1165
rect 2476 1161 2480 1165
rect 820 1155 824 1159
rect 876 1155 880 1159
rect 932 1155 936 1159
rect 988 1155 992 1159
rect 444 1141 448 1145
rect 500 1141 504 1145
rect 556 1139 560 1143
rect 612 1141 616 1145
rect 668 1141 672 1145
rect 724 1139 728 1143
rect 780 1141 784 1145
rect 836 1141 840 1145
rect 892 1139 896 1143
rect 948 1141 952 1145
rect 1004 1139 1008 1143
rect 1404 1103 1408 1107
rect 1484 1103 1488 1107
rect 1572 1103 1576 1107
rect 1668 1103 1672 1107
rect 1756 1103 1760 1107
rect 1844 1103 1848 1107
rect 1932 1103 1936 1107
rect 2020 1103 2024 1107
rect 2108 1103 2112 1107
rect 2196 1103 2200 1107
rect 2292 1103 2296 1107
rect 2396 1103 2400 1107
rect 2476 1103 2480 1107
rect 1388 1087 1392 1091
rect 1468 1089 1472 1093
rect 1556 1087 1560 1091
rect 1652 1087 1656 1091
rect 1740 1089 1744 1093
rect 1828 1089 1832 1093
rect 1916 1087 1920 1091
rect 2004 1089 2008 1093
rect 2092 1089 2096 1093
rect 2180 1087 2184 1091
rect 2276 1089 2280 1093
rect 2380 1089 2384 1093
rect 2460 1087 2464 1091
rect 260 1083 264 1087
rect 348 1083 352 1087
rect 436 1083 440 1087
rect 532 1083 536 1087
rect 628 1083 632 1087
rect 716 1083 720 1087
rect 804 1083 808 1087
rect 884 1083 888 1087
rect 964 1083 968 1087
rect 1052 1083 1056 1087
rect 1140 1083 1144 1087
rect 244 1067 248 1071
rect 332 1069 336 1073
rect 420 1069 424 1073
rect 516 1069 520 1073
rect 612 1067 616 1071
rect 700 1067 704 1071
rect 788 1069 792 1073
rect 868 1069 872 1073
rect 948 1067 952 1071
rect 1036 1067 1040 1071
rect 1124 1069 1128 1073
rect 1436 1059 1440 1063
rect 1500 1059 1504 1063
rect 1572 1059 1576 1063
rect 1644 1059 1648 1063
rect 1708 1059 1712 1063
rect 1772 1059 1776 1063
rect 1844 1061 1848 1065
rect 1924 1059 1928 1063
rect 2012 1059 2016 1063
rect 2116 1059 2120 1063
rect 2236 1059 2240 1063
rect 2356 1059 2360 1063
rect 2460 1059 2464 1063
rect 156 1045 160 1049
rect 212 1043 216 1047
rect 308 1043 312 1047
rect 420 1043 424 1047
rect 540 1043 544 1047
rect 660 1043 664 1047
rect 772 1043 776 1047
rect 884 1043 888 1047
rect 988 1043 992 1047
rect 1100 1045 1104 1049
rect 1212 1043 1216 1047
rect 1452 1045 1456 1049
rect 1516 1045 1520 1049
rect 1588 1045 1592 1049
rect 1660 1043 1664 1047
rect 1724 1045 1728 1049
rect 1788 1043 1792 1047
rect 1860 1045 1864 1049
rect 1940 1045 1944 1049
rect 2028 1043 2032 1047
rect 2132 1045 2136 1049
rect 2252 1045 2256 1049
rect 2372 1043 2376 1047
rect 2476 1043 2480 1047
rect 172 1029 176 1033
rect 228 1029 232 1033
rect 324 1027 328 1031
rect 436 1029 440 1033
rect 556 1029 560 1033
rect 676 1027 680 1031
rect 788 1029 792 1033
rect 900 1029 904 1033
rect 1004 1027 1008 1031
rect 1116 1029 1120 1033
rect 1228 1027 1232 1031
rect 1548 983 1552 987
rect 1604 983 1608 987
rect 1660 983 1664 987
rect 1716 983 1720 987
rect 1772 983 1776 987
rect 1844 983 1848 987
rect 1924 983 1928 987
rect 2020 983 2024 987
rect 2132 983 2136 987
rect 2252 983 2256 987
rect 2372 983 2376 987
rect 2476 983 2480 987
rect 172 971 176 975
rect 252 971 256 975
rect 364 971 368 975
rect 476 971 480 975
rect 588 971 592 975
rect 700 971 704 975
rect 796 971 800 975
rect 884 971 888 975
rect 972 971 976 975
rect 1052 971 1056 975
rect 1124 971 1128 975
rect 1204 971 1208 975
rect 1260 971 1264 975
rect 1532 967 1536 971
rect 1588 969 1592 973
rect 1644 967 1648 971
rect 1700 967 1704 971
rect 1756 969 1760 973
rect 1828 969 1832 973
rect 1908 967 1912 971
rect 2004 969 2008 973
rect 2116 969 2120 973
rect 2236 969 2240 973
rect 2356 967 2360 971
rect 2460 967 2464 971
rect 156 957 160 961
rect 236 955 240 959
rect 348 955 352 959
rect 460 957 464 961
rect 572 957 576 961
rect 684 955 688 959
rect 780 957 784 961
rect 868 955 872 959
rect 956 955 960 959
rect 1036 957 1040 961
rect 1108 955 1112 959
rect 1188 955 1192 959
rect 1244 957 1248 961
rect 156 935 160 939
rect 212 935 216 939
rect 300 935 304 939
rect 404 935 408 939
rect 516 935 520 939
rect 628 935 632 939
rect 740 937 744 941
rect 836 935 840 939
rect 932 935 936 939
rect 1020 935 1024 939
rect 1100 935 1104 939
rect 1180 935 1184 939
rect 1244 935 1248 939
rect 1372 933 1376 937
rect 1444 933 1448 937
rect 1532 931 1536 935
rect 1620 931 1624 935
rect 1700 931 1704 935
rect 1796 931 1800 935
rect 1900 931 1904 935
rect 2020 931 2024 935
rect 2156 931 2160 935
rect 2300 931 2304 935
rect 2444 931 2448 935
rect 172 921 176 925
rect 228 921 232 925
rect 316 921 320 925
rect 420 921 424 925
rect 532 919 536 923
rect 644 921 648 925
rect 756 921 760 925
rect 852 919 856 923
rect 948 921 952 925
rect 1036 921 1040 925
rect 1116 919 1120 923
rect 1196 919 1200 923
rect 1260 919 1264 923
rect 1388 917 1392 921
rect 1460 917 1464 921
rect 1548 915 1552 919
rect 1636 915 1640 919
rect 1716 917 1720 921
rect 1812 917 1816 921
rect 1916 917 1920 921
rect 2036 917 2040 921
rect 2172 917 2176 921
rect 2316 915 2320 919
rect 2460 915 2464 919
rect 284 863 288 867
rect 380 863 384 867
rect 476 863 480 867
rect 580 863 584 867
rect 684 863 688 867
rect 780 863 784 867
rect 876 863 880 867
rect 964 863 968 867
rect 1044 863 1048 867
rect 1124 863 1128 867
rect 1204 863 1208 867
rect 1260 863 1264 867
rect 1524 855 1528 859
rect 1596 855 1600 859
rect 1660 855 1664 859
rect 1724 855 1728 859
rect 1788 855 1792 859
rect 1852 855 1856 859
rect 1924 855 1928 859
rect 2012 855 2016 859
rect 2116 855 2120 859
rect 2236 855 2240 859
rect 2356 855 2360 859
rect 2476 855 2480 859
rect 268 847 272 851
rect 364 849 368 853
rect 460 849 464 853
rect 564 849 568 853
rect 668 849 672 853
rect 764 847 768 851
rect 860 847 864 851
rect 948 849 952 853
rect 1028 849 1032 853
rect 1108 849 1112 853
rect 1188 849 1192 853
rect 1244 849 1248 853
rect 1508 839 1512 843
rect 1580 839 1584 843
rect 1644 841 1648 845
rect 1708 841 1712 845
rect 1772 839 1776 843
rect 1836 839 1840 843
rect 1908 841 1912 845
rect 1996 841 2000 845
rect 2100 841 2104 845
rect 2220 841 2224 845
rect 2340 841 2344 845
rect 2460 839 2464 843
rect 244 825 248 829
rect 308 823 312 827
rect 388 823 392 827
rect 468 823 472 827
rect 556 823 560 827
rect 644 823 648 827
rect 732 823 736 827
rect 812 823 816 827
rect 900 823 904 827
rect 988 823 992 827
rect 1076 823 1080 827
rect 1444 813 1448 817
rect 260 809 264 813
rect 324 807 328 811
rect 404 807 408 811
rect 484 809 488 813
rect 572 809 576 813
rect 660 809 664 813
rect 748 809 752 813
rect 828 809 832 813
rect 916 809 920 813
rect 1004 809 1008 813
rect 1516 811 1520 815
rect 1596 811 1600 815
rect 1676 813 1680 817
rect 1764 811 1768 815
rect 1852 811 1856 815
rect 1940 813 1944 817
rect 2028 811 2032 815
rect 2116 811 2120 815
rect 2204 811 2208 815
rect 2292 811 2296 815
rect 2388 811 2392 815
rect 2460 811 2464 815
rect 1092 807 1096 811
rect 1460 797 1464 801
rect 1532 797 1536 801
rect 1612 795 1616 799
rect 1692 797 1696 801
rect 1780 797 1784 801
rect 1868 797 1872 801
rect 1956 797 1960 801
rect 2044 797 2048 801
rect 2132 797 2136 801
rect 2220 797 2224 801
rect 2308 795 2312 799
rect 2404 795 2408 799
rect 2476 795 2480 799
rect 188 751 192 755
rect 284 751 288 755
rect 380 751 384 755
rect 476 751 480 755
rect 564 751 568 755
rect 644 751 648 755
rect 716 751 720 755
rect 788 751 792 755
rect 860 751 864 755
rect 932 751 936 755
rect 1012 751 1016 755
rect 172 735 176 739
rect 268 737 272 741
rect 364 735 368 739
rect 460 735 464 739
rect 548 737 552 741
rect 628 735 632 739
rect 700 737 704 741
rect 772 737 776 741
rect 844 737 848 741
rect 916 737 920 741
rect 996 737 1000 741
rect 1388 739 1392 743
rect 1484 739 1488 743
rect 1604 739 1608 743
rect 1724 739 1728 743
rect 1844 739 1848 743
rect 1964 739 1968 743
rect 2076 739 2080 743
rect 2180 739 2184 743
rect 2284 739 2288 743
rect 2388 739 2392 743
rect 2476 739 2480 743
rect 1372 725 1376 729
rect 1468 725 1472 729
rect 1588 723 1592 727
rect 1708 725 1712 729
rect 1828 723 1832 727
rect 1948 723 1952 727
rect 2060 725 2064 729
rect 2164 725 2168 729
rect 2268 725 2272 729
rect 2372 723 2376 727
rect 2460 723 2464 727
rect 180 711 184 715
rect 268 711 272 715
rect 348 711 352 715
rect 428 713 432 717
rect 508 711 512 715
rect 580 711 584 715
rect 644 711 648 715
rect 708 711 712 715
rect 772 711 776 715
rect 844 711 848 715
rect 916 711 920 715
rect 196 695 200 699
rect 284 697 288 701
rect 364 695 368 699
rect 444 697 448 701
rect 524 695 528 699
rect 596 695 600 699
rect 660 697 664 701
rect 724 697 728 701
rect 788 697 792 701
rect 860 697 864 701
rect 1372 699 1376 703
rect 1436 699 1440 703
rect 1540 699 1544 703
rect 1644 699 1648 703
rect 1756 699 1760 703
rect 1868 699 1872 703
rect 1972 699 1976 703
rect 2068 699 2072 703
rect 2156 699 2160 703
rect 2236 699 2240 703
rect 2316 699 2320 703
rect 2396 699 2400 703
rect 2460 699 2464 703
rect 932 695 936 699
rect 1388 685 1392 689
rect 1452 685 1456 689
rect 1556 685 1560 689
rect 1660 683 1664 687
rect 1772 685 1776 689
rect 1884 683 1888 687
rect 1988 685 1992 689
rect 2084 685 2088 689
rect 2172 685 2176 689
rect 2252 683 2256 687
rect 2332 685 2336 689
rect 2412 683 2416 687
rect 2476 683 2480 687
rect 252 643 256 647
rect 332 643 336 647
rect 412 643 416 647
rect 492 643 496 647
rect 564 643 568 647
rect 628 643 632 647
rect 692 643 696 647
rect 756 643 760 647
rect 820 643 824 647
rect 884 643 888 647
rect 956 643 960 647
rect 236 627 240 631
rect 316 629 320 633
rect 396 627 400 631
rect 476 629 480 633
rect 548 627 552 631
rect 612 629 616 633
rect 676 627 680 631
rect 740 629 744 633
rect 804 627 808 631
rect 868 627 872 631
rect 940 629 944 633
rect 1516 623 1520 627
rect 1596 623 1600 627
rect 1684 623 1688 627
rect 1772 623 1776 627
rect 1868 623 1872 627
rect 1956 623 1960 627
rect 2044 623 2048 627
rect 2124 623 2128 627
rect 2204 623 2208 627
rect 2276 623 2280 627
rect 2348 623 2352 627
rect 2420 623 2424 627
rect 2476 623 2480 627
rect 212 603 216 607
rect 308 603 312 607
rect 412 603 416 607
rect 508 603 512 607
rect 604 603 608 607
rect 692 605 696 609
rect 772 603 776 607
rect 852 603 856 607
rect 932 605 936 609
rect 1500 607 1504 611
rect 1580 609 1584 613
rect 1668 609 1672 613
rect 1756 607 1760 611
rect 1852 609 1856 613
rect 1940 607 1944 611
rect 2028 607 2032 611
rect 2108 609 2112 613
rect 2188 607 2192 611
rect 2260 607 2264 611
rect 2332 609 2336 613
rect 2404 607 2408 611
rect 2460 607 2464 611
rect 1012 603 1016 607
rect 1092 603 1096 607
rect 228 587 232 591
rect 324 589 328 593
rect 428 587 432 591
rect 524 589 528 593
rect 620 587 624 591
rect 708 589 712 593
rect 788 589 792 593
rect 868 587 872 591
rect 948 589 952 593
rect 1028 589 1032 593
rect 1108 587 1112 591
rect 1460 583 1464 587
rect 1564 583 1568 587
rect 1676 583 1680 587
rect 1780 583 1784 587
rect 1884 583 1888 587
rect 1988 585 1992 589
rect 2092 583 2096 587
rect 2188 583 2192 587
rect 2284 583 2288 587
rect 2380 583 2384 587
rect 2460 583 2464 587
rect 1476 567 1480 571
rect 1580 569 1584 573
rect 1692 569 1696 573
rect 1796 569 1800 573
rect 1900 567 1904 571
rect 2004 569 2008 573
rect 2108 567 2112 571
rect 2204 569 2208 573
rect 2300 567 2304 571
rect 2396 567 2400 571
rect 2476 567 2480 571
rect 212 531 216 535
rect 308 531 312 535
rect 412 531 416 535
rect 524 531 528 535
rect 628 531 632 535
rect 732 531 736 535
rect 828 531 832 535
rect 916 531 920 535
rect 1004 531 1008 535
rect 1092 531 1096 535
rect 1188 531 1192 535
rect 196 515 200 519
rect 292 515 296 519
rect 396 517 400 521
rect 508 515 512 519
rect 612 517 616 521
rect 716 517 720 521
rect 812 515 816 519
rect 900 517 904 521
rect 988 517 992 521
rect 1076 515 1080 519
rect 1172 517 1176 521
rect 1404 511 1408 515
rect 1484 511 1488 515
rect 1564 511 1568 515
rect 1652 511 1656 515
rect 1748 511 1752 515
rect 1836 511 1840 515
rect 1924 511 1928 515
rect 2012 511 2016 515
rect 2100 511 2104 515
rect 2188 511 2192 515
rect 2284 511 2288 515
rect 2380 511 2384 515
rect 2476 511 2480 515
rect 156 491 160 495
rect 252 491 256 495
rect 372 491 376 495
rect 492 491 496 495
rect 620 491 624 495
rect 740 491 744 495
rect 852 493 856 497
rect 1388 495 1392 499
rect 1468 495 1472 499
rect 1548 497 1552 501
rect 1636 495 1640 499
rect 1732 497 1736 501
rect 1820 497 1824 501
rect 1908 495 1912 499
rect 1996 497 2000 501
rect 2084 497 2088 501
rect 2172 495 2176 499
rect 2268 497 2272 501
rect 2364 497 2368 501
rect 2460 495 2464 499
rect 956 491 960 495
rect 1060 491 1064 495
rect 1164 491 1168 495
rect 1244 491 1248 495
rect 172 475 176 479
rect 268 477 272 481
rect 388 477 392 481
rect 508 475 512 479
rect 636 475 640 479
rect 756 477 760 481
rect 868 477 872 481
rect 972 477 976 481
rect 1076 475 1080 479
rect 1180 475 1184 479
rect 1260 477 1264 481
rect 1372 473 1376 477
rect 1436 471 1440 475
rect 1524 471 1528 475
rect 1620 471 1624 475
rect 1716 471 1720 475
rect 1820 473 1824 477
rect 1932 471 1936 475
rect 2060 471 2064 475
rect 2196 471 2200 475
rect 2340 471 2344 475
rect 2460 471 2464 475
rect 1388 457 1392 461
rect 1452 457 1456 461
rect 1540 455 1544 459
rect 1636 457 1640 461
rect 1732 455 1736 459
rect 1836 457 1840 461
rect 1948 455 1952 459
rect 2076 455 2080 459
rect 2212 457 2216 461
rect 2356 455 2360 459
rect 2476 455 2480 459
rect 172 419 176 423
rect 228 419 232 423
rect 284 419 288 423
rect 340 419 344 423
rect 420 419 424 423
rect 508 419 512 423
rect 604 419 608 423
rect 708 419 712 423
rect 820 419 824 423
rect 932 419 936 423
rect 1044 419 1048 423
rect 1164 419 1168 423
rect 1260 419 1264 423
rect 156 403 160 407
rect 212 405 216 409
rect 268 403 272 407
rect 324 405 328 409
rect 404 405 408 409
rect 492 403 496 407
rect 588 403 592 407
rect 692 405 696 409
rect 804 405 808 409
rect 916 405 920 409
rect 1028 403 1032 407
rect 1148 405 1152 409
rect 1244 405 1248 409
rect 1388 399 1392 403
rect 1460 399 1464 403
rect 1548 399 1552 403
rect 1636 399 1640 403
rect 1716 399 1720 403
rect 1812 399 1816 403
rect 1924 399 1928 403
rect 2052 399 2056 403
rect 2196 399 2200 403
rect 2348 399 2352 403
rect 2476 399 2480 403
rect 1372 385 1376 389
rect 1444 383 1448 387
rect 1532 385 1536 389
rect 1620 383 1624 387
rect 1700 383 1704 387
rect 1796 385 1800 389
rect 1908 383 1912 387
rect 2036 383 2040 387
rect 2180 385 2184 389
rect 2332 385 2336 389
rect 2460 383 2464 387
rect 156 377 160 381
rect 212 375 216 379
rect 284 375 288 379
rect 364 377 368 381
rect 436 375 440 379
rect 516 375 520 379
rect 596 375 600 379
rect 676 375 680 379
rect 756 377 760 381
rect 828 375 832 379
rect 900 375 904 379
rect 972 375 976 379
rect 1044 375 1048 379
rect 1116 375 1120 379
rect 1188 375 1192 379
rect 1244 375 1248 379
rect 172 359 176 363
rect 228 361 232 365
rect 300 359 304 363
rect 380 361 384 365
rect 452 361 456 365
rect 532 359 536 363
rect 612 359 616 363
rect 692 361 696 365
rect 772 361 776 365
rect 844 359 848 363
rect 916 361 920 365
rect 988 359 992 363
rect 1060 361 1064 365
rect 1132 361 1136 365
rect 1204 359 1208 363
rect 1260 361 1264 365
rect 1684 359 1688 363
rect 1740 359 1744 363
rect 1812 359 1816 363
rect 1908 359 1912 363
rect 2028 359 2032 363
rect 2164 359 2168 363
rect 2308 359 2312 363
rect 2460 359 2464 363
rect 1700 345 1704 349
rect 1756 343 1760 347
rect 1828 345 1832 349
rect 1924 345 1928 349
rect 2044 345 2048 349
rect 2180 345 2184 349
rect 2324 343 2328 347
rect 2476 343 2480 347
rect 172 299 176 303
rect 236 299 240 303
rect 324 299 328 303
rect 412 299 416 303
rect 492 299 496 303
rect 580 299 584 303
rect 668 299 672 303
rect 764 299 768 303
rect 860 299 864 303
rect 964 299 968 303
rect 1068 299 1072 303
rect 1172 299 1176 303
rect 1260 299 1264 303
rect 1388 291 1392 295
rect 1468 291 1472 295
rect 1564 291 1568 295
rect 1660 291 1664 295
rect 1748 291 1752 295
rect 1844 291 1848 295
rect 1948 291 1952 295
rect 2060 291 2064 295
rect 2188 291 2192 295
rect 2324 291 2328 295
rect 2460 291 2464 295
rect 156 283 160 287
rect 220 285 224 289
rect 308 285 312 289
rect 396 283 400 287
rect 476 285 480 289
rect 564 283 568 287
rect 652 283 656 287
rect 748 285 752 289
rect 844 285 848 289
rect 948 285 952 289
rect 1052 285 1056 289
rect 1156 283 1160 287
rect 1244 283 1248 287
rect 1372 275 1376 279
rect 1452 277 1456 281
rect 1548 277 1552 281
rect 1644 277 1648 281
rect 1732 275 1736 279
rect 1828 275 1832 279
rect 1932 277 1936 281
rect 2044 277 2048 281
rect 2172 277 2176 281
rect 2308 277 2312 281
rect 2444 275 2448 279
rect 156 257 160 261
rect 236 255 240 259
rect 332 255 336 259
rect 428 257 432 261
rect 524 255 528 259
rect 620 255 624 259
rect 716 257 720 261
rect 812 255 816 259
rect 908 255 912 259
rect 1012 255 1016 259
rect 1116 255 1120 259
rect 1220 255 1224 259
rect 1372 253 1376 257
rect 1444 251 1448 255
rect 1540 251 1544 255
rect 1636 253 1640 257
rect 1732 251 1736 255
rect 1820 251 1824 255
rect 1908 253 1912 257
rect 2004 251 2008 255
rect 2108 251 2112 255
rect 2220 251 2224 255
rect 2340 251 2344 255
rect 2460 251 2464 255
rect 172 241 176 245
rect 252 239 256 243
rect 348 239 352 243
rect 444 241 448 245
rect 540 239 544 243
rect 636 239 640 243
rect 732 241 736 245
rect 828 239 832 243
rect 924 239 928 243
rect 1028 241 1032 245
rect 1132 241 1136 245
rect 1236 239 1240 243
rect 1388 237 1392 241
rect 1460 237 1464 241
rect 1556 235 1560 239
rect 1652 237 1656 241
rect 1748 237 1752 241
rect 1836 237 1840 241
rect 1924 237 1928 241
rect 2020 237 2024 241
rect 2124 237 2128 241
rect 2236 237 2240 241
rect 2356 235 2360 239
rect 2476 235 2480 239
rect 196 179 200 183
rect 276 179 280 183
rect 364 179 368 183
rect 452 179 456 183
rect 548 179 552 183
rect 644 179 648 183
rect 732 179 736 183
rect 820 179 824 183
rect 908 179 912 183
rect 996 179 1000 183
rect 1084 179 1088 183
rect 1172 179 1176 183
rect 1428 179 1432 183
rect 1532 179 1536 183
rect 1636 179 1640 183
rect 1748 179 1752 183
rect 1852 179 1856 183
rect 1956 179 1960 183
rect 2052 179 2056 183
rect 2148 179 2152 183
rect 2236 179 2240 183
rect 2324 179 2328 183
rect 2412 179 2416 183
rect 2476 179 2480 183
rect 180 163 184 167
rect 260 163 264 167
rect 348 165 352 169
rect 436 163 440 167
rect 532 165 536 169
rect 628 165 632 169
rect 716 163 720 167
rect 804 165 808 169
rect 892 163 896 167
rect 980 165 984 169
rect 1068 165 1072 169
rect 1156 163 1160 167
rect 1412 163 1416 167
rect 1516 165 1520 169
rect 1620 163 1624 167
rect 1732 165 1736 169
rect 1836 163 1840 167
rect 1940 163 1944 167
rect 2036 165 2040 169
rect 2132 165 2136 169
rect 2220 165 2224 169
rect 2308 163 2312 167
rect 2396 165 2400 169
rect 2460 163 2464 167
rect 156 125 160 129
rect 212 123 216 127
rect 268 123 272 127
rect 324 123 328 127
rect 380 123 384 127
rect 436 123 440 127
rect 492 123 496 127
rect 556 123 560 127
rect 628 123 632 127
rect 692 125 696 129
rect 756 123 760 127
rect 820 123 824 127
rect 884 123 888 127
rect 948 123 952 127
rect 1012 123 1016 127
rect 1076 123 1080 127
rect 1140 123 1144 127
rect 1204 123 1208 127
rect 1372 125 1376 129
rect 1428 123 1432 127
rect 1484 123 1488 127
rect 1540 123 1544 127
rect 1596 123 1600 127
rect 1652 123 1656 127
rect 1708 123 1712 127
rect 1764 123 1768 127
rect 1820 123 1824 127
rect 1876 125 1880 129
rect 1932 123 1936 127
rect 1988 123 1992 127
rect 2044 123 2048 127
rect 2100 123 2104 127
rect 2164 123 2168 127
rect 2228 123 2232 127
rect 2292 123 2296 127
rect 2348 123 2352 127
rect 2404 123 2408 127
rect 2460 123 2464 127
rect 172 109 176 113
rect 228 109 232 113
rect 284 109 288 113
rect 340 109 344 113
rect 396 109 400 113
rect 452 109 456 113
rect 508 109 512 113
rect 572 109 576 113
rect 644 107 648 111
rect 708 109 712 113
rect 772 109 776 113
rect 836 109 840 113
rect 900 109 904 113
rect 964 109 968 113
rect 1028 109 1032 113
rect 1092 109 1096 113
rect 1156 109 1160 113
rect 1220 107 1224 111
rect 1388 109 1392 113
rect 1444 109 1448 113
rect 1500 109 1504 113
rect 1556 109 1560 113
rect 1612 109 1616 113
rect 1668 109 1672 113
rect 1724 109 1728 113
rect 1780 109 1784 113
rect 1836 107 1840 111
rect 1892 109 1896 113
rect 1948 109 1952 113
rect 2004 109 2008 113
rect 2060 109 2064 113
rect 2116 109 2120 113
rect 2180 109 2184 113
rect 2244 109 2248 113
rect 2308 109 2312 113
rect 2364 107 2368 111
rect 2476 109 2480 113
<< m2 >>
rect 779 2571 785 2572
rect 779 2570 780 2571
rect 756 2568 780 2570
rect 756 2562 758 2568
rect 779 2567 780 2568
rect 784 2567 785 2571
rect 835 2571 841 2572
rect 835 2570 836 2571
rect 779 2566 785 2567
rect 800 2568 836 2570
rect 800 2562 802 2568
rect 835 2567 836 2568
rect 840 2567 841 2571
rect 891 2571 897 2572
rect 891 2570 892 2571
rect 835 2566 841 2567
rect 872 2568 892 2570
rect 872 2562 874 2568
rect 891 2567 892 2568
rect 896 2567 897 2571
rect 947 2571 953 2572
rect 947 2570 948 2571
rect 891 2566 897 2567
rect 924 2568 948 2570
rect 924 2562 926 2568
rect 947 2567 948 2568
rect 952 2567 953 2571
rect 947 2566 953 2567
rect 740 2560 758 2562
rect 796 2560 802 2562
rect 852 2560 874 2562
rect 908 2560 926 2562
rect 740 2558 742 2560
rect 796 2558 798 2560
rect 852 2558 854 2560
rect 908 2558 910 2560
rect 718 2557 724 2558
rect 110 2556 116 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 718 2553 719 2557
rect 723 2553 724 2557
rect 718 2552 724 2553
rect 739 2557 745 2558
rect 739 2553 740 2557
rect 744 2553 745 2557
rect 739 2552 745 2553
rect 774 2557 780 2558
rect 774 2553 775 2557
rect 779 2553 780 2557
rect 774 2552 780 2553
rect 795 2557 801 2558
rect 795 2553 796 2557
rect 800 2553 801 2557
rect 795 2552 801 2553
rect 830 2557 836 2558
rect 830 2553 831 2557
rect 835 2553 836 2557
rect 830 2552 836 2553
rect 851 2557 857 2558
rect 851 2553 852 2557
rect 856 2553 857 2557
rect 851 2552 857 2553
rect 886 2557 892 2558
rect 886 2553 887 2557
rect 891 2553 892 2557
rect 886 2552 892 2553
rect 907 2557 913 2558
rect 907 2553 908 2557
rect 912 2553 913 2557
rect 907 2552 913 2553
rect 942 2557 948 2558
rect 942 2553 943 2557
rect 947 2553 948 2557
rect 1286 2556 1292 2557
rect 942 2552 948 2553
rect 950 2555 956 2556
rect 110 2551 116 2552
rect 950 2551 951 2555
rect 955 2554 956 2555
rect 963 2555 969 2556
rect 963 2554 964 2555
rect 955 2552 964 2554
rect 955 2551 956 2552
rect 950 2550 956 2551
rect 963 2551 964 2552
rect 968 2551 969 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1710 2555 1716 2556
rect 1710 2554 1711 2555
rect 1286 2551 1292 2552
rect 1404 2552 1711 2554
rect 963 2550 969 2551
rect 1404 2550 1406 2552
rect 1710 2551 1711 2552
rect 1715 2551 1716 2555
rect 1710 2550 1716 2551
rect 1403 2549 1409 2550
rect 1403 2545 1404 2549
rect 1408 2545 1409 2549
rect 1459 2547 1465 2548
rect 1459 2546 1460 2547
rect 1403 2544 1409 2545
rect 1424 2544 1460 2546
rect 110 2539 116 2540
rect 110 2535 111 2539
rect 115 2535 116 2539
rect 1286 2539 1292 2540
rect 110 2534 116 2535
rect 702 2536 708 2537
rect 702 2532 703 2536
rect 707 2532 708 2536
rect 702 2531 708 2532
rect 758 2536 764 2537
rect 758 2532 759 2536
rect 763 2532 764 2536
rect 758 2531 764 2532
rect 814 2536 820 2537
rect 814 2532 815 2536
rect 819 2532 820 2536
rect 814 2531 820 2532
rect 870 2536 876 2537
rect 870 2532 871 2536
rect 875 2532 876 2536
rect 870 2531 876 2532
rect 926 2536 932 2537
rect 926 2532 927 2536
rect 931 2532 932 2536
rect 1286 2535 1287 2539
rect 1291 2535 1292 2539
rect 1424 2538 1426 2544
rect 1459 2543 1460 2544
rect 1464 2543 1465 2547
rect 1515 2547 1521 2548
rect 1515 2546 1516 2547
rect 1459 2542 1465 2543
rect 1480 2544 1516 2546
rect 1480 2538 1482 2544
rect 1515 2543 1516 2544
rect 1520 2543 1521 2547
rect 1571 2547 1577 2548
rect 1571 2546 1572 2547
rect 1515 2542 1521 2543
rect 1548 2544 1572 2546
rect 1548 2538 1550 2544
rect 1571 2543 1572 2544
rect 1576 2543 1577 2547
rect 1627 2547 1633 2548
rect 1627 2546 1628 2547
rect 1571 2542 1577 2543
rect 1604 2544 1628 2546
rect 1604 2538 1606 2544
rect 1627 2543 1628 2544
rect 1632 2543 1633 2547
rect 1683 2547 1689 2548
rect 1683 2546 1684 2547
rect 1627 2542 1633 2543
rect 1656 2544 1684 2546
rect 1656 2538 1658 2544
rect 1683 2543 1684 2544
rect 1688 2543 1689 2547
rect 1739 2547 1745 2548
rect 1739 2546 1740 2547
rect 1683 2542 1689 2543
rect 1704 2544 1740 2546
rect 1704 2538 1706 2544
rect 1739 2543 1740 2544
rect 1744 2543 1745 2547
rect 1795 2547 1801 2548
rect 1795 2546 1796 2547
rect 1739 2542 1745 2543
rect 1768 2544 1796 2546
rect 1768 2538 1770 2544
rect 1795 2543 1796 2544
rect 1800 2543 1801 2547
rect 1851 2547 1857 2548
rect 1851 2546 1852 2547
rect 1795 2542 1801 2543
rect 1812 2544 1852 2546
rect 1286 2534 1292 2535
rect 1420 2536 1426 2538
rect 1476 2536 1482 2538
rect 1532 2536 1550 2538
rect 1588 2536 1606 2538
rect 1644 2536 1658 2538
rect 1700 2536 1706 2538
rect 1756 2536 1770 2538
rect 1420 2534 1422 2536
rect 1476 2534 1478 2536
rect 1532 2534 1534 2536
rect 1588 2534 1590 2536
rect 1644 2534 1646 2536
rect 1700 2534 1702 2536
rect 1756 2534 1758 2536
rect 1812 2534 1814 2544
rect 1851 2543 1852 2544
rect 1856 2543 1857 2547
rect 1907 2547 1913 2548
rect 1907 2546 1908 2547
rect 1851 2542 1857 2543
rect 1884 2544 1908 2546
rect 1884 2538 1886 2544
rect 1907 2543 1908 2544
rect 1912 2543 1913 2547
rect 1963 2547 1969 2548
rect 1963 2546 1964 2547
rect 1907 2542 1913 2543
rect 1940 2544 1964 2546
rect 1940 2538 1942 2544
rect 1963 2543 1964 2544
rect 1968 2543 1969 2547
rect 2019 2547 2025 2548
rect 2019 2546 2020 2547
rect 1963 2542 1969 2543
rect 1999 2544 2020 2546
rect 1999 2538 2001 2544
rect 2019 2543 2020 2544
rect 2024 2543 2025 2547
rect 2075 2547 2081 2548
rect 2075 2546 2076 2547
rect 2019 2542 2025 2543
rect 2052 2544 2076 2546
rect 2052 2538 2054 2544
rect 2075 2543 2076 2544
rect 2080 2543 2081 2547
rect 2131 2547 2137 2548
rect 2131 2546 2132 2547
rect 2075 2542 2081 2543
rect 2108 2544 2132 2546
rect 2108 2538 2110 2544
rect 2131 2543 2132 2544
rect 2136 2543 2137 2547
rect 2187 2547 2193 2548
rect 2187 2546 2188 2547
rect 2131 2542 2137 2543
rect 2164 2544 2188 2546
rect 2164 2538 2166 2544
rect 2187 2543 2188 2544
rect 2192 2543 2193 2547
rect 2187 2542 2193 2543
rect 1868 2536 1886 2538
rect 1924 2536 1942 2538
rect 1980 2536 2001 2538
rect 2036 2536 2054 2538
rect 2092 2536 2110 2538
rect 2148 2536 2166 2538
rect 1868 2534 1870 2536
rect 1924 2534 1926 2536
rect 1980 2534 1982 2536
rect 2036 2534 2038 2536
rect 2092 2534 2094 2536
rect 2148 2534 2150 2536
rect 1398 2533 1404 2534
rect 926 2531 932 2532
rect 1326 2532 1332 2533
rect 1326 2528 1327 2532
rect 1331 2528 1332 2532
rect 1398 2529 1399 2533
rect 1403 2529 1404 2533
rect 1398 2528 1404 2529
rect 1419 2533 1425 2534
rect 1419 2529 1420 2533
rect 1424 2529 1425 2533
rect 1419 2528 1425 2529
rect 1454 2533 1460 2534
rect 1454 2529 1455 2533
rect 1459 2529 1460 2533
rect 1454 2528 1460 2529
rect 1475 2533 1481 2534
rect 1475 2529 1476 2533
rect 1480 2529 1481 2533
rect 1475 2528 1481 2529
rect 1510 2533 1516 2534
rect 1510 2529 1511 2533
rect 1515 2529 1516 2533
rect 1510 2528 1516 2529
rect 1531 2533 1537 2534
rect 1531 2529 1532 2533
rect 1536 2529 1537 2533
rect 1531 2528 1537 2529
rect 1566 2533 1572 2534
rect 1566 2529 1567 2533
rect 1571 2529 1572 2533
rect 1566 2528 1572 2529
rect 1587 2533 1593 2534
rect 1587 2529 1588 2533
rect 1592 2529 1593 2533
rect 1587 2528 1593 2529
rect 1622 2533 1628 2534
rect 1622 2529 1623 2533
rect 1627 2529 1628 2533
rect 1622 2528 1628 2529
rect 1643 2533 1649 2534
rect 1643 2529 1644 2533
rect 1648 2529 1649 2533
rect 1643 2528 1649 2529
rect 1678 2533 1684 2534
rect 1678 2529 1679 2533
rect 1683 2529 1684 2533
rect 1678 2528 1684 2529
rect 1699 2533 1705 2534
rect 1699 2529 1700 2533
rect 1704 2529 1705 2533
rect 1699 2528 1705 2529
rect 1734 2533 1740 2534
rect 1734 2529 1735 2533
rect 1739 2529 1740 2533
rect 1734 2528 1740 2529
rect 1755 2533 1761 2534
rect 1755 2529 1756 2533
rect 1760 2529 1761 2533
rect 1755 2528 1761 2529
rect 1790 2533 1796 2534
rect 1790 2529 1791 2533
rect 1795 2529 1796 2533
rect 1790 2528 1796 2529
rect 1811 2533 1817 2534
rect 1811 2529 1812 2533
rect 1816 2529 1817 2533
rect 1811 2528 1817 2529
rect 1846 2533 1852 2534
rect 1846 2529 1847 2533
rect 1851 2529 1852 2533
rect 1846 2528 1852 2529
rect 1867 2533 1873 2534
rect 1867 2529 1868 2533
rect 1872 2529 1873 2533
rect 1867 2528 1873 2529
rect 1902 2533 1908 2534
rect 1902 2529 1903 2533
rect 1907 2529 1908 2533
rect 1902 2528 1908 2529
rect 1923 2533 1929 2534
rect 1923 2529 1924 2533
rect 1928 2529 1929 2533
rect 1923 2528 1929 2529
rect 1958 2533 1964 2534
rect 1958 2529 1959 2533
rect 1963 2529 1964 2533
rect 1958 2528 1964 2529
rect 1979 2533 1985 2534
rect 1979 2529 1980 2533
rect 1984 2529 1985 2533
rect 1979 2528 1985 2529
rect 2014 2533 2020 2534
rect 2014 2529 2015 2533
rect 2019 2529 2020 2533
rect 2014 2528 2020 2529
rect 2035 2533 2041 2534
rect 2035 2529 2036 2533
rect 2040 2529 2041 2533
rect 2035 2528 2041 2529
rect 2070 2533 2076 2534
rect 2070 2529 2071 2533
rect 2075 2529 2076 2533
rect 2070 2528 2076 2529
rect 2091 2533 2097 2534
rect 2091 2529 2092 2533
rect 2096 2529 2097 2533
rect 2091 2528 2097 2529
rect 2126 2533 2132 2534
rect 2126 2529 2127 2533
rect 2131 2529 2132 2533
rect 2126 2528 2132 2529
rect 2147 2533 2153 2534
rect 2147 2529 2148 2533
rect 2152 2529 2153 2533
rect 2147 2528 2153 2529
rect 2182 2533 2188 2534
rect 2182 2529 2183 2533
rect 2187 2529 2188 2533
rect 2502 2532 2508 2533
rect 2182 2528 2188 2529
rect 2190 2531 2196 2532
rect 1326 2527 1332 2528
rect 2190 2527 2191 2531
rect 2195 2530 2196 2531
rect 2203 2531 2209 2532
rect 2203 2530 2204 2531
rect 2195 2528 2204 2530
rect 2195 2527 2196 2528
rect 2190 2526 2196 2527
rect 2203 2527 2204 2528
rect 2208 2527 2209 2531
rect 2502 2528 2503 2532
rect 2507 2528 2508 2532
rect 2502 2527 2508 2528
rect 2203 2526 2209 2527
rect 166 2524 172 2525
rect 110 2521 116 2522
rect 110 2517 111 2521
rect 115 2517 116 2521
rect 166 2520 167 2524
rect 171 2520 172 2524
rect 166 2519 172 2520
rect 222 2524 228 2525
rect 222 2520 223 2524
rect 227 2520 228 2524
rect 222 2519 228 2520
rect 278 2524 284 2525
rect 278 2520 279 2524
rect 283 2520 284 2524
rect 278 2519 284 2520
rect 342 2524 348 2525
rect 342 2520 343 2524
rect 347 2520 348 2524
rect 342 2519 348 2520
rect 406 2524 412 2525
rect 406 2520 407 2524
rect 411 2520 412 2524
rect 406 2519 412 2520
rect 478 2524 484 2525
rect 478 2520 479 2524
rect 483 2520 484 2524
rect 478 2519 484 2520
rect 558 2524 564 2525
rect 558 2520 559 2524
rect 563 2520 564 2524
rect 558 2519 564 2520
rect 638 2524 644 2525
rect 638 2520 639 2524
rect 643 2520 644 2524
rect 638 2519 644 2520
rect 718 2524 724 2525
rect 718 2520 719 2524
rect 723 2520 724 2524
rect 718 2519 724 2520
rect 798 2524 804 2525
rect 798 2520 799 2524
rect 803 2520 804 2524
rect 798 2519 804 2520
rect 878 2524 884 2525
rect 878 2520 879 2524
rect 883 2520 884 2524
rect 878 2519 884 2520
rect 958 2524 964 2525
rect 958 2520 959 2524
rect 963 2520 964 2524
rect 958 2519 964 2520
rect 1038 2524 1044 2525
rect 1038 2520 1039 2524
rect 1043 2520 1044 2524
rect 1038 2519 1044 2520
rect 1286 2521 1292 2522
rect 110 2516 116 2517
rect 1286 2517 1287 2521
rect 1291 2517 1292 2521
rect 1286 2516 1292 2517
rect 1326 2515 1332 2516
rect 1326 2511 1327 2515
rect 1331 2511 1332 2515
rect 2502 2515 2508 2516
rect 1326 2510 1332 2511
rect 1382 2512 1388 2513
rect 1382 2508 1383 2512
rect 1387 2508 1388 2512
rect 1382 2507 1388 2508
rect 1438 2512 1444 2513
rect 1438 2508 1439 2512
rect 1443 2508 1444 2512
rect 1438 2507 1444 2508
rect 1494 2512 1500 2513
rect 1494 2508 1495 2512
rect 1499 2508 1500 2512
rect 1494 2507 1500 2508
rect 1550 2512 1556 2513
rect 1550 2508 1551 2512
rect 1555 2508 1556 2512
rect 1550 2507 1556 2508
rect 1606 2512 1612 2513
rect 1606 2508 1607 2512
rect 1611 2508 1612 2512
rect 1606 2507 1612 2508
rect 1662 2512 1668 2513
rect 1662 2508 1663 2512
rect 1667 2508 1668 2512
rect 1662 2507 1668 2508
rect 1718 2512 1724 2513
rect 1718 2508 1719 2512
rect 1723 2508 1724 2512
rect 1718 2507 1724 2508
rect 1774 2512 1780 2513
rect 1774 2508 1775 2512
rect 1779 2508 1780 2512
rect 1774 2507 1780 2508
rect 1830 2512 1836 2513
rect 1830 2508 1831 2512
rect 1835 2508 1836 2512
rect 1830 2507 1836 2508
rect 1886 2512 1892 2513
rect 1886 2508 1887 2512
rect 1891 2508 1892 2512
rect 1886 2507 1892 2508
rect 1942 2512 1948 2513
rect 1942 2508 1943 2512
rect 1947 2508 1948 2512
rect 1942 2507 1948 2508
rect 1998 2512 2004 2513
rect 1998 2508 1999 2512
rect 2003 2508 2004 2512
rect 1998 2507 2004 2508
rect 2054 2512 2060 2513
rect 2054 2508 2055 2512
rect 2059 2508 2060 2512
rect 2054 2507 2060 2508
rect 2110 2512 2116 2513
rect 2110 2508 2111 2512
rect 2115 2508 2116 2512
rect 2110 2507 2116 2508
rect 2166 2512 2172 2513
rect 2166 2508 2167 2512
rect 2171 2508 2172 2512
rect 2502 2511 2503 2515
rect 2507 2511 2508 2515
rect 2502 2510 2508 2511
rect 2166 2507 2172 2508
rect 110 2504 116 2505
rect 1286 2504 1292 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 110 2499 116 2500
rect 182 2503 188 2504
rect 182 2499 183 2503
rect 187 2499 188 2503
rect 182 2498 188 2499
rect 203 2503 209 2504
rect 203 2499 204 2503
rect 208 2502 209 2503
rect 238 2503 244 2504
rect 208 2500 234 2502
rect 208 2499 209 2500
rect 203 2498 209 2499
rect 232 2490 234 2500
rect 238 2499 239 2503
rect 243 2499 244 2503
rect 238 2498 244 2499
rect 254 2503 265 2504
rect 254 2499 255 2503
rect 259 2499 260 2503
rect 264 2499 265 2503
rect 254 2498 265 2499
rect 294 2503 300 2504
rect 294 2499 295 2503
rect 299 2499 300 2503
rect 315 2503 321 2504
rect 315 2502 316 2503
rect 294 2498 300 2499
rect 304 2500 316 2502
rect 304 2494 306 2500
rect 315 2499 316 2500
rect 320 2499 321 2503
rect 315 2498 321 2499
rect 358 2503 364 2504
rect 358 2499 359 2503
rect 363 2499 364 2503
rect 358 2498 364 2499
rect 379 2503 385 2504
rect 379 2499 380 2503
rect 384 2499 385 2503
rect 379 2498 385 2499
rect 422 2503 428 2504
rect 422 2499 423 2503
rect 427 2499 428 2503
rect 443 2503 449 2504
rect 443 2502 444 2503
rect 422 2498 428 2499
rect 432 2500 444 2502
rect 381 2494 383 2498
rect 432 2494 434 2500
rect 443 2499 444 2500
rect 448 2499 449 2503
rect 443 2498 449 2499
rect 494 2503 500 2504
rect 494 2499 495 2503
rect 499 2499 500 2503
rect 515 2503 521 2504
rect 515 2502 516 2503
rect 494 2498 500 2499
rect 504 2500 516 2502
rect 504 2494 506 2500
rect 515 2499 516 2500
rect 520 2499 521 2503
rect 515 2498 521 2499
rect 574 2503 580 2504
rect 574 2499 575 2503
rect 579 2499 580 2503
rect 574 2498 580 2499
rect 590 2503 601 2504
rect 590 2499 591 2503
rect 595 2499 596 2503
rect 600 2499 601 2503
rect 590 2498 601 2499
rect 654 2503 660 2504
rect 654 2499 655 2503
rect 659 2499 660 2503
rect 675 2503 681 2504
rect 675 2502 676 2503
rect 654 2498 660 2499
rect 664 2500 676 2502
rect 664 2494 666 2500
rect 675 2499 676 2500
rect 680 2499 681 2503
rect 675 2498 681 2499
rect 734 2503 740 2504
rect 734 2499 735 2503
rect 739 2499 740 2503
rect 734 2498 740 2499
rect 755 2503 761 2504
rect 755 2499 756 2503
rect 760 2502 761 2503
rect 814 2503 820 2504
rect 760 2500 810 2502
rect 760 2499 761 2500
rect 755 2498 761 2499
rect 252 2492 306 2494
rect 319 2492 383 2494
rect 388 2492 434 2494
rect 436 2492 506 2494
rect 580 2492 666 2494
rect 232 2489 249 2490
rect 232 2488 244 2489
rect 187 2487 193 2488
rect 187 2483 188 2487
rect 192 2486 193 2487
rect 192 2484 238 2486
rect 243 2485 244 2488
rect 248 2485 249 2489
rect 243 2484 249 2485
rect 192 2483 193 2484
rect 187 2482 193 2483
rect 236 2482 238 2484
rect 252 2482 254 2492
rect 299 2487 305 2488
rect 299 2483 300 2487
rect 304 2486 305 2487
rect 319 2486 321 2492
rect 388 2490 390 2492
rect 436 2490 438 2492
rect 580 2490 582 2492
rect 808 2490 810 2500
rect 814 2499 815 2503
rect 819 2499 820 2503
rect 814 2498 820 2499
rect 835 2503 841 2504
rect 835 2499 836 2503
rect 840 2502 841 2503
rect 894 2503 900 2504
rect 840 2500 890 2502
rect 840 2499 841 2500
rect 835 2498 841 2499
rect 888 2490 890 2500
rect 894 2499 895 2503
rect 899 2499 900 2503
rect 894 2498 900 2499
rect 915 2503 921 2504
rect 915 2499 916 2503
rect 920 2502 921 2503
rect 974 2503 980 2504
rect 920 2500 970 2502
rect 920 2499 921 2500
rect 915 2498 921 2499
rect 968 2490 970 2500
rect 974 2499 975 2503
rect 979 2499 980 2503
rect 974 2498 980 2499
rect 995 2503 1001 2504
rect 995 2499 996 2503
rect 1000 2502 1001 2503
rect 1054 2503 1060 2504
rect 1000 2500 1046 2502
rect 1000 2499 1001 2500
rect 995 2498 1001 2499
rect 1044 2490 1046 2500
rect 1054 2499 1055 2503
rect 1059 2499 1060 2503
rect 1054 2498 1060 2499
rect 1070 2503 1081 2504
rect 1070 2499 1071 2503
rect 1075 2499 1076 2503
rect 1080 2499 1081 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1798 2499 1804 2500
rect 1070 2498 1081 2499
rect 1798 2495 1799 2499
rect 1803 2498 1804 2499
rect 2190 2499 2196 2500
rect 2190 2498 2191 2499
rect 1803 2496 2191 2498
rect 1803 2495 1804 2496
rect 1798 2494 1804 2495
rect 2190 2495 2191 2496
rect 2195 2495 2196 2499
rect 2190 2494 2196 2495
rect 1350 2492 1356 2493
rect 304 2484 321 2486
rect 363 2489 390 2490
rect 363 2485 364 2489
rect 368 2488 390 2489
rect 427 2489 438 2490
rect 368 2485 369 2488
rect 363 2484 369 2485
rect 427 2485 428 2489
rect 432 2488 438 2489
rect 579 2489 585 2490
rect 432 2485 433 2488
rect 427 2484 433 2485
rect 499 2487 505 2488
rect 304 2483 305 2484
rect 299 2482 305 2483
rect 499 2483 500 2487
rect 504 2486 505 2487
rect 504 2484 550 2486
rect 579 2485 580 2489
rect 584 2485 585 2489
rect 808 2489 825 2490
rect 808 2488 820 2489
rect 579 2484 585 2485
rect 622 2487 628 2488
rect 504 2483 505 2484
rect 499 2482 505 2483
rect 548 2482 550 2484
rect 590 2483 596 2484
rect 590 2482 591 2483
rect 236 2480 254 2482
rect 548 2480 591 2482
rect 590 2479 591 2480
rect 595 2479 596 2483
rect 622 2483 623 2487
rect 627 2486 628 2487
rect 659 2487 665 2488
rect 659 2486 660 2487
rect 627 2484 660 2486
rect 627 2483 628 2484
rect 622 2482 628 2483
rect 659 2483 660 2484
rect 664 2483 665 2487
rect 659 2482 665 2483
rect 739 2487 745 2488
rect 739 2483 740 2487
rect 744 2486 745 2487
rect 744 2484 814 2486
rect 819 2485 820 2488
rect 824 2485 825 2489
rect 888 2489 905 2490
rect 888 2488 900 2489
rect 819 2484 825 2485
rect 899 2485 900 2488
rect 904 2485 905 2489
rect 968 2489 985 2490
rect 968 2488 980 2489
rect 899 2484 905 2485
rect 979 2485 980 2488
rect 984 2485 985 2489
rect 1044 2489 1065 2490
rect 1044 2488 1060 2489
rect 979 2484 985 2485
rect 1059 2485 1060 2488
rect 1064 2485 1065 2489
rect 1059 2484 1065 2485
rect 1326 2489 1332 2490
rect 1326 2485 1327 2489
rect 1331 2485 1332 2489
rect 1350 2488 1351 2492
rect 1355 2488 1356 2492
rect 1350 2487 1356 2488
rect 1422 2492 1428 2493
rect 1422 2488 1423 2492
rect 1427 2488 1428 2492
rect 1422 2487 1428 2488
rect 1510 2492 1516 2493
rect 1510 2488 1511 2492
rect 1515 2488 1516 2492
rect 1510 2487 1516 2488
rect 1598 2492 1604 2493
rect 1598 2488 1599 2492
rect 1603 2488 1604 2492
rect 1598 2487 1604 2488
rect 1686 2492 1692 2493
rect 1686 2488 1687 2492
rect 1691 2488 1692 2492
rect 1686 2487 1692 2488
rect 1774 2492 1780 2493
rect 1774 2488 1775 2492
rect 1779 2488 1780 2492
rect 1774 2487 1780 2488
rect 1862 2492 1868 2493
rect 1862 2488 1863 2492
rect 1867 2488 1868 2492
rect 1862 2487 1868 2488
rect 1950 2492 1956 2493
rect 1950 2488 1951 2492
rect 1955 2488 1956 2492
rect 1950 2487 1956 2488
rect 2038 2492 2044 2493
rect 2038 2488 2039 2492
rect 2043 2488 2044 2492
rect 2038 2487 2044 2488
rect 2126 2492 2132 2493
rect 2126 2488 2127 2492
rect 2131 2488 2132 2492
rect 2126 2487 2132 2488
rect 2502 2489 2508 2490
rect 1326 2484 1332 2485
rect 2502 2485 2503 2489
rect 2507 2485 2508 2489
rect 2502 2484 2508 2485
rect 744 2483 745 2484
rect 739 2482 745 2483
rect 812 2482 814 2484
rect 950 2483 956 2484
rect 950 2482 951 2483
rect 812 2480 951 2482
rect 590 2478 596 2479
rect 950 2479 951 2480
rect 955 2479 956 2483
rect 950 2478 956 2479
rect 434 2475 440 2476
rect 434 2474 435 2475
rect 188 2472 435 2474
rect 188 2470 190 2472
rect 434 2471 435 2472
rect 439 2471 440 2475
rect 714 2475 720 2476
rect 714 2474 715 2475
rect 434 2470 440 2471
rect 508 2472 715 2474
rect 508 2470 510 2472
rect 714 2471 715 2472
rect 719 2471 720 2475
rect 1070 2475 1076 2476
rect 1070 2474 1071 2475
rect 714 2470 720 2471
rect 796 2472 1071 2474
rect 796 2470 798 2472
rect 1070 2471 1071 2472
rect 1075 2471 1076 2475
rect 1070 2470 1076 2471
rect 1326 2472 1332 2473
rect 2502 2472 2508 2473
rect 187 2469 193 2470
rect 187 2465 188 2469
rect 192 2465 193 2469
rect 507 2469 513 2470
rect 187 2464 193 2465
rect 251 2467 260 2468
rect 251 2463 252 2467
rect 259 2463 260 2467
rect 331 2467 337 2468
rect 331 2466 332 2467
rect 251 2462 260 2463
rect 319 2464 332 2466
rect 319 2454 321 2464
rect 331 2463 332 2464
rect 336 2463 337 2467
rect 419 2467 425 2468
rect 419 2466 420 2467
rect 331 2462 337 2463
rect 352 2464 420 2466
rect 352 2454 354 2464
rect 419 2463 420 2464
rect 424 2463 425 2467
rect 507 2465 508 2469
rect 512 2465 513 2469
rect 795 2469 801 2470
rect 603 2467 609 2468
rect 603 2466 604 2467
rect 507 2464 513 2465
rect 524 2464 604 2466
rect 419 2462 425 2463
rect 524 2454 526 2464
rect 603 2463 604 2464
rect 608 2463 609 2467
rect 603 2462 609 2463
rect 699 2467 705 2468
rect 699 2463 700 2467
rect 704 2466 705 2467
rect 762 2467 768 2468
rect 762 2466 763 2467
rect 704 2464 763 2466
rect 704 2463 705 2464
rect 699 2462 705 2463
rect 762 2463 763 2464
rect 767 2463 768 2467
rect 795 2465 796 2469
rect 800 2465 801 2469
rect 1326 2468 1327 2472
rect 1331 2468 1332 2472
rect 883 2467 889 2468
rect 883 2466 884 2467
rect 795 2464 801 2465
rect 816 2464 884 2466
rect 762 2462 768 2463
rect 816 2458 818 2464
rect 883 2463 884 2464
rect 888 2463 889 2467
rect 971 2467 977 2468
rect 971 2466 972 2467
rect 883 2462 889 2463
rect 936 2464 972 2466
rect 936 2458 938 2464
rect 971 2463 972 2464
rect 976 2463 977 2467
rect 1067 2467 1073 2468
rect 1067 2466 1068 2467
rect 971 2462 977 2463
rect 992 2464 1068 2466
rect 812 2456 818 2458
rect 900 2456 938 2458
rect 812 2454 814 2456
rect 900 2454 902 2456
rect 992 2454 994 2464
rect 1067 2463 1068 2464
rect 1072 2463 1073 2467
rect 1163 2467 1169 2468
rect 1326 2467 1332 2468
rect 1366 2471 1372 2472
rect 1366 2467 1367 2471
rect 1371 2467 1372 2471
rect 1163 2466 1164 2467
rect 1067 2462 1073 2463
rect 1159 2464 1164 2466
rect 1159 2458 1161 2464
rect 1163 2463 1164 2464
rect 1168 2463 1169 2467
rect 1366 2466 1372 2467
rect 1387 2471 1393 2472
rect 1387 2467 1388 2471
rect 1392 2470 1393 2471
rect 1438 2471 1444 2472
rect 1392 2468 1434 2470
rect 1392 2467 1393 2468
rect 1387 2466 1393 2467
rect 1163 2462 1169 2463
rect 1084 2456 1161 2458
rect 1432 2458 1434 2468
rect 1438 2467 1439 2471
rect 1443 2467 1444 2471
rect 1438 2466 1444 2467
rect 1459 2471 1465 2472
rect 1459 2467 1460 2471
rect 1464 2470 1465 2471
rect 1526 2471 1532 2472
rect 1464 2468 1522 2470
rect 1464 2467 1465 2468
rect 1459 2466 1465 2467
rect 1520 2458 1522 2468
rect 1526 2467 1527 2471
rect 1531 2467 1532 2471
rect 1526 2466 1532 2467
rect 1547 2471 1553 2472
rect 1547 2467 1548 2471
rect 1552 2470 1553 2471
rect 1614 2471 1620 2472
rect 1552 2468 1594 2470
rect 1552 2467 1553 2468
rect 1547 2466 1553 2467
rect 1592 2458 1594 2468
rect 1614 2467 1615 2471
rect 1619 2467 1620 2471
rect 1614 2466 1620 2467
rect 1635 2471 1641 2472
rect 1635 2467 1636 2471
rect 1640 2470 1641 2471
rect 1702 2471 1708 2472
rect 1640 2468 1698 2470
rect 1640 2467 1641 2468
rect 1635 2466 1641 2467
rect 1696 2458 1698 2468
rect 1702 2467 1703 2471
rect 1707 2467 1708 2471
rect 1702 2466 1708 2467
rect 1710 2471 1716 2472
rect 1710 2467 1711 2471
rect 1715 2470 1716 2471
rect 1723 2471 1729 2472
rect 1723 2470 1724 2471
rect 1715 2468 1724 2470
rect 1715 2467 1716 2468
rect 1710 2466 1716 2467
rect 1723 2467 1724 2468
rect 1728 2467 1729 2471
rect 1723 2466 1729 2467
rect 1790 2471 1796 2472
rect 1790 2467 1791 2471
rect 1795 2467 1796 2471
rect 1790 2466 1796 2467
rect 1811 2471 1817 2472
rect 1811 2467 1812 2471
rect 1816 2470 1817 2471
rect 1878 2471 1884 2472
rect 1816 2468 1874 2470
rect 1816 2467 1817 2468
rect 1811 2466 1817 2467
rect 1872 2458 1874 2468
rect 1878 2467 1879 2471
rect 1883 2467 1884 2471
rect 1878 2466 1884 2467
rect 1899 2471 1905 2472
rect 1899 2467 1900 2471
rect 1904 2470 1905 2471
rect 1966 2471 1972 2472
rect 1904 2468 1946 2470
rect 1904 2467 1905 2468
rect 1899 2466 1905 2467
rect 1944 2458 1946 2468
rect 1966 2467 1967 2471
rect 1971 2467 1972 2471
rect 1966 2466 1972 2467
rect 1987 2471 1993 2472
rect 1987 2467 1988 2471
rect 1992 2470 1993 2471
rect 2054 2471 2060 2472
rect 1992 2468 2001 2470
rect 1992 2467 1993 2468
rect 1987 2466 1993 2467
rect 1999 2458 2001 2468
rect 2054 2467 2055 2471
rect 2059 2467 2060 2471
rect 2054 2466 2060 2467
rect 2075 2471 2081 2472
rect 2075 2467 2076 2471
rect 2080 2470 2081 2471
rect 2142 2471 2148 2472
rect 2080 2468 2134 2470
rect 2080 2467 2081 2468
rect 2075 2466 2081 2467
rect 2132 2458 2134 2468
rect 2142 2467 2143 2471
rect 2147 2467 2148 2471
rect 2142 2466 2148 2467
rect 2150 2471 2156 2472
rect 2150 2467 2151 2471
rect 2155 2470 2156 2471
rect 2163 2471 2169 2472
rect 2163 2470 2164 2471
rect 2155 2468 2164 2470
rect 2155 2467 2156 2468
rect 2150 2466 2156 2467
rect 2163 2467 2164 2468
rect 2168 2467 2169 2471
rect 2502 2468 2503 2472
rect 2507 2468 2508 2472
rect 2502 2467 2508 2468
rect 2163 2466 2169 2467
rect 1432 2457 1449 2458
rect 1432 2456 1444 2457
rect 1084 2454 1086 2456
rect 1371 2455 1377 2456
rect 182 2453 188 2454
rect 110 2452 116 2453
rect 110 2448 111 2452
rect 115 2448 116 2452
rect 182 2449 183 2453
rect 187 2449 188 2453
rect 246 2453 252 2454
rect 182 2448 188 2449
rect 190 2451 196 2452
rect 110 2447 116 2448
rect 190 2447 191 2451
rect 195 2450 196 2451
rect 203 2451 209 2452
rect 203 2450 204 2451
rect 195 2448 204 2450
rect 195 2447 196 2448
rect 190 2446 196 2447
rect 203 2447 204 2448
rect 208 2447 209 2451
rect 246 2449 247 2453
rect 251 2449 252 2453
rect 246 2448 252 2449
rect 267 2453 321 2454
rect 267 2449 268 2453
rect 272 2452 321 2453
rect 326 2453 332 2454
rect 272 2449 273 2452
rect 267 2448 273 2449
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 347 2453 354 2454
rect 347 2449 348 2453
rect 352 2452 354 2453
rect 414 2453 420 2454
rect 352 2449 353 2452
rect 347 2448 353 2449
rect 414 2449 415 2453
rect 419 2449 420 2453
rect 502 2453 508 2454
rect 414 2448 420 2449
rect 434 2451 441 2452
rect 203 2446 209 2447
rect 434 2447 435 2451
rect 440 2447 441 2451
rect 502 2449 503 2453
rect 507 2449 508 2453
rect 502 2448 508 2449
rect 523 2453 529 2454
rect 523 2449 524 2453
rect 528 2449 529 2453
rect 523 2448 529 2449
rect 598 2453 604 2454
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 694 2453 700 2454
rect 598 2448 604 2449
rect 619 2451 628 2452
rect 434 2446 441 2447
rect 619 2447 620 2451
rect 627 2447 628 2451
rect 694 2449 695 2453
rect 699 2449 700 2453
rect 790 2453 796 2454
rect 694 2448 700 2449
rect 714 2451 721 2452
rect 619 2446 628 2447
rect 714 2447 715 2451
rect 720 2447 721 2451
rect 790 2449 791 2453
rect 795 2449 796 2453
rect 790 2448 796 2449
rect 811 2453 817 2454
rect 811 2449 812 2453
rect 816 2449 817 2453
rect 811 2448 817 2449
rect 878 2453 884 2454
rect 878 2449 879 2453
rect 883 2449 884 2453
rect 878 2448 884 2449
rect 899 2453 905 2454
rect 899 2449 900 2453
rect 904 2449 905 2453
rect 899 2448 905 2449
rect 966 2453 972 2454
rect 966 2449 967 2453
rect 971 2449 972 2453
rect 966 2448 972 2449
rect 987 2453 994 2454
rect 987 2449 988 2453
rect 992 2452 994 2453
rect 1062 2453 1068 2454
rect 992 2449 993 2452
rect 987 2448 993 2449
rect 1062 2449 1063 2453
rect 1067 2449 1068 2453
rect 1062 2448 1068 2449
rect 1083 2453 1089 2454
rect 1083 2449 1084 2453
rect 1088 2449 1089 2453
rect 1083 2448 1089 2449
rect 1158 2453 1164 2454
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1286 2452 1292 2453
rect 1158 2448 1164 2449
rect 1179 2451 1188 2452
rect 714 2446 721 2447
rect 1179 2447 1180 2451
rect 1187 2447 1188 2451
rect 1286 2448 1287 2452
rect 1291 2448 1292 2452
rect 1371 2451 1372 2455
rect 1376 2454 1377 2455
rect 1376 2452 1438 2454
rect 1443 2453 1444 2456
rect 1448 2453 1449 2457
rect 1520 2457 1537 2458
rect 1520 2456 1532 2457
rect 1443 2452 1449 2453
rect 1531 2453 1532 2456
rect 1536 2453 1537 2457
rect 1592 2457 1625 2458
rect 1592 2456 1620 2457
rect 1531 2452 1537 2453
rect 1619 2453 1620 2456
rect 1624 2453 1625 2457
rect 1696 2457 1713 2458
rect 1696 2456 1708 2457
rect 1619 2452 1625 2453
rect 1707 2453 1708 2456
rect 1712 2453 1713 2457
rect 1872 2457 1889 2458
rect 1872 2456 1884 2457
rect 1707 2452 1713 2453
rect 1795 2455 1804 2456
rect 1376 2451 1377 2452
rect 1371 2450 1377 2451
rect 1436 2450 1438 2452
rect 1658 2451 1664 2452
rect 1658 2450 1659 2451
rect 1436 2448 1659 2450
rect 1286 2447 1292 2448
rect 1658 2447 1659 2448
rect 1663 2447 1664 2451
rect 1795 2451 1796 2455
rect 1803 2451 1804 2455
rect 1883 2453 1884 2456
rect 1888 2453 1889 2457
rect 1944 2457 1977 2458
rect 1944 2456 1972 2457
rect 1883 2452 1889 2453
rect 1971 2453 1972 2456
rect 1976 2453 1977 2457
rect 1999 2457 2065 2458
rect 1999 2456 2060 2457
rect 1971 2452 1977 2453
rect 2059 2453 2060 2456
rect 2064 2453 2065 2457
rect 2132 2457 2153 2458
rect 2132 2456 2148 2457
rect 2059 2452 2065 2453
rect 2147 2453 2148 2456
rect 2152 2453 2153 2457
rect 2147 2452 2153 2453
rect 1795 2450 1804 2451
rect 1179 2446 1188 2447
rect 1658 2446 1664 2447
rect 110 2435 116 2436
rect 110 2431 111 2435
rect 115 2431 116 2435
rect 1286 2435 1292 2436
rect 110 2430 116 2431
rect 166 2432 172 2433
rect 166 2428 167 2432
rect 171 2428 172 2432
rect 166 2427 172 2428
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 486 2432 492 2433
rect 486 2428 487 2432
rect 491 2428 492 2432
rect 486 2427 492 2428
rect 582 2432 588 2433
rect 582 2428 583 2432
rect 587 2428 588 2432
rect 582 2427 588 2428
rect 678 2432 684 2433
rect 678 2428 679 2432
rect 683 2428 684 2432
rect 678 2427 684 2428
rect 774 2432 780 2433
rect 774 2428 775 2432
rect 779 2428 780 2432
rect 774 2427 780 2428
rect 862 2432 868 2433
rect 862 2428 863 2432
rect 867 2428 868 2432
rect 862 2427 868 2428
rect 950 2432 956 2433
rect 950 2428 951 2432
rect 955 2428 956 2432
rect 950 2427 956 2428
rect 1046 2432 1052 2433
rect 1046 2428 1047 2432
rect 1051 2428 1052 2432
rect 1046 2427 1052 2428
rect 1142 2432 1148 2433
rect 1142 2428 1143 2432
rect 1147 2428 1148 2432
rect 1286 2431 1287 2435
rect 1291 2431 1292 2435
rect 1286 2430 1292 2431
rect 1142 2427 1148 2428
rect 1371 2427 1380 2428
rect 1371 2423 1372 2427
rect 1379 2423 1380 2427
rect 1443 2427 1449 2428
rect 1443 2426 1444 2427
rect 1371 2422 1380 2423
rect 1388 2424 1444 2426
rect 150 2416 156 2417
rect 110 2413 116 2414
rect 110 2409 111 2413
rect 115 2409 116 2413
rect 150 2412 151 2416
rect 155 2412 156 2416
rect 150 2411 156 2412
rect 230 2416 236 2417
rect 230 2412 231 2416
rect 235 2412 236 2416
rect 230 2411 236 2412
rect 318 2416 324 2417
rect 318 2412 319 2416
rect 323 2412 324 2416
rect 318 2411 324 2412
rect 414 2416 420 2417
rect 414 2412 415 2416
rect 419 2412 420 2416
rect 414 2411 420 2412
rect 518 2416 524 2417
rect 518 2412 519 2416
rect 523 2412 524 2416
rect 518 2411 524 2412
rect 622 2416 628 2417
rect 622 2412 623 2416
rect 627 2412 628 2416
rect 622 2411 628 2412
rect 726 2416 732 2417
rect 726 2412 727 2416
rect 731 2412 732 2416
rect 726 2411 732 2412
rect 830 2416 836 2417
rect 830 2412 831 2416
rect 835 2412 836 2416
rect 830 2411 836 2412
rect 934 2416 940 2417
rect 934 2412 935 2416
rect 939 2412 940 2416
rect 934 2411 940 2412
rect 1038 2416 1044 2417
rect 1038 2412 1039 2416
rect 1043 2412 1044 2416
rect 1038 2411 1044 2412
rect 1150 2416 1156 2417
rect 1150 2412 1151 2416
rect 1155 2412 1156 2416
rect 1388 2414 1390 2424
rect 1443 2423 1444 2424
rect 1448 2423 1449 2427
rect 1547 2427 1553 2428
rect 1547 2426 1548 2427
rect 1443 2422 1449 2423
rect 1460 2424 1548 2426
rect 1460 2414 1462 2424
rect 1547 2423 1548 2424
rect 1552 2423 1553 2427
rect 1643 2427 1649 2428
rect 1643 2426 1644 2427
rect 1547 2422 1553 2423
rect 1564 2424 1644 2426
rect 1564 2414 1566 2424
rect 1643 2423 1644 2424
rect 1648 2423 1649 2427
rect 1643 2422 1649 2423
rect 1739 2427 1745 2428
rect 1739 2423 1740 2427
rect 1744 2426 1745 2427
rect 1827 2427 1833 2428
rect 1744 2424 1814 2426
rect 1744 2423 1745 2424
rect 1739 2422 1745 2423
rect 1812 2418 1814 2424
rect 1827 2423 1828 2427
rect 1832 2426 1833 2427
rect 1915 2427 1921 2428
rect 1832 2424 1910 2426
rect 1832 2423 1833 2424
rect 1827 2422 1833 2423
rect 1908 2418 1910 2424
rect 1915 2423 1916 2427
rect 1920 2426 1921 2427
rect 2011 2427 2017 2428
rect 1920 2424 2001 2426
rect 1920 2423 1921 2424
rect 1915 2422 1921 2423
rect 1999 2418 2001 2424
rect 2011 2423 2012 2427
rect 2016 2426 2017 2427
rect 2107 2427 2113 2428
rect 2016 2424 2102 2426
rect 2016 2423 2017 2424
rect 2011 2422 2017 2423
rect 2100 2418 2102 2424
rect 2107 2423 2108 2427
rect 2112 2426 2113 2427
rect 2150 2427 2156 2428
rect 2150 2426 2151 2427
rect 2112 2424 2151 2426
rect 2112 2423 2113 2424
rect 2107 2422 2113 2423
rect 2150 2423 2151 2424
rect 2155 2423 2156 2427
rect 2150 2422 2156 2423
rect 1812 2416 1846 2418
rect 1908 2416 1934 2418
rect 1999 2416 2030 2418
rect 2100 2416 2126 2418
rect 1844 2414 1846 2416
rect 1932 2414 1934 2416
rect 2028 2414 2030 2416
rect 2124 2414 2126 2416
rect 1150 2411 1156 2412
rect 1286 2413 1292 2414
rect 1366 2413 1372 2414
rect 110 2408 116 2409
rect 1286 2409 1287 2413
rect 1291 2409 1292 2413
rect 1286 2408 1292 2409
rect 1326 2412 1332 2413
rect 1326 2408 1327 2412
rect 1331 2408 1332 2412
rect 1366 2409 1367 2413
rect 1371 2409 1372 2413
rect 1366 2408 1372 2409
rect 1387 2413 1393 2414
rect 1387 2409 1388 2413
rect 1392 2409 1393 2413
rect 1387 2408 1393 2409
rect 1438 2413 1444 2414
rect 1438 2409 1439 2413
rect 1443 2409 1444 2413
rect 1438 2408 1444 2409
rect 1459 2413 1465 2414
rect 1459 2409 1460 2413
rect 1464 2409 1465 2413
rect 1459 2408 1465 2409
rect 1542 2413 1548 2414
rect 1542 2409 1543 2413
rect 1547 2409 1548 2413
rect 1542 2408 1548 2409
rect 1563 2413 1569 2414
rect 1563 2409 1564 2413
rect 1568 2409 1569 2413
rect 1563 2408 1569 2409
rect 1638 2413 1644 2414
rect 1638 2409 1639 2413
rect 1643 2409 1644 2413
rect 1734 2413 1740 2414
rect 1638 2408 1644 2409
rect 1658 2411 1665 2412
rect 1326 2407 1332 2408
rect 1658 2407 1659 2411
rect 1664 2407 1665 2411
rect 1734 2409 1735 2413
rect 1739 2409 1740 2413
rect 1822 2413 1828 2414
rect 1734 2408 1740 2409
rect 1755 2411 1764 2412
rect 1658 2406 1665 2407
rect 1755 2407 1756 2411
rect 1763 2407 1764 2411
rect 1822 2409 1823 2413
rect 1827 2409 1828 2413
rect 1822 2408 1828 2409
rect 1843 2413 1849 2414
rect 1843 2409 1844 2413
rect 1848 2409 1849 2413
rect 1843 2408 1849 2409
rect 1910 2413 1916 2414
rect 1910 2409 1911 2413
rect 1915 2409 1916 2413
rect 1910 2408 1916 2409
rect 1931 2413 1937 2414
rect 1931 2409 1932 2413
rect 1936 2409 1937 2413
rect 1931 2408 1937 2409
rect 2006 2413 2012 2414
rect 2006 2409 2007 2413
rect 2011 2409 2012 2413
rect 2006 2408 2012 2409
rect 2027 2413 2033 2414
rect 2027 2409 2028 2413
rect 2032 2409 2033 2413
rect 2027 2408 2033 2409
rect 2102 2413 2108 2414
rect 2102 2409 2103 2413
rect 2107 2409 2108 2413
rect 2102 2408 2108 2409
rect 2123 2413 2129 2414
rect 2123 2409 2124 2413
rect 2128 2409 2129 2413
rect 2123 2408 2129 2409
rect 2502 2412 2508 2413
rect 2502 2408 2503 2412
rect 2507 2408 2508 2412
rect 2502 2407 2508 2408
rect 1755 2406 1764 2407
rect 110 2396 116 2397
rect 1286 2396 1292 2397
rect 110 2392 111 2396
rect 115 2392 116 2396
rect 110 2391 116 2392
rect 166 2395 172 2396
rect 166 2391 167 2395
rect 171 2391 172 2395
rect 166 2390 172 2391
rect 187 2395 193 2396
rect 187 2391 188 2395
rect 192 2394 193 2395
rect 246 2395 252 2396
rect 192 2392 230 2394
rect 192 2391 193 2392
rect 187 2390 193 2391
rect 228 2382 230 2392
rect 246 2391 247 2395
rect 251 2391 252 2395
rect 246 2390 252 2391
rect 267 2395 273 2396
rect 267 2391 268 2395
rect 272 2394 273 2395
rect 334 2395 340 2396
rect 272 2392 321 2394
rect 272 2391 273 2392
rect 267 2390 273 2391
rect 319 2382 321 2392
rect 334 2391 335 2395
rect 339 2391 340 2395
rect 334 2390 340 2391
rect 355 2395 361 2396
rect 355 2391 356 2395
rect 360 2394 361 2395
rect 430 2395 436 2396
rect 360 2392 426 2394
rect 360 2391 361 2392
rect 355 2390 361 2391
rect 424 2382 426 2392
rect 430 2391 431 2395
rect 435 2391 436 2395
rect 430 2390 436 2391
rect 438 2395 444 2396
rect 438 2391 439 2395
rect 443 2394 444 2395
rect 451 2395 457 2396
rect 451 2394 452 2395
rect 443 2392 452 2394
rect 443 2391 444 2392
rect 438 2390 444 2391
rect 451 2391 452 2392
rect 456 2391 457 2395
rect 451 2390 457 2391
rect 534 2395 540 2396
rect 534 2391 535 2395
rect 539 2391 540 2395
rect 534 2390 540 2391
rect 555 2395 561 2396
rect 555 2391 556 2395
rect 560 2394 561 2395
rect 638 2395 644 2396
rect 560 2392 630 2394
rect 560 2391 561 2392
rect 555 2390 561 2391
rect 628 2382 630 2392
rect 638 2391 639 2395
rect 643 2391 644 2395
rect 638 2390 644 2391
rect 659 2395 665 2396
rect 659 2391 660 2395
rect 664 2394 665 2395
rect 742 2395 748 2396
rect 664 2392 738 2394
rect 664 2391 665 2392
rect 659 2390 665 2391
rect 736 2382 738 2392
rect 742 2391 743 2395
rect 747 2391 748 2395
rect 742 2390 748 2391
rect 762 2395 769 2396
rect 762 2391 763 2395
rect 768 2391 769 2395
rect 762 2390 769 2391
rect 846 2395 852 2396
rect 846 2391 847 2395
rect 851 2391 852 2395
rect 846 2390 852 2391
rect 867 2395 873 2396
rect 867 2391 868 2395
rect 872 2391 873 2395
rect 867 2390 873 2391
rect 950 2395 956 2396
rect 950 2391 951 2395
rect 955 2391 956 2395
rect 950 2390 956 2391
rect 971 2395 977 2396
rect 971 2391 972 2395
rect 976 2394 977 2395
rect 1054 2395 1060 2396
rect 976 2392 1050 2394
rect 976 2391 977 2392
rect 971 2390 977 2391
rect 869 2382 871 2390
rect 1048 2382 1050 2392
rect 1054 2391 1055 2395
rect 1059 2391 1060 2395
rect 1054 2390 1060 2391
rect 1075 2395 1081 2396
rect 1075 2391 1076 2395
rect 1080 2394 1081 2395
rect 1166 2395 1172 2396
rect 1080 2392 1161 2394
rect 1080 2391 1081 2392
rect 1075 2390 1081 2391
rect 1159 2382 1161 2392
rect 1166 2391 1167 2395
rect 1171 2391 1172 2395
rect 1166 2390 1172 2391
rect 1174 2395 1180 2396
rect 1174 2391 1175 2395
rect 1179 2394 1180 2395
rect 1187 2395 1193 2396
rect 1187 2394 1188 2395
rect 1179 2392 1188 2394
rect 1179 2391 1180 2392
rect 1174 2390 1180 2391
rect 1187 2391 1188 2392
rect 1192 2391 1193 2395
rect 1286 2392 1287 2396
rect 1291 2392 1292 2396
rect 1286 2391 1292 2392
rect 1326 2395 1332 2396
rect 1326 2391 1327 2395
rect 1331 2391 1332 2395
rect 2502 2395 2508 2396
rect 1187 2390 1193 2391
rect 1326 2390 1332 2391
rect 1350 2392 1356 2393
rect 1350 2388 1351 2392
rect 1355 2388 1356 2392
rect 1350 2387 1356 2388
rect 1422 2392 1428 2393
rect 1422 2388 1423 2392
rect 1427 2388 1428 2392
rect 1422 2387 1428 2388
rect 1526 2392 1532 2393
rect 1526 2388 1527 2392
rect 1531 2388 1532 2392
rect 1526 2387 1532 2388
rect 1622 2392 1628 2393
rect 1622 2388 1623 2392
rect 1627 2388 1628 2392
rect 1622 2387 1628 2388
rect 1718 2392 1724 2393
rect 1718 2388 1719 2392
rect 1723 2388 1724 2392
rect 1718 2387 1724 2388
rect 1806 2392 1812 2393
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1894 2392 1900 2393
rect 1894 2388 1895 2392
rect 1899 2388 1900 2392
rect 1894 2387 1900 2388
rect 1990 2392 1996 2393
rect 1990 2388 1991 2392
rect 1995 2388 1996 2392
rect 1990 2387 1996 2388
rect 2086 2392 2092 2393
rect 2086 2388 2087 2392
rect 2091 2388 2092 2392
rect 2502 2391 2503 2395
rect 2507 2391 2508 2395
rect 2502 2390 2508 2391
rect 2086 2387 2092 2388
rect 228 2381 257 2382
rect 228 2380 252 2381
rect 171 2379 177 2380
rect 171 2375 172 2379
rect 176 2378 177 2379
rect 190 2379 196 2380
rect 190 2378 191 2379
rect 176 2376 191 2378
rect 176 2375 177 2376
rect 171 2374 177 2375
rect 190 2375 191 2376
rect 195 2375 196 2379
rect 251 2377 252 2380
rect 256 2377 257 2381
rect 319 2381 345 2382
rect 319 2380 340 2381
rect 251 2376 257 2377
rect 339 2377 340 2380
rect 344 2377 345 2381
rect 424 2381 441 2382
rect 424 2380 436 2381
rect 339 2376 345 2377
rect 435 2377 436 2380
rect 440 2377 441 2381
rect 628 2381 649 2382
rect 628 2380 644 2381
rect 435 2376 441 2377
rect 539 2379 545 2380
rect 190 2374 196 2375
rect 539 2375 540 2379
rect 544 2378 545 2379
rect 544 2376 630 2378
rect 643 2377 644 2380
rect 648 2377 649 2381
rect 736 2381 753 2382
rect 736 2380 748 2381
rect 643 2376 649 2377
rect 747 2377 748 2380
rect 752 2377 753 2381
rect 869 2381 961 2382
rect 869 2380 956 2381
rect 747 2376 753 2377
rect 851 2379 857 2380
rect 544 2375 545 2376
rect 539 2374 545 2375
rect 628 2375 636 2376
rect 628 2372 631 2375
rect 630 2371 631 2372
rect 635 2371 636 2375
rect 851 2375 852 2379
rect 856 2378 857 2379
rect 856 2376 950 2378
rect 955 2377 956 2380
rect 960 2377 961 2381
rect 1048 2381 1065 2382
rect 1048 2380 1060 2381
rect 955 2376 961 2377
rect 1059 2377 1060 2380
rect 1064 2377 1065 2381
rect 1159 2381 1177 2382
rect 1159 2380 1172 2381
rect 1059 2376 1065 2377
rect 1171 2377 1172 2380
rect 1176 2377 1177 2381
rect 1171 2376 1177 2377
rect 856 2375 857 2376
rect 851 2374 857 2375
rect 948 2374 950 2376
rect 1182 2375 1188 2376
rect 1182 2374 1183 2375
rect 948 2372 1183 2374
rect 630 2370 636 2371
rect 1182 2371 1183 2372
rect 1187 2371 1188 2375
rect 1182 2370 1188 2371
rect 1350 2372 1356 2373
rect 1326 2369 1332 2370
rect 438 2367 444 2368
rect 438 2366 439 2367
rect 180 2364 439 2366
rect 180 2362 182 2364
rect 438 2363 439 2364
rect 443 2363 444 2367
rect 1146 2367 1152 2368
rect 1146 2366 1147 2367
rect 438 2362 444 2363
rect 876 2364 1147 2366
rect 876 2362 878 2364
rect 1146 2363 1147 2364
rect 1151 2363 1152 2367
rect 1326 2365 1327 2369
rect 1331 2365 1332 2369
rect 1350 2368 1351 2372
rect 1355 2368 1356 2372
rect 1350 2367 1356 2368
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1494 2372 1500 2373
rect 1494 2368 1495 2372
rect 1499 2368 1500 2372
rect 1494 2367 1500 2368
rect 1582 2372 1588 2373
rect 1582 2368 1583 2372
rect 1587 2368 1588 2372
rect 1582 2367 1588 2368
rect 1670 2372 1676 2373
rect 1670 2368 1671 2372
rect 1675 2368 1676 2372
rect 1670 2367 1676 2368
rect 1750 2372 1756 2373
rect 1750 2368 1751 2372
rect 1755 2368 1756 2372
rect 1750 2367 1756 2368
rect 1830 2372 1836 2373
rect 1830 2368 1831 2372
rect 1835 2368 1836 2372
rect 1830 2367 1836 2368
rect 1918 2372 1924 2373
rect 1918 2368 1919 2372
rect 1923 2368 1924 2372
rect 1918 2367 1924 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2094 2372 2100 2373
rect 2094 2368 2095 2372
rect 2099 2368 2100 2372
rect 2094 2367 2100 2368
rect 2502 2369 2508 2370
rect 1326 2364 1332 2365
rect 2502 2365 2503 2369
rect 2507 2365 2508 2369
rect 2502 2364 2508 2365
rect 1146 2362 1152 2363
rect 179 2361 185 2362
rect 179 2357 180 2361
rect 184 2357 185 2361
rect 875 2361 881 2362
rect 283 2359 289 2360
rect 283 2358 284 2359
rect 179 2356 185 2357
rect 196 2356 284 2358
rect 196 2346 198 2356
rect 283 2355 284 2356
rect 288 2355 289 2359
rect 395 2359 401 2360
rect 395 2358 396 2359
rect 283 2354 289 2355
rect 319 2356 396 2358
rect 319 2350 321 2356
rect 395 2355 396 2356
rect 400 2355 401 2359
rect 507 2359 513 2360
rect 507 2358 508 2359
rect 395 2354 401 2355
rect 412 2356 508 2358
rect 300 2348 321 2350
rect 300 2346 302 2348
rect 412 2346 414 2356
rect 507 2355 508 2356
rect 512 2355 513 2359
rect 507 2354 513 2355
rect 627 2359 633 2360
rect 627 2355 628 2359
rect 632 2358 633 2359
rect 747 2359 753 2360
rect 632 2356 742 2358
rect 632 2355 633 2356
rect 627 2354 633 2355
rect 740 2350 742 2356
rect 747 2355 748 2359
rect 752 2358 753 2359
rect 770 2359 776 2360
rect 770 2358 771 2359
rect 752 2356 771 2358
rect 752 2355 753 2356
rect 747 2354 753 2355
rect 770 2355 771 2356
rect 775 2355 776 2359
rect 875 2357 876 2361
rect 880 2357 881 2361
rect 1003 2359 1009 2360
rect 1003 2358 1004 2359
rect 875 2356 881 2357
rect 892 2356 1004 2358
rect 770 2354 776 2355
rect 740 2348 766 2350
rect 764 2346 766 2348
rect 892 2346 894 2356
rect 1003 2355 1004 2356
rect 1008 2355 1009 2359
rect 1003 2354 1009 2355
rect 1131 2359 1137 2360
rect 1131 2355 1132 2359
rect 1136 2358 1137 2359
rect 1174 2359 1180 2360
rect 1174 2358 1175 2359
rect 1136 2356 1175 2358
rect 1136 2355 1137 2356
rect 1131 2354 1137 2355
rect 1174 2355 1175 2356
rect 1179 2355 1180 2359
rect 1174 2354 1180 2355
rect 1326 2352 1332 2353
rect 2502 2352 2508 2353
rect 1326 2348 1327 2352
rect 1331 2348 1332 2352
rect 1326 2347 1332 2348
rect 1366 2351 1372 2352
rect 1366 2347 1367 2351
rect 1371 2347 1372 2351
rect 1366 2346 1372 2347
rect 1374 2351 1380 2352
rect 1374 2347 1375 2351
rect 1379 2350 1380 2351
rect 1387 2351 1393 2352
rect 1387 2350 1388 2351
rect 1379 2348 1388 2350
rect 1379 2347 1380 2348
rect 1374 2346 1380 2347
rect 1387 2347 1388 2348
rect 1392 2347 1393 2351
rect 1387 2346 1393 2347
rect 1422 2351 1428 2352
rect 1422 2347 1423 2351
rect 1427 2347 1428 2351
rect 1443 2351 1449 2352
rect 1443 2350 1444 2351
rect 1422 2346 1428 2347
rect 1432 2348 1444 2350
rect 174 2345 180 2346
rect 110 2344 116 2345
rect 110 2340 111 2344
rect 115 2340 116 2344
rect 174 2341 175 2345
rect 179 2341 180 2345
rect 174 2340 180 2341
rect 195 2345 201 2346
rect 195 2341 196 2345
rect 200 2341 201 2345
rect 195 2340 201 2341
rect 278 2345 284 2346
rect 278 2341 279 2345
rect 283 2341 284 2345
rect 278 2340 284 2341
rect 299 2345 305 2346
rect 299 2341 300 2345
rect 304 2341 305 2345
rect 299 2340 305 2341
rect 390 2345 396 2346
rect 390 2341 391 2345
rect 395 2341 396 2345
rect 390 2340 396 2341
rect 411 2345 417 2346
rect 411 2341 412 2345
rect 416 2341 417 2345
rect 411 2340 417 2341
rect 502 2345 508 2346
rect 502 2341 503 2345
rect 507 2341 508 2345
rect 622 2345 628 2346
rect 502 2340 508 2341
rect 510 2343 516 2344
rect 110 2339 116 2340
rect 510 2339 511 2343
rect 515 2342 516 2343
rect 523 2343 529 2344
rect 523 2342 524 2343
rect 515 2340 524 2342
rect 515 2339 516 2340
rect 510 2338 516 2339
rect 523 2339 524 2340
rect 528 2339 529 2343
rect 622 2341 623 2345
rect 627 2341 628 2345
rect 742 2345 748 2346
rect 622 2340 628 2341
rect 630 2343 636 2344
rect 523 2338 529 2339
rect 630 2339 631 2343
rect 635 2342 636 2343
rect 643 2343 649 2344
rect 643 2342 644 2343
rect 635 2340 644 2342
rect 635 2339 636 2340
rect 630 2338 636 2339
rect 643 2339 644 2340
rect 648 2339 649 2343
rect 742 2341 743 2345
rect 747 2341 748 2345
rect 742 2340 748 2341
rect 763 2345 769 2346
rect 763 2341 764 2345
rect 768 2341 769 2345
rect 763 2340 769 2341
rect 870 2345 876 2346
rect 870 2341 871 2345
rect 875 2341 876 2345
rect 870 2340 876 2341
rect 891 2345 897 2346
rect 891 2341 892 2345
rect 896 2341 897 2345
rect 891 2340 897 2341
rect 998 2345 1004 2346
rect 998 2341 999 2345
rect 1003 2341 1004 2345
rect 1126 2345 1132 2346
rect 998 2340 1004 2341
rect 1014 2343 1025 2344
rect 643 2338 649 2339
rect 1014 2339 1015 2343
rect 1019 2339 1020 2343
rect 1024 2339 1025 2343
rect 1126 2341 1127 2345
rect 1131 2341 1132 2345
rect 1286 2344 1292 2345
rect 1126 2340 1132 2341
rect 1146 2343 1153 2344
rect 1014 2338 1025 2339
rect 1146 2339 1147 2343
rect 1152 2339 1153 2343
rect 1286 2340 1287 2344
rect 1291 2340 1292 2344
rect 1432 2342 1434 2348
rect 1443 2347 1444 2348
rect 1448 2347 1449 2351
rect 1443 2346 1449 2347
rect 1510 2351 1516 2352
rect 1510 2347 1511 2351
rect 1515 2347 1516 2351
rect 1531 2351 1537 2352
rect 1531 2350 1532 2351
rect 1510 2346 1516 2347
rect 1520 2348 1532 2350
rect 1520 2342 1522 2348
rect 1531 2347 1532 2348
rect 1536 2347 1537 2351
rect 1531 2346 1537 2347
rect 1598 2351 1604 2352
rect 1598 2347 1599 2351
rect 1603 2347 1604 2351
rect 1598 2346 1604 2347
rect 1619 2351 1625 2352
rect 1619 2347 1620 2351
rect 1624 2350 1625 2351
rect 1686 2351 1692 2352
rect 1624 2348 1678 2350
rect 1624 2347 1625 2348
rect 1619 2346 1625 2347
rect 1286 2339 1292 2340
rect 1372 2340 1434 2342
rect 1436 2340 1522 2342
rect 1146 2338 1153 2339
rect 1372 2338 1374 2340
rect 1436 2338 1438 2340
rect 1371 2337 1377 2338
rect 1371 2333 1372 2337
rect 1376 2333 1377 2337
rect 1371 2332 1377 2333
rect 1427 2337 1438 2338
rect 1427 2333 1428 2337
rect 1432 2336 1438 2337
rect 1676 2338 1678 2348
rect 1686 2347 1687 2351
rect 1691 2347 1692 2351
rect 1686 2346 1692 2347
rect 1694 2351 1700 2352
rect 1694 2347 1695 2351
rect 1699 2350 1700 2351
rect 1707 2351 1713 2352
rect 1707 2350 1708 2351
rect 1699 2348 1708 2350
rect 1699 2347 1700 2348
rect 1694 2346 1700 2347
rect 1707 2347 1708 2348
rect 1712 2347 1713 2351
rect 1707 2346 1713 2347
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2347 1772 2351
rect 1766 2346 1772 2347
rect 1787 2351 1793 2352
rect 1787 2347 1788 2351
rect 1792 2350 1793 2351
rect 1846 2351 1852 2352
rect 1792 2348 1842 2350
rect 1792 2347 1793 2348
rect 1787 2346 1793 2347
rect 1840 2338 1842 2348
rect 1846 2347 1847 2351
rect 1851 2347 1852 2351
rect 1846 2346 1852 2347
rect 1867 2351 1873 2352
rect 1867 2347 1868 2351
rect 1872 2350 1873 2351
rect 1934 2351 1940 2352
rect 1872 2348 1926 2350
rect 1872 2347 1873 2348
rect 1867 2346 1873 2347
rect 1924 2338 1926 2348
rect 1934 2347 1935 2351
rect 1939 2347 1940 2351
rect 1934 2346 1940 2347
rect 1955 2351 1961 2352
rect 1955 2347 1956 2351
rect 1960 2350 1961 2351
rect 2022 2351 2028 2352
rect 1960 2348 2001 2350
rect 1960 2347 1961 2348
rect 1955 2346 1961 2347
rect 1999 2338 2001 2348
rect 2022 2347 2023 2351
rect 2027 2347 2028 2351
rect 2022 2346 2028 2347
rect 2043 2351 2049 2352
rect 2043 2347 2044 2351
rect 2048 2350 2049 2351
rect 2110 2351 2116 2352
rect 2048 2348 2102 2350
rect 2048 2347 2049 2348
rect 2043 2346 2049 2347
rect 2100 2338 2102 2348
rect 2110 2347 2111 2351
rect 2115 2347 2116 2351
rect 2110 2346 2116 2347
rect 2118 2351 2124 2352
rect 2118 2347 2119 2351
rect 2123 2350 2124 2351
rect 2131 2351 2137 2352
rect 2131 2350 2132 2351
rect 2123 2348 2132 2350
rect 2123 2347 2124 2348
rect 2118 2346 2124 2347
rect 2131 2347 2132 2348
rect 2136 2347 2137 2351
rect 2502 2348 2503 2352
rect 2507 2348 2508 2352
rect 2502 2347 2508 2348
rect 2131 2346 2137 2347
rect 1676 2337 1697 2338
rect 1676 2336 1692 2337
rect 1432 2333 1433 2336
rect 1427 2332 1433 2333
rect 1515 2335 1521 2336
rect 1515 2331 1516 2335
rect 1520 2334 1521 2335
rect 1566 2335 1572 2336
rect 1520 2332 1562 2334
rect 1520 2331 1521 2332
rect 1515 2330 1521 2331
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 1286 2327 1292 2328
rect 110 2322 116 2323
rect 158 2324 164 2325
rect 158 2320 159 2324
rect 163 2320 164 2324
rect 158 2319 164 2320
rect 262 2324 268 2325
rect 262 2320 263 2324
rect 267 2320 268 2324
rect 262 2319 268 2320
rect 374 2324 380 2325
rect 374 2320 375 2324
rect 379 2320 380 2324
rect 374 2319 380 2320
rect 486 2324 492 2325
rect 486 2320 487 2324
rect 491 2320 492 2324
rect 486 2319 492 2320
rect 606 2324 612 2325
rect 606 2320 607 2324
rect 611 2320 612 2324
rect 606 2319 612 2320
rect 726 2324 732 2325
rect 726 2320 727 2324
rect 731 2320 732 2324
rect 726 2319 732 2320
rect 854 2324 860 2325
rect 854 2320 855 2324
rect 859 2320 860 2324
rect 854 2319 860 2320
rect 982 2324 988 2325
rect 982 2320 983 2324
rect 987 2320 988 2324
rect 982 2319 988 2320
rect 1110 2324 1116 2325
rect 1110 2320 1111 2324
rect 1115 2320 1116 2324
rect 1286 2323 1287 2327
rect 1291 2323 1292 2327
rect 1560 2326 1562 2332
rect 1566 2331 1567 2335
rect 1571 2334 1572 2335
rect 1603 2335 1609 2336
rect 1603 2334 1604 2335
rect 1571 2332 1604 2334
rect 1571 2331 1572 2332
rect 1566 2330 1572 2331
rect 1603 2331 1604 2332
rect 1608 2331 1609 2335
rect 1691 2333 1692 2336
rect 1696 2333 1697 2337
rect 1840 2337 1857 2338
rect 1840 2336 1852 2337
rect 1691 2332 1697 2333
rect 1758 2335 1764 2336
rect 1603 2330 1609 2331
rect 1758 2331 1759 2335
rect 1763 2334 1764 2335
rect 1771 2335 1777 2336
rect 1771 2334 1772 2335
rect 1763 2332 1772 2334
rect 1763 2331 1764 2332
rect 1758 2330 1764 2331
rect 1771 2331 1772 2332
rect 1776 2331 1777 2335
rect 1851 2333 1852 2336
rect 1856 2333 1857 2337
rect 1924 2337 1945 2338
rect 1924 2336 1940 2337
rect 1851 2332 1857 2333
rect 1939 2333 1940 2336
rect 1944 2333 1945 2337
rect 1999 2337 2033 2338
rect 1999 2336 2028 2337
rect 1939 2332 1945 2333
rect 2027 2333 2028 2336
rect 2032 2333 2033 2337
rect 2100 2337 2121 2338
rect 2100 2336 2116 2337
rect 2027 2332 2033 2333
rect 2115 2333 2116 2336
rect 2120 2333 2121 2337
rect 2115 2332 2121 2333
rect 1771 2330 1777 2331
rect 1694 2327 1700 2328
rect 1694 2326 1695 2327
rect 1560 2324 1695 2326
rect 1286 2322 1292 2323
rect 1694 2323 1695 2324
rect 1699 2323 1700 2327
rect 1694 2322 1700 2323
rect 1110 2319 1116 2320
rect 1658 2319 1664 2320
rect 1658 2318 1659 2319
rect 1372 2316 1659 2318
rect 1372 2314 1374 2316
rect 1658 2315 1659 2316
rect 1663 2315 1664 2319
rect 2118 2319 2124 2320
rect 2118 2318 2119 2319
rect 1658 2314 1664 2315
rect 1836 2316 2119 2318
rect 1836 2314 1838 2316
rect 2118 2315 2119 2316
rect 2123 2315 2124 2319
rect 2118 2314 2124 2315
rect 1371 2313 1377 2314
rect 1371 2309 1372 2313
rect 1376 2309 1377 2313
rect 1835 2313 1841 2314
rect 1459 2311 1465 2312
rect 1459 2310 1460 2311
rect 206 2308 212 2309
rect 110 2305 116 2306
rect 110 2301 111 2305
rect 115 2301 116 2305
rect 206 2304 207 2308
rect 211 2304 212 2308
rect 206 2303 212 2304
rect 286 2308 292 2309
rect 286 2304 287 2308
rect 291 2304 292 2308
rect 286 2303 292 2304
rect 374 2308 380 2309
rect 374 2304 375 2308
rect 379 2304 380 2308
rect 374 2303 380 2304
rect 470 2308 476 2309
rect 470 2304 471 2308
rect 475 2304 476 2308
rect 470 2303 476 2304
rect 558 2308 564 2309
rect 558 2304 559 2308
rect 563 2304 564 2308
rect 558 2303 564 2304
rect 646 2308 652 2309
rect 646 2304 647 2308
rect 651 2304 652 2308
rect 646 2303 652 2304
rect 734 2308 740 2309
rect 734 2304 735 2308
rect 739 2304 740 2308
rect 734 2303 740 2304
rect 814 2308 820 2309
rect 814 2304 815 2308
rect 819 2304 820 2308
rect 814 2303 820 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 990 2308 996 2309
rect 990 2304 991 2308
rect 995 2304 996 2308
rect 990 2303 996 2304
rect 1078 2308 1084 2309
rect 1371 2308 1377 2309
rect 1388 2308 1460 2310
rect 1078 2304 1079 2308
rect 1083 2304 1084 2308
rect 1078 2303 1084 2304
rect 1286 2305 1292 2306
rect 110 2300 116 2301
rect 1286 2301 1287 2305
rect 1291 2301 1292 2305
rect 1286 2300 1292 2301
rect 1388 2298 1390 2308
rect 1459 2307 1460 2308
rect 1464 2307 1465 2311
rect 1547 2311 1553 2312
rect 1547 2310 1548 2311
rect 1459 2306 1465 2307
rect 1476 2308 1548 2310
rect 1476 2298 1478 2308
rect 1547 2307 1548 2308
rect 1552 2307 1553 2311
rect 1547 2306 1553 2307
rect 1643 2311 1649 2312
rect 1643 2307 1644 2311
rect 1648 2310 1649 2311
rect 1739 2311 1745 2312
rect 1648 2308 1734 2310
rect 1648 2307 1649 2308
rect 1643 2306 1649 2307
rect 1732 2302 1734 2308
rect 1739 2307 1740 2311
rect 1744 2310 1745 2311
rect 1822 2311 1828 2312
rect 1822 2310 1823 2311
rect 1744 2308 1823 2310
rect 1744 2307 1745 2308
rect 1739 2306 1745 2307
rect 1822 2307 1823 2308
rect 1827 2307 1828 2311
rect 1835 2309 1836 2313
rect 1840 2309 1841 2313
rect 1931 2311 1937 2312
rect 1931 2310 1932 2311
rect 1835 2308 1841 2309
rect 1852 2308 1932 2310
rect 1822 2306 1828 2307
rect 1732 2300 1758 2302
rect 1756 2298 1758 2300
rect 1852 2298 1854 2308
rect 1931 2307 1932 2308
rect 1936 2307 1937 2311
rect 2019 2311 2025 2312
rect 2019 2310 2020 2311
rect 1931 2306 1937 2307
rect 1999 2308 2020 2310
rect 1999 2302 2001 2308
rect 2019 2307 2020 2308
rect 2024 2307 2025 2311
rect 2115 2311 2121 2312
rect 2115 2310 2116 2311
rect 2019 2306 2025 2307
rect 2036 2308 2116 2310
rect 1948 2300 2001 2302
rect 1948 2298 1950 2300
rect 2036 2298 2038 2308
rect 2115 2307 2116 2308
rect 2120 2307 2121 2311
rect 2211 2311 2217 2312
rect 2211 2310 2212 2311
rect 2115 2306 2121 2307
rect 2132 2308 2212 2310
rect 2132 2298 2134 2308
rect 2211 2307 2212 2308
rect 2216 2307 2217 2311
rect 2211 2306 2217 2307
rect 1366 2297 1372 2298
rect 1326 2296 1332 2297
rect 1326 2292 1327 2296
rect 1331 2292 1332 2296
rect 1366 2293 1367 2297
rect 1371 2293 1372 2297
rect 1366 2292 1372 2293
rect 1387 2297 1393 2298
rect 1387 2293 1388 2297
rect 1392 2293 1393 2297
rect 1387 2292 1393 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1475 2297 1481 2298
rect 1475 2293 1476 2297
rect 1480 2293 1481 2297
rect 1475 2292 1481 2293
rect 1542 2297 1548 2298
rect 1542 2293 1543 2297
rect 1547 2293 1548 2297
rect 1638 2297 1644 2298
rect 1542 2292 1548 2293
rect 1563 2295 1572 2296
rect 1326 2291 1332 2292
rect 1563 2291 1564 2295
rect 1571 2291 1572 2295
rect 1638 2293 1639 2297
rect 1643 2293 1644 2297
rect 1734 2297 1740 2298
rect 1638 2292 1644 2293
rect 1658 2295 1665 2296
rect 1563 2290 1572 2291
rect 1658 2291 1659 2295
rect 1664 2291 1665 2295
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1755 2297 1761 2298
rect 1755 2293 1756 2297
rect 1760 2293 1761 2297
rect 1755 2292 1761 2293
rect 1830 2297 1836 2298
rect 1830 2293 1831 2297
rect 1835 2293 1836 2297
rect 1830 2292 1836 2293
rect 1851 2297 1857 2298
rect 1851 2293 1852 2297
rect 1856 2293 1857 2297
rect 1851 2292 1857 2293
rect 1926 2297 1932 2298
rect 1926 2293 1927 2297
rect 1931 2293 1932 2297
rect 1926 2292 1932 2293
rect 1947 2297 1953 2298
rect 1947 2293 1948 2297
rect 1952 2293 1953 2297
rect 1947 2292 1953 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2035 2297 2041 2298
rect 2035 2293 2036 2297
rect 2040 2293 2041 2297
rect 2035 2292 2041 2293
rect 2110 2297 2116 2298
rect 2110 2293 2111 2297
rect 2115 2293 2116 2297
rect 2110 2292 2116 2293
rect 2131 2297 2137 2298
rect 2131 2293 2132 2297
rect 2136 2293 2137 2297
rect 2131 2292 2137 2293
rect 2206 2297 2212 2298
rect 2206 2293 2207 2297
rect 2211 2293 2212 2297
rect 2502 2296 2508 2297
rect 2206 2292 2212 2293
rect 2222 2295 2233 2296
rect 1658 2290 1665 2291
rect 2222 2291 2223 2295
rect 2227 2291 2228 2295
rect 2232 2291 2233 2295
rect 2502 2292 2503 2296
rect 2507 2292 2508 2296
rect 2502 2291 2508 2292
rect 2222 2290 2233 2291
rect 110 2288 116 2289
rect 1286 2288 1292 2289
rect 110 2284 111 2288
rect 115 2284 116 2288
rect 110 2283 116 2284
rect 222 2287 228 2288
rect 222 2283 223 2287
rect 227 2283 228 2287
rect 222 2282 228 2283
rect 243 2287 249 2288
rect 243 2283 244 2287
rect 248 2283 249 2287
rect 243 2282 249 2283
rect 302 2287 308 2288
rect 302 2283 303 2287
rect 307 2283 308 2287
rect 302 2282 308 2283
rect 323 2287 329 2288
rect 323 2283 324 2287
rect 328 2286 329 2287
rect 390 2287 396 2288
rect 328 2284 382 2286
rect 328 2283 329 2284
rect 323 2282 329 2283
rect 245 2274 247 2282
rect 380 2274 382 2284
rect 390 2283 391 2287
rect 395 2283 396 2287
rect 390 2282 396 2283
rect 411 2287 417 2288
rect 411 2283 412 2287
rect 416 2286 417 2287
rect 486 2287 492 2288
rect 416 2284 482 2286
rect 416 2283 417 2284
rect 411 2282 417 2283
rect 480 2274 482 2284
rect 486 2283 487 2287
rect 491 2283 492 2287
rect 486 2282 492 2283
rect 494 2287 500 2288
rect 494 2283 495 2287
rect 499 2286 500 2287
rect 507 2287 513 2288
rect 507 2286 508 2287
rect 499 2284 508 2286
rect 499 2283 500 2284
rect 494 2282 500 2283
rect 507 2283 508 2284
rect 512 2283 513 2287
rect 507 2282 513 2283
rect 574 2287 580 2288
rect 574 2283 575 2287
rect 579 2283 580 2287
rect 574 2282 580 2283
rect 595 2287 601 2288
rect 595 2283 596 2287
rect 600 2286 601 2287
rect 662 2287 668 2288
rect 600 2284 646 2286
rect 600 2283 601 2284
rect 595 2282 601 2283
rect 644 2274 646 2284
rect 662 2283 663 2287
rect 667 2283 668 2287
rect 662 2282 668 2283
rect 683 2287 689 2288
rect 683 2283 684 2287
rect 688 2286 689 2287
rect 750 2287 756 2288
rect 688 2284 742 2286
rect 688 2283 689 2284
rect 683 2282 689 2283
rect 740 2274 742 2284
rect 750 2283 751 2287
rect 755 2283 756 2287
rect 750 2282 756 2283
rect 770 2287 777 2288
rect 770 2283 771 2287
rect 776 2283 777 2287
rect 770 2282 777 2283
rect 830 2287 836 2288
rect 830 2283 831 2287
rect 835 2283 836 2287
rect 830 2282 836 2283
rect 851 2287 857 2288
rect 851 2283 852 2287
rect 856 2286 857 2287
rect 918 2287 924 2288
rect 856 2284 910 2286
rect 856 2283 857 2284
rect 851 2282 857 2283
rect 908 2274 910 2284
rect 918 2283 919 2287
rect 923 2283 924 2287
rect 918 2282 924 2283
rect 939 2287 945 2288
rect 939 2283 940 2287
rect 944 2286 945 2287
rect 974 2287 980 2288
rect 974 2286 975 2287
rect 944 2284 975 2286
rect 944 2283 945 2284
rect 939 2282 945 2283
rect 974 2283 975 2284
rect 979 2283 980 2287
rect 974 2282 980 2283
rect 1006 2287 1012 2288
rect 1006 2283 1007 2287
rect 1011 2283 1012 2287
rect 1006 2282 1012 2283
rect 1027 2287 1033 2288
rect 1027 2283 1028 2287
rect 1032 2286 1033 2287
rect 1094 2287 1100 2288
rect 1032 2284 1086 2286
rect 1032 2283 1033 2284
rect 1027 2282 1033 2283
rect 1084 2274 1086 2284
rect 1094 2283 1095 2287
rect 1099 2283 1100 2287
rect 1094 2282 1100 2283
rect 1102 2287 1108 2288
rect 1102 2283 1103 2287
rect 1107 2286 1108 2287
rect 1115 2287 1121 2288
rect 1115 2286 1116 2287
rect 1107 2284 1116 2286
rect 1107 2283 1108 2284
rect 1102 2282 1108 2283
rect 1115 2283 1116 2284
rect 1120 2283 1121 2287
rect 1286 2284 1287 2288
rect 1291 2284 1292 2288
rect 1286 2283 1292 2284
rect 1115 2282 1121 2283
rect 1326 2279 1332 2280
rect 1326 2275 1327 2279
rect 1331 2275 1332 2279
rect 2502 2279 2508 2280
rect 1326 2274 1332 2275
rect 1350 2276 1356 2277
rect 245 2273 313 2274
rect 245 2272 308 2273
rect 227 2271 233 2272
rect 227 2267 228 2271
rect 232 2270 233 2271
rect 232 2268 278 2270
rect 307 2269 308 2272
rect 312 2269 313 2273
rect 380 2273 401 2274
rect 380 2272 396 2273
rect 307 2268 313 2269
rect 395 2269 396 2272
rect 400 2269 401 2273
rect 480 2273 497 2274
rect 480 2272 492 2273
rect 395 2268 401 2269
rect 491 2269 492 2272
rect 496 2269 497 2273
rect 644 2273 673 2274
rect 644 2272 668 2273
rect 491 2268 497 2269
rect 579 2271 588 2272
rect 232 2267 233 2268
rect 227 2266 233 2267
rect 276 2266 278 2268
rect 510 2267 516 2268
rect 510 2266 511 2267
rect 276 2264 511 2266
rect 510 2263 511 2264
rect 515 2263 516 2267
rect 579 2267 580 2271
rect 587 2267 588 2271
rect 667 2269 668 2272
rect 672 2269 673 2273
rect 740 2273 761 2274
rect 740 2272 756 2273
rect 667 2268 673 2269
rect 755 2269 756 2272
rect 760 2269 761 2273
rect 908 2273 929 2274
rect 908 2272 924 2273
rect 755 2268 761 2269
rect 835 2271 841 2272
rect 579 2266 588 2267
rect 835 2267 836 2271
rect 840 2270 841 2271
rect 840 2268 918 2270
rect 923 2269 924 2272
rect 928 2269 929 2273
rect 1084 2273 1105 2274
rect 1084 2272 1100 2273
rect 923 2268 929 2269
rect 1011 2271 1020 2272
rect 840 2267 841 2268
rect 835 2266 841 2267
rect 510 2262 516 2263
rect 916 2262 918 2268
rect 1011 2267 1012 2271
rect 1019 2267 1020 2271
rect 1099 2269 1100 2272
rect 1104 2269 1105 2273
rect 1350 2272 1351 2276
rect 1355 2272 1356 2276
rect 1350 2271 1356 2272
rect 1438 2276 1444 2277
rect 1438 2272 1439 2276
rect 1443 2272 1444 2276
rect 1438 2271 1444 2272
rect 1526 2276 1532 2277
rect 1526 2272 1527 2276
rect 1531 2272 1532 2276
rect 1526 2271 1532 2272
rect 1622 2276 1628 2277
rect 1622 2272 1623 2276
rect 1627 2272 1628 2276
rect 1622 2271 1628 2272
rect 1718 2276 1724 2277
rect 1718 2272 1719 2276
rect 1723 2272 1724 2276
rect 1718 2271 1724 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1814 2271 1820 2272
rect 1822 2271 1828 2272
rect 1099 2268 1105 2269
rect 1011 2266 1020 2267
rect 1822 2267 1823 2271
rect 1827 2270 1828 2271
rect 1874 2271 1880 2272
rect 1910 2271 1916 2272
rect 1998 2276 2004 2277
rect 1998 2272 1999 2276
rect 2003 2272 2004 2276
rect 1998 2271 2004 2272
rect 2094 2276 2100 2277
rect 2094 2272 2095 2276
rect 2099 2272 2100 2276
rect 2094 2271 2100 2272
rect 2190 2276 2196 2277
rect 2190 2272 2191 2276
rect 2195 2272 2196 2276
rect 2502 2275 2503 2279
rect 2507 2275 2508 2279
rect 2502 2274 2508 2275
rect 2190 2271 2196 2272
rect 1874 2270 1875 2271
rect 1827 2268 1875 2270
rect 1827 2267 1828 2268
rect 1822 2266 1828 2267
rect 1874 2267 1875 2268
rect 1879 2267 1880 2271
rect 1874 2266 1880 2267
rect 1454 2264 1460 2265
rect 1102 2263 1108 2264
rect 1102 2262 1103 2263
rect 916 2260 1103 2262
rect 1102 2259 1103 2260
rect 1107 2259 1108 2263
rect 1102 2258 1108 2259
rect 1326 2261 1332 2262
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1454 2260 1455 2264
rect 1459 2260 1460 2264
rect 1454 2259 1460 2260
rect 1542 2264 1548 2265
rect 1542 2260 1543 2264
rect 1547 2260 1548 2264
rect 1542 2259 1548 2260
rect 1638 2264 1644 2265
rect 1638 2260 1639 2264
rect 1643 2260 1644 2264
rect 1638 2259 1644 2260
rect 1734 2264 1740 2265
rect 1734 2260 1735 2264
rect 1739 2260 1740 2264
rect 1734 2259 1740 2260
rect 1838 2264 1844 2265
rect 1838 2260 1839 2264
rect 1843 2260 1844 2264
rect 1838 2259 1844 2260
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 1934 2259 1940 2260
rect 2030 2264 2036 2265
rect 2030 2260 2031 2264
rect 2035 2260 2036 2264
rect 2030 2259 2036 2260
rect 2118 2264 2124 2265
rect 2118 2260 2119 2264
rect 2123 2260 2124 2264
rect 2118 2259 2124 2260
rect 2214 2264 2220 2265
rect 2214 2260 2215 2264
rect 2219 2260 2220 2264
rect 2214 2259 2220 2260
rect 2310 2264 2316 2265
rect 2310 2260 2311 2264
rect 2315 2260 2316 2264
rect 2310 2259 2316 2260
rect 2502 2261 2508 2262
rect 1326 2256 1332 2257
rect 2502 2257 2503 2261
rect 2507 2257 2508 2261
rect 2502 2256 2508 2257
rect 494 2255 500 2256
rect 494 2254 495 2255
rect 268 2252 495 2254
rect 268 2250 270 2252
rect 494 2251 495 2252
rect 499 2251 500 2255
rect 1130 2255 1136 2256
rect 1130 2254 1131 2255
rect 494 2250 500 2251
rect 924 2252 1131 2254
rect 924 2250 926 2252
rect 1130 2251 1131 2252
rect 1135 2251 1136 2255
rect 1130 2250 1136 2251
rect 267 2249 273 2250
rect 267 2245 268 2249
rect 272 2245 273 2249
rect 923 2249 929 2250
rect 323 2247 329 2248
rect 323 2246 324 2247
rect 267 2244 273 2245
rect 284 2244 324 2246
rect 284 2234 286 2244
rect 323 2243 324 2244
rect 328 2243 329 2247
rect 387 2247 393 2248
rect 387 2246 388 2247
rect 323 2242 329 2243
rect 340 2244 388 2246
rect 340 2234 342 2244
rect 387 2243 388 2244
rect 392 2243 393 2247
rect 451 2247 457 2248
rect 451 2246 452 2247
rect 387 2242 393 2243
rect 404 2244 452 2246
rect 404 2234 406 2244
rect 451 2243 452 2244
rect 456 2243 457 2247
rect 507 2247 513 2248
rect 507 2246 508 2247
rect 451 2242 457 2243
rect 468 2244 508 2246
rect 468 2234 470 2244
rect 507 2243 508 2244
rect 512 2243 513 2247
rect 507 2242 513 2243
rect 563 2247 569 2248
rect 563 2243 564 2247
rect 568 2246 569 2247
rect 619 2247 625 2248
rect 568 2244 614 2246
rect 568 2243 569 2244
rect 563 2242 569 2243
rect 612 2238 614 2244
rect 619 2243 620 2247
rect 624 2246 625 2247
rect 675 2247 681 2248
rect 624 2244 670 2246
rect 624 2243 625 2244
rect 619 2242 625 2243
rect 668 2238 670 2244
rect 675 2243 676 2247
rect 680 2246 681 2247
rect 731 2247 737 2248
rect 680 2244 726 2246
rect 680 2243 681 2244
rect 675 2242 681 2243
rect 724 2238 726 2244
rect 731 2243 732 2247
rect 736 2246 737 2247
rect 795 2247 801 2248
rect 736 2244 786 2246
rect 736 2243 737 2244
rect 731 2242 737 2243
rect 784 2238 786 2244
rect 795 2243 796 2247
rect 800 2246 801 2247
rect 859 2247 865 2248
rect 800 2244 846 2246
rect 800 2243 801 2244
rect 795 2242 801 2243
rect 844 2238 846 2244
rect 859 2243 860 2247
rect 864 2246 865 2247
rect 864 2244 918 2246
rect 923 2245 924 2249
rect 928 2245 929 2249
rect 923 2244 929 2245
rect 974 2247 980 2248
rect 864 2243 865 2244
rect 859 2242 865 2243
rect 916 2238 918 2244
rect 974 2243 975 2247
rect 979 2246 980 2247
rect 987 2247 993 2248
rect 987 2246 988 2247
rect 979 2244 988 2246
rect 979 2243 980 2244
rect 974 2242 980 2243
rect 987 2243 988 2244
rect 992 2243 993 2247
rect 1051 2247 1057 2248
rect 1051 2246 1052 2247
rect 987 2242 993 2243
rect 1004 2244 1052 2246
rect 612 2236 638 2238
rect 668 2236 695 2238
rect 724 2236 750 2238
rect 784 2236 814 2238
rect 844 2236 878 2238
rect 916 2236 942 2238
rect 636 2234 638 2236
rect 693 2234 695 2236
rect 748 2234 750 2236
rect 812 2234 814 2236
rect 876 2234 878 2236
rect 940 2234 942 2236
rect 1004 2234 1006 2244
rect 1051 2243 1052 2244
rect 1056 2243 1057 2247
rect 1115 2247 1121 2248
rect 1115 2246 1116 2247
rect 1051 2242 1057 2243
rect 1068 2244 1116 2246
rect 1068 2234 1070 2244
rect 1115 2243 1116 2244
rect 1120 2243 1121 2247
rect 1115 2242 1121 2243
rect 1326 2244 1332 2245
rect 2502 2244 2508 2245
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1326 2239 1332 2240
rect 1470 2243 1476 2244
rect 1470 2239 1471 2243
rect 1475 2239 1476 2243
rect 1470 2238 1476 2239
rect 1491 2243 1497 2244
rect 1491 2239 1492 2243
rect 1496 2242 1497 2243
rect 1558 2243 1564 2244
rect 1496 2240 1550 2242
rect 1496 2239 1497 2240
rect 1491 2238 1497 2239
rect 262 2233 268 2234
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 262 2229 263 2233
rect 267 2229 268 2233
rect 262 2228 268 2229
rect 283 2233 289 2234
rect 283 2229 284 2233
rect 288 2229 289 2233
rect 283 2228 289 2229
rect 318 2233 324 2234
rect 318 2229 319 2233
rect 323 2229 324 2233
rect 318 2228 324 2229
rect 339 2233 345 2234
rect 339 2229 340 2233
rect 344 2229 345 2233
rect 339 2228 345 2229
rect 382 2233 388 2234
rect 382 2229 383 2233
rect 387 2229 388 2233
rect 382 2228 388 2229
rect 403 2233 409 2234
rect 403 2229 404 2233
rect 408 2229 409 2233
rect 403 2228 409 2229
rect 446 2233 452 2234
rect 446 2229 447 2233
rect 451 2229 452 2233
rect 446 2228 452 2229
rect 467 2233 473 2234
rect 467 2229 468 2233
rect 472 2229 473 2233
rect 467 2228 473 2229
rect 502 2233 508 2234
rect 502 2229 503 2233
rect 507 2229 508 2233
rect 558 2233 564 2234
rect 502 2228 508 2229
rect 510 2231 516 2232
rect 110 2227 116 2228
rect 510 2227 511 2231
rect 515 2230 516 2231
rect 523 2231 529 2232
rect 523 2230 524 2231
rect 515 2228 524 2230
rect 515 2227 516 2228
rect 510 2226 516 2227
rect 523 2227 524 2228
rect 528 2227 529 2231
rect 558 2229 559 2233
rect 563 2229 564 2233
rect 614 2233 620 2234
rect 558 2228 564 2229
rect 579 2231 588 2232
rect 523 2226 529 2227
rect 579 2227 580 2231
rect 587 2227 588 2231
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 635 2233 641 2234
rect 635 2229 636 2233
rect 640 2229 641 2233
rect 635 2228 641 2229
rect 670 2233 676 2234
rect 670 2229 671 2233
rect 675 2229 676 2233
rect 670 2228 676 2229
rect 691 2233 697 2234
rect 691 2229 692 2233
rect 696 2229 697 2233
rect 691 2228 697 2229
rect 726 2233 732 2234
rect 726 2229 727 2233
rect 731 2229 732 2233
rect 726 2228 732 2229
rect 747 2233 753 2234
rect 747 2229 748 2233
rect 752 2229 753 2233
rect 747 2228 753 2229
rect 790 2233 796 2234
rect 790 2229 791 2233
rect 795 2229 796 2233
rect 790 2228 796 2229
rect 811 2233 817 2234
rect 811 2229 812 2233
rect 816 2229 817 2233
rect 811 2228 817 2229
rect 854 2233 860 2234
rect 854 2229 855 2233
rect 859 2229 860 2233
rect 854 2228 860 2229
rect 875 2233 881 2234
rect 875 2229 876 2233
rect 880 2229 881 2233
rect 875 2228 881 2229
rect 918 2233 924 2234
rect 918 2229 919 2233
rect 923 2229 924 2233
rect 918 2228 924 2229
rect 939 2233 945 2234
rect 939 2229 940 2233
rect 944 2229 945 2233
rect 939 2228 945 2229
rect 982 2233 988 2234
rect 982 2229 983 2233
rect 987 2229 988 2233
rect 982 2228 988 2229
rect 1003 2233 1009 2234
rect 1003 2229 1004 2233
rect 1008 2229 1009 2233
rect 1003 2228 1009 2229
rect 1046 2233 1052 2234
rect 1046 2229 1047 2233
rect 1051 2229 1052 2233
rect 1046 2228 1052 2229
rect 1067 2233 1073 2234
rect 1067 2229 1068 2233
rect 1072 2229 1073 2233
rect 1067 2228 1073 2229
rect 1110 2233 1116 2234
rect 1110 2229 1111 2233
rect 1115 2229 1116 2233
rect 1286 2232 1292 2233
rect 1110 2228 1116 2229
rect 1130 2231 1137 2232
rect 579 2226 588 2227
rect 1130 2227 1131 2231
rect 1136 2227 1137 2231
rect 1286 2228 1287 2232
rect 1291 2228 1292 2232
rect 1548 2230 1550 2240
rect 1558 2239 1559 2243
rect 1563 2239 1564 2243
rect 1558 2238 1564 2239
rect 1579 2243 1585 2244
rect 1579 2239 1580 2243
rect 1584 2242 1585 2243
rect 1654 2243 1660 2244
rect 1584 2240 1650 2242
rect 1584 2239 1585 2240
rect 1579 2238 1585 2239
rect 1648 2230 1650 2240
rect 1654 2239 1655 2243
rect 1659 2239 1660 2243
rect 1654 2238 1660 2239
rect 1675 2243 1681 2244
rect 1675 2239 1676 2243
rect 1680 2242 1681 2243
rect 1750 2243 1756 2244
rect 1680 2240 1746 2242
rect 1680 2239 1681 2240
rect 1675 2238 1681 2239
rect 1744 2230 1746 2240
rect 1750 2239 1751 2243
rect 1755 2239 1756 2243
rect 1750 2238 1756 2239
rect 1771 2243 1777 2244
rect 1771 2239 1772 2243
rect 1776 2242 1777 2243
rect 1854 2243 1860 2244
rect 1776 2240 1850 2242
rect 1776 2239 1777 2240
rect 1771 2238 1777 2239
rect 1848 2230 1850 2240
rect 1854 2239 1855 2243
rect 1859 2239 1860 2243
rect 1854 2238 1860 2239
rect 1874 2243 1881 2244
rect 1874 2239 1875 2243
rect 1880 2239 1881 2243
rect 1874 2238 1881 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 1971 2243 1977 2244
rect 1971 2239 1972 2243
rect 1976 2242 1977 2243
rect 2046 2243 2052 2244
rect 1976 2240 2001 2242
rect 1976 2239 1977 2240
rect 1971 2238 1977 2239
rect 1999 2230 2001 2240
rect 2046 2239 2047 2243
rect 2051 2239 2052 2243
rect 2046 2238 2052 2239
rect 2067 2243 2073 2244
rect 2067 2239 2068 2243
rect 2072 2242 2073 2243
rect 2134 2243 2140 2244
rect 2072 2240 2126 2242
rect 2072 2239 2073 2240
rect 2067 2238 2073 2239
rect 2124 2230 2126 2240
rect 2134 2239 2135 2243
rect 2139 2239 2140 2243
rect 2134 2238 2140 2239
rect 2155 2243 2161 2244
rect 2155 2239 2156 2243
rect 2160 2242 2161 2243
rect 2230 2243 2236 2244
rect 2160 2240 2226 2242
rect 2160 2239 2161 2240
rect 2155 2238 2161 2239
rect 2224 2230 2226 2240
rect 2230 2239 2231 2243
rect 2235 2239 2236 2243
rect 2230 2238 2236 2239
rect 2251 2243 2257 2244
rect 2251 2239 2252 2243
rect 2256 2242 2257 2243
rect 2326 2243 2332 2244
rect 2256 2240 2318 2242
rect 2256 2239 2257 2240
rect 2251 2238 2257 2239
rect 2316 2230 2318 2240
rect 2326 2239 2327 2243
rect 2331 2239 2332 2243
rect 2326 2238 2332 2239
rect 2334 2243 2340 2244
rect 2334 2239 2335 2243
rect 2339 2242 2340 2243
rect 2347 2243 2353 2244
rect 2347 2242 2348 2243
rect 2339 2240 2348 2242
rect 2339 2239 2340 2240
rect 2334 2238 2340 2239
rect 2347 2239 2348 2240
rect 2352 2239 2353 2243
rect 2502 2240 2503 2244
rect 2507 2240 2508 2244
rect 2502 2239 2508 2240
rect 2347 2238 2353 2239
rect 1548 2229 1569 2230
rect 1548 2228 1564 2229
rect 1286 2227 1292 2228
rect 1475 2227 1481 2228
rect 1130 2226 1137 2227
rect 1475 2223 1476 2227
rect 1480 2226 1481 2227
rect 1480 2224 1558 2226
rect 1563 2225 1564 2228
rect 1568 2225 1569 2229
rect 1648 2229 1665 2230
rect 1648 2228 1660 2229
rect 1563 2224 1569 2225
rect 1659 2225 1660 2228
rect 1664 2225 1665 2229
rect 1744 2229 1761 2230
rect 1744 2228 1756 2229
rect 1659 2224 1665 2225
rect 1755 2225 1756 2228
rect 1760 2225 1761 2229
rect 1848 2229 1865 2230
rect 1848 2228 1860 2229
rect 1755 2224 1761 2225
rect 1859 2225 1860 2228
rect 1864 2225 1865 2229
rect 1999 2229 2057 2230
rect 1999 2228 2052 2229
rect 1859 2224 1865 2225
rect 1955 2227 1961 2228
rect 1480 2223 1481 2224
rect 1475 2222 1481 2223
rect 1556 2222 1558 2224
rect 1586 2223 1592 2224
rect 1586 2222 1587 2223
rect 1556 2220 1587 2222
rect 1586 2219 1587 2220
rect 1591 2219 1592 2223
rect 1955 2223 1956 2227
rect 1960 2226 1961 2227
rect 1960 2224 2001 2226
rect 2051 2225 2052 2228
rect 2056 2225 2057 2229
rect 2124 2229 2145 2230
rect 2124 2228 2140 2229
rect 2051 2224 2057 2225
rect 2139 2225 2140 2228
rect 2144 2225 2145 2229
rect 2224 2229 2241 2230
rect 2224 2228 2236 2229
rect 2139 2224 2145 2225
rect 2235 2225 2236 2228
rect 2240 2225 2241 2229
rect 2316 2229 2337 2230
rect 2316 2228 2332 2229
rect 2235 2224 2241 2225
rect 2331 2225 2332 2228
rect 2336 2225 2337 2229
rect 2331 2224 2337 2225
rect 1960 2223 1961 2224
rect 1955 2222 1961 2223
rect 1999 2222 2001 2224
rect 2222 2223 2228 2224
rect 2222 2222 2223 2223
rect 1999 2220 2223 2222
rect 1586 2218 1592 2219
rect 2222 2219 2223 2220
rect 2227 2219 2228 2223
rect 2222 2218 2228 2219
rect 110 2215 116 2216
rect 110 2211 111 2215
rect 115 2211 116 2215
rect 1286 2215 1292 2216
rect 110 2210 116 2211
rect 246 2212 252 2213
rect 246 2208 247 2212
rect 251 2208 252 2212
rect 246 2207 252 2208
rect 302 2212 308 2213
rect 302 2208 303 2212
rect 307 2208 308 2212
rect 302 2207 308 2208
rect 366 2212 372 2213
rect 366 2208 367 2212
rect 371 2208 372 2212
rect 366 2207 372 2208
rect 430 2212 436 2213
rect 430 2208 431 2212
rect 435 2208 436 2212
rect 430 2207 436 2208
rect 486 2212 492 2213
rect 486 2208 487 2212
rect 491 2208 492 2212
rect 486 2207 492 2208
rect 542 2212 548 2213
rect 542 2208 543 2212
rect 547 2208 548 2212
rect 542 2207 548 2208
rect 598 2212 604 2213
rect 598 2208 599 2212
rect 603 2208 604 2212
rect 598 2207 604 2208
rect 654 2212 660 2213
rect 654 2208 655 2212
rect 659 2208 660 2212
rect 654 2207 660 2208
rect 710 2212 716 2213
rect 710 2208 711 2212
rect 715 2208 716 2212
rect 710 2207 716 2208
rect 774 2212 780 2213
rect 774 2208 775 2212
rect 779 2208 780 2212
rect 774 2207 780 2208
rect 838 2212 844 2213
rect 838 2208 839 2212
rect 843 2208 844 2212
rect 838 2207 844 2208
rect 902 2212 908 2213
rect 902 2208 903 2212
rect 907 2208 908 2212
rect 902 2207 908 2208
rect 966 2212 972 2213
rect 966 2208 967 2212
rect 971 2208 972 2212
rect 966 2207 972 2208
rect 1030 2212 1036 2213
rect 1030 2208 1031 2212
rect 1035 2208 1036 2212
rect 1030 2207 1036 2208
rect 1094 2212 1100 2213
rect 1094 2208 1095 2212
rect 1099 2208 1100 2212
rect 1286 2211 1287 2215
rect 1291 2211 1292 2215
rect 1286 2210 1292 2211
rect 1890 2211 1896 2212
rect 1890 2210 1891 2211
rect 1094 2207 1100 2208
rect 1748 2208 1891 2210
rect 1748 2206 1750 2208
rect 1890 2207 1891 2208
rect 1895 2207 1896 2211
rect 2334 2211 2340 2212
rect 2334 2210 2335 2211
rect 1890 2206 1896 2207
rect 1932 2208 2335 2210
rect 1932 2206 1934 2208
rect 2334 2207 2335 2208
rect 2339 2207 2340 2211
rect 2334 2206 2340 2207
rect 1747 2205 1753 2206
rect 358 2203 364 2204
rect 358 2199 359 2203
rect 363 2202 364 2203
rect 510 2203 516 2204
rect 510 2202 511 2203
rect 363 2200 511 2202
rect 363 2199 364 2200
rect 358 2198 364 2199
rect 510 2199 511 2200
rect 515 2199 516 2203
rect 510 2198 516 2199
rect 1571 2203 1577 2204
rect 1571 2199 1572 2203
rect 1576 2202 1577 2203
rect 1627 2203 1633 2204
rect 1576 2200 1622 2202
rect 1576 2199 1577 2200
rect 1571 2198 1577 2199
rect 334 2196 340 2197
rect 110 2193 116 2194
rect 110 2189 111 2193
rect 115 2189 116 2193
rect 334 2192 335 2196
rect 339 2192 340 2196
rect 334 2191 340 2192
rect 390 2196 396 2197
rect 390 2192 391 2196
rect 395 2192 396 2196
rect 390 2191 396 2192
rect 446 2196 452 2197
rect 446 2192 447 2196
rect 451 2192 452 2196
rect 446 2191 452 2192
rect 502 2196 508 2197
rect 502 2192 503 2196
rect 507 2192 508 2196
rect 502 2191 508 2192
rect 558 2196 564 2197
rect 558 2192 559 2196
rect 563 2192 564 2196
rect 1620 2194 1622 2200
rect 1627 2199 1628 2203
rect 1632 2202 1633 2203
rect 1683 2203 1689 2204
rect 1632 2200 1678 2202
rect 1632 2199 1633 2200
rect 1627 2198 1633 2199
rect 1676 2194 1678 2200
rect 1683 2199 1684 2203
rect 1688 2202 1689 2203
rect 1688 2200 1742 2202
rect 1747 2201 1748 2205
rect 1752 2201 1753 2205
rect 1931 2205 1937 2206
rect 1747 2200 1753 2201
rect 1811 2203 1817 2204
rect 1688 2199 1689 2200
rect 1683 2198 1689 2199
rect 1740 2194 1742 2200
rect 1811 2199 1812 2203
rect 1816 2202 1817 2203
rect 1826 2203 1832 2204
rect 1826 2202 1827 2203
rect 1816 2200 1827 2202
rect 1816 2199 1817 2200
rect 1811 2198 1817 2199
rect 1826 2199 1827 2200
rect 1831 2199 1832 2203
rect 1875 2203 1881 2204
rect 1875 2202 1876 2203
rect 1826 2198 1832 2199
rect 1852 2200 1876 2202
rect 1852 2194 1854 2200
rect 1875 2199 1876 2200
rect 1880 2199 1881 2203
rect 1931 2201 1932 2205
rect 1936 2201 1937 2205
rect 1987 2203 1993 2204
rect 1987 2202 1988 2203
rect 1931 2200 1937 2201
rect 1964 2200 1988 2202
rect 1875 2198 1881 2199
rect 1964 2194 1966 2200
rect 1987 2199 1988 2200
rect 1992 2199 1993 2203
rect 2043 2203 2049 2204
rect 2043 2202 2044 2203
rect 1987 2198 1993 2199
rect 2004 2200 2044 2202
rect 558 2191 564 2192
rect 1286 2193 1292 2194
rect 110 2188 116 2189
rect 1286 2189 1287 2193
rect 1291 2189 1292 2193
rect 1620 2192 1646 2194
rect 1676 2192 1702 2194
rect 1740 2192 1766 2194
rect 1644 2190 1646 2192
rect 1700 2190 1702 2192
rect 1764 2190 1766 2192
rect 1828 2192 1854 2194
rect 1948 2192 1966 2194
rect 1828 2190 1830 2192
rect 1948 2190 1950 2192
rect 2004 2190 2006 2200
rect 2043 2199 2044 2200
rect 2048 2199 2049 2203
rect 2099 2203 2105 2204
rect 2099 2202 2100 2203
rect 2043 2198 2049 2199
rect 2072 2200 2100 2202
rect 2072 2194 2074 2200
rect 2099 2199 2100 2200
rect 2104 2199 2105 2203
rect 2163 2203 2169 2204
rect 2163 2202 2164 2203
rect 2099 2198 2105 2199
rect 2116 2200 2164 2202
rect 2060 2192 2074 2194
rect 2060 2190 2062 2192
rect 2116 2190 2118 2200
rect 2163 2199 2164 2200
rect 2168 2199 2169 2203
rect 2227 2203 2233 2204
rect 2227 2202 2228 2203
rect 2163 2198 2169 2199
rect 2180 2200 2228 2202
rect 2180 2190 2182 2200
rect 2227 2199 2228 2200
rect 2232 2199 2233 2203
rect 2291 2203 2297 2204
rect 2291 2202 2292 2203
rect 2227 2198 2233 2199
rect 2248 2200 2292 2202
rect 2248 2194 2250 2200
rect 2291 2199 2292 2200
rect 2296 2199 2297 2203
rect 2347 2203 2353 2204
rect 2347 2202 2348 2203
rect 2291 2198 2297 2199
rect 2312 2200 2348 2202
rect 2312 2194 2314 2200
rect 2347 2199 2348 2200
rect 2352 2199 2353 2203
rect 2403 2203 2409 2204
rect 2403 2202 2404 2203
rect 2347 2198 2353 2199
rect 2368 2200 2404 2202
rect 2368 2194 2370 2200
rect 2403 2199 2404 2200
rect 2408 2199 2409 2203
rect 2459 2203 2465 2204
rect 2459 2202 2460 2203
rect 2403 2198 2409 2199
rect 2424 2200 2460 2202
rect 2424 2194 2426 2200
rect 2459 2199 2460 2200
rect 2464 2199 2465 2203
rect 2459 2198 2465 2199
rect 2244 2192 2250 2194
rect 2308 2192 2314 2194
rect 2364 2192 2370 2194
rect 2420 2192 2426 2194
rect 2244 2190 2246 2192
rect 2308 2190 2310 2192
rect 2364 2190 2366 2192
rect 2420 2190 2422 2192
rect 1566 2189 1572 2190
rect 1286 2188 1292 2189
rect 1326 2188 1332 2189
rect 1326 2184 1327 2188
rect 1331 2184 1332 2188
rect 1566 2185 1567 2189
rect 1571 2185 1572 2189
rect 1622 2189 1628 2190
rect 1566 2184 1572 2185
rect 1586 2187 1593 2188
rect 1326 2183 1332 2184
rect 1586 2183 1587 2187
rect 1592 2183 1593 2187
rect 1622 2185 1623 2189
rect 1627 2185 1628 2189
rect 1622 2184 1628 2185
rect 1643 2189 1649 2190
rect 1643 2185 1644 2189
rect 1648 2185 1649 2189
rect 1643 2184 1649 2185
rect 1678 2189 1684 2190
rect 1678 2185 1679 2189
rect 1683 2185 1684 2189
rect 1678 2184 1684 2185
rect 1699 2189 1705 2190
rect 1699 2185 1700 2189
rect 1704 2185 1705 2189
rect 1699 2184 1705 2185
rect 1742 2189 1748 2190
rect 1742 2185 1743 2189
rect 1747 2185 1748 2189
rect 1742 2184 1748 2185
rect 1763 2189 1769 2190
rect 1763 2185 1764 2189
rect 1768 2185 1769 2189
rect 1763 2184 1769 2185
rect 1806 2189 1812 2190
rect 1806 2185 1807 2189
rect 1811 2185 1812 2189
rect 1806 2184 1812 2185
rect 1827 2189 1833 2190
rect 1827 2185 1828 2189
rect 1832 2185 1833 2189
rect 1827 2184 1833 2185
rect 1870 2189 1876 2190
rect 1870 2185 1871 2189
rect 1875 2185 1876 2189
rect 1926 2189 1932 2190
rect 1870 2184 1876 2185
rect 1890 2187 1897 2188
rect 1586 2182 1593 2183
rect 1890 2183 1891 2187
rect 1896 2183 1897 2187
rect 1926 2185 1927 2189
rect 1931 2185 1932 2189
rect 1926 2184 1932 2185
rect 1947 2189 1953 2190
rect 1947 2185 1948 2189
rect 1952 2185 1953 2189
rect 1947 2184 1953 2185
rect 1982 2189 1988 2190
rect 1982 2185 1983 2189
rect 1987 2185 1988 2189
rect 1982 2184 1988 2185
rect 2003 2189 2009 2190
rect 2003 2185 2004 2189
rect 2008 2185 2009 2189
rect 2003 2184 2009 2185
rect 2038 2189 2044 2190
rect 2038 2185 2039 2189
rect 2043 2185 2044 2189
rect 2038 2184 2044 2185
rect 2059 2189 2065 2190
rect 2059 2185 2060 2189
rect 2064 2185 2065 2189
rect 2059 2184 2065 2185
rect 2094 2189 2100 2190
rect 2094 2185 2095 2189
rect 2099 2185 2100 2189
rect 2094 2184 2100 2185
rect 2115 2189 2121 2190
rect 2115 2185 2116 2189
rect 2120 2185 2121 2189
rect 2115 2184 2121 2185
rect 2158 2189 2164 2190
rect 2158 2185 2159 2189
rect 2163 2185 2164 2189
rect 2158 2184 2164 2185
rect 2179 2189 2185 2190
rect 2179 2185 2180 2189
rect 2184 2185 2185 2189
rect 2179 2184 2185 2185
rect 2222 2189 2228 2190
rect 2222 2185 2223 2189
rect 2227 2185 2228 2189
rect 2222 2184 2228 2185
rect 2243 2189 2249 2190
rect 2243 2185 2244 2189
rect 2248 2185 2249 2189
rect 2243 2184 2249 2185
rect 2286 2189 2292 2190
rect 2286 2185 2287 2189
rect 2291 2185 2292 2189
rect 2286 2184 2292 2185
rect 2307 2189 2313 2190
rect 2307 2185 2308 2189
rect 2312 2185 2313 2189
rect 2307 2184 2313 2185
rect 2342 2189 2348 2190
rect 2342 2185 2343 2189
rect 2347 2185 2348 2189
rect 2342 2184 2348 2185
rect 2363 2189 2369 2190
rect 2363 2185 2364 2189
rect 2368 2185 2369 2189
rect 2363 2184 2369 2185
rect 2398 2189 2404 2190
rect 2398 2185 2399 2189
rect 2403 2185 2404 2189
rect 2398 2184 2404 2185
rect 2419 2189 2425 2190
rect 2419 2185 2420 2189
rect 2424 2185 2425 2189
rect 2419 2184 2425 2185
rect 2454 2189 2460 2190
rect 2454 2185 2455 2189
rect 2459 2185 2460 2189
rect 2502 2188 2508 2189
rect 2454 2184 2460 2185
rect 2470 2187 2481 2188
rect 1890 2182 1897 2183
rect 2470 2183 2471 2187
rect 2475 2183 2476 2187
rect 2480 2183 2481 2187
rect 2502 2184 2503 2188
rect 2507 2184 2508 2188
rect 2502 2183 2508 2184
rect 2470 2182 2481 2183
rect 110 2176 116 2177
rect 1286 2176 1292 2177
rect 110 2172 111 2176
rect 115 2172 116 2176
rect 110 2171 116 2172
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 350 2170 356 2171
rect 371 2175 377 2176
rect 371 2171 372 2175
rect 376 2174 377 2175
rect 406 2175 412 2176
rect 376 2172 402 2174
rect 376 2171 377 2172
rect 371 2170 377 2171
rect 400 2162 402 2172
rect 406 2171 407 2175
rect 411 2171 412 2175
rect 406 2170 412 2171
rect 427 2175 433 2176
rect 427 2171 428 2175
rect 432 2174 433 2175
rect 462 2175 468 2176
rect 432 2172 458 2174
rect 432 2171 433 2172
rect 427 2170 433 2171
rect 456 2162 458 2172
rect 462 2171 463 2175
rect 467 2171 468 2175
rect 462 2170 468 2171
rect 483 2175 489 2176
rect 483 2171 484 2175
rect 488 2174 489 2175
rect 518 2175 524 2176
rect 488 2172 514 2174
rect 488 2171 489 2172
rect 483 2170 489 2171
rect 512 2162 514 2172
rect 518 2171 519 2175
rect 523 2171 524 2175
rect 518 2170 524 2171
rect 539 2175 545 2176
rect 539 2171 540 2175
rect 544 2174 545 2175
rect 574 2175 580 2176
rect 544 2172 570 2174
rect 544 2171 545 2172
rect 539 2170 545 2171
rect 568 2162 570 2172
rect 574 2171 575 2175
rect 579 2171 580 2175
rect 574 2170 580 2171
rect 582 2175 588 2176
rect 582 2171 583 2175
rect 587 2174 588 2175
rect 595 2175 601 2176
rect 595 2174 596 2175
rect 587 2172 596 2174
rect 587 2171 588 2172
rect 582 2170 588 2171
rect 595 2171 596 2172
rect 600 2171 601 2175
rect 1286 2172 1287 2176
rect 1291 2172 1292 2176
rect 1286 2171 1292 2172
rect 1326 2171 1332 2172
rect 595 2170 601 2171
rect 1326 2167 1327 2171
rect 1331 2167 1332 2171
rect 2502 2171 2508 2172
rect 1326 2166 1332 2167
rect 1550 2168 1556 2169
rect 1550 2164 1551 2168
rect 1555 2164 1556 2168
rect 1550 2163 1556 2164
rect 1606 2168 1612 2169
rect 1606 2164 1607 2168
rect 1611 2164 1612 2168
rect 1606 2163 1612 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1726 2168 1732 2169
rect 1726 2164 1727 2168
rect 1731 2164 1732 2168
rect 1726 2163 1732 2164
rect 1790 2168 1796 2169
rect 1790 2164 1791 2168
rect 1795 2164 1796 2168
rect 1790 2163 1796 2164
rect 1854 2168 1860 2169
rect 1854 2164 1855 2168
rect 1859 2164 1860 2168
rect 1854 2163 1860 2164
rect 1910 2168 1916 2169
rect 1910 2164 1911 2168
rect 1915 2164 1916 2168
rect 1910 2163 1916 2164
rect 1966 2168 1972 2169
rect 1966 2164 1967 2168
rect 1971 2164 1972 2168
rect 1966 2163 1972 2164
rect 2022 2168 2028 2169
rect 2022 2164 2023 2168
rect 2027 2164 2028 2168
rect 2022 2163 2028 2164
rect 2078 2168 2084 2169
rect 2078 2164 2079 2168
rect 2083 2164 2084 2168
rect 2078 2163 2084 2164
rect 2142 2168 2148 2169
rect 2142 2164 2143 2168
rect 2147 2164 2148 2168
rect 2142 2163 2148 2164
rect 2206 2168 2212 2169
rect 2206 2164 2207 2168
rect 2211 2164 2212 2168
rect 2206 2163 2212 2164
rect 2270 2168 2276 2169
rect 2270 2164 2271 2168
rect 2275 2164 2276 2168
rect 2270 2163 2276 2164
rect 2326 2168 2332 2169
rect 2326 2164 2327 2168
rect 2331 2164 2332 2168
rect 2326 2163 2332 2164
rect 2382 2168 2388 2169
rect 2382 2164 2383 2168
rect 2387 2164 2388 2168
rect 2382 2163 2388 2164
rect 2438 2168 2444 2169
rect 2438 2164 2439 2168
rect 2443 2164 2444 2168
rect 2502 2167 2503 2171
rect 2507 2167 2508 2171
rect 2502 2166 2508 2167
rect 2438 2163 2444 2164
rect 400 2161 417 2162
rect 400 2160 412 2161
rect 355 2159 364 2160
rect 355 2155 356 2159
rect 363 2155 364 2159
rect 411 2157 412 2160
rect 416 2157 417 2161
rect 456 2161 473 2162
rect 456 2160 468 2161
rect 411 2156 417 2157
rect 467 2157 468 2160
rect 472 2157 473 2161
rect 512 2161 529 2162
rect 512 2160 524 2161
rect 467 2156 473 2157
rect 523 2157 524 2160
rect 528 2157 529 2161
rect 568 2161 585 2162
rect 568 2160 580 2161
rect 523 2156 529 2157
rect 579 2157 580 2160
rect 584 2157 585 2161
rect 579 2156 585 2157
rect 355 2154 364 2155
rect 582 2147 588 2148
rect 582 2146 583 2147
rect 420 2144 583 2146
rect 420 2142 422 2144
rect 582 2143 583 2144
rect 587 2143 588 2147
rect 1126 2147 1132 2148
rect 1126 2146 1127 2147
rect 582 2142 588 2143
rect 932 2144 1127 2146
rect 932 2142 934 2144
rect 1126 2143 1127 2144
rect 1131 2143 1132 2147
rect 1126 2142 1132 2143
rect 1662 2144 1668 2145
rect 419 2141 425 2142
rect 419 2137 420 2141
rect 424 2137 425 2141
rect 931 2141 937 2142
rect 515 2139 521 2140
rect 515 2138 516 2139
rect 419 2136 425 2137
rect 436 2136 516 2138
rect 436 2126 438 2136
rect 515 2135 516 2136
rect 520 2135 521 2139
rect 611 2139 617 2140
rect 611 2138 612 2139
rect 515 2134 521 2135
rect 533 2136 612 2138
rect 533 2126 535 2136
rect 611 2135 612 2136
rect 616 2135 617 2139
rect 715 2139 721 2140
rect 715 2138 716 2139
rect 611 2134 617 2135
rect 628 2136 716 2138
rect 628 2126 630 2136
rect 715 2135 716 2136
rect 720 2135 721 2139
rect 819 2139 825 2140
rect 819 2138 820 2139
rect 715 2134 721 2135
rect 732 2136 820 2138
rect 732 2126 734 2136
rect 819 2135 820 2136
rect 824 2135 825 2139
rect 931 2137 932 2141
rect 936 2137 937 2141
rect 1326 2141 1332 2142
rect 931 2136 937 2137
rect 1043 2139 1049 2140
rect 819 2134 825 2135
rect 1043 2135 1044 2139
rect 1048 2135 1049 2139
rect 1155 2139 1161 2140
rect 1155 2138 1156 2139
rect 1043 2134 1049 2135
rect 1072 2136 1156 2138
rect 1045 2130 1047 2134
rect 948 2128 1047 2130
rect 948 2126 950 2128
rect 1072 2126 1074 2136
rect 1155 2135 1156 2136
rect 1160 2135 1161 2139
rect 1243 2139 1249 2140
rect 1243 2138 1244 2139
rect 1155 2134 1161 2135
rect 1212 2136 1244 2138
rect 1212 2126 1214 2136
rect 1243 2135 1244 2136
rect 1248 2135 1249 2139
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1718 2144 1724 2145
rect 1718 2140 1719 2144
rect 1723 2140 1724 2144
rect 1718 2139 1724 2140
rect 1790 2144 1796 2145
rect 1790 2140 1791 2144
rect 1795 2140 1796 2144
rect 1790 2139 1796 2140
rect 1870 2144 1876 2145
rect 1870 2140 1871 2144
rect 1875 2140 1876 2144
rect 1870 2139 1876 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2078 2144 2084 2145
rect 2078 2140 2079 2144
rect 2083 2140 2084 2144
rect 2078 2139 2084 2140
rect 2198 2144 2204 2145
rect 2198 2140 2199 2144
rect 2203 2140 2204 2144
rect 2198 2139 2204 2140
rect 2326 2144 2332 2145
rect 2326 2140 2327 2144
rect 2331 2140 2332 2144
rect 2326 2139 2332 2140
rect 2438 2144 2444 2145
rect 2438 2140 2439 2144
rect 2443 2140 2444 2144
rect 2438 2139 2444 2140
rect 2502 2141 2508 2142
rect 1326 2136 1332 2137
rect 2502 2137 2503 2141
rect 2507 2137 2508 2141
rect 2502 2136 2508 2137
rect 1243 2134 1249 2135
rect 414 2125 420 2126
rect 110 2124 116 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 414 2121 415 2125
rect 419 2121 420 2125
rect 414 2120 420 2121
rect 435 2125 441 2126
rect 435 2121 436 2125
rect 440 2121 441 2125
rect 435 2120 441 2121
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 531 2125 537 2126
rect 531 2121 532 2125
rect 536 2121 537 2125
rect 531 2120 537 2121
rect 606 2125 612 2126
rect 606 2121 607 2125
rect 611 2121 612 2125
rect 606 2120 612 2121
rect 627 2125 633 2126
rect 627 2121 628 2125
rect 632 2121 633 2125
rect 627 2120 633 2121
rect 710 2125 716 2126
rect 710 2121 711 2125
rect 715 2121 716 2125
rect 710 2120 716 2121
rect 731 2125 737 2126
rect 731 2121 732 2125
rect 736 2121 737 2125
rect 731 2120 737 2121
rect 814 2125 820 2126
rect 814 2121 815 2125
rect 819 2121 820 2125
rect 926 2125 932 2126
rect 814 2120 820 2121
rect 822 2123 828 2124
rect 110 2119 116 2120
rect 822 2119 823 2123
rect 827 2122 828 2123
rect 835 2123 841 2124
rect 835 2122 836 2123
rect 827 2120 836 2122
rect 827 2119 828 2120
rect 822 2118 828 2119
rect 835 2119 836 2120
rect 840 2119 841 2123
rect 926 2121 927 2125
rect 931 2121 932 2125
rect 926 2120 932 2121
rect 947 2125 953 2126
rect 947 2121 948 2125
rect 952 2121 953 2125
rect 947 2120 953 2121
rect 1038 2125 1044 2126
rect 1038 2121 1039 2125
rect 1043 2121 1044 2125
rect 1038 2120 1044 2121
rect 1059 2125 1074 2126
rect 1059 2121 1060 2125
rect 1064 2124 1074 2125
rect 1150 2125 1156 2126
rect 1064 2121 1065 2124
rect 1059 2120 1065 2121
rect 1150 2121 1151 2125
rect 1155 2121 1156 2125
rect 1150 2120 1156 2121
rect 1171 2125 1214 2126
rect 1171 2121 1172 2125
rect 1176 2124 1214 2125
rect 1238 2125 1244 2126
rect 1176 2121 1177 2124
rect 1171 2120 1177 2121
rect 1238 2121 1239 2125
rect 1243 2121 1244 2125
rect 1286 2124 1292 2125
rect 1238 2120 1244 2121
rect 1254 2123 1265 2124
rect 835 2118 841 2119
rect 1254 2119 1255 2123
rect 1259 2119 1260 2123
rect 1264 2119 1265 2123
rect 1286 2120 1287 2124
rect 1291 2120 1292 2124
rect 1286 2119 1292 2120
rect 1326 2124 1332 2125
rect 2502 2124 2508 2125
rect 1326 2120 1327 2124
rect 1331 2120 1332 2124
rect 1326 2119 1332 2120
rect 1678 2123 1684 2124
rect 1678 2119 1679 2123
rect 1683 2119 1684 2123
rect 1254 2118 1265 2119
rect 1678 2118 1684 2119
rect 1699 2123 1705 2124
rect 1699 2119 1700 2123
rect 1704 2122 1705 2123
rect 1734 2123 1740 2124
rect 1704 2120 1730 2122
rect 1704 2119 1705 2120
rect 1699 2118 1705 2119
rect 1728 2110 1730 2120
rect 1734 2119 1735 2123
rect 1739 2119 1740 2123
rect 1734 2118 1740 2119
rect 1755 2123 1761 2124
rect 1755 2119 1756 2123
rect 1760 2122 1761 2123
rect 1806 2123 1812 2124
rect 1760 2120 1802 2122
rect 1760 2119 1761 2120
rect 1755 2118 1761 2119
rect 1800 2110 1802 2120
rect 1806 2119 1807 2123
rect 1811 2119 1812 2123
rect 1806 2118 1812 2119
rect 1826 2123 1833 2124
rect 1826 2119 1827 2123
rect 1832 2119 1833 2123
rect 1826 2118 1833 2119
rect 1886 2123 1892 2124
rect 1886 2119 1887 2123
rect 1891 2119 1892 2123
rect 1907 2123 1913 2124
rect 1907 2122 1908 2123
rect 1886 2118 1892 2119
rect 1896 2120 1908 2122
rect 1896 2114 1898 2120
rect 1907 2119 1908 2120
rect 1912 2119 1913 2123
rect 1907 2118 1913 2119
rect 1982 2123 1988 2124
rect 1982 2119 1983 2123
rect 1987 2119 1988 2123
rect 1982 2118 1988 2119
rect 1990 2123 1996 2124
rect 1990 2119 1991 2123
rect 1995 2122 1996 2123
rect 2003 2123 2009 2124
rect 2003 2122 2004 2123
rect 1995 2120 2004 2122
rect 1995 2119 1996 2120
rect 1990 2118 1996 2119
rect 2003 2119 2004 2120
rect 2008 2119 2009 2123
rect 2003 2118 2009 2119
rect 2094 2123 2100 2124
rect 2094 2119 2095 2123
rect 2099 2119 2100 2123
rect 2115 2123 2121 2124
rect 2115 2122 2116 2123
rect 2094 2118 2100 2119
rect 2104 2120 2116 2122
rect 2104 2114 2106 2120
rect 2115 2119 2116 2120
rect 2120 2119 2121 2123
rect 2115 2118 2121 2119
rect 2214 2123 2220 2124
rect 2214 2119 2215 2123
rect 2219 2119 2220 2123
rect 2235 2123 2241 2124
rect 2235 2122 2236 2123
rect 2214 2118 2220 2119
rect 2224 2120 2236 2122
rect 2224 2114 2226 2120
rect 2235 2119 2236 2120
rect 2240 2119 2241 2123
rect 2235 2118 2241 2119
rect 2342 2123 2348 2124
rect 2342 2119 2343 2123
rect 2347 2119 2348 2123
rect 2342 2118 2348 2119
rect 2363 2123 2369 2124
rect 2363 2119 2364 2123
rect 2368 2122 2369 2123
rect 2454 2123 2460 2124
rect 2368 2120 2450 2122
rect 2368 2119 2369 2120
rect 2363 2118 2369 2119
rect 1820 2112 1898 2114
rect 1988 2112 2106 2114
rect 2108 2112 2226 2114
rect 1728 2109 1745 2110
rect 1728 2108 1740 2109
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 1286 2107 1292 2108
rect 110 2102 116 2103
rect 398 2104 404 2105
rect 398 2100 399 2104
rect 403 2100 404 2104
rect 398 2099 404 2100
rect 494 2104 500 2105
rect 494 2100 495 2104
rect 499 2100 500 2104
rect 494 2099 500 2100
rect 590 2104 596 2105
rect 590 2100 591 2104
rect 595 2100 596 2104
rect 590 2099 596 2100
rect 694 2104 700 2105
rect 694 2100 695 2104
rect 699 2100 700 2104
rect 694 2099 700 2100
rect 798 2104 804 2105
rect 798 2100 799 2104
rect 803 2100 804 2104
rect 798 2099 804 2100
rect 910 2104 916 2105
rect 910 2100 911 2104
rect 915 2100 916 2104
rect 910 2099 916 2100
rect 1022 2104 1028 2105
rect 1022 2100 1023 2104
rect 1027 2100 1028 2104
rect 1022 2099 1028 2100
rect 1134 2104 1140 2105
rect 1134 2100 1135 2104
rect 1139 2100 1140 2104
rect 1134 2099 1140 2100
rect 1222 2104 1228 2105
rect 1222 2100 1223 2104
rect 1227 2100 1228 2104
rect 1286 2103 1287 2107
rect 1291 2103 1292 2107
rect 1286 2102 1292 2103
rect 1683 2107 1689 2108
rect 1683 2103 1684 2107
rect 1688 2106 1689 2107
rect 1688 2104 1734 2106
rect 1739 2105 1740 2108
rect 1744 2105 1745 2109
rect 1800 2109 1817 2110
rect 1800 2108 1812 2109
rect 1739 2104 1745 2105
rect 1811 2105 1812 2108
rect 1816 2105 1817 2109
rect 1811 2104 1817 2105
rect 1688 2103 1689 2104
rect 1683 2102 1689 2103
rect 1732 2102 1734 2104
rect 1820 2102 1822 2112
rect 1988 2110 1990 2112
rect 2108 2110 2110 2112
rect 1987 2109 1993 2110
rect 1891 2107 1897 2108
rect 1891 2103 1892 2107
rect 1896 2106 1897 2107
rect 1896 2104 1946 2106
rect 1987 2105 1988 2109
rect 1992 2105 1993 2109
rect 1987 2104 1993 2105
rect 2099 2109 2110 2110
rect 2099 2105 2100 2109
rect 2104 2108 2110 2109
rect 2448 2110 2450 2120
rect 2454 2119 2455 2123
rect 2459 2119 2460 2123
rect 2454 2118 2460 2119
rect 2462 2123 2468 2124
rect 2462 2119 2463 2123
rect 2467 2122 2468 2123
rect 2475 2123 2481 2124
rect 2475 2122 2476 2123
rect 2467 2120 2476 2122
rect 2467 2119 2468 2120
rect 2462 2118 2468 2119
rect 2475 2119 2476 2120
rect 2480 2119 2481 2123
rect 2502 2120 2503 2124
rect 2507 2120 2508 2124
rect 2502 2119 2508 2120
rect 2475 2118 2481 2119
rect 2448 2109 2465 2110
rect 2448 2108 2460 2109
rect 2104 2105 2105 2108
rect 2099 2104 2105 2105
rect 2219 2107 2225 2108
rect 1896 2103 1897 2104
rect 1891 2102 1897 2103
rect 1944 2102 1946 2104
rect 2219 2103 2220 2107
rect 2224 2106 2225 2107
rect 2334 2107 2340 2108
rect 2334 2106 2335 2107
rect 2224 2104 2335 2106
rect 2224 2103 2225 2104
rect 2219 2102 2225 2103
rect 2334 2103 2335 2104
rect 2339 2103 2340 2107
rect 2334 2102 2340 2103
rect 2347 2107 2353 2108
rect 2347 2103 2348 2107
rect 2352 2106 2353 2107
rect 2352 2104 2414 2106
rect 2459 2105 2460 2108
rect 2464 2105 2465 2109
rect 2459 2104 2465 2105
rect 2352 2103 2353 2104
rect 2347 2102 2353 2103
rect 2412 2102 2414 2104
rect 2470 2103 2476 2104
rect 2470 2102 2471 2103
rect 1732 2100 1822 2102
rect 1944 2100 1994 2102
rect 2412 2100 2471 2102
rect 1222 2099 1228 2100
rect 1990 2099 1996 2100
rect 1990 2095 1991 2099
rect 1995 2095 1996 2099
rect 2470 2099 2471 2100
rect 2475 2099 2476 2103
rect 2470 2098 2476 2099
rect 1990 2094 1996 2095
rect 374 2092 380 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 446 2092 452 2093
rect 446 2088 447 2092
rect 451 2088 452 2092
rect 446 2087 452 2088
rect 518 2092 524 2093
rect 518 2088 519 2092
rect 523 2088 524 2092
rect 518 2087 524 2088
rect 598 2092 604 2093
rect 598 2088 599 2092
rect 603 2088 604 2092
rect 598 2087 604 2088
rect 678 2092 684 2093
rect 678 2088 679 2092
rect 683 2088 684 2092
rect 678 2087 684 2088
rect 758 2092 764 2093
rect 758 2088 759 2092
rect 763 2088 764 2092
rect 758 2087 764 2088
rect 830 2092 836 2093
rect 830 2088 831 2092
rect 835 2088 836 2092
rect 830 2087 836 2088
rect 902 2092 908 2093
rect 902 2088 903 2092
rect 907 2088 908 2092
rect 902 2087 908 2088
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 1030 2092 1036 2093
rect 1030 2088 1031 2092
rect 1035 2088 1036 2092
rect 1030 2087 1036 2088
rect 1102 2092 1108 2093
rect 1102 2088 1103 2092
rect 1107 2088 1108 2092
rect 1102 2087 1108 2088
rect 1166 2092 1172 2093
rect 1166 2088 1167 2092
rect 1171 2088 1172 2092
rect 1166 2087 1172 2088
rect 1222 2092 1228 2093
rect 1222 2088 1223 2092
rect 1227 2088 1228 2092
rect 1222 2087 1228 2088
rect 1286 2089 1292 2090
rect 110 2084 116 2085
rect 1286 2085 1287 2089
rect 1291 2085 1292 2089
rect 1286 2084 1292 2085
rect 1858 2083 1864 2084
rect 1858 2082 1859 2083
rect 1788 2080 1859 2082
rect 1788 2078 1790 2080
rect 1858 2079 1859 2080
rect 1863 2079 1864 2083
rect 1858 2078 1864 2079
rect 1260 2077 1377 2078
rect 1260 2076 1372 2077
rect 1260 2074 1262 2076
rect 1259 2073 1265 2074
rect 1371 2073 1372 2076
rect 1376 2073 1377 2077
rect 1787 2077 1793 2078
rect 1427 2075 1433 2076
rect 1427 2074 1428 2075
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 390 2071 396 2072
rect 390 2067 391 2071
rect 395 2067 396 2071
rect 390 2066 396 2067
rect 411 2071 417 2072
rect 411 2067 412 2071
rect 416 2070 417 2071
rect 454 2071 460 2072
rect 454 2070 455 2071
rect 416 2068 455 2070
rect 416 2067 417 2068
rect 411 2066 417 2067
rect 454 2067 455 2068
rect 459 2067 460 2071
rect 454 2066 460 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 478 2071 489 2072
rect 478 2067 479 2071
rect 483 2067 484 2071
rect 488 2067 489 2071
rect 478 2066 489 2067
rect 534 2071 540 2072
rect 534 2067 535 2071
rect 539 2067 540 2071
rect 555 2071 561 2072
rect 555 2070 556 2071
rect 534 2066 540 2067
rect 544 2068 556 2070
rect 544 2062 546 2068
rect 555 2067 556 2068
rect 560 2067 561 2071
rect 555 2066 561 2067
rect 614 2071 620 2072
rect 614 2067 615 2071
rect 619 2067 620 2071
rect 614 2066 620 2067
rect 630 2071 641 2072
rect 630 2067 631 2071
rect 635 2067 636 2071
rect 640 2067 641 2071
rect 630 2066 641 2067
rect 694 2071 700 2072
rect 694 2067 695 2071
rect 699 2067 700 2071
rect 715 2071 721 2072
rect 715 2070 716 2071
rect 694 2066 700 2067
rect 704 2068 716 2070
rect 704 2062 706 2068
rect 715 2067 716 2068
rect 720 2067 721 2071
rect 715 2066 721 2067
rect 774 2071 780 2072
rect 774 2067 775 2071
rect 779 2067 780 2071
rect 774 2066 780 2067
rect 795 2071 801 2072
rect 795 2067 796 2071
rect 800 2070 801 2071
rect 846 2071 852 2072
rect 800 2068 842 2070
rect 800 2067 801 2068
rect 795 2066 801 2067
rect 822 2063 828 2064
rect 822 2062 823 2063
rect 468 2060 546 2062
rect 620 2060 706 2062
rect 708 2060 823 2062
rect 468 2058 470 2060
rect 620 2058 622 2060
rect 708 2058 710 2060
rect 822 2059 823 2060
rect 827 2059 828 2063
rect 822 2058 828 2059
rect 840 2058 842 2068
rect 846 2067 847 2071
rect 851 2067 852 2071
rect 846 2066 852 2067
rect 867 2071 873 2072
rect 867 2067 868 2071
rect 872 2067 873 2071
rect 867 2066 873 2067
rect 918 2071 924 2072
rect 918 2067 919 2071
rect 923 2067 924 2071
rect 918 2066 924 2067
rect 939 2071 945 2072
rect 939 2067 940 2071
rect 944 2070 945 2071
rect 982 2071 988 2072
rect 944 2068 974 2070
rect 944 2067 945 2068
rect 939 2066 945 2067
rect 869 2058 871 2066
rect 972 2058 974 2068
rect 982 2067 983 2071
rect 987 2067 988 2071
rect 982 2066 988 2067
rect 1003 2071 1009 2072
rect 1003 2067 1004 2071
rect 1008 2070 1009 2071
rect 1046 2071 1052 2072
rect 1008 2068 1038 2070
rect 1008 2067 1009 2068
rect 1003 2066 1009 2067
rect 1036 2058 1038 2068
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1067 2071 1073 2072
rect 1067 2067 1068 2071
rect 1072 2070 1073 2071
rect 1118 2071 1124 2072
rect 1072 2068 1114 2070
rect 1072 2067 1073 2068
rect 1067 2066 1073 2067
rect 1112 2058 1114 2068
rect 1118 2067 1119 2071
rect 1123 2067 1124 2071
rect 1118 2066 1124 2067
rect 1126 2071 1132 2072
rect 1126 2067 1127 2071
rect 1131 2070 1132 2071
rect 1139 2071 1145 2072
rect 1139 2070 1140 2071
rect 1131 2068 1140 2070
rect 1131 2067 1132 2068
rect 1126 2066 1132 2067
rect 1139 2067 1140 2068
rect 1144 2067 1145 2071
rect 1139 2066 1145 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 1203 2071 1209 2072
rect 1203 2067 1204 2071
rect 1208 2070 1209 2071
rect 1238 2071 1244 2072
rect 1208 2068 1234 2070
rect 1208 2067 1209 2068
rect 1203 2066 1209 2067
rect 1232 2058 1234 2068
rect 1238 2067 1239 2071
rect 1243 2067 1244 2071
rect 1259 2069 1260 2073
rect 1264 2069 1265 2073
rect 1259 2068 1265 2069
rect 1286 2072 1292 2073
rect 1371 2072 1377 2073
rect 1388 2072 1428 2074
rect 1286 2068 1287 2072
rect 1291 2068 1292 2072
rect 1286 2067 1292 2068
rect 1238 2066 1244 2067
rect 1388 2062 1390 2072
rect 1427 2071 1428 2072
rect 1432 2071 1433 2075
rect 1507 2075 1513 2076
rect 1507 2074 1508 2075
rect 1427 2070 1433 2071
rect 1444 2072 1508 2074
rect 1444 2062 1446 2072
rect 1507 2071 1508 2072
rect 1512 2071 1513 2075
rect 1595 2075 1601 2076
rect 1595 2074 1596 2075
rect 1507 2070 1513 2071
rect 1524 2072 1596 2074
rect 1524 2062 1526 2072
rect 1595 2071 1596 2072
rect 1600 2071 1601 2075
rect 1683 2075 1689 2076
rect 1683 2074 1684 2075
rect 1595 2070 1601 2071
rect 1612 2072 1684 2074
rect 1612 2062 1614 2072
rect 1683 2071 1684 2072
rect 1688 2071 1689 2075
rect 1787 2073 1788 2077
rect 1792 2073 1793 2077
rect 1899 2075 1905 2076
rect 1899 2074 1900 2075
rect 1787 2072 1793 2073
rect 1804 2072 1900 2074
rect 1683 2070 1689 2071
rect 1804 2062 1806 2072
rect 1899 2071 1900 2072
rect 1904 2071 1905 2075
rect 2027 2075 2033 2076
rect 2027 2074 2028 2075
rect 1899 2070 1905 2071
rect 1916 2072 2028 2074
rect 1916 2062 1918 2072
rect 2027 2071 2028 2072
rect 2032 2071 2033 2075
rect 2171 2075 2177 2076
rect 2171 2074 2172 2075
rect 2027 2070 2033 2071
rect 2044 2072 2172 2074
rect 2044 2062 2046 2072
rect 2171 2071 2172 2072
rect 2176 2071 2177 2075
rect 2323 2075 2329 2076
rect 2323 2074 2324 2075
rect 2171 2070 2177 2071
rect 2188 2072 2324 2074
rect 2188 2062 2190 2072
rect 2323 2071 2324 2072
rect 2328 2071 2329 2075
rect 2323 2070 2329 2071
rect 2459 2075 2468 2076
rect 2459 2071 2460 2075
rect 2467 2071 2468 2075
rect 2459 2070 2468 2071
rect 1366 2061 1372 2062
rect 1326 2060 1332 2061
rect 467 2057 473 2058
rect 395 2055 401 2056
rect 395 2051 396 2055
rect 400 2054 401 2055
rect 400 2052 442 2054
rect 467 2053 468 2057
rect 472 2053 473 2057
rect 619 2057 625 2058
rect 467 2052 473 2053
rect 539 2055 545 2056
rect 400 2051 401 2052
rect 395 2050 401 2051
rect 440 2050 442 2052
rect 478 2051 484 2052
rect 478 2050 479 2051
rect 440 2048 479 2050
rect 478 2047 479 2048
rect 483 2047 484 2051
rect 539 2051 540 2055
rect 544 2054 545 2055
rect 544 2052 590 2054
rect 619 2053 620 2057
rect 624 2053 625 2057
rect 619 2052 625 2053
rect 699 2057 710 2058
rect 699 2053 700 2057
rect 704 2056 710 2057
rect 840 2057 857 2058
rect 840 2056 852 2057
rect 704 2053 705 2056
rect 699 2052 705 2053
rect 779 2055 785 2056
rect 544 2051 545 2052
rect 539 2050 545 2051
rect 588 2050 590 2052
rect 630 2051 636 2052
rect 630 2050 631 2051
rect 588 2048 631 2050
rect 478 2046 484 2047
rect 630 2047 631 2048
rect 635 2047 636 2051
rect 779 2051 780 2055
rect 784 2054 785 2055
rect 784 2052 846 2054
rect 851 2053 852 2056
rect 856 2053 857 2057
rect 869 2057 929 2058
rect 869 2056 924 2057
rect 851 2052 857 2053
rect 923 2053 924 2056
rect 928 2053 929 2057
rect 972 2057 993 2058
rect 972 2056 988 2057
rect 923 2052 929 2053
rect 987 2053 988 2056
rect 992 2053 993 2057
rect 1036 2057 1057 2058
rect 1036 2056 1052 2057
rect 987 2052 993 2053
rect 1051 2053 1052 2056
rect 1056 2053 1057 2057
rect 1112 2057 1129 2058
rect 1112 2056 1124 2057
rect 1051 2052 1057 2053
rect 1123 2053 1124 2056
rect 1128 2053 1129 2057
rect 1232 2057 1249 2058
rect 1232 2056 1244 2057
rect 1123 2052 1129 2053
rect 1187 2055 1193 2056
rect 784 2051 785 2052
rect 779 2050 785 2051
rect 844 2050 846 2052
rect 1082 2051 1088 2052
rect 1082 2050 1083 2051
rect 844 2048 1083 2050
rect 630 2046 636 2047
rect 1082 2047 1083 2048
rect 1087 2047 1088 2051
rect 1187 2051 1188 2055
rect 1192 2054 1193 2055
rect 1192 2052 1226 2054
rect 1243 2053 1244 2056
rect 1248 2053 1249 2057
rect 1326 2056 1327 2060
rect 1331 2056 1332 2060
rect 1366 2057 1367 2061
rect 1371 2057 1372 2061
rect 1366 2056 1372 2057
rect 1387 2061 1393 2062
rect 1387 2057 1388 2061
rect 1392 2057 1393 2061
rect 1387 2056 1393 2057
rect 1422 2061 1428 2062
rect 1422 2057 1423 2061
rect 1427 2057 1428 2061
rect 1422 2056 1428 2057
rect 1443 2061 1449 2062
rect 1443 2057 1444 2061
rect 1448 2057 1449 2061
rect 1443 2056 1449 2057
rect 1502 2061 1508 2062
rect 1502 2057 1503 2061
rect 1507 2057 1508 2061
rect 1502 2056 1508 2057
rect 1523 2061 1529 2062
rect 1523 2057 1524 2061
rect 1528 2057 1529 2061
rect 1523 2056 1529 2057
rect 1590 2061 1596 2062
rect 1590 2057 1591 2061
rect 1595 2057 1596 2061
rect 1590 2056 1596 2057
rect 1611 2061 1617 2062
rect 1611 2057 1612 2061
rect 1616 2057 1617 2061
rect 1611 2056 1617 2057
rect 1678 2061 1684 2062
rect 1678 2057 1679 2061
rect 1683 2057 1684 2061
rect 1782 2061 1788 2062
rect 1678 2056 1684 2057
rect 1686 2059 1692 2060
rect 1326 2055 1332 2056
rect 1686 2055 1687 2059
rect 1691 2058 1692 2059
rect 1699 2059 1705 2060
rect 1699 2058 1700 2059
rect 1691 2056 1700 2058
rect 1691 2055 1692 2056
rect 1686 2054 1692 2055
rect 1699 2055 1700 2056
rect 1704 2055 1705 2059
rect 1782 2057 1783 2061
rect 1787 2057 1788 2061
rect 1782 2056 1788 2057
rect 1803 2061 1809 2062
rect 1803 2057 1804 2061
rect 1808 2057 1809 2061
rect 1803 2056 1809 2057
rect 1894 2061 1900 2062
rect 1894 2057 1895 2061
rect 1899 2057 1900 2061
rect 1894 2056 1900 2057
rect 1915 2061 1921 2062
rect 1915 2057 1916 2061
rect 1920 2057 1921 2061
rect 1915 2056 1921 2057
rect 2022 2061 2028 2062
rect 2022 2057 2023 2061
rect 2027 2057 2028 2061
rect 2022 2056 2028 2057
rect 2043 2061 2049 2062
rect 2043 2057 2044 2061
rect 2048 2057 2049 2061
rect 2043 2056 2049 2057
rect 2166 2061 2172 2062
rect 2166 2057 2167 2061
rect 2171 2057 2172 2061
rect 2166 2056 2172 2057
rect 2187 2061 2193 2062
rect 2187 2057 2188 2061
rect 2192 2057 2193 2061
rect 2187 2056 2193 2057
rect 2318 2061 2324 2062
rect 2318 2057 2319 2061
rect 2323 2057 2324 2061
rect 2454 2061 2460 2062
rect 2318 2056 2324 2057
rect 2334 2059 2345 2060
rect 1699 2054 1705 2055
rect 2334 2055 2335 2059
rect 2339 2055 2340 2059
rect 2344 2055 2345 2059
rect 2454 2057 2455 2061
rect 2459 2057 2460 2061
rect 2502 2060 2508 2061
rect 2454 2056 2460 2057
rect 2470 2059 2481 2060
rect 2334 2054 2345 2055
rect 2470 2055 2471 2059
rect 2475 2055 2476 2059
rect 2480 2055 2481 2059
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2470 2054 2481 2055
rect 1243 2052 1249 2053
rect 1192 2051 1193 2052
rect 1187 2050 1193 2051
rect 1224 2050 1226 2052
rect 1254 2051 1260 2052
rect 1254 2050 1255 2051
rect 1224 2048 1255 2050
rect 1082 2046 1088 2047
rect 1254 2047 1255 2048
rect 1259 2047 1260 2051
rect 1254 2046 1260 2047
rect 1326 2043 1332 2044
rect 658 2039 664 2040
rect 658 2038 659 2039
rect 300 2036 659 2038
rect 300 2034 302 2036
rect 658 2035 659 2036
rect 663 2035 664 2039
rect 1326 2039 1327 2043
rect 1331 2039 1332 2043
rect 2502 2043 2508 2044
rect 1326 2038 1332 2039
rect 1350 2040 1356 2041
rect 1350 2036 1351 2040
rect 1355 2036 1356 2040
rect 1350 2035 1356 2036
rect 1406 2040 1412 2041
rect 1406 2036 1407 2040
rect 1411 2036 1412 2040
rect 1406 2035 1412 2036
rect 1486 2040 1492 2041
rect 1486 2036 1487 2040
rect 1491 2036 1492 2040
rect 1486 2035 1492 2036
rect 1574 2040 1580 2041
rect 1574 2036 1575 2040
rect 1579 2036 1580 2040
rect 1574 2035 1580 2036
rect 1662 2040 1668 2041
rect 1662 2036 1663 2040
rect 1667 2036 1668 2040
rect 1662 2035 1668 2036
rect 1766 2040 1772 2041
rect 1766 2036 1767 2040
rect 1771 2036 1772 2040
rect 1766 2035 1772 2036
rect 1878 2040 1884 2041
rect 1878 2036 1879 2040
rect 1883 2036 1884 2040
rect 1878 2035 1884 2036
rect 2006 2040 2012 2041
rect 2006 2036 2007 2040
rect 2011 2036 2012 2040
rect 2006 2035 2012 2036
rect 2150 2040 2156 2041
rect 2150 2036 2151 2040
rect 2155 2036 2156 2040
rect 2150 2035 2156 2036
rect 2302 2040 2308 2041
rect 2302 2036 2303 2040
rect 2307 2036 2308 2040
rect 2302 2035 2308 2036
rect 2438 2040 2444 2041
rect 2438 2036 2439 2040
rect 2443 2036 2444 2040
rect 2502 2039 2503 2043
rect 2507 2039 2508 2043
rect 2502 2038 2508 2039
rect 2438 2035 2444 2036
rect 658 2034 664 2035
rect 299 2033 305 2034
rect 299 2029 300 2033
rect 304 2029 305 2033
rect 379 2031 385 2032
rect 379 2030 380 2031
rect 299 2028 305 2029
rect 319 2028 380 2030
rect 319 2018 321 2028
rect 379 2027 380 2028
rect 384 2027 385 2031
rect 379 2026 385 2027
rect 454 2031 460 2032
rect 454 2027 455 2031
rect 459 2030 460 2031
rect 467 2031 473 2032
rect 467 2030 468 2031
rect 459 2028 468 2030
rect 459 2027 460 2028
rect 454 2026 460 2027
rect 467 2027 468 2028
rect 472 2027 473 2031
rect 555 2031 561 2032
rect 555 2030 556 2031
rect 467 2026 473 2027
rect 484 2028 556 2030
rect 484 2018 486 2028
rect 555 2027 556 2028
rect 560 2027 561 2031
rect 643 2031 649 2032
rect 643 2030 644 2031
rect 555 2026 561 2027
rect 572 2028 644 2030
rect 572 2018 574 2028
rect 643 2027 644 2028
rect 648 2027 649 2031
rect 643 2026 649 2027
rect 723 2031 732 2032
rect 723 2027 724 2031
rect 731 2027 732 2031
rect 803 2031 809 2032
rect 803 2030 804 2031
rect 723 2026 732 2027
rect 740 2028 804 2030
rect 740 2018 742 2028
rect 803 2027 804 2028
rect 808 2027 809 2031
rect 891 2031 897 2032
rect 891 2030 892 2031
rect 803 2026 809 2027
rect 820 2028 892 2030
rect 820 2018 822 2028
rect 891 2027 892 2028
rect 896 2027 897 2031
rect 979 2031 985 2032
rect 979 2030 980 2031
rect 891 2026 897 2027
rect 908 2028 980 2030
rect 908 2018 910 2028
rect 979 2027 980 2028
rect 984 2027 985 2031
rect 1067 2031 1073 2032
rect 1067 2030 1068 2031
rect 979 2026 985 2027
rect 996 2028 1068 2030
rect 996 2018 998 2028
rect 1067 2027 1068 2028
rect 1072 2027 1073 2031
rect 1067 2026 1073 2027
rect 1350 2028 1356 2029
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1350 2024 1351 2028
rect 1355 2024 1356 2028
rect 1350 2023 1356 2024
rect 1422 2028 1428 2029
rect 1422 2024 1423 2028
rect 1427 2024 1428 2028
rect 1422 2023 1428 2024
rect 1518 2028 1524 2029
rect 1518 2024 1519 2028
rect 1523 2024 1524 2028
rect 1518 2023 1524 2024
rect 1614 2028 1620 2029
rect 1614 2024 1615 2028
rect 1619 2024 1620 2028
rect 1614 2023 1620 2024
rect 1718 2028 1724 2029
rect 1718 2024 1719 2028
rect 1723 2024 1724 2028
rect 1718 2023 1724 2024
rect 1822 2028 1828 2029
rect 1822 2024 1823 2028
rect 1827 2024 1828 2028
rect 1822 2023 1828 2024
rect 1934 2028 1940 2029
rect 1934 2024 1935 2028
rect 1939 2024 1940 2028
rect 1934 2023 1940 2024
rect 2054 2028 2060 2029
rect 2054 2024 2055 2028
rect 2059 2024 2060 2028
rect 2054 2023 2060 2024
rect 2182 2028 2188 2029
rect 2182 2024 2183 2028
rect 2187 2024 2188 2028
rect 2182 2023 2188 2024
rect 2318 2028 2324 2029
rect 2318 2024 2319 2028
rect 2323 2024 2324 2028
rect 2318 2023 2324 2024
rect 2438 2028 2444 2029
rect 2438 2024 2439 2028
rect 2443 2024 2444 2028
rect 2438 2023 2444 2024
rect 2502 2025 2508 2026
rect 1326 2020 1332 2021
rect 2502 2021 2503 2025
rect 2507 2021 2508 2025
rect 2502 2020 2508 2021
rect 294 2017 300 2018
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 294 2013 295 2017
rect 299 2013 300 2017
rect 294 2012 300 2013
rect 315 2017 321 2018
rect 315 2013 316 2017
rect 320 2013 321 2017
rect 315 2012 321 2013
rect 374 2017 380 2018
rect 374 2013 375 2017
rect 379 2013 380 2017
rect 462 2017 468 2018
rect 374 2012 380 2013
rect 395 2015 401 2016
rect 110 2011 116 2012
rect 395 2011 396 2015
rect 400 2014 401 2015
rect 406 2015 412 2016
rect 406 2014 407 2015
rect 400 2012 407 2014
rect 400 2011 401 2012
rect 395 2010 401 2011
rect 406 2011 407 2012
rect 411 2011 412 2015
rect 462 2013 463 2017
rect 467 2013 468 2017
rect 462 2012 468 2013
rect 483 2017 489 2018
rect 483 2013 484 2017
rect 488 2013 489 2017
rect 483 2012 489 2013
rect 550 2017 556 2018
rect 550 2013 551 2017
rect 555 2013 556 2017
rect 550 2012 556 2013
rect 571 2017 577 2018
rect 571 2013 572 2017
rect 576 2013 577 2017
rect 571 2012 577 2013
rect 638 2017 644 2018
rect 638 2013 639 2017
rect 643 2013 644 2017
rect 718 2017 724 2018
rect 638 2012 644 2013
rect 658 2015 665 2016
rect 406 2010 412 2011
rect 658 2011 659 2015
rect 664 2011 665 2015
rect 718 2013 719 2017
rect 723 2013 724 2017
rect 718 2012 724 2013
rect 739 2017 745 2018
rect 739 2013 740 2017
rect 744 2013 745 2017
rect 739 2012 745 2013
rect 798 2017 804 2018
rect 798 2013 799 2017
rect 803 2013 804 2017
rect 798 2012 804 2013
rect 819 2017 825 2018
rect 819 2013 820 2017
rect 824 2013 825 2017
rect 819 2012 825 2013
rect 886 2017 892 2018
rect 886 2013 887 2017
rect 891 2013 892 2017
rect 886 2012 892 2013
rect 907 2017 913 2018
rect 907 2013 908 2017
rect 912 2013 913 2017
rect 907 2012 913 2013
rect 974 2017 980 2018
rect 974 2013 975 2017
rect 979 2013 980 2017
rect 974 2012 980 2013
rect 995 2017 1001 2018
rect 995 2013 996 2017
rect 1000 2013 1001 2017
rect 995 2012 1001 2013
rect 1062 2017 1068 2018
rect 1062 2013 1063 2017
rect 1067 2013 1068 2017
rect 1286 2016 1292 2017
rect 1062 2012 1068 2013
rect 1082 2015 1089 2016
rect 658 2010 665 2011
rect 1082 2011 1083 2015
rect 1088 2011 1089 2015
rect 1286 2012 1287 2016
rect 1291 2012 1292 2016
rect 1286 2011 1292 2012
rect 1082 2010 1089 2011
rect 1326 2008 1332 2009
rect 2502 2008 2508 2009
rect 1326 2004 1327 2008
rect 1331 2004 1332 2008
rect 1326 2003 1332 2004
rect 1366 2007 1372 2008
rect 1366 2003 1367 2007
rect 1371 2003 1372 2007
rect 1366 2002 1372 2003
rect 1387 2007 1393 2008
rect 1387 2003 1388 2007
rect 1392 2006 1393 2007
rect 1438 2007 1444 2008
rect 1392 2004 1434 2006
rect 1392 2003 1393 2004
rect 1387 2002 1393 2003
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 1286 1999 1292 2000
rect 110 1994 116 1995
rect 278 1996 284 1997
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 358 1996 364 1997
rect 358 1992 359 1996
rect 363 1992 364 1996
rect 358 1991 364 1992
rect 446 1996 452 1997
rect 446 1992 447 1996
rect 451 1992 452 1996
rect 446 1991 452 1992
rect 534 1996 540 1997
rect 534 1992 535 1996
rect 539 1992 540 1996
rect 534 1991 540 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 702 1996 708 1997
rect 702 1992 703 1996
rect 707 1992 708 1996
rect 702 1991 708 1992
rect 782 1996 788 1997
rect 782 1992 783 1996
rect 787 1992 788 1996
rect 782 1991 788 1992
rect 870 1996 876 1997
rect 870 1992 871 1996
rect 875 1992 876 1996
rect 870 1991 876 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1286 1995 1287 1999
rect 1291 1995 1292 1999
rect 1286 1994 1292 1995
rect 1432 1994 1434 2004
rect 1438 2003 1439 2007
rect 1443 2003 1444 2007
rect 1438 2002 1444 2003
rect 1459 2007 1465 2008
rect 1459 2003 1460 2007
rect 1464 2006 1465 2007
rect 1534 2007 1540 2008
rect 1464 2004 1530 2006
rect 1464 2003 1465 2004
rect 1459 2002 1465 2003
rect 1528 1994 1530 2004
rect 1534 2003 1535 2007
rect 1539 2003 1540 2007
rect 1534 2002 1540 2003
rect 1555 2007 1561 2008
rect 1555 2003 1556 2007
rect 1560 2006 1561 2007
rect 1630 2007 1636 2008
rect 1560 2004 1626 2006
rect 1560 2003 1561 2004
rect 1555 2002 1561 2003
rect 1624 1994 1626 2004
rect 1630 2003 1631 2007
rect 1635 2003 1636 2007
rect 1630 2002 1636 2003
rect 1651 2007 1657 2008
rect 1651 2003 1652 2007
rect 1656 2006 1657 2007
rect 1734 2007 1740 2008
rect 1656 2004 1730 2006
rect 1656 2003 1657 2004
rect 1651 2002 1657 2003
rect 1728 1994 1730 2004
rect 1734 2003 1735 2007
rect 1739 2003 1740 2007
rect 1734 2002 1740 2003
rect 1742 2007 1748 2008
rect 1742 2003 1743 2007
rect 1747 2006 1748 2007
rect 1755 2007 1761 2008
rect 1755 2006 1756 2007
rect 1747 2004 1756 2006
rect 1747 2003 1748 2004
rect 1742 2002 1748 2003
rect 1755 2003 1756 2004
rect 1760 2003 1761 2007
rect 1755 2002 1761 2003
rect 1838 2007 1844 2008
rect 1838 2003 1839 2007
rect 1843 2003 1844 2007
rect 1838 2002 1844 2003
rect 1858 2007 1865 2008
rect 1858 2003 1859 2007
rect 1864 2003 1865 2007
rect 1858 2002 1865 2003
rect 1950 2007 1956 2008
rect 1950 2003 1951 2007
rect 1955 2003 1956 2007
rect 1950 2002 1956 2003
rect 1966 2007 1977 2008
rect 1966 2003 1967 2007
rect 1971 2003 1972 2007
rect 1976 2003 1977 2007
rect 1966 2002 1977 2003
rect 2070 2007 2076 2008
rect 2070 2003 2071 2007
rect 2075 2003 2076 2007
rect 2091 2007 2097 2008
rect 2091 2006 2092 2007
rect 2070 2002 2076 2003
rect 2080 2004 2092 2006
rect 2080 1998 2082 2004
rect 2091 2003 2092 2004
rect 2096 2003 2097 2007
rect 2091 2002 2097 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2219 2007 2225 2008
rect 2219 2003 2220 2007
rect 2224 2006 2225 2007
rect 2334 2007 2340 2008
rect 2224 2004 2326 2006
rect 2224 2003 2225 2004
rect 2219 2002 2225 2003
rect 1956 1996 2082 1998
rect 2114 1999 2120 2000
rect 1956 1994 1958 1996
rect 2114 1995 2115 1999
rect 2119 1998 2120 1999
rect 2310 1999 2316 2000
rect 2310 1998 2311 1999
rect 2119 1996 2311 1998
rect 2119 1995 2120 1996
rect 2114 1994 2120 1995
rect 2310 1995 2311 1996
rect 2315 1995 2316 1999
rect 2310 1994 2316 1995
rect 2324 1994 2326 2004
rect 2334 2003 2335 2007
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2342 2007 2348 2008
rect 2342 2003 2343 2007
rect 2347 2006 2348 2007
rect 2355 2007 2361 2008
rect 2355 2006 2356 2007
rect 2347 2004 2356 2006
rect 2347 2003 2348 2004
rect 2342 2002 2348 2003
rect 2355 2003 2356 2004
rect 2360 2003 2361 2007
rect 2355 2002 2361 2003
rect 2454 2007 2460 2008
rect 2454 2003 2455 2007
rect 2459 2003 2460 2007
rect 2454 2002 2460 2003
rect 2462 2007 2468 2008
rect 2462 2003 2463 2007
rect 2467 2006 2468 2007
rect 2475 2007 2481 2008
rect 2475 2006 2476 2007
rect 2467 2004 2476 2006
rect 2467 2003 2468 2004
rect 2462 2002 2468 2003
rect 2475 2003 2476 2004
rect 2480 2003 2481 2007
rect 2502 2004 2503 2008
rect 2507 2004 2508 2008
rect 2502 2003 2508 2004
rect 2475 2002 2481 2003
rect 1432 1993 1449 1994
rect 1432 1992 1444 1993
rect 1046 1991 1052 1992
rect 1371 1991 1377 1992
rect 1371 1987 1372 1991
rect 1376 1990 1377 1991
rect 1376 1988 1438 1990
rect 1443 1989 1444 1992
rect 1448 1989 1449 1993
rect 1528 1993 1545 1994
rect 1528 1992 1540 1993
rect 1443 1988 1449 1989
rect 1539 1989 1540 1992
rect 1544 1989 1545 1993
rect 1624 1993 1641 1994
rect 1624 1992 1636 1993
rect 1539 1988 1545 1989
rect 1635 1989 1636 1992
rect 1640 1989 1641 1993
rect 1728 1993 1745 1994
rect 1728 1992 1740 1993
rect 1635 1988 1641 1989
rect 1739 1989 1740 1992
rect 1744 1989 1745 1993
rect 1955 1993 1961 1994
rect 1739 1988 1745 1989
rect 1843 1991 1849 1992
rect 1376 1987 1377 1988
rect 1371 1986 1377 1987
rect 1436 1986 1438 1988
rect 1686 1987 1692 1988
rect 1686 1986 1687 1987
rect 1436 1984 1687 1986
rect 1686 1983 1687 1984
rect 1691 1983 1692 1987
rect 1843 1987 1844 1991
rect 1848 1990 1849 1991
rect 1848 1988 1910 1990
rect 1955 1989 1956 1993
rect 1960 1989 1961 1993
rect 2324 1993 2345 1994
rect 2324 1992 2340 1993
rect 1955 1988 1961 1989
rect 2075 1991 2081 1992
rect 1848 1987 1849 1988
rect 1843 1986 1849 1987
rect 1908 1986 1910 1988
rect 1966 1987 1972 1988
rect 1966 1986 1967 1987
rect 1908 1984 1967 1986
rect 1686 1982 1692 1983
rect 1966 1983 1967 1984
rect 1971 1983 1972 1987
rect 2075 1987 2076 1991
rect 2080 1990 2081 1991
rect 2174 1991 2180 1992
rect 2080 1988 2170 1990
rect 2080 1987 2081 1988
rect 2075 1986 2081 1987
rect 1966 1982 1972 1983
rect 2168 1982 2170 1988
rect 2174 1987 2175 1991
rect 2179 1990 2180 1991
rect 2203 1991 2209 1992
rect 2203 1990 2204 1991
rect 2179 1988 2204 1990
rect 2179 1987 2180 1988
rect 2174 1986 2180 1987
rect 2203 1987 2204 1988
rect 2208 1987 2209 1991
rect 2339 1989 2340 1992
rect 2344 1989 2345 1993
rect 2339 1988 2345 1989
rect 2459 1991 2465 1992
rect 2203 1986 2209 1987
rect 2459 1987 2460 1991
rect 2464 1990 2465 1991
rect 2470 1991 2476 1992
rect 2470 1990 2471 1991
rect 2464 1988 2471 1990
rect 2464 1987 2465 1988
rect 2459 1986 2465 1987
rect 2470 1987 2471 1988
rect 2475 1987 2476 1991
rect 2470 1986 2476 1987
rect 2342 1983 2348 1984
rect 2342 1982 2343 1983
rect 134 1980 140 1981
rect 110 1977 116 1978
rect 110 1973 111 1977
rect 115 1973 116 1977
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 206 1980 212 1981
rect 206 1976 207 1980
rect 211 1976 212 1980
rect 206 1975 212 1976
rect 286 1980 292 1981
rect 286 1976 287 1980
rect 291 1976 292 1980
rect 286 1975 292 1976
rect 382 1980 388 1981
rect 382 1976 383 1980
rect 387 1976 388 1980
rect 382 1975 388 1976
rect 486 1980 492 1981
rect 486 1976 487 1980
rect 491 1976 492 1980
rect 486 1975 492 1976
rect 590 1980 596 1981
rect 590 1976 591 1980
rect 595 1976 596 1980
rect 590 1975 596 1976
rect 694 1980 700 1981
rect 694 1976 695 1980
rect 699 1976 700 1980
rect 694 1975 700 1976
rect 798 1980 804 1981
rect 798 1976 799 1980
rect 803 1976 804 1980
rect 798 1975 804 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1014 1980 1020 1981
rect 2168 1980 2343 1982
rect 1014 1976 1015 1980
rect 1019 1976 1020 1980
rect 2342 1979 2343 1980
rect 2347 1979 2348 1983
rect 2342 1978 2348 1979
rect 1014 1975 1020 1976
rect 1286 1977 1292 1978
rect 110 1972 116 1973
rect 1286 1973 1287 1977
rect 1291 1973 1292 1977
rect 1742 1975 1748 1976
rect 1742 1974 1743 1975
rect 1286 1972 1292 1973
rect 1460 1972 1743 1974
rect 1460 1970 1462 1972
rect 1742 1971 1743 1972
rect 1747 1971 1748 1975
rect 2114 1975 2120 1976
rect 2114 1974 2115 1975
rect 1742 1970 1748 1971
rect 1948 1972 2115 1974
rect 1948 1970 1950 1972
rect 2114 1971 2115 1972
rect 2119 1971 2120 1975
rect 2114 1970 2120 1971
rect 1459 1969 1465 1970
rect 1459 1965 1460 1969
rect 1464 1965 1465 1969
rect 1947 1969 1953 1970
rect 1547 1967 1553 1968
rect 1547 1966 1548 1967
rect 1459 1964 1465 1965
rect 1476 1964 1548 1966
rect 110 1960 116 1961
rect 1286 1960 1292 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 110 1955 116 1956
rect 150 1959 156 1960
rect 150 1955 151 1959
rect 155 1955 156 1959
rect 150 1954 156 1955
rect 171 1959 177 1960
rect 171 1955 172 1959
rect 176 1958 177 1959
rect 222 1959 228 1960
rect 176 1956 210 1958
rect 176 1955 177 1956
rect 171 1954 177 1955
rect 208 1946 210 1956
rect 222 1955 223 1959
rect 227 1955 228 1959
rect 222 1954 228 1955
rect 243 1959 249 1960
rect 243 1955 244 1959
rect 248 1955 249 1959
rect 243 1954 249 1955
rect 302 1959 308 1960
rect 302 1955 303 1959
rect 307 1955 308 1959
rect 302 1954 308 1955
rect 323 1959 329 1960
rect 323 1955 324 1959
rect 328 1958 329 1959
rect 366 1959 372 1960
rect 366 1958 367 1959
rect 328 1956 367 1958
rect 328 1955 329 1956
rect 323 1954 329 1955
rect 366 1955 367 1956
rect 371 1955 372 1959
rect 366 1954 372 1955
rect 398 1959 404 1960
rect 398 1955 399 1959
rect 403 1955 404 1959
rect 398 1954 404 1955
rect 419 1959 425 1960
rect 419 1955 420 1959
rect 424 1958 425 1959
rect 502 1959 508 1960
rect 424 1956 498 1958
rect 424 1955 425 1956
rect 419 1954 425 1955
rect 245 1946 247 1954
rect 496 1946 498 1956
rect 502 1955 503 1959
rect 507 1955 508 1959
rect 502 1954 508 1955
rect 523 1959 529 1960
rect 523 1955 524 1959
rect 528 1958 529 1959
rect 606 1959 612 1960
rect 528 1956 602 1958
rect 528 1955 529 1956
rect 523 1954 529 1955
rect 600 1946 602 1956
rect 606 1955 607 1959
rect 611 1955 612 1959
rect 606 1954 612 1955
rect 614 1959 620 1960
rect 614 1955 615 1959
rect 619 1958 620 1959
rect 627 1959 633 1960
rect 627 1958 628 1959
rect 619 1956 628 1958
rect 619 1955 620 1956
rect 614 1954 620 1955
rect 627 1955 628 1956
rect 632 1955 633 1959
rect 627 1954 633 1955
rect 710 1959 716 1960
rect 710 1955 711 1959
rect 715 1955 716 1959
rect 710 1954 716 1955
rect 726 1959 737 1960
rect 726 1955 727 1959
rect 731 1955 732 1959
rect 736 1955 737 1959
rect 726 1954 737 1955
rect 814 1959 820 1960
rect 814 1955 815 1959
rect 819 1955 820 1959
rect 835 1959 841 1960
rect 835 1958 836 1959
rect 814 1954 820 1955
rect 824 1956 836 1958
rect 824 1950 826 1956
rect 835 1955 836 1956
rect 840 1955 841 1959
rect 835 1954 841 1955
rect 918 1959 924 1960
rect 918 1955 919 1959
rect 923 1955 924 1959
rect 918 1954 924 1955
rect 939 1959 945 1960
rect 939 1955 940 1959
rect 944 1958 945 1959
rect 1030 1959 1036 1960
rect 944 1956 1026 1958
rect 944 1955 945 1956
rect 939 1954 945 1955
rect 716 1948 826 1950
rect 716 1946 718 1948
rect 1024 1946 1026 1956
rect 1030 1955 1031 1959
rect 1035 1955 1036 1959
rect 1030 1954 1036 1955
rect 1038 1959 1044 1960
rect 1038 1955 1039 1959
rect 1043 1958 1044 1959
rect 1051 1959 1057 1960
rect 1051 1958 1052 1959
rect 1043 1956 1052 1958
rect 1043 1955 1044 1956
rect 1038 1954 1044 1955
rect 1051 1955 1052 1956
rect 1056 1955 1057 1959
rect 1286 1956 1287 1960
rect 1291 1956 1292 1960
rect 1286 1955 1292 1956
rect 1051 1954 1057 1955
rect 1476 1954 1478 1964
rect 1547 1963 1548 1964
rect 1552 1963 1553 1967
rect 1643 1967 1649 1968
rect 1643 1966 1644 1967
rect 1547 1962 1553 1963
rect 1564 1964 1644 1966
rect 1564 1954 1566 1964
rect 1643 1963 1644 1964
rect 1648 1963 1649 1967
rect 1739 1967 1745 1968
rect 1739 1966 1740 1967
rect 1643 1962 1649 1963
rect 1660 1964 1740 1966
rect 1660 1954 1662 1964
rect 1739 1963 1740 1964
rect 1744 1963 1745 1967
rect 1843 1967 1849 1968
rect 1843 1966 1844 1967
rect 1739 1962 1745 1963
rect 1756 1964 1844 1966
rect 1756 1954 1758 1964
rect 1843 1963 1844 1964
rect 1848 1963 1849 1967
rect 1947 1965 1948 1969
rect 1952 1965 1953 1969
rect 2051 1967 2057 1968
rect 2051 1966 2052 1967
rect 1947 1964 1953 1965
rect 1999 1964 2052 1966
rect 1843 1962 1849 1963
rect 1999 1958 2001 1964
rect 2051 1963 2052 1964
rect 2056 1963 2057 1967
rect 2155 1967 2161 1968
rect 2155 1966 2156 1967
rect 2051 1962 2057 1963
rect 2068 1964 2156 1966
rect 1964 1956 2001 1958
rect 1964 1954 1966 1956
rect 2068 1954 2070 1964
rect 2155 1963 2156 1964
rect 2160 1963 2161 1967
rect 2155 1962 2161 1963
rect 2246 1967 2252 1968
rect 2246 1963 2247 1967
rect 2251 1966 2252 1967
rect 2259 1967 2265 1968
rect 2259 1966 2260 1967
rect 2251 1964 2260 1966
rect 2251 1963 2252 1964
rect 2246 1962 2252 1963
rect 2259 1963 2260 1964
rect 2264 1963 2265 1967
rect 2371 1967 2377 1968
rect 2371 1966 2372 1967
rect 2259 1962 2265 1963
rect 2276 1964 2372 1966
rect 2276 1954 2278 1964
rect 2371 1963 2372 1964
rect 2376 1963 2377 1967
rect 2371 1962 2377 1963
rect 2459 1967 2468 1968
rect 2459 1963 2460 1967
rect 2467 1963 2468 1967
rect 2459 1962 2468 1963
rect 2310 1959 2316 1960
rect 2310 1955 2311 1959
rect 2315 1958 2316 1959
rect 2315 1956 2390 1958
rect 2315 1955 2316 1956
rect 2310 1954 2316 1955
rect 2388 1954 2390 1956
rect 1454 1953 1460 1954
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1475 1953 1481 1954
rect 1475 1949 1476 1953
rect 1480 1949 1481 1953
rect 1475 1948 1481 1949
rect 1542 1953 1548 1954
rect 1542 1949 1543 1953
rect 1547 1949 1548 1953
rect 1542 1948 1548 1949
rect 1563 1953 1569 1954
rect 1563 1949 1564 1953
rect 1568 1949 1569 1953
rect 1563 1948 1569 1949
rect 1638 1953 1644 1954
rect 1638 1949 1639 1953
rect 1643 1949 1644 1953
rect 1638 1948 1644 1949
rect 1659 1953 1665 1954
rect 1659 1949 1660 1953
rect 1664 1949 1665 1953
rect 1659 1948 1665 1949
rect 1734 1953 1740 1954
rect 1734 1949 1735 1953
rect 1739 1949 1740 1953
rect 1734 1948 1740 1949
rect 1755 1953 1761 1954
rect 1755 1949 1756 1953
rect 1760 1949 1761 1953
rect 1755 1948 1761 1949
rect 1838 1953 1844 1954
rect 1838 1949 1839 1953
rect 1843 1949 1844 1953
rect 1942 1953 1948 1954
rect 1838 1948 1844 1949
rect 1846 1951 1852 1952
rect 1326 1947 1332 1948
rect 1846 1947 1847 1951
rect 1851 1950 1852 1951
rect 1859 1951 1865 1952
rect 1859 1950 1860 1951
rect 1851 1948 1860 1950
rect 1851 1947 1852 1948
rect 1846 1946 1852 1947
rect 1859 1947 1860 1948
rect 1864 1947 1865 1951
rect 1942 1949 1943 1953
rect 1947 1949 1948 1953
rect 1942 1948 1948 1949
rect 1963 1953 1969 1954
rect 1963 1949 1964 1953
rect 1968 1949 1969 1953
rect 1963 1948 1969 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2046 1948 2052 1949
rect 2067 1953 2073 1954
rect 2067 1949 2068 1953
rect 2072 1949 2073 1953
rect 2067 1948 2073 1949
rect 2150 1953 2156 1954
rect 2150 1949 2151 1953
rect 2155 1949 2156 1953
rect 2254 1953 2260 1954
rect 2150 1948 2156 1949
rect 2171 1951 2180 1952
rect 1859 1946 1865 1947
rect 2171 1947 2172 1951
rect 2179 1947 2180 1951
rect 2254 1949 2255 1953
rect 2259 1949 2260 1953
rect 2254 1948 2260 1949
rect 2275 1953 2281 1954
rect 2275 1949 2276 1953
rect 2280 1949 2281 1953
rect 2275 1948 2281 1949
rect 2366 1953 2372 1954
rect 2366 1949 2367 1953
rect 2371 1949 2372 1953
rect 2366 1948 2372 1949
rect 2387 1953 2393 1954
rect 2387 1949 2388 1953
rect 2392 1949 2393 1953
rect 2387 1948 2393 1949
rect 2454 1953 2460 1954
rect 2454 1949 2455 1953
rect 2459 1949 2460 1953
rect 2502 1952 2508 1953
rect 2454 1948 2460 1949
rect 2462 1951 2468 1952
rect 2171 1946 2180 1947
rect 2462 1947 2463 1951
rect 2467 1950 2468 1951
rect 2475 1951 2481 1952
rect 2475 1950 2476 1951
rect 2467 1948 2476 1950
rect 2467 1947 2468 1948
rect 2462 1946 2468 1947
rect 2475 1947 2476 1948
rect 2480 1947 2481 1951
rect 2502 1948 2503 1952
rect 2507 1948 2508 1952
rect 2502 1947 2508 1948
rect 2475 1946 2481 1947
rect 208 1945 233 1946
rect 208 1944 228 1945
rect 155 1943 161 1944
rect 155 1939 156 1943
rect 160 1939 161 1943
rect 227 1941 228 1944
rect 232 1941 233 1945
rect 245 1945 313 1946
rect 245 1944 308 1945
rect 227 1940 233 1941
rect 307 1941 308 1944
rect 312 1941 313 1945
rect 496 1945 513 1946
rect 496 1944 508 1945
rect 307 1940 313 1941
rect 403 1943 412 1944
rect 155 1938 161 1939
rect 403 1939 404 1943
rect 411 1939 412 1943
rect 507 1941 508 1944
rect 512 1941 513 1945
rect 600 1945 617 1946
rect 600 1944 612 1945
rect 507 1940 513 1941
rect 611 1941 612 1944
rect 616 1941 617 1945
rect 611 1940 617 1941
rect 715 1945 721 1946
rect 715 1941 716 1945
rect 720 1941 721 1945
rect 1024 1945 1041 1946
rect 1024 1944 1036 1945
rect 715 1940 721 1941
rect 819 1943 825 1944
rect 403 1938 412 1939
rect 819 1939 820 1943
rect 824 1942 825 1943
rect 886 1943 892 1944
rect 824 1940 882 1942
rect 824 1939 825 1940
rect 819 1938 825 1939
rect 157 1934 159 1938
rect 614 1935 620 1936
rect 614 1934 615 1935
rect 157 1932 615 1934
rect 614 1931 615 1932
rect 619 1931 620 1935
rect 880 1934 882 1940
rect 886 1939 887 1943
rect 891 1942 892 1943
rect 923 1943 929 1944
rect 923 1942 924 1943
rect 891 1940 924 1942
rect 891 1939 892 1940
rect 886 1938 892 1939
rect 923 1939 924 1940
rect 928 1939 929 1943
rect 1035 1941 1036 1944
rect 1040 1941 1041 1945
rect 1035 1940 1041 1941
rect 923 1938 929 1939
rect 1038 1935 1044 1936
rect 1038 1934 1039 1935
rect 880 1932 1039 1934
rect 614 1930 620 1931
rect 1038 1931 1039 1932
rect 1043 1931 1044 1935
rect 1038 1930 1044 1931
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 2502 1935 2508 1936
rect 1326 1930 1332 1931
rect 1438 1932 1444 1933
rect 1438 1928 1439 1932
rect 1443 1928 1444 1932
rect 1438 1927 1444 1928
rect 1526 1932 1532 1933
rect 1526 1928 1527 1932
rect 1531 1928 1532 1932
rect 1526 1927 1532 1928
rect 1622 1932 1628 1933
rect 1622 1928 1623 1932
rect 1627 1928 1628 1932
rect 1622 1927 1628 1928
rect 1718 1932 1724 1933
rect 1718 1928 1719 1932
rect 1723 1928 1724 1932
rect 1718 1927 1724 1928
rect 1822 1932 1828 1933
rect 1822 1928 1823 1932
rect 1827 1928 1828 1932
rect 1822 1927 1828 1928
rect 1926 1932 1932 1933
rect 1926 1928 1927 1932
rect 1931 1928 1932 1932
rect 1926 1927 1932 1928
rect 2030 1932 2036 1933
rect 2030 1928 2031 1932
rect 2035 1928 2036 1932
rect 2030 1927 2036 1928
rect 2134 1932 2140 1933
rect 2134 1928 2135 1932
rect 2139 1928 2140 1932
rect 2134 1927 2140 1928
rect 2238 1932 2244 1933
rect 2238 1928 2239 1932
rect 2243 1928 2244 1932
rect 2238 1927 2244 1928
rect 2350 1932 2356 1933
rect 2350 1928 2351 1932
rect 2355 1928 2356 1932
rect 2350 1927 2356 1928
rect 2438 1932 2444 1933
rect 2438 1928 2439 1932
rect 2443 1928 2444 1932
rect 2502 1931 2503 1935
rect 2507 1931 2508 1935
rect 2502 1930 2508 1931
rect 2438 1927 2444 1928
rect 702 1923 708 1924
rect 702 1922 703 1923
rect 319 1920 703 1922
rect 319 1918 321 1920
rect 702 1919 703 1920
rect 707 1919 708 1923
rect 702 1918 708 1919
rect 243 1917 321 1918
rect 155 1915 161 1916
rect 155 1911 156 1915
rect 160 1911 161 1915
rect 243 1913 244 1917
rect 248 1916 321 1917
rect 1526 1916 1532 1917
rect 248 1913 249 1916
rect 243 1912 249 1913
rect 366 1915 372 1916
rect 155 1910 161 1911
rect 366 1911 367 1915
rect 371 1914 372 1915
rect 379 1915 385 1916
rect 379 1914 380 1915
rect 371 1912 380 1914
rect 371 1911 372 1912
rect 366 1910 372 1911
rect 379 1911 380 1912
rect 384 1911 385 1915
rect 379 1910 385 1911
rect 531 1915 537 1916
rect 531 1911 532 1915
rect 536 1911 537 1915
rect 691 1915 697 1916
rect 691 1914 692 1915
rect 531 1910 537 1911
rect 552 1912 692 1914
rect 157 1906 159 1910
rect 533 1906 535 1910
rect 552 1906 554 1912
rect 691 1911 692 1912
rect 696 1911 697 1915
rect 691 1910 697 1911
rect 867 1915 873 1916
rect 867 1911 868 1915
rect 872 1911 873 1915
rect 867 1910 873 1911
rect 1043 1915 1049 1916
rect 1043 1911 1044 1915
rect 1048 1914 1049 1915
rect 1074 1915 1080 1916
rect 1074 1914 1075 1915
rect 1048 1912 1075 1914
rect 1048 1911 1049 1912
rect 1043 1910 1049 1911
rect 1074 1911 1075 1912
rect 1079 1911 1080 1915
rect 1074 1910 1080 1911
rect 1326 1913 1332 1914
rect 157 1904 263 1906
rect 261 1902 263 1904
rect 396 1904 535 1906
rect 548 1904 554 1906
rect 869 1906 871 1910
rect 1326 1909 1327 1913
rect 1331 1909 1332 1913
rect 1526 1912 1527 1916
rect 1531 1912 1532 1916
rect 1526 1911 1532 1912
rect 1614 1916 1620 1917
rect 1614 1912 1615 1916
rect 1619 1912 1620 1916
rect 1614 1911 1620 1912
rect 1710 1916 1716 1917
rect 1710 1912 1711 1916
rect 1715 1912 1716 1916
rect 1710 1911 1716 1912
rect 1814 1916 1820 1917
rect 1814 1912 1815 1916
rect 1819 1912 1820 1916
rect 1814 1911 1820 1912
rect 1918 1916 1924 1917
rect 1918 1912 1919 1916
rect 1923 1912 1924 1916
rect 1918 1911 1924 1912
rect 2014 1916 2020 1917
rect 2014 1912 2015 1916
rect 2019 1912 2020 1916
rect 2014 1911 2020 1912
rect 2110 1916 2116 1917
rect 2110 1912 2111 1916
rect 2115 1912 2116 1916
rect 2110 1911 2116 1912
rect 2198 1916 2204 1917
rect 2198 1912 2199 1916
rect 2203 1912 2204 1916
rect 2198 1911 2204 1912
rect 2286 1916 2292 1917
rect 2286 1912 2287 1916
rect 2291 1912 2292 1916
rect 2286 1911 2292 1912
rect 2374 1916 2380 1917
rect 2374 1912 2375 1916
rect 2379 1912 2380 1916
rect 2374 1911 2380 1912
rect 2438 1916 2444 1917
rect 2438 1912 2439 1916
rect 2443 1912 2444 1916
rect 2438 1911 2444 1912
rect 2502 1913 2508 1914
rect 1326 1908 1332 1909
rect 2502 1909 2503 1913
rect 2507 1909 2508 1913
rect 2502 1908 2508 1909
rect 869 1904 1062 1906
rect 396 1902 398 1904
rect 548 1902 550 1904
rect 1060 1902 1062 1904
rect 150 1901 156 1902
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 150 1897 151 1901
rect 155 1897 156 1901
rect 238 1901 244 1902
rect 150 1896 156 1897
rect 171 1899 177 1900
rect 110 1895 116 1896
rect 171 1895 172 1899
rect 176 1898 177 1899
rect 198 1899 204 1900
rect 198 1898 199 1899
rect 176 1896 199 1898
rect 176 1895 177 1896
rect 171 1894 177 1895
rect 198 1895 199 1896
rect 203 1895 204 1899
rect 238 1897 239 1901
rect 243 1897 244 1901
rect 238 1896 244 1897
rect 259 1901 265 1902
rect 259 1897 260 1901
rect 264 1897 265 1901
rect 259 1896 265 1897
rect 374 1901 380 1902
rect 374 1897 375 1901
rect 379 1897 380 1901
rect 374 1896 380 1897
rect 395 1901 401 1902
rect 395 1897 396 1901
rect 400 1897 401 1901
rect 395 1896 401 1897
rect 526 1901 532 1902
rect 526 1897 527 1901
rect 531 1897 532 1901
rect 526 1896 532 1897
rect 547 1901 553 1902
rect 547 1897 548 1901
rect 552 1897 553 1901
rect 547 1896 553 1897
rect 686 1901 692 1902
rect 686 1897 687 1901
rect 691 1897 692 1901
rect 862 1901 868 1902
rect 686 1896 692 1897
rect 702 1899 713 1900
rect 198 1894 204 1895
rect 702 1895 703 1899
rect 707 1895 708 1899
rect 712 1895 713 1899
rect 862 1897 863 1901
rect 867 1897 868 1901
rect 1038 1901 1044 1902
rect 862 1896 868 1897
rect 883 1899 892 1900
rect 702 1894 713 1895
rect 883 1895 884 1899
rect 891 1895 892 1899
rect 1038 1897 1039 1901
rect 1043 1897 1044 1901
rect 1038 1896 1044 1897
rect 1059 1901 1065 1902
rect 1059 1897 1060 1901
rect 1064 1897 1065 1901
rect 1059 1896 1065 1897
rect 1286 1900 1292 1901
rect 1286 1896 1287 1900
rect 1291 1896 1292 1900
rect 1286 1895 1292 1896
rect 1326 1896 1332 1897
rect 2502 1896 2508 1897
rect 883 1894 892 1895
rect 1326 1892 1327 1896
rect 1331 1892 1332 1896
rect 1326 1891 1332 1892
rect 1542 1895 1548 1896
rect 1542 1891 1543 1895
rect 1547 1891 1548 1895
rect 1542 1890 1548 1891
rect 1563 1895 1569 1896
rect 1563 1891 1564 1895
rect 1568 1891 1569 1895
rect 1563 1890 1569 1891
rect 1630 1895 1636 1896
rect 1630 1891 1631 1895
rect 1635 1891 1636 1895
rect 1630 1890 1636 1891
rect 1651 1895 1657 1896
rect 1651 1891 1652 1895
rect 1656 1891 1657 1895
rect 1651 1890 1657 1891
rect 1726 1895 1732 1896
rect 1726 1891 1727 1895
rect 1731 1891 1732 1895
rect 1726 1890 1732 1891
rect 1747 1895 1753 1896
rect 1747 1891 1748 1895
rect 1752 1894 1753 1895
rect 1830 1895 1836 1896
rect 1752 1892 1822 1894
rect 1752 1891 1753 1892
rect 1747 1890 1753 1891
rect 110 1883 116 1884
rect 110 1879 111 1883
rect 115 1879 116 1883
rect 1286 1883 1292 1884
rect 110 1878 116 1879
rect 134 1880 140 1881
rect 134 1876 135 1880
rect 139 1876 140 1880
rect 134 1875 140 1876
rect 222 1880 228 1881
rect 222 1876 223 1880
rect 227 1876 228 1880
rect 222 1875 228 1876
rect 358 1880 364 1881
rect 358 1876 359 1880
rect 363 1876 364 1880
rect 358 1875 364 1876
rect 510 1880 516 1881
rect 510 1876 511 1880
rect 515 1876 516 1880
rect 510 1875 516 1876
rect 670 1880 676 1881
rect 670 1876 671 1880
rect 675 1876 676 1880
rect 670 1875 676 1876
rect 846 1880 852 1881
rect 846 1876 847 1880
rect 851 1876 852 1880
rect 846 1875 852 1876
rect 1022 1880 1028 1881
rect 1022 1876 1023 1880
rect 1027 1876 1028 1880
rect 1286 1879 1287 1883
rect 1291 1879 1292 1883
rect 1565 1882 1567 1890
rect 1653 1882 1655 1890
rect 1820 1882 1822 1892
rect 1830 1891 1831 1895
rect 1835 1891 1836 1895
rect 1830 1890 1836 1891
rect 1851 1895 1857 1896
rect 1851 1891 1852 1895
rect 1856 1894 1857 1895
rect 1934 1895 1940 1896
rect 1856 1892 1930 1894
rect 1856 1891 1857 1892
rect 1851 1890 1857 1891
rect 1928 1882 1930 1892
rect 1934 1891 1935 1895
rect 1939 1891 1940 1895
rect 1934 1890 1940 1891
rect 1955 1895 1961 1896
rect 1955 1891 1956 1895
rect 1960 1894 1961 1895
rect 1974 1895 1980 1896
rect 1974 1894 1975 1895
rect 1960 1892 1975 1894
rect 1960 1891 1961 1892
rect 1955 1890 1961 1891
rect 1974 1891 1975 1892
rect 1979 1891 1980 1895
rect 1974 1890 1980 1891
rect 2030 1895 2036 1896
rect 2030 1891 2031 1895
rect 2035 1891 2036 1895
rect 2030 1890 2036 1891
rect 2051 1895 2057 1896
rect 2051 1891 2052 1895
rect 2056 1894 2057 1895
rect 2126 1895 2132 1896
rect 2056 1892 2122 1894
rect 2056 1891 2057 1892
rect 2051 1890 2057 1891
rect 2120 1882 2122 1892
rect 2126 1891 2127 1895
rect 2131 1891 2132 1895
rect 2126 1890 2132 1891
rect 2147 1895 2153 1896
rect 2147 1891 2148 1895
rect 2152 1894 2153 1895
rect 2214 1895 2220 1896
rect 2152 1892 2206 1894
rect 2152 1891 2153 1892
rect 2147 1890 2153 1891
rect 2204 1882 2206 1892
rect 2214 1891 2215 1895
rect 2219 1891 2220 1895
rect 2214 1890 2220 1891
rect 2235 1895 2241 1896
rect 2235 1891 2236 1895
rect 2240 1894 2241 1895
rect 2246 1895 2252 1896
rect 2246 1894 2247 1895
rect 2240 1892 2247 1894
rect 2240 1891 2241 1892
rect 2235 1890 2241 1891
rect 2246 1891 2247 1892
rect 2251 1891 2252 1895
rect 2246 1890 2252 1891
rect 2302 1895 2308 1896
rect 2302 1891 2303 1895
rect 2307 1891 2308 1895
rect 2302 1890 2308 1891
rect 2318 1895 2329 1896
rect 2318 1891 2319 1895
rect 2323 1891 2324 1895
rect 2328 1891 2329 1895
rect 2318 1890 2329 1891
rect 2390 1895 2396 1896
rect 2390 1891 2391 1895
rect 2395 1891 2396 1895
rect 2411 1895 2417 1896
rect 2411 1894 2412 1895
rect 2390 1890 2396 1891
rect 2400 1892 2412 1894
rect 2400 1886 2402 1892
rect 2411 1891 2412 1892
rect 2416 1891 2417 1895
rect 2411 1890 2417 1891
rect 2454 1895 2460 1896
rect 2454 1891 2455 1895
rect 2459 1891 2460 1895
rect 2454 1890 2460 1891
rect 2475 1895 2481 1896
rect 2475 1891 2476 1895
rect 2480 1894 2481 1895
rect 2486 1895 2492 1896
rect 2486 1894 2487 1895
rect 2480 1892 2487 1894
rect 2480 1891 2481 1892
rect 2475 1890 2481 1891
rect 2486 1891 2487 1892
rect 2491 1891 2492 1895
rect 2502 1892 2503 1896
rect 2507 1892 2508 1896
rect 2502 1891 2508 1892
rect 2486 1890 2492 1891
rect 2308 1884 2402 1886
rect 2308 1882 2310 1884
rect 1565 1881 1641 1882
rect 1565 1880 1636 1881
rect 1286 1878 1292 1879
rect 1547 1879 1553 1880
rect 1022 1875 1028 1876
rect 1547 1875 1548 1879
rect 1552 1878 1553 1879
rect 1552 1876 1630 1878
rect 1635 1877 1636 1880
rect 1640 1877 1641 1881
rect 1653 1881 1737 1882
rect 1653 1880 1732 1881
rect 1635 1876 1641 1877
rect 1731 1877 1732 1880
rect 1736 1877 1737 1881
rect 1820 1881 1841 1882
rect 1820 1880 1836 1881
rect 1731 1876 1737 1877
rect 1835 1877 1836 1880
rect 1840 1877 1841 1881
rect 1928 1881 1945 1882
rect 1928 1880 1940 1881
rect 1835 1876 1841 1877
rect 1939 1877 1940 1880
rect 1944 1877 1945 1881
rect 2120 1881 2137 1882
rect 2120 1880 2132 1881
rect 1939 1876 1945 1877
rect 2035 1879 2041 1880
rect 1552 1875 1553 1876
rect 1547 1874 1553 1875
rect 1628 1874 1630 1876
rect 1846 1875 1852 1876
rect 1846 1874 1847 1875
rect 1628 1872 1847 1874
rect 1846 1871 1847 1872
rect 1851 1871 1852 1875
rect 2035 1875 2036 1879
rect 2040 1878 2041 1879
rect 2040 1876 2126 1878
rect 2131 1877 2132 1880
rect 2136 1877 2137 1881
rect 2204 1881 2225 1882
rect 2204 1880 2220 1881
rect 2131 1876 2137 1877
rect 2219 1877 2220 1880
rect 2224 1877 2225 1881
rect 2219 1876 2225 1877
rect 2307 1881 2313 1882
rect 2307 1877 2308 1881
rect 2312 1877 2313 1881
rect 2307 1876 2313 1877
rect 2395 1879 2401 1880
rect 2040 1875 2041 1876
rect 2035 1874 2041 1875
rect 2124 1874 2126 1876
rect 2318 1875 2324 1876
rect 2318 1874 2319 1875
rect 2124 1872 2319 1874
rect 1846 1870 1852 1871
rect 2318 1871 2319 1872
rect 2323 1871 2324 1875
rect 2395 1875 2396 1879
rect 2400 1878 2401 1879
rect 2459 1879 2468 1880
rect 2400 1876 2454 1878
rect 2400 1875 2401 1876
rect 2395 1874 2401 1875
rect 2318 1870 2324 1871
rect 2452 1870 2454 1876
rect 2459 1875 2460 1879
rect 2467 1875 2468 1879
rect 2459 1874 2468 1875
rect 2474 1871 2480 1872
rect 2474 1870 2475 1871
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 190 1868 196 1869
rect 190 1864 191 1868
rect 195 1864 196 1868
rect 190 1863 196 1864
rect 262 1868 268 1869
rect 262 1864 263 1868
rect 267 1864 268 1868
rect 262 1863 268 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 406 1868 412 1869
rect 406 1864 407 1868
rect 411 1864 412 1868
rect 406 1863 412 1864
rect 478 1868 484 1869
rect 478 1864 479 1868
rect 483 1864 484 1868
rect 478 1863 484 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 614 1868 620 1869
rect 614 1864 615 1868
rect 619 1864 620 1868
rect 614 1863 620 1864
rect 678 1868 684 1869
rect 678 1864 679 1868
rect 683 1864 684 1868
rect 678 1863 684 1864
rect 742 1868 748 1869
rect 742 1864 743 1868
rect 747 1864 748 1868
rect 742 1863 748 1864
rect 814 1868 820 1869
rect 814 1864 815 1868
rect 819 1864 820 1868
rect 814 1863 820 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 958 1868 964 1869
rect 958 1864 959 1868
rect 963 1864 964 1868
rect 958 1863 964 1864
rect 1038 1868 1044 1869
rect 2452 1868 2475 1870
rect 1038 1864 1039 1868
rect 1043 1864 1044 1868
rect 1802 1867 1808 1868
rect 1802 1866 1803 1867
rect 1038 1863 1044 1864
rect 1286 1865 1292 1866
rect 110 1860 116 1861
rect 1286 1861 1287 1865
rect 1291 1861 1292 1865
rect 1540 1864 1803 1866
rect 1540 1862 1542 1864
rect 1802 1863 1803 1864
rect 1807 1863 1808 1867
rect 2474 1867 2475 1868
rect 2479 1867 2480 1871
rect 2474 1866 2480 1867
rect 1802 1862 1808 1863
rect 1286 1860 1292 1861
rect 1539 1861 1545 1862
rect 1539 1857 1540 1861
rect 1544 1857 1545 1861
rect 1611 1859 1617 1860
rect 1611 1858 1612 1859
rect 1539 1856 1545 1857
rect 1557 1856 1612 1858
rect 110 1848 116 1849
rect 1286 1848 1292 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 150 1847 156 1848
rect 150 1843 151 1847
rect 155 1843 156 1847
rect 150 1842 156 1843
rect 158 1847 164 1848
rect 158 1843 159 1847
rect 163 1846 164 1847
rect 171 1847 177 1848
rect 171 1846 172 1847
rect 163 1844 172 1846
rect 163 1843 164 1844
rect 158 1842 164 1843
rect 171 1843 172 1844
rect 176 1843 177 1847
rect 171 1842 177 1843
rect 206 1847 212 1848
rect 206 1843 207 1847
rect 211 1843 212 1847
rect 206 1842 212 1843
rect 227 1847 233 1848
rect 227 1843 228 1847
rect 232 1843 233 1847
rect 227 1842 233 1843
rect 278 1847 284 1848
rect 278 1843 279 1847
rect 283 1843 284 1847
rect 278 1842 284 1843
rect 299 1847 305 1848
rect 299 1843 300 1847
rect 304 1846 305 1847
rect 350 1847 356 1848
rect 304 1844 321 1846
rect 304 1843 305 1844
rect 299 1842 305 1843
rect 229 1834 231 1842
rect 319 1834 321 1844
rect 350 1843 351 1847
rect 355 1843 356 1847
rect 350 1842 356 1843
rect 358 1847 364 1848
rect 358 1843 359 1847
rect 363 1846 364 1847
rect 371 1847 377 1848
rect 371 1846 372 1847
rect 363 1844 372 1846
rect 363 1843 364 1844
rect 358 1842 364 1843
rect 371 1843 372 1844
rect 376 1843 377 1847
rect 371 1842 377 1843
rect 422 1847 428 1848
rect 422 1843 423 1847
rect 427 1843 428 1847
rect 422 1842 428 1843
rect 443 1847 449 1848
rect 443 1843 444 1847
rect 448 1846 449 1847
rect 494 1847 500 1848
rect 448 1844 490 1846
rect 448 1843 449 1844
rect 443 1842 449 1843
rect 488 1834 490 1844
rect 494 1843 495 1847
rect 499 1843 500 1847
rect 494 1842 500 1843
rect 515 1847 521 1848
rect 515 1843 516 1847
rect 520 1843 521 1847
rect 515 1842 521 1843
rect 566 1847 572 1848
rect 566 1843 567 1847
rect 571 1843 572 1847
rect 566 1842 572 1843
rect 587 1847 593 1848
rect 587 1843 588 1847
rect 592 1846 593 1847
rect 630 1847 636 1848
rect 592 1844 622 1846
rect 592 1843 593 1844
rect 587 1842 593 1843
rect 517 1834 519 1842
rect 620 1834 622 1844
rect 630 1843 631 1847
rect 635 1843 636 1847
rect 630 1842 636 1843
rect 651 1847 657 1848
rect 651 1843 652 1847
rect 656 1846 657 1847
rect 694 1847 700 1848
rect 656 1844 686 1846
rect 656 1843 657 1844
rect 651 1842 657 1843
rect 684 1834 686 1844
rect 694 1843 695 1847
rect 699 1843 700 1847
rect 694 1842 700 1843
rect 715 1847 721 1848
rect 715 1843 716 1847
rect 720 1843 721 1847
rect 715 1842 721 1843
rect 758 1847 764 1848
rect 758 1843 759 1847
rect 763 1843 764 1847
rect 758 1842 764 1843
rect 779 1847 785 1848
rect 779 1843 780 1847
rect 784 1846 785 1847
rect 830 1847 836 1848
rect 784 1844 826 1846
rect 784 1843 785 1844
rect 779 1842 785 1843
rect 717 1834 719 1842
rect 824 1838 826 1844
rect 830 1843 831 1847
rect 835 1843 836 1847
rect 830 1842 836 1843
rect 851 1847 857 1848
rect 851 1843 852 1847
rect 856 1846 857 1847
rect 902 1847 908 1848
rect 856 1844 898 1846
rect 856 1843 857 1844
rect 851 1842 857 1843
rect 824 1836 839 1838
rect 837 1834 839 1836
rect 896 1834 898 1844
rect 902 1843 903 1847
rect 907 1843 908 1847
rect 902 1842 908 1843
rect 923 1847 929 1848
rect 923 1843 924 1847
rect 928 1843 929 1847
rect 923 1842 929 1843
rect 974 1847 980 1848
rect 974 1843 975 1847
rect 979 1843 980 1847
rect 974 1842 980 1843
rect 982 1847 988 1848
rect 982 1843 983 1847
rect 987 1846 988 1847
rect 995 1847 1001 1848
rect 995 1846 996 1847
rect 987 1844 996 1846
rect 987 1843 988 1844
rect 982 1842 988 1843
rect 995 1843 996 1844
rect 1000 1843 1001 1847
rect 995 1842 1001 1843
rect 1054 1847 1060 1848
rect 1054 1843 1055 1847
rect 1059 1843 1060 1847
rect 1054 1842 1060 1843
rect 1074 1847 1081 1848
rect 1074 1843 1075 1847
rect 1080 1843 1081 1847
rect 1286 1844 1287 1848
rect 1291 1844 1292 1848
rect 1557 1846 1559 1856
rect 1611 1855 1612 1856
rect 1616 1855 1617 1859
rect 1691 1859 1697 1860
rect 1691 1858 1692 1859
rect 1611 1854 1617 1855
rect 1661 1856 1692 1858
rect 1661 1850 1663 1856
rect 1691 1855 1692 1856
rect 1696 1855 1697 1859
rect 1691 1854 1697 1855
rect 1787 1859 1793 1860
rect 1787 1855 1788 1859
rect 1792 1858 1793 1859
rect 1883 1859 1889 1860
rect 1792 1856 1874 1858
rect 1792 1855 1793 1856
rect 1787 1854 1793 1855
rect 1628 1848 1663 1850
rect 1872 1850 1874 1856
rect 1883 1855 1884 1859
rect 1888 1858 1889 1859
rect 1974 1859 1980 1860
rect 1888 1856 1946 1858
rect 1888 1855 1889 1856
rect 1883 1854 1889 1855
rect 1944 1850 1946 1856
rect 1974 1855 1975 1859
rect 1979 1858 1980 1859
rect 1987 1859 1993 1860
rect 1987 1858 1988 1859
rect 1979 1856 1988 1858
rect 1979 1855 1980 1856
rect 1974 1854 1980 1855
rect 1987 1855 1988 1856
rect 1992 1855 1993 1859
rect 1987 1854 1993 1855
rect 2083 1859 2089 1860
rect 2083 1855 2084 1859
rect 2088 1858 2089 1859
rect 2166 1859 2172 1860
rect 2166 1858 2167 1859
rect 2088 1856 2167 1858
rect 2088 1855 2089 1856
rect 2083 1854 2089 1855
rect 2166 1855 2167 1856
rect 2171 1855 2172 1859
rect 2166 1854 2172 1855
rect 2179 1859 2185 1860
rect 2179 1855 2180 1859
rect 2184 1855 2185 1859
rect 2179 1854 2185 1855
rect 2275 1859 2281 1860
rect 2275 1855 2276 1859
rect 2280 1855 2281 1859
rect 2371 1859 2377 1860
rect 2371 1858 2372 1859
rect 2275 1854 2281 1855
rect 2296 1856 2372 1858
rect 2181 1850 2183 1854
rect 2277 1850 2279 1854
rect 2296 1850 2298 1856
rect 2371 1855 2372 1856
rect 2376 1855 2377 1859
rect 2371 1854 2377 1855
rect 2459 1859 2465 1860
rect 2459 1855 2460 1859
rect 2464 1855 2465 1859
rect 2459 1854 2465 1855
rect 2461 1850 2463 1854
rect 1872 1848 1902 1850
rect 1944 1848 2007 1850
rect 1628 1846 1630 1848
rect 1900 1846 1902 1848
rect 2005 1846 2007 1848
rect 2100 1848 2183 1850
rect 2196 1848 2279 1850
rect 2292 1848 2298 1850
rect 2389 1848 2463 1850
rect 2100 1846 2102 1848
rect 2196 1846 2198 1848
rect 2292 1846 2294 1848
rect 2389 1846 2391 1848
rect 1534 1845 1540 1846
rect 1286 1843 1292 1844
rect 1326 1844 1332 1845
rect 1074 1842 1081 1843
rect 925 1834 927 1842
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1534 1841 1535 1845
rect 1539 1841 1540 1845
rect 1534 1840 1540 1841
rect 1555 1845 1561 1846
rect 1555 1841 1556 1845
rect 1560 1841 1561 1845
rect 1555 1840 1561 1841
rect 1606 1845 1612 1846
rect 1606 1841 1607 1845
rect 1611 1841 1612 1845
rect 1606 1840 1612 1841
rect 1627 1845 1633 1846
rect 1627 1841 1628 1845
rect 1632 1841 1633 1845
rect 1627 1840 1633 1841
rect 1686 1845 1692 1846
rect 1686 1841 1687 1845
rect 1691 1841 1692 1845
rect 1782 1845 1788 1846
rect 1686 1840 1692 1841
rect 1694 1843 1700 1844
rect 1326 1839 1332 1840
rect 1694 1839 1695 1843
rect 1699 1842 1700 1843
rect 1707 1843 1713 1844
rect 1707 1842 1708 1843
rect 1699 1840 1708 1842
rect 1699 1839 1700 1840
rect 1694 1838 1700 1839
rect 1707 1839 1708 1840
rect 1712 1839 1713 1843
rect 1782 1841 1783 1845
rect 1787 1841 1788 1845
rect 1878 1845 1884 1846
rect 1782 1840 1788 1841
rect 1802 1843 1809 1844
rect 1707 1838 1713 1839
rect 1802 1839 1803 1843
rect 1808 1839 1809 1843
rect 1878 1841 1879 1845
rect 1883 1841 1884 1845
rect 1878 1840 1884 1841
rect 1899 1845 1905 1846
rect 1899 1841 1900 1845
rect 1904 1841 1905 1845
rect 1899 1840 1905 1841
rect 1982 1845 1988 1846
rect 1982 1841 1983 1845
rect 1987 1841 1988 1845
rect 1982 1840 1988 1841
rect 2003 1845 2009 1846
rect 2003 1841 2004 1845
rect 2008 1841 2009 1845
rect 2003 1840 2009 1841
rect 2078 1845 2084 1846
rect 2078 1841 2079 1845
rect 2083 1841 2084 1845
rect 2078 1840 2084 1841
rect 2099 1845 2105 1846
rect 2099 1841 2100 1845
rect 2104 1841 2105 1845
rect 2099 1840 2105 1841
rect 2174 1845 2180 1846
rect 2174 1841 2175 1845
rect 2179 1841 2180 1845
rect 2174 1840 2180 1841
rect 2195 1845 2201 1846
rect 2195 1841 2196 1845
rect 2200 1841 2201 1845
rect 2195 1840 2201 1841
rect 2270 1845 2276 1846
rect 2270 1841 2271 1845
rect 2275 1841 2276 1845
rect 2270 1840 2276 1841
rect 2291 1845 2297 1846
rect 2291 1841 2292 1845
rect 2296 1841 2297 1845
rect 2291 1840 2297 1841
rect 2366 1845 2372 1846
rect 2366 1841 2367 1845
rect 2371 1841 2372 1845
rect 2366 1840 2372 1841
rect 2387 1845 2393 1846
rect 2387 1841 2388 1845
rect 2392 1841 2393 1845
rect 2387 1840 2393 1841
rect 2454 1845 2460 1846
rect 2454 1841 2455 1845
rect 2459 1841 2460 1845
rect 2502 1844 2508 1845
rect 2454 1840 2460 1841
rect 2474 1843 2481 1844
rect 1802 1838 1809 1839
rect 2474 1839 2475 1843
rect 2480 1839 2481 1843
rect 2502 1840 2503 1844
rect 2507 1840 2508 1844
rect 2502 1839 2508 1840
rect 2474 1838 2481 1839
rect 229 1833 289 1834
rect 229 1832 284 1833
rect 155 1831 161 1832
rect 155 1827 156 1831
rect 160 1827 161 1831
rect 155 1826 161 1827
rect 198 1831 204 1832
rect 198 1827 199 1831
rect 203 1830 204 1831
rect 211 1831 217 1832
rect 211 1830 212 1831
rect 203 1828 212 1830
rect 203 1827 204 1828
rect 198 1826 204 1827
rect 211 1827 212 1828
rect 216 1827 217 1831
rect 283 1829 284 1832
rect 288 1829 289 1833
rect 319 1833 361 1834
rect 319 1832 356 1833
rect 283 1828 289 1829
rect 355 1829 356 1832
rect 360 1829 361 1833
rect 488 1833 505 1834
rect 488 1832 500 1833
rect 355 1828 361 1829
rect 427 1831 433 1832
rect 211 1826 217 1827
rect 427 1827 428 1831
rect 432 1830 433 1831
rect 458 1831 464 1832
rect 458 1830 459 1831
rect 432 1828 459 1830
rect 432 1827 433 1828
rect 427 1826 433 1827
rect 458 1827 459 1828
rect 463 1827 464 1831
rect 499 1829 500 1832
rect 504 1829 505 1833
rect 517 1833 577 1834
rect 517 1832 572 1833
rect 499 1828 505 1829
rect 571 1829 572 1832
rect 576 1829 577 1833
rect 620 1833 641 1834
rect 620 1832 636 1833
rect 571 1828 577 1829
rect 635 1829 636 1832
rect 640 1829 641 1833
rect 684 1833 705 1834
rect 684 1832 700 1833
rect 635 1828 641 1829
rect 699 1829 700 1832
rect 704 1829 705 1833
rect 717 1833 769 1834
rect 717 1832 764 1833
rect 699 1828 705 1829
rect 763 1829 764 1832
rect 768 1829 769 1833
rect 763 1828 769 1829
rect 835 1833 841 1834
rect 835 1829 836 1833
rect 840 1829 841 1833
rect 896 1833 913 1834
rect 896 1832 908 1833
rect 835 1828 841 1829
rect 907 1829 908 1832
rect 912 1829 913 1833
rect 925 1833 985 1834
rect 925 1832 980 1833
rect 907 1828 913 1829
rect 979 1829 980 1832
rect 984 1829 985 1833
rect 979 1828 985 1829
rect 1059 1831 1068 1832
rect 458 1826 464 1827
rect 1059 1827 1060 1831
rect 1067 1827 1068 1831
rect 1059 1826 1068 1827
rect 1326 1827 1332 1828
rect 157 1822 159 1826
rect 358 1823 364 1824
rect 358 1822 359 1823
rect 157 1820 359 1822
rect 358 1819 359 1820
rect 363 1819 364 1823
rect 1326 1823 1327 1827
rect 1331 1823 1332 1827
rect 2502 1827 2508 1828
rect 1326 1822 1332 1823
rect 1518 1824 1524 1825
rect 1518 1820 1519 1824
rect 1523 1820 1524 1824
rect 1518 1819 1524 1820
rect 1590 1824 1596 1825
rect 1590 1820 1591 1824
rect 1595 1820 1596 1824
rect 1590 1819 1596 1820
rect 1670 1824 1676 1825
rect 1670 1820 1671 1824
rect 1675 1820 1676 1824
rect 1670 1819 1676 1820
rect 1766 1824 1772 1825
rect 1766 1820 1767 1824
rect 1771 1820 1772 1824
rect 1766 1819 1772 1820
rect 1862 1824 1868 1825
rect 1862 1820 1863 1824
rect 1867 1820 1868 1824
rect 1862 1819 1868 1820
rect 1966 1824 1972 1825
rect 1966 1820 1967 1824
rect 1971 1820 1972 1824
rect 1966 1819 1972 1820
rect 2062 1824 2068 1825
rect 2062 1820 2063 1824
rect 2067 1820 2068 1824
rect 2062 1819 2068 1820
rect 2158 1824 2164 1825
rect 2158 1820 2159 1824
rect 2163 1820 2164 1824
rect 2158 1819 2164 1820
rect 2254 1824 2260 1825
rect 2254 1820 2255 1824
rect 2259 1820 2260 1824
rect 2254 1819 2260 1820
rect 2350 1824 2356 1825
rect 2350 1820 2351 1824
rect 2355 1820 2356 1824
rect 2350 1819 2356 1820
rect 2438 1824 2444 1825
rect 2438 1820 2439 1824
rect 2443 1820 2444 1824
rect 2502 1823 2503 1827
rect 2507 1823 2508 1827
rect 2502 1822 2508 1823
rect 2438 1819 2444 1820
rect 358 1818 364 1819
rect 650 1811 656 1812
rect 650 1810 651 1811
rect 444 1808 651 1810
rect 444 1806 446 1808
rect 650 1807 651 1808
rect 655 1807 656 1811
rect 982 1811 988 1812
rect 982 1810 983 1811
rect 650 1806 656 1807
rect 724 1808 983 1810
rect 724 1806 726 1808
rect 982 1807 983 1808
rect 987 1807 988 1811
rect 982 1806 988 1807
rect 1462 1808 1468 1809
rect 443 1805 449 1806
rect 155 1803 164 1804
rect 155 1799 156 1803
rect 163 1799 164 1803
rect 235 1803 241 1804
rect 235 1802 236 1803
rect 155 1798 164 1799
rect 173 1800 236 1802
rect 173 1790 175 1800
rect 235 1799 236 1800
rect 240 1799 241 1803
rect 339 1803 345 1804
rect 339 1802 340 1803
rect 235 1798 241 1799
rect 319 1800 340 1802
rect 319 1790 321 1800
rect 339 1799 340 1800
rect 344 1799 345 1803
rect 443 1801 444 1805
rect 448 1801 449 1805
rect 723 1805 729 1806
rect 443 1800 449 1801
rect 498 1803 504 1804
rect 339 1798 345 1799
rect 498 1799 499 1803
rect 503 1802 504 1803
rect 539 1803 545 1804
rect 539 1802 540 1803
rect 503 1800 540 1802
rect 503 1799 504 1800
rect 498 1798 504 1799
rect 539 1799 540 1800
rect 544 1799 545 1803
rect 635 1803 641 1804
rect 635 1802 636 1803
rect 539 1798 545 1799
rect 556 1800 636 1802
rect 556 1790 558 1800
rect 635 1799 636 1800
rect 640 1799 641 1803
rect 723 1801 724 1805
rect 728 1801 729 1805
rect 1326 1805 1332 1806
rect 723 1800 729 1801
rect 803 1803 809 1804
rect 635 1798 641 1799
rect 803 1799 804 1803
rect 808 1799 809 1803
rect 803 1798 809 1799
rect 883 1803 889 1804
rect 883 1799 884 1803
rect 888 1799 889 1803
rect 883 1798 889 1799
rect 963 1803 969 1804
rect 963 1799 964 1803
rect 968 1799 969 1803
rect 963 1798 969 1799
rect 1043 1803 1049 1804
rect 1043 1799 1044 1803
rect 1048 1802 1049 1803
rect 1123 1803 1129 1804
rect 1048 1800 1118 1802
rect 1048 1799 1049 1800
rect 1043 1798 1049 1799
rect 805 1794 807 1798
rect 885 1794 887 1798
rect 965 1794 967 1798
rect 740 1792 807 1794
rect 821 1792 887 1794
rect 900 1792 967 1794
rect 1116 1794 1118 1800
rect 1123 1799 1124 1803
rect 1128 1802 1129 1803
rect 1138 1803 1144 1804
rect 1138 1802 1139 1803
rect 1128 1800 1139 1802
rect 1128 1799 1129 1800
rect 1123 1798 1129 1799
rect 1138 1799 1139 1800
rect 1143 1799 1144 1803
rect 1326 1801 1327 1805
rect 1331 1801 1332 1805
rect 1462 1804 1463 1808
rect 1467 1804 1468 1808
rect 1462 1803 1468 1804
rect 1558 1808 1564 1809
rect 1558 1804 1559 1808
rect 1563 1804 1564 1808
rect 1558 1803 1564 1804
rect 1662 1808 1668 1809
rect 1662 1804 1663 1808
rect 1667 1804 1668 1808
rect 1662 1803 1668 1804
rect 1766 1808 1772 1809
rect 1766 1804 1767 1808
rect 1771 1804 1772 1808
rect 1766 1803 1772 1804
rect 1878 1808 1884 1809
rect 1878 1804 1879 1808
rect 1883 1804 1884 1808
rect 1878 1803 1884 1804
rect 1982 1808 1988 1809
rect 1982 1804 1983 1808
rect 1987 1804 1988 1808
rect 1982 1803 1988 1804
rect 2086 1808 2092 1809
rect 2086 1804 2087 1808
rect 2091 1804 2092 1808
rect 2086 1803 2092 1804
rect 2182 1808 2188 1809
rect 2182 1804 2183 1808
rect 2187 1804 2188 1808
rect 2182 1803 2188 1804
rect 2270 1808 2276 1809
rect 2270 1804 2271 1808
rect 2275 1804 2276 1808
rect 2270 1803 2276 1804
rect 2366 1808 2372 1809
rect 2366 1804 2367 1808
rect 2371 1804 2372 1808
rect 2366 1803 2372 1804
rect 2438 1808 2444 1809
rect 2438 1804 2439 1808
rect 2443 1804 2444 1808
rect 2438 1803 2444 1804
rect 2502 1805 2508 1806
rect 1326 1800 1332 1801
rect 2502 1801 2503 1805
rect 2507 1801 2508 1805
rect 2502 1800 2508 1801
rect 1138 1798 1144 1799
rect 1116 1792 1143 1794
rect 740 1790 742 1792
rect 821 1790 823 1792
rect 900 1790 902 1792
rect 1141 1790 1143 1792
rect 150 1789 156 1790
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 150 1785 151 1789
rect 155 1785 156 1789
rect 150 1784 156 1785
rect 171 1789 177 1790
rect 171 1785 172 1789
rect 176 1785 177 1789
rect 171 1784 177 1785
rect 230 1789 236 1790
rect 230 1785 231 1789
rect 235 1785 236 1789
rect 230 1784 236 1785
rect 251 1789 321 1790
rect 251 1785 252 1789
rect 256 1788 321 1789
rect 334 1789 340 1790
rect 256 1785 257 1788
rect 251 1784 257 1785
rect 334 1785 335 1789
rect 339 1785 340 1789
rect 438 1789 444 1790
rect 334 1784 340 1785
rect 355 1787 364 1788
rect 110 1783 116 1784
rect 355 1783 356 1787
rect 363 1783 364 1787
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 534 1789 540 1790
rect 438 1784 444 1785
rect 458 1787 465 1788
rect 355 1782 364 1783
rect 458 1783 459 1787
rect 464 1783 465 1787
rect 534 1785 535 1789
rect 539 1785 540 1789
rect 534 1784 540 1785
rect 555 1789 561 1790
rect 555 1785 556 1789
rect 560 1785 561 1789
rect 555 1784 561 1785
rect 630 1789 636 1790
rect 630 1785 631 1789
rect 635 1785 636 1789
rect 718 1789 724 1790
rect 630 1784 636 1785
rect 650 1787 657 1788
rect 458 1782 465 1783
rect 650 1783 651 1787
rect 656 1783 657 1787
rect 718 1785 719 1789
rect 723 1785 724 1789
rect 718 1784 724 1785
rect 739 1789 745 1790
rect 739 1785 740 1789
rect 744 1785 745 1789
rect 739 1784 745 1785
rect 798 1789 804 1790
rect 798 1785 799 1789
rect 803 1785 804 1789
rect 798 1784 804 1785
rect 819 1789 825 1790
rect 819 1785 820 1789
rect 824 1785 825 1789
rect 819 1784 825 1785
rect 878 1789 884 1790
rect 878 1785 879 1789
rect 883 1785 884 1789
rect 878 1784 884 1785
rect 899 1789 905 1790
rect 899 1785 900 1789
rect 904 1785 905 1789
rect 899 1784 905 1785
rect 958 1789 964 1790
rect 958 1785 959 1789
rect 963 1785 964 1789
rect 1038 1789 1044 1790
rect 958 1784 964 1785
rect 979 1787 985 1788
rect 650 1782 657 1783
rect 979 1783 980 1787
rect 984 1786 985 1787
rect 998 1787 1004 1788
rect 998 1786 999 1787
rect 984 1784 999 1786
rect 984 1783 985 1784
rect 979 1782 985 1783
rect 998 1783 999 1784
rect 1003 1783 1004 1787
rect 1038 1785 1039 1789
rect 1043 1785 1044 1789
rect 1118 1789 1124 1790
rect 1038 1784 1044 1785
rect 1059 1787 1068 1788
rect 998 1782 1004 1783
rect 1059 1783 1060 1787
rect 1067 1783 1068 1787
rect 1118 1785 1119 1789
rect 1123 1785 1124 1789
rect 1118 1784 1124 1785
rect 1139 1789 1145 1790
rect 1139 1785 1140 1789
rect 1144 1785 1145 1789
rect 1139 1784 1145 1785
rect 1286 1788 1292 1789
rect 1286 1784 1287 1788
rect 1291 1784 1292 1788
rect 1286 1783 1292 1784
rect 1326 1788 1332 1789
rect 2502 1788 2508 1789
rect 1326 1784 1327 1788
rect 1331 1784 1332 1788
rect 1326 1783 1332 1784
rect 1478 1787 1484 1788
rect 1478 1783 1479 1787
rect 1483 1783 1484 1787
rect 1059 1782 1068 1783
rect 1478 1782 1484 1783
rect 1499 1787 1505 1788
rect 1499 1783 1500 1787
rect 1504 1786 1505 1787
rect 1558 1787 1564 1788
rect 1558 1786 1559 1787
rect 1504 1784 1559 1786
rect 1504 1783 1505 1784
rect 1499 1782 1505 1783
rect 1558 1783 1559 1784
rect 1563 1783 1564 1787
rect 1558 1782 1564 1783
rect 1574 1787 1580 1788
rect 1574 1783 1575 1787
rect 1579 1783 1580 1787
rect 1595 1787 1601 1788
rect 1595 1786 1596 1787
rect 1574 1782 1580 1783
rect 1584 1784 1596 1786
rect 1584 1778 1586 1784
rect 1595 1783 1596 1784
rect 1600 1783 1601 1787
rect 1595 1782 1601 1783
rect 1678 1787 1684 1788
rect 1678 1783 1679 1787
rect 1683 1783 1684 1787
rect 1678 1782 1684 1783
rect 1699 1787 1705 1788
rect 1699 1783 1700 1787
rect 1704 1786 1705 1787
rect 1782 1787 1788 1788
rect 1704 1784 1778 1786
rect 1704 1783 1705 1784
rect 1699 1782 1705 1783
rect 1484 1776 1586 1778
rect 1484 1774 1486 1776
rect 1776 1774 1778 1784
rect 1782 1783 1783 1787
rect 1787 1783 1788 1787
rect 1782 1782 1788 1783
rect 1803 1787 1809 1788
rect 1803 1783 1804 1787
rect 1808 1786 1809 1787
rect 1894 1787 1900 1788
rect 1808 1784 1890 1786
rect 1808 1783 1809 1784
rect 1803 1782 1809 1783
rect 1888 1774 1890 1784
rect 1894 1783 1895 1787
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1902 1787 1908 1788
rect 1902 1783 1903 1787
rect 1907 1786 1908 1787
rect 1915 1787 1921 1788
rect 1915 1786 1916 1787
rect 1907 1784 1916 1786
rect 1907 1783 1908 1784
rect 1902 1782 1908 1783
rect 1915 1783 1916 1784
rect 1920 1783 1921 1787
rect 1915 1782 1921 1783
rect 1998 1787 2004 1788
rect 1998 1783 1999 1787
rect 2003 1783 2004 1787
rect 1998 1782 2004 1783
rect 2019 1787 2025 1788
rect 2019 1783 2020 1787
rect 2024 1786 2025 1787
rect 2102 1787 2108 1788
rect 2024 1784 2086 1786
rect 2024 1783 2025 1784
rect 2019 1782 2025 1783
rect 2084 1774 2086 1784
rect 2102 1783 2103 1787
rect 2107 1783 2108 1787
rect 2102 1782 2108 1783
rect 2123 1787 2129 1788
rect 2123 1783 2124 1787
rect 2128 1786 2129 1787
rect 2198 1787 2204 1788
rect 2128 1784 2190 1786
rect 2128 1783 2129 1784
rect 2123 1782 2129 1783
rect 2188 1774 2190 1784
rect 2198 1783 2199 1787
rect 2203 1783 2204 1787
rect 2198 1782 2204 1783
rect 2219 1787 2225 1788
rect 2219 1783 2220 1787
rect 2224 1786 2225 1787
rect 2286 1787 2292 1788
rect 2224 1784 2278 1786
rect 2224 1783 2225 1784
rect 2219 1782 2225 1783
rect 2276 1774 2278 1784
rect 2286 1783 2287 1787
rect 2291 1783 2292 1787
rect 2286 1782 2292 1783
rect 2307 1787 2313 1788
rect 2307 1783 2308 1787
rect 2312 1786 2313 1787
rect 2382 1787 2388 1788
rect 2312 1784 2378 1786
rect 2312 1783 2313 1784
rect 2307 1782 2313 1783
rect 2376 1774 2378 1784
rect 2382 1783 2383 1787
rect 2387 1783 2388 1787
rect 2382 1782 2388 1783
rect 2402 1787 2409 1788
rect 2402 1783 2403 1787
rect 2408 1783 2409 1787
rect 2402 1782 2409 1783
rect 2454 1787 2460 1788
rect 2454 1783 2455 1787
rect 2459 1783 2460 1787
rect 2454 1782 2460 1783
rect 2462 1787 2468 1788
rect 2462 1783 2463 1787
rect 2467 1786 2468 1787
rect 2475 1787 2481 1788
rect 2475 1786 2476 1787
rect 2467 1784 2476 1786
rect 2467 1783 2468 1784
rect 2462 1782 2468 1783
rect 2475 1783 2476 1784
rect 2480 1783 2481 1787
rect 2502 1784 2503 1788
rect 2507 1784 2508 1788
rect 2502 1783 2508 1784
rect 2475 1782 2481 1783
rect 1483 1773 1489 1774
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 1286 1771 1292 1772
rect 110 1766 116 1767
rect 134 1768 140 1769
rect 134 1764 135 1768
rect 139 1764 140 1768
rect 134 1763 140 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 318 1768 324 1769
rect 318 1764 319 1768
rect 323 1764 324 1768
rect 318 1763 324 1764
rect 422 1768 428 1769
rect 422 1764 423 1768
rect 427 1764 428 1768
rect 422 1763 428 1764
rect 518 1768 524 1769
rect 518 1764 519 1768
rect 523 1764 524 1768
rect 518 1763 524 1764
rect 614 1768 620 1769
rect 614 1764 615 1768
rect 619 1764 620 1768
rect 614 1763 620 1764
rect 702 1768 708 1769
rect 702 1764 703 1768
rect 707 1764 708 1768
rect 702 1763 708 1764
rect 782 1768 788 1769
rect 782 1764 783 1768
rect 787 1764 788 1768
rect 782 1763 788 1764
rect 862 1768 868 1769
rect 862 1764 863 1768
rect 867 1764 868 1768
rect 862 1763 868 1764
rect 942 1768 948 1769
rect 942 1764 943 1768
rect 947 1764 948 1768
rect 942 1763 948 1764
rect 1022 1768 1028 1769
rect 1022 1764 1023 1768
rect 1027 1764 1028 1768
rect 1022 1763 1028 1764
rect 1102 1768 1108 1769
rect 1102 1764 1103 1768
rect 1107 1764 1108 1768
rect 1286 1767 1287 1771
rect 1291 1767 1292 1771
rect 1483 1769 1484 1773
rect 1488 1769 1489 1773
rect 1776 1773 1793 1774
rect 1776 1772 1788 1773
rect 1483 1768 1489 1769
rect 1579 1771 1585 1772
rect 1286 1766 1292 1767
rect 1579 1767 1580 1771
rect 1584 1770 1585 1771
rect 1683 1771 1689 1772
rect 1584 1768 1678 1770
rect 1584 1767 1585 1768
rect 1579 1766 1585 1767
rect 1102 1763 1108 1764
rect 1676 1762 1678 1768
rect 1683 1767 1684 1771
rect 1688 1770 1689 1771
rect 1694 1771 1700 1772
rect 1694 1770 1695 1771
rect 1688 1768 1695 1770
rect 1688 1767 1689 1768
rect 1683 1766 1689 1767
rect 1694 1767 1695 1768
rect 1699 1767 1700 1771
rect 1787 1769 1788 1772
rect 1792 1769 1793 1773
rect 1888 1773 1905 1774
rect 1888 1772 1900 1773
rect 1787 1768 1793 1769
rect 1899 1769 1900 1772
rect 1904 1769 1905 1773
rect 2084 1773 2113 1774
rect 2084 1772 2108 1773
rect 1899 1768 1905 1769
rect 2003 1771 2009 1772
rect 1694 1766 1700 1767
rect 2003 1767 2004 1771
rect 2008 1767 2009 1771
rect 2107 1769 2108 1772
rect 2112 1769 2113 1773
rect 2188 1773 2209 1774
rect 2188 1772 2204 1773
rect 2107 1768 2113 1769
rect 2203 1769 2204 1772
rect 2208 1769 2209 1773
rect 2276 1773 2297 1774
rect 2276 1772 2292 1773
rect 2203 1768 2209 1769
rect 2291 1769 2292 1772
rect 2296 1769 2297 1773
rect 2376 1773 2393 1774
rect 2376 1772 2388 1773
rect 2291 1768 2297 1769
rect 2387 1769 2388 1772
rect 2392 1769 2393 1773
rect 2387 1768 2393 1769
rect 2459 1771 2465 1772
rect 2003 1766 2009 1767
rect 2370 1767 2376 1768
rect 2370 1766 2371 1767
rect 2005 1764 2371 1766
rect 1902 1763 1908 1764
rect 1902 1762 1903 1763
rect 1676 1760 1903 1762
rect 1902 1759 1903 1760
rect 1907 1759 1908 1763
rect 2370 1763 2371 1764
rect 2375 1763 2376 1767
rect 2459 1767 2460 1771
rect 2464 1770 2465 1771
rect 2486 1771 2492 1772
rect 2486 1770 2487 1771
rect 2464 1768 2487 1770
rect 2464 1767 2465 1768
rect 2459 1766 2465 1767
rect 2486 1767 2487 1768
rect 2491 1767 2492 1771
rect 2486 1766 2492 1767
rect 2370 1762 2376 1763
rect 1902 1758 1908 1759
rect 1794 1755 1800 1756
rect 1794 1754 1795 1755
rect 134 1752 140 1753
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 134 1748 135 1752
rect 139 1748 140 1752
rect 134 1747 140 1748
rect 238 1752 244 1753
rect 238 1748 239 1752
rect 243 1748 244 1752
rect 238 1747 244 1748
rect 350 1752 356 1753
rect 350 1748 351 1752
rect 355 1748 356 1752
rect 350 1747 356 1748
rect 462 1752 468 1753
rect 462 1748 463 1752
rect 467 1748 468 1752
rect 462 1747 468 1748
rect 574 1752 580 1753
rect 574 1748 575 1752
rect 579 1748 580 1752
rect 574 1747 580 1748
rect 678 1752 684 1753
rect 678 1748 679 1752
rect 683 1748 684 1752
rect 678 1747 684 1748
rect 782 1752 788 1753
rect 782 1748 783 1752
rect 787 1748 788 1752
rect 782 1747 788 1748
rect 886 1752 892 1753
rect 886 1748 887 1752
rect 891 1748 892 1752
rect 886 1747 892 1748
rect 990 1752 996 1753
rect 990 1748 991 1752
rect 995 1748 996 1752
rect 990 1747 996 1748
rect 1102 1752 1108 1753
rect 1102 1748 1103 1752
rect 1107 1748 1108 1752
rect 1477 1752 1795 1754
rect 1477 1750 1479 1752
rect 1794 1751 1795 1752
rect 1799 1751 1800 1755
rect 2342 1755 2348 1756
rect 2342 1754 2343 1755
rect 1794 1750 1800 1751
rect 1892 1752 2343 1754
rect 1892 1750 1894 1752
rect 2342 1751 2343 1752
rect 2347 1751 2348 1755
rect 2342 1750 2348 1751
rect 1102 1747 1108 1748
rect 1286 1749 1292 1750
rect 110 1744 116 1745
rect 1286 1745 1287 1749
rect 1291 1745 1292 1749
rect 1475 1749 1481 1750
rect 1286 1744 1292 1745
rect 1379 1747 1385 1748
rect 1379 1743 1380 1747
rect 1384 1746 1385 1747
rect 1384 1744 1471 1746
rect 1475 1745 1476 1749
rect 1480 1745 1481 1749
rect 1891 1749 1897 1750
rect 1475 1744 1481 1745
rect 1558 1747 1564 1748
rect 1384 1743 1385 1744
rect 1379 1742 1385 1743
rect 1469 1738 1471 1744
rect 1558 1743 1559 1747
rect 1563 1746 1564 1747
rect 1571 1747 1577 1748
rect 1571 1746 1572 1747
rect 1563 1744 1572 1746
rect 1563 1743 1564 1744
rect 1558 1742 1564 1743
rect 1571 1743 1572 1744
rect 1576 1743 1577 1747
rect 1675 1747 1681 1748
rect 1675 1746 1676 1747
rect 1571 1742 1577 1743
rect 1588 1744 1676 1746
rect 1469 1736 1494 1738
rect 1492 1734 1494 1736
rect 1588 1734 1590 1744
rect 1675 1743 1676 1744
rect 1680 1743 1681 1747
rect 1779 1747 1785 1748
rect 1779 1746 1780 1747
rect 1675 1742 1681 1743
rect 1692 1744 1780 1746
rect 1692 1734 1694 1744
rect 1779 1743 1780 1744
rect 1784 1743 1785 1747
rect 1891 1745 1892 1749
rect 1896 1745 1897 1749
rect 2003 1747 2009 1748
rect 2003 1746 2004 1747
rect 1891 1744 1897 1745
rect 1999 1744 2004 1746
rect 1779 1742 1785 1743
rect 1999 1738 2001 1744
rect 2003 1743 2004 1744
rect 2008 1743 2009 1747
rect 2115 1747 2121 1748
rect 2115 1746 2116 1747
rect 2003 1742 2009 1743
rect 2020 1744 2116 1746
rect 1908 1736 2001 1738
rect 1908 1734 1910 1736
rect 2020 1734 2022 1744
rect 2115 1743 2116 1744
rect 2120 1743 2121 1747
rect 2235 1747 2241 1748
rect 2235 1746 2236 1747
rect 2115 1742 2121 1743
rect 2132 1744 2236 1746
rect 2132 1734 2134 1744
rect 2235 1743 2236 1744
rect 2240 1743 2241 1747
rect 2355 1747 2361 1748
rect 2355 1746 2356 1747
rect 2235 1742 2241 1743
rect 2252 1744 2356 1746
rect 2252 1734 2254 1744
rect 2355 1743 2356 1744
rect 2360 1743 2361 1747
rect 2355 1742 2361 1743
rect 2459 1747 2468 1748
rect 2459 1743 2460 1747
rect 2467 1743 2468 1747
rect 2459 1742 2468 1743
rect 1374 1733 1380 1734
rect 110 1732 116 1733
rect 1286 1732 1292 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 150 1731 156 1732
rect 150 1727 151 1731
rect 155 1727 156 1731
rect 150 1726 156 1727
rect 171 1731 177 1732
rect 171 1727 172 1731
rect 176 1730 177 1731
rect 182 1731 188 1732
rect 182 1730 183 1731
rect 176 1728 183 1730
rect 176 1727 177 1728
rect 171 1726 177 1727
rect 182 1727 183 1728
rect 187 1727 188 1731
rect 182 1726 188 1727
rect 254 1731 260 1732
rect 254 1727 255 1731
rect 259 1727 260 1731
rect 275 1731 281 1732
rect 275 1730 276 1731
rect 254 1726 260 1727
rect 264 1728 276 1730
rect 264 1722 266 1728
rect 275 1727 276 1728
rect 280 1727 281 1731
rect 275 1726 281 1727
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 387 1731 393 1732
rect 387 1730 388 1731
rect 366 1726 372 1727
rect 376 1728 388 1730
rect 376 1722 378 1728
rect 387 1727 388 1728
rect 392 1727 393 1731
rect 387 1726 393 1727
rect 478 1731 484 1732
rect 478 1727 479 1731
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 498 1731 505 1732
rect 498 1727 499 1731
rect 504 1727 505 1731
rect 498 1726 505 1727
rect 590 1731 596 1732
rect 590 1727 591 1731
rect 595 1727 596 1731
rect 590 1726 596 1727
rect 611 1731 617 1732
rect 611 1727 612 1731
rect 616 1727 617 1731
rect 611 1726 617 1727
rect 694 1731 700 1732
rect 694 1727 695 1731
rect 699 1727 700 1731
rect 694 1726 700 1727
rect 715 1731 721 1732
rect 715 1727 716 1731
rect 720 1730 721 1731
rect 734 1731 740 1732
rect 734 1730 735 1731
rect 720 1728 735 1730
rect 720 1727 721 1728
rect 715 1726 721 1727
rect 734 1727 735 1728
rect 739 1727 740 1731
rect 734 1726 740 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 819 1731 825 1732
rect 819 1727 820 1731
rect 824 1727 825 1731
rect 819 1726 825 1727
rect 902 1731 908 1732
rect 902 1727 903 1731
rect 907 1727 908 1731
rect 902 1726 908 1727
rect 918 1731 929 1732
rect 918 1727 919 1731
rect 923 1727 924 1731
rect 928 1727 929 1731
rect 918 1726 929 1727
rect 1006 1731 1012 1732
rect 1006 1727 1007 1731
rect 1011 1727 1012 1731
rect 1027 1731 1033 1732
rect 1027 1730 1028 1731
rect 1006 1726 1012 1727
rect 1016 1728 1028 1730
rect 613 1722 615 1726
rect 821 1722 823 1726
rect 1016 1722 1018 1728
rect 1027 1727 1028 1728
rect 1032 1727 1033 1731
rect 1027 1726 1033 1727
rect 1118 1731 1124 1732
rect 1118 1727 1119 1731
rect 1123 1727 1124 1731
rect 1118 1726 1124 1727
rect 1138 1731 1145 1732
rect 1138 1727 1139 1731
rect 1144 1727 1145 1731
rect 1286 1728 1287 1732
rect 1291 1728 1292 1732
rect 1286 1727 1292 1728
rect 1326 1732 1332 1733
rect 1326 1728 1327 1732
rect 1331 1728 1332 1732
rect 1374 1729 1375 1733
rect 1379 1729 1380 1733
rect 1470 1733 1476 1734
rect 1374 1728 1380 1729
rect 1395 1731 1401 1732
rect 1326 1727 1332 1728
rect 1395 1727 1396 1731
rect 1400 1730 1401 1731
rect 1438 1731 1444 1732
rect 1438 1730 1439 1731
rect 1400 1728 1439 1730
rect 1400 1727 1401 1728
rect 1138 1726 1145 1727
rect 1395 1726 1401 1727
rect 1438 1727 1439 1728
rect 1443 1727 1444 1731
rect 1470 1729 1471 1733
rect 1475 1729 1476 1733
rect 1470 1728 1476 1729
rect 1491 1733 1497 1734
rect 1491 1729 1492 1733
rect 1496 1729 1497 1733
rect 1491 1728 1497 1729
rect 1566 1733 1572 1734
rect 1566 1729 1567 1733
rect 1571 1729 1572 1733
rect 1566 1728 1572 1729
rect 1587 1733 1593 1734
rect 1587 1729 1588 1733
rect 1592 1729 1593 1733
rect 1587 1728 1593 1729
rect 1670 1733 1676 1734
rect 1670 1729 1671 1733
rect 1675 1729 1676 1733
rect 1670 1728 1676 1729
rect 1691 1733 1697 1734
rect 1691 1729 1692 1733
rect 1696 1729 1697 1733
rect 1691 1728 1697 1729
rect 1774 1733 1780 1734
rect 1774 1729 1775 1733
rect 1779 1729 1780 1733
rect 1886 1733 1892 1734
rect 1774 1728 1780 1729
rect 1794 1731 1801 1732
rect 1438 1726 1444 1727
rect 1794 1727 1795 1731
rect 1800 1727 1801 1731
rect 1886 1729 1887 1733
rect 1891 1729 1892 1733
rect 1886 1728 1892 1729
rect 1907 1733 1913 1734
rect 1907 1729 1908 1733
rect 1912 1729 1913 1733
rect 1907 1728 1913 1729
rect 1998 1733 2004 1734
rect 1998 1729 1999 1733
rect 2003 1729 2004 1733
rect 1998 1728 2004 1729
rect 2019 1733 2025 1734
rect 2019 1729 2020 1733
rect 2024 1729 2025 1733
rect 2019 1728 2025 1729
rect 2110 1733 2116 1734
rect 2110 1729 2111 1733
rect 2115 1729 2116 1733
rect 2110 1728 2116 1729
rect 2131 1733 2137 1734
rect 2131 1729 2132 1733
rect 2136 1729 2137 1733
rect 2131 1728 2137 1729
rect 2230 1733 2236 1734
rect 2230 1729 2231 1733
rect 2235 1729 2236 1733
rect 2230 1728 2236 1729
rect 2251 1733 2257 1734
rect 2251 1729 2252 1733
rect 2256 1729 2257 1733
rect 2251 1728 2257 1729
rect 2350 1733 2356 1734
rect 2350 1729 2351 1733
rect 2355 1729 2356 1733
rect 2454 1733 2460 1734
rect 2350 1728 2356 1729
rect 2370 1731 2377 1732
rect 1794 1726 1801 1727
rect 2370 1727 2371 1731
rect 2376 1727 2377 1731
rect 2454 1729 2455 1733
rect 2459 1729 2460 1733
rect 2502 1732 2508 1733
rect 2454 1728 2460 1729
rect 2470 1731 2481 1732
rect 2370 1726 2377 1727
rect 2470 1727 2471 1731
rect 2475 1727 2476 1731
rect 2480 1727 2481 1731
rect 2502 1728 2503 1732
rect 2507 1728 2508 1732
rect 2502 1727 2508 1728
rect 2470 1726 2481 1727
rect 157 1720 266 1722
rect 319 1720 378 1722
rect 484 1720 615 1722
rect 701 1720 823 1722
rect 908 1720 1018 1722
rect 157 1718 159 1720
rect 319 1718 321 1720
rect 484 1718 486 1720
rect 701 1718 703 1720
rect 908 1718 910 1720
rect 155 1717 161 1718
rect 155 1713 156 1717
rect 160 1713 161 1717
rect 155 1712 161 1713
rect 259 1717 321 1718
rect 259 1713 260 1717
rect 264 1716 321 1717
rect 483 1717 489 1718
rect 264 1713 265 1716
rect 259 1712 265 1713
rect 358 1715 364 1716
rect 358 1711 359 1715
rect 363 1714 364 1715
rect 371 1715 377 1716
rect 371 1714 372 1715
rect 363 1712 372 1714
rect 363 1711 364 1712
rect 358 1710 364 1711
rect 371 1711 372 1712
rect 376 1711 377 1715
rect 483 1713 484 1717
rect 488 1713 489 1717
rect 699 1717 705 1718
rect 483 1712 489 1713
rect 595 1715 601 1716
rect 371 1710 377 1711
rect 595 1711 596 1715
rect 600 1714 601 1715
rect 658 1715 664 1716
rect 658 1714 659 1715
rect 600 1712 659 1714
rect 600 1711 601 1712
rect 595 1710 601 1711
rect 658 1711 659 1712
rect 663 1711 664 1715
rect 699 1713 700 1717
rect 704 1713 705 1717
rect 907 1717 913 1718
rect 699 1712 705 1713
rect 803 1715 809 1716
rect 658 1710 664 1711
rect 803 1711 804 1715
rect 808 1711 809 1715
rect 907 1713 908 1717
rect 912 1713 913 1717
rect 907 1712 913 1713
rect 998 1715 1004 1716
rect 803 1710 809 1711
rect 918 1711 924 1712
rect 918 1710 919 1711
rect 805 1708 919 1710
rect 918 1707 919 1708
rect 923 1707 924 1711
rect 998 1711 999 1715
rect 1003 1714 1004 1715
rect 1011 1715 1017 1716
rect 1011 1714 1012 1715
rect 1003 1712 1012 1714
rect 1003 1711 1004 1712
rect 998 1710 1004 1711
rect 1011 1711 1012 1712
rect 1016 1711 1017 1715
rect 1011 1710 1017 1711
rect 1123 1715 1129 1716
rect 1123 1711 1124 1715
rect 1128 1714 1129 1715
rect 1194 1715 1200 1716
rect 1194 1714 1195 1715
rect 1128 1712 1195 1714
rect 1128 1711 1129 1712
rect 1123 1710 1129 1711
rect 1194 1711 1195 1712
rect 1199 1711 1200 1715
rect 1194 1710 1200 1711
rect 1326 1715 1332 1716
rect 1326 1711 1327 1715
rect 1331 1711 1332 1715
rect 2502 1715 2508 1716
rect 1326 1710 1332 1711
rect 1358 1712 1364 1713
rect 1358 1708 1359 1712
rect 1363 1708 1364 1712
rect 1358 1707 1364 1708
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1550 1712 1556 1713
rect 1550 1708 1551 1712
rect 1555 1708 1556 1712
rect 1550 1707 1556 1708
rect 1654 1712 1660 1713
rect 1654 1708 1655 1712
rect 1659 1708 1660 1712
rect 1654 1707 1660 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1870 1712 1876 1713
rect 1870 1708 1871 1712
rect 1875 1708 1876 1712
rect 1870 1707 1876 1708
rect 1982 1712 1988 1713
rect 1982 1708 1983 1712
rect 1987 1708 1988 1712
rect 1982 1707 1988 1708
rect 2094 1712 2100 1713
rect 2094 1708 2095 1712
rect 2099 1708 2100 1712
rect 2094 1707 2100 1708
rect 2214 1712 2220 1713
rect 2214 1708 2215 1712
rect 2219 1708 2220 1712
rect 2214 1707 2220 1708
rect 2334 1712 2340 1713
rect 2334 1708 2335 1712
rect 2339 1708 2340 1712
rect 2334 1707 2340 1708
rect 2438 1712 2444 1713
rect 2438 1708 2439 1712
rect 2443 1708 2444 1712
rect 2502 1711 2503 1715
rect 2507 1711 2508 1715
rect 2502 1710 2508 1711
rect 2438 1707 2444 1708
rect 918 1706 924 1707
rect 1350 1700 1356 1701
rect 1326 1697 1332 1698
rect 1326 1693 1327 1697
rect 1331 1693 1332 1697
rect 1350 1696 1351 1700
rect 1355 1696 1356 1700
rect 1350 1695 1356 1696
rect 1430 1700 1436 1701
rect 1430 1696 1431 1700
rect 1435 1696 1436 1700
rect 1430 1695 1436 1696
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1646 1700 1652 1701
rect 1646 1696 1647 1700
rect 1651 1696 1652 1700
rect 1646 1695 1652 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 2014 1700 2020 1701
rect 2014 1696 2015 1700
rect 2019 1696 2020 1700
rect 2014 1695 2020 1696
rect 2158 1700 2164 1701
rect 2158 1696 2159 1700
rect 2163 1696 2164 1700
rect 2158 1695 2164 1696
rect 2310 1700 2316 1701
rect 2310 1696 2311 1700
rect 2315 1696 2316 1700
rect 2310 1695 2316 1696
rect 2438 1700 2444 1701
rect 2438 1696 2439 1700
rect 2443 1696 2444 1700
rect 2438 1695 2444 1696
rect 2502 1697 2508 1698
rect 1326 1692 1332 1693
rect 2502 1693 2503 1697
rect 2507 1693 2508 1697
rect 2502 1692 2508 1693
rect 182 1691 188 1692
rect 182 1687 183 1691
rect 187 1690 188 1691
rect 195 1691 201 1692
rect 195 1690 196 1691
rect 187 1688 196 1690
rect 187 1687 188 1688
rect 182 1686 188 1687
rect 195 1687 196 1688
rect 200 1687 201 1691
rect 275 1691 281 1692
rect 275 1690 276 1691
rect 195 1686 201 1687
rect 245 1688 276 1690
rect 245 1682 247 1688
rect 275 1687 276 1688
rect 280 1687 281 1691
rect 355 1691 361 1692
rect 355 1690 356 1691
rect 275 1686 281 1687
rect 319 1688 356 1690
rect 319 1682 321 1688
rect 355 1687 356 1688
rect 360 1687 361 1691
rect 355 1686 361 1687
rect 443 1691 452 1692
rect 443 1687 444 1691
rect 451 1687 452 1691
rect 539 1691 545 1692
rect 539 1690 540 1691
rect 443 1686 452 1687
rect 460 1688 540 1690
rect 212 1680 247 1682
rect 292 1680 321 1682
rect 212 1678 214 1680
rect 292 1678 294 1680
rect 460 1678 462 1688
rect 539 1687 540 1688
rect 544 1687 545 1691
rect 643 1691 649 1692
rect 643 1690 644 1691
rect 539 1686 545 1687
rect 564 1688 644 1690
rect 564 1682 566 1688
rect 643 1687 644 1688
rect 648 1687 649 1691
rect 643 1686 649 1687
rect 734 1691 740 1692
rect 734 1687 735 1691
rect 739 1690 740 1691
rect 747 1691 753 1692
rect 747 1690 748 1691
rect 739 1688 748 1690
rect 739 1687 740 1688
rect 734 1686 740 1687
rect 747 1687 748 1688
rect 752 1687 753 1691
rect 851 1691 857 1692
rect 851 1690 852 1691
rect 747 1686 753 1687
rect 788 1688 852 1690
rect 556 1680 566 1682
rect 556 1678 558 1680
rect 788 1678 790 1688
rect 851 1687 852 1688
rect 856 1687 857 1691
rect 955 1691 961 1692
rect 955 1690 956 1691
rect 851 1686 857 1687
rect 869 1688 956 1690
rect 869 1678 871 1688
rect 955 1687 956 1688
rect 960 1687 961 1691
rect 955 1686 961 1687
rect 1067 1691 1073 1692
rect 1067 1687 1068 1691
rect 1072 1690 1073 1691
rect 1090 1691 1096 1692
rect 1090 1690 1091 1691
rect 1072 1688 1091 1690
rect 1072 1687 1073 1688
rect 1067 1686 1073 1687
rect 1090 1687 1091 1688
rect 1095 1687 1096 1691
rect 1179 1691 1185 1692
rect 1179 1690 1180 1691
rect 1090 1686 1096 1687
rect 1159 1688 1180 1690
rect 1159 1682 1161 1688
rect 1179 1687 1180 1688
rect 1184 1687 1185 1691
rect 1179 1686 1185 1687
rect 1084 1680 1161 1682
rect 1326 1680 1332 1681
rect 2502 1680 2508 1681
rect 1084 1678 1086 1680
rect 190 1677 196 1678
rect 110 1676 116 1677
rect 110 1672 111 1676
rect 115 1672 116 1676
rect 190 1673 191 1677
rect 195 1673 196 1677
rect 190 1672 196 1673
rect 211 1677 217 1678
rect 211 1673 212 1677
rect 216 1673 217 1677
rect 211 1672 217 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 291 1677 297 1678
rect 291 1673 292 1677
rect 296 1673 297 1677
rect 291 1672 297 1673
rect 350 1677 356 1678
rect 350 1673 351 1677
rect 355 1673 356 1677
rect 438 1677 444 1678
rect 350 1672 356 1673
rect 358 1675 364 1676
rect 110 1671 116 1672
rect 358 1671 359 1675
rect 363 1674 364 1675
rect 371 1675 377 1676
rect 371 1674 372 1675
rect 363 1672 372 1674
rect 363 1671 364 1672
rect 358 1670 364 1671
rect 371 1671 372 1672
rect 376 1671 377 1675
rect 438 1673 439 1677
rect 443 1673 444 1677
rect 438 1672 444 1673
rect 459 1677 465 1678
rect 459 1673 460 1677
rect 464 1673 465 1677
rect 459 1672 465 1673
rect 534 1677 540 1678
rect 534 1673 535 1677
rect 539 1673 540 1677
rect 534 1672 540 1673
rect 555 1677 561 1678
rect 555 1673 556 1677
rect 560 1673 561 1677
rect 555 1672 561 1673
rect 638 1677 644 1678
rect 638 1673 639 1677
rect 643 1673 644 1677
rect 742 1677 748 1678
rect 638 1672 644 1673
rect 658 1675 665 1676
rect 371 1670 377 1671
rect 658 1671 659 1675
rect 664 1671 665 1675
rect 742 1673 743 1677
rect 747 1673 748 1677
rect 742 1672 748 1673
rect 763 1677 790 1678
rect 763 1673 764 1677
rect 768 1676 790 1677
rect 846 1677 852 1678
rect 768 1673 769 1676
rect 763 1672 769 1673
rect 846 1673 847 1677
rect 851 1673 852 1677
rect 846 1672 852 1673
rect 867 1677 873 1678
rect 867 1673 868 1677
rect 872 1673 873 1677
rect 867 1672 873 1673
rect 950 1677 956 1678
rect 950 1673 951 1677
rect 955 1673 956 1677
rect 1062 1677 1068 1678
rect 950 1672 956 1673
rect 966 1675 977 1676
rect 658 1670 665 1671
rect 966 1671 967 1675
rect 971 1671 972 1675
rect 976 1671 977 1675
rect 1062 1673 1063 1677
rect 1067 1673 1068 1677
rect 1062 1672 1068 1673
rect 1083 1677 1089 1678
rect 1083 1673 1084 1677
rect 1088 1673 1089 1677
rect 1083 1672 1089 1673
rect 1174 1677 1180 1678
rect 1174 1673 1175 1677
rect 1179 1673 1180 1677
rect 1286 1676 1292 1677
rect 1174 1672 1180 1673
rect 1194 1675 1201 1676
rect 966 1670 977 1671
rect 1194 1671 1195 1675
rect 1200 1671 1201 1675
rect 1286 1672 1287 1676
rect 1291 1672 1292 1676
rect 1326 1676 1327 1680
rect 1331 1676 1332 1680
rect 1326 1675 1332 1676
rect 1366 1679 1372 1680
rect 1366 1675 1367 1679
rect 1371 1675 1372 1679
rect 1366 1674 1372 1675
rect 1374 1679 1380 1680
rect 1374 1675 1375 1679
rect 1379 1678 1380 1679
rect 1387 1679 1393 1680
rect 1387 1678 1388 1679
rect 1379 1676 1388 1678
rect 1379 1675 1380 1676
rect 1374 1674 1380 1675
rect 1387 1675 1388 1676
rect 1392 1675 1393 1679
rect 1387 1674 1393 1675
rect 1446 1679 1452 1680
rect 1446 1675 1447 1679
rect 1451 1675 1452 1679
rect 1446 1674 1452 1675
rect 1467 1679 1473 1680
rect 1467 1675 1468 1679
rect 1472 1675 1473 1679
rect 1467 1674 1473 1675
rect 1550 1679 1556 1680
rect 1550 1675 1551 1679
rect 1555 1675 1556 1679
rect 1550 1674 1556 1675
rect 1571 1679 1577 1680
rect 1571 1675 1572 1679
rect 1576 1678 1577 1679
rect 1662 1679 1668 1680
rect 1576 1676 1654 1678
rect 1576 1675 1577 1676
rect 1571 1674 1577 1675
rect 1286 1671 1292 1672
rect 1194 1670 1201 1671
rect 1469 1666 1471 1674
rect 1652 1666 1654 1676
rect 1662 1675 1663 1679
rect 1667 1675 1668 1679
rect 1662 1674 1668 1675
rect 1670 1679 1676 1680
rect 1670 1675 1671 1679
rect 1675 1678 1676 1679
rect 1683 1679 1689 1680
rect 1683 1678 1684 1679
rect 1675 1676 1684 1678
rect 1675 1675 1676 1676
rect 1670 1674 1676 1675
rect 1683 1675 1684 1676
rect 1688 1675 1689 1679
rect 1683 1674 1689 1675
rect 1774 1679 1780 1680
rect 1774 1675 1775 1679
rect 1779 1675 1780 1679
rect 1774 1674 1780 1675
rect 1795 1679 1801 1680
rect 1795 1675 1796 1679
rect 1800 1678 1801 1679
rect 1894 1679 1900 1680
rect 1800 1676 1890 1678
rect 1800 1675 1801 1676
rect 1795 1674 1801 1675
rect 1888 1666 1890 1676
rect 1894 1675 1895 1679
rect 1899 1675 1900 1679
rect 1894 1674 1900 1675
rect 1915 1679 1921 1680
rect 1915 1675 1916 1679
rect 1920 1678 1921 1679
rect 2030 1679 2036 1680
rect 1920 1676 2001 1678
rect 1920 1675 1921 1676
rect 1915 1674 1921 1675
rect 1999 1666 2001 1676
rect 2030 1675 2031 1679
rect 2035 1675 2036 1679
rect 2030 1674 2036 1675
rect 2051 1679 2057 1680
rect 2051 1675 2052 1679
rect 2056 1678 2057 1679
rect 2174 1679 2180 1680
rect 2056 1676 2170 1678
rect 2056 1675 2057 1676
rect 2051 1674 2057 1675
rect 2168 1670 2170 1676
rect 2174 1675 2175 1679
rect 2179 1675 2180 1679
rect 2174 1674 2180 1675
rect 2195 1679 2201 1680
rect 2195 1675 2196 1679
rect 2200 1678 2201 1679
rect 2326 1679 2332 1680
rect 2200 1676 2322 1678
rect 2200 1675 2201 1676
rect 2195 1674 2201 1675
rect 2168 1668 2183 1670
rect 2181 1666 2183 1668
rect 2320 1666 2322 1676
rect 2326 1675 2327 1679
rect 2331 1675 2332 1679
rect 2326 1674 2332 1675
rect 2342 1679 2353 1680
rect 2342 1675 2343 1679
rect 2347 1675 2348 1679
rect 2352 1675 2353 1679
rect 2342 1674 2353 1675
rect 2454 1679 2460 1680
rect 2454 1675 2455 1679
rect 2459 1675 2460 1679
rect 2454 1674 2460 1675
rect 2462 1679 2468 1680
rect 2462 1675 2463 1679
rect 2467 1678 2468 1679
rect 2475 1679 2481 1680
rect 2475 1678 2476 1679
rect 2467 1676 2476 1678
rect 2467 1675 2468 1676
rect 2462 1674 2468 1675
rect 2475 1675 2476 1676
rect 2480 1675 2481 1679
rect 2502 1676 2503 1680
rect 2507 1676 2508 1680
rect 2502 1675 2508 1676
rect 2475 1674 2481 1675
rect 1469 1665 1561 1666
rect 1469 1664 1556 1665
rect 1371 1663 1377 1664
rect 110 1659 116 1660
rect 110 1655 111 1659
rect 115 1655 116 1659
rect 1286 1659 1292 1660
rect 110 1654 116 1655
rect 174 1656 180 1657
rect 174 1652 175 1656
rect 179 1652 180 1656
rect 174 1651 180 1652
rect 254 1656 260 1657
rect 254 1652 255 1656
rect 259 1652 260 1656
rect 254 1651 260 1652
rect 334 1656 340 1657
rect 334 1652 335 1656
rect 339 1652 340 1656
rect 334 1651 340 1652
rect 422 1656 428 1657
rect 422 1652 423 1656
rect 427 1652 428 1656
rect 422 1651 428 1652
rect 518 1656 524 1657
rect 518 1652 519 1656
rect 523 1652 524 1656
rect 518 1651 524 1652
rect 622 1656 628 1657
rect 622 1652 623 1656
rect 627 1652 628 1656
rect 622 1651 628 1652
rect 726 1656 732 1657
rect 726 1652 727 1656
rect 731 1652 732 1656
rect 726 1651 732 1652
rect 830 1656 836 1657
rect 830 1652 831 1656
rect 835 1652 836 1656
rect 830 1651 836 1652
rect 934 1656 940 1657
rect 934 1652 935 1656
rect 939 1652 940 1656
rect 934 1651 940 1652
rect 1046 1656 1052 1657
rect 1046 1652 1047 1656
rect 1051 1652 1052 1656
rect 1046 1651 1052 1652
rect 1158 1656 1164 1657
rect 1158 1652 1159 1656
rect 1163 1652 1164 1656
rect 1286 1655 1287 1659
rect 1291 1655 1292 1659
rect 1371 1659 1372 1663
rect 1376 1662 1377 1663
rect 1382 1663 1388 1664
rect 1382 1662 1383 1663
rect 1376 1660 1383 1662
rect 1376 1659 1377 1660
rect 1371 1658 1377 1659
rect 1382 1659 1383 1660
rect 1387 1659 1388 1663
rect 1382 1658 1388 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1662 1444 1663
rect 1451 1663 1457 1664
rect 1451 1662 1452 1663
rect 1443 1660 1452 1662
rect 1443 1659 1444 1660
rect 1438 1658 1444 1659
rect 1451 1659 1452 1660
rect 1456 1659 1457 1663
rect 1555 1661 1556 1664
rect 1560 1661 1561 1665
rect 1652 1665 1673 1666
rect 1652 1664 1668 1665
rect 1555 1660 1561 1661
rect 1667 1661 1668 1664
rect 1672 1661 1673 1665
rect 1888 1665 1905 1666
rect 1888 1664 1900 1665
rect 1667 1660 1673 1661
rect 1779 1663 1785 1664
rect 1451 1658 1457 1659
rect 1779 1659 1780 1663
rect 1784 1662 1785 1663
rect 1784 1660 1894 1662
rect 1899 1661 1900 1664
rect 1904 1661 1905 1665
rect 1999 1665 2041 1666
rect 1999 1664 2036 1665
rect 1899 1660 1905 1661
rect 2035 1661 2036 1664
rect 2040 1661 2041 1665
rect 2035 1660 2041 1661
rect 2179 1665 2185 1666
rect 2179 1661 2180 1665
rect 2184 1661 2185 1665
rect 2320 1665 2337 1666
rect 2320 1664 2332 1665
rect 2179 1660 2185 1661
rect 2331 1661 2332 1664
rect 2336 1661 2337 1665
rect 2331 1660 2337 1661
rect 2459 1663 2465 1664
rect 1784 1659 1785 1660
rect 1779 1658 1785 1659
rect 1892 1658 1894 1660
rect 2346 1659 2352 1660
rect 2346 1658 2347 1659
rect 1892 1656 2347 1658
rect 1286 1654 1292 1655
rect 2346 1655 2347 1656
rect 2351 1655 2352 1659
rect 2459 1659 2460 1663
rect 2464 1662 2465 1663
rect 2470 1663 2476 1664
rect 2470 1662 2471 1663
rect 2464 1660 2471 1662
rect 2464 1659 2465 1660
rect 2459 1658 2465 1659
rect 2470 1659 2471 1660
rect 2475 1659 2476 1663
rect 2470 1658 2476 1659
rect 2346 1654 2352 1655
rect 1158 1651 1164 1652
rect 214 1644 220 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 270 1644 276 1645
rect 270 1640 271 1644
rect 275 1640 276 1644
rect 270 1639 276 1640
rect 334 1644 340 1645
rect 334 1640 335 1644
rect 339 1640 340 1644
rect 334 1639 340 1640
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 478 1644 484 1645
rect 478 1640 479 1644
rect 483 1640 484 1644
rect 478 1639 484 1640
rect 558 1644 564 1645
rect 558 1640 559 1644
rect 563 1640 564 1644
rect 558 1639 564 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 742 1644 748 1645
rect 742 1640 743 1644
rect 747 1640 748 1644
rect 742 1639 748 1640
rect 838 1644 844 1645
rect 838 1640 839 1644
rect 843 1640 844 1644
rect 838 1639 844 1640
rect 942 1644 948 1645
rect 942 1640 943 1644
rect 947 1640 948 1644
rect 942 1639 948 1640
rect 1054 1644 1060 1645
rect 1054 1640 1055 1644
rect 1059 1640 1060 1644
rect 1054 1639 1060 1640
rect 1174 1644 1180 1645
rect 1174 1640 1175 1644
rect 1179 1640 1180 1644
rect 2138 1643 2144 1644
rect 2138 1642 2139 1643
rect 1174 1639 1180 1640
rect 1286 1641 1292 1642
rect 110 1636 116 1637
rect 1286 1637 1287 1641
rect 1291 1637 1292 1641
rect 1604 1640 2139 1642
rect 1604 1638 1606 1640
rect 2138 1639 2139 1640
rect 2143 1639 2144 1643
rect 2138 1638 2144 1639
rect 1286 1636 1292 1637
rect 1603 1637 1609 1638
rect 1371 1635 1380 1636
rect 1371 1631 1372 1635
rect 1379 1631 1380 1635
rect 1435 1635 1441 1636
rect 1435 1634 1436 1635
rect 1371 1630 1380 1631
rect 1389 1632 1436 1634
rect 110 1624 116 1625
rect 1286 1624 1292 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 230 1623 236 1624
rect 230 1619 231 1623
rect 235 1619 236 1623
rect 230 1618 236 1619
rect 251 1623 257 1624
rect 251 1619 252 1623
rect 256 1622 257 1623
rect 286 1623 292 1624
rect 256 1620 282 1622
rect 256 1619 257 1620
rect 251 1618 257 1619
rect 280 1610 282 1620
rect 286 1619 287 1623
rect 291 1619 292 1623
rect 286 1618 292 1619
rect 294 1623 300 1624
rect 294 1619 295 1623
rect 299 1622 300 1623
rect 307 1623 313 1624
rect 307 1622 308 1623
rect 299 1620 308 1622
rect 299 1619 300 1620
rect 294 1618 300 1619
rect 307 1619 308 1620
rect 312 1619 313 1623
rect 307 1618 313 1619
rect 350 1623 356 1624
rect 350 1619 351 1623
rect 355 1619 356 1623
rect 371 1623 377 1624
rect 371 1622 372 1623
rect 350 1618 356 1619
rect 360 1620 372 1622
rect 360 1614 362 1620
rect 371 1619 372 1620
rect 376 1619 377 1623
rect 371 1618 377 1619
rect 422 1623 428 1624
rect 422 1619 423 1623
rect 427 1619 428 1623
rect 422 1618 428 1619
rect 443 1623 452 1624
rect 443 1619 444 1623
rect 451 1619 452 1623
rect 443 1618 452 1619
rect 494 1623 500 1624
rect 494 1619 495 1623
rect 499 1619 500 1623
rect 515 1623 521 1624
rect 515 1622 516 1623
rect 494 1618 500 1619
rect 504 1620 516 1622
rect 504 1614 506 1620
rect 515 1619 516 1620
rect 520 1619 521 1623
rect 515 1618 521 1619
rect 574 1623 580 1624
rect 574 1619 575 1623
rect 579 1619 580 1623
rect 595 1623 601 1624
rect 595 1622 596 1623
rect 574 1618 580 1619
rect 584 1620 596 1622
rect 584 1614 586 1620
rect 595 1619 596 1620
rect 600 1619 601 1623
rect 595 1618 601 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 683 1623 689 1624
rect 683 1619 684 1623
rect 688 1622 689 1623
rect 758 1623 764 1624
rect 688 1620 750 1622
rect 688 1619 689 1620
rect 683 1618 689 1619
rect 319 1612 362 1614
rect 428 1612 506 1614
rect 520 1612 586 1614
rect 280 1609 297 1610
rect 280 1608 292 1609
rect 235 1607 241 1608
rect 235 1603 236 1607
rect 240 1606 241 1607
rect 240 1604 278 1606
rect 291 1605 292 1608
rect 296 1605 297 1609
rect 291 1604 297 1605
rect 240 1603 241 1604
rect 235 1602 241 1603
rect 276 1602 278 1604
rect 319 1602 321 1612
rect 428 1610 430 1612
rect 520 1610 522 1612
rect 427 1609 433 1610
rect 355 1607 364 1608
rect 355 1603 356 1607
rect 363 1603 364 1607
rect 427 1605 428 1609
rect 432 1605 433 1609
rect 427 1604 433 1605
rect 499 1609 522 1610
rect 499 1605 500 1609
rect 504 1608 522 1609
rect 748 1610 750 1620
rect 758 1619 759 1623
rect 763 1619 764 1623
rect 758 1618 764 1619
rect 779 1623 785 1624
rect 779 1619 780 1623
rect 784 1622 785 1623
rect 806 1623 812 1624
rect 806 1622 807 1623
rect 784 1620 807 1622
rect 784 1619 785 1620
rect 779 1618 785 1619
rect 806 1619 807 1620
rect 811 1619 812 1623
rect 806 1618 812 1619
rect 854 1623 860 1624
rect 854 1619 855 1623
rect 859 1619 860 1623
rect 854 1618 860 1619
rect 870 1623 881 1624
rect 870 1619 871 1623
rect 875 1619 876 1623
rect 880 1619 881 1623
rect 870 1618 881 1619
rect 958 1623 964 1624
rect 958 1619 959 1623
rect 963 1619 964 1623
rect 979 1623 985 1624
rect 979 1622 980 1623
rect 958 1618 964 1619
rect 968 1620 980 1622
rect 968 1614 970 1620
rect 979 1619 980 1620
rect 984 1619 985 1623
rect 979 1618 985 1619
rect 1070 1623 1076 1624
rect 1070 1619 1071 1623
rect 1075 1619 1076 1623
rect 1070 1618 1076 1619
rect 1090 1623 1097 1624
rect 1090 1619 1091 1623
rect 1096 1619 1097 1623
rect 1090 1618 1097 1619
rect 1190 1623 1196 1624
rect 1190 1619 1191 1623
rect 1195 1619 1196 1623
rect 1211 1623 1217 1624
rect 1211 1622 1212 1623
rect 1190 1618 1196 1619
rect 1200 1620 1212 1622
rect 1200 1614 1202 1620
rect 1211 1619 1212 1620
rect 1216 1619 1217 1623
rect 1286 1620 1287 1624
rect 1291 1620 1292 1624
rect 1389 1622 1391 1632
rect 1435 1631 1436 1632
rect 1440 1631 1441 1635
rect 1523 1635 1529 1636
rect 1523 1634 1524 1635
rect 1435 1630 1441 1631
rect 1452 1632 1524 1634
rect 1452 1622 1454 1632
rect 1523 1631 1524 1632
rect 1528 1631 1529 1635
rect 1603 1633 1604 1637
rect 1608 1633 1609 1637
rect 1683 1635 1689 1636
rect 1683 1634 1684 1635
rect 1603 1632 1609 1633
rect 1620 1632 1684 1634
rect 1523 1630 1529 1631
rect 1620 1622 1622 1632
rect 1683 1631 1684 1632
rect 1688 1631 1689 1635
rect 1755 1635 1761 1636
rect 1755 1634 1756 1635
rect 1683 1630 1689 1631
rect 1700 1632 1756 1634
rect 1700 1622 1702 1632
rect 1755 1631 1756 1632
rect 1760 1631 1761 1635
rect 1843 1635 1849 1636
rect 1843 1634 1844 1635
rect 1755 1630 1761 1631
rect 1772 1632 1844 1634
rect 1772 1622 1774 1632
rect 1843 1631 1844 1632
rect 1848 1631 1849 1635
rect 1939 1635 1945 1636
rect 1939 1634 1940 1635
rect 1843 1630 1849 1631
rect 1861 1632 1940 1634
rect 1861 1622 1863 1632
rect 1939 1631 1940 1632
rect 1944 1631 1945 1635
rect 2059 1635 2065 1636
rect 2059 1634 2060 1635
rect 1939 1630 1945 1631
rect 1956 1632 2060 1634
rect 1956 1622 1958 1632
rect 2059 1631 2060 1632
rect 2064 1631 2065 1635
rect 2187 1635 2193 1636
rect 2187 1634 2188 1635
rect 2059 1630 2065 1631
rect 2076 1632 2188 1634
rect 2076 1622 2078 1632
rect 2187 1631 2188 1632
rect 2192 1631 2193 1635
rect 2331 1635 2337 1636
rect 2331 1634 2332 1635
rect 2187 1630 2193 1631
rect 2204 1632 2332 1634
rect 2204 1622 2206 1632
rect 2331 1631 2332 1632
rect 2336 1631 2337 1635
rect 2331 1630 2337 1631
rect 2459 1635 2468 1636
rect 2459 1631 2460 1635
rect 2467 1631 2468 1635
rect 2459 1630 2468 1631
rect 1366 1621 1372 1622
rect 1286 1619 1292 1620
rect 1326 1620 1332 1621
rect 1211 1618 1217 1619
rect 1326 1616 1327 1620
rect 1331 1616 1332 1620
rect 1366 1617 1367 1621
rect 1371 1617 1372 1621
rect 1366 1616 1372 1617
rect 1387 1621 1393 1622
rect 1387 1617 1388 1621
rect 1392 1617 1393 1621
rect 1387 1616 1393 1617
rect 1430 1621 1436 1622
rect 1430 1617 1431 1621
rect 1435 1617 1436 1621
rect 1430 1616 1436 1617
rect 1451 1621 1457 1622
rect 1451 1617 1452 1621
rect 1456 1617 1457 1621
rect 1451 1616 1457 1617
rect 1518 1621 1524 1622
rect 1518 1617 1519 1621
rect 1523 1617 1524 1621
rect 1598 1621 1604 1622
rect 1518 1616 1524 1617
rect 1534 1619 1545 1620
rect 1326 1615 1332 1616
rect 1534 1615 1535 1619
rect 1539 1615 1540 1619
rect 1544 1615 1545 1619
rect 1598 1617 1599 1621
rect 1603 1617 1604 1621
rect 1598 1616 1604 1617
rect 1619 1621 1625 1622
rect 1619 1617 1620 1621
rect 1624 1617 1625 1621
rect 1619 1616 1625 1617
rect 1678 1621 1684 1622
rect 1678 1617 1679 1621
rect 1683 1617 1684 1621
rect 1678 1616 1684 1617
rect 1699 1621 1705 1622
rect 1699 1617 1700 1621
rect 1704 1617 1705 1621
rect 1699 1616 1705 1617
rect 1750 1621 1756 1622
rect 1750 1617 1751 1621
rect 1755 1617 1756 1621
rect 1750 1616 1756 1617
rect 1771 1621 1777 1622
rect 1771 1617 1772 1621
rect 1776 1617 1777 1621
rect 1771 1616 1777 1617
rect 1838 1621 1844 1622
rect 1838 1617 1839 1621
rect 1843 1617 1844 1621
rect 1838 1616 1844 1617
rect 1859 1621 1865 1622
rect 1859 1617 1860 1621
rect 1864 1617 1865 1621
rect 1859 1616 1865 1617
rect 1934 1621 1940 1622
rect 1934 1617 1935 1621
rect 1939 1617 1940 1621
rect 1934 1616 1940 1617
rect 1955 1621 1961 1622
rect 1955 1617 1956 1621
rect 1960 1617 1961 1621
rect 1955 1616 1961 1617
rect 2054 1621 2060 1622
rect 2054 1617 2055 1621
rect 2059 1617 2060 1621
rect 2054 1616 2060 1617
rect 2075 1621 2081 1622
rect 2075 1617 2076 1621
rect 2080 1617 2081 1621
rect 2075 1616 2081 1617
rect 2182 1621 2188 1622
rect 2182 1617 2183 1621
rect 2187 1617 2188 1621
rect 2182 1616 2188 1617
rect 2203 1621 2209 1622
rect 2203 1617 2204 1621
rect 2208 1617 2209 1621
rect 2203 1616 2209 1617
rect 2326 1621 2332 1622
rect 2326 1617 2327 1621
rect 2331 1617 2332 1621
rect 2454 1621 2460 1622
rect 2326 1616 2332 1617
rect 2346 1619 2353 1620
rect 1534 1614 1545 1615
rect 2346 1615 2347 1619
rect 2352 1615 2353 1619
rect 2454 1617 2455 1621
rect 2459 1617 2460 1621
rect 2502 1620 2508 1621
rect 2454 1616 2460 1617
rect 2462 1619 2468 1620
rect 2346 1614 2353 1615
rect 2462 1615 2463 1619
rect 2467 1618 2468 1619
rect 2475 1619 2481 1620
rect 2475 1618 2476 1619
rect 2467 1616 2476 1618
rect 2467 1615 2468 1616
rect 2462 1614 2468 1615
rect 2475 1615 2476 1616
rect 2480 1615 2481 1619
rect 2502 1616 2503 1620
rect 2507 1616 2508 1620
rect 2502 1615 2508 1616
rect 2475 1614 2481 1615
rect 860 1612 970 1614
rect 1076 1612 1202 1614
rect 860 1610 862 1612
rect 1076 1610 1078 1612
rect 748 1609 769 1610
rect 748 1608 764 1609
rect 504 1605 505 1608
rect 499 1604 505 1605
rect 526 1607 532 1608
rect 355 1602 364 1603
rect 526 1603 527 1607
rect 531 1606 532 1607
rect 579 1607 585 1608
rect 579 1606 580 1607
rect 531 1604 580 1606
rect 531 1603 532 1604
rect 526 1602 532 1603
rect 579 1603 580 1604
rect 584 1603 585 1607
rect 579 1602 585 1603
rect 667 1607 673 1608
rect 667 1603 668 1607
rect 672 1606 673 1607
rect 672 1604 758 1606
rect 763 1605 764 1608
rect 768 1605 769 1609
rect 763 1604 769 1605
rect 859 1609 865 1610
rect 859 1605 860 1609
rect 864 1605 865 1609
rect 1075 1609 1081 1610
rect 859 1604 865 1605
rect 963 1607 972 1608
rect 672 1603 673 1604
rect 667 1602 673 1603
rect 756 1602 758 1604
rect 870 1603 876 1604
rect 870 1602 871 1603
rect 276 1600 321 1602
rect 756 1600 871 1602
rect 870 1599 871 1600
rect 875 1599 876 1603
rect 963 1603 964 1607
rect 971 1603 972 1607
rect 1075 1605 1076 1609
rect 1080 1605 1081 1609
rect 1075 1604 1081 1605
rect 1195 1607 1201 1608
rect 963 1602 972 1603
rect 1195 1603 1196 1607
rect 1200 1606 1201 1607
rect 1210 1607 1216 1608
rect 1210 1606 1211 1607
rect 1200 1604 1211 1606
rect 1200 1603 1201 1604
rect 1195 1602 1201 1603
rect 1210 1603 1211 1604
rect 1215 1603 1216 1607
rect 1210 1602 1216 1603
rect 1326 1603 1332 1604
rect 870 1598 876 1599
rect 1326 1599 1327 1603
rect 1331 1599 1332 1603
rect 2502 1603 2508 1604
rect 1326 1598 1332 1599
rect 1350 1600 1356 1601
rect 1350 1596 1351 1600
rect 1355 1596 1356 1600
rect 1350 1595 1356 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1502 1600 1508 1601
rect 1502 1596 1503 1600
rect 1507 1596 1508 1600
rect 1502 1595 1508 1596
rect 1582 1600 1588 1601
rect 1582 1596 1583 1600
rect 1587 1596 1588 1600
rect 1582 1595 1588 1596
rect 1662 1600 1668 1601
rect 1662 1596 1663 1600
rect 1667 1596 1668 1600
rect 1662 1595 1668 1596
rect 1734 1600 1740 1601
rect 1734 1596 1735 1600
rect 1739 1596 1740 1600
rect 1734 1595 1740 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1918 1600 1924 1601
rect 1918 1596 1919 1600
rect 1923 1596 1924 1600
rect 1918 1595 1924 1596
rect 2038 1600 2044 1601
rect 2038 1596 2039 1600
rect 2043 1596 2044 1600
rect 2038 1595 2044 1596
rect 2166 1600 2172 1601
rect 2166 1596 2167 1600
rect 2171 1596 2172 1600
rect 2166 1595 2172 1596
rect 2310 1600 2316 1601
rect 2310 1596 2311 1600
rect 2315 1596 2316 1600
rect 2310 1595 2316 1596
rect 2438 1600 2444 1601
rect 2438 1596 2439 1600
rect 2443 1596 2444 1600
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2438 1595 2444 1596
rect 291 1587 300 1588
rect 291 1583 292 1587
rect 299 1583 300 1587
rect 355 1587 361 1588
rect 355 1586 356 1587
rect 291 1582 300 1583
rect 319 1584 356 1586
rect 319 1574 321 1584
rect 355 1583 356 1584
rect 360 1583 361 1587
rect 427 1587 433 1588
rect 427 1586 428 1587
rect 355 1582 361 1583
rect 388 1584 428 1586
rect 388 1578 390 1584
rect 427 1583 428 1584
rect 432 1583 433 1587
rect 427 1582 433 1583
rect 507 1587 513 1588
rect 507 1583 508 1587
rect 512 1583 513 1587
rect 507 1582 513 1583
rect 603 1587 609 1588
rect 603 1583 604 1587
rect 608 1586 609 1587
rect 618 1587 624 1588
rect 618 1586 619 1587
rect 608 1584 619 1586
rect 608 1583 609 1584
rect 603 1582 609 1583
rect 618 1583 619 1584
rect 623 1583 624 1587
rect 707 1587 713 1588
rect 707 1586 708 1587
rect 618 1582 624 1583
rect 629 1584 708 1586
rect 509 1578 511 1582
rect 629 1578 631 1584
rect 707 1583 708 1584
rect 712 1583 713 1587
rect 707 1582 713 1583
rect 806 1587 812 1588
rect 806 1583 807 1587
rect 811 1586 812 1587
rect 819 1587 825 1588
rect 819 1586 820 1587
rect 811 1584 820 1586
rect 811 1583 812 1584
rect 806 1582 812 1583
rect 819 1583 820 1584
rect 824 1583 825 1587
rect 819 1582 825 1583
rect 939 1587 945 1588
rect 939 1583 940 1587
rect 944 1583 945 1587
rect 939 1582 945 1583
rect 990 1587 996 1588
rect 990 1583 991 1587
rect 995 1586 996 1587
rect 1067 1587 1073 1588
rect 1067 1586 1068 1587
rect 995 1584 1068 1586
rect 995 1583 996 1584
rect 990 1582 996 1583
rect 1067 1583 1068 1584
rect 1072 1583 1073 1587
rect 1195 1587 1201 1588
rect 1195 1586 1196 1587
rect 1067 1582 1073 1583
rect 1159 1584 1196 1586
rect 941 1578 943 1582
rect 1159 1578 1161 1584
rect 1195 1583 1196 1584
rect 1200 1583 1201 1587
rect 1195 1582 1201 1583
rect 1350 1584 1356 1585
rect 372 1576 390 1578
rect 444 1576 511 1578
rect 620 1576 631 1578
rect 837 1576 943 1578
rect 1084 1576 1161 1578
rect 1326 1581 1332 1582
rect 1326 1577 1327 1581
rect 1331 1577 1332 1581
rect 1350 1580 1351 1584
rect 1355 1580 1356 1584
rect 1350 1579 1356 1580
rect 1422 1584 1428 1585
rect 1422 1580 1423 1584
rect 1427 1580 1428 1584
rect 1422 1579 1428 1580
rect 1526 1584 1532 1585
rect 1526 1580 1527 1584
rect 1531 1580 1532 1584
rect 1526 1579 1532 1580
rect 1646 1584 1652 1585
rect 1646 1580 1647 1584
rect 1651 1580 1652 1584
rect 1646 1579 1652 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1934 1584 1940 1585
rect 1934 1580 1935 1584
rect 1939 1580 1940 1584
rect 1934 1579 1940 1580
rect 2102 1584 2108 1585
rect 2102 1580 2103 1584
rect 2107 1580 2108 1584
rect 2102 1579 2108 1580
rect 2278 1584 2284 1585
rect 2278 1580 2279 1584
rect 2283 1580 2284 1584
rect 2278 1579 2284 1580
rect 2438 1584 2444 1585
rect 2438 1580 2439 1584
rect 2443 1580 2444 1584
rect 2438 1579 2444 1580
rect 2502 1581 2508 1582
rect 1326 1576 1332 1577
rect 2502 1577 2503 1581
rect 2507 1577 2508 1581
rect 2502 1576 2508 1577
rect 372 1574 374 1576
rect 444 1574 446 1576
rect 620 1574 622 1576
rect 837 1574 839 1576
rect 1084 1574 1086 1576
rect 286 1573 292 1574
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 286 1569 287 1573
rect 291 1569 292 1573
rect 286 1568 292 1569
rect 307 1573 321 1574
rect 307 1569 308 1573
rect 312 1572 321 1573
rect 350 1573 356 1574
rect 312 1569 313 1572
rect 307 1568 313 1569
rect 350 1569 351 1573
rect 355 1569 356 1573
rect 350 1568 356 1569
rect 371 1573 377 1574
rect 371 1569 372 1573
rect 376 1569 377 1573
rect 371 1568 377 1569
rect 422 1573 428 1574
rect 422 1569 423 1573
rect 427 1569 428 1573
rect 422 1568 428 1569
rect 443 1573 449 1574
rect 443 1569 444 1573
rect 448 1569 449 1573
rect 443 1568 449 1569
rect 502 1573 508 1574
rect 502 1569 503 1573
rect 507 1569 508 1573
rect 598 1573 604 1574
rect 502 1568 508 1569
rect 523 1571 532 1572
rect 110 1567 116 1568
rect 523 1567 524 1571
rect 531 1567 532 1571
rect 598 1569 599 1573
rect 603 1569 604 1573
rect 598 1568 604 1569
rect 619 1573 625 1574
rect 619 1569 620 1573
rect 624 1569 625 1573
rect 619 1568 625 1569
rect 702 1573 708 1574
rect 702 1569 703 1573
rect 707 1569 708 1573
rect 814 1573 820 1574
rect 702 1568 708 1569
rect 723 1571 729 1572
rect 523 1566 532 1567
rect 723 1567 724 1571
rect 728 1570 729 1571
rect 742 1571 748 1572
rect 742 1570 743 1571
rect 728 1568 743 1570
rect 728 1567 729 1568
rect 723 1566 729 1567
rect 742 1567 743 1568
rect 747 1567 748 1571
rect 814 1569 815 1573
rect 819 1569 820 1573
rect 814 1568 820 1569
rect 835 1573 841 1574
rect 835 1569 836 1573
rect 840 1569 841 1573
rect 835 1568 841 1569
rect 934 1573 940 1574
rect 934 1569 935 1573
rect 939 1569 940 1573
rect 1062 1573 1068 1574
rect 934 1568 940 1569
rect 954 1571 961 1572
rect 742 1566 748 1567
rect 954 1567 955 1571
rect 960 1567 961 1571
rect 1062 1569 1063 1573
rect 1067 1569 1068 1573
rect 1062 1568 1068 1569
rect 1083 1573 1089 1574
rect 1083 1569 1084 1573
rect 1088 1569 1089 1573
rect 1083 1568 1089 1569
rect 1190 1573 1196 1574
rect 1190 1569 1191 1573
rect 1195 1569 1196 1573
rect 1286 1572 1292 1573
rect 1190 1568 1196 1569
rect 1210 1571 1217 1572
rect 954 1566 961 1567
rect 1210 1567 1211 1571
rect 1216 1567 1217 1571
rect 1286 1568 1287 1572
rect 1291 1568 1292 1572
rect 1286 1567 1292 1568
rect 1210 1566 1217 1567
rect 1326 1564 1332 1565
rect 2502 1564 2508 1565
rect 1326 1560 1327 1564
rect 1331 1560 1332 1564
rect 1326 1559 1332 1560
rect 1366 1563 1372 1564
rect 1366 1559 1367 1563
rect 1371 1559 1372 1563
rect 1366 1558 1372 1559
rect 1374 1563 1380 1564
rect 1374 1559 1375 1563
rect 1379 1562 1380 1563
rect 1387 1563 1393 1564
rect 1387 1562 1388 1563
rect 1379 1560 1388 1562
rect 1379 1559 1380 1560
rect 1374 1558 1380 1559
rect 1387 1559 1388 1560
rect 1392 1559 1393 1563
rect 1387 1558 1393 1559
rect 1438 1563 1444 1564
rect 1438 1559 1439 1563
rect 1443 1559 1444 1563
rect 1459 1563 1465 1564
rect 1459 1562 1460 1563
rect 1438 1558 1444 1559
rect 1448 1560 1460 1562
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 1286 1555 1292 1556
rect 110 1550 116 1551
rect 270 1552 276 1553
rect 270 1548 271 1552
rect 275 1548 276 1552
rect 270 1547 276 1548
rect 334 1552 340 1553
rect 334 1548 335 1552
rect 339 1548 340 1552
rect 334 1547 340 1548
rect 406 1552 412 1553
rect 406 1548 407 1552
rect 411 1548 412 1552
rect 406 1547 412 1548
rect 486 1552 492 1553
rect 486 1548 487 1552
rect 491 1548 492 1552
rect 486 1547 492 1548
rect 582 1552 588 1553
rect 582 1548 583 1552
rect 587 1548 588 1552
rect 582 1547 588 1548
rect 686 1552 692 1553
rect 686 1548 687 1552
rect 691 1548 692 1552
rect 686 1547 692 1548
rect 798 1552 804 1553
rect 798 1548 799 1552
rect 803 1548 804 1552
rect 798 1547 804 1548
rect 918 1552 924 1553
rect 918 1548 919 1552
rect 923 1548 924 1552
rect 918 1547 924 1548
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1174 1552 1180 1553
rect 1174 1548 1175 1552
rect 1179 1548 1180 1552
rect 1286 1551 1287 1555
rect 1291 1551 1292 1555
rect 1448 1554 1450 1560
rect 1459 1559 1460 1560
rect 1464 1559 1465 1563
rect 1459 1558 1465 1559
rect 1542 1563 1548 1564
rect 1542 1559 1543 1563
rect 1547 1559 1548 1563
rect 1542 1558 1548 1559
rect 1563 1563 1569 1564
rect 1563 1559 1564 1563
rect 1568 1559 1569 1563
rect 1563 1558 1569 1559
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1559 1668 1563
rect 1662 1558 1668 1559
rect 1683 1563 1689 1564
rect 1683 1559 1684 1563
rect 1688 1562 1689 1563
rect 1798 1563 1804 1564
rect 1688 1560 1790 1562
rect 1688 1559 1689 1560
rect 1683 1558 1689 1559
rect 1286 1550 1292 1551
rect 1372 1552 1450 1554
rect 1372 1550 1374 1552
rect 1565 1550 1567 1558
rect 1788 1550 1790 1560
rect 1798 1559 1799 1563
rect 1803 1559 1804 1563
rect 1798 1558 1804 1559
rect 1819 1563 1825 1564
rect 1819 1559 1820 1563
rect 1824 1562 1825 1563
rect 1950 1563 1956 1564
rect 1824 1560 1946 1562
rect 1824 1559 1825 1560
rect 1819 1558 1825 1559
rect 1944 1550 1946 1560
rect 1950 1559 1951 1563
rect 1955 1559 1956 1563
rect 1950 1558 1956 1559
rect 1971 1563 1977 1564
rect 1971 1559 1972 1563
rect 1976 1562 1977 1563
rect 2118 1563 2124 1564
rect 1976 1560 2001 1562
rect 1976 1559 1977 1560
rect 1971 1558 1977 1559
rect 1999 1550 2001 1560
rect 2118 1559 2119 1563
rect 2123 1559 2124 1563
rect 2118 1558 2124 1559
rect 2138 1563 2145 1564
rect 2138 1559 2139 1563
rect 2144 1559 2145 1563
rect 2138 1558 2145 1559
rect 2294 1563 2300 1564
rect 2294 1559 2295 1563
rect 2299 1559 2300 1563
rect 2294 1558 2300 1559
rect 2310 1563 2321 1564
rect 2310 1559 2311 1563
rect 2315 1559 2316 1563
rect 2320 1559 2321 1563
rect 2310 1558 2321 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 2470 1563 2481 1564
rect 2470 1559 2471 1563
rect 2475 1559 2476 1563
rect 2480 1559 2481 1563
rect 2502 1560 2503 1564
rect 2507 1560 2508 1564
rect 2502 1559 2508 1560
rect 2470 1558 2481 1559
rect 1174 1547 1180 1548
rect 1371 1549 1377 1550
rect 1371 1545 1372 1549
rect 1376 1545 1377 1549
rect 1565 1549 1673 1550
rect 1565 1548 1668 1549
rect 1371 1544 1377 1545
rect 1443 1547 1449 1548
rect 1443 1543 1444 1547
rect 1448 1546 1449 1547
rect 1534 1547 1540 1548
rect 1534 1546 1535 1547
rect 1448 1544 1535 1546
rect 1448 1543 1449 1544
rect 1443 1542 1449 1543
rect 1534 1543 1535 1544
rect 1539 1543 1540 1547
rect 1534 1542 1540 1543
rect 1547 1547 1553 1548
rect 1547 1543 1548 1547
rect 1552 1546 1553 1547
rect 1552 1544 1663 1546
rect 1667 1545 1668 1548
rect 1672 1545 1673 1549
rect 1788 1549 1809 1550
rect 1788 1548 1804 1549
rect 1667 1544 1673 1545
rect 1803 1545 1804 1548
rect 1808 1545 1809 1549
rect 1944 1549 1961 1550
rect 1944 1548 1956 1549
rect 1803 1544 1809 1545
rect 1955 1545 1956 1548
rect 1960 1545 1961 1549
rect 1999 1549 2129 1550
rect 1999 1548 2124 1549
rect 1955 1544 1961 1545
rect 2123 1545 2124 1548
rect 2128 1545 2129 1549
rect 2123 1544 2129 1545
rect 2270 1547 2276 1548
rect 1552 1543 1553 1544
rect 1547 1542 1553 1543
rect 1661 1542 1663 1544
rect 1874 1543 1880 1544
rect 1874 1542 1875 1543
rect 1661 1540 1875 1542
rect 1874 1539 1875 1540
rect 1879 1539 1880 1543
rect 2270 1543 2271 1547
rect 2275 1546 2276 1547
rect 2299 1547 2305 1548
rect 2299 1546 2300 1547
rect 2275 1544 2300 1546
rect 2275 1543 2276 1544
rect 2270 1542 2276 1543
rect 2299 1543 2300 1544
rect 2304 1543 2305 1547
rect 2459 1547 2468 1548
rect 2299 1542 2305 1543
rect 2310 1543 2316 1544
rect 1874 1538 1880 1539
rect 2310 1539 2311 1543
rect 2315 1539 2316 1543
rect 2459 1543 2460 1547
rect 2467 1543 2468 1547
rect 2459 1542 2468 1543
rect 2310 1538 2316 1539
rect 1999 1536 2314 1538
rect 470 1532 476 1533
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 470 1528 471 1532
rect 475 1528 476 1532
rect 470 1527 476 1528
rect 550 1532 556 1533
rect 550 1528 551 1532
rect 555 1528 556 1532
rect 550 1527 556 1528
rect 638 1532 644 1533
rect 638 1528 639 1532
rect 643 1528 644 1532
rect 638 1527 644 1528
rect 734 1532 740 1533
rect 734 1528 735 1532
rect 739 1528 740 1532
rect 734 1527 740 1528
rect 838 1532 844 1533
rect 838 1528 839 1532
rect 843 1528 844 1532
rect 838 1527 844 1528
rect 950 1532 956 1533
rect 950 1528 951 1532
rect 955 1528 956 1532
rect 950 1527 956 1528
rect 1062 1532 1068 1533
rect 1062 1528 1063 1532
rect 1067 1528 1068 1532
rect 1062 1527 1068 1528
rect 1174 1532 1180 1533
rect 1174 1528 1175 1532
rect 1179 1528 1180 1532
rect 1999 1530 2001 1536
rect 2362 1535 2368 1536
rect 2362 1534 2363 1535
rect 2156 1532 2363 1534
rect 2156 1530 2158 1532
rect 2362 1531 2363 1532
rect 2367 1531 2368 1535
rect 2362 1530 2368 1531
rect 1174 1527 1180 1528
rect 1286 1529 1292 1530
rect 110 1524 116 1525
rect 1286 1525 1287 1529
rect 1291 1525 1292 1529
rect 1963 1529 2001 1530
rect 1286 1524 1292 1525
rect 1371 1527 1380 1528
rect 1371 1523 1372 1527
rect 1379 1523 1380 1527
rect 1443 1527 1449 1528
rect 1443 1526 1444 1527
rect 1371 1522 1380 1523
rect 1389 1524 1444 1526
rect 1389 1514 1391 1524
rect 1443 1523 1444 1524
rect 1448 1523 1449 1527
rect 1547 1527 1553 1528
rect 1547 1526 1548 1527
rect 1443 1522 1449 1523
rect 1460 1524 1548 1526
rect 1460 1514 1462 1524
rect 1547 1523 1548 1524
rect 1552 1523 1553 1527
rect 1547 1522 1553 1523
rect 1651 1527 1660 1528
rect 1651 1523 1652 1527
rect 1659 1523 1660 1527
rect 1651 1522 1660 1523
rect 1755 1527 1761 1528
rect 1755 1523 1756 1527
rect 1760 1523 1761 1527
rect 1755 1522 1761 1523
rect 1859 1527 1865 1528
rect 1859 1523 1860 1527
rect 1864 1523 1865 1527
rect 1963 1525 1964 1529
rect 1968 1528 2001 1529
rect 2155 1529 2161 1530
rect 1968 1525 1969 1528
rect 2059 1527 2065 1528
rect 2059 1526 2060 1527
rect 1963 1524 1969 1525
rect 1999 1524 2060 1526
rect 1859 1522 1865 1523
rect 1470 1519 1476 1520
rect 1470 1515 1471 1519
rect 1475 1518 1476 1519
rect 1757 1518 1759 1522
rect 1861 1518 1863 1522
rect 1475 1516 1567 1518
rect 1475 1515 1476 1516
rect 1470 1514 1476 1515
rect 1565 1514 1567 1516
rect 1668 1516 1759 1518
rect 1772 1516 1863 1518
rect 1668 1514 1670 1516
rect 1772 1514 1774 1516
rect 1999 1514 2001 1524
rect 2059 1523 2060 1524
rect 2064 1523 2065 1527
rect 2155 1525 2156 1529
rect 2160 1525 2161 1529
rect 2251 1527 2257 1528
rect 2251 1526 2252 1527
rect 2155 1524 2161 1525
rect 2173 1524 2252 1526
rect 2059 1522 2065 1523
rect 2173 1514 2175 1524
rect 2251 1523 2252 1524
rect 2256 1523 2257 1527
rect 2251 1522 2257 1523
rect 2347 1527 2356 1528
rect 2347 1523 2348 1527
rect 2355 1523 2356 1527
rect 2347 1522 2356 1523
rect 2443 1527 2449 1528
rect 2443 1523 2444 1527
rect 2448 1526 2449 1527
rect 2470 1527 2476 1528
rect 2470 1526 2471 1527
rect 2448 1524 2471 1526
rect 2448 1523 2449 1524
rect 2443 1522 2449 1523
rect 2470 1523 2471 1524
rect 2475 1523 2476 1527
rect 2470 1522 2476 1523
rect 1366 1513 1372 1514
rect 110 1512 116 1513
rect 1286 1512 1292 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 486 1511 492 1512
rect 486 1507 487 1511
rect 491 1507 492 1511
rect 486 1506 492 1507
rect 507 1511 513 1512
rect 507 1507 508 1511
rect 512 1507 513 1511
rect 507 1506 513 1507
rect 566 1511 572 1512
rect 566 1507 567 1511
rect 571 1507 572 1511
rect 566 1506 572 1507
rect 587 1511 593 1512
rect 587 1507 588 1511
rect 592 1510 593 1511
rect 654 1511 660 1512
rect 592 1508 646 1510
rect 592 1507 593 1508
rect 587 1506 593 1507
rect 509 1498 511 1506
rect 644 1498 646 1508
rect 654 1507 655 1511
rect 659 1507 660 1511
rect 654 1506 660 1507
rect 662 1511 668 1512
rect 662 1507 663 1511
rect 667 1510 668 1511
rect 675 1511 681 1512
rect 675 1510 676 1511
rect 667 1508 676 1510
rect 667 1507 668 1508
rect 662 1506 668 1507
rect 675 1507 676 1508
rect 680 1507 681 1511
rect 675 1506 681 1507
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 771 1511 777 1512
rect 771 1507 772 1511
rect 776 1510 777 1511
rect 854 1511 860 1512
rect 776 1508 850 1510
rect 776 1507 777 1508
rect 771 1506 777 1507
rect 848 1498 850 1508
rect 854 1507 855 1511
rect 859 1507 860 1511
rect 854 1506 860 1507
rect 870 1511 881 1512
rect 870 1507 871 1511
rect 875 1507 876 1511
rect 880 1507 881 1511
rect 870 1506 881 1507
rect 966 1511 972 1512
rect 966 1507 967 1511
rect 971 1507 972 1511
rect 966 1506 972 1507
rect 987 1511 996 1512
rect 987 1507 988 1511
rect 995 1507 996 1511
rect 987 1506 996 1507
rect 1078 1511 1084 1512
rect 1078 1507 1079 1511
rect 1083 1507 1084 1511
rect 1078 1506 1084 1507
rect 1094 1511 1105 1512
rect 1094 1507 1095 1511
rect 1099 1507 1100 1511
rect 1104 1507 1105 1511
rect 1094 1506 1105 1507
rect 1190 1511 1196 1512
rect 1190 1507 1191 1511
rect 1195 1507 1196 1511
rect 1211 1511 1217 1512
rect 1211 1510 1212 1511
rect 1190 1506 1196 1507
rect 1200 1508 1212 1510
rect 1200 1502 1202 1508
rect 1211 1507 1212 1508
rect 1216 1507 1217 1511
rect 1286 1508 1287 1512
rect 1291 1508 1292 1512
rect 1286 1507 1292 1508
rect 1326 1512 1332 1513
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1366 1509 1367 1513
rect 1371 1509 1372 1513
rect 1366 1508 1372 1509
rect 1387 1513 1393 1514
rect 1387 1509 1388 1513
rect 1392 1509 1393 1513
rect 1387 1508 1393 1509
rect 1438 1513 1444 1514
rect 1438 1509 1439 1513
rect 1443 1509 1444 1513
rect 1438 1508 1444 1509
rect 1459 1513 1465 1514
rect 1459 1509 1460 1513
rect 1464 1509 1465 1513
rect 1459 1508 1465 1509
rect 1542 1513 1548 1514
rect 1542 1509 1543 1513
rect 1547 1509 1548 1513
rect 1542 1508 1548 1509
rect 1563 1513 1569 1514
rect 1563 1509 1564 1513
rect 1568 1509 1569 1513
rect 1563 1508 1569 1509
rect 1646 1513 1652 1514
rect 1646 1509 1647 1513
rect 1651 1509 1652 1513
rect 1646 1508 1652 1509
rect 1667 1513 1673 1514
rect 1667 1509 1668 1513
rect 1672 1509 1673 1513
rect 1667 1508 1673 1509
rect 1750 1513 1756 1514
rect 1750 1509 1751 1513
rect 1755 1509 1756 1513
rect 1750 1508 1756 1509
rect 1771 1513 1777 1514
rect 1771 1509 1772 1513
rect 1776 1509 1777 1513
rect 1771 1508 1777 1509
rect 1854 1513 1860 1514
rect 1854 1509 1855 1513
rect 1859 1509 1860 1513
rect 1958 1513 1964 1514
rect 1854 1508 1860 1509
rect 1874 1511 1881 1512
rect 1326 1507 1332 1508
rect 1874 1507 1875 1511
rect 1880 1507 1881 1511
rect 1958 1509 1959 1513
rect 1963 1509 1964 1513
rect 1958 1508 1964 1509
rect 1979 1513 2001 1514
rect 1979 1509 1980 1513
rect 1984 1512 2001 1513
rect 2054 1513 2060 1514
rect 1984 1509 1985 1512
rect 1979 1508 1985 1509
rect 2054 1509 2055 1513
rect 2059 1509 2060 1513
rect 2150 1513 2156 1514
rect 2054 1508 2060 1509
rect 2075 1511 2081 1512
rect 1211 1506 1217 1507
rect 1874 1506 1881 1507
rect 2075 1507 2076 1511
rect 2080 1510 2081 1511
rect 2142 1511 2148 1512
rect 2142 1510 2143 1511
rect 2080 1508 2143 1510
rect 2080 1507 2081 1508
rect 2075 1506 2081 1507
rect 2142 1507 2143 1508
rect 2147 1507 2148 1511
rect 2150 1509 2151 1513
rect 2155 1509 2156 1513
rect 2150 1508 2156 1509
rect 2171 1513 2177 1514
rect 2171 1509 2172 1513
rect 2176 1509 2177 1513
rect 2171 1508 2177 1509
rect 2246 1513 2252 1514
rect 2246 1509 2247 1513
rect 2251 1509 2252 1513
rect 2342 1513 2348 1514
rect 2246 1508 2252 1509
rect 2267 1511 2276 1512
rect 2142 1506 2148 1507
rect 2267 1507 2268 1511
rect 2275 1507 2276 1511
rect 2342 1509 2343 1513
rect 2347 1509 2348 1513
rect 2438 1513 2444 1514
rect 2342 1508 2348 1509
rect 2362 1511 2369 1512
rect 2267 1506 2276 1507
rect 2362 1507 2363 1511
rect 2368 1507 2369 1511
rect 2438 1509 2439 1513
rect 2443 1509 2444 1513
rect 2502 1512 2508 1513
rect 2438 1508 2444 1509
rect 2459 1511 2468 1512
rect 2362 1506 2369 1507
rect 2459 1507 2460 1511
rect 2467 1507 2468 1511
rect 2502 1508 2503 1512
rect 2507 1508 2508 1512
rect 2502 1507 2508 1508
rect 2459 1506 2468 1507
rect 1084 1500 1202 1502
rect 1084 1498 1086 1500
rect 509 1497 577 1498
rect 509 1496 572 1497
rect 491 1495 497 1496
rect 491 1491 492 1495
rect 496 1494 497 1495
rect 496 1492 566 1494
rect 571 1493 572 1496
rect 576 1493 577 1497
rect 644 1497 665 1498
rect 644 1496 660 1497
rect 571 1492 577 1493
rect 659 1493 660 1496
rect 664 1493 665 1497
rect 848 1497 865 1498
rect 848 1496 860 1497
rect 659 1492 665 1493
rect 742 1495 748 1496
rect 496 1491 497 1492
rect 491 1490 497 1491
rect 564 1486 566 1492
rect 742 1491 743 1495
rect 747 1494 748 1495
rect 755 1495 761 1496
rect 755 1494 756 1495
rect 747 1492 756 1494
rect 747 1491 748 1492
rect 742 1490 748 1491
rect 755 1491 756 1492
rect 760 1491 761 1495
rect 859 1493 860 1496
rect 864 1493 865 1497
rect 1083 1497 1089 1498
rect 859 1492 865 1493
rect 971 1495 977 1496
rect 755 1490 761 1491
rect 870 1491 876 1492
rect 870 1487 871 1491
rect 875 1487 876 1491
rect 971 1491 972 1495
rect 976 1494 977 1495
rect 976 1492 1039 1494
rect 1083 1493 1084 1497
rect 1088 1493 1089 1497
rect 1083 1492 1089 1493
rect 1195 1495 1204 1496
rect 976 1491 977 1492
rect 971 1490 977 1491
rect 1037 1490 1039 1492
rect 1094 1491 1100 1492
rect 1094 1490 1095 1491
rect 1037 1488 1095 1490
rect 870 1486 876 1487
rect 1094 1487 1095 1488
rect 1099 1487 1100 1491
rect 1195 1491 1196 1495
rect 1203 1491 1204 1495
rect 1195 1490 1204 1491
rect 1326 1495 1332 1496
rect 1326 1491 1327 1495
rect 1331 1491 1332 1495
rect 2502 1495 2508 1496
rect 1326 1490 1332 1491
rect 1350 1492 1356 1493
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1422 1492 1428 1493
rect 1422 1488 1423 1492
rect 1427 1488 1428 1492
rect 1422 1487 1428 1488
rect 1526 1492 1532 1493
rect 1526 1488 1527 1492
rect 1531 1488 1532 1492
rect 1526 1487 1532 1488
rect 1630 1492 1636 1493
rect 1630 1488 1631 1492
rect 1635 1488 1636 1492
rect 1630 1487 1636 1488
rect 1734 1492 1740 1493
rect 1734 1488 1735 1492
rect 1739 1488 1740 1492
rect 1734 1487 1740 1488
rect 1838 1492 1844 1493
rect 1838 1488 1839 1492
rect 1843 1488 1844 1492
rect 1838 1487 1844 1488
rect 1942 1492 1948 1493
rect 1942 1488 1943 1492
rect 1947 1488 1948 1492
rect 1942 1487 1948 1488
rect 2038 1492 2044 1493
rect 2038 1488 2039 1492
rect 2043 1488 2044 1492
rect 2038 1487 2044 1488
rect 2134 1492 2140 1493
rect 2134 1488 2135 1492
rect 2139 1488 2140 1492
rect 2134 1487 2140 1488
rect 2230 1492 2236 1493
rect 2230 1488 2231 1492
rect 2235 1488 2236 1492
rect 2230 1487 2236 1488
rect 2326 1492 2332 1493
rect 2326 1488 2327 1492
rect 2331 1488 2332 1492
rect 2326 1487 2332 1488
rect 2422 1492 2428 1493
rect 2422 1488 2423 1492
rect 2427 1488 2428 1492
rect 2502 1491 2503 1495
rect 2507 1491 2508 1495
rect 2502 1490 2508 1491
rect 2422 1487 2428 1488
rect 1094 1486 1100 1487
rect 564 1484 874 1486
rect 1122 1483 1128 1484
rect 1122 1482 1123 1483
rect 380 1480 774 1482
rect 860 1480 1123 1482
rect 380 1478 382 1480
rect 770 1479 776 1480
rect 379 1477 385 1478
rect 379 1473 380 1477
rect 384 1473 385 1477
rect 467 1475 473 1476
rect 467 1474 468 1475
rect 379 1472 385 1473
rect 396 1472 468 1474
rect 396 1462 398 1472
rect 467 1471 468 1472
rect 472 1471 473 1475
rect 563 1475 569 1476
rect 563 1474 564 1475
rect 467 1470 473 1471
rect 484 1472 564 1474
rect 484 1462 486 1472
rect 563 1471 564 1472
rect 568 1471 569 1475
rect 563 1470 569 1471
rect 659 1475 668 1476
rect 659 1471 660 1475
rect 667 1471 668 1475
rect 755 1475 761 1476
rect 755 1474 756 1475
rect 659 1470 668 1471
rect 676 1472 756 1474
rect 676 1462 678 1472
rect 755 1471 756 1472
rect 760 1471 761 1475
rect 770 1475 771 1479
rect 775 1475 776 1479
rect 860 1478 862 1480
rect 1122 1479 1123 1480
rect 1127 1479 1128 1483
rect 1122 1478 1128 1479
rect 770 1474 776 1475
rect 859 1477 865 1478
rect 859 1473 860 1477
rect 864 1473 865 1477
rect 1350 1476 1356 1477
rect 859 1472 865 1473
rect 963 1475 969 1476
rect 755 1470 761 1471
rect 963 1471 964 1475
rect 968 1471 969 1475
rect 1067 1475 1073 1476
rect 1067 1474 1068 1475
rect 963 1470 969 1471
rect 988 1472 1068 1474
rect 965 1466 967 1470
rect 988 1466 990 1472
rect 1067 1471 1068 1472
rect 1072 1471 1073 1475
rect 1171 1475 1177 1476
rect 1171 1474 1172 1475
rect 1067 1470 1073 1471
rect 1159 1472 1172 1474
rect 1159 1466 1161 1472
rect 1171 1471 1172 1472
rect 1176 1471 1177 1475
rect 1171 1470 1177 1471
rect 1326 1473 1332 1474
rect 1326 1469 1327 1473
rect 1331 1469 1332 1473
rect 1350 1472 1351 1476
rect 1355 1472 1356 1476
rect 1350 1471 1356 1472
rect 1422 1476 1428 1477
rect 1422 1472 1423 1476
rect 1427 1472 1428 1476
rect 1422 1471 1428 1472
rect 1518 1476 1524 1477
rect 1518 1472 1519 1476
rect 1523 1472 1524 1476
rect 1518 1471 1524 1472
rect 1614 1476 1620 1477
rect 1614 1472 1615 1476
rect 1619 1472 1620 1476
rect 1614 1471 1620 1472
rect 1710 1476 1716 1477
rect 1710 1472 1711 1476
rect 1715 1472 1716 1476
rect 1710 1471 1716 1472
rect 1814 1476 1820 1477
rect 1814 1472 1815 1476
rect 1819 1472 1820 1476
rect 1814 1471 1820 1472
rect 1926 1476 1932 1477
rect 1926 1472 1927 1476
rect 1931 1472 1932 1476
rect 1926 1471 1932 1472
rect 2046 1476 2052 1477
rect 2046 1472 2047 1476
rect 2051 1472 2052 1476
rect 2046 1471 2052 1472
rect 2174 1476 2180 1477
rect 2174 1472 2175 1476
rect 2179 1472 2180 1476
rect 2174 1471 2180 1472
rect 2302 1476 2308 1477
rect 2302 1472 2303 1476
rect 2307 1472 2308 1476
rect 2302 1471 2308 1472
rect 2438 1476 2444 1477
rect 2438 1472 2439 1476
rect 2443 1472 2444 1476
rect 2438 1471 2444 1472
rect 2502 1473 2508 1474
rect 1326 1468 1332 1469
rect 2502 1469 2503 1473
rect 2507 1469 2508 1473
rect 2502 1468 2508 1469
rect 876 1464 967 1466
rect 980 1464 990 1466
rect 1084 1464 1161 1466
rect 876 1462 878 1464
rect 980 1462 982 1464
rect 1084 1462 1086 1464
rect 374 1461 380 1462
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 374 1457 375 1461
rect 379 1457 380 1461
rect 374 1456 380 1457
rect 395 1461 401 1462
rect 395 1457 396 1461
rect 400 1457 401 1461
rect 395 1456 401 1457
rect 462 1461 468 1462
rect 462 1457 463 1461
rect 467 1457 468 1461
rect 462 1456 468 1457
rect 483 1461 489 1462
rect 483 1457 484 1461
rect 488 1457 489 1461
rect 483 1456 489 1457
rect 558 1461 564 1462
rect 558 1457 559 1461
rect 563 1457 564 1461
rect 654 1461 660 1462
rect 558 1456 564 1457
rect 579 1459 585 1460
rect 110 1455 116 1456
rect 579 1455 580 1459
rect 584 1458 585 1459
rect 622 1459 628 1460
rect 622 1458 623 1459
rect 584 1456 623 1458
rect 584 1455 585 1456
rect 579 1454 585 1455
rect 622 1455 623 1456
rect 627 1455 628 1459
rect 654 1457 655 1461
rect 659 1457 660 1461
rect 654 1456 660 1457
rect 675 1461 681 1462
rect 675 1457 676 1461
rect 680 1457 681 1461
rect 675 1456 681 1457
rect 750 1461 756 1462
rect 750 1457 751 1461
rect 755 1457 756 1461
rect 854 1461 860 1462
rect 750 1456 756 1457
rect 770 1459 777 1460
rect 622 1454 628 1455
rect 770 1455 771 1459
rect 776 1455 777 1459
rect 854 1457 855 1461
rect 859 1457 860 1461
rect 854 1456 860 1457
rect 875 1461 881 1462
rect 875 1457 876 1461
rect 880 1457 881 1461
rect 875 1456 881 1457
rect 958 1461 964 1462
rect 958 1457 959 1461
rect 963 1457 964 1461
rect 958 1456 964 1457
rect 979 1461 985 1462
rect 979 1457 980 1461
rect 984 1457 985 1461
rect 979 1456 985 1457
rect 1062 1461 1068 1462
rect 1062 1457 1063 1461
rect 1067 1457 1068 1461
rect 1062 1456 1068 1457
rect 1083 1461 1089 1462
rect 1083 1457 1084 1461
rect 1088 1457 1089 1461
rect 1083 1456 1089 1457
rect 1166 1461 1172 1462
rect 1166 1457 1167 1461
rect 1171 1457 1172 1461
rect 1286 1460 1292 1461
rect 1166 1456 1172 1457
rect 1187 1459 1193 1460
rect 770 1454 777 1455
rect 1187 1455 1188 1459
rect 1192 1458 1193 1459
rect 1198 1459 1204 1460
rect 1198 1458 1199 1459
rect 1192 1456 1199 1458
rect 1192 1455 1193 1456
rect 1187 1454 1193 1455
rect 1198 1455 1199 1456
rect 1203 1455 1204 1459
rect 1286 1456 1287 1460
rect 1291 1456 1292 1460
rect 1286 1455 1292 1456
rect 1326 1456 1332 1457
rect 2502 1456 2508 1457
rect 1198 1454 1204 1455
rect 1326 1452 1327 1456
rect 1331 1452 1332 1456
rect 1326 1451 1332 1452
rect 1366 1455 1372 1456
rect 1366 1451 1367 1455
rect 1371 1451 1372 1455
rect 1366 1450 1372 1451
rect 1387 1455 1393 1456
rect 1387 1451 1388 1455
rect 1392 1454 1393 1455
rect 1414 1455 1420 1456
rect 1414 1454 1415 1455
rect 1392 1452 1415 1454
rect 1392 1451 1393 1452
rect 1387 1450 1393 1451
rect 1414 1451 1415 1452
rect 1419 1451 1420 1455
rect 1414 1450 1420 1451
rect 1438 1455 1444 1456
rect 1438 1451 1439 1455
rect 1443 1451 1444 1455
rect 1459 1455 1465 1456
rect 1459 1454 1460 1455
rect 1438 1450 1444 1451
rect 1448 1452 1460 1454
rect 1448 1446 1450 1452
rect 1459 1451 1460 1452
rect 1464 1451 1465 1455
rect 1459 1450 1465 1451
rect 1534 1455 1540 1456
rect 1534 1451 1535 1455
rect 1539 1451 1540 1455
rect 1534 1450 1540 1451
rect 1555 1455 1561 1456
rect 1555 1451 1556 1455
rect 1560 1451 1561 1455
rect 1555 1450 1561 1451
rect 1630 1455 1636 1456
rect 1630 1451 1631 1455
rect 1635 1451 1636 1455
rect 1630 1450 1636 1451
rect 1651 1455 1660 1456
rect 1651 1451 1652 1455
rect 1659 1451 1660 1455
rect 1651 1450 1660 1451
rect 1726 1455 1732 1456
rect 1726 1451 1727 1455
rect 1731 1451 1732 1455
rect 1747 1455 1753 1456
rect 1747 1454 1748 1455
rect 1726 1450 1732 1451
rect 1736 1452 1748 1454
rect 1372 1444 1450 1446
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 1286 1443 1292 1444
rect 110 1438 116 1439
rect 358 1440 364 1441
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 446 1440 452 1441
rect 446 1436 447 1440
rect 451 1436 452 1440
rect 446 1435 452 1436
rect 542 1440 548 1441
rect 542 1436 543 1440
rect 547 1436 548 1440
rect 542 1435 548 1436
rect 638 1440 644 1441
rect 638 1436 639 1440
rect 643 1436 644 1440
rect 638 1435 644 1436
rect 734 1440 740 1441
rect 734 1436 735 1440
rect 739 1436 740 1440
rect 734 1435 740 1436
rect 838 1440 844 1441
rect 838 1436 839 1440
rect 843 1436 844 1440
rect 838 1435 844 1436
rect 942 1440 948 1441
rect 942 1436 943 1440
rect 947 1436 948 1440
rect 942 1435 948 1436
rect 1046 1440 1052 1441
rect 1046 1436 1047 1440
rect 1051 1436 1052 1440
rect 1046 1435 1052 1436
rect 1150 1440 1156 1441
rect 1150 1436 1151 1440
rect 1155 1436 1156 1440
rect 1286 1439 1287 1443
rect 1291 1439 1292 1443
rect 1372 1442 1374 1444
rect 1557 1442 1559 1450
rect 1736 1446 1738 1452
rect 1747 1451 1748 1452
rect 1752 1451 1753 1455
rect 1747 1450 1753 1451
rect 1830 1455 1836 1456
rect 1830 1451 1831 1455
rect 1835 1451 1836 1455
rect 1830 1450 1836 1451
rect 1838 1455 1844 1456
rect 1838 1451 1839 1455
rect 1843 1454 1844 1455
rect 1851 1455 1857 1456
rect 1851 1454 1852 1455
rect 1843 1452 1852 1454
rect 1843 1451 1844 1452
rect 1838 1450 1844 1451
rect 1851 1451 1852 1452
rect 1856 1451 1857 1455
rect 1851 1450 1857 1451
rect 1942 1455 1948 1456
rect 1942 1451 1943 1455
rect 1947 1451 1948 1455
rect 1942 1450 1948 1451
rect 1958 1455 1969 1456
rect 1958 1451 1959 1455
rect 1963 1451 1964 1455
rect 1968 1451 1969 1455
rect 1958 1450 1969 1451
rect 2062 1455 2068 1456
rect 2062 1451 2063 1455
rect 2067 1451 2068 1455
rect 2083 1455 2089 1456
rect 2083 1454 2084 1455
rect 2062 1450 2068 1451
rect 2072 1452 2084 1454
rect 2072 1446 2074 1452
rect 2083 1451 2084 1452
rect 2088 1451 2089 1455
rect 2083 1450 2089 1451
rect 2190 1455 2196 1456
rect 2190 1451 2191 1455
rect 2195 1451 2196 1455
rect 2211 1455 2217 1456
rect 2211 1454 2212 1455
rect 2190 1450 2196 1451
rect 2200 1452 2212 1454
rect 2200 1446 2202 1452
rect 2211 1451 2212 1452
rect 2216 1451 2217 1455
rect 2211 1450 2217 1451
rect 2318 1455 2324 1456
rect 2318 1451 2319 1455
rect 2323 1451 2324 1455
rect 2318 1450 2324 1451
rect 2339 1455 2345 1456
rect 2339 1451 2340 1455
rect 2344 1454 2345 1455
rect 2350 1455 2356 1456
rect 2350 1454 2351 1455
rect 2344 1452 2351 1454
rect 2344 1451 2345 1452
rect 2339 1450 2345 1451
rect 2350 1451 2351 1452
rect 2355 1451 2356 1455
rect 2350 1450 2356 1451
rect 2454 1455 2460 1456
rect 2454 1451 2455 1455
rect 2459 1451 2460 1455
rect 2454 1450 2460 1451
rect 2470 1455 2481 1456
rect 2470 1451 2471 1455
rect 2475 1451 2476 1455
rect 2480 1451 2481 1455
rect 2502 1452 2503 1456
rect 2507 1452 2508 1456
rect 2502 1451 2508 1452
rect 2470 1450 2481 1451
rect 1644 1444 1738 1446
rect 1948 1444 2074 1446
rect 2076 1444 2202 1446
rect 1286 1438 1292 1439
rect 1371 1441 1377 1442
rect 1371 1437 1372 1441
rect 1376 1437 1377 1441
rect 1557 1441 1641 1442
rect 1557 1440 1636 1441
rect 1371 1436 1377 1437
rect 1443 1439 1449 1440
rect 1150 1435 1156 1436
rect 1443 1435 1444 1439
rect 1448 1438 1449 1439
rect 1470 1439 1476 1440
rect 1470 1438 1471 1439
rect 1448 1436 1471 1438
rect 1448 1435 1449 1436
rect 1443 1434 1449 1435
rect 1470 1435 1471 1436
rect 1475 1435 1476 1439
rect 1470 1434 1476 1435
rect 1539 1439 1545 1440
rect 1539 1435 1540 1439
rect 1544 1438 1545 1439
rect 1544 1436 1559 1438
rect 1635 1437 1636 1440
rect 1640 1437 1641 1441
rect 1635 1436 1641 1437
rect 1544 1435 1545 1436
rect 1539 1434 1545 1435
rect 1557 1434 1559 1436
rect 1644 1434 1646 1444
rect 1948 1442 1950 1444
rect 2076 1442 2078 1444
rect 1947 1441 1953 1442
rect 1702 1439 1708 1440
rect 1702 1435 1703 1439
rect 1707 1438 1708 1439
rect 1731 1439 1737 1440
rect 1731 1438 1732 1439
rect 1707 1436 1732 1438
rect 1707 1435 1708 1436
rect 1702 1434 1708 1435
rect 1731 1435 1732 1436
rect 1736 1435 1737 1439
rect 1731 1434 1737 1435
rect 1835 1439 1841 1440
rect 1835 1435 1836 1439
rect 1840 1438 1841 1439
rect 1840 1436 1902 1438
rect 1947 1437 1948 1441
rect 1952 1437 1953 1441
rect 1947 1436 1953 1437
rect 2067 1441 2078 1442
rect 2067 1437 2068 1441
rect 2072 1440 2078 1441
rect 2072 1437 2073 1440
rect 2067 1436 2073 1437
rect 2142 1439 2148 1440
rect 1840 1435 1841 1436
rect 1835 1434 1841 1435
rect 1900 1434 1902 1436
rect 1958 1435 1964 1436
rect 1958 1434 1959 1435
rect 1557 1432 1646 1434
rect 1900 1432 1959 1434
rect 1958 1431 1959 1432
rect 1963 1431 1964 1435
rect 2142 1435 2143 1439
rect 2147 1438 2148 1439
rect 2195 1439 2201 1440
rect 2195 1438 2196 1439
rect 2147 1436 2196 1438
rect 2147 1435 2148 1436
rect 2142 1434 2148 1435
rect 2195 1435 2196 1436
rect 2200 1435 2201 1439
rect 2195 1434 2201 1435
rect 2254 1439 2260 1440
rect 2254 1435 2255 1439
rect 2259 1438 2260 1439
rect 2323 1439 2329 1440
rect 2323 1438 2324 1439
rect 2259 1436 2324 1438
rect 2259 1435 2260 1436
rect 2254 1434 2260 1435
rect 2323 1435 2324 1436
rect 2328 1435 2329 1439
rect 2323 1434 2329 1435
rect 2459 1439 2468 1440
rect 2459 1435 2460 1439
rect 2467 1435 2468 1439
rect 2459 1434 2468 1435
rect 1958 1430 1964 1431
rect 230 1428 236 1429
rect 110 1425 116 1426
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 230 1424 231 1428
rect 235 1424 236 1428
rect 230 1423 236 1424
rect 318 1428 324 1429
rect 318 1424 319 1428
rect 323 1424 324 1428
rect 318 1423 324 1424
rect 414 1428 420 1429
rect 414 1424 415 1428
rect 419 1424 420 1428
rect 414 1423 420 1424
rect 510 1428 516 1429
rect 510 1424 511 1428
rect 515 1424 516 1428
rect 510 1423 516 1424
rect 614 1428 620 1429
rect 614 1424 615 1428
rect 619 1424 620 1428
rect 614 1423 620 1424
rect 710 1428 716 1429
rect 710 1424 711 1428
rect 715 1424 716 1428
rect 710 1423 716 1424
rect 806 1428 812 1429
rect 806 1424 807 1428
rect 811 1424 812 1428
rect 806 1423 812 1424
rect 894 1428 900 1429
rect 894 1424 895 1428
rect 899 1424 900 1428
rect 894 1423 900 1424
rect 990 1428 996 1429
rect 990 1424 991 1428
rect 995 1424 996 1428
rect 990 1423 996 1424
rect 1086 1428 1092 1429
rect 1086 1424 1087 1428
rect 1091 1424 1092 1428
rect 1086 1423 1092 1424
rect 1286 1425 1292 1426
rect 110 1420 116 1421
rect 1286 1421 1287 1425
rect 1291 1421 1292 1425
rect 1602 1423 1608 1424
rect 1602 1422 1603 1423
rect 1286 1420 1292 1421
rect 1508 1420 1603 1422
rect 1508 1418 1510 1420
rect 1602 1419 1603 1420
rect 1607 1419 1608 1423
rect 1838 1423 1844 1424
rect 1838 1422 1839 1423
rect 1602 1418 1608 1419
rect 1780 1420 1839 1422
rect 1780 1418 1782 1420
rect 1838 1419 1839 1420
rect 1843 1419 1844 1423
rect 1838 1418 1844 1419
rect 1507 1417 1513 1418
rect 1371 1415 1377 1416
rect 1371 1411 1372 1415
rect 1376 1414 1377 1415
rect 1414 1415 1420 1416
rect 1376 1412 1410 1414
rect 1376 1411 1377 1412
rect 1371 1410 1377 1411
rect 110 1408 116 1409
rect 1286 1408 1292 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 246 1407 252 1408
rect 246 1403 247 1407
rect 251 1403 252 1407
rect 246 1402 252 1403
rect 267 1407 273 1408
rect 267 1403 268 1407
rect 272 1406 273 1407
rect 334 1407 340 1408
rect 272 1404 321 1406
rect 272 1403 273 1404
rect 267 1402 273 1403
rect 319 1394 321 1404
rect 334 1403 335 1407
rect 339 1403 340 1407
rect 334 1402 340 1403
rect 355 1407 361 1408
rect 355 1403 356 1407
rect 360 1406 361 1407
rect 430 1407 436 1408
rect 360 1404 426 1406
rect 360 1403 361 1404
rect 355 1402 361 1403
rect 424 1394 426 1404
rect 430 1403 431 1407
rect 435 1403 436 1407
rect 430 1402 436 1403
rect 451 1407 457 1408
rect 451 1403 452 1407
rect 456 1406 457 1407
rect 502 1407 508 1408
rect 502 1406 503 1407
rect 456 1404 503 1406
rect 456 1403 457 1404
rect 451 1402 457 1403
rect 502 1403 503 1404
rect 507 1403 508 1407
rect 502 1402 508 1403
rect 526 1407 532 1408
rect 526 1403 527 1407
rect 531 1403 532 1407
rect 526 1402 532 1403
rect 542 1407 553 1408
rect 542 1403 543 1407
rect 547 1403 548 1407
rect 552 1403 553 1407
rect 542 1402 553 1403
rect 630 1407 636 1408
rect 630 1403 631 1407
rect 635 1403 636 1407
rect 651 1407 657 1408
rect 651 1406 652 1407
rect 630 1402 636 1403
rect 640 1404 652 1406
rect 640 1398 642 1404
rect 651 1403 652 1404
rect 656 1403 657 1407
rect 651 1402 657 1403
rect 726 1407 732 1408
rect 726 1403 727 1407
rect 731 1403 732 1407
rect 726 1402 732 1403
rect 747 1407 753 1408
rect 747 1403 748 1407
rect 752 1406 753 1407
rect 822 1407 828 1408
rect 752 1404 818 1406
rect 752 1403 753 1404
rect 747 1402 753 1403
rect 533 1396 642 1398
rect 533 1394 535 1396
rect 816 1394 818 1404
rect 822 1403 823 1407
rect 827 1403 828 1407
rect 822 1402 828 1403
rect 843 1407 849 1408
rect 843 1403 844 1407
rect 848 1406 849 1407
rect 910 1407 916 1408
rect 848 1404 902 1406
rect 848 1403 849 1404
rect 843 1402 849 1403
rect 900 1394 902 1404
rect 910 1403 911 1407
rect 915 1403 916 1407
rect 910 1402 916 1403
rect 931 1407 937 1408
rect 931 1403 932 1407
rect 936 1406 937 1407
rect 1006 1407 1012 1408
rect 936 1404 998 1406
rect 936 1403 937 1404
rect 931 1402 937 1403
rect 996 1394 998 1404
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1027 1407 1033 1408
rect 1027 1403 1028 1407
rect 1032 1406 1033 1407
rect 1102 1407 1108 1408
rect 1032 1404 1098 1406
rect 1032 1403 1033 1404
rect 1027 1402 1033 1403
rect 1096 1394 1098 1404
rect 1102 1403 1103 1407
rect 1107 1403 1108 1407
rect 1102 1402 1108 1403
rect 1122 1407 1129 1408
rect 1122 1403 1123 1407
rect 1128 1403 1129 1407
rect 1286 1404 1287 1408
rect 1291 1404 1292 1408
rect 1408 1406 1410 1412
rect 1414 1411 1415 1415
rect 1419 1414 1420 1415
rect 1427 1415 1433 1416
rect 1427 1414 1428 1415
rect 1419 1412 1428 1414
rect 1419 1411 1420 1412
rect 1414 1410 1420 1411
rect 1427 1411 1428 1412
rect 1432 1411 1433 1415
rect 1507 1413 1508 1417
rect 1512 1413 1513 1417
rect 1779 1417 1785 1418
rect 1595 1415 1601 1416
rect 1595 1414 1596 1415
rect 1507 1412 1513 1413
rect 1524 1412 1596 1414
rect 1427 1410 1433 1411
rect 1408 1404 1446 1406
rect 1286 1403 1292 1404
rect 1122 1402 1129 1403
rect 1444 1402 1446 1404
rect 1524 1402 1526 1412
rect 1595 1411 1596 1412
rect 1600 1411 1601 1415
rect 1683 1415 1689 1416
rect 1683 1414 1684 1415
rect 1595 1410 1601 1411
rect 1612 1412 1684 1414
rect 1612 1402 1614 1412
rect 1683 1411 1684 1412
rect 1688 1411 1689 1415
rect 1779 1413 1780 1417
rect 1784 1413 1785 1417
rect 1883 1415 1889 1416
rect 1883 1414 1884 1415
rect 1779 1412 1785 1413
rect 1796 1412 1884 1414
rect 1683 1410 1689 1411
rect 1796 1402 1798 1412
rect 1883 1411 1884 1412
rect 1888 1411 1889 1415
rect 1995 1415 2001 1416
rect 1995 1414 1996 1415
rect 1883 1410 1889 1411
rect 1900 1412 1996 1414
rect 1900 1402 1902 1412
rect 1995 1411 1996 1412
rect 2000 1411 2001 1415
rect 2115 1415 2121 1416
rect 2115 1414 2116 1415
rect 1995 1410 2001 1411
rect 2012 1412 2116 1414
rect 2012 1402 2014 1412
rect 2115 1411 2116 1412
rect 2120 1411 2121 1415
rect 2115 1410 2121 1411
rect 2235 1415 2241 1416
rect 2235 1411 2236 1415
rect 2240 1414 2241 1415
rect 2355 1415 2364 1416
rect 2240 1412 2350 1414
rect 2240 1411 2241 1412
rect 2235 1410 2241 1411
rect 2348 1406 2350 1412
rect 2355 1411 2356 1415
rect 2363 1411 2364 1415
rect 2355 1410 2364 1411
rect 2459 1415 2465 1416
rect 2459 1411 2460 1415
rect 2464 1414 2465 1415
rect 2470 1415 2476 1416
rect 2470 1414 2471 1415
rect 2464 1412 2471 1414
rect 2464 1411 2465 1412
rect 2459 1410 2465 1411
rect 2470 1411 2471 1412
rect 2475 1411 2476 1415
rect 2470 1410 2476 1411
rect 2348 1404 2374 1406
rect 2372 1402 2374 1404
rect 1366 1401 1372 1402
rect 1326 1400 1332 1401
rect 1326 1396 1327 1400
rect 1331 1396 1332 1400
rect 1366 1397 1367 1401
rect 1371 1397 1372 1401
rect 1422 1401 1428 1402
rect 1366 1396 1372 1397
rect 1374 1399 1380 1400
rect 1326 1395 1332 1396
rect 1374 1395 1375 1399
rect 1379 1398 1380 1399
rect 1387 1399 1393 1400
rect 1387 1398 1388 1399
rect 1379 1396 1388 1398
rect 1379 1395 1380 1396
rect 1374 1394 1380 1395
rect 1387 1395 1388 1396
rect 1392 1395 1393 1399
rect 1422 1397 1423 1401
rect 1427 1397 1428 1401
rect 1422 1396 1428 1397
rect 1443 1401 1449 1402
rect 1443 1397 1444 1401
rect 1448 1397 1449 1401
rect 1443 1396 1449 1397
rect 1502 1401 1508 1402
rect 1502 1397 1503 1401
rect 1507 1397 1508 1401
rect 1502 1396 1508 1397
rect 1523 1401 1529 1402
rect 1523 1397 1524 1401
rect 1528 1397 1529 1401
rect 1523 1396 1529 1397
rect 1590 1401 1596 1402
rect 1590 1397 1591 1401
rect 1595 1397 1596 1401
rect 1590 1396 1596 1397
rect 1611 1401 1617 1402
rect 1611 1397 1612 1401
rect 1616 1397 1617 1401
rect 1611 1396 1617 1397
rect 1678 1401 1684 1402
rect 1678 1397 1679 1401
rect 1683 1397 1684 1401
rect 1774 1401 1780 1402
rect 1678 1396 1684 1397
rect 1699 1399 1708 1400
rect 1387 1394 1393 1395
rect 1699 1395 1700 1399
rect 1707 1395 1708 1399
rect 1774 1397 1775 1401
rect 1779 1397 1780 1401
rect 1774 1396 1780 1397
rect 1795 1401 1801 1402
rect 1795 1397 1796 1401
rect 1800 1397 1801 1401
rect 1795 1396 1801 1397
rect 1878 1401 1884 1402
rect 1878 1397 1879 1401
rect 1883 1397 1884 1401
rect 1878 1396 1884 1397
rect 1899 1401 1905 1402
rect 1899 1397 1900 1401
rect 1904 1397 1905 1401
rect 1899 1396 1905 1397
rect 1990 1401 1996 1402
rect 1990 1397 1991 1401
rect 1995 1397 1996 1401
rect 1990 1396 1996 1397
rect 2011 1401 2017 1402
rect 2011 1397 2012 1401
rect 2016 1397 2017 1401
rect 2011 1396 2017 1397
rect 2110 1401 2116 1402
rect 2110 1397 2111 1401
rect 2115 1397 2116 1401
rect 2230 1401 2236 1402
rect 2110 1396 2116 1397
rect 2118 1399 2124 1400
rect 1699 1394 1708 1395
rect 2118 1395 2119 1399
rect 2123 1398 2124 1399
rect 2131 1399 2137 1400
rect 2131 1398 2132 1399
rect 2123 1396 2132 1398
rect 2123 1395 2124 1396
rect 2118 1394 2124 1395
rect 2131 1395 2132 1396
rect 2136 1395 2137 1399
rect 2230 1397 2231 1401
rect 2235 1397 2236 1401
rect 2350 1401 2356 1402
rect 2230 1396 2236 1397
rect 2251 1399 2260 1400
rect 2131 1394 2137 1395
rect 2251 1395 2252 1399
rect 2259 1395 2260 1399
rect 2350 1397 2351 1401
rect 2355 1397 2356 1401
rect 2350 1396 2356 1397
rect 2371 1401 2377 1402
rect 2371 1397 2372 1401
rect 2376 1397 2377 1401
rect 2371 1396 2377 1397
rect 2454 1401 2460 1402
rect 2454 1397 2455 1401
rect 2459 1397 2460 1401
rect 2502 1400 2508 1401
rect 2454 1396 2460 1397
rect 2462 1399 2468 1400
rect 2251 1394 2260 1395
rect 2462 1395 2463 1399
rect 2467 1398 2468 1399
rect 2475 1399 2481 1400
rect 2475 1398 2476 1399
rect 2467 1396 2476 1398
rect 2467 1395 2468 1396
rect 2462 1394 2468 1395
rect 2475 1395 2476 1396
rect 2480 1395 2481 1399
rect 2502 1396 2503 1400
rect 2507 1396 2508 1400
rect 2502 1395 2508 1396
rect 2475 1394 2481 1395
rect 319 1393 345 1394
rect 319 1392 340 1393
rect 251 1391 257 1392
rect 251 1387 252 1391
rect 256 1390 257 1391
rect 256 1388 321 1390
rect 339 1389 340 1392
rect 344 1389 345 1393
rect 424 1393 441 1394
rect 424 1392 436 1393
rect 339 1388 345 1389
rect 435 1389 436 1392
rect 440 1389 441 1393
rect 435 1388 441 1389
rect 531 1393 537 1394
rect 531 1389 532 1393
rect 536 1389 537 1393
rect 816 1393 833 1394
rect 816 1392 828 1393
rect 531 1388 537 1389
rect 622 1391 628 1392
rect 256 1387 257 1388
rect 251 1386 257 1387
rect 319 1386 321 1388
rect 542 1387 548 1388
rect 542 1386 543 1387
rect 319 1384 543 1386
rect 542 1383 543 1384
rect 547 1383 548 1387
rect 622 1387 623 1391
rect 627 1390 628 1391
rect 635 1391 641 1392
rect 635 1390 636 1391
rect 627 1388 636 1390
rect 627 1387 628 1388
rect 622 1386 628 1387
rect 635 1387 636 1388
rect 640 1387 641 1391
rect 635 1386 641 1387
rect 731 1391 737 1392
rect 731 1387 732 1391
rect 736 1387 737 1391
rect 827 1389 828 1392
rect 832 1389 833 1393
rect 900 1393 921 1394
rect 900 1392 916 1393
rect 827 1388 833 1389
rect 915 1389 916 1392
rect 920 1389 921 1393
rect 996 1393 1017 1394
rect 996 1392 1012 1393
rect 915 1388 921 1389
rect 1011 1389 1012 1392
rect 1016 1389 1017 1393
rect 1096 1393 1113 1394
rect 1096 1392 1108 1393
rect 1011 1388 1017 1389
rect 1107 1389 1108 1392
rect 1112 1389 1113 1393
rect 1107 1388 1113 1389
rect 731 1386 737 1387
rect 1022 1387 1028 1388
rect 1022 1386 1023 1387
rect 733 1384 1023 1386
rect 542 1382 548 1383
rect 1022 1383 1023 1384
rect 1027 1383 1028 1387
rect 1022 1382 1028 1383
rect 1326 1383 1332 1384
rect 902 1379 908 1380
rect 902 1378 903 1379
rect 613 1376 903 1378
rect 613 1374 615 1376
rect 902 1375 903 1376
rect 907 1375 908 1379
rect 1326 1379 1327 1383
rect 1331 1379 1332 1383
rect 2502 1383 2508 1384
rect 1326 1378 1332 1379
rect 1350 1380 1356 1381
rect 1350 1376 1351 1380
rect 1355 1376 1356 1380
rect 1350 1375 1356 1376
rect 1406 1380 1412 1381
rect 1406 1376 1407 1380
rect 1411 1376 1412 1380
rect 1406 1375 1412 1376
rect 1486 1380 1492 1381
rect 1486 1376 1487 1380
rect 1491 1376 1492 1380
rect 1486 1375 1492 1376
rect 1574 1380 1580 1381
rect 1574 1376 1575 1380
rect 1579 1376 1580 1380
rect 1574 1375 1580 1376
rect 1662 1380 1668 1381
rect 1662 1376 1663 1380
rect 1667 1376 1668 1380
rect 1662 1375 1668 1376
rect 1758 1380 1764 1381
rect 1758 1376 1759 1380
rect 1763 1376 1764 1380
rect 1758 1375 1764 1376
rect 1862 1380 1868 1381
rect 1862 1376 1863 1380
rect 1867 1376 1868 1380
rect 1862 1375 1868 1376
rect 1974 1380 1980 1381
rect 1974 1376 1975 1380
rect 1979 1376 1980 1380
rect 1974 1375 1980 1376
rect 2094 1380 2100 1381
rect 2094 1376 2095 1380
rect 2099 1376 2100 1380
rect 2094 1375 2100 1376
rect 2214 1380 2220 1381
rect 2214 1376 2215 1380
rect 2219 1376 2220 1380
rect 2214 1375 2220 1376
rect 2334 1380 2340 1381
rect 2334 1376 2335 1380
rect 2339 1376 2340 1380
rect 2334 1375 2340 1376
rect 2438 1380 2444 1381
rect 2438 1376 2439 1380
rect 2443 1376 2444 1380
rect 2502 1379 2503 1383
rect 2507 1379 2508 1383
rect 2502 1378 2508 1379
rect 2438 1375 2444 1376
rect 902 1374 908 1375
rect 611 1373 617 1374
rect 155 1371 161 1372
rect 155 1367 156 1371
rect 160 1367 161 1371
rect 155 1366 161 1367
rect 219 1371 225 1372
rect 219 1367 220 1371
rect 224 1370 225 1371
rect 315 1371 321 1372
rect 224 1368 274 1370
rect 224 1367 225 1368
rect 219 1366 225 1367
rect 157 1362 159 1366
rect 272 1362 274 1368
rect 315 1367 316 1371
rect 320 1370 321 1371
rect 411 1371 417 1372
rect 320 1368 407 1370
rect 320 1367 321 1368
rect 315 1366 321 1367
rect 405 1362 407 1368
rect 411 1367 412 1371
rect 416 1370 417 1371
rect 502 1371 508 1372
rect 416 1368 486 1370
rect 416 1367 417 1368
rect 411 1366 417 1367
rect 484 1362 486 1368
rect 502 1367 503 1371
rect 507 1370 508 1371
rect 515 1371 521 1372
rect 515 1370 516 1371
rect 507 1368 516 1370
rect 507 1367 508 1368
rect 502 1366 508 1367
rect 515 1367 516 1368
rect 520 1367 521 1371
rect 611 1369 612 1373
rect 616 1369 617 1373
rect 707 1371 713 1372
rect 707 1370 708 1371
rect 611 1368 617 1369
rect 629 1368 708 1370
rect 515 1366 521 1367
rect 157 1360 238 1362
rect 272 1360 335 1362
rect 405 1360 430 1362
rect 484 1360 535 1362
rect 236 1358 238 1360
rect 333 1358 335 1360
rect 428 1358 430 1360
rect 533 1358 535 1360
rect 629 1358 631 1368
rect 707 1367 708 1368
rect 712 1367 713 1371
rect 803 1371 809 1372
rect 803 1370 804 1371
rect 707 1366 713 1367
rect 724 1368 804 1370
rect 724 1358 726 1368
rect 803 1367 804 1368
rect 808 1367 809 1371
rect 899 1371 905 1372
rect 899 1370 900 1371
rect 803 1366 809 1367
rect 821 1368 900 1370
rect 821 1358 823 1368
rect 899 1367 900 1368
rect 904 1367 905 1371
rect 1003 1371 1009 1372
rect 1003 1370 1004 1371
rect 899 1366 905 1367
rect 916 1368 1004 1370
rect 916 1358 918 1368
rect 1003 1367 1004 1368
rect 1008 1367 1009 1371
rect 1003 1366 1009 1367
rect 1350 1364 1356 1365
rect 1326 1361 1332 1362
rect 150 1357 156 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 150 1353 151 1357
rect 155 1353 156 1357
rect 214 1357 220 1358
rect 150 1352 156 1353
rect 158 1355 164 1356
rect 110 1351 116 1352
rect 158 1351 159 1355
rect 163 1354 164 1355
rect 171 1355 177 1356
rect 171 1354 172 1355
rect 163 1352 172 1354
rect 163 1351 164 1352
rect 158 1350 164 1351
rect 171 1351 172 1352
rect 176 1351 177 1355
rect 214 1353 215 1357
rect 219 1353 220 1357
rect 214 1352 220 1353
rect 235 1357 241 1358
rect 235 1353 236 1357
rect 240 1353 241 1357
rect 235 1352 241 1353
rect 310 1357 316 1358
rect 310 1353 311 1357
rect 315 1353 316 1357
rect 310 1352 316 1353
rect 331 1357 337 1358
rect 331 1353 332 1357
rect 336 1353 337 1357
rect 331 1352 337 1353
rect 406 1357 412 1358
rect 406 1353 407 1357
rect 411 1353 412 1357
rect 406 1352 412 1353
rect 427 1357 433 1358
rect 427 1353 428 1357
rect 432 1353 433 1357
rect 427 1352 433 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 531 1357 537 1358
rect 531 1353 532 1357
rect 536 1353 537 1357
rect 531 1352 537 1353
rect 606 1357 612 1358
rect 606 1353 607 1357
rect 611 1353 612 1357
rect 606 1352 612 1353
rect 627 1357 633 1358
rect 627 1353 628 1357
rect 632 1353 633 1357
rect 627 1352 633 1353
rect 702 1357 708 1358
rect 702 1353 703 1357
rect 707 1353 708 1357
rect 702 1352 708 1353
rect 723 1357 729 1358
rect 723 1353 724 1357
rect 728 1353 729 1357
rect 723 1352 729 1353
rect 798 1357 804 1358
rect 798 1353 799 1357
rect 803 1353 804 1357
rect 798 1352 804 1353
rect 819 1357 825 1358
rect 819 1353 820 1357
rect 824 1353 825 1357
rect 819 1352 825 1353
rect 894 1357 900 1358
rect 894 1353 895 1357
rect 899 1353 900 1357
rect 894 1352 900 1353
rect 915 1357 921 1358
rect 915 1353 916 1357
rect 920 1353 921 1357
rect 915 1352 921 1353
rect 998 1357 1004 1358
rect 1326 1357 1327 1361
rect 1331 1357 1332 1361
rect 1350 1360 1351 1364
rect 1355 1360 1356 1364
rect 1350 1359 1356 1360
rect 1406 1364 1412 1365
rect 1406 1360 1407 1364
rect 1411 1360 1412 1364
rect 1406 1359 1412 1360
rect 1478 1364 1484 1365
rect 1478 1360 1479 1364
rect 1483 1360 1484 1364
rect 1478 1359 1484 1360
rect 1566 1364 1572 1365
rect 1566 1360 1567 1364
rect 1571 1360 1572 1364
rect 1566 1359 1572 1360
rect 1654 1364 1660 1365
rect 1654 1360 1655 1364
rect 1659 1360 1660 1364
rect 1654 1359 1660 1360
rect 1750 1364 1756 1365
rect 1750 1360 1751 1364
rect 1755 1360 1756 1364
rect 1750 1359 1756 1360
rect 1854 1364 1860 1365
rect 1854 1360 1855 1364
rect 1859 1360 1860 1364
rect 1854 1359 1860 1360
rect 1966 1364 1972 1365
rect 1966 1360 1967 1364
rect 1971 1360 1972 1364
rect 1966 1359 1972 1360
rect 2078 1364 2084 1365
rect 2078 1360 2079 1364
rect 2083 1360 2084 1364
rect 2078 1359 2084 1360
rect 2198 1364 2204 1365
rect 2198 1360 2199 1364
rect 2203 1360 2204 1364
rect 2198 1359 2204 1360
rect 2326 1364 2332 1365
rect 2326 1360 2327 1364
rect 2331 1360 2332 1364
rect 2326 1359 2332 1360
rect 2438 1364 2444 1365
rect 2438 1360 2439 1364
rect 2443 1360 2444 1364
rect 2438 1359 2444 1360
rect 2502 1361 2508 1362
rect 998 1353 999 1357
rect 1003 1353 1004 1357
rect 1286 1356 1292 1357
rect 1326 1356 1332 1357
rect 2502 1357 2503 1361
rect 2507 1357 2508 1361
rect 2502 1356 2508 1357
rect 998 1352 1004 1353
rect 1019 1355 1028 1356
rect 171 1350 177 1351
rect 1019 1351 1020 1355
rect 1027 1351 1028 1355
rect 1286 1352 1287 1356
rect 1291 1352 1292 1356
rect 1286 1351 1292 1352
rect 1019 1350 1028 1351
rect 1326 1344 1332 1345
rect 2502 1344 2508 1345
rect 1326 1340 1327 1344
rect 1331 1340 1332 1344
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 1286 1339 1292 1340
rect 1326 1339 1332 1340
rect 1366 1343 1372 1344
rect 1366 1339 1367 1343
rect 1371 1339 1372 1343
rect 110 1334 116 1335
rect 134 1336 140 1337
rect 134 1332 135 1336
rect 139 1332 140 1336
rect 134 1331 140 1332
rect 198 1336 204 1337
rect 198 1332 199 1336
rect 203 1332 204 1336
rect 198 1331 204 1332
rect 294 1336 300 1337
rect 294 1332 295 1336
rect 299 1332 300 1336
rect 294 1331 300 1332
rect 390 1336 396 1337
rect 390 1332 391 1336
rect 395 1332 396 1336
rect 390 1331 396 1332
rect 494 1336 500 1337
rect 494 1332 495 1336
rect 499 1332 500 1336
rect 494 1331 500 1332
rect 590 1336 596 1337
rect 590 1332 591 1336
rect 595 1332 596 1336
rect 590 1331 596 1332
rect 686 1336 692 1337
rect 686 1332 687 1336
rect 691 1332 692 1336
rect 686 1331 692 1332
rect 782 1336 788 1337
rect 782 1332 783 1336
rect 787 1332 788 1336
rect 782 1331 788 1332
rect 878 1336 884 1337
rect 878 1332 879 1336
rect 883 1332 884 1336
rect 878 1331 884 1332
rect 982 1336 988 1337
rect 982 1332 983 1336
rect 987 1332 988 1336
rect 1286 1335 1287 1339
rect 1291 1335 1292 1339
rect 1366 1338 1372 1339
rect 1387 1343 1393 1344
rect 1387 1339 1388 1343
rect 1392 1339 1393 1343
rect 1387 1338 1393 1339
rect 1422 1343 1428 1344
rect 1422 1339 1423 1343
rect 1427 1339 1428 1343
rect 1422 1338 1428 1339
rect 1443 1343 1449 1344
rect 1443 1339 1444 1343
rect 1448 1342 1449 1343
rect 1494 1343 1500 1344
rect 1448 1340 1490 1342
rect 1448 1339 1449 1340
rect 1443 1338 1449 1339
rect 1286 1334 1292 1335
rect 982 1331 988 1332
rect 1389 1330 1391 1338
rect 1488 1330 1490 1340
rect 1494 1339 1495 1343
rect 1499 1339 1500 1343
rect 1494 1338 1500 1339
rect 1515 1343 1521 1344
rect 1515 1339 1516 1343
rect 1520 1342 1521 1343
rect 1526 1343 1532 1344
rect 1526 1342 1527 1343
rect 1520 1340 1527 1342
rect 1520 1339 1521 1340
rect 1515 1338 1521 1339
rect 1526 1339 1527 1340
rect 1531 1339 1532 1343
rect 1526 1338 1532 1339
rect 1582 1343 1588 1344
rect 1582 1339 1583 1343
rect 1587 1339 1588 1343
rect 1582 1338 1588 1339
rect 1602 1343 1609 1344
rect 1602 1339 1603 1343
rect 1608 1339 1609 1343
rect 1602 1338 1609 1339
rect 1670 1343 1676 1344
rect 1670 1339 1671 1343
rect 1675 1339 1676 1343
rect 1691 1343 1697 1344
rect 1691 1342 1692 1343
rect 1670 1338 1676 1339
rect 1680 1340 1692 1342
rect 1680 1334 1682 1340
rect 1691 1339 1692 1340
rect 1696 1339 1697 1343
rect 1691 1338 1697 1339
rect 1766 1343 1772 1344
rect 1766 1339 1767 1343
rect 1771 1339 1772 1343
rect 1787 1343 1793 1344
rect 1787 1342 1788 1343
rect 1766 1338 1772 1339
rect 1776 1340 1788 1342
rect 1776 1334 1778 1340
rect 1787 1339 1788 1340
rect 1792 1339 1793 1343
rect 1787 1338 1793 1339
rect 1870 1343 1876 1344
rect 1870 1339 1871 1343
rect 1875 1339 1876 1343
rect 1870 1338 1876 1339
rect 1891 1343 1897 1344
rect 1891 1339 1892 1343
rect 1896 1342 1897 1343
rect 1982 1343 1988 1344
rect 1896 1340 1978 1342
rect 1896 1339 1897 1340
rect 1891 1338 1897 1339
rect 1588 1332 1682 1334
rect 1684 1332 1778 1334
rect 1588 1330 1590 1332
rect 1684 1330 1686 1332
rect 1389 1329 1433 1330
rect 1389 1328 1428 1329
rect 1371 1327 1380 1328
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 414 1324 420 1325
rect 414 1320 415 1324
rect 419 1320 420 1324
rect 414 1319 420 1320
rect 510 1324 516 1325
rect 510 1320 511 1324
rect 515 1320 516 1324
rect 510 1319 516 1320
rect 598 1324 604 1325
rect 598 1320 599 1324
rect 603 1320 604 1324
rect 598 1319 604 1320
rect 686 1324 692 1325
rect 686 1320 687 1324
rect 691 1320 692 1324
rect 686 1319 692 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 878 1324 884 1325
rect 878 1320 879 1324
rect 883 1320 884 1324
rect 1371 1323 1372 1327
rect 1379 1323 1380 1327
rect 1427 1325 1428 1328
rect 1432 1325 1433 1329
rect 1488 1329 1505 1330
rect 1488 1328 1500 1329
rect 1427 1324 1433 1325
rect 1499 1325 1500 1328
rect 1504 1325 1505 1329
rect 1499 1324 1505 1325
rect 1587 1329 1593 1330
rect 1587 1325 1588 1329
rect 1592 1325 1593 1329
rect 1587 1324 1593 1325
rect 1675 1329 1686 1330
rect 1675 1325 1676 1329
rect 1680 1328 1686 1329
rect 1976 1330 1978 1340
rect 1982 1339 1983 1343
rect 1987 1339 1988 1343
rect 1982 1338 1988 1339
rect 2003 1343 2009 1344
rect 2003 1339 2004 1343
rect 2008 1339 2009 1343
rect 2003 1338 2009 1339
rect 2094 1343 2100 1344
rect 2094 1339 2095 1343
rect 2099 1339 2100 1343
rect 2094 1338 2100 1339
rect 2115 1343 2121 1344
rect 2115 1339 2116 1343
rect 2120 1342 2121 1343
rect 2214 1343 2220 1344
rect 2120 1340 2210 1342
rect 2120 1339 2121 1340
rect 2115 1338 2121 1339
rect 2005 1330 2007 1338
rect 2208 1330 2210 1340
rect 2214 1339 2215 1343
rect 2219 1339 2220 1343
rect 2214 1338 2220 1339
rect 2222 1343 2228 1344
rect 2222 1339 2223 1343
rect 2227 1342 2228 1343
rect 2235 1343 2241 1344
rect 2235 1342 2236 1343
rect 2227 1340 2236 1342
rect 2227 1339 2228 1340
rect 2222 1338 2228 1339
rect 2235 1339 2236 1340
rect 2240 1339 2241 1343
rect 2235 1338 2241 1339
rect 2342 1343 2348 1344
rect 2342 1339 2343 1343
rect 2347 1339 2348 1343
rect 2342 1338 2348 1339
rect 2358 1343 2369 1344
rect 2358 1339 2359 1343
rect 2363 1339 2364 1343
rect 2368 1339 2369 1343
rect 2358 1338 2369 1339
rect 2454 1343 2460 1344
rect 2454 1339 2455 1343
rect 2459 1339 2460 1343
rect 2454 1338 2460 1339
rect 2470 1343 2481 1344
rect 2470 1339 2471 1343
rect 2475 1339 2476 1343
rect 2480 1339 2481 1343
rect 2502 1340 2503 1344
rect 2507 1340 2508 1344
rect 2502 1339 2508 1340
rect 2470 1338 2481 1339
rect 1976 1329 1993 1330
rect 1976 1328 1988 1329
rect 1680 1325 1681 1328
rect 1675 1324 1681 1325
rect 1742 1327 1748 1328
rect 1371 1322 1380 1323
rect 1742 1323 1743 1327
rect 1747 1326 1748 1327
rect 1771 1327 1777 1328
rect 1771 1326 1772 1327
rect 1747 1324 1772 1326
rect 1747 1323 1748 1324
rect 1742 1322 1748 1323
rect 1771 1323 1772 1324
rect 1776 1323 1777 1327
rect 1771 1322 1777 1323
rect 1875 1327 1881 1328
rect 1875 1323 1876 1327
rect 1880 1326 1881 1327
rect 1880 1324 1942 1326
rect 1987 1325 1988 1328
rect 1992 1325 1993 1329
rect 2005 1329 2105 1330
rect 2005 1328 2100 1329
rect 1987 1324 1993 1325
rect 2099 1325 2100 1328
rect 2104 1325 2105 1329
rect 2208 1329 2225 1330
rect 2208 1328 2220 1329
rect 2099 1324 2105 1325
rect 2219 1325 2220 1328
rect 2224 1325 2225 1329
rect 2219 1324 2225 1325
rect 2347 1327 2356 1328
rect 1880 1323 1881 1324
rect 1875 1322 1881 1323
rect 1940 1322 1942 1324
rect 2118 1323 2124 1324
rect 2118 1322 2119 1323
rect 878 1319 884 1320
rect 1286 1321 1292 1322
rect 110 1316 116 1317
rect 1286 1317 1287 1321
rect 1291 1317 1292 1321
rect 1940 1320 2119 1322
rect 2118 1319 2119 1320
rect 2123 1319 2124 1323
rect 2347 1323 2348 1327
rect 2355 1323 2356 1327
rect 2347 1322 2356 1323
rect 2459 1327 2468 1328
rect 2459 1323 2460 1327
rect 2467 1323 2468 1327
rect 2459 1322 2468 1323
rect 2118 1318 2124 1319
rect 1286 1316 1292 1317
rect 1842 1307 1848 1308
rect 1842 1306 1843 1307
rect 110 1304 116 1305
rect 1286 1304 1292 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 150 1303 156 1304
rect 150 1299 151 1303
rect 155 1299 156 1303
rect 150 1298 156 1299
rect 171 1303 177 1304
rect 171 1299 172 1303
rect 176 1299 177 1303
rect 171 1298 177 1299
rect 230 1303 236 1304
rect 230 1299 231 1303
rect 235 1299 236 1303
rect 230 1298 236 1299
rect 251 1303 257 1304
rect 251 1299 252 1303
rect 256 1302 257 1303
rect 334 1303 340 1304
rect 256 1300 321 1302
rect 256 1299 257 1300
rect 251 1298 257 1299
rect 173 1290 175 1298
rect 319 1290 321 1300
rect 334 1299 335 1303
rect 339 1299 340 1303
rect 334 1298 340 1299
rect 355 1303 361 1304
rect 355 1299 356 1303
rect 360 1302 361 1303
rect 430 1303 436 1304
rect 360 1300 426 1302
rect 360 1299 361 1300
rect 355 1298 361 1299
rect 424 1290 426 1300
rect 430 1299 431 1303
rect 435 1299 436 1303
rect 430 1298 436 1299
rect 446 1303 457 1304
rect 446 1299 447 1303
rect 451 1299 452 1303
rect 456 1299 457 1303
rect 446 1298 457 1299
rect 526 1303 532 1304
rect 526 1299 527 1303
rect 531 1299 532 1303
rect 526 1298 532 1299
rect 547 1303 553 1304
rect 547 1299 548 1303
rect 552 1302 553 1303
rect 614 1303 620 1304
rect 552 1300 606 1302
rect 552 1299 553 1300
rect 547 1298 553 1299
rect 604 1290 606 1300
rect 614 1299 615 1303
rect 619 1299 620 1303
rect 614 1298 620 1299
rect 635 1303 641 1304
rect 635 1299 636 1303
rect 640 1302 641 1303
rect 702 1303 708 1304
rect 640 1300 694 1302
rect 640 1299 641 1300
rect 635 1298 641 1299
rect 692 1290 694 1300
rect 702 1299 703 1303
rect 707 1299 708 1303
rect 702 1298 708 1299
rect 723 1303 729 1304
rect 723 1299 724 1303
rect 728 1302 729 1303
rect 798 1303 804 1304
rect 728 1300 794 1302
rect 728 1299 729 1300
rect 723 1298 729 1299
rect 792 1290 794 1300
rect 798 1299 799 1303
rect 803 1299 804 1303
rect 798 1298 804 1299
rect 819 1303 825 1304
rect 819 1299 820 1303
rect 824 1299 825 1303
rect 819 1298 825 1299
rect 894 1303 900 1304
rect 894 1299 895 1303
rect 899 1299 900 1303
rect 894 1298 900 1299
rect 902 1303 908 1304
rect 902 1299 903 1303
rect 907 1302 908 1303
rect 915 1303 921 1304
rect 915 1302 916 1303
rect 907 1300 916 1302
rect 907 1299 908 1300
rect 902 1298 908 1299
rect 915 1299 916 1300
rect 920 1299 921 1303
rect 1286 1300 1287 1304
rect 1291 1300 1292 1304
rect 1620 1304 1843 1306
rect 1620 1302 1622 1304
rect 1842 1303 1843 1304
rect 1847 1303 1848 1307
rect 2222 1307 2228 1308
rect 2222 1306 2223 1307
rect 1842 1302 1848 1303
rect 1924 1304 2223 1306
rect 1924 1302 1926 1304
rect 2222 1303 2223 1304
rect 2227 1303 2228 1307
rect 2470 1307 2476 1308
rect 2470 1306 2471 1307
rect 2222 1302 2228 1303
rect 2404 1304 2471 1306
rect 2404 1302 2406 1304
rect 2470 1303 2471 1304
rect 2475 1303 2476 1307
rect 2470 1302 2476 1303
rect 1619 1301 1625 1302
rect 1286 1299 1292 1300
rect 1371 1299 1377 1300
rect 915 1298 921 1299
rect 821 1290 823 1298
rect 1371 1295 1372 1299
rect 1376 1298 1377 1299
rect 1427 1299 1433 1300
rect 1376 1296 1422 1298
rect 1376 1295 1377 1296
rect 1371 1294 1377 1295
rect 1246 1291 1252 1292
rect 173 1289 241 1290
rect 173 1288 236 1289
rect 155 1287 164 1288
rect 155 1283 156 1287
rect 163 1283 164 1287
rect 235 1285 236 1288
rect 240 1285 241 1289
rect 319 1289 345 1290
rect 319 1288 340 1289
rect 235 1284 241 1285
rect 339 1285 340 1288
rect 344 1285 345 1289
rect 424 1289 441 1290
rect 424 1288 436 1289
rect 339 1284 345 1285
rect 435 1285 436 1288
rect 440 1285 441 1289
rect 604 1289 625 1290
rect 604 1288 620 1289
rect 435 1284 441 1285
rect 531 1287 537 1288
rect 155 1282 164 1283
rect 531 1283 532 1287
rect 536 1283 537 1287
rect 619 1285 620 1288
rect 624 1285 625 1289
rect 692 1289 713 1290
rect 692 1288 708 1289
rect 619 1284 625 1285
rect 707 1285 708 1288
rect 712 1285 713 1289
rect 792 1289 809 1290
rect 792 1288 804 1289
rect 707 1284 713 1285
rect 803 1285 804 1288
rect 808 1285 809 1289
rect 821 1289 905 1290
rect 821 1288 900 1289
rect 803 1284 809 1285
rect 899 1285 900 1288
rect 904 1285 905 1289
rect 1246 1287 1247 1291
rect 1251 1290 1252 1291
rect 1420 1290 1422 1296
rect 1427 1295 1428 1299
rect 1432 1298 1433 1299
rect 1523 1299 1532 1300
rect 1432 1296 1521 1298
rect 1432 1295 1433 1296
rect 1427 1294 1433 1295
rect 1519 1290 1521 1296
rect 1523 1295 1524 1299
rect 1531 1295 1532 1299
rect 1619 1297 1620 1301
rect 1624 1297 1625 1301
rect 1923 1301 1929 1302
rect 1723 1299 1729 1300
rect 1723 1298 1724 1299
rect 1619 1296 1625 1297
rect 1636 1296 1724 1298
rect 1523 1294 1532 1295
rect 1251 1288 1391 1290
rect 1420 1288 1446 1290
rect 1519 1288 1542 1290
rect 1251 1287 1252 1288
rect 1246 1286 1252 1287
rect 1389 1286 1391 1288
rect 1444 1286 1446 1288
rect 1540 1286 1542 1288
rect 1636 1286 1638 1296
rect 1723 1295 1724 1296
rect 1728 1295 1729 1299
rect 1723 1294 1729 1295
rect 1827 1299 1833 1300
rect 1827 1295 1828 1299
rect 1832 1298 1833 1299
rect 1850 1299 1856 1300
rect 1850 1298 1851 1299
rect 1832 1296 1851 1298
rect 1832 1295 1833 1296
rect 1827 1294 1833 1295
rect 1850 1295 1851 1296
rect 1855 1295 1856 1299
rect 1923 1297 1924 1301
rect 1928 1297 1929 1301
rect 2403 1301 2409 1302
rect 2019 1299 2025 1300
rect 2019 1298 2020 1299
rect 1923 1296 1929 1297
rect 1999 1296 2020 1298
rect 1850 1294 1856 1295
rect 1999 1290 2001 1296
rect 2019 1295 2020 1296
rect 2024 1295 2025 1299
rect 2107 1299 2113 1300
rect 2107 1298 2108 1299
rect 2019 1294 2025 1295
rect 2036 1296 2108 1298
rect 1940 1288 2001 1290
rect 1940 1286 1942 1288
rect 2036 1286 2038 1296
rect 2107 1295 2108 1296
rect 2112 1295 2113 1299
rect 2187 1299 2193 1300
rect 2187 1298 2188 1299
rect 2107 1294 2113 1295
rect 2124 1296 2188 1298
rect 2124 1286 2126 1296
rect 2187 1295 2188 1296
rect 2192 1295 2193 1299
rect 2259 1299 2265 1300
rect 2259 1298 2260 1299
rect 2187 1294 2193 1295
rect 2204 1296 2260 1298
rect 2204 1286 2206 1296
rect 2259 1295 2260 1296
rect 2264 1295 2265 1299
rect 2259 1294 2265 1295
rect 2331 1299 2337 1300
rect 2331 1295 2332 1299
rect 2336 1298 2337 1299
rect 2336 1296 2398 1298
rect 2403 1297 2404 1301
rect 2408 1297 2409 1301
rect 2403 1296 2409 1297
rect 2459 1299 2465 1300
rect 2336 1295 2337 1296
rect 2331 1294 2337 1295
rect 2396 1290 2398 1296
rect 2459 1295 2460 1299
rect 2464 1295 2465 1299
rect 2459 1294 2465 1295
rect 2410 1291 2416 1292
rect 2410 1290 2411 1291
rect 2396 1288 2411 1290
rect 2410 1287 2411 1288
rect 2415 1287 2416 1291
rect 2461 1290 2463 1294
rect 2410 1286 2416 1287
rect 2420 1288 2463 1290
rect 2420 1286 2422 1288
rect 1366 1285 1372 1286
rect 899 1284 905 1285
rect 1326 1284 1332 1285
rect 531 1282 537 1283
rect 1114 1283 1120 1284
rect 1114 1282 1115 1283
rect 533 1280 1115 1282
rect 1114 1279 1115 1280
rect 1119 1279 1120 1283
rect 1326 1280 1327 1284
rect 1331 1280 1332 1284
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 1387 1285 1393 1286
rect 1387 1281 1388 1285
rect 1392 1281 1393 1285
rect 1387 1280 1393 1281
rect 1422 1285 1428 1286
rect 1422 1281 1423 1285
rect 1427 1281 1428 1285
rect 1422 1280 1428 1281
rect 1443 1285 1449 1286
rect 1443 1281 1444 1285
rect 1448 1281 1449 1285
rect 1443 1280 1449 1281
rect 1518 1285 1524 1286
rect 1518 1281 1519 1285
rect 1523 1281 1524 1285
rect 1518 1280 1524 1281
rect 1539 1285 1545 1286
rect 1539 1281 1540 1285
rect 1544 1281 1545 1285
rect 1539 1280 1545 1281
rect 1614 1285 1620 1286
rect 1614 1281 1615 1285
rect 1619 1281 1620 1285
rect 1614 1280 1620 1281
rect 1635 1285 1641 1286
rect 1635 1281 1636 1285
rect 1640 1281 1641 1285
rect 1635 1280 1641 1281
rect 1718 1285 1724 1286
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1822 1285 1828 1286
rect 1718 1280 1724 1281
rect 1739 1283 1748 1284
rect 1326 1279 1332 1280
rect 1739 1279 1740 1283
rect 1747 1279 1748 1283
rect 1822 1281 1823 1285
rect 1827 1281 1828 1285
rect 1918 1285 1924 1286
rect 1822 1280 1828 1281
rect 1842 1283 1849 1284
rect 1114 1278 1120 1279
rect 1739 1278 1748 1279
rect 1842 1279 1843 1283
rect 1848 1279 1849 1283
rect 1918 1281 1919 1285
rect 1923 1281 1924 1285
rect 1918 1280 1924 1281
rect 1939 1285 1945 1286
rect 1939 1281 1940 1285
rect 1944 1281 1945 1285
rect 1939 1280 1945 1281
rect 2014 1285 2020 1286
rect 2014 1281 2015 1285
rect 2019 1281 2020 1285
rect 2014 1280 2020 1281
rect 2035 1285 2041 1286
rect 2035 1281 2036 1285
rect 2040 1281 2041 1285
rect 2035 1280 2041 1281
rect 2102 1285 2108 1286
rect 2102 1281 2103 1285
rect 2107 1281 2108 1285
rect 2102 1280 2108 1281
rect 2123 1285 2129 1286
rect 2123 1281 2124 1285
rect 2128 1281 2129 1285
rect 2123 1280 2129 1281
rect 2182 1285 2188 1286
rect 2182 1281 2183 1285
rect 2187 1281 2188 1285
rect 2182 1280 2188 1281
rect 2203 1285 2209 1286
rect 2203 1281 2204 1285
rect 2208 1281 2209 1285
rect 2203 1280 2209 1281
rect 2254 1285 2260 1286
rect 2254 1281 2255 1285
rect 2259 1281 2260 1285
rect 2326 1285 2332 1286
rect 2254 1280 2260 1281
rect 2262 1283 2268 1284
rect 1842 1278 1849 1279
rect 2262 1279 2263 1283
rect 2267 1282 2268 1283
rect 2275 1283 2281 1284
rect 2275 1282 2276 1283
rect 2267 1280 2276 1282
rect 2267 1279 2268 1280
rect 2262 1278 2268 1279
rect 2275 1279 2276 1280
rect 2280 1279 2281 1283
rect 2326 1281 2327 1285
rect 2331 1281 2332 1285
rect 2398 1285 2404 1286
rect 2326 1280 2332 1281
rect 2347 1283 2356 1284
rect 2275 1278 2281 1279
rect 2347 1279 2348 1283
rect 2355 1279 2356 1283
rect 2398 1281 2399 1285
rect 2403 1281 2404 1285
rect 2398 1280 2404 1281
rect 2419 1285 2425 1286
rect 2419 1281 2420 1285
rect 2424 1281 2425 1285
rect 2419 1280 2425 1281
rect 2454 1285 2460 1286
rect 2454 1281 2455 1285
rect 2459 1281 2460 1285
rect 2502 1284 2508 1285
rect 2454 1280 2460 1281
rect 2462 1283 2468 1284
rect 2347 1278 2356 1279
rect 2462 1279 2463 1283
rect 2467 1282 2468 1283
rect 2475 1283 2481 1284
rect 2475 1282 2476 1283
rect 2467 1280 2476 1282
rect 2467 1279 2468 1280
rect 2462 1278 2468 1279
rect 2475 1279 2476 1280
rect 2480 1279 2481 1283
rect 2502 1280 2503 1284
rect 2507 1280 2508 1284
rect 2502 1279 2508 1280
rect 2475 1278 2481 1279
rect 446 1275 452 1276
rect 446 1274 447 1275
rect 196 1272 447 1274
rect 196 1270 198 1272
rect 446 1271 447 1272
rect 451 1271 452 1275
rect 446 1270 452 1271
rect 195 1269 201 1270
rect 195 1265 196 1269
rect 200 1265 201 1269
rect 251 1267 257 1268
rect 251 1266 252 1267
rect 195 1264 201 1265
rect 232 1264 252 1266
rect 232 1258 234 1264
rect 251 1263 252 1264
rect 256 1263 257 1267
rect 251 1262 257 1263
rect 307 1267 313 1268
rect 307 1263 308 1267
rect 312 1263 313 1267
rect 371 1267 377 1268
rect 371 1266 372 1267
rect 307 1262 313 1263
rect 325 1264 372 1266
rect 309 1258 311 1262
rect 212 1256 234 1258
rect 268 1256 311 1258
rect 212 1254 214 1256
rect 268 1254 270 1256
rect 325 1254 327 1264
rect 371 1263 372 1264
rect 376 1263 377 1267
rect 443 1267 449 1268
rect 443 1266 444 1267
rect 371 1262 377 1263
rect 388 1264 444 1266
rect 388 1254 390 1264
rect 443 1263 444 1264
rect 448 1263 449 1267
rect 443 1262 449 1263
rect 531 1267 537 1268
rect 531 1263 532 1267
rect 536 1263 537 1267
rect 531 1262 537 1263
rect 643 1267 649 1268
rect 643 1263 644 1267
rect 648 1266 649 1267
rect 654 1267 660 1268
rect 654 1266 655 1267
rect 648 1264 655 1266
rect 648 1263 649 1264
rect 643 1262 649 1263
rect 654 1263 655 1264
rect 659 1263 660 1267
rect 779 1267 785 1268
rect 779 1266 780 1267
rect 654 1262 660 1263
rect 664 1264 780 1266
rect 533 1258 535 1262
rect 664 1258 666 1264
rect 779 1263 780 1264
rect 784 1263 785 1267
rect 931 1267 937 1268
rect 931 1266 932 1267
rect 779 1262 785 1263
rect 796 1264 932 1266
rect 460 1256 535 1258
rect 660 1256 666 1258
rect 460 1254 462 1256
rect 660 1254 662 1256
rect 796 1254 798 1264
rect 931 1263 932 1264
rect 936 1263 937 1267
rect 1099 1267 1105 1268
rect 1099 1266 1100 1267
rect 931 1262 937 1263
rect 949 1264 1100 1266
rect 949 1254 951 1264
rect 1099 1263 1100 1264
rect 1104 1263 1105 1267
rect 1099 1262 1105 1263
rect 1243 1267 1252 1268
rect 1243 1263 1244 1267
rect 1251 1263 1252 1267
rect 1243 1262 1252 1263
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1263 1332 1267
rect 2502 1267 2508 1268
rect 1326 1262 1332 1263
rect 1350 1264 1356 1265
rect 1350 1260 1351 1264
rect 1355 1260 1356 1264
rect 1350 1259 1356 1260
rect 1406 1264 1412 1265
rect 1406 1260 1407 1264
rect 1411 1260 1412 1264
rect 1406 1259 1412 1260
rect 1502 1264 1508 1265
rect 1502 1260 1503 1264
rect 1507 1260 1508 1264
rect 1502 1259 1508 1260
rect 1598 1264 1604 1265
rect 1598 1260 1599 1264
rect 1603 1260 1604 1264
rect 1598 1259 1604 1260
rect 1702 1264 1708 1265
rect 1702 1260 1703 1264
rect 1707 1260 1708 1264
rect 1702 1259 1708 1260
rect 1806 1264 1812 1265
rect 1806 1260 1807 1264
rect 1811 1260 1812 1264
rect 1806 1259 1812 1260
rect 1902 1264 1908 1265
rect 1902 1260 1903 1264
rect 1907 1260 1908 1264
rect 1902 1259 1908 1260
rect 1998 1264 2004 1265
rect 1998 1260 1999 1264
rect 2003 1260 2004 1264
rect 1998 1259 2004 1260
rect 2086 1264 2092 1265
rect 2086 1260 2087 1264
rect 2091 1260 2092 1264
rect 2086 1259 2092 1260
rect 2166 1264 2172 1265
rect 2166 1260 2167 1264
rect 2171 1260 2172 1264
rect 2166 1259 2172 1260
rect 2238 1264 2244 1265
rect 2238 1260 2239 1264
rect 2243 1260 2244 1264
rect 2238 1259 2244 1260
rect 2310 1264 2316 1265
rect 2310 1260 2311 1264
rect 2315 1260 2316 1264
rect 2310 1259 2316 1260
rect 2382 1264 2388 1265
rect 2382 1260 2383 1264
rect 2387 1260 2388 1264
rect 2382 1259 2388 1260
rect 2438 1264 2444 1265
rect 2438 1260 2439 1264
rect 2443 1260 2444 1264
rect 2502 1263 2503 1267
rect 2507 1263 2508 1267
rect 2502 1262 2508 1263
rect 2438 1259 2444 1260
rect 190 1253 196 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 190 1249 191 1253
rect 195 1249 196 1253
rect 190 1248 196 1249
rect 211 1253 217 1254
rect 211 1249 212 1253
rect 216 1249 217 1253
rect 211 1248 217 1249
rect 246 1253 252 1254
rect 246 1249 247 1253
rect 251 1249 252 1253
rect 246 1248 252 1249
rect 267 1253 273 1254
rect 267 1249 268 1253
rect 272 1249 273 1253
rect 267 1248 273 1249
rect 302 1253 308 1254
rect 302 1249 303 1253
rect 307 1249 308 1253
rect 302 1248 308 1249
rect 323 1253 329 1254
rect 323 1249 324 1253
rect 328 1249 329 1253
rect 323 1248 329 1249
rect 366 1253 372 1254
rect 366 1249 367 1253
rect 371 1249 372 1253
rect 366 1248 372 1249
rect 387 1253 393 1254
rect 387 1249 388 1253
rect 392 1249 393 1253
rect 387 1248 393 1249
rect 438 1253 444 1254
rect 438 1249 439 1253
rect 443 1249 444 1253
rect 438 1248 444 1249
rect 459 1253 465 1254
rect 459 1249 460 1253
rect 464 1249 465 1253
rect 459 1248 465 1249
rect 526 1253 532 1254
rect 526 1249 527 1253
rect 531 1249 532 1253
rect 638 1253 644 1254
rect 526 1248 532 1249
rect 547 1251 556 1252
rect 110 1247 116 1248
rect 547 1247 548 1251
rect 555 1247 556 1251
rect 638 1249 639 1253
rect 643 1249 644 1253
rect 638 1248 644 1249
rect 659 1253 665 1254
rect 659 1249 660 1253
rect 664 1249 665 1253
rect 659 1248 665 1249
rect 774 1253 780 1254
rect 774 1249 775 1253
rect 779 1249 780 1253
rect 774 1248 780 1249
rect 795 1253 801 1254
rect 795 1249 796 1253
rect 800 1249 801 1253
rect 795 1248 801 1249
rect 926 1253 932 1254
rect 926 1249 927 1253
rect 931 1249 932 1253
rect 926 1248 932 1249
rect 947 1253 953 1254
rect 947 1249 948 1253
rect 952 1249 953 1253
rect 947 1248 953 1249
rect 1094 1253 1100 1254
rect 1094 1249 1095 1253
rect 1099 1249 1100 1253
rect 1238 1253 1244 1254
rect 1094 1248 1100 1249
rect 1114 1251 1121 1252
rect 547 1246 556 1247
rect 1114 1247 1115 1251
rect 1120 1247 1121 1251
rect 1238 1249 1239 1253
rect 1243 1249 1244 1253
rect 1286 1252 1292 1253
rect 1238 1248 1244 1249
rect 1259 1251 1265 1252
rect 1114 1246 1121 1247
rect 1259 1247 1260 1251
rect 1264 1250 1265 1251
rect 1278 1251 1284 1252
rect 1278 1250 1279 1251
rect 1264 1248 1279 1250
rect 1264 1247 1265 1248
rect 1259 1246 1265 1247
rect 1278 1247 1279 1248
rect 1283 1247 1284 1251
rect 1286 1248 1287 1252
rect 1291 1248 1292 1252
rect 1286 1247 1292 1248
rect 1278 1246 1284 1247
rect 1350 1236 1356 1237
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 1286 1235 1292 1236
rect 110 1230 116 1231
rect 174 1232 180 1233
rect 174 1228 175 1232
rect 179 1228 180 1232
rect 174 1227 180 1228
rect 230 1232 236 1233
rect 230 1228 231 1232
rect 235 1228 236 1232
rect 230 1227 236 1228
rect 286 1232 292 1233
rect 286 1228 287 1232
rect 291 1228 292 1232
rect 286 1227 292 1228
rect 350 1232 356 1233
rect 350 1228 351 1232
rect 355 1228 356 1232
rect 350 1227 356 1228
rect 422 1232 428 1233
rect 422 1228 423 1232
rect 427 1228 428 1232
rect 422 1227 428 1228
rect 510 1232 516 1233
rect 510 1228 511 1232
rect 515 1228 516 1232
rect 510 1227 516 1228
rect 622 1232 628 1233
rect 622 1228 623 1232
rect 627 1228 628 1232
rect 622 1227 628 1228
rect 758 1232 764 1233
rect 758 1228 759 1232
rect 763 1228 764 1232
rect 758 1227 764 1228
rect 910 1232 916 1233
rect 910 1228 911 1232
rect 915 1228 916 1232
rect 910 1227 916 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1222 1232 1228 1233
rect 1222 1228 1223 1232
rect 1227 1228 1228 1232
rect 1286 1231 1287 1235
rect 1291 1231 1292 1235
rect 1286 1230 1292 1231
rect 1326 1233 1332 1234
rect 1326 1229 1327 1233
rect 1331 1229 1332 1233
rect 1350 1232 1351 1236
rect 1355 1232 1356 1236
rect 1350 1231 1356 1232
rect 1446 1236 1452 1237
rect 1446 1232 1447 1236
rect 1451 1232 1452 1236
rect 1446 1231 1452 1232
rect 1574 1236 1580 1237
rect 1574 1232 1575 1236
rect 1579 1232 1580 1236
rect 1574 1231 1580 1232
rect 1694 1236 1700 1237
rect 1694 1232 1695 1236
rect 1699 1232 1700 1236
rect 1694 1231 1700 1232
rect 1814 1236 1820 1237
rect 1814 1232 1815 1236
rect 1819 1232 1820 1236
rect 1814 1231 1820 1232
rect 1926 1236 1932 1237
rect 1926 1232 1927 1236
rect 1931 1232 1932 1236
rect 1926 1231 1932 1232
rect 2030 1236 2036 1237
rect 2030 1232 2031 1236
rect 2035 1232 2036 1236
rect 2030 1231 2036 1232
rect 2126 1236 2132 1237
rect 2126 1232 2127 1236
rect 2131 1232 2132 1236
rect 2126 1231 2132 1232
rect 2214 1236 2220 1237
rect 2214 1232 2215 1236
rect 2219 1232 2220 1236
rect 2214 1231 2220 1232
rect 2294 1236 2300 1237
rect 2294 1232 2295 1236
rect 2299 1232 2300 1236
rect 2294 1231 2300 1232
rect 2374 1236 2380 1237
rect 2374 1232 2375 1236
rect 2379 1232 2380 1236
rect 2374 1231 2380 1232
rect 2438 1236 2444 1237
rect 2438 1232 2439 1236
rect 2443 1232 2444 1236
rect 2438 1231 2444 1232
rect 2502 1233 2508 1234
rect 1326 1228 1332 1229
rect 2502 1229 2503 1233
rect 2507 1229 2508 1233
rect 2502 1228 2508 1229
rect 1222 1227 1228 1228
rect 350 1220 356 1221
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 350 1216 351 1220
rect 355 1216 356 1220
rect 350 1215 356 1216
rect 406 1220 412 1221
rect 406 1216 407 1220
rect 411 1216 412 1220
rect 406 1215 412 1216
rect 462 1220 468 1221
rect 462 1216 463 1220
rect 467 1216 468 1220
rect 462 1215 468 1216
rect 518 1220 524 1221
rect 518 1216 519 1220
rect 523 1216 524 1220
rect 518 1215 524 1216
rect 574 1220 580 1221
rect 574 1216 575 1220
rect 579 1216 580 1220
rect 574 1215 580 1216
rect 630 1220 636 1221
rect 630 1216 631 1220
rect 635 1216 636 1220
rect 630 1215 636 1216
rect 686 1220 692 1221
rect 686 1216 687 1220
rect 691 1216 692 1220
rect 686 1215 692 1216
rect 742 1220 748 1221
rect 742 1216 743 1220
rect 747 1216 748 1220
rect 742 1215 748 1216
rect 798 1220 804 1221
rect 798 1216 799 1220
rect 803 1216 804 1220
rect 798 1215 804 1216
rect 854 1220 860 1221
rect 854 1216 855 1220
rect 859 1216 860 1220
rect 854 1215 860 1216
rect 910 1220 916 1221
rect 910 1216 911 1220
rect 915 1216 916 1220
rect 910 1215 916 1216
rect 1286 1217 1292 1218
rect 110 1212 116 1213
rect 1286 1213 1287 1217
rect 1291 1213 1292 1217
rect 1286 1212 1292 1213
rect 1326 1216 1332 1217
rect 2502 1216 2508 1217
rect 1326 1212 1327 1216
rect 1331 1212 1332 1216
rect 1326 1211 1332 1212
rect 1366 1215 1372 1216
rect 1366 1211 1367 1215
rect 1371 1211 1372 1215
rect 1366 1210 1372 1211
rect 1387 1215 1393 1216
rect 1387 1211 1388 1215
rect 1392 1211 1393 1215
rect 1387 1210 1393 1211
rect 1462 1215 1468 1216
rect 1462 1211 1463 1215
rect 1467 1211 1468 1215
rect 1462 1210 1468 1211
rect 1478 1215 1489 1216
rect 1478 1211 1479 1215
rect 1483 1211 1484 1215
rect 1488 1211 1489 1215
rect 1478 1210 1489 1211
rect 1590 1215 1596 1216
rect 1590 1211 1591 1215
rect 1595 1211 1596 1215
rect 1590 1210 1596 1211
rect 1611 1215 1617 1216
rect 1611 1211 1612 1215
rect 1616 1214 1617 1215
rect 1710 1215 1716 1216
rect 1616 1212 1706 1214
rect 1616 1211 1617 1212
rect 1611 1210 1617 1211
rect 1278 1207 1284 1208
rect 1278 1203 1279 1207
rect 1283 1206 1284 1207
rect 1283 1204 1374 1206
rect 1283 1203 1284 1204
rect 1278 1202 1284 1203
rect 1372 1202 1374 1204
rect 1389 1202 1391 1210
rect 1704 1202 1706 1212
rect 1710 1211 1711 1215
rect 1715 1211 1716 1215
rect 1710 1210 1716 1211
rect 1731 1215 1737 1216
rect 1731 1211 1732 1215
rect 1736 1214 1737 1215
rect 1830 1215 1836 1216
rect 1736 1212 1826 1214
rect 1736 1211 1737 1212
rect 1731 1210 1737 1211
rect 1824 1202 1826 1212
rect 1830 1211 1831 1215
rect 1835 1211 1836 1215
rect 1830 1210 1836 1211
rect 1850 1215 1857 1216
rect 1850 1211 1851 1215
rect 1856 1211 1857 1215
rect 1850 1210 1857 1211
rect 1942 1215 1948 1216
rect 1942 1211 1943 1215
rect 1947 1211 1948 1215
rect 1942 1210 1948 1211
rect 1963 1215 1969 1216
rect 1963 1211 1964 1215
rect 1968 1214 1969 1215
rect 2046 1215 2052 1216
rect 1968 1212 2001 1214
rect 1968 1211 1969 1212
rect 1963 1210 1969 1211
rect 1999 1202 2001 1212
rect 2046 1211 2047 1215
rect 2051 1211 2052 1215
rect 2046 1210 2052 1211
rect 2067 1215 2073 1216
rect 2067 1211 2068 1215
rect 2072 1211 2073 1215
rect 2067 1210 2073 1211
rect 2142 1215 2148 1216
rect 2142 1211 2143 1215
rect 2147 1211 2148 1215
rect 2142 1210 2148 1211
rect 2163 1215 2169 1216
rect 2163 1211 2164 1215
rect 2168 1214 2169 1215
rect 2230 1215 2236 1216
rect 2168 1212 2222 1214
rect 2168 1211 2169 1212
rect 2163 1210 2169 1211
rect 2069 1202 2071 1210
rect 2220 1202 2222 1212
rect 2230 1211 2231 1215
rect 2235 1211 2236 1215
rect 2230 1210 2236 1211
rect 2251 1215 2257 1216
rect 2251 1211 2252 1215
rect 2256 1214 2257 1215
rect 2310 1215 2316 1216
rect 2256 1212 2306 1214
rect 2256 1211 2257 1212
rect 2251 1210 2257 1211
rect 2304 1202 2306 1212
rect 2310 1211 2311 1215
rect 2315 1211 2316 1215
rect 2310 1210 2316 1211
rect 2331 1215 2337 1216
rect 2331 1211 2332 1215
rect 2336 1214 2337 1215
rect 2374 1215 2380 1216
rect 2374 1214 2375 1215
rect 2336 1212 2375 1214
rect 2336 1211 2337 1212
rect 2331 1210 2337 1211
rect 2374 1211 2375 1212
rect 2379 1211 2380 1215
rect 2374 1210 2380 1211
rect 2390 1215 2396 1216
rect 2390 1211 2391 1215
rect 2395 1211 2396 1215
rect 2390 1210 2396 1211
rect 2410 1215 2417 1216
rect 2410 1211 2411 1215
rect 2416 1211 2417 1215
rect 2410 1210 2417 1211
rect 2454 1215 2460 1216
rect 2454 1211 2455 1215
rect 2459 1211 2460 1215
rect 2454 1210 2460 1211
rect 2470 1215 2481 1216
rect 2470 1211 2471 1215
rect 2475 1211 2476 1215
rect 2480 1211 2481 1215
rect 2502 1212 2503 1216
rect 2507 1212 2508 1216
rect 2502 1211 2508 1212
rect 2470 1210 2481 1211
rect 1371 1201 1377 1202
rect 110 1200 116 1201
rect 1286 1200 1292 1201
rect 110 1196 111 1200
rect 115 1196 116 1200
rect 110 1195 116 1196
rect 366 1199 372 1200
rect 366 1195 367 1199
rect 371 1195 372 1199
rect 366 1194 372 1195
rect 387 1199 393 1200
rect 387 1195 388 1199
rect 392 1198 393 1199
rect 422 1199 428 1200
rect 392 1196 418 1198
rect 392 1195 393 1196
rect 387 1194 393 1195
rect 416 1186 418 1196
rect 422 1195 423 1199
rect 427 1195 428 1199
rect 422 1194 428 1195
rect 443 1199 449 1200
rect 443 1195 444 1199
rect 448 1198 449 1199
rect 478 1199 484 1200
rect 448 1196 474 1198
rect 448 1195 449 1196
rect 443 1194 449 1195
rect 472 1186 474 1196
rect 478 1195 479 1199
rect 483 1195 484 1199
rect 478 1194 484 1195
rect 499 1199 505 1200
rect 499 1195 500 1199
rect 504 1198 505 1199
rect 534 1199 540 1200
rect 504 1196 526 1198
rect 504 1195 505 1196
rect 499 1194 505 1195
rect 524 1186 526 1196
rect 534 1195 535 1199
rect 539 1195 540 1199
rect 534 1194 540 1195
rect 555 1199 561 1200
rect 555 1195 556 1199
rect 560 1198 561 1199
rect 590 1199 596 1200
rect 560 1196 586 1198
rect 560 1195 561 1196
rect 555 1194 561 1195
rect 584 1186 586 1196
rect 590 1195 591 1199
rect 595 1195 596 1199
rect 590 1194 596 1195
rect 611 1199 617 1200
rect 611 1195 612 1199
rect 616 1198 617 1199
rect 638 1199 644 1200
rect 638 1198 639 1199
rect 616 1196 639 1198
rect 616 1195 617 1196
rect 611 1194 617 1195
rect 638 1195 639 1196
rect 643 1195 644 1199
rect 638 1194 644 1195
rect 646 1199 652 1200
rect 646 1195 647 1199
rect 651 1195 652 1199
rect 646 1194 652 1195
rect 654 1199 660 1200
rect 654 1195 655 1199
rect 659 1198 660 1199
rect 667 1199 673 1200
rect 667 1198 668 1199
rect 659 1196 668 1198
rect 659 1195 660 1196
rect 654 1194 660 1195
rect 667 1195 668 1196
rect 672 1195 673 1199
rect 667 1194 673 1195
rect 702 1199 708 1200
rect 702 1195 703 1199
rect 707 1195 708 1199
rect 723 1199 729 1200
rect 723 1198 724 1199
rect 702 1194 708 1195
rect 712 1196 724 1198
rect 712 1190 714 1196
rect 723 1195 724 1196
rect 728 1195 729 1199
rect 723 1194 729 1195
rect 758 1199 764 1200
rect 758 1195 759 1199
rect 763 1195 764 1199
rect 758 1194 764 1195
rect 774 1199 785 1200
rect 774 1195 775 1199
rect 779 1195 780 1199
rect 784 1195 785 1199
rect 774 1194 785 1195
rect 814 1199 820 1200
rect 814 1195 815 1199
rect 819 1195 820 1199
rect 814 1194 820 1195
rect 835 1199 841 1200
rect 835 1195 836 1199
rect 840 1195 841 1199
rect 835 1194 841 1195
rect 870 1199 876 1200
rect 870 1195 871 1199
rect 875 1195 876 1199
rect 870 1194 876 1195
rect 886 1199 897 1200
rect 886 1195 887 1199
rect 891 1195 892 1199
rect 896 1195 897 1199
rect 886 1194 897 1195
rect 926 1199 932 1200
rect 926 1195 927 1199
rect 931 1195 932 1199
rect 926 1194 932 1195
rect 947 1199 953 1200
rect 947 1195 948 1199
rect 952 1195 953 1199
rect 1286 1196 1287 1200
rect 1291 1196 1292 1200
rect 1371 1197 1372 1201
rect 1376 1197 1377 1201
rect 1389 1201 1473 1202
rect 1389 1200 1468 1201
rect 1371 1196 1377 1197
rect 1467 1197 1468 1200
rect 1472 1197 1473 1201
rect 1704 1201 1721 1202
rect 1704 1200 1716 1201
rect 1467 1196 1473 1197
rect 1595 1199 1601 1200
rect 1286 1195 1292 1196
rect 1595 1195 1596 1199
rect 1600 1198 1601 1199
rect 1600 1196 1710 1198
rect 1715 1197 1716 1200
rect 1720 1197 1721 1201
rect 1824 1201 1841 1202
rect 1824 1200 1836 1201
rect 1715 1196 1721 1197
rect 1835 1197 1836 1200
rect 1840 1197 1841 1201
rect 1999 1201 2057 1202
rect 1999 1200 2052 1201
rect 1835 1196 1841 1197
rect 1947 1199 1956 1200
rect 1600 1195 1601 1196
rect 947 1194 953 1195
rect 1595 1194 1601 1195
rect 1708 1194 1710 1196
rect 1754 1195 1760 1196
rect 1754 1194 1755 1195
rect 837 1190 839 1194
rect 949 1190 951 1194
rect 1708 1192 1755 1194
rect 1754 1191 1755 1192
rect 1759 1191 1760 1195
rect 1947 1195 1948 1199
rect 1955 1195 1956 1199
rect 2051 1197 2052 1200
rect 2056 1197 2057 1201
rect 2069 1201 2153 1202
rect 2069 1200 2148 1201
rect 2051 1196 2057 1197
rect 2147 1197 2148 1200
rect 2152 1197 2153 1201
rect 2220 1201 2241 1202
rect 2220 1200 2236 1201
rect 2147 1196 2153 1197
rect 2235 1197 2236 1200
rect 2240 1197 2241 1201
rect 2304 1201 2321 1202
rect 2304 1200 2316 1201
rect 2235 1196 2241 1197
rect 2315 1197 2316 1200
rect 2320 1197 2321 1201
rect 2315 1196 2321 1197
rect 2395 1199 2401 1200
rect 1947 1194 1956 1195
rect 2395 1195 2396 1199
rect 2400 1198 2401 1199
rect 2434 1199 2440 1200
rect 2434 1198 2435 1199
rect 2400 1196 2435 1198
rect 2400 1195 2401 1196
rect 2395 1194 2401 1195
rect 2434 1195 2435 1196
rect 2439 1195 2440 1199
rect 2434 1194 2440 1195
rect 2459 1199 2468 1200
rect 2459 1195 2460 1199
rect 2467 1195 2468 1199
rect 2459 1194 2468 1195
rect 1754 1190 1760 1191
rect 652 1188 714 1190
rect 764 1188 839 1190
rect 876 1188 951 1190
rect 652 1186 654 1188
rect 764 1186 766 1188
rect 876 1186 878 1188
rect 1478 1187 1484 1188
rect 1478 1186 1479 1187
rect 416 1185 433 1186
rect 416 1184 428 1185
rect 371 1183 377 1184
rect 371 1179 372 1183
rect 376 1182 377 1183
rect 376 1180 423 1182
rect 427 1181 428 1184
rect 432 1181 433 1185
rect 472 1185 489 1186
rect 472 1184 484 1185
rect 427 1180 433 1181
rect 483 1181 484 1184
rect 488 1181 489 1185
rect 524 1185 545 1186
rect 524 1184 540 1185
rect 483 1180 489 1181
rect 539 1181 540 1184
rect 544 1181 545 1185
rect 584 1185 601 1186
rect 584 1184 596 1185
rect 539 1180 545 1181
rect 595 1181 596 1184
rect 600 1181 601 1185
rect 595 1180 601 1181
rect 651 1185 657 1186
rect 651 1181 652 1185
rect 656 1181 657 1185
rect 763 1185 769 1186
rect 651 1180 657 1181
rect 707 1183 713 1184
rect 376 1179 377 1180
rect 371 1178 377 1179
rect 421 1178 423 1180
rect 550 1179 556 1180
rect 550 1178 551 1179
rect 421 1176 551 1178
rect 550 1175 551 1176
rect 555 1175 556 1179
rect 707 1179 708 1183
rect 712 1182 713 1183
rect 712 1180 746 1182
rect 763 1181 764 1185
rect 768 1181 769 1185
rect 875 1185 881 1186
rect 763 1180 769 1181
rect 819 1183 825 1184
rect 712 1179 713 1180
rect 707 1178 713 1179
rect 744 1178 746 1180
rect 774 1179 780 1180
rect 774 1178 775 1179
rect 744 1176 775 1178
rect 550 1174 556 1175
rect 774 1175 775 1176
rect 779 1175 780 1179
rect 819 1179 820 1183
rect 824 1179 825 1183
rect 875 1181 876 1185
rect 880 1181 881 1185
rect 1372 1184 1479 1186
rect 875 1180 881 1181
rect 894 1183 900 1184
rect 819 1178 825 1179
rect 886 1179 892 1180
rect 886 1178 887 1179
rect 821 1176 887 1178
rect 774 1174 780 1175
rect 886 1175 887 1176
rect 891 1175 892 1179
rect 894 1179 895 1183
rect 899 1182 900 1183
rect 931 1183 937 1184
rect 931 1182 932 1183
rect 899 1180 932 1182
rect 899 1179 900 1180
rect 894 1178 900 1179
rect 931 1179 932 1180
rect 936 1179 937 1183
rect 1372 1182 1374 1184
rect 1478 1183 1479 1184
rect 1483 1183 1484 1187
rect 2210 1187 2216 1188
rect 2210 1186 2211 1187
rect 1478 1182 1484 1183
rect 1988 1184 2211 1186
rect 1988 1182 1990 1184
rect 2210 1183 2211 1184
rect 2215 1183 2216 1187
rect 2210 1182 2216 1183
rect 931 1178 937 1179
rect 1371 1181 1377 1182
rect 1371 1177 1372 1181
rect 1376 1177 1377 1181
rect 1987 1181 1993 1182
rect 1371 1176 1377 1177
rect 1475 1179 1481 1180
rect 886 1174 892 1175
rect 1475 1175 1476 1179
rect 1480 1175 1481 1179
rect 1603 1179 1609 1180
rect 1603 1178 1604 1179
rect 1475 1174 1481 1175
rect 1548 1176 1604 1178
rect 1477 1170 1479 1174
rect 1389 1168 1479 1170
rect 722 1167 728 1168
rect 722 1166 723 1167
rect 428 1164 590 1166
rect 428 1162 430 1164
rect 427 1161 433 1162
rect 427 1157 428 1161
rect 432 1157 433 1161
rect 483 1159 489 1160
rect 483 1158 484 1159
rect 427 1156 433 1157
rect 444 1156 484 1158
rect 444 1146 446 1156
rect 483 1155 484 1156
rect 488 1155 489 1159
rect 539 1159 545 1160
rect 539 1158 540 1159
rect 483 1154 489 1155
rect 500 1156 540 1158
rect 500 1146 502 1156
rect 539 1155 540 1156
rect 544 1155 545 1159
rect 539 1154 545 1155
rect 588 1150 590 1164
rect 596 1164 723 1166
rect 596 1162 598 1164
rect 722 1163 723 1164
rect 727 1163 728 1167
rect 1002 1167 1008 1168
rect 1002 1166 1003 1167
rect 722 1162 728 1163
rect 764 1164 1003 1166
rect 764 1162 766 1164
rect 1002 1163 1003 1164
rect 1007 1163 1008 1167
rect 1389 1166 1391 1168
rect 1548 1166 1550 1176
rect 1603 1175 1604 1176
rect 1608 1175 1609 1179
rect 1603 1174 1609 1175
rect 1739 1179 1745 1180
rect 1739 1175 1740 1179
rect 1744 1175 1745 1179
rect 1739 1174 1745 1175
rect 1854 1179 1860 1180
rect 1854 1175 1855 1179
rect 1859 1178 1860 1179
rect 1867 1179 1873 1180
rect 1867 1178 1868 1179
rect 1859 1176 1868 1178
rect 1859 1175 1860 1176
rect 1854 1174 1860 1175
rect 1867 1175 1868 1176
rect 1872 1175 1873 1179
rect 1987 1177 1988 1181
rect 1992 1177 1993 1181
rect 1987 1176 1993 1177
rect 2091 1179 2097 1180
rect 1867 1174 1873 1175
rect 2091 1175 2092 1179
rect 2096 1175 2097 1179
rect 2091 1174 2097 1175
rect 2195 1179 2201 1180
rect 2195 1175 2196 1179
rect 2200 1178 2201 1179
rect 2291 1179 2297 1180
rect 2200 1176 2282 1178
rect 2200 1175 2201 1176
rect 2195 1174 2201 1175
rect 1741 1170 1743 1174
rect 2093 1170 2095 1174
rect 1741 1168 1886 1170
rect 1884 1166 1886 1168
rect 2005 1168 2095 1170
rect 2280 1170 2282 1176
rect 2291 1175 2292 1179
rect 2296 1178 2297 1179
rect 2374 1179 2380 1180
rect 2296 1176 2370 1178
rect 2296 1175 2297 1176
rect 2291 1174 2297 1175
rect 2368 1170 2370 1176
rect 2374 1175 2375 1179
rect 2379 1178 2380 1179
rect 2387 1179 2393 1180
rect 2387 1178 2388 1179
rect 2379 1176 2388 1178
rect 2379 1175 2380 1176
rect 2374 1174 2380 1175
rect 2387 1175 2388 1176
rect 2392 1175 2393 1179
rect 2387 1174 2393 1175
rect 2459 1179 2465 1180
rect 2459 1175 2460 1179
rect 2464 1178 2465 1179
rect 2478 1179 2484 1180
rect 2478 1178 2479 1179
rect 2464 1176 2479 1178
rect 2464 1175 2465 1176
rect 2459 1174 2465 1175
rect 2478 1175 2479 1176
rect 2483 1175 2484 1179
rect 2478 1174 2484 1175
rect 2434 1171 2440 1172
rect 2280 1168 2310 1170
rect 2368 1168 2406 1170
rect 2005 1166 2007 1168
rect 2308 1166 2310 1168
rect 2404 1166 2406 1168
rect 2434 1167 2435 1171
rect 2439 1170 2440 1171
rect 2439 1168 2479 1170
rect 2439 1167 2440 1168
rect 2434 1166 2440 1167
rect 2477 1166 2479 1168
rect 1366 1165 1372 1166
rect 1002 1162 1008 1163
rect 1326 1164 1332 1165
rect 595 1161 601 1162
rect 595 1157 596 1161
rect 600 1157 601 1161
rect 763 1161 769 1162
rect 595 1156 601 1157
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1158 644 1159
rect 651 1159 657 1160
rect 651 1158 652 1159
rect 643 1156 652 1158
rect 643 1155 644 1156
rect 638 1154 644 1155
rect 651 1155 652 1156
rect 656 1155 657 1159
rect 707 1159 713 1160
rect 707 1158 708 1159
rect 651 1154 657 1155
rect 668 1156 708 1158
rect 588 1148 615 1150
rect 613 1146 615 1148
rect 668 1146 670 1156
rect 707 1155 708 1156
rect 712 1155 713 1159
rect 763 1157 764 1161
rect 768 1157 769 1161
rect 1326 1160 1327 1164
rect 1331 1160 1332 1164
rect 1366 1161 1367 1165
rect 1371 1161 1372 1165
rect 1366 1160 1372 1161
rect 1387 1165 1393 1166
rect 1387 1161 1388 1165
rect 1392 1161 1393 1165
rect 1387 1160 1393 1161
rect 1470 1165 1476 1166
rect 1470 1161 1471 1165
rect 1475 1161 1476 1165
rect 1470 1160 1476 1161
rect 1491 1165 1550 1166
rect 1491 1161 1492 1165
rect 1496 1164 1550 1165
rect 1598 1165 1604 1166
rect 1496 1161 1497 1164
rect 1491 1160 1497 1161
rect 1598 1161 1599 1165
rect 1603 1161 1604 1165
rect 1734 1165 1740 1166
rect 1598 1160 1604 1161
rect 1606 1163 1612 1164
rect 763 1156 769 1157
rect 819 1159 825 1160
rect 707 1154 713 1155
rect 819 1155 820 1159
rect 824 1155 825 1159
rect 875 1159 881 1160
rect 875 1158 876 1159
rect 819 1154 825 1155
rect 837 1156 876 1158
rect 821 1150 823 1154
rect 780 1148 823 1150
rect 780 1146 782 1148
rect 837 1146 839 1156
rect 875 1155 876 1156
rect 880 1155 881 1159
rect 875 1154 881 1155
rect 886 1159 892 1160
rect 886 1155 887 1159
rect 891 1158 892 1159
rect 931 1159 937 1160
rect 931 1158 932 1159
rect 891 1156 932 1158
rect 891 1155 892 1156
rect 886 1154 892 1155
rect 931 1155 932 1156
rect 936 1155 937 1159
rect 987 1159 993 1160
rect 1326 1159 1332 1160
rect 1606 1159 1607 1163
rect 1611 1162 1612 1163
rect 1619 1163 1625 1164
rect 1619 1162 1620 1163
rect 1611 1160 1620 1162
rect 1611 1159 1612 1160
rect 987 1158 988 1159
rect 931 1154 937 1155
rect 949 1156 988 1158
rect 949 1146 951 1156
rect 987 1155 988 1156
rect 992 1155 993 1159
rect 1606 1158 1612 1159
rect 1619 1159 1620 1160
rect 1624 1159 1625 1163
rect 1734 1161 1735 1165
rect 1739 1161 1740 1165
rect 1862 1165 1868 1166
rect 1734 1160 1740 1161
rect 1754 1163 1761 1164
rect 1619 1158 1625 1159
rect 1754 1159 1755 1163
rect 1760 1159 1761 1163
rect 1862 1161 1863 1165
rect 1867 1161 1868 1165
rect 1862 1160 1868 1161
rect 1883 1165 1889 1166
rect 1883 1161 1884 1165
rect 1888 1161 1889 1165
rect 1883 1160 1889 1161
rect 1982 1165 1988 1166
rect 1982 1161 1983 1165
rect 1987 1161 1988 1165
rect 1982 1160 1988 1161
rect 2003 1165 2009 1166
rect 2003 1161 2004 1165
rect 2008 1161 2009 1165
rect 2003 1160 2009 1161
rect 2086 1165 2092 1166
rect 2086 1161 2087 1165
rect 2091 1161 2092 1165
rect 2190 1165 2196 1166
rect 2086 1160 2092 1161
rect 2107 1163 2113 1164
rect 1754 1158 1761 1159
rect 2107 1159 2108 1163
rect 2112 1162 2113 1163
rect 2166 1163 2172 1164
rect 2166 1162 2167 1163
rect 2112 1160 2167 1162
rect 2112 1159 2113 1160
rect 2107 1158 2113 1159
rect 2166 1159 2167 1160
rect 2171 1159 2172 1163
rect 2190 1161 2191 1165
rect 2195 1161 2196 1165
rect 2286 1165 2292 1166
rect 2190 1160 2196 1161
rect 2210 1163 2217 1164
rect 2166 1158 2172 1159
rect 2210 1159 2211 1163
rect 2216 1159 2217 1163
rect 2286 1161 2287 1165
rect 2291 1161 2292 1165
rect 2286 1160 2292 1161
rect 2307 1165 2313 1166
rect 2307 1161 2308 1165
rect 2312 1161 2313 1165
rect 2307 1160 2313 1161
rect 2382 1165 2388 1166
rect 2382 1161 2383 1165
rect 2387 1161 2388 1165
rect 2382 1160 2388 1161
rect 2403 1165 2409 1166
rect 2403 1161 2404 1165
rect 2408 1161 2409 1165
rect 2403 1160 2409 1161
rect 2454 1165 2460 1166
rect 2454 1161 2455 1165
rect 2459 1161 2460 1165
rect 2454 1160 2460 1161
rect 2475 1165 2481 1166
rect 2475 1161 2476 1165
rect 2480 1161 2481 1165
rect 2475 1160 2481 1161
rect 2502 1164 2508 1165
rect 2502 1160 2503 1164
rect 2507 1160 2508 1164
rect 2502 1159 2508 1160
rect 2210 1158 2217 1159
rect 987 1154 993 1155
rect 1326 1147 1332 1148
rect 422 1145 428 1146
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 422 1141 423 1145
rect 427 1141 428 1145
rect 422 1140 428 1141
rect 443 1145 449 1146
rect 443 1141 444 1145
rect 448 1141 449 1145
rect 443 1140 449 1141
rect 478 1145 484 1146
rect 478 1141 479 1145
rect 483 1141 484 1145
rect 478 1140 484 1141
rect 499 1145 505 1146
rect 499 1141 500 1145
rect 504 1141 505 1145
rect 499 1140 505 1141
rect 534 1145 540 1146
rect 534 1141 535 1145
rect 539 1141 540 1145
rect 590 1145 596 1146
rect 534 1140 540 1141
rect 555 1143 561 1144
rect 110 1139 116 1140
rect 555 1139 556 1143
rect 560 1142 561 1143
rect 582 1143 588 1144
rect 582 1142 583 1143
rect 560 1140 583 1142
rect 560 1139 561 1140
rect 555 1138 561 1139
rect 582 1139 583 1140
rect 587 1139 588 1143
rect 590 1141 591 1145
rect 595 1141 596 1145
rect 590 1140 596 1141
rect 611 1145 617 1146
rect 611 1141 612 1145
rect 616 1141 617 1145
rect 611 1140 617 1141
rect 646 1145 652 1146
rect 646 1141 647 1145
rect 651 1141 652 1145
rect 646 1140 652 1141
rect 667 1145 673 1146
rect 667 1141 668 1145
rect 672 1141 673 1145
rect 667 1140 673 1141
rect 702 1145 708 1146
rect 702 1141 703 1145
rect 707 1141 708 1145
rect 758 1145 764 1146
rect 702 1140 708 1141
rect 722 1143 729 1144
rect 582 1138 588 1139
rect 722 1139 723 1143
rect 728 1139 729 1143
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 779 1145 785 1146
rect 779 1141 780 1145
rect 784 1141 785 1145
rect 779 1140 785 1141
rect 814 1145 820 1146
rect 814 1141 815 1145
rect 819 1141 820 1145
rect 814 1140 820 1141
rect 835 1145 841 1146
rect 835 1141 836 1145
rect 840 1141 841 1145
rect 835 1140 841 1141
rect 870 1145 876 1146
rect 870 1141 871 1145
rect 875 1141 876 1145
rect 926 1145 932 1146
rect 870 1140 876 1141
rect 891 1143 900 1144
rect 722 1138 729 1139
rect 891 1139 892 1143
rect 899 1139 900 1143
rect 926 1141 927 1145
rect 931 1141 932 1145
rect 926 1140 932 1141
rect 947 1145 953 1146
rect 947 1141 948 1145
rect 952 1141 953 1145
rect 947 1140 953 1141
rect 982 1145 988 1146
rect 982 1141 983 1145
rect 987 1141 988 1145
rect 1286 1144 1292 1145
rect 982 1140 988 1141
rect 1002 1143 1009 1144
rect 891 1138 900 1139
rect 1002 1139 1003 1143
rect 1008 1139 1009 1143
rect 1286 1140 1287 1144
rect 1291 1140 1292 1144
rect 1326 1143 1327 1147
rect 1331 1143 1332 1147
rect 2502 1147 2508 1148
rect 1326 1142 1332 1143
rect 1350 1144 1356 1145
rect 1286 1139 1292 1140
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1454 1144 1460 1145
rect 1454 1140 1455 1144
rect 1459 1140 1460 1144
rect 1454 1139 1460 1140
rect 1582 1144 1588 1145
rect 1582 1140 1583 1144
rect 1587 1140 1588 1144
rect 1582 1139 1588 1140
rect 1718 1144 1724 1145
rect 1718 1140 1719 1144
rect 1723 1140 1724 1144
rect 1718 1139 1724 1140
rect 1846 1144 1852 1145
rect 1846 1140 1847 1144
rect 1851 1140 1852 1144
rect 1846 1139 1852 1140
rect 1966 1144 1972 1145
rect 1966 1140 1967 1144
rect 1971 1140 1972 1144
rect 1966 1139 1972 1140
rect 2070 1144 2076 1145
rect 2070 1140 2071 1144
rect 2075 1140 2076 1144
rect 2070 1139 2076 1140
rect 2174 1144 2180 1145
rect 2174 1140 2175 1144
rect 2179 1140 2180 1144
rect 2174 1139 2180 1140
rect 2270 1144 2276 1145
rect 2270 1140 2271 1144
rect 2275 1140 2276 1144
rect 2270 1139 2276 1140
rect 2366 1144 2372 1145
rect 2366 1140 2367 1144
rect 2371 1140 2372 1144
rect 2366 1139 2372 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2502 1143 2503 1147
rect 2507 1143 2508 1147
rect 2502 1142 2508 1143
rect 2438 1139 2444 1140
rect 1002 1138 1009 1139
rect 1366 1128 1372 1129
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 1286 1127 1292 1128
rect 110 1122 116 1123
rect 406 1124 412 1125
rect 406 1120 407 1124
rect 411 1120 412 1124
rect 406 1119 412 1120
rect 462 1124 468 1125
rect 462 1120 463 1124
rect 467 1120 468 1124
rect 462 1119 468 1120
rect 518 1124 524 1125
rect 518 1120 519 1124
rect 523 1120 524 1124
rect 518 1119 524 1120
rect 574 1124 580 1125
rect 574 1120 575 1124
rect 579 1120 580 1124
rect 574 1119 580 1120
rect 630 1124 636 1125
rect 630 1120 631 1124
rect 635 1120 636 1124
rect 630 1119 636 1120
rect 686 1124 692 1125
rect 686 1120 687 1124
rect 691 1120 692 1124
rect 686 1119 692 1120
rect 742 1124 748 1125
rect 742 1120 743 1124
rect 747 1120 748 1124
rect 742 1119 748 1120
rect 798 1124 804 1125
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 798 1119 804 1120
rect 854 1124 860 1125
rect 854 1120 855 1124
rect 859 1120 860 1124
rect 854 1119 860 1120
rect 910 1124 916 1125
rect 910 1120 911 1124
rect 915 1120 916 1124
rect 910 1119 916 1120
rect 966 1124 972 1125
rect 966 1120 967 1124
rect 971 1120 972 1124
rect 1286 1123 1287 1127
rect 1291 1123 1292 1127
rect 1286 1122 1292 1123
rect 1326 1125 1332 1126
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1366 1124 1367 1128
rect 1371 1124 1372 1128
rect 1366 1123 1372 1124
rect 1446 1128 1452 1129
rect 1446 1124 1447 1128
rect 1451 1124 1452 1128
rect 1446 1123 1452 1124
rect 1534 1128 1540 1129
rect 1534 1124 1535 1128
rect 1539 1124 1540 1128
rect 1534 1123 1540 1124
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1806 1128 1812 1129
rect 1806 1124 1807 1128
rect 1811 1124 1812 1128
rect 1806 1123 1812 1124
rect 1894 1128 1900 1129
rect 1894 1124 1895 1128
rect 1899 1124 1900 1128
rect 1894 1123 1900 1124
rect 1982 1128 1988 1129
rect 1982 1124 1983 1128
rect 1987 1124 1988 1128
rect 1982 1123 1988 1124
rect 2070 1128 2076 1129
rect 2070 1124 2071 1128
rect 2075 1124 2076 1128
rect 2070 1123 2076 1124
rect 2158 1128 2164 1129
rect 2158 1124 2159 1128
rect 2163 1124 2164 1128
rect 2158 1123 2164 1124
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 2438 1128 2444 1129
rect 2438 1124 2439 1128
rect 2443 1124 2444 1128
rect 2438 1123 2444 1124
rect 2502 1125 2508 1126
rect 1326 1120 1332 1121
rect 2502 1121 2503 1125
rect 2507 1121 2508 1125
rect 2502 1120 2508 1121
rect 966 1119 972 1120
rect 222 1108 228 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 222 1104 223 1108
rect 227 1104 228 1108
rect 222 1103 228 1104
rect 310 1108 316 1109
rect 310 1104 311 1108
rect 315 1104 316 1108
rect 310 1103 316 1104
rect 398 1108 404 1109
rect 398 1104 399 1108
rect 403 1104 404 1108
rect 398 1103 404 1104
rect 494 1108 500 1109
rect 494 1104 495 1108
rect 499 1104 500 1108
rect 494 1103 500 1104
rect 590 1108 596 1109
rect 590 1104 591 1108
rect 595 1104 596 1108
rect 590 1103 596 1104
rect 678 1108 684 1109
rect 678 1104 679 1108
rect 683 1104 684 1108
rect 678 1103 684 1104
rect 766 1108 772 1109
rect 766 1104 767 1108
rect 771 1104 772 1108
rect 766 1103 772 1104
rect 846 1108 852 1109
rect 846 1104 847 1108
rect 851 1104 852 1108
rect 846 1103 852 1104
rect 926 1108 932 1109
rect 926 1104 927 1108
rect 931 1104 932 1108
rect 926 1103 932 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1102 1108 1108 1109
rect 1102 1104 1103 1108
rect 1107 1104 1108 1108
rect 1326 1108 1332 1109
rect 2502 1108 2508 1109
rect 1102 1103 1108 1104
rect 1286 1105 1292 1106
rect 110 1100 116 1101
rect 1286 1101 1287 1105
rect 1291 1101 1292 1105
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1326 1103 1332 1104
rect 1382 1107 1388 1108
rect 1382 1103 1383 1107
rect 1387 1103 1388 1107
rect 1382 1102 1388 1103
rect 1403 1107 1409 1108
rect 1403 1103 1404 1107
rect 1408 1106 1409 1107
rect 1422 1107 1428 1108
rect 1422 1106 1423 1107
rect 1408 1104 1423 1106
rect 1408 1103 1409 1104
rect 1403 1102 1409 1103
rect 1422 1103 1423 1104
rect 1427 1103 1428 1107
rect 1422 1102 1428 1103
rect 1462 1107 1468 1108
rect 1462 1103 1463 1107
rect 1467 1103 1468 1107
rect 1462 1102 1468 1103
rect 1478 1107 1489 1108
rect 1478 1103 1479 1107
rect 1483 1103 1484 1107
rect 1488 1103 1489 1107
rect 1478 1102 1489 1103
rect 1550 1107 1556 1108
rect 1550 1103 1551 1107
rect 1555 1103 1556 1107
rect 1571 1107 1577 1108
rect 1571 1106 1572 1107
rect 1550 1102 1556 1103
rect 1560 1104 1572 1106
rect 1286 1100 1292 1101
rect 1560 1098 1562 1104
rect 1571 1103 1572 1104
rect 1576 1103 1577 1107
rect 1571 1102 1577 1103
rect 1646 1107 1652 1108
rect 1646 1103 1647 1107
rect 1651 1103 1652 1107
rect 1646 1102 1652 1103
rect 1667 1107 1673 1108
rect 1667 1103 1668 1107
rect 1672 1106 1673 1107
rect 1734 1107 1740 1108
rect 1672 1104 1730 1106
rect 1672 1103 1673 1104
rect 1667 1102 1673 1103
rect 1468 1096 1562 1098
rect 1468 1094 1470 1096
rect 1728 1094 1730 1104
rect 1734 1103 1735 1107
rect 1739 1103 1740 1107
rect 1734 1102 1740 1103
rect 1755 1107 1761 1108
rect 1755 1103 1756 1107
rect 1760 1103 1761 1107
rect 1755 1102 1761 1103
rect 1822 1107 1828 1108
rect 1822 1103 1823 1107
rect 1827 1103 1828 1107
rect 1822 1102 1828 1103
rect 1843 1107 1849 1108
rect 1843 1103 1844 1107
rect 1848 1106 1849 1107
rect 1854 1107 1860 1108
rect 1854 1106 1855 1107
rect 1848 1104 1855 1106
rect 1848 1103 1849 1104
rect 1843 1102 1849 1103
rect 1854 1103 1855 1104
rect 1859 1103 1860 1107
rect 1854 1102 1860 1103
rect 1910 1107 1916 1108
rect 1910 1103 1911 1107
rect 1915 1103 1916 1107
rect 1910 1102 1916 1103
rect 1931 1107 1937 1108
rect 1931 1103 1932 1107
rect 1936 1106 1937 1107
rect 1998 1107 2004 1108
rect 1936 1104 1990 1106
rect 1936 1103 1937 1104
rect 1931 1102 1937 1103
rect 1757 1098 1759 1102
rect 1757 1096 1830 1098
rect 1828 1094 1830 1096
rect 1988 1094 1990 1104
rect 1998 1103 1999 1107
rect 2003 1103 2004 1107
rect 1998 1102 2004 1103
rect 2019 1107 2025 1108
rect 2019 1103 2020 1107
rect 2024 1106 2025 1107
rect 2086 1107 2092 1108
rect 2024 1104 2082 1106
rect 2024 1103 2025 1104
rect 2019 1102 2025 1103
rect 2080 1098 2082 1104
rect 2086 1103 2087 1107
rect 2091 1103 2092 1107
rect 2086 1102 2092 1103
rect 2107 1107 2113 1108
rect 2107 1103 2108 1107
rect 2112 1106 2113 1107
rect 2118 1107 2124 1108
rect 2118 1106 2119 1107
rect 2112 1104 2119 1106
rect 2112 1103 2113 1104
rect 2107 1102 2113 1103
rect 2118 1103 2119 1104
rect 2123 1103 2124 1107
rect 2118 1102 2124 1103
rect 2174 1107 2180 1108
rect 2174 1103 2175 1107
rect 2179 1103 2180 1107
rect 2174 1102 2180 1103
rect 2195 1107 2201 1108
rect 2195 1103 2196 1107
rect 2200 1106 2201 1107
rect 2270 1107 2276 1108
rect 2200 1104 2266 1106
rect 2200 1103 2201 1104
rect 2195 1102 2201 1103
rect 2264 1098 2266 1104
rect 2270 1103 2271 1107
rect 2275 1103 2276 1107
rect 2270 1102 2276 1103
rect 2291 1107 2297 1108
rect 2291 1103 2292 1107
rect 2296 1106 2297 1107
rect 2374 1107 2380 1108
rect 2296 1104 2370 1106
rect 2296 1103 2297 1104
rect 2291 1102 2297 1103
rect 2368 1098 2370 1104
rect 2374 1103 2375 1107
rect 2379 1103 2380 1107
rect 2374 1102 2380 1103
rect 2382 1107 2388 1108
rect 2382 1103 2383 1107
rect 2387 1106 2388 1107
rect 2395 1107 2401 1108
rect 2395 1106 2396 1107
rect 2387 1104 2396 1106
rect 2387 1103 2388 1104
rect 2382 1102 2388 1103
rect 2395 1103 2396 1104
rect 2400 1103 2401 1107
rect 2395 1102 2401 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2462 1107 2468 1108
rect 2462 1103 2463 1107
rect 2467 1106 2468 1107
rect 2475 1107 2481 1108
rect 2475 1106 2476 1107
rect 2467 1104 2476 1106
rect 2467 1103 2468 1104
rect 2462 1102 2468 1103
rect 2475 1103 2476 1104
rect 2480 1103 2481 1107
rect 2502 1104 2503 1108
rect 2507 1104 2508 1108
rect 2502 1103 2508 1104
rect 2475 1102 2481 1103
rect 2080 1096 2095 1098
rect 2264 1096 2278 1098
rect 2368 1096 2383 1098
rect 2093 1094 2095 1096
rect 2276 1094 2278 1096
rect 2381 1094 2383 1096
rect 1467 1093 1473 1094
rect 1387 1091 1393 1092
rect 110 1088 116 1089
rect 1286 1088 1292 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 238 1087 244 1088
rect 238 1083 239 1087
rect 243 1083 244 1087
rect 238 1082 244 1083
rect 259 1087 265 1088
rect 259 1083 260 1087
rect 264 1086 265 1087
rect 326 1087 332 1088
rect 264 1084 321 1086
rect 264 1083 265 1084
rect 259 1082 265 1083
rect 319 1074 321 1084
rect 326 1083 327 1087
rect 331 1083 332 1087
rect 326 1082 332 1083
rect 347 1087 353 1088
rect 347 1083 348 1087
rect 352 1083 353 1087
rect 347 1082 353 1083
rect 414 1087 420 1088
rect 414 1083 415 1087
rect 419 1083 420 1087
rect 414 1082 420 1083
rect 422 1087 428 1088
rect 422 1083 423 1087
rect 427 1086 428 1087
rect 435 1087 441 1088
rect 435 1086 436 1087
rect 427 1084 436 1086
rect 427 1083 428 1084
rect 422 1082 428 1083
rect 435 1083 436 1084
rect 440 1083 441 1087
rect 435 1082 441 1083
rect 510 1087 516 1088
rect 510 1083 511 1087
rect 515 1083 516 1087
rect 510 1082 516 1083
rect 526 1087 537 1088
rect 526 1083 527 1087
rect 531 1083 532 1087
rect 536 1083 537 1087
rect 526 1082 537 1083
rect 606 1087 612 1088
rect 606 1083 607 1087
rect 611 1083 612 1087
rect 627 1087 633 1088
rect 627 1086 628 1087
rect 606 1082 612 1083
rect 616 1084 628 1086
rect 349 1074 351 1082
rect 616 1078 618 1084
rect 627 1083 628 1084
rect 632 1083 633 1087
rect 627 1082 633 1083
rect 694 1087 700 1088
rect 694 1083 695 1087
rect 699 1083 700 1087
rect 694 1082 700 1083
rect 715 1087 721 1088
rect 715 1083 716 1087
rect 720 1086 721 1087
rect 782 1087 788 1088
rect 720 1084 774 1086
rect 720 1083 721 1084
rect 715 1082 721 1083
rect 516 1076 618 1078
rect 516 1074 518 1076
rect 772 1074 774 1084
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 803 1087 809 1088
rect 803 1083 804 1087
rect 808 1086 809 1087
rect 862 1087 868 1088
rect 808 1084 858 1086
rect 808 1083 809 1084
rect 803 1082 809 1083
rect 856 1074 858 1084
rect 862 1083 863 1087
rect 867 1083 868 1087
rect 862 1082 868 1083
rect 883 1087 892 1088
rect 883 1083 884 1087
rect 891 1083 892 1087
rect 883 1082 892 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 963 1087 969 1088
rect 963 1086 964 1087
rect 942 1082 948 1083
rect 952 1084 964 1086
rect 952 1078 954 1084
rect 963 1083 964 1084
rect 968 1083 969 1087
rect 963 1082 969 1083
rect 1030 1087 1036 1088
rect 1030 1083 1031 1087
rect 1035 1083 1036 1087
rect 1030 1082 1036 1083
rect 1051 1087 1057 1088
rect 1051 1083 1052 1087
rect 1056 1086 1057 1087
rect 1118 1087 1124 1088
rect 1056 1084 1110 1086
rect 1056 1083 1057 1084
rect 1051 1082 1057 1083
rect 876 1076 954 1078
rect 319 1073 337 1074
rect 319 1072 332 1073
rect 243 1071 249 1072
rect 243 1067 244 1071
rect 248 1070 249 1071
rect 248 1068 321 1070
rect 331 1069 332 1072
rect 336 1069 337 1073
rect 349 1073 425 1074
rect 349 1072 420 1073
rect 331 1068 337 1069
rect 419 1069 420 1072
rect 424 1069 425 1073
rect 419 1068 425 1069
rect 515 1073 521 1074
rect 515 1069 516 1073
rect 520 1069 521 1073
rect 772 1073 793 1074
rect 772 1072 788 1073
rect 515 1068 521 1069
rect 582 1071 588 1072
rect 248 1067 249 1068
rect 243 1066 249 1067
rect 319 1066 321 1068
rect 526 1067 532 1068
rect 526 1066 527 1067
rect 319 1064 527 1066
rect 526 1063 527 1064
rect 531 1063 532 1067
rect 582 1067 583 1071
rect 587 1070 588 1071
rect 611 1071 617 1072
rect 611 1070 612 1071
rect 587 1068 612 1070
rect 587 1067 588 1068
rect 582 1066 588 1067
rect 611 1067 612 1068
rect 616 1067 617 1071
rect 611 1066 617 1067
rect 699 1071 705 1072
rect 699 1067 700 1071
rect 704 1070 705 1071
rect 704 1068 782 1070
rect 787 1069 788 1072
rect 792 1069 793 1073
rect 856 1073 873 1074
rect 856 1072 868 1073
rect 787 1068 793 1069
rect 867 1069 868 1072
rect 872 1069 873 1073
rect 867 1068 873 1069
rect 704 1067 705 1068
rect 699 1066 705 1067
rect 780 1066 782 1068
rect 876 1066 878 1076
rect 1108 1074 1110 1084
rect 1118 1083 1119 1087
rect 1123 1083 1124 1087
rect 1118 1082 1124 1083
rect 1126 1087 1132 1088
rect 1126 1083 1127 1087
rect 1131 1086 1132 1087
rect 1139 1087 1145 1088
rect 1139 1086 1140 1087
rect 1131 1084 1140 1086
rect 1131 1083 1132 1084
rect 1126 1082 1132 1083
rect 1139 1083 1140 1084
rect 1144 1083 1145 1087
rect 1286 1084 1287 1088
rect 1291 1084 1292 1088
rect 1387 1087 1388 1091
rect 1392 1087 1393 1091
rect 1467 1089 1468 1093
rect 1472 1089 1473 1093
rect 1728 1093 1745 1094
rect 1728 1092 1740 1093
rect 1467 1088 1473 1089
rect 1555 1091 1561 1092
rect 1387 1086 1393 1087
rect 1478 1087 1484 1088
rect 1478 1086 1479 1087
rect 1389 1084 1479 1086
rect 1286 1083 1292 1084
rect 1478 1083 1479 1084
rect 1483 1083 1484 1087
rect 1555 1087 1556 1091
rect 1560 1090 1561 1091
rect 1606 1091 1612 1092
rect 1606 1090 1607 1091
rect 1560 1088 1607 1090
rect 1560 1087 1561 1088
rect 1555 1086 1561 1087
rect 1606 1087 1607 1088
rect 1611 1087 1612 1091
rect 1606 1086 1612 1087
rect 1651 1091 1657 1092
rect 1651 1087 1652 1091
rect 1656 1087 1657 1091
rect 1739 1089 1740 1092
rect 1744 1089 1745 1093
rect 1739 1088 1745 1089
rect 1827 1093 1833 1094
rect 1827 1089 1828 1093
rect 1832 1089 1833 1093
rect 1988 1093 2009 1094
rect 1988 1092 2004 1093
rect 1827 1088 1833 1089
rect 1915 1091 1921 1092
rect 1651 1086 1657 1087
rect 1786 1087 1792 1088
rect 1786 1086 1787 1087
rect 1653 1084 1787 1086
rect 1139 1082 1145 1083
rect 1478 1082 1484 1083
rect 1786 1083 1787 1084
rect 1791 1083 1792 1087
rect 1915 1087 1916 1091
rect 1920 1090 1921 1091
rect 1958 1091 1964 1092
rect 1958 1090 1959 1091
rect 1920 1088 1959 1090
rect 1920 1087 1921 1088
rect 1915 1086 1921 1087
rect 1958 1087 1959 1088
rect 1963 1087 1964 1091
rect 2003 1089 2004 1092
rect 2008 1089 2009 1093
rect 2003 1088 2009 1089
rect 2091 1093 2097 1094
rect 2091 1089 2092 1093
rect 2096 1089 2097 1093
rect 2275 1093 2281 1094
rect 2091 1088 2097 1089
rect 2166 1091 2172 1092
rect 1958 1086 1964 1087
rect 2166 1087 2167 1091
rect 2171 1090 2172 1091
rect 2179 1091 2185 1092
rect 2179 1090 2180 1091
rect 2171 1088 2180 1090
rect 2171 1087 2172 1088
rect 2166 1086 2172 1087
rect 2179 1087 2180 1088
rect 2184 1087 2185 1091
rect 2275 1089 2276 1093
rect 2280 1089 2281 1093
rect 2275 1088 2281 1089
rect 2379 1093 2385 1094
rect 2379 1089 2380 1093
rect 2384 1089 2385 1093
rect 2379 1088 2385 1089
rect 2459 1091 2465 1092
rect 2179 1086 2185 1087
rect 2459 1087 2460 1091
rect 2464 1090 2465 1091
rect 2470 1091 2476 1092
rect 2470 1090 2471 1091
rect 2464 1088 2471 1090
rect 2464 1087 2465 1088
rect 2459 1086 2465 1087
rect 2470 1087 2471 1088
rect 2475 1087 2476 1091
rect 2470 1086 2476 1087
rect 1786 1082 1792 1083
rect 1108 1073 1129 1074
rect 1108 1072 1124 1073
rect 947 1071 953 1072
rect 947 1067 948 1071
rect 952 1070 953 1071
rect 1006 1071 1012 1072
rect 952 1068 1002 1070
rect 952 1067 953 1068
rect 947 1066 953 1067
rect 780 1064 878 1066
rect 526 1062 532 1063
rect 1000 1062 1002 1068
rect 1006 1067 1007 1071
rect 1011 1070 1012 1071
rect 1035 1071 1041 1072
rect 1035 1070 1036 1071
rect 1011 1068 1036 1070
rect 1011 1067 1012 1068
rect 1006 1066 1012 1067
rect 1035 1067 1036 1068
rect 1040 1067 1041 1071
rect 1123 1069 1124 1072
rect 1128 1069 1129 1073
rect 2366 1071 2372 1072
rect 2366 1070 2367 1071
rect 1123 1068 1129 1069
rect 1845 1068 2367 1070
rect 1035 1066 1041 1067
rect 1845 1066 1847 1068
rect 2366 1067 2367 1068
rect 2371 1067 2372 1071
rect 2366 1066 2372 1067
rect 1843 1065 1849 1066
rect 1126 1063 1132 1064
rect 1126 1062 1127 1063
rect 1000 1060 1127 1062
rect 1126 1059 1127 1060
rect 1131 1059 1132 1063
rect 1126 1058 1132 1059
rect 1422 1063 1428 1064
rect 1422 1059 1423 1063
rect 1427 1062 1428 1063
rect 1435 1063 1441 1064
rect 1435 1062 1436 1063
rect 1427 1060 1436 1062
rect 1427 1059 1428 1060
rect 1422 1058 1428 1059
rect 1435 1059 1436 1060
rect 1440 1059 1441 1063
rect 1499 1063 1505 1064
rect 1499 1062 1500 1063
rect 1435 1058 1441 1059
rect 1452 1060 1500 1062
rect 674 1055 680 1056
rect 674 1054 675 1055
rect 156 1052 675 1054
rect 156 1050 158 1052
rect 674 1051 675 1052
rect 679 1051 680 1055
rect 674 1050 680 1051
rect 798 1055 804 1056
rect 798 1051 799 1055
rect 803 1054 804 1055
rect 803 1052 1102 1054
rect 803 1051 804 1052
rect 798 1050 804 1051
rect 1100 1050 1102 1052
rect 1452 1050 1454 1060
rect 1499 1059 1500 1060
rect 1504 1059 1505 1063
rect 1499 1058 1505 1059
rect 1571 1063 1577 1064
rect 1571 1059 1572 1063
rect 1576 1059 1577 1063
rect 1643 1063 1649 1064
rect 1643 1062 1644 1063
rect 1571 1058 1577 1059
rect 1588 1060 1644 1062
rect 1516 1056 1575 1058
rect 1516 1050 1518 1056
rect 1588 1050 1590 1060
rect 1643 1059 1644 1060
rect 1648 1059 1649 1063
rect 1643 1058 1649 1059
rect 1707 1063 1716 1064
rect 1707 1059 1708 1063
rect 1715 1059 1716 1063
rect 1771 1063 1777 1064
rect 1771 1062 1772 1063
rect 1707 1058 1716 1059
rect 1724 1060 1772 1062
rect 1724 1050 1726 1060
rect 1771 1059 1772 1060
rect 1776 1059 1777 1063
rect 1843 1061 1844 1065
rect 1848 1061 1849 1065
rect 1843 1060 1849 1061
rect 1923 1063 1929 1064
rect 1771 1058 1777 1059
rect 1923 1059 1924 1063
rect 1928 1059 1929 1063
rect 2011 1063 2017 1064
rect 2011 1062 2012 1063
rect 1923 1058 1929 1059
rect 1999 1060 2012 1062
rect 1860 1056 1927 1058
rect 1860 1050 1862 1056
rect 1999 1054 2001 1060
rect 2011 1059 2012 1060
rect 2016 1059 2017 1063
rect 2011 1058 2017 1059
rect 2115 1063 2124 1064
rect 2115 1059 2116 1063
rect 2123 1059 2124 1063
rect 2115 1058 2124 1059
rect 2235 1063 2241 1064
rect 2235 1059 2236 1063
rect 2240 1059 2241 1063
rect 2235 1058 2241 1059
rect 2355 1063 2361 1064
rect 2355 1059 2356 1063
rect 2360 1059 2361 1063
rect 2355 1058 2361 1059
rect 2459 1063 2468 1064
rect 2459 1059 2460 1063
rect 2467 1059 2468 1063
rect 2459 1058 2468 1059
rect 1940 1052 2001 1054
rect 2132 1056 2239 1058
rect 2252 1056 2359 1058
rect 1940 1050 1942 1052
rect 2132 1050 2134 1056
rect 2252 1050 2254 1056
rect 155 1049 161 1050
rect 155 1045 156 1049
rect 160 1045 161 1049
rect 1099 1049 1105 1050
rect 1430 1049 1436 1050
rect 211 1047 217 1048
rect 211 1046 212 1047
rect 155 1044 161 1045
rect 173 1044 212 1046
rect 173 1034 175 1044
rect 211 1043 212 1044
rect 216 1043 217 1047
rect 307 1047 313 1048
rect 307 1046 308 1047
rect 211 1042 217 1043
rect 228 1044 308 1046
rect 228 1034 230 1044
rect 307 1043 308 1044
rect 312 1043 313 1047
rect 307 1042 313 1043
rect 419 1047 428 1048
rect 419 1043 420 1047
rect 427 1043 428 1047
rect 419 1042 428 1043
rect 539 1047 545 1048
rect 539 1043 540 1047
rect 544 1043 545 1047
rect 659 1047 665 1048
rect 659 1046 660 1047
rect 539 1042 545 1043
rect 556 1044 660 1046
rect 541 1038 543 1042
rect 436 1036 543 1038
rect 436 1034 438 1036
rect 556 1034 558 1044
rect 659 1043 660 1044
rect 664 1043 665 1047
rect 659 1042 665 1043
rect 771 1047 780 1048
rect 771 1043 772 1047
rect 779 1043 780 1047
rect 883 1047 889 1048
rect 883 1046 884 1047
rect 771 1042 780 1043
rect 788 1044 884 1046
rect 788 1034 790 1044
rect 883 1043 884 1044
rect 888 1043 889 1047
rect 987 1047 993 1048
rect 987 1046 988 1047
rect 883 1042 889 1043
rect 900 1044 988 1046
rect 900 1034 902 1044
rect 987 1043 988 1044
rect 992 1043 993 1047
rect 1099 1045 1100 1049
rect 1104 1045 1105 1049
rect 1326 1048 1332 1049
rect 1211 1047 1217 1048
rect 1211 1046 1212 1047
rect 1099 1044 1105 1045
rect 1159 1044 1212 1046
rect 987 1042 993 1043
rect 1159 1038 1161 1044
rect 1211 1043 1212 1044
rect 1216 1043 1217 1047
rect 1326 1044 1327 1048
rect 1331 1044 1332 1048
rect 1430 1045 1431 1049
rect 1435 1045 1436 1049
rect 1430 1044 1436 1045
rect 1451 1049 1457 1050
rect 1451 1045 1452 1049
rect 1456 1045 1457 1049
rect 1451 1044 1457 1045
rect 1494 1049 1500 1050
rect 1494 1045 1495 1049
rect 1499 1045 1500 1049
rect 1494 1044 1500 1045
rect 1515 1049 1521 1050
rect 1515 1045 1516 1049
rect 1520 1045 1521 1049
rect 1515 1044 1521 1045
rect 1566 1049 1572 1050
rect 1566 1045 1567 1049
rect 1571 1045 1572 1049
rect 1566 1044 1572 1045
rect 1587 1049 1593 1050
rect 1587 1045 1588 1049
rect 1592 1045 1593 1049
rect 1587 1044 1593 1045
rect 1638 1049 1644 1050
rect 1638 1045 1639 1049
rect 1643 1045 1644 1049
rect 1702 1049 1708 1050
rect 1638 1044 1644 1045
rect 1646 1047 1652 1048
rect 1326 1043 1332 1044
rect 1646 1043 1647 1047
rect 1651 1046 1652 1047
rect 1659 1047 1665 1048
rect 1659 1046 1660 1047
rect 1651 1044 1660 1046
rect 1651 1043 1652 1044
rect 1211 1042 1217 1043
rect 1646 1042 1652 1043
rect 1659 1043 1660 1044
rect 1664 1043 1665 1047
rect 1702 1045 1703 1049
rect 1707 1045 1708 1049
rect 1702 1044 1708 1045
rect 1723 1049 1729 1050
rect 1723 1045 1724 1049
rect 1728 1045 1729 1049
rect 1723 1044 1729 1045
rect 1766 1049 1772 1050
rect 1766 1045 1767 1049
rect 1771 1045 1772 1049
rect 1838 1049 1844 1050
rect 1766 1044 1772 1045
rect 1786 1047 1793 1048
rect 1659 1042 1665 1043
rect 1786 1043 1787 1047
rect 1792 1043 1793 1047
rect 1838 1045 1839 1049
rect 1843 1045 1844 1049
rect 1838 1044 1844 1045
rect 1859 1049 1865 1050
rect 1859 1045 1860 1049
rect 1864 1045 1865 1049
rect 1859 1044 1865 1045
rect 1918 1049 1924 1050
rect 1918 1045 1919 1049
rect 1923 1045 1924 1049
rect 1918 1044 1924 1045
rect 1939 1049 1945 1050
rect 1939 1045 1940 1049
rect 1944 1045 1945 1049
rect 1939 1044 1945 1045
rect 2006 1049 2012 1050
rect 2006 1045 2007 1049
rect 2011 1045 2012 1049
rect 2110 1049 2116 1050
rect 2006 1044 2012 1045
rect 2014 1047 2020 1048
rect 1786 1042 1793 1043
rect 2014 1043 2015 1047
rect 2019 1046 2020 1047
rect 2027 1047 2033 1048
rect 2027 1046 2028 1047
rect 2019 1044 2028 1046
rect 2019 1043 2020 1044
rect 2014 1042 2020 1043
rect 2027 1043 2028 1044
rect 2032 1043 2033 1047
rect 2110 1045 2111 1049
rect 2115 1045 2116 1049
rect 2110 1044 2116 1045
rect 2131 1049 2137 1050
rect 2131 1045 2132 1049
rect 2136 1045 2137 1049
rect 2131 1044 2137 1045
rect 2230 1049 2236 1050
rect 2230 1045 2231 1049
rect 2235 1045 2236 1049
rect 2230 1044 2236 1045
rect 2251 1049 2257 1050
rect 2251 1045 2252 1049
rect 2256 1045 2257 1049
rect 2251 1044 2257 1045
rect 2350 1049 2356 1050
rect 2350 1045 2351 1049
rect 2355 1045 2356 1049
rect 2454 1049 2460 1050
rect 2350 1044 2356 1045
rect 2366 1047 2377 1048
rect 2027 1042 2033 1043
rect 2366 1043 2367 1047
rect 2371 1043 2372 1047
rect 2376 1043 2377 1047
rect 2454 1045 2455 1049
rect 2459 1045 2460 1049
rect 2502 1048 2508 1049
rect 2454 1044 2460 1045
rect 2462 1047 2468 1048
rect 2366 1042 2377 1043
rect 2462 1043 2463 1047
rect 2467 1046 2468 1047
rect 2475 1047 2481 1048
rect 2475 1046 2476 1047
rect 2467 1044 2476 1046
rect 2467 1043 2468 1044
rect 2462 1042 2468 1043
rect 2475 1043 2476 1044
rect 2480 1043 2481 1047
rect 2502 1044 2503 1048
rect 2507 1044 2508 1048
rect 2502 1043 2508 1044
rect 2475 1042 2481 1043
rect 1116 1036 1161 1038
rect 1116 1034 1118 1036
rect 150 1033 156 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 150 1029 151 1033
rect 155 1029 156 1033
rect 150 1028 156 1029
rect 171 1033 177 1034
rect 171 1029 172 1033
rect 176 1029 177 1033
rect 171 1028 177 1029
rect 206 1033 212 1034
rect 206 1029 207 1033
rect 211 1029 212 1033
rect 206 1028 212 1029
rect 227 1033 233 1034
rect 227 1029 228 1033
rect 232 1029 233 1033
rect 227 1028 233 1029
rect 302 1033 308 1034
rect 302 1029 303 1033
rect 307 1029 308 1033
rect 414 1033 420 1034
rect 302 1028 308 1029
rect 323 1031 329 1032
rect 110 1027 116 1028
rect 323 1027 324 1031
rect 328 1030 329 1031
rect 334 1031 340 1032
rect 334 1030 335 1031
rect 328 1028 335 1030
rect 328 1027 329 1028
rect 323 1026 329 1027
rect 334 1027 335 1028
rect 339 1027 340 1031
rect 414 1029 415 1033
rect 419 1029 420 1033
rect 414 1028 420 1029
rect 435 1033 441 1034
rect 435 1029 436 1033
rect 440 1029 441 1033
rect 435 1028 441 1029
rect 534 1033 540 1034
rect 534 1029 535 1033
rect 539 1029 540 1033
rect 534 1028 540 1029
rect 555 1033 561 1034
rect 555 1029 556 1033
rect 560 1029 561 1033
rect 555 1028 561 1029
rect 654 1033 660 1034
rect 654 1029 655 1033
rect 659 1029 660 1033
rect 766 1033 772 1034
rect 654 1028 660 1029
rect 674 1031 681 1032
rect 334 1026 340 1027
rect 674 1027 675 1031
rect 680 1027 681 1031
rect 766 1029 767 1033
rect 771 1029 772 1033
rect 766 1028 772 1029
rect 787 1033 793 1034
rect 787 1029 788 1033
rect 792 1029 793 1033
rect 787 1028 793 1029
rect 878 1033 884 1034
rect 878 1029 879 1033
rect 883 1029 884 1033
rect 878 1028 884 1029
rect 899 1033 905 1034
rect 899 1029 900 1033
rect 904 1029 905 1033
rect 899 1028 905 1029
rect 982 1033 988 1034
rect 982 1029 983 1033
rect 987 1029 988 1033
rect 1094 1033 1100 1034
rect 982 1028 988 1029
rect 1003 1031 1012 1032
rect 674 1026 681 1027
rect 1003 1027 1004 1031
rect 1011 1027 1012 1031
rect 1094 1029 1095 1033
rect 1099 1029 1100 1033
rect 1094 1028 1100 1029
rect 1115 1033 1121 1034
rect 1115 1029 1116 1033
rect 1120 1029 1121 1033
rect 1115 1028 1121 1029
rect 1206 1033 1212 1034
rect 1206 1029 1207 1033
rect 1211 1029 1212 1033
rect 1286 1032 1292 1033
rect 1206 1028 1212 1029
rect 1226 1031 1233 1032
rect 1003 1026 1012 1027
rect 1226 1027 1227 1031
rect 1232 1027 1233 1031
rect 1286 1028 1287 1032
rect 1291 1028 1292 1032
rect 1286 1027 1292 1028
rect 1326 1031 1332 1032
rect 1326 1027 1327 1031
rect 1331 1027 1332 1031
rect 2502 1031 2508 1032
rect 1226 1026 1233 1027
rect 1326 1026 1332 1027
rect 1414 1028 1420 1029
rect 1414 1024 1415 1028
rect 1419 1024 1420 1028
rect 1414 1023 1420 1024
rect 1478 1028 1484 1029
rect 1478 1024 1479 1028
rect 1483 1024 1484 1028
rect 1478 1023 1484 1024
rect 1550 1028 1556 1029
rect 1550 1024 1551 1028
rect 1555 1024 1556 1028
rect 1550 1023 1556 1024
rect 1622 1028 1628 1029
rect 1622 1024 1623 1028
rect 1627 1024 1628 1028
rect 1622 1023 1628 1024
rect 1686 1028 1692 1029
rect 1686 1024 1687 1028
rect 1691 1024 1692 1028
rect 1686 1023 1692 1024
rect 1750 1028 1756 1029
rect 1750 1024 1751 1028
rect 1755 1024 1756 1028
rect 1750 1023 1756 1024
rect 1822 1028 1828 1029
rect 1822 1024 1823 1028
rect 1827 1024 1828 1028
rect 1822 1023 1828 1024
rect 1902 1028 1908 1029
rect 1902 1024 1903 1028
rect 1907 1024 1908 1028
rect 1902 1023 1908 1024
rect 1990 1028 1996 1029
rect 1990 1024 1991 1028
rect 1995 1024 1996 1028
rect 1990 1023 1996 1024
rect 2094 1028 2100 1029
rect 2094 1024 2095 1028
rect 2099 1024 2100 1028
rect 2094 1023 2100 1024
rect 2214 1028 2220 1029
rect 2214 1024 2215 1028
rect 2219 1024 2220 1028
rect 2214 1023 2220 1024
rect 2334 1028 2340 1029
rect 2334 1024 2335 1028
rect 2339 1024 2340 1028
rect 2334 1023 2340 1024
rect 2438 1028 2444 1029
rect 2438 1024 2439 1028
rect 2443 1024 2444 1028
rect 2502 1027 2503 1031
rect 2507 1027 2508 1031
rect 2502 1026 2508 1027
rect 2438 1023 2444 1024
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 1286 1015 1292 1016
rect 110 1010 116 1011
rect 134 1012 140 1013
rect 134 1008 135 1012
rect 139 1008 140 1012
rect 134 1007 140 1008
rect 190 1012 196 1013
rect 190 1008 191 1012
rect 195 1008 196 1012
rect 190 1007 196 1008
rect 286 1012 292 1013
rect 286 1008 287 1012
rect 291 1008 292 1012
rect 286 1007 292 1008
rect 398 1012 404 1013
rect 398 1008 399 1012
rect 403 1008 404 1012
rect 398 1007 404 1008
rect 518 1012 524 1013
rect 518 1008 519 1012
rect 523 1008 524 1012
rect 518 1007 524 1008
rect 638 1012 644 1013
rect 638 1008 639 1012
rect 643 1008 644 1012
rect 638 1007 644 1008
rect 750 1012 756 1013
rect 750 1008 751 1012
rect 755 1008 756 1012
rect 750 1007 756 1008
rect 862 1012 868 1013
rect 862 1008 863 1012
rect 867 1008 868 1012
rect 862 1007 868 1008
rect 966 1012 972 1013
rect 966 1008 967 1012
rect 971 1008 972 1012
rect 966 1007 972 1008
rect 1078 1012 1084 1013
rect 1078 1008 1079 1012
rect 1083 1008 1084 1012
rect 1078 1007 1084 1008
rect 1190 1012 1196 1013
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1286 1011 1287 1015
rect 1291 1011 1292 1015
rect 1286 1010 1292 1011
rect 1190 1007 1196 1008
rect 1510 1008 1516 1009
rect 1326 1005 1332 1006
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1566 1008 1572 1009
rect 1566 1004 1567 1008
rect 1571 1004 1572 1008
rect 1566 1003 1572 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1734 1008 1740 1009
rect 1734 1004 1735 1008
rect 1739 1004 1740 1008
rect 1734 1003 1740 1004
rect 1806 1008 1812 1009
rect 1806 1004 1807 1008
rect 1811 1004 1812 1008
rect 1806 1003 1812 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1982 1008 1988 1009
rect 1982 1004 1983 1008
rect 1987 1004 1988 1008
rect 1982 1003 1988 1004
rect 2094 1008 2100 1009
rect 2094 1004 2095 1008
rect 2099 1004 2100 1008
rect 2094 1003 2100 1004
rect 2214 1008 2220 1009
rect 2214 1004 2215 1008
rect 2219 1004 2220 1008
rect 2214 1003 2220 1004
rect 2334 1008 2340 1009
rect 2334 1004 2335 1008
rect 2339 1004 2340 1008
rect 2334 1003 2340 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 2502 1005 2508 1006
rect 1326 1000 1332 1001
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 134 996 140 997
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 134 992 135 996
rect 139 992 140 996
rect 134 991 140 992
rect 214 996 220 997
rect 214 992 215 996
rect 219 992 220 996
rect 214 991 220 992
rect 326 996 332 997
rect 326 992 327 996
rect 331 992 332 996
rect 326 991 332 992
rect 438 996 444 997
rect 438 992 439 996
rect 443 992 444 996
rect 438 991 444 992
rect 550 996 556 997
rect 550 992 551 996
rect 555 992 556 996
rect 550 991 556 992
rect 662 996 668 997
rect 662 992 663 996
rect 667 992 668 996
rect 662 991 668 992
rect 758 996 764 997
rect 758 992 759 996
rect 763 992 764 996
rect 758 991 764 992
rect 846 996 852 997
rect 846 992 847 996
rect 851 992 852 996
rect 846 991 852 992
rect 934 996 940 997
rect 934 992 935 996
rect 939 992 940 996
rect 934 991 940 992
rect 1014 996 1020 997
rect 1014 992 1015 996
rect 1019 992 1020 996
rect 1014 991 1020 992
rect 1086 996 1092 997
rect 1086 992 1087 996
rect 1091 992 1092 996
rect 1086 991 1092 992
rect 1166 996 1172 997
rect 1166 992 1167 996
rect 1171 992 1172 996
rect 1166 991 1172 992
rect 1222 996 1228 997
rect 1222 992 1223 996
rect 1227 992 1228 996
rect 1222 991 1228 992
rect 1286 993 1292 994
rect 110 988 116 989
rect 1286 989 1287 993
rect 1291 989 1292 993
rect 1286 988 1292 989
rect 1326 988 1332 989
rect 2502 988 2508 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1526 982 1532 983
rect 1534 987 1540 988
rect 1534 983 1535 987
rect 1539 986 1540 987
rect 1547 987 1553 988
rect 1547 986 1548 987
rect 1539 984 1548 986
rect 1539 983 1540 984
rect 1534 982 1540 983
rect 1547 983 1548 984
rect 1552 983 1553 987
rect 1547 982 1553 983
rect 1582 987 1588 988
rect 1582 983 1583 987
rect 1587 983 1588 987
rect 1582 982 1588 983
rect 1598 987 1609 988
rect 1598 983 1599 987
rect 1603 983 1604 987
rect 1608 983 1609 987
rect 1598 982 1609 983
rect 1638 987 1644 988
rect 1638 983 1639 987
rect 1643 983 1644 987
rect 1659 987 1665 988
rect 1659 986 1660 987
rect 1638 982 1644 983
rect 1648 984 1660 986
rect 1648 978 1650 984
rect 1659 983 1660 984
rect 1664 983 1665 987
rect 1659 982 1665 983
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1710 987 1721 988
rect 1710 983 1711 987
rect 1715 983 1716 987
rect 1720 983 1721 987
rect 1710 982 1721 983
rect 1750 987 1756 988
rect 1750 983 1751 987
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1771 987 1777 988
rect 1771 983 1772 987
rect 1776 986 1777 987
rect 1782 987 1788 988
rect 1782 986 1783 987
rect 1776 984 1783 986
rect 1776 983 1777 984
rect 1771 982 1777 983
rect 1782 983 1783 984
rect 1787 983 1788 987
rect 1782 982 1788 983
rect 1822 987 1828 988
rect 1822 983 1823 987
rect 1827 983 1828 987
rect 1822 982 1828 983
rect 1843 987 1849 988
rect 1843 983 1844 987
rect 1848 983 1849 987
rect 1843 982 1849 983
rect 1902 987 1908 988
rect 1902 983 1903 987
rect 1907 983 1908 987
rect 1902 982 1908 983
rect 1923 987 1929 988
rect 1923 983 1924 987
rect 1928 983 1929 987
rect 1923 982 1929 983
rect 1998 987 2004 988
rect 1998 983 1999 987
rect 2003 983 2004 987
rect 1998 982 2004 983
rect 2019 987 2025 988
rect 2019 983 2020 987
rect 2024 983 2025 987
rect 2019 982 2025 983
rect 2110 987 2116 988
rect 2110 983 2111 987
rect 2115 983 2116 987
rect 2110 982 2116 983
rect 2131 987 2137 988
rect 2131 983 2132 987
rect 2136 986 2137 987
rect 2230 987 2236 988
rect 2136 984 2226 986
rect 2136 983 2137 984
rect 2131 982 2137 983
rect 1845 978 1847 982
rect 1925 978 1927 982
rect 110 976 116 977
rect 1286 976 1292 977
rect 110 972 111 976
rect 115 972 116 976
rect 110 971 116 972
rect 150 975 156 976
rect 150 971 151 975
rect 155 971 156 975
rect 150 970 156 971
rect 158 975 164 976
rect 158 971 159 975
rect 163 974 164 975
rect 171 975 177 976
rect 171 974 172 975
rect 163 972 172 974
rect 163 971 164 972
rect 158 970 164 971
rect 171 971 172 972
rect 176 971 177 975
rect 171 970 177 971
rect 230 975 236 976
rect 230 971 231 975
rect 235 971 236 975
rect 230 970 236 971
rect 251 975 257 976
rect 251 971 252 975
rect 256 971 257 975
rect 251 970 257 971
rect 342 975 348 976
rect 342 971 343 975
rect 347 971 348 975
rect 342 970 348 971
rect 363 975 369 976
rect 363 971 364 975
rect 368 974 369 975
rect 454 975 460 976
rect 368 972 446 974
rect 368 971 369 972
rect 363 970 369 971
rect 253 966 255 970
rect 156 964 255 966
rect 156 962 158 964
rect 444 962 446 972
rect 454 971 455 975
rect 459 971 460 975
rect 454 970 460 971
rect 475 975 481 976
rect 475 971 476 975
rect 480 974 481 975
rect 566 975 572 976
rect 480 972 562 974
rect 480 971 481 972
rect 475 970 481 971
rect 560 962 562 972
rect 566 971 567 975
rect 571 971 572 975
rect 566 970 572 971
rect 574 975 580 976
rect 574 971 575 975
rect 579 974 580 975
rect 587 975 593 976
rect 587 974 588 975
rect 579 972 588 974
rect 579 971 580 972
rect 574 970 580 971
rect 587 971 588 972
rect 592 971 593 975
rect 587 970 593 971
rect 678 975 684 976
rect 678 971 679 975
rect 683 971 684 975
rect 678 970 684 971
rect 699 975 705 976
rect 699 971 700 975
rect 704 974 705 975
rect 774 975 780 976
rect 704 972 770 974
rect 704 971 705 972
rect 699 970 705 971
rect 768 962 770 972
rect 774 971 775 975
rect 779 971 780 975
rect 774 970 780 971
rect 795 975 804 976
rect 795 971 796 975
rect 803 971 804 975
rect 795 970 804 971
rect 862 975 868 976
rect 862 971 863 975
rect 867 971 868 975
rect 862 970 868 971
rect 883 975 889 976
rect 883 971 884 975
rect 888 974 889 975
rect 918 975 924 976
rect 918 974 919 975
rect 888 972 919 974
rect 888 971 889 972
rect 883 970 889 971
rect 918 971 919 972
rect 923 971 924 975
rect 918 970 924 971
rect 950 975 956 976
rect 950 971 951 975
rect 955 971 956 975
rect 971 975 977 976
rect 971 974 972 975
rect 950 970 956 971
rect 960 972 972 974
rect 960 966 962 972
rect 971 971 972 972
rect 976 971 977 975
rect 971 970 977 971
rect 1030 975 1036 976
rect 1030 971 1031 975
rect 1035 971 1036 975
rect 1030 970 1036 971
rect 1046 975 1057 976
rect 1046 971 1047 975
rect 1051 971 1052 975
rect 1056 971 1057 975
rect 1046 970 1057 971
rect 1102 975 1108 976
rect 1102 971 1103 975
rect 1107 971 1108 975
rect 1123 975 1129 976
rect 1123 974 1124 975
rect 1102 970 1108 971
rect 1112 972 1124 974
rect 1112 966 1114 972
rect 1123 971 1124 972
rect 1128 971 1129 975
rect 1123 970 1129 971
rect 1182 975 1188 976
rect 1182 971 1183 975
rect 1187 971 1188 975
rect 1182 970 1188 971
rect 1203 975 1209 976
rect 1203 971 1204 975
rect 1208 974 1209 975
rect 1238 975 1244 976
rect 1208 972 1234 974
rect 1208 971 1209 972
rect 1203 970 1209 971
rect 788 964 962 966
rect 1036 964 1114 966
rect 155 961 161 962
rect 155 957 156 961
rect 160 957 161 961
rect 444 961 465 962
rect 444 960 460 961
rect 155 956 161 957
rect 235 959 241 960
rect 235 955 236 959
rect 240 958 241 959
rect 334 959 340 960
rect 240 956 321 958
rect 240 955 241 956
rect 235 954 241 955
rect 319 950 321 956
rect 334 955 335 959
rect 339 958 340 959
rect 347 959 353 960
rect 347 958 348 959
rect 339 956 348 958
rect 339 955 340 956
rect 334 954 340 955
rect 347 955 348 956
rect 352 955 353 959
rect 459 957 460 960
rect 464 957 465 961
rect 560 961 577 962
rect 560 960 572 961
rect 459 956 465 957
rect 571 957 572 960
rect 576 957 577 961
rect 768 961 785 962
rect 768 960 780 961
rect 571 956 577 957
rect 683 959 689 960
rect 347 954 353 955
rect 683 955 684 959
rect 688 958 689 959
rect 688 956 774 958
rect 779 957 780 960
rect 784 957 785 961
rect 779 956 785 957
rect 688 955 689 956
rect 683 954 689 955
rect 772 954 774 956
rect 788 954 790 964
rect 1036 962 1038 964
rect 1232 962 1234 972
rect 1238 971 1239 975
rect 1243 971 1244 975
rect 1238 970 1244 971
rect 1246 975 1252 976
rect 1246 971 1247 975
rect 1251 974 1252 975
rect 1259 975 1265 976
rect 1259 974 1260 975
rect 1251 972 1260 974
rect 1251 971 1252 972
rect 1246 970 1252 971
rect 1259 971 1260 972
rect 1264 971 1265 975
rect 1286 972 1287 976
rect 1291 972 1292 976
rect 1588 976 1650 978
rect 1757 976 1847 978
rect 1852 976 1927 978
rect 1588 974 1590 976
rect 1757 974 1759 976
rect 1852 974 1854 976
rect 2006 975 2012 976
rect 2006 974 2007 975
rect 1587 973 1593 974
rect 1286 971 1292 972
rect 1531 971 1537 972
rect 1259 970 1265 971
rect 1531 967 1532 971
rect 1536 970 1537 971
rect 1536 968 1570 970
rect 1587 969 1588 973
rect 1592 969 1593 973
rect 1755 973 1761 974
rect 1587 968 1593 969
rect 1643 971 1652 972
rect 1536 967 1537 968
rect 1531 966 1537 967
rect 1568 966 1570 968
rect 1598 967 1604 968
rect 1598 966 1599 967
rect 1568 964 1599 966
rect 1598 963 1599 964
rect 1603 963 1604 967
rect 1643 967 1644 971
rect 1651 967 1652 971
rect 1643 966 1652 967
rect 1654 971 1660 972
rect 1654 967 1655 971
rect 1659 970 1660 971
rect 1699 971 1705 972
rect 1699 970 1700 971
rect 1659 968 1700 970
rect 1659 967 1660 968
rect 1654 966 1660 967
rect 1699 967 1700 968
rect 1704 967 1705 971
rect 1755 969 1756 973
rect 1760 969 1761 973
rect 1755 968 1761 969
rect 1827 973 1854 974
rect 1827 969 1828 973
rect 1832 972 1854 973
rect 2003 973 2007 974
rect 1832 969 1833 972
rect 1827 968 1833 969
rect 1907 971 1913 972
rect 1699 966 1705 967
rect 1907 967 1908 971
rect 1912 970 1913 971
rect 1912 968 2001 970
rect 2003 969 2004 973
rect 2011 971 2012 975
rect 2021 974 2023 982
rect 2224 974 2226 984
rect 2230 983 2231 987
rect 2235 983 2236 987
rect 2230 982 2236 983
rect 2246 987 2257 988
rect 2246 983 2247 987
rect 2251 983 2252 987
rect 2256 983 2257 987
rect 2246 982 2257 983
rect 2350 987 2356 988
rect 2350 983 2351 987
rect 2355 983 2356 987
rect 2350 982 2356 983
rect 2371 987 2377 988
rect 2371 983 2372 987
rect 2376 986 2377 987
rect 2430 987 2436 988
rect 2430 986 2431 987
rect 2376 984 2431 986
rect 2376 983 2377 984
rect 2371 982 2377 983
rect 2430 983 2431 984
rect 2435 983 2436 987
rect 2430 982 2436 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2454 982 2460 983
rect 2475 987 2484 988
rect 2475 983 2476 987
rect 2483 983 2484 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2475 982 2484 983
rect 2021 973 2121 974
rect 2021 972 2116 973
rect 2008 970 2012 971
rect 2008 969 2009 970
rect 2003 968 2009 969
rect 2115 969 2116 972
rect 2120 969 2121 973
rect 2224 973 2241 974
rect 2224 972 2236 973
rect 2115 968 2121 969
rect 2235 969 2236 972
rect 2240 969 2241 973
rect 2235 968 2241 969
rect 2355 971 2361 972
rect 1912 967 1913 968
rect 1907 966 1913 967
rect 1999 966 2001 968
rect 2246 967 2252 968
rect 2246 966 2247 967
rect 1999 964 2247 966
rect 1598 962 1604 963
rect 2246 963 2247 964
rect 2251 963 2252 967
rect 2355 967 2356 971
rect 2360 970 2361 971
rect 2446 971 2452 972
rect 2446 970 2447 971
rect 2360 968 2447 970
rect 2360 967 2361 968
rect 2355 966 2361 967
rect 2446 967 2447 968
rect 2451 967 2452 971
rect 2446 966 2452 967
rect 2459 971 2468 972
rect 2459 967 2460 971
rect 2467 967 2468 971
rect 2459 966 2468 967
rect 2246 962 2252 963
rect 1035 961 1041 962
rect 854 959 860 960
rect 854 955 855 959
rect 859 958 860 959
rect 867 959 873 960
rect 867 958 868 959
rect 859 956 868 958
rect 859 955 860 956
rect 854 954 860 955
rect 867 955 868 956
rect 872 955 873 959
rect 867 954 873 955
rect 955 959 961 960
rect 955 955 956 959
rect 960 958 961 959
rect 960 956 1006 958
rect 1035 957 1036 961
rect 1040 957 1041 961
rect 1232 961 1249 962
rect 1232 960 1244 961
rect 1035 956 1041 957
rect 1107 959 1113 960
rect 960 955 961 956
rect 955 954 961 955
rect 1004 954 1006 956
rect 1046 955 1052 956
rect 1046 954 1047 955
rect 772 952 790 954
rect 1004 952 1047 954
rect 574 951 580 952
rect 574 950 575 951
rect 319 948 575 950
rect 574 947 575 948
rect 579 947 580 951
rect 1046 951 1047 952
rect 1051 951 1052 955
rect 1107 955 1108 959
rect 1112 958 1113 959
rect 1187 959 1196 960
rect 1112 956 1161 958
rect 1112 955 1113 956
rect 1107 954 1113 955
rect 1046 950 1052 951
rect 1159 950 1161 956
rect 1187 955 1188 959
rect 1195 955 1196 959
rect 1243 957 1244 960
rect 1248 957 1249 961
rect 1243 956 1249 957
rect 1187 954 1196 955
rect 1246 951 1252 952
rect 1246 950 1247 951
rect 1159 948 1247 950
rect 574 946 580 947
rect 766 947 772 948
rect 766 946 767 947
rect 740 944 767 946
rect 740 942 742 944
rect 766 943 767 944
rect 771 943 772 947
rect 1246 947 1247 948
rect 1251 947 1252 951
rect 1246 946 1252 947
rect 766 942 772 943
rect 1534 943 1540 944
rect 1534 942 1535 943
rect 739 941 745 942
rect 155 939 164 940
rect 155 935 156 939
rect 163 935 164 939
rect 211 939 217 940
rect 211 938 212 939
rect 155 934 164 935
rect 173 936 212 938
rect 173 926 175 936
rect 211 935 212 936
rect 216 935 217 939
rect 299 939 305 940
rect 299 938 300 939
rect 211 934 217 935
rect 228 936 300 938
rect 228 926 230 936
rect 299 935 300 936
rect 304 935 305 939
rect 403 939 409 940
rect 403 938 404 939
rect 299 934 305 935
rect 319 936 404 938
rect 319 926 321 936
rect 403 935 404 936
rect 408 935 409 939
rect 515 939 521 940
rect 515 938 516 939
rect 403 934 409 935
rect 420 936 516 938
rect 420 926 422 936
rect 515 935 516 936
rect 520 935 521 939
rect 515 934 521 935
rect 534 939 540 940
rect 534 935 535 939
rect 539 938 540 939
rect 627 939 633 940
rect 627 938 628 939
rect 539 936 628 938
rect 539 935 540 936
rect 534 934 540 935
rect 627 935 628 936
rect 632 935 633 939
rect 739 937 740 941
rect 744 937 745 941
rect 1444 940 1535 942
rect 835 939 841 940
rect 835 938 836 939
rect 739 936 745 937
rect 756 936 836 938
rect 627 934 633 935
rect 430 931 436 932
rect 430 927 431 931
rect 435 930 436 931
rect 435 928 646 930
rect 435 927 436 928
rect 430 926 436 927
rect 644 926 646 928
rect 756 926 758 936
rect 835 935 836 936
rect 840 935 841 939
rect 835 934 841 935
rect 918 939 924 940
rect 918 935 919 939
rect 923 938 924 939
rect 931 939 937 940
rect 931 938 932 939
rect 923 936 932 938
rect 923 935 924 936
rect 918 934 924 935
rect 931 935 932 936
rect 936 935 937 939
rect 1019 939 1025 940
rect 1019 938 1020 939
rect 931 934 937 935
rect 988 936 1020 938
rect 988 930 990 936
rect 1019 935 1020 936
rect 1024 935 1025 939
rect 1099 939 1105 940
rect 1099 938 1100 939
rect 1019 934 1025 935
rect 1036 936 1100 938
rect 948 928 990 930
rect 948 926 950 928
rect 1036 926 1038 936
rect 1099 935 1100 936
rect 1104 935 1105 939
rect 1099 934 1105 935
rect 1179 939 1185 940
rect 1179 935 1180 939
rect 1184 938 1185 939
rect 1243 939 1252 940
rect 1184 936 1239 938
rect 1184 935 1185 936
rect 1179 934 1185 935
rect 1237 930 1239 936
rect 1243 935 1244 939
rect 1251 935 1252 939
rect 1243 934 1252 935
rect 1262 939 1268 940
rect 1262 935 1263 939
rect 1267 938 1268 939
rect 1444 938 1446 940
rect 1534 939 1535 940
rect 1539 939 1540 943
rect 1534 938 1540 939
rect 1267 937 1377 938
rect 1267 936 1372 937
rect 1267 935 1268 936
rect 1262 934 1268 935
rect 1371 933 1372 936
rect 1376 933 1377 937
rect 1371 932 1377 933
rect 1443 937 1449 938
rect 1443 933 1444 937
rect 1448 933 1449 937
rect 1531 935 1537 936
rect 1531 934 1532 935
rect 1443 932 1449 933
rect 1461 932 1532 934
rect 1237 928 1366 930
rect 1364 926 1366 928
rect 150 925 156 926
rect 110 924 116 925
rect 110 920 111 924
rect 115 920 116 924
rect 150 921 151 925
rect 155 921 156 925
rect 150 920 156 921
rect 171 925 177 926
rect 171 921 172 925
rect 176 921 177 925
rect 171 920 177 921
rect 206 925 212 926
rect 206 921 207 925
rect 211 921 212 925
rect 206 920 212 921
rect 227 925 233 926
rect 227 921 228 925
rect 232 921 233 925
rect 227 920 233 921
rect 294 925 300 926
rect 294 921 295 925
rect 299 921 300 925
rect 294 920 300 921
rect 315 925 321 926
rect 315 921 316 925
rect 320 921 321 925
rect 315 920 321 921
rect 398 925 404 926
rect 398 921 399 925
rect 403 921 404 925
rect 398 920 404 921
rect 419 925 425 926
rect 419 921 420 925
rect 424 921 425 925
rect 419 920 425 921
rect 510 925 516 926
rect 510 921 511 925
rect 515 921 516 925
rect 622 925 628 926
rect 510 920 516 921
rect 531 923 540 924
rect 110 919 116 920
rect 531 919 532 923
rect 539 919 540 923
rect 622 921 623 925
rect 627 921 628 925
rect 622 920 628 921
rect 643 925 649 926
rect 643 921 644 925
rect 648 921 649 925
rect 643 920 649 921
rect 734 925 740 926
rect 734 921 735 925
rect 739 921 740 925
rect 734 920 740 921
rect 755 925 761 926
rect 755 921 756 925
rect 760 921 761 925
rect 755 920 761 921
rect 830 925 836 926
rect 830 921 831 925
rect 835 921 836 925
rect 926 925 932 926
rect 830 920 836 921
rect 851 923 860 924
rect 531 918 540 919
rect 851 919 852 923
rect 859 919 860 923
rect 926 921 927 925
rect 931 921 932 925
rect 926 920 932 921
rect 947 925 953 926
rect 947 921 948 925
rect 952 921 953 925
rect 947 920 953 921
rect 1014 925 1020 926
rect 1014 921 1015 925
rect 1019 921 1020 925
rect 1014 920 1020 921
rect 1035 925 1041 926
rect 1035 921 1036 925
rect 1040 921 1041 925
rect 1035 920 1041 921
rect 1094 925 1100 926
rect 1094 921 1095 925
rect 1099 921 1100 925
rect 1174 925 1180 926
rect 1094 920 1100 921
rect 1115 923 1124 924
rect 851 918 860 919
rect 1115 919 1116 923
rect 1123 919 1124 923
rect 1174 921 1175 925
rect 1179 921 1180 925
rect 1238 925 1244 926
rect 1174 920 1180 921
rect 1190 923 1201 924
rect 1115 918 1124 919
rect 1190 919 1191 923
rect 1195 919 1196 923
rect 1200 919 1201 923
rect 1238 921 1239 925
rect 1243 921 1244 925
rect 1286 924 1292 925
rect 1364 924 1391 926
rect 1238 920 1244 921
rect 1259 923 1268 924
rect 1190 918 1201 919
rect 1259 919 1260 923
rect 1267 919 1268 923
rect 1286 920 1287 924
rect 1291 920 1292 924
rect 1389 922 1391 924
rect 1461 922 1463 932
rect 1531 931 1532 932
rect 1536 931 1537 935
rect 1531 930 1537 931
rect 1619 935 1625 936
rect 1619 931 1620 935
rect 1624 934 1625 935
rect 1699 935 1705 936
rect 1624 932 1694 934
rect 1624 931 1625 932
rect 1619 930 1625 931
rect 1692 926 1694 932
rect 1699 931 1700 935
rect 1704 934 1705 935
rect 1722 935 1728 936
rect 1722 934 1723 935
rect 1704 932 1723 934
rect 1704 931 1705 932
rect 1699 930 1705 931
rect 1722 931 1723 932
rect 1727 931 1728 935
rect 1722 930 1728 931
rect 1782 935 1788 936
rect 1782 931 1783 935
rect 1787 934 1788 935
rect 1795 935 1801 936
rect 1795 934 1796 935
rect 1787 932 1796 934
rect 1787 931 1788 932
rect 1782 930 1788 931
rect 1795 931 1796 932
rect 1800 931 1801 935
rect 1899 935 1905 936
rect 1899 934 1900 935
rect 1795 930 1801 931
rect 1812 932 1900 934
rect 1692 924 1718 926
rect 1716 922 1718 924
rect 1812 922 1814 932
rect 1899 931 1900 932
rect 1904 931 1905 935
rect 2019 935 2025 936
rect 2019 934 2020 935
rect 1899 930 1905 931
rect 1999 932 2020 934
rect 1999 926 2001 932
rect 2019 931 2020 932
rect 2024 931 2025 935
rect 2155 935 2161 936
rect 2155 934 2156 935
rect 2019 930 2025 931
rect 2036 932 2156 934
rect 1916 924 2001 926
rect 1916 922 1918 924
rect 2036 922 2038 932
rect 2155 931 2156 932
rect 2160 931 2161 935
rect 2299 935 2305 936
rect 2299 934 2300 935
rect 2155 930 2161 931
rect 2172 932 2300 934
rect 2172 922 2174 932
rect 2299 931 2300 932
rect 2304 931 2305 935
rect 2299 930 2305 931
rect 2406 935 2412 936
rect 2406 931 2407 935
rect 2411 934 2412 935
rect 2443 935 2449 936
rect 2443 934 2444 935
rect 2411 932 2444 934
rect 2411 931 2412 932
rect 2406 930 2412 931
rect 2443 931 2444 932
rect 2448 931 2449 935
rect 2443 930 2449 931
rect 1366 921 1372 922
rect 1286 919 1292 920
rect 1326 920 1332 921
rect 1259 918 1268 919
rect 1326 916 1327 920
rect 1331 916 1332 920
rect 1366 917 1367 921
rect 1371 917 1372 921
rect 1366 916 1372 917
rect 1387 921 1393 922
rect 1387 917 1388 921
rect 1392 917 1393 921
rect 1387 916 1393 917
rect 1438 921 1444 922
rect 1438 917 1439 921
rect 1443 917 1444 921
rect 1438 916 1444 917
rect 1459 921 1465 922
rect 1459 917 1460 921
rect 1464 917 1465 921
rect 1459 916 1465 917
rect 1526 921 1532 922
rect 1526 917 1527 921
rect 1531 917 1532 921
rect 1614 921 1620 922
rect 1526 916 1532 917
rect 1547 919 1553 920
rect 1326 915 1332 916
rect 1547 915 1548 919
rect 1552 918 1553 919
rect 1566 919 1572 920
rect 1566 918 1567 919
rect 1552 916 1567 918
rect 1552 915 1553 916
rect 1547 914 1553 915
rect 1566 915 1567 916
rect 1571 915 1572 919
rect 1614 917 1615 921
rect 1619 917 1620 921
rect 1694 921 1700 922
rect 1614 916 1620 917
rect 1635 919 1641 920
rect 1566 914 1572 915
rect 1635 915 1636 919
rect 1640 918 1641 919
rect 1654 919 1660 920
rect 1654 918 1655 919
rect 1640 916 1655 918
rect 1640 915 1641 916
rect 1635 914 1641 915
rect 1654 915 1655 916
rect 1659 915 1660 919
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1715 921 1721 922
rect 1715 917 1716 921
rect 1720 917 1721 921
rect 1715 916 1721 917
rect 1790 921 1796 922
rect 1790 917 1791 921
rect 1795 917 1796 921
rect 1790 916 1796 917
rect 1811 921 1817 922
rect 1811 917 1812 921
rect 1816 917 1817 921
rect 1811 916 1817 917
rect 1894 921 1900 922
rect 1894 917 1895 921
rect 1899 917 1900 921
rect 1894 916 1900 917
rect 1915 921 1921 922
rect 1915 917 1916 921
rect 1920 917 1921 921
rect 1915 916 1921 917
rect 2014 921 2020 922
rect 2014 917 2015 921
rect 2019 917 2020 921
rect 2014 916 2020 917
rect 2035 921 2041 922
rect 2035 917 2036 921
rect 2040 917 2041 921
rect 2035 916 2041 917
rect 2150 921 2156 922
rect 2150 917 2151 921
rect 2155 917 2156 921
rect 2150 916 2156 917
rect 2171 921 2177 922
rect 2171 917 2172 921
rect 2176 917 2177 921
rect 2171 916 2177 917
rect 2294 921 2300 922
rect 2294 917 2295 921
rect 2299 917 2300 921
rect 2438 921 2444 922
rect 2294 916 2300 917
rect 2302 919 2308 920
rect 1654 914 1660 915
rect 2302 915 2303 919
rect 2307 918 2308 919
rect 2315 919 2321 920
rect 2315 918 2316 919
rect 2307 916 2316 918
rect 2307 915 2308 916
rect 2302 914 2308 915
rect 2315 915 2316 916
rect 2320 915 2321 919
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2502 920 2508 921
rect 2438 916 2444 917
rect 2446 919 2452 920
rect 2315 914 2321 915
rect 2446 915 2447 919
rect 2451 918 2452 919
rect 2459 919 2465 920
rect 2459 918 2460 919
rect 2451 916 2460 918
rect 2451 915 2452 916
rect 2446 914 2452 915
rect 2459 915 2460 916
rect 2464 915 2465 919
rect 2502 916 2503 920
rect 2507 916 2508 920
rect 2502 915 2508 916
rect 2459 914 2465 915
rect 110 907 116 908
rect 110 903 111 907
rect 115 903 116 907
rect 1286 907 1292 908
rect 110 902 116 903
rect 134 904 140 905
rect 134 900 135 904
rect 139 900 140 904
rect 134 899 140 900
rect 190 904 196 905
rect 190 900 191 904
rect 195 900 196 904
rect 190 899 196 900
rect 278 904 284 905
rect 278 900 279 904
rect 283 900 284 904
rect 278 899 284 900
rect 382 904 388 905
rect 382 900 383 904
rect 387 900 388 904
rect 382 899 388 900
rect 494 904 500 905
rect 494 900 495 904
rect 499 900 500 904
rect 494 899 500 900
rect 606 904 612 905
rect 606 900 607 904
rect 611 900 612 904
rect 606 899 612 900
rect 718 904 724 905
rect 718 900 719 904
rect 723 900 724 904
rect 718 899 724 900
rect 814 904 820 905
rect 814 900 815 904
rect 819 900 820 904
rect 814 899 820 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 998 904 1004 905
rect 998 900 999 904
rect 1003 900 1004 904
rect 998 899 1004 900
rect 1078 904 1084 905
rect 1078 900 1079 904
rect 1083 900 1084 904
rect 1078 899 1084 900
rect 1158 904 1164 905
rect 1158 900 1159 904
rect 1163 900 1164 904
rect 1158 899 1164 900
rect 1222 904 1228 905
rect 1222 900 1223 904
rect 1227 900 1228 904
rect 1286 903 1287 907
rect 1291 903 1292 907
rect 1286 902 1292 903
rect 1326 903 1332 904
rect 1222 899 1228 900
rect 1326 899 1327 903
rect 1331 899 1332 903
rect 2502 903 2508 904
rect 1326 898 1332 899
rect 1350 900 1356 901
rect 1350 896 1351 900
rect 1355 896 1356 900
rect 1350 895 1356 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1510 900 1516 901
rect 1510 896 1511 900
rect 1515 896 1516 900
rect 1510 895 1516 896
rect 1598 900 1604 901
rect 1598 896 1599 900
rect 1603 896 1604 900
rect 1598 895 1604 896
rect 1678 900 1684 901
rect 1678 896 1679 900
rect 1683 896 1684 900
rect 1678 895 1684 896
rect 1774 900 1780 901
rect 1774 896 1775 900
rect 1779 896 1780 900
rect 1774 895 1780 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1998 900 2004 901
rect 1998 896 1999 900
rect 2003 896 2004 900
rect 1998 895 2004 896
rect 2134 900 2140 901
rect 2134 896 2135 900
rect 2139 896 2140 900
rect 2134 895 2140 896
rect 2278 900 2284 901
rect 2278 896 2279 900
rect 2283 896 2284 900
rect 2278 895 2284 896
rect 2422 900 2428 901
rect 2422 896 2423 900
rect 2427 896 2428 900
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2422 895 2428 896
rect 246 888 252 889
rect 110 885 116 886
rect 110 881 111 885
rect 115 881 116 885
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 342 888 348 889
rect 342 884 343 888
rect 347 884 348 888
rect 342 883 348 884
rect 438 888 444 889
rect 438 884 439 888
rect 443 884 444 888
rect 438 883 444 884
rect 542 888 548 889
rect 542 884 543 888
rect 547 884 548 888
rect 542 883 548 884
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 742 888 748 889
rect 742 884 743 888
rect 747 884 748 888
rect 742 883 748 884
rect 838 888 844 889
rect 838 884 839 888
rect 843 884 844 888
rect 838 883 844 884
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 1006 888 1012 889
rect 1006 884 1007 888
rect 1011 884 1012 888
rect 1006 883 1012 884
rect 1086 888 1092 889
rect 1086 884 1087 888
rect 1091 884 1092 888
rect 1086 883 1092 884
rect 1166 888 1172 889
rect 1166 884 1167 888
rect 1171 884 1172 888
rect 1166 883 1172 884
rect 1222 888 1228 889
rect 1222 884 1223 888
rect 1227 884 1228 888
rect 1222 883 1228 884
rect 1286 885 1292 886
rect 110 880 116 881
rect 1286 881 1287 885
rect 1291 881 1292 885
rect 1286 880 1292 881
rect 1486 880 1492 881
rect 1326 877 1332 878
rect 1326 873 1327 877
rect 1331 873 1332 877
rect 1486 876 1487 880
rect 1491 876 1492 880
rect 1486 875 1492 876
rect 1558 880 1564 881
rect 1558 876 1559 880
rect 1563 876 1564 880
rect 1558 875 1564 876
rect 1622 880 1628 881
rect 1622 876 1623 880
rect 1627 876 1628 880
rect 1622 875 1628 876
rect 1686 880 1692 881
rect 1686 876 1687 880
rect 1691 876 1692 880
rect 1686 875 1692 876
rect 1750 880 1756 881
rect 1750 876 1751 880
rect 1755 876 1756 880
rect 1750 875 1756 876
rect 1814 880 1820 881
rect 1814 876 1815 880
rect 1819 876 1820 880
rect 1814 875 1820 876
rect 1886 880 1892 881
rect 1886 876 1887 880
rect 1891 876 1892 880
rect 1886 875 1892 876
rect 1974 880 1980 881
rect 1974 876 1975 880
rect 1979 876 1980 880
rect 1974 875 1980 876
rect 2078 880 2084 881
rect 2078 876 2079 880
rect 2083 876 2084 880
rect 2078 875 2084 876
rect 2198 880 2204 881
rect 2198 876 2199 880
rect 2203 876 2204 880
rect 2198 875 2204 876
rect 2318 880 2324 881
rect 2318 876 2319 880
rect 2323 876 2324 880
rect 2318 875 2324 876
rect 2438 880 2444 881
rect 2438 876 2439 880
rect 2443 876 2444 880
rect 2438 875 2444 876
rect 2502 877 2508 878
rect 1326 872 1332 873
rect 2502 873 2503 877
rect 2507 873 2508 877
rect 2502 872 2508 873
rect 110 868 116 869
rect 1286 868 1292 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 262 867 268 868
rect 262 863 263 867
rect 267 863 268 867
rect 262 862 268 863
rect 283 867 289 868
rect 283 863 284 867
rect 288 866 289 867
rect 358 867 364 868
rect 288 864 321 866
rect 288 863 289 864
rect 283 862 289 863
rect 319 854 321 864
rect 358 863 359 867
rect 363 863 364 867
rect 358 862 364 863
rect 379 867 385 868
rect 379 863 380 867
rect 384 866 385 867
rect 454 867 460 868
rect 384 864 450 866
rect 384 863 385 864
rect 379 862 385 863
rect 448 854 450 864
rect 454 863 455 867
rect 459 863 460 867
rect 454 862 460 863
rect 475 867 481 868
rect 475 863 476 867
rect 480 866 481 867
rect 558 867 564 868
rect 480 864 554 866
rect 480 863 481 864
rect 475 862 481 863
rect 552 854 554 864
rect 558 863 559 867
rect 563 863 564 867
rect 558 862 564 863
rect 579 867 585 868
rect 579 863 580 867
rect 584 866 585 867
rect 662 867 668 868
rect 584 864 658 866
rect 584 863 585 864
rect 579 862 585 863
rect 656 854 658 864
rect 662 863 663 867
rect 667 863 668 867
rect 662 862 668 863
rect 670 867 676 868
rect 670 863 671 867
rect 675 866 676 867
rect 683 867 689 868
rect 683 866 684 867
rect 675 864 684 866
rect 675 863 676 864
rect 670 862 676 863
rect 683 863 684 864
rect 688 863 689 867
rect 683 862 689 863
rect 758 867 764 868
rect 758 863 759 867
rect 763 863 764 867
rect 758 862 764 863
rect 766 867 772 868
rect 766 863 767 867
rect 771 866 772 867
rect 779 867 785 868
rect 779 866 780 867
rect 771 864 780 866
rect 771 863 772 864
rect 766 862 772 863
rect 779 863 780 864
rect 784 863 785 867
rect 779 862 785 863
rect 854 867 860 868
rect 854 863 855 867
rect 859 863 860 867
rect 854 862 860 863
rect 875 867 881 868
rect 875 863 876 867
rect 880 866 881 867
rect 942 867 948 868
rect 880 864 934 866
rect 880 863 881 864
rect 875 862 881 863
rect 932 854 934 864
rect 942 863 943 867
rect 947 863 948 867
rect 942 862 948 863
rect 963 867 969 868
rect 963 863 964 867
rect 968 866 969 867
rect 1022 867 1028 868
rect 968 864 1018 866
rect 968 863 969 864
rect 963 862 969 863
rect 1016 854 1018 864
rect 1022 863 1023 867
rect 1027 863 1028 867
rect 1022 862 1028 863
rect 1043 867 1049 868
rect 1043 863 1044 867
rect 1048 866 1049 867
rect 1102 867 1108 868
rect 1048 864 1098 866
rect 1048 863 1049 864
rect 1043 862 1049 863
rect 1096 854 1098 864
rect 1102 863 1103 867
rect 1107 863 1108 867
rect 1102 862 1108 863
rect 1123 867 1129 868
rect 1123 863 1124 867
rect 1128 866 1129 867
rect 1182 867 1188 868
rect 1128 864 1161 866
rect 1128 863 1129 864
rect 1123 862 1129 863
rect 1159 854 1161 864
rect 1182 863 1183 867
rect 1187 863 1188 867
rect 1182 862 1188 863
rect 1203 867 1209 868
rect 1203 863 1204 867
rect 1208 866 1209 867
rect 1238 867 1244 868
rect 1208 864 1234 866
rect 1208 863 1209 864
rect 1203 862 1209 863
rect 1232 854 1234 864
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 1238 862 1244 863
rect 1246 867 1252 868
rect 1246 863 1247 867
rect 1251 866 1252 867
rect 1259 867 1265 868
rect 1259 866 1260 867
rect 1251 864 1260 866
rect 1251 863 1252 864
rect 1246 862 1252 863
rect 1259 863 1260 864
rect 1264 863 1265 867
rect 1286 864 1287 868
rect 1291 864 1292 868
rect 1286 863 1292 864
rect 1259 862 1265 863
rect 1326 860 1332 861
rect 2502 860 2508 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1502 859 1508 860
rect 1502 855 1503 859
rect 1507 855 1508 859
rect 1502 854 1508 855
rect 1518 859 1529 860
rect 1518 855 1519 859
rect 1523 855 1524 859
rect 1528 855 1529 859
rect 1518 854 1529 855
rect 1574 859 1580 860
rect 1574 855 1575 859
rect 1579 855 1580 859
rect 1574 854 1580 855
rect 1595 859 1601 860
rect 1595 855 1596 859
rect 1600 858 1601 859
rect 1638 859 1644 860
rect 1600 856 1626 858
rect 1600 855 1601 856
rect 1595 854 1601 855
rect 319 853 369 854
rect 319 852 364 853
rect 267 851 273 852
rect 267 847 268 851
rect 272 850 273 851
rect 272 848 321 850
rect 363 849 364 852
rect 368 849 369 853
rect 448 853 465 854
rect 448 852 460 853
rect 363 848 369 849
rect 459 849 460 852
rect 464 849 465 853
rect 552 853 569 854
rect 552 852 564 853
rect 459 848 465 849
rect 563 849 564 852
rect 568 849 569 853
rect 656 853 673 854
rect 656 852 668 853
rect 563 848 569 849
rect 667 849 668 852
rect 672 849 673 853
rect 932 853 953 854
rect 932 852 948 853
rect 667 848 673 849
rect 763 851 769 852
rect 272 847 273 848
rect 267 846 273 847
rect 319 846 321 848
rect 430 847 436 848
rect 430 846 431 847
rect 319 844 431 846
rect 430 843 431 844
rect 435 843 436 847
rect 763 847 764 851
rect 768 850 769 851
rect 859 851 865 852
rect 768 848 854 850
rect 768 847 769 848
rect 763 846 769 847
rect 430 842 436 843
rect 852 838 854 848
rect 859 847 860 851
rect 864 850 865 851
rect 864 848 942 850
rect 947 849 948 852
rect 952 849 953 853
rect 1016 853 1033 854
rect 1016 852 1028 853
rect 947 848 953 849
rect 1027 849 1028 852
rect 1032 849 1033 853
rect 1096 853 1113 854
rect 1096 852 1108 853
rect 1027 848 1033 849
rect 1107 849 1108 852
rect 1112 849 1113 853
rect 1159 853 1193 854
rect 1159 852 1188 853
rect 1107 848 1113 849
rect 1187 849 1188 852
rect 1192 849 1193 853
rect 1232 853 1249 854
rect 1232 852 1244 853
rect 1187 848 1193 849
rect 1243 849 1244 852
rect 1248 849 1249 853
rect 1243 848 1249 849
rect 864 847 865 848
rect 859 846 865 847
rect 940 846 942 848
rect 1118 847 1124 848
rect 1118 846 1119 847
rect 940 844 1119 846
rect 1118 843 1119 844
rect 1123 843 1124 847
rect 1624 846 1626 856
rect 1638 855 1639 859
rect 1643 855 1644 859
rect 1638 854 1644 855
rect 1646 859 1652 860
rect 1646 855 1647 859
rect 1651 858 1652 859
rect 1659 859 1665 860
rect 1659 858 1660 859
rect 1651 856 1660 858
rect 1651 855 1652 856
rect 1646 854 1652 855
rect 1659 855 1660 856
rect 1664 855 1665 859
rect 1659 854 1665 855
rect 1702 859 1708 860
rect 1702 855 1703 859
rect 1707 855 1708 859
rect 1702 854 1708 855
rect 1722 859 1729 860
rect 1722 855 1723 859
rect 1728 855 1729 859
rect 1722 854 1729 855
rect 1766 859 1772 860
rect 1766 855 1767 859
rect 1771 855 1772 859
rect 1787 859 1793 860
rect 1787 858 1788 859
rect 1766 854 1772 855
rect 1776 856 1788 858
rect 1776 850 1778 856
rect 1787 855 1788 856
rect 1792 855 1793 859
rect 1787 854 1793 855
rect 1830 859 1836 860
rect 1830 855 1831 859
rect 1835 855 1836 859
rect 1830 854 1836 855
rect 1851 859 1857 860
rect 1851 855 1852 859
rect 1856 858 1857 859
rect 1902 859 1908 860
rect 1856 856 1898 858
rect 1856 855 1857 856
rect 1851 854 1857 855
rect 1708 848 1778 850
rect 1708 846 1710 848
rect 1896 846 1898 856
rect 1902 855 1903 859
rect 1907 855 1908 859
rect 1902 854 1908 855
rect 1923 859 1929 860
rect 1923 855 1924 859
rect 1928 855 1929 859
rect 1923 854 1929 855
rect 1990 859 1996 860
rect 1990 855 1991 859
rect 1995 855 1996 859
rect 1990 854 1996 855
rect 2011 859 2017 860
rect 2011 855 2012 859
rect 2016 858 2017 859
rect 2094 859 2100 860
rect 2016 856 2090 858
rect 2016 855 2017 856
rect 2011 854 2017 855
rect 1925 846 1927 854
rect 2088 846 2090 856
rect 2094 855 2095 859
rect 2099 855 2100 859
rect 2094 854 2100 855
rect 2115 859 2121 860
rect 2115 855 2116 859
rect 2120 858 2121 859
rect 2214 859 2220 860
rect 2120 856 2210 858
rect 2120 855 2121 856
rect 2115 854 2121 855
rect 2208 846 2210 856
rect 2214 855 2215 859
rect 2219 855 2220 859
rect 2214 854 2220 855
rect 2235 859 2241 860
rect 2235 855 2236 859
rect 2240 855 2241 859
rect 2235 854 2241 855
rect 2334 859 2340 860
rect 2334 855 2335 859
rect 2339 855 2340 859
rect 2334 854 2340 855
rect 2342 859 2348 860
rect 2342 855 2343 859
rect 2347 858 2348 859
rect 2355 859 2361 860
rect 2355 858 2356 859
rect 2347 856 2356 858
rect 2347 855 2348 856
rect 2342 854 2348 855
rect 2355 855 2356 856
rect 2360 855 2361 859
rect 2355 854 2361 855
rect 2454 859 2460 860
rect 2454 855 2455 859
rect 2459 855 2460 859
rect 2454 854 2460 855
rect 2462 859 2468 860
rect 2462 855 2463 859
rect 2467 858 2468 859
rect 2475 859 2481 860
rect 2475 858 2476 859
rect 2467 856 2476 858
rect 2467 855 2468 856
rect 2462 854 2468 855
rect 2475 855 2476 856
rect 2480 855 2481 859
rect 2502 856 2503 860
rect 2507 856 2508 860
rect 2502 855 2508 856
rect 2475 854 2481 855
rect 2237 846 2239 854
rect 1624 845 1649 846
rect 1624 844 1644 845
rect 1118 842 1124 843
rect 1507 843 1513 844
rect 1090 839 1096 840
rect 1090 838 1091 839
rect 852 836 1091 838
rect 402 835 408 836
rect 402 834 403 835
rect 244 832 403 834
rect 244 830 246 832
rect 402 831 403 832
rect 407 831 408 835
rect 1090 835 1091 836
rect 1095 835 1096 839
rect 1507 839 1508 843
rect 1512 842 1513 843
rect 1566 843 1572 844
rect 1512 840 1562 842
rect 1512 839 1513 840
rect 1507 838 1513 839
rect 1090 834 1096 835
rect 1560 834 1562 840
rect 1566 839 1567 843
rect 1571 842 1572 843
rect 1579 843 1585 844
rect 1579 842 1580 843
rect 1571 840 1580 842
rect 1571 839 1572 840
rect 1566 838 1572 839
rect 1579 839 1580 840
rect 1584 839 1585 843
rect 1643 841 1644 844
rect 1648 841 1649 845
rect 1643 840 1649 841
rect 1707 845 1713 846
rect 1707 841 1708 845
rect 1712 841 1713 845
rect 1896 845 1913 846
rect 1896 844 1908 845
rect 1707 840 1713 841
rect 1771 843 1777 844
rect 1579 838 1585 839
rect 1771 839 1772 843
rect 1776 842 1777 843
rect 1818 843 1824 844
rect 1818 842 1819 843
rect 1776 840 1819 842
rect 1776 839 1777 840
rect 1771 838 1777 839
rect 1818 839 1819 840
rect 1823 839 1824 843
rect 1818 838 1824 839
rect 1835 843 1844 844
rect 1835 839 1836 843
rect 1843 839 1844 843
rect 1907 841 1908 844
rect 1912 841 1913 845
rect 1925 845 2001 846
rect 1925 844 1996 845
rect 1907 840 1913 841
rect 1995 841 1996 844
rect 2000 841 2001 845
rect 2088 845 2105 846
rect 2088 844 2100 845
rect 1995 840 2001 841
rect 2099 841 2100 844
rect 2104 841 2105 845
rect 2208 845 2225 846
rect 2208 844 2220 845
rect 2099 840 2105 841
rect 2219 841 2220 844
rect 2224 841 2225 845
rect 2237 845 2345 846
rect 2237 844 2340 845
rect 2219 840 2225 841
rect 2339 841 2340 844
rect 2344 841 2345 845
rect 2339 840 2345 841
rect 2430 843 2436 844
rect 1835 838 1844 839
rect 2430 839 2431 843
rect 2435 842 2436 843
rect 2459 843 2465 844
rect 2459 842 2460 843
rect 2435 840 2460 842
rect 2435 839 2436 840
rect 2430 838 2436 839
rect 2459 839 2460 840
rect 2464 839 2465 843
rect 2459 838 2465 839
rect 1646 835 1652 836
rect 1646 834 1647 835
rect 1560 832 1647 834
rect 402 830 408 831
rect 1646 831 1647 832
rect 1651 831 1652 835
rect 1646 830 1652 831
rect 243 829 249 830
rect 243 825 244 829
rect 248 825 249 829
rect 307 827 313 828
rect 307 826 308 827
rect 243 824 249 825
rect 284 824 308 826
rect 284 814 286 824
rect 307 823 308 824
rect 312 823 313 827
rect 307 822 313 823
rect 387 827 393 828
rect 387 823 388 827
rect 392 826 393 827
rect 467 827 473 828
rect 392 824 462 826
rect 392 823 393 824
rect 387 822 393 823
rect 460 818 462 824
rect 467 823 468 827
rect 472 826 473 827
rect 555 827 561 828
rect 472 824 550 826
rect 472 823 473 824
rect 467 822 473 823
rect 548 818 550 824
rect 555 823 556 827
rect 560 826 561 827
rect 643 827 649 828
rect 560 824 638 826
rect 560 823 561 824
rect 555 822 561 823
rect 636 818 638 824
rect 643 823 644 827
rect 648 826 649 827
rect 670 827 676 828
rect 670 826 671 827
rect 648 824 671 826
rect 648 823 649 824
rect 643 822 649 823
rect 670 823 671 824
rect 675 823 676 827
rect 670 822 676 823
rect 731 827 737 828
rect 731 823 732 827
rect 736 826 737 827
rect 762 827 768 828
rect 762 826 763 827
rect 736 824 763 826
rect 736 823 737 824
rect 731 822 737 823
rect 762 823 763 824
rect 767 823 768 827
rect 811 827 817 828
rect 811 826 812 827
rect 762 822 768 823
rect 772 824 812 826
rect 772 818 774 824
rect 811 823 812 824
rect 816 823 817 827
rect 899 827 905 828
rect 899 826 900 827
rect 811 822 817 823
rect 829 824 900 826
rect 460 816 486 818
rect 548 816 574 818
rect 636 816 662 818
rect 484 814 486 816
rect 572 814 574 816
rect 660 814 662 816
rect 748 816 774 818
rect 748 814 750 816
rect 829 814 831 824
rect 899 823 900 824
rect 904 823 905 827
rect 987 827 993 828
rect 987 826 988 827
rect 899 822 905 823
rect 916 824 988 826
rect 916 814 918 824
rect 987 823 988 824
rect 992 823 993 827
rect 1075 827 1081 828
rect 1075 826 1076 827
rect 987 822 993 823
rect 1004 824 1076 826
rect 1004 814 1006 824
rect 1075 823 1076 824
rect 1080 823 1081 827
rect 1075 822 1081 823
rect 1518 823 1524 824
rect 1518 822 1519 823
rect 1444 820 1519 822
rect 1444 818 1446 820
rect 1518 819 1519 820
rect 1523 819 1524 823
rect 1722 823 1728 824
rect 1722 822 1723 823
rect 1518 818 1524 819
rect 1676 820 1723 822
rect 1676 818 1678 820
rect 1722 819 1723 820
rect 1727 819 1728 823
rect 2342 823 2348 824
rect 2342 822 2343 823
rect 1722 818 1728 819
rect 1940 820 2343 822
rect 1940 818 1942 820
rect 2342 819 2343 820
rect 2347 819 2348 823
rect 2342 818 2348 819
rect 1443 817 1449 818
rect 238 813 244 814
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 238 809 239 813
rect 243 809 244 813
rect 238 808 244 809
rect 259 813 286 814
rect 259 809 260 813
rect 264 812 286 813
rect 302 813 308 814
rect 264 809 265 812
rect 259 808 265 809
rect 302 809 303 813
rect 307 809 308 813
rect 382 813 388 814
rect 302 808 308 809
rect 323 811 329 812
rect 110 807 116 808
rect 323 807 324 811
rect 328 810 329 811
rect 350 811 356 812
rect 350 810 351 811
rect 328 808 351 810
rect 328 807 329 808
rect 323 806 329 807
rect 350 807 351 808
rect 355 807 356 811
rect 382 809 383 813
rect 387 809 388 813
rect 462 813 468 814
rect 382 808 388 809
rect 402 811 409 812
rect 350 806 356 807
rect 402 807 403 811
rect 408 807 409 811
rect 462 809 463 813
rect 467 809 468 813
rect 462 808 468 809
rect 483 813 489 814
rect 483 809 484 813
rect 488 809 489 813
rect 483 808 489 809
rect 550 813 556 814
rect 550 809 551 813
rect 555 809 556 813
rect 550 808 556 809
rect 571 813 577 814
rect 571 809 572 813
rect 576 809 577 813
rect 571 808 577 809
rect 638 813 644 814
rect 638 809 639 813
rect 643 809 644 813
rect 638 808 644 809
rect 659 813 665 814
rect 659 809 660 813
rect 664 809 665 813
rect 659 808 665 809
rect 726 813 732 814
rect 726 809 727 813
rect 731 809 732 813
rect 726 808 732 809
rect 747 813 753 814
rect 747 809 748 813
rect 752 809 753 813
rect 747 808 753 809
rect 806 813 812 814
rect 806 809 807 813
rect 811 809 812 813
rect 806 808 812 809
rect 827 813 833 814
rect 827 809 828 813
rect 832 809 833 813
rect 827 808 833 809
rect 894 813 900 814
rect 894 809 895 813
rect 899 809 900 813
rect 894 808 900 809
rect 915 813 921 814
rect 915 809 916 813
rect 920 809 921 813
rect 915 808 921 809
rect 982 813 988 814
rect 982 809 983 813
rect 987 809 988 813
rect 982 808 988 809
rect 1003 813 1009 814
rect 1003 809 1004 813
rect 1008 809 1009 813
rect 1003 808 1009 809
rect 1070 813 1076 814
rect 1443 813 1444 817
rect 1448 813 1449 817
rect 1675 817 1681 818
rect 1515 815 1521 816
rect 1515 814 1516 815
rect 1070 809 1071 813
rect 1075 809 1076 813
rect 1286 812 1292 813
rect 1443 812 1449 813
rect 1461 812 1516 814
rect 1070 808 1076 809
rect 1090 811 1097 812
rect 402 806 409 807
rect 1090 807 1091 811
rect 1096 807 1097 811
rect 1286 808 1287 812
rect 1291 808 1292 812
rect 1286 807 1292 808
rect 1090 806 1097 807
rect 1461 802 1463 812
rect 1515 811 1516 812
rect 1520 811 1521 815
rect 1595 815 1601 816
rect 1595 814 1596 815
rect 1515 810 1521 811
rect 1532 812 1596 814
rect 1532 802 1534 812
rect 1595 811 1596 812
rect 1600 811 1601 815
rect 1675 813 1676 817
rect 1680 813 1681 817
rect 1939 817 1945 818
rect 1763 815 1769 816
rect 1763 814 1764 815
rect 1675 812 1681 813
rect 1692 812 1764 814
rect 1595 810 1601 811
rect 1692 802 1694 812
rect 1763 811 1764 812
rect 1768 811 1769 815
rect 1851 815 1857 816
rect 1851 814 1852 815
rect 1763 810 1769 811
rect 1780 812 1852 814
rect 1780 802 1782 812
rect 1851 811 1852 812
rect 1856 811 1857 815
rect 1939 813 1940 817
rect 1944 813 1945 817
rect 2027 815 2033 816
rect 2027 814 2028 815
rect 1939 812 1945 813
rect 1999 812 2028 814
rect 1851 810 1857 811
rect 1818 807 1824 808
rect 1818 803 1819 807
rect 1823 806 1824 807
rect 1999 806 2001 812
rect 2027 811 2028 812
rect 2032 811 2033 815
rect 2115 815 2121 816
rect 2115 814 2116 815
rect 2027 810 2033 811
rect 2044 812 2116 814
rect 1823 804 1870 806
rect 1823 803 1824 804
rect 1818 802 1824 803
rect 1868 802 1870 804
rect 1956 804 2001 806
rect 1956 802 1958 804
rect 2044 802 2046 812
rect 2115 811 2116 812
rect 2120 811 2121 815
rect 2203 815 2209 816
rect 2203 814 2204 815
rect 2115 810 2121 811
rect 2132 812 2204 814
rect 2132 802 2134 812
rect 2203 811 2204 812
rect 2208 811 2209 815
rect 2203 810 2209 811
rect 2291 815 2297 816
rect 2291 811 2292 815
rect 2296 811 2297 815
rect 2291 810 2297 811
rect 2387 815 2396 816
rect 2387 811 2388 815
rect 2395 811 2396 815
rect 2387 810 2396 811
rect 2459 815 2468 816
rect 2459 811 2460 815
rect 2467 811 2468 815
rect 2459 810 2468 811
rect 2293 806 2295 810
rect 2220 804 2295 806
rect 2220 802 2222 804
rect 1438 801 1444 802
rect 1326 800 1332 801
rect 1326 796 1327 800
rect 1331 796 1332 800
rect 1438 797 1439 801
rect 1443 797 1444 801
rect 1438 796 1444 797
rect 1459 801 1465 802
rect 1459 797 1460 801
rect 1464 797 1465 801
rect 1459 796 1465 797
rect 1510 801 1516 802
rect 1510 797 1511 801
rect 1515 797 1516 801
rect 1510 796 1516 797
rect 1531 801 1537 802
rect 1531 797 1532 801
rect 1536 797 1537 801
rect 1531 796 1537 797
rect 1590 801 1596 802
rect 1590 797 1591 801
rect 1595 797 1596 801
rect 1670 801 1676 802
rect 1590 796 1596 797
rect 1598 799 1604 800
rect 110 795 116 796
rect 110 791 111 795
rect 115 791 116 795
rect 1286 795 1292 796
rect 1326 795 1332 796
rect 1598 795 1599 799
rect 1603 798 1604 799
rect 1611 799 1617 800
rect 1611 798 1612 799
rect 1603 796 1612 798
rect 1603 795 1604 796
rect 110 790 116 791
rect 222 792 228 793
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 286 792 292 793
rect 286 788 287 792
rect 291 788 292 792
rect 286 787 292 788
rect 366 792 372 793
rect 366 788 367 792
rect 371 788 372 792
rect 366 787 372 788
rect 446 792 452 793
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 534 792 540 793
rect 534 788 535 792
rect 539 788 540 792
rect 534 787 540 788
rect 622 792 628 793
rect 622 788 623 792
rect 627 788 628 792
rect 622 787 628 788
rect 710 792 716 793
rect 710 788 711 792
rect 715 788 716 792
rect 710 787 716 788
rect 790 792 796 793
rect 790 788 791 792
rect 795 788 796 792
rect 790 787 796 788
rect 878 792 884 793
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 966 792 972 793
rect 966 788 967 792
rect 971 788 972 792
rect 966 787 972 788
rect 1054 792 1060 793
rect 1054 788 1055 792
rect 1059 788 1060 792
rect 1286 791 1287 795
rect 1291 791 1292 795
rect 1598 794 1604 795
rect 1611 795 1612 796
rect 1616 795 1617 799
rect 1670 797 1671 801
rect 1675 797 1676 801
rect 1670 796 1676 797
rect 1691 801 1697 802
rect 1691 797 1692 801
rect 1696 797 1697 801
rect 1691 796 1697 797
rect 1758 801 1764 802
rect 1758 797 1759 801
rect 1763 797 1764 801
rect 1758 796 1764 797
rect 1779 801 1785 802
rect 1779 797 1780 801
rect 1784 797 1785 801
rect 1779 796 1785 797
rect 1846 801 1852 802
rect 1846 797 1847 801
rect 1851 797 1852 801
rect 1846 796 1852 797
rect 1867 801 1873 802
rect 1867 797 1868 801
rect 1872 797 1873 801
rect 1867 796 1873 797
rect 1934 801 1940 802
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 1955 801 1961 802
rect 1955 797 1956 801
rect 1960 797 1961 801
rect 1955 796 1961 797
rect 2022 801 2028 802
rect 2022 797 2023 801
rect 2027 797 2028 801
rect 2022 796 2028 797
rect 2043 801 2049 802
rect 2043 797 2044 801
rect 2048 797 2049 801
rect 2043 796 2049 797
rect 2110 801 2116 802
rect 2110 797 2111 801
rect 2115 797 2116 801
rect 2110 796 2116 797
rect 2131 801 2137 802
rect 2131 797 2132 801
rect 2136 797 2137 801
rect 2131 796 2137 797
rect 2198 801 2204 802
rect 2198 797 2199 801
rect 2203 797 2204 801
rect 2198 796 2204 797
rect 2219 801 2225 802
rect 2219 797 2220 801
rect 2224 797 2225 801
rect 2219 796 2225 797
rect 2286 801 2292 802
rect 2286 797 2287 801
rect 2291 797 2292 801
rect 2382 801 2388 802
rect 2286 796 2292 797
rect 2294 799 2300 800
rect 1611 794 1617 795
rect 2294 795 2295 799
rect 2299 798 2300 799
rect 2307 799 2313 800
rect 2307 798 2308 799
rect 2299 796 2308 798
rect 2299 795 2300 796
rect 2294 794 2300 795
rect 2307 795 2308 796
rect 2312 795 2313 799
rect 2382 797 2383 801
rect 2387 797 2388 801
rect 2454 801 2460 802
rect 2382 796 2388 797
rect 2403 799 2412 800
rect 2307 794 2313 795
rect 2403 795 2404 799
rect 2411 795 2412 799
rect 2454 797 2455 801
rect 2459 797 2460 801
rect 2502 800 2508 801
rect 2454 796 2460 797
rect 2470 799 2481 800
rect 2403 794 2412 795
rect 2470 795 2471 799
rect 2475 795 2476 799
rect 2480 795 2481 799
rect 2502 796 2503 800
rect 2507 796 2508 800
rect 2502 795 2508 796
rect 2470 794 2481 795
rect 1286 790 1292 791
rect 1054 787 1060 788
rect 762 783 768 784
rect 762 779 763 783
rect 767 782 768 783
rect 1010 783 1016 784
rect 1010 782 1011 783
rect 767 780 1011 782
rect 767 779 768 780
rect 762 778 768 779
rect 1010 779 1011 780
rect 1015 779 1016 783
rect 1010 778 1016 779
rect 1326 783 1332 784
rect 1326 779 1327 783
rect 1331 779 1332 783
rect 2502 783 2508 784
rect 1326 778 1332 779
rect 1422 780 1428 781
rect 150 776 156 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 150 772 151 776
rect 155 772 156 776
rect 150 771 156 772
rect 246 776 252 777
rect 246 772 247 776
rect 251 772 252 776
rect 246 771 252 772
rect 342 776 348 777
rect 342 772 343 776
rect 347 772 348 776
rect 342 771 348 772
rect 438 776 444 777
rect 438 772 439 776
rect 443 772 444 776
rect 438 771 444 772
rect 526 776 532 777
rect 526 772 527 776
rect 531 772 532 776
rect 526 771 532 772
rect 606 776 612 777
rect 606 772 607 776
rect 611 772 612 776
rect 606 771 612 772
rect 678 776 684 777
rect 678 772 679 776
rect 683 772 684 776
rect 678 771 684 772
rect 750 776 756 777
rect 750 772 751 776
rect 755 772 756 776
rect 750 771 756 772
rect 822 776 828 777
rect 822 772 823 776
rect 827 772 828 776
rect 822 771 828 772
rect 894 776 900 777
rect 894 772 895 776
rect 899 772 900 776
rect 894 771 900 772
rect 974 776 980 777
rect 974 772 975 776
rect 979 772 980 776
rect 1422 776 1423 780
rect 1427 776 1428 780
rect 1422 775 1428 776
rect 1494 780 1500 781
rect 1494 776 1495 780
rect 1499 776 1500 780
rect 1494 775 1500 776
rect 1574 780 1580 781
rect 1574 776 1575 780
rect 1579 776 1580 780
rect 1574 775 1580 776
rect 1654 780 1660 781
rect 1654 776 1655 780
rect 1659 776 1660 780
rect 1654 775 1660 776
rect 1742 780 1748 781
rect 1742 776 1743 780
rect 1747 776 1748 780
rect 1742 775 1748 776
rect 1830 780 1836 781
rect 1830 776 1831 780
rect 1835 776 1836 780
rect 1830 775 1836 776
rect 1918 780 1924 781
rect 1918 776 1919 780
rect 1923 776 1924 780
rect 1918 775 1924 776
rect 2006 780 2012 781
rect 2006 776 2007 780
rect 2011 776 2012 780
rect 2006 775 2012 776
rect 2094 780 2100 781
rect 2094 776 2095 780
rect 2099 776 2100 780
rect 2094 775 2100 776
rect 2182 780 2188 781
rect 2182 776 2183 780
rect 2187 776 2188 780
rect 2182 775 2188 776
rect 2270 780 2276 781
rect 2270 776 2271 780
rect 2275 776 2276 780
rect 2270 775 2276 776
rect 2366 780 2372 781
rect 2366 776 2367 780
rect 2371 776 2372 780
rect 2366 775 2372 776
rect 2438 780 2444 781
rect 2438 776 2439 780
rect 2443 776 2444 780
rect 2502 779 2503 783
rect 2507 779 2508 783
rect 2502 778 2508 779
rect 2438 775 2444 776
rect 974 771 980 772
rect 1286 773 1292 774
rect 110 768 116 769
rect 1286 769 1287 773
rect 1291 769 1292 773
rect 1286 768 1292 769
rect 1350 764 1356 765
rect 1326 761 1332 762
rect 1326 757 1327 761
rect 1331 757 1332 761
rect 1350 760 1351 764
rect 1355 760 1356 764
rect 1350 759 1356 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1566 764 1572 765
rect 1566 760 1567 764
rect 1571 760 1572 764
rect 1566 759 1572 760
rect 1686 764 1692 765
rect 1686 760 1687 764
rect 1691 760 1692 764
rect 1686 759 1692 760
rect 1806 764 1812 765
rect 1806 760 1807 764
rect 1811 760 1812 764
rect 1806 759 1812 760
rect 1926 764 1932 765
rect 1926 760 1927 764
rect 1931 760 1932 764
rect 1926 759 1932 760
rect 2038 764 2044 765
rect 2038 760 2039 764
rect 2043 760 2044 764
rect 2038 759 2044 760
rect 2142 764 2148 765
rect 2142 760 2143 764
rect 2147 760 2148 764
rect 2142 759 2148 760
rect 2246 764 2252 765
rect 2246 760 2247 764
rect 2251 760 2252 764
rect 2246 759 2252 760
rect 2350 764 2356 765
rect 2350 760 2351 764
rect 2355 760 2356 764
rect 2350 759 2356 760
rect 2438 764 2444 765
rect 2438 760 2439 764
rect 2443 760 2444 764
rect 2438 759 2444 760
rect 2502 761 2508 762
rect 110 756 116 757
rect 1286 756 1292 757
rect 1326 756 1332 757
rect 2502 757 2503 761
rect 2507 757 2508 761
rect 2502 756 2508 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 166 750 172 751
rect 182 755 193 756
rect 182 751 183 755
rect 187 751 188 755
rect 192 751 193 755
rect 182 750 193 751
rect 262 755 268 756
rect 262 751 263 755
rect 267 751 268 755
rect 262 750 268 751
rect 278 755 289 756
rect 278 751 279 755
rect 283 751 284 755
rect 288 751 289 755
rect 278 750 289 751
rect 358 755 364 756
rect 358 751 359 755
rect 363 751 364 755
rect 379 755 385 756
rect 379 754 380 755
rect 358 750 364 751
rect 368 752 380 754
rect 368 746 370 752
rect 379 751 380 752
rect 384 751 385 755
rect 379 750 385 751
rect 454 755 460 756
rect 454 751 455 755
rect 459 751 460 755
rect 454 750 460 751
rect 475 755 481 756
rect 475 751 476 755
rect 480 754 481 755
rect 542 755 548 756
rect 480 752 534 754
rect 480 751 481 752
rect 475 750 481 751
rect 268 744 370 746
rect 268 742 270 744
rect 532 742 534 752
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 563 755 572 756
rect 563 751 564 755
rect 571 751 572 755
rect 563 750 572 751
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 643 755 649 756
rect 643 751 644 755
rect 648 754 649 755
rect 694 755 700 756
rect 648 752 690 754
rect 648 751 649 752
rect 643 750 649 751
rect 688 742 690 752
rect 694 751 695 755
rect 699 751 700 755
rect 694 750 700 751
rect 715 755 721 756
rect 715 751 716 755
rect 720 754 721 755
rect 766 755 772 756
rect 720 752 762 754
rect 720 751 721 752
rect 715 750 721 751
rect 760 742 762 752
rect 766 751 767 755
rect 771 751 772 755
rect 766 750 772 751
rect 787 755 793 756
rect 787 751 788 755
rect 792 754 793 755
rect 838 755 844 756
rect 792 752 830 754
rect 792 751 793 752
rect 787 750 793 751
rect 828 742 830 752
rect 838 751 839 755
rect 843 751 844 755
rect 838 750 844 751
rect 859 755 865 756
rect 859 751 860 755
rect 864 754 865 755
rect 910 755 916 756
rect 864 752 906 754
rect 864 751 865 752
rect 859 750 865 751
rect 904 742 906 752
rect 910 751 911 755
rect 915 751 916 755
rect 910 750 916 751
rect 931 755 937 756
rect 931 751 932 755
rect 936 754 937 755
rect 990 755 996 756
rect 936 752 978 754
rect 936 751 937 752
rect 931 750 937 751
rect 976 742 978 752
rect 990 751 991 755
rect 995 751 996 755
rect 990 750 996 751
rect 1010 755 1017 756
rect 1010 751 1011 755
rect 1016 751 1017 755
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1010 750 1017 751
rect 1326 744 1332 745
rect 2502 744 2508 745
rect 267 741 273 742
rect 171 739 177 740
rect 171 735 172 739
rect 176 735 177 739
rect 267 737 268 741
rect 272 737 273 741
rect 532 741 553 742
rect 532 740 548 741
rect 267 736 273 737
rect 350 739 356 740
rect 171 734 177 735
rect 278 735 284 736
rect 278 734 279 735
rect 173 732 279 734
rect 278 731 279 732
rect 283 731 284 735
rect 350 735 351 739
rect 355 738 356 739
rect 363 739 369 740
rect 363 738 364 739
rect 355 736 364 738
rect 355 735 356 736
rect 350 734 356 735
rect 363 735 364 736
rect 368 735 369 739
rect 363 734 369 735
rect 374 739 380 740
rect 374 735 375 739
rect 379 738 380 739
rect 459 739 465 740
rect 459 738 460 739
rect 379 736 460 738
rect 379 735 380 736
rect 374 734 380 735
rect 459 735 460 736
rect 464 735 465 739
rect 547 737 548 740
rect 552 737 553 741
rect 688 741 705 742
rect 688 740 700 741
rect 547 736 553 737
rect 627 739 633 740
rect 459 734 465 735
rect 627 735 628 739
rect 632 738 633 739
rect 632 736 694 738
rect 699 737 700 740
rect 704 737 705 741
rect 760 741 777 742
rect 760 740 772 741
rect 699 736 705 737
rect 771 737 772 740
rect 776 737 777 741
rect 828 741 849 742
rect 828 740 844 741
rect 771 736 777 737
rect 843 737 844 740
rect 848 737 849 741
rect 904 741 921 742
rect 904 740 916 741
rect 843 736 849 737
rect 915 737 916 740
rect 920 737 921 741
rect 976 741 1001 742
rect 976 740 996 741
rect 915 736 921 737
rect 995 737 996 740
rect 1000 737 1001 741
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 1326 739 1332 740
rect 1366 743 1372 744
rect 1366 739 1367 743
rect 1371 739 1372 743
rect 1366 738 1372 739
rect 1374 743 1380 744
rect 1374 739 1375 743
rect 1379 742 1380 743
rect 1387 743 1393 744
rect 1387 742 1388 743
rect 1379 740 1388 742
rect 1379 739 1380 740
rect 1374 738 1380 739
rect 1387 739 1388 740
rect 1392 739 1393 743
rect 1387 738 1393 739
rect 1462 743 1468 744
rect 1462 739 1463 743
rect 1467 739 1468 743
rect 1462 738 1468 739
rect 1483 743 1489 744
rect 1483 739 1484 743
rect 1488 739 1489 743
rect 1483 738 1489 739
rect 1582 743 1588 744
rect 1582 739 1583 743
rect 1587 739 1588 743
rect 1603 743 1609 744
rect 1603 742 1604 743
rect 1582 738 1588 739
rect 1592 740 1604 742
rect 995 736 1001 737
rect 632 735 633 736
rect 627 734 633 735
rect 692 734 694 736
rect 930 735 936 736
rect 930 734 931 735
rect 692 732 931 734
rect 278 730 284 731
rect 930 731 931 732
rect 935 731 936 735
rect 1485 734 1487 738
rect 1592 734 1594 740
rect 1603 739 1604 740
rect 1608 739 1609 743
rect 1603 738 1609 739
rect 1702 743 1708 744
rect 1702 739 1703 743
rect 1707 739 1708 743
rect 1702 738 1708 739
rect 1722 743 1729 744
rect 1722 739 1723 743
rect 1728 739 1729 743
rect 1722 738 1729 739
rect 1822 743 1828 744
rect 1822 739 1823 743
rect 1827 739 1828 743
rect 1822 738 1828 739
rect 1843 743 1849 744
rect 1843 739 1844 743
rect 1848 739 1849 743
rect 1843 738 1849 739
rect 1942 743 1948 744
rect 1942 739 1943 743
rect 1947 739 1948 743
rect 1942 738 1948 739
rect 1963 743 1969 744
rect 1963 739 1964 743
rect 1968 742 1969 743
rect 2054 743 2060 744
rect 1968 740 2001 742
rect 1968 739 1969 740
rect 1963 738 1969 739
rect 1845 734 1847 738
rect 930 730 936 731
rect 1372 732 1487 734
rect 1492 732 1594 734
rect 1708 732 1847 734
rect 1372 730 1374 732
rect 1492 730 1494 732
rect 1708 730 1710 732
rect 1999 730 2001 740
rect 2054 739 2055 743
rect 2059 739 2060 743
rect 2054 738 2060 739
rect 2075 743 2081 744
rect 2075 739 2076 743
rect 2080 742 2081 743
rect 2158 743 2164 744
rect 2080 740 2134 742
rect 2080 739 2081 740
rect 2075 738 2081 739
rect 2132 730 2134 740
rect 2158 739 2159 743
rect 2163 739 2164 743
rect 2158 738 2164 739
rect 2179 743 2185 744
rect 2179 739 2180 743
rect 2184 742 2185 743
rect 2262 743 2268 744
rect 2184 740 2254 742
rect 2184 739 2185 740
rect 2179 738 2185 739
rect 2252 730 2254 740
rect 2262 739 2263 743
rect 2267 739 2268 743
rect 2262 738 2268 739
rect 2270 743 2276 744
rect 2270 739 2271 743
rect 2275 742 2276 743
rect 2283 743 2289 744
rect 2283 742 2284 743
rect 2275 740 2284 742
rect 2275 739 2276 740
rect 2270 738 2276 739
rect 2283 739 2284 740
rect 2288 739 2289 743
rect 2283 738 2289 739
rect 2366 743 2372 744
rect 2366 739 2367 743
rect 2371 739 2372 743
rect 2366 738 2372 739
rect 2387 743 2396 744
rect 2387 739 2388 743
rect 2395 739 2396 743
rect 2387 738 2396 739
rect 2454 743 2460 744
rect 2454 739 2455 743
rect 2459 739 2460 743
rect 2454 738 2460 739
rect 2462 743 2468 744
rect 2462 739 2463 743
rect 2467 742 2468 743
rect 2475 743 2481 744
rect 2475 742 2476 743
rect 2467 740 2476 742
rect 2467 739 2468 740
rect 2462 738 2468 739
rect 2475 739 2476 740
rect 2480 739 2481 743
rect 2502 740 2503 744
rect 2507 740 2508 744
rect 2502 739 2508 740
rect 2475 738 2481 739
rect 1371 729 1377 730
rect 1371 725 1372 729
rect 1376 725 1377 729
rect 1371 724 1377 725
rect 1467 729 1494 730
rect 1467 725 1468 729
rect 1472 728 1494 729
rect 1707 729 1713 730
rect 1472 725 1473 728
rect 1467 724 1473 725
rect 1587 727 1593 728
rect 594 723 600 724
rect 594 722 595 723
rect 428 720 595 722
rect 428 718 430 720
rect 594 719 595 720
rect 599 719 600 723
rect 1587 723 1588 727
rect 1592 726 1593 727
rect 1598 727 1604 728
rect 1598 726 1599 727
rect 1592 724 1599 726
rect 1592 723 1593 724
rect 1587 722 1593 723
rect 1598 723 1599 724
rect 1603 723 1604 727
rect 1707 725 1708 729
rect 1712 725 1713 729
rect 1999 729 2065 730
rect 1999 728 2060 729
rect 1707 724 1713 725
rect 1827 727 1833 728
rect 1598 722 1604 723
rect 1827 723 1828 727
rect 1832 726 1833 727
rect 1882 727 1888 728
rect 1882 726 1883 727
rect 1832 724 1883 726
rect 1832 723 1833 724
rect 1827 722 1833 723
rect 1882 723 1883 724
rect 1887 723 1888 727
rect 1882 722 1888 723
rect 1947 727 1953 728
rect 1947 723 1948 727
rect 1952 726 1953 727
rect 1952 724 2001 726
rect 2059 725 2060 728
rect 2064 725 2065 729
rect 2132 729 2169 730
rect 2132 728 2164 729
rect 2059 724 2065 725
rect 2163 725 2164 728
rect 2168 725 2169 729
rect 2252 729 2273 730
rect 2252 728 2268 729
rect 2163 724 2169 725
rect 2267 725 2268 728
rect 2272 725 2273 729
rect 2267 724 2273 725
rect 2371 727 2377 728
rect 1952 723 1953 724
rect 1947 722 1953 723
rect 1999 722 2001 724
rect 2294 723 2300 724
rect 2294 722 2295 723
rect 1999 720 2295 722
rect 594 718 600 719
rect 2294 719 2295 720
rect 2299 719 2300 723
rect 2371 723 2372 727
rect 2376 726 2377 727
rect 2410 727 2416 728
rect 2410 726 2411 727
rect 2376 724 2411 726
rect 2376 723 2377 724
rect 2371 722 2377 723
rect 2410 723 2411 724
rect 2415 723 2416 727
rect 2410 722 2416 723
rect 2459 727 2465 728
rect 2459 723 2460 727
rect 2464 726 2465 727
rect 2470 727 2476 728
rect 2470 726 2471 727
rect 2464 724 2471 726
rect 2464 723 2465 724
rect 2459 722 2465 723
rect 2470 723 2471 724
rect 2475 723 2476 727
rect 2470 722 2476 723
rect 2294 718 2300 719
rect 427 717 433 718
rect 179 715 188 716
rect 179 711 180 715
rect 187 711 188 715
rect 179 710 188 711
rect 267 715 273 716
rect 267 711 268 715
rect 272 714 273 715
rect 310 715 316 716
rect 310 714 311 715
rect 272 712 311 714
rect 272 711 273 712
rect 267 710 273 711
rect 310 711 311 712
rect 315 711 316 715
rect 347 715 353 716
rect 347 714 348 715
rect 310 710 316 711
rect 319 712 348 714
rect 319 706 321 712
rect 347 711 348 712
rect 352 711 353 715
rect 427 713 428 717
rect 432 713 433 717
rect 507 715 513 716
rect 507 714 508 715
rect 427 712 433 713
rect 445 712 508 714
rect 347 710 353 711
rect 284 704 321 706
rect 284 702 286 704
rect 445 702 447 712
rect 507 711 508 712
rect 512 711 513 715
rect 507 710 513 711
rect 566 715 572 716
rect 566 711 567 715
rect 571 714 572 715
rect 579 715 585 716
rect 579 714 580 715
rect 571 712 580 714
rect 571 711 572 712
rect 566 710 572 711
rect 579 711 580 712
rect 584 711 585 715
rect 579 710 585 711
rect 630 715 636 716
rect 630 711 631 715
rect 635 714 636 715
rect 643 715 649 716
rect 643 714 644 715
rect 635 712 644 714
rect 635 711 636 712
rect 630 710 636 711
rect 643 711 644 712
rect 648 711 649 715
rect 707 715 713 716
rect 707 714 708 715
rect 643 710 649 711
rect 684 712 708 714
rect 684 706 686 712
rect 707 711 708 712
rect 712 711 713 715
rect 771 715 777 716
rect 771 714 772 715
rect 707 710 713 711
rect 724 712 772 714
rect 660 704 686 706
rect 660 702 662 704
rect 724 702 726 712
rect 771 711 772 712
rect 776 711 777 715
rect 843 715 849 716
rect 843 714 844 715
rect 771 710 777 711
rect 800 712 844 714
rect 800 706 802 712
rect 843 711 844 712
rect 848 711 849 715
rect 915 715 921 716
rect 915 714 916 715
rect 843 710 849 711
rect 860 712 916 714
rect 788 704 802 706
rect 788 702 790 704
rect 860 702 862 712
rect 915 711 916 712
rect 920 711 921 715
rect 915 710 921 711
rect 1371 703 1380 704
rect 174 701 180 702
rect 110 700 116 701
rect 110 696 111 700
rect 115 696 116 700
rect 174 697 175 701
rect 179 697 180 701
rect 262 701 268 702
rect 174 696 180 697
rect 195 699 201 700
rect 110 695 116 696
rect 195 695 196 699
rect 200 698 201 699
rect 222 699 228 700
rect 222 698 223 699
rect 200 696 223 698
rect 200 695 201 696
rect 195 694 201 695
rect 222 695 223 696
rect 227 695 228 699
rect 262 697 263 701
rect 267 697 268 701
rect 262 696 268 697
rect 283 701 289 702
rect 283 697 284 701
rect 288 697 289 701
rect 283 696 289 697
rect 342 701 348 702
rect 342 697 343 701
rect 347 697 348 701
rect 422 701 428 702
rect 342 696 348 697
rect 363 699 369 700
rect 222 694 228 695
rect 363 695 364 699
rect 368 698 369 699
rect 374 699 380 700
rect 374 698 375 699
rect 368 696 375 698
rect 368 695 369 696
rect 363 694 369 695
rect 374 695 375 696
rect 379 695 380 699
rect 422 697 423 701
rect 427 697 428 701
rect 422 696 428 697
rect 443 701 449 702
rect 443 697 444 701
rect 448 697 449 701
rect 443 696 449 697
rect 502 701 508 702
rect 502 697 503 701
rect 507 697 508 701
rect 574 701 580 702
rect 502 696 508 697
rect 523 699 529 700
rect 374 694 380 695
rect 523 695 524 699
rect 528 698 529 699
rect 534 699 540 700
rect 534 698 535 699
rect 528 696 535 698
rect 528 695 529 696
rect 523 694 529 695
rect 534 695 535 696
rect 539 695 540 699
rect 574 697 575 701
rect 579 697 580 701
rect 638 701 644 702
rect 574 696 580 697
rect 594 699 601 700
rect 534 694 540 695
rect 594 695 595 699
rect 600 695 601 699
rect 638 697 639 701
rect 643 697 644 701
rect 638 696 644 697
rect 659 701 665 702
rect 659 697 660 701
rect 664 697 665 701
rect 659 696 665 697
rect 702 701 708 702
rect 702 697 703 701
rect 707 697 708 701
rect 702 696 708 697
rect 723 701 729 702
rect 723 697 724 701
rect 728 697 729 701
rect 723 696 729 697
rect 766 701 772 702
rect 766 697 767 701
rect 771 697 772 701
rect 766 696 772 697
rect 787 701 793 702
rect 787 697 788 701
rect 792 697 793 701
rect 787 696 793 697
rect 838 701 844 702
rect 838 697 839 701
rect 843 697 844 701
rect 838 696 844 697
rect 859 701 865 702
rect 859 697 860 701
rect 864 697 865 701
rect 859 696 865 697
rect 910 701 916 702
rect 910 697 911 701
rect 915 697 916 701
rect 1286 700 1292 701
rect 910 696 916 697
rect 930 699 937 700
rect 594 694 601 695
rect 930 695 931 699
rect 936 695 937 699
rect 1286 696 1287 700
rect 1291 696 1292 700
rect 1371 699 1372 703
rect 1379 699 1380 703
rect 1435 703 1441 704
rect 1435 702 1436 703
rect 1371 698 1380 699
rect 1389 700 1436 702
rect 1286 695 1292 696
rect 930 694 937 695
rect 1389 690 1391 700
rect 1435 699 1436 700
rect 1440 699 1441 703
rect 1539 703 1545 704
rect 1539 702 1540 703
rect 1435 698 1441 699
rect 1452 700 1540 702
rect 1452 690 1454 700
rect 1539 699 1540 700
rect 1544 699 1545 703
rect 1643 703 1649 704
rect 1643 702 1644 703
rect 1539 698 1545 699
rect 1557 700 1644 702
rect 1557 690 1559 700
rect 1643 699 1644 700
rect 1648 699 1649 703
rect 1643 698 1649 699
rect 1755 703 1764 704
rect 1755 699 1756 703
rect 1763 699 1764 703
rect 1867 703 1873 704
rect 1867 702 1868 703
rect 1755 698 1764 699
rect 1772 700 1868 702
rect 1772 690 1774 700
rect 1867 699 1868 700
rect 1872 699 1873 703
rect 1867 698 1873 699
rect 1971 703 1980 704
rect 1971 699 1972 703
rect 1979 699 1980 703
rect 2067 703 2073 704
rect 2067 702 2068 703
rect 1971 698 1980 699
rect 1999 700 2068 702
rect 1999 694 2001 700
rect 2067 699 2068 700
rect 2072 699 2073 703
rect 2155 703 2161 704
rect 2155 702 2156 703
rect 2067 698 2073 699
rect 2084 700 2156 702
rect 1988 692 2001 694
rect 1988 690 1990 692
rect 2084 690 2086 700
rect 2155 699 2156 700
rect 2160 699 2161 703
rect 2155 698 2161 699
rect 2235 703 2241 704
rect 2235 699 2236 703
rect 2240 702 2241 703
rect 2274 703 2280 704
rect 2274 702 2275 703
rect 2240 700 2275 702
rect 2240 699 2241 700
rect 2235 698 2241 699
rect 2274 699 2275 700
rect 2279 699 2280 703
rect 2315 703 2321 704
rect 2315 702 2316 703
rect 2274 698 2280 699
rect 2284 700 2316 702
rect 2284 694 2286 700
rect 2315 699 2316 700
rect 2320 699 2321 703
rect 2315 698 2321 699
rect 2395 703 2401 704
rect 2395 699 2396 703
rect 2400 699 2401 703
rect 2395 698 2401 699
rect 2459 703 2468 704
rect 2459 699 2460 703
rect 2467 699 2468 703
rect 2459 698 2468 699
rect 2397 694 2399 698
rect 2172 692 2286 694
rect 2332 692 2399 694
rect 2172 690 2174 692
rect 2332 690 2334 692
rect 1366 689 1372 690
rect 1326 688 1332 689
rect 1326 684 1327 688
rect 1331 684 1332 688
rect 1366 685 1367 689
rect 1371 685 1372 689
rect 1366 684 1372 685
rect 1387 689 1393 690
rect 1387 685 1388 689
rect 1392 685 1393 689
rect 1387 684 1393 685
rect 1430 689 1436 690
rect 1430 685 1431 689
rect 1435 685 1436 689
rect 1430 684 1436 685
rect 1451 689 1457 690
rect 1451 685 1452 689
rect 1456 685 1457 689
rect 1451 684 1457 685
rect 1534 689 1540 690
rect 1534 685 1535 689
rect 1539 685 1540 689
rect 1534 684 1540 685
rect 1555 689 1561 690
rect 1555 685 1556 689
rect 1560 685 1561 689
rect 1555 684 1561 685
rect 1638 689 1644 690
rect 1638 685 1639 689
rect 1643 685 1644 689
rect 1750 689 1756 690
rect 1638 684 1644 685
rect 1654 687 1665 688
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 1286 683 1292 684
rect 1326 683 1332 684
rect 1654 683 1655 687
rect 1659 683 1660 687
rect 1664 683 1665 687
rect 1750 685 1751 689
rect 1755 685 1756 689
rect 1750 684 1756 685
rect 1771 689 1777 690
rect 1771 685 1772 689
rect 1776 685 1777 689
rect 1771 684 1777 685
rect 1862 689 1868 690
rect 1862 685 1863 689
rect 1867 685 1868 689
rect 1966 689 1972 690
rect 1862 684 1868 685
rect 1882 687 1889 688
rect 110 678 116 679
rect 158 680 164 681
rect 158 676 159 680
rect 163 676 164 680
rect 158 675 164 676
rect 246 680 252 681
rect 246 676 247 680
rect 251 676 252 680
rect 246 675 252 676
rect 326 680 332 681
rect 326 676 327 680
rect 331 676 332 680
rect 326 675 332 676
rect 406 680 412 681
rect 406 676 407 680
rect 411 676 412 680
rect 406 675 412 676
rect 486 680 492 681
rect 486 676 487 680
rect 491 676 492 680
rect 486 675 492 676
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 686 680 692 681
rect 686 676 687 680
rect 691 676 692 680
rect 686 675 692 676
rect 750 680 756 681
rect 750 676 751 680
rect 755 676 756 680
rect 750 675 756 676
rect 822 680 828 681
rect 822 676 823 680
rect 827 676 828 680
rect 822 675 828 676
rect 894 680 900 681
rect 894 676 895 680
rect 899 676 900 680
rect 1286 679 1287 683
rect 1291 679 1292 683
rect 1654 682 1665 683
rect 1882 683 1883 687
rect 1888 683 1889 687
rect 1966 685 1967 689
rect 1971 685 1972 689
rect 1966 684 1972 685
rect 1987 689 1993 690
rect 1987 685 1988 689
rect 1992 685 1993 689
rect 1987 684 1993 685
rect 2062 689 2068 690
rect 2062 685 2063 689
rect 2067 685 2068 689
rect 2062 684 2068 685
rect 2083 689 2089 690
rect 2083 685 2084 689
rect 2088 685 2089 689
rect 2083 684 2089 685
rect 2150 689 2156 690
rect 2150 685 2151 689
rect 2155 685 2156 689
rect 2150 684 2156 685
rect 2171 689 2177 690
rect 2171 685 2172 689
rect 2176 685 2177 689
rect 2171 684 2177 685
rect 2230 689 2236 690
rect 2230 685 2231 689
rect 2235 685 2236 689
rect 2310 689 2316 690
rect 2230 684 2236 685
rect 2246 687 2257 688
rect 1882 682 1889 683
rect 2246 683 2247 687
rect 2251 683 2252 687
rect 2256 683 2257 687
rect 2310 685 2311 689
rect 2315 685 2316 689
rect 2310 684 2316 685
rect 2331 689 2337 690
rect 2331 685 2332 689
rect 2336 685 2337 689
rect 2331 684 2337 685
rect 2390 689 2396 690
rect 2390 685 2391 689
rect 2395 685 2396 689
rect 2454 689 2460 690
rect 2390 684 2396 685
rect 2410 687 2417 688
rect 2246 682 2257 683
rect 2410 683 2411 687
rect 2416 683 2417 687
rect 2454 685 2455 689
rect 2459 685 2460 689
rect 2502 688 2508 689
rect 2454 684 2460 685
rect 2470 687 2481 688
rect 2410 682 2417 683
rect 2470 683 2471 687
rect 2475 683 2476 687
rect 2480 683 2481 687
rect 2502 684 2503 688
rect 2507 684 2508 688
rect 2502 683 2508 684
rect 2470 682 2481 683
rect 1286 678 1292 679
rect 894 675 900 676
rect 1326 671 1332 672
rect 214 668 220 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 214 664 215 668
rect 219 664 220 668
rect 214 663 220 664
rect 294 668 300 669
rect 294 664 295 668
rect 299 664 300 668
rect 294 663 300 664
rect 374 668 380 669
rect 374 664 375 668
rect 379 664 380 668
rect 374 663 380 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 526 668 532 669
rect 526 664 527 668
rect 531 664 532 668
rect 526 663 532 664
rect 590 668 596 669
rect 590 664 591 668
rect 595 664 596 668
rect 590 663 596 664
rect 654 668 660 669
rect 654 664 655 668
rect 659 664 660 668
rect 654 663 660 664
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 782 668 788 669
rect 782 664 783 668
rect 787 664 788 668
rect 782 663 788 664
rect 846 668 852 669
rect 846 664 847 668
rect 851 664 852 668
rect 846 663 852 664
rect 918 668 924 669
rect 918 664 919 668
rect 923 664 924 668
rect 1326 667 1327 671
rect 1331 667 1332 671
rect 2502 671 2508 672
rect 1326 666 1332 667
rect 1350 668 1356 669
rect 918 663 924 664
rect 1286 665 1292 666
rect 110 660 116 661
rect 1286 661 1287 665
rect 1291 661 1292 665
rect 1350 664 1351 668
rect 1355 664 1356 668
rect 1350 663 1356 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1414 663 1420 664
rect 1518 668 1524 669
rect 1518 664 1519 668
rect 1523 664 1524 668
rect 1518 663 1524 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1734 668 1740 669
rect 1734 664 1735 668
rect 1739 664 1740 668
rect 1734 663 1740 664
rect 1846 668 1852 669
rect 1846 664 1847 668
rect 1851 664 1852 668
rect 1846 663 1852 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2134 668 2140 669
rect 2134 664 2135 668
rect 2139 664 2140 668
rect 2134 663 2140 664
rect 2214 668 2220 669
rect 2214 664 2215 668
rect 2219 664 2220 668
rect 2214 663 2220 664
rect 2294 668 2300 669
rect 2294 664 2295 668
rect 2299 664 2300 668
rect 2294 663 2300 664
rect 2374 668 2380 669
rect 2374 664 2375 668
rect 2379 664 2380 668
rect 2374 663 2380 664
rect 2438 668 2444 669
rect 2438 664 2439 668
rect 2443 664 2444 668
rect 2502 667 2503 671
rect 2507 667 2508 671
rect 2502 666 2508 667
rect 2438 663 2444 664
rect 1286 660 1292 661
rect 110 648 116 649
rect 1286 648 1292 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 230 647 236 648
rect 230 643 231 647
rect 235 643 236 647
rect 230 642 236 643
rect 251 647 257 648
rect 251 643 252 647
rect 256 646 257 647
rect 294 647 300 648
rect 294 646 295 647
rect 256 644 295 646
rect 256 643 257 644
rect 251 642 257 643
rect 294 643 295 644
rect 299 643 300 647
rect 294 642 300 643
rect 310 647 316 648
rect 310 643 311 647
rect 315 643 316 647
rect 310 642 316 643
rect 318 647 324 648
rect 318 643 319 647
rect 323 646 324 647
rect 331 647 337 648
rect 331 646 332 647
rect 323 644 332 646
rect 323 643 324 644
rect 318 642 324 643
rect 331 643 332 644
rect 336 643 337 647
rect 331 642 337 643
rect 390 647 396 648
rect 390 643 391 647
rect 395 643 396 647
rect 411 647 417 648
rect 411 646 412 647
rect 390 642 396 643
rect 400 644 412 646
rect 400 638 402 644
rect 411 643 412 644
rect 416 643 417 647
rect 411 642 417 643
rect 470 647 476 648
rect 470 643 471 647
rect 475 643 476 647
rect 470 642 476 643
rect 491 647 500 648
rect 491 643 492 647
rect 499 643 500 647
rect 491 642 500 643
rect 542 647 548 648
rect 542 643 543 647
rect 547 643 548 647
rect 563 647 569 648
rect 563 646 564 647
rect 542 642 548 643
rect 552 644 564 646
rect 552 638 554 644
rect 563 643 564 644
rect 568 643 569 647
rect 563 642 569 643
rect 606 647 612 648
rect 606 643 607 647
rect 611 643 612 647
rect 606 642 612 643
rect 627 647 636 648
rect 627 643 628 647
rect 635 643 636 647
rect 627 642 636 643
rect 670 647 676 648
rect 670 643 671 647
rect 675 643 676 647
rect 691 647 697 648
rect 691 646 692 647
rect 670 642 676 643
rect 680 644 692 646
rect 680 638 682 644
rect 691 643 692 644
rect 696 643 697 647
rect 691 642 697 643
rect 734 647 740 648
rect 734 643 735 647
rect 739 643 740 647
rect 734 642 740 643
rect 750 647 761 648
rect 750 643 751 647
rect 755 643 756 647
rect 760 643 761 647
rect 750 642 761 643
rect 798 647 804 648
rect 798 643 799 647
rect 803 643 804 647
rect 819 647 825 648
rect 819 646 820 647
rect 798 642 804 643
rect 808 644 820 646
rect 808 638 810 644
rect 819 643 820 644
rect 824 643 825 647
rect 819 642 825 643
rect 862 647 868 648
rect 862 643 863 647
rect 867 643 868 647
rect 862 642 868 643
rect 883 647 889 648
rect 883 643 884 647
rect 888 646 889 647
rect 934 647 940 648
rect 888 644 926 646
rect 888 643 889 644
rect 883 642 889 643
rect 319 636 402 638
rect 476 636 554 638
rect 612 636 682 638
rect 740 636 810 638
rect 319 634 321 636
rect 476 634 478 636
rect 612 634 614 636
rect 740 634 742 636
rect 924 634 926 644
rect 934 643 935 647
rect 939 643 940 647
rect 934 642 940 643
rect 942 647 948 648
rect 942 643 943 647
rect 947 646 948 647
rect 955 647 961 648
rect 955 646 956 647
rect 947 644 956 646
rect 947 643 948 644
rect 942 642 948 643
rect 955 643 956 644
rect 960 643 961 647
rect 1286 644 1287 648
rect 1291 644 1292 648
rect 1478 648 1484 649
rect 1286 643 1292 644
rect 1326 645 1332 646
rect 955 642 961 643
rect 1326 641 1327 645
rect 1331 641 1332 645
rect 1478 644 1479 648
rect 1483 644 1484 648
rect 1478 643 1484 644
rect 1558 648 1564 649
rect 1558 644 1559 648
rect 1563 644 1564 648
rect 1558 643 1564 644
rect 1646 648 1652 649
rect 1646 644 1647 648
rect 1651 644 1652 648
rect 1646 643 1652 644
rect 1734 648 1740 649
rect 1734 644 1735 648
rect 1739 644 1740 648
rect 1734 643 1740 644
rect 1830 648 1836 649
rect 1830 644 1831 648
rect 1835 644 1836 648
rect 1830 643 1836 644
rect 1918 648 1924 649
rect 1918 644 1919 648
rect 1923 644 1924 648
rect 1918 643 1924 644
rect 2006 648 2012 649
rect 2006 644 2007 648
rect 2011 644 2012 648
rect 2006 643 2012 644
rect 2086 648 2092 649
rect 2086 644 2087 648
rect 2091 644 2092 648
rect 2086 643 2092 644
rect 2166 648 2172 649
rect 2166 644 2167 648
rect 2171 644 2172 648
rect 2166 643 2172 644
rect 2238 648 2244 649
rect 2238 644 2239 648
rect 2243 644 2244 648
rect 2238 643 2244 644
rect 2310 648 2316 649
rect 2310 644 2311 648
rect 2315 644 2316 648
rect 2310 643 2316 644
rect 2382 648 2388 649
rect 2382 644 2383 648
rect 2387 644 2388 648
rect 2382 643 2388 644
rect 2438 648 2444 649
rect 2438 644 2439 648
rect 2443 644 2444 648
rect 2438 643 2444 644
rect 2502 645 2508 646
rect 1326 640 1332 641
rect 2502 641 2503 645
rect 2507 641 2508 645
rect 2502 640 2508 641
rect 315 633 321 634
rect 222 631 228 632
rect 222 627 223 631
rect 227 630 228 631
rect 235 631 241 632
rect 235 630 236 631
rect 227 628 236 630
rect 227 627 228 628
rect 222 626 228 627
rect 235 627 236 628
rect 240 627 241 631
rect 315 629 316 633
rect 320 629 321 633
rect 475 633 481 634
rect 315 628 321 629
rect 395 631 401 632
rect 235 626 241 627
rect 395 627 396 631
rect 400 630 401 631
rect 426 631 432 632
rect 426 630 427 631
rect 400 628 427 630
rect 400 627 401 628
rect 395 626 401 627
rect 426 627 427 628
rect 431 627 432 631
rect 475 629 476 633
rect 480 629 481 633
rect 611 633 617 634
rect 475 628 481 629
rect 534 631 540 632
rect 426 626 432 627
rect 534 627 535 631
rect 539 630 540 631
rect 547 631 553 632
rect 547 630 548 631
rect 539 628 548 630
rect 539 627 540 628
rect 534 626 540 627
rect 547 627 548 628
rect 552 627 553 631
rect 611 629 612 633
rect 616 629 617 633
rect 739 633 745 634
rect 611 628 617 629
rect 675 631 681 632
rect 547 626 553 627
rect 675 627 676 631
rect 680 630 681 631
rect 680 628 718 630
rect 739 629 740 633
rect 744 629 745 633
rect 924 633 945 634
rect 924 632 940 633
rect 739 628 745 629
rect 803 631 809 632
rect 680 627 681 628
rect 675 626 681 627
rect 716 626 718 628
rect 750 627 756 628
rect 750 626 751 627
rect 716 624 751 626
rect 750 623 751 624
rect 755 623 756 627
rect 803 627 804 631
rect 808 630 809 631
rect 867 631 876 632
rect 808 628 862 630
rect 808 627 809 628
rect 803 626 809 627
rect 750 622 756 623
rect 860 622 862 628
rect 867 627 868 631
rect 875 627 876 631
rect 939 629 940 632
rect 944 629 945 633
rect 939 628 945 629
rect 1326 628 1332 629
rect 2502 628 2508 629
rect 867 626 876 627
rect 1326 624 1327 628
rect 1331 624 1332 628
rect 942 623 948 624
rect 1326 623 1332 624
rect 1494 627 1500 628
rect 1494 623 1495 627
rect 1499 623 1500 627
rect 942 622 943 623
rect 860 620 943 622
rect 942 619 943 620
rect 947 619 948 623
rect 1494 622 1500 623
rect 1515 627 1521 628
rect 1515 623 1516 627
rect 1520 626 1521 627
rect 1574 627 1580 628
rect 1520 624 1566 626
rect 1520 623 1521 624
rect 1515 622 1521 623
rect 942 618 948 619
rect 1106 615 1112 616
rect 1106 614 1107 615
rect 692 612 926 614
rect 692 610 694 612
rect 691 609 697 610
rect 211 607 217 608
rect 211 603 212 607
rect 216 606 217 607
rect 294 607 300 608
rect 216 604 270 606
rect 216 603 217 604
rect 211 602 217 603
rect 268 598 270 604
rect 294 603 295 607
rect 299 606 300 607
rect 307 607 313 608
rect 307 606 308 607
rect 299 604 308 606
rect 299 603 300 604
rect 294 602 300 603
rect 307 603 308 604
rect 312 603 313 607
rect 307 602 313 603
rect 411 607 420 608
rect 411 603 412 607
rect 419 603 420 607
rect 411 602 420 603
rect 494 607 500 608
rect 494 603 495 607
rect 499 606 500 607
rect 507 607 513 608
rect 507 606 508 607
rect 499 604 508 606
rect 499 603 500 604
rect 494 602 500 603
rect 507 603 508 604
rect 512 603 513 607
rect 603 607 609 608
rect 603 606 604 607
rect 507 602 513 603
rect 524 604 604 606
rect 268 596 321 598
rect 319 594 321 596
rect 524 594 526 604
rect 603 603 604 604
rect 608 603 609 607
rect 691 605 692 609
rect 696 605 697 609
rect 771 607 777 608
rect 771 606 772 607
rect 691 604 697 605
rect 708 604 772 606
rect 603 602 609 603
rect 708 594 710 604
rect 771 603 772 604
rect 776 603 777 607
rect 851 607 857 608
rect 851 606 852 607
rect 771 602 777 603
rect 788 604 852 606
rect 788 594 790 604
rect 851 603 852 604
rect 856 603 857 607
rect 851 602 857 603
rect 924 598 926 612
rect 932 612 1107 614
rect 932 610 934 612
rect 1106 611 1107 612
rect 1111 611 1112 615
rect 1564 614 1566 624
rect 1574 623 1575 627
rect 1579 623 1580 627
rect 1574 622 1580 623
rect 1595 627 1601 628
rect 1595 623 1596 627
rect 1600 626 1601 627
rect 1662 627 1668 628
rect 1600 624 1654 626
rect 1600 623 1601 624
rect 1595 622 1601 623
rect 1652 618 1654 624
rect 1662 623 1663 627
rect 1667 623 1668 627
rect 1662 622 1668 623
rect 1678 627 1689 628
rect 1678 623 1679 627
rect 1683 623 1684 627
rect 1688 623 1689 627
rect 1678 622 1689 623
rect 1750 627 1756 628
rect 1750 623 1751 627
rect 1755 623 1756 627
rect 1750 622 1756 623
rect 1758 627 1764 628
rect 1758 623 1759 627
rect 1763 626 1764 627
rect 1771 627 1777 628
rect 1771 626 1772 627
rect 1763 624 1772 626
rect 1763 623 1764 624
rect 1758 622 1764 623
rect 1771 623 1772 624
rect 1776 623 1777 627
rect 1771 622 1777 623
rect 1846 627 1852 628
rect 1846 623 1847 627
rect 1851 623 1852 627
rect 1846 622 1852 623
rect 1862 627 1873 628
rect 1862 623 1863 627
rect 1867 623 1868 627
rect 1872 623 1873 627
rect 1862 622 1873 623
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 1955 627 1961 628
rect 1955 626 1956 627
rect 1934 622 1940 623
rect 1944 624 1956 626
rect 1944 618 1946 624
rect 1955 623 1956 624
rect 1960 623 1961 627
rect 1955 622 1961 623
rect 2022 627 2028 628
rect 2022 623 2023 627
rect 2027 623 2028 627
rect 2022 622 2028 623
rect 2043 627 2049 628
rect 2043 623 2044 627
rect 2048 626 2049 627
rect 2102 627 2108 628
rect 2048 624 2094 626
rect 2048 623 2049 624
rect 2043 622 2049 623
rect 1652 616 1671 618
rect 1669 614 1671 616
rect 1852 616 1946 618
rect 1852 614 1854 616
rect 2092 614 2094 624
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2123 627 2129 628
rect 2123 623 2124 627
rect 2128 626 2129 627
rect 2174 627 2180 628
rect 2174 626 2175 627
rect 2128 624 2175 626
rect 2128 623 2129 624
rect 2123 622 2129 623
rect 2174 623 2175 624
rect 2179 623 2180 627
rect 2174 622 2180 623
rect 2182 627 2188 628
rect 2182 623 2183 627
rect 2187 623 2188 627
rect 2203 627 2209 628
rect 2203 626 2204 627
rect 2182 622 2188 623
rect 2192 624 2204 626
rect 2192 618 2194 624
rect 2203 623 2204 624
rect 2208 623 2209 627
rect 2203 622 2209 623
rect 2254 627 2260 628
rect 2254 623 2255 627
rect 2259 623 2260 627
rect 2254 622 2260 623
rect 2274 627 2281 628
rect 2274 623 2275 627
rect 2280 623 2281 627
rect 2274 622 2281 623
rect 2326 627 2332 628
rect 2326 623 2327 627
rect 2331 623 2332 627
rect 2326 622 2332 623
rect 2342 627 2353 628
rect 2342 623 2343 627
rect 2347 623 2348 627
rect 2352 623 2353 627
rect 2342 622 2353 623
rect 2398 627 2404 628
rect 2398 623 2399 627
rect 2403 623 2404 627
rect 2419 627 2425 628
rect 2419 626 2420 627
rect 2398 622 2404 623
rect 2408 624 2420 626
rect 2408 618 2410 624
rect 2419 623 2420 624
rect 2424 623 2425 627
rect 2419 622 2425 623
rect 2454 627 2460 628
rect 2454 623 2455 627
rect 2459 623 2460 627
rect 2454 622 2460 623
rect 2462 627 2468 628
rect 2462 623 2463 627
rect 2467 626 2468 627
rect 2475 627 2481 628
rect 2475 626 2476 627
rect 2467 624 2476 626
rect 2467 623 2468 624
rect 2462 622 2468 623
rect 2475 623 2476 624
rect 2480 623 2481 627
rect 2502 624 2503 628
rect 2507 624 2508 628
rect 2502 623 2508 624
rect 2475 622 2481 623
rect 2116 616 2194 618
rect 2332 616 2410 618
rect 1564 613 1585 614
rect 1564 612 1580 613
rect 1106 610 1112 611
rect 1499 611 1505 612
rect 931 609 937 610
rect 931 605 932 609
rect 936 605 937 609
rect 931 604 937 605
rect 1011 607 1020 608
rect 1011 603 1012 607
rect 1019 603 1020 607
rect 1091 607 1097 608
rect 1091 606 1092 607
rect 1011 602 1020 603
rect 1029 604 1092 606
rect 924 596 950 598
rect 948 594 950 596
rect 1029 594 1031 604
rect 1091 603 1092 604
rect 1096 603 1097 607
rect 1499 607 1500 611
rect 1504 610 1505 611
rect 1504 608 1575 610
rect 1579 609 1580 612
rect 1584 609 1585 613
rect 1579 608 1585 609
rect 1667 613 1673 614
rect 1667 609 1668 613
rect 1672 609 1673 613
rect 1851 613 1857 614
rect 1667 608 1673 609
rect 1755 611 1761 612
rect 1504 607 1505 608
rect 1499 606 1505 607
rect 1573 606 1575 608
rect 1654 607 1660 608
rect 1654 606 1655 607
rect 1573 604 1655 606
rect 1091 602 1097 603
rect 1654 603 1655 604
rect 1659 603 1660 607
rect 1755 607 1756 611
rect 1760 607 1761 611
rect 1851 609 1852 613
rect 1856 609 1857 613
rect 2092 613 2113 614
rect 2092 612 2108 613
rect 1851 608 1857 609
rect 1902 611 1908 612
rect 1755 606 1761 607
rect 1862 607 1868 608
rect 1862 606 1863 607
rect 1757 604 1863 606
rect 1654 602 1660 603
rect 1862 603 1863 604
rect 1867 603 1868 607
rect 1902 607 1903 611
rect 1907 610 1908 611
rect 1939 611 1945 612
rect 1939 610 1940 611
rect 1907 608 1940 610
rect 1907 607 1908 608
rect 1902 606 1908 607
rect 1939 607 1940 608
rect 1944 607 1945 611
rect 1939 606 1945 607
rect 2027 611 2033 612
rect 2027 607 2028 611
rect 2032 610 2033 611
rect 2032 608 2102 610
rect 2107 609 2108 612
rect 2112 609 2113 613
rect 2107 608 2113 609
rect 2032 607 2033 608
rect 2027 606 2033 607
rect 2100 606 2102 608
rect 2116 606 2118 616
rect 2332 614 2334 616
rect 2331 613 2337 614
rect 2187 611 2193 612
rect 2187 607 2188 611
rect 2192 610 2193 611
rect 2246 611 2252 612
rect 2246 610 2247 611
rect 2192 608 2247 610
rect 2192 607 2193 608
rect 2187 606 2193 607
rect 2246 607 2247 608
rect 2251 607 2252 611
rect 2246 606 2252 607
rect 2259 611 2265 612
rect 2259 607 2260 611
rect 2264 610 2265 611
rect 2264 608 2306 610
rect 2331 609 2332 613
rect 2336 609 2337 613
rect 2331 608 2337 609
rect 2403 611 2412 612
rect 2264 607 2265 608
rect 2259 606 2265 607
rect 2304 606 2306 608
rect 2342 607 2348 608
rect 2342 606 2343 607
rect 2100 604 2118 606
rect 2304 604 2343 606
rect 1862 602 1868 603
rect 2342 603 2343 604
rect 2347 603 2348 607
rect 2403 607 2404 611
rect 2411 607 2412 611
rect 2403 606 2412 607
rect 2459 611 2465 612
rect 2459 607 2460 611
rect 2464 610 2465 611
rect 2470 611 2476 612
rect 2470 610 2471 611
rect 2464 608 2471 610
rect 2464 607 2465 608
rect 2459 606 2465 607
rect 2470 607 2471 608
rect 2475 607 2476 611
rect 2470 606 2476 607
rect 2342 602 2348 603
rect 2298 595 2304 596
rect 2298 594 2299 595
rect 206 593 212 594
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 206 589 207 593
rect 211 589 212 593
rect 302 593 308 594
rect 206 588 212 589
rect 214 591 220 592
rect 110 587 116 588
rect 214 587 215 591
rect 219 590 220 591
rect 227 591 233 592
rect 227 590 228 591
rect 219 588 228 590
rect 219 587 220 588
rect 214 586 220 587
rect 227 587 228 588
rect 232 587 233 591
rect 302 589 303 593
rect 307 589 308 593
rect 319 593 329 594
rect 319 592 324 593
rect 302 588 308 589
rect 323 589 324 592
rect 328 589 329 593
rect 323 588 329 589
rect 406 593 412 594
rect 406 589 407 593
rect 411 589 412 593
rect 502 593 508 594
rect 406 588 412 589
rect 426 591 433 592
rect 227 586 233 587
rect 426 587 427 591
rect 432 587 433 591
rect 502 589 503 593
rect 507 589 508 593
rect 502 588 508 589
rect 523 593 529 594
rect 523 589 524 593
rect 528 589 529 593
rect 523 588 529 589
rect 598 593 604 594
rect 598 589 599 593
rect 603 589 604 593
rect 686 593 692 594
rect 598 588 604 589
rect 619 591 628 592
rect 426 586 433 587
rect 619 587 620 591
rect 627 587 628 591
rect 686 589 687 593
rect 691 589 692 593
rect 686 588 692 589
rect 707 593 713 594
rect 707 589 708 593
rect 712 589 713 593
rect 707 588 713 589
rect 766 593 772 594
rect 766 589 767 593
rect 771 589 772 593
rect 766 588 772 589
rect 787 593 793 594
rect 787 589 788 593
rect 792 589 793 593
rect 787 588 793 589
rect 846 593 852 594
rect 846 589 847 593
rect 851 589 852 593
rect 926 593 932 594
rect 846 588 852 589
rect 867 591 876 592
rect 619 586 628 587
rect 867 587 868 591
rect 875 587 876 591
rect 926 589 927 593
rect 931 589 932 593
rect 926 588 932 589
rect 947 593 953 594
rect 947 589 948 593
rect 952 589 953 593
rect 947 588 953 589
rect 1006 593 1012 594
rect 1006 589 1007 593
rect 1011 589 1012 593
rect 1006 588 1012 589
rect 1027 593 1033 594
rect 1027 589 1028 593
rect 1032 589 1033 593
rect 1027 588 1033 589
rect 1086 593 1092 594
rect 1086 589 1087 593
rect 1091 589 1092 593
rect 1286 592 1292 593
rect 1086 588 1092 589
rect 1106 591 1113 592
rect 867 586 876 587
rect 1106 587 1107 591
rect 1112 587 1113 591
rect 1286 588 1287 592
rect 1291 588 1292 592
rect 1988 592 2299 594
rect 1988 590 1990 592
rect 2298 591 2299 592
rect 2303 591 2304 595
rect 2298 590 2304 591
rect 1987 589 1993 590
rect 1286 587 1292 588
rect 1459 587 1465 588
rect 1106 586 1113 587
rect 1459 583 1460 587
rect 1464 583 1465 587
rect 1459 582 1465 583
rect 1563 587 1569 588
rect 1563 583 1564 587
rect 1568 586 1569 587
rect 1675 587 1684 588
rect 1568 584 1671 586
rect 1568 583 1569 584
rect 1563 582 1569 583
rect 1461 578 1463 582
rect 1669 578 1671 584
rect 1675 583 1676 587
rect 1683 583 1684 587
rect 1675 582 1684 583
rect 1779 587 1785 588
rect 1779 583 1780 587
rect 1784 586 1785 587
rect 1834 587 1840 588
rect 1834 586 1835 587
rect 1784 584 1835 586
rect 1784 583 1785 584
rect 1779 582 1785 583
rect 1834 583 1835 584
rect 1839 583 1840 587
rect 1883 587 1889 588
rect 1883 586 1884 587
rect 1834 582 1840 583
rect 1844 584 1884 586
rect 1844 578 1846 584
rect 1883 583 1884 584
rect 1888 583 1889 587
rect 1987 585 1988 589
rect 1992 585 1993 589
rect 1987 584 1993 585
rect 2091 587 2097 588
rect 1883 582 1889 583
rect 2091 583 2092 587
rect 2096 583 2097 587
rect 2091 582 2097 583
rect 2174 587 2180 588
rect 2174 583 2175 587
rect 2179 586 2180 587
rect 2187 587 2193 588
rect 2187 586 2188 587
rect 2179 584 2188 586
rect 2179 583 2180 584
rect 2174 582 2180 583
rect 2187 583 2188 584
rect 2192 583 2193 587
rect 2283 587 2289 588
rect 2283 586 2284 587
rect 2187 582 2193 583
rect 2204 584 2284 586
rect 2093 578 2095 582
rect 1461 576 1582 578
rect 1669 576 1694 578
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 1286 575 1292 576
rect 110 570 116 571
rect 190 572 196 573
rect 190 568 191 572
rect 195 568 196 572
rect 190 567 196 568
rect 286 572 292 573
rect 286 568 287 572
rect 291 568 292 572
rect 286 567 292 568
rect 390 572 396 573
rect 390 568 391 572
rect 395 568 396 572
rect 390 567 396 568
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 670 572 676 573
rect 670 568 671 572
rect 675 568 676 572
rect 670 567 676 568
rect 750 572 756 573
rect 750 568 751 572
rect 755 568 756 572
rect 750 567 756 568
rect 830 572 836 573
rect 830 568 831 572
rect 835 568 836 572
rect 830 567 836 568
rect 910 572 916 573
rect 910 568 911 572
rect 915 568 916 572
rect 910 567 916 568
rect 990 572 996 573
rect 990 568 991 572
rect 995 568 996 572
rect 990 567 996 568
rect 1070 572 1076 573
rect 1070 568 1071 572
rect 1075 568 1076 572
rect 1286 571 1287 575
rect 1291 571 1292 575
rect 1580 574 1582 576
rect 1692 574 1694 576
rect 1796 576 1846 578
rect 2004 576 2095 578
rect 1796 574 1798 576
rect 2004 574 2006 576
rect 2204 574 2206 584
rect 2283 583 2284 584
rect 2288 583 2289 587
rect 2283 582 2289 583
rect 2379 587 2388 588
rect 2379 583 2380 587
rect 2387 583 2388 587
rect 2379 582 2388 583
rect 2459 587 2468 588
rect 2459 583 2460 587
rect 2467 583 2468 587
rect 2459 582 2468 583
rect 1454 573 1460 574
rect 1286 570 1292 571
rect 1326 572 1332 573
rect 1070 567 1076 568
rect 1326 568 1327 572
rect 1331 568 1332 572
rect 1454 569 1455 573
rect 1459 569 1460 573
rect 1558 573 1564 574
rect 1454 568 1460 569
rect 1470 571 1481 572
rect 1326 567 1332 568
rect 1470 567 1471 571
rect 1475 567 1476 571
rect 1480 567 1481 571
rect 1558 569 1559 573
rect 1563 569 1564 573
rect 1558 568 1564 569
rect 1579 573 1585 574
rect 1579 569 1580 573
rect 1584 569 1585 573
rect 1579 568 1585 569
rect 1670 573 1676 574
rect 1670 569 1671 573
rect 1675 569 1676 573
rect 1670 568 1676 569
rect 1691 573 1697 574
rect 1691 569 1692 573
rect 1696 569 1697 573
rect 1691 568 1697 569
rect 1774 573 1780 574
rect 1774 569 1775 573
rect 1779 569 1780 573
rect 1774 568 1780 569
rect 1795 573 1801 574
rect 1795 569 1796 573
rect 1800 569 1801 573
rect 1795 568 1801 569
rect 1878 573 1884 574
rect 1878 569 1879 573
rect 1883 569 1884 573
rect 1982 573 1988 574
rect 1878 568 1884 569
rect 1899 571 1908 572
rect 1470 566 1481 567
rect 1899 567 1900 571
rect 1907 567 1908 571
rect 1982 569 1983 573
rect 1987 569 1988 573
rect 1982 568 1988 569
rect 2003 573 2009 574
rect 2003 569 2004 573
rect 2008 569 2009 573
rect 2003 568 2009 569
rect 2086 573 2092 574
rect 2086 569 2087 573
rect 2091 569 2092 573
rect 2182 573 2188 574
rect 2086 568 2092 569
rect 2107 571 2113 572
rect 1899 566 1908 567
rect 2107 567 2108 571
rect 2112 570 2113 571
rect 2158 571 2164 572
rect 2158 570 2159 571
rect 2112 568 2159 570
rect 2112 567 2113 568
rect 2107 566 2113 567
rect 2158 567 2159 568
rect 2163 567 2164 571
rect 2182 569 2183 573
rect 2187 569 2188 573
rect 2182 568 2188 569
rect 2203 573 2209 574
rect 2203 569 2204 573
rect 2208 569 2209 573
rect 2203 568 2209 569
rect 2278 573 2284 574
rect 2278 569 2279 573
rect 2283 569 2284 573
rect 2374 573 2380 574
rect 2278 568 2284 569
rect 2298 571 2305 572
rect 2158 566 2164 567
rect 2298 567 2299 571
rect 2304 567 2305 571
rect 2374 569 2375 573
rect 2379 569 2380 573
rect 2454 573 2460 574
rect 2374 568 2380 569
rect 2395 571 2401 572
rect 2298 566 2305 567
rect 2395 567 2396 571
rect 2400 570 2401 571
rect 2406 571 2412 572
rect 2406 570 2407 571
rect 2400 568 2407 570
rect 2400 567 2401 568
rect 2395 566 2401 567
rect 2406 567 2407 568
rect 2411 567 2412 571
rect 2454 569 2455 573
rect 2459 569 2460 573
rect 2502 572 2508 573
rect 2454 568 2460 569
rect 2462 571 2468 572
rect 2406 566 2412 567
rect 2462 567 2463 571
rect 2467 570 2468 571
rect 2475 571 2481 572
rect 2475 570 2476 571
rect 2467 568 2476 570
rect 2467 567 2468 568
rect 2462 566 2468 567
rect 2475 567 2476 568
rect 2480 567 2481 571
rect 2502 568 2503 572
rect 2507 568 2508 572
rect 2502 567 2508 568
rect 2475 566 2481 567
rect 174 556 180 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 270 556 276 557
rect 270 552 271 556
rect 275 552 276 556
rect 270 551 276 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 486 556 492 557
rect 486 552 487 556
rect 491 552 492 556
rect 486 551 492 552
rect 590 556 596 557
rect 590 552 591 556
rect 595 552 596 556
rect 590 551 596 552
rect 694 556 700 557
rect 694 552 695 556
rect 699 552 700 556
rect 694 551 700 552
rect 790 556 796 557
rect 790 552 791 556
rect 795 552 796 556
rect 790 551 796 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 966 556 972 557
rect 966 552 967 556
rect 971 552 972 556
rect 966 551 972 552
rect 1054 556 1060 557
rect 1054 552 1055 556
rect 1059 552 1060 556
rect 1054 551 1060 552
rect 1150 556 1156 557
rect 1150 552 1151 556
rect 1155 552 1156 556
rect 1326 555 1332 556
rect 1150 551 1156 552
rect 1286 553 1292 554
rect 110 548 116 549
rect 1286 549 1287 553
rect 1291 549 1292 553
rect 1326 551 1327 555
rect 1331 551 1332 555
rect 2502 555 2508 556
rect 1326 550 1332 551
rect 1438 552 1444 553
rect 1286 548 1292 549
rect 1438 548 1439 552
rect 1443 548 1444 552
rect 1438 547 1444 548
rect 1542 552 1548 553
rect 1542 548 1543 552
rect 1547 548 1548 552
rect 1542 547 1548 548
rect 1654 552 1660 553
rect 1654 548 1655 552
rect 1659 548 1660 552
rect 1654 547 1660 548
rect 1758 552 1764 553
rect 1758 548 1759 552
rect 1763 548 1764 552
rect 1758 547 1764 548
rect 1862 552 1868 553
rect 1862 548 1863 552
rect 1867 548 1868 552
rect 1862 547 1868 548
rect 1966 552 1972 553
rect 1966 548 1967 552
rect 1971 548 1972 552
rect 1966 547 1972 548
rect 2070 552 2076 553
rect 2070 548 2071 552
rect 2075 548 2076 552
rect 2070 547 2076 548
rect 2166 552 2172 553
rect 2166 548 2167 552
rect 2171 548 2172 552
rect 2166 547 2172 548
rect 2262 552 2268 553
rect 2262 548 2263 552
rect 2267 548 2268 552
rect 2262 547 2268 548
rect 2358 552 2364 553
rect 2358 548 2359 552
rect 2363 548 2364 552
rect 2358 547 2364 548
rect 2438 552 2444 553
rect 2438 548 2439 552
rect 2443 548 2444 552
rect 2502 551 2503 555
rect 2507 551 2508 555
rect 2502 550 2508 551
rect 2438 547 2444 548
rect 110 536 116 537
rect 1286 536 1292 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 190 535 196 536
rect 190 531 191 535
rect 195 531 196 535
rect 190 530 196 531
rect 211 535 217 536
rect 211 531 212 535
rect 216 534 217 535
rect 238 535 244 536
rect 238 534 239 535
rect 216 532 239 534
rect 216 531 217 532
rect 211 530 217 531
rect 238 531 239 532
rect 243 531 244 535
rect 238 530 244 531
rect 286 535 292 536
rect 286 531 287 535
rect 291 531 292 535
rect 286 530 292 531
rect 307 535 313 536
rect 307 531 308 535
rect 312 534 313 535
rect 390 535 396 536
rect 312 532 321 534
rect 312 531 313 532
rect 307 530 313 531
rect 319 522 321 532
rect 390 531 391 535
rect 395 531 396 535
rect 390 530 396 531
rect 411 535 420 536
rect 411 531 412 535
rect 419 531 420 535
rect 411 530 420 531
rect 502 535 508 536
rect 502 531 503 535
rect 507 531 508 535
rect 502 530 508 531
rect 523 535 529 536
rect 523 531 524 535
rect 528 534 529 535
rect 606 535 612 536
rect 528 532 598 534
rect 528 531 529 532
rect 523 530 529 531
rect 596 522 598 532
rect 606 531 607 535
rect 611 531 612 535
rect 606 530 612 531
rect 627 535 633 536
rect 627 531 628 535
rect 632 534 633 535
rect 710 535 716 536
rect 632 532 702 534
rect 632 531 633 532
rect 627 530 633 531
rect 700 522 702 532
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 731 535 737 536
rect 731 531 732 535
rect 736 534 737 535
rect 742 535 748 536
rect 742 534 743 535
rect 736 532 743 534
rect 736 531 737 532
rect 731 530 737 531
rect 742 531 743 532
rect 747 531 748 535
rect 742 530 748 531
rect 806 535 812 536
rect 806 531 807 535
rect 811 531 812 535
rect 806 530 812 531
rect 827 535 833 536
rect 827 531 828 535
rect 832 531 833 535
rect 827 530 833 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 915 535 921 536
rect 915 531 916 535
rect 920 534 921 535
rect 982 535 988 536
rect 920 532 974 534
rect 920 531 921 532
rect 915 530 921 531
rect 829 522 831 530
rect 972 522 974 532
rect 982 531 983 535
rect 987 531 988 535
rect 982 530 988 531
rect 1003 535 1009 536
rect 1003 531 1004 535
rect 1008 534 1009 535
rect 1014 535 1020 536
rect 1014 534 1015 535
rect 1008 532 1015 534
rect 1008 531 1009 532
rect 1003 530 1009 531
rect 1014 531 1015 532
rect 1019 531 1020 535
rect 1014 530 1020 531
rect 1070 535 1076 536
rect 1070 531 1071 535
rect 1075 531 1076 535
rect 1070 530 1076 531
rect 1091 535 1097 536
rect 1091 531 1092 535
rect 1096 534 1097 535
rect 1166 535 1172 536
rect 1096 532 1161 534
rect 1096 531 1097 532
rect 1091 530 1097 531
rect 1159 522 1161 532
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1166 530 1172 531
rect 1174 535 1180 536
rect 1174 531 1175 535
rect 1179 534 1180 535
rect 1187 535 1193 536
rect 1187 534 1188 535
rect 1179 532 1188 534
rect 1179 531 1180 532
rect 1174 530 1180 531
rect 1187 531 1188 532
rect 1192 531 1193 535
rect 1286 532 1287 536
rect 1291 532 1292 536
rect 1366 536 1372 537
rect 1286 531 1292 532
rect 1326 533 1332 534
rect 1187 530 1193 531
rect 1326 529 1327 533
rect 1331 529 1332 533
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1446 536 1452 537
rect 1446 532 1447 536
rect 1451 532 1452 536
rect 1446 531 1452 532
rect 1526 536 1532 537
rect 1526 532 1527 536
rect 1531 532 1532 536
rect 1526 531 1532 532
rect 1614 536 1620 537
rect 1614 532 1615 536
rect 1619 532 1620 536
rect 1614 531 1620 532
rect 1710 536 1716 537
rect 1710 532 1711 536
rect 1715 532 1716 536
rect 1710 531 1716 532
rect 1798 536 1804 537
rect 1798 532 1799 536
rect 1803 532 1804 536
rect 1798 531 1804 532
rect 1886 536 1892 537
rect 1886 532 1887 536
rect 1891 532 1892 536
rect 1886 531 1892 532
rect 1974 536 1980 537
rect 1974 532 1975 536
rect 1979 532 1980 536
rect 1974 531 1980 532
rect 2062 536 2068 537
rect 2062 532 2063 536
rect 2067 532 2068 536
rect 2062 531 2068 532
rect 2150 536 2156 537
rect 2150 532 2151 536
rect 2155 532 2156 536
rect 2150 531 2156 532
rect 2246 536 2252 537
rect 2246 532 2247 536
rect 2251 532 2252 536
rect 2246 531 2252 532
rect 2342 536 2348 537
rect 2342 532 2343 536
rect 2347 532 2348 536
rect 2342 531 2348 532
rect 2438 536 2444 537
rect 2438 532 2439 536
rect 2443 532 2444 536
rect 2438 531 2444 532
rect 2502 533 2508 534
rect 1326 528 1332 529
rect 2502 529 2503 533
rect 2507 529 2508 533
rect 2502 528 2508 529
rect 319 521 401 522
rect 319 520 396 521
rect 195 519 201 520
rect 195 515 196 519
rect 200 518 201 519
rect 214 519 220 520
rect 214 518 215 519
rect 200 516 215 518
rect 200 515 201 516
rect 195 514 201 515
rect 214 515 215 516
rect 219 515 220 519
rect 214 514 220 515
rect 291 519 297 520
rect 291 515 292 519
rect 296 518 297 519
rect 296 516 321 518
rect 395 517 396 520
rect 400 517 401 521
rect 596 521 617 522
rect 596 520 612 521
rect 395 516 401 517
rect 507 519 513 520
rect 296 515 297 516
rect 291 514 297 515
rect 319 514 321 516
rect 494 515 500 516
rect 494 514 495 515
rect 319 512 495 514
rect 494 511 495 512
rect 499 511 500 515
rect 507 515 508 519
rect 512 518 513 519
rect 512 516 566 518
rect 611 517 612 520
rect 616 517 617 521
rect 700 521 721 522
rect 700 520 716 521
rect 611 516 617 517
rect 715 517 716 520
rect 720 517 721 521
rect 829 521 905 522
rect 829 520 900 521
rect 715 516 721 517
rect 811 519 817 520
rect 512 515 513 516
rect 507 514 513 515
rect 564 514 566 516
rect 622 515 628 516
rect 622 514 623 515
rect 564 512 623 514
rect 494 510 500 511
rect 622 511 623 512
rect 627 511 628 515
rect 811 515 812 519
rect 816 518 817 519
rect 816 516 894 518
rect 899 517 900 520
rect 904 517 905 521
rect 972 521 993 522
rect 972 520 988 521
rect 899 516 905 517
rect 987 517 988 520
rect 992 517 993 521
rect 1159 521 1177 522
rect 1159 520 1172 521
rect 987 516 993 517
rect 1075 519 1084 520
rect 816 515 817 516
rect 811 514 817 515
rect 622 510 628 511
rect 892 510 894 516
rect 1075 515 1076 519
rect 1083 515 1084 519
rect 1171 517 1172 520
rect 1176 517 1177 521
rect 1171 516 1177 517
rect 1326 516 1332 517
rect 2502 516 2508 517
rect 1075 514 1084 515
rect 1326 512 1327 516
rect 1331 512 1332 516
rect 1174 511 1180 512
rect 1326 511 1332 512
rect 1382 515 1388 516
rect 1382 511 1383 515
rect 1387 511 1388 515
rect 1174 510 1175 511
rect 892 508 1175 510
rect 1174 507 1175 508
rect 1179 507 1180 511
rect 1382 510 1388 511
rect 1390 515 1396 516
rect 1390 511 1391 515
rect 1395 514 1396 515
rect 1403 515 1409 516
rect 1403 514 1404 515
rect 1395 512 1404 514
rect 1395 511 1396 512
rect 1390 510 1396 511
rect 1403 511 1404 512
rect 1408 511 1409 515
rect 1403 510 1409 511
rect 1462 515 1468 516
rect 1462 511 1463 515
rect 1467 511 1468 515
rect 1462 510 1468 511
rect 1483 515 1489 516
rect 1483 511 1484 515
rect 1488 511 1489 515
rect 1483 510 1489 511
rect 1542 515 1548 516
rect 1542 511 1543 515
rect 1547 511 1548 515
rect 1542 510 1548 511
rect 1550 515 1556 516
rect 1550 511 1551 515
rect 1555 514 1556 515
rect 1563 515 1569 516
rect 1563 514 1564 515
rect 1555 512 1564 514
rect 1555 511 1556 512
rect 1550 510 1556 511
rect 1563 511 1564 512
rect 1568 511 1569 515
rect 1563 510 1569 511
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 1651 515 1657 516
rect 1651 511 1652 515
rect 1656 511 1657 515
rect 1651 510 1657 511
rect 1726 515 1732 516
rect 1726 511 1727 515
rect 1731 511 1732 515
rect 1726 510 1732 511
rect 1747 515 1753 516
rect 1747 511 1748 515
rect 1752 511 1753 515
rect 1747 510 1753 511
rect 1814 515 1820 516
rect 1814 511 1815 515
rect 1819 511 1820 515
rect 1814 510 1820 511
rect 1834 515 1841 516
rect 1834 511 1835 515
rect 1840 511 1841 515
rect 1834 510 1841 511
rect 1902 515 1908 516
rect 1902 511 1903 515
rect 1907 511 1908 515
rect 1902 510 1908 511
rect 1923 515 1929 516
rect 1923 511 1924 515
rect 1928 511 1929 515
rect 1923 510 1929 511
rect 1990 515 1996 516
rect 1990 511 1991 515
rect 1995 511 1996 515
rect 1990 510 1996 511
rect 2011 515 2017 516
rect 2011 511 2012 515
rect 2016 514 2017 515
rect 2078 515 2084 516
rect 2016 512 2070 514
rect 2016 511 2017 512
rect 2011 510 2017 511
rect 1174 506 1180 507
rect 1178 503 1184 504
rect 1178 502 1179 503
rect 852 500 1179 502
rect 852 498 854 500
rect 1178 499 1179 500
rect 1183 499 1184 503
rect 1485 502 1487 510
rect 1653 502 1655 510
rect 1749 502 1751 510
rect 1925 502 1927 510
rect 2068 502 2070 512
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2099 515 2105 516
rect 2099 511 2100 515
rect 2104 514 2105 515
rect 2150 515 2156 516
rect 2150 514 2151 515
rect 2104 512 2151 514
rect 2104 511 2105 512
rect 2099 510 2105 511
rect 2150 511 2151 512
rect 2155 511 2156 515
rect 2150 510 2156 511
rect 2166 515 2172 516
rect 2166 511 2167 515
rect 2171 511 2172 515
rect 2166 510 2172 511
rect 2187 515 2193 516
rect 2187 511 2188 515
rect 2192 514 2193 515
rect 2262 515 2268 516
rect 2192 512 2258 514
rect 2192 511 2193 512
rect 2187 510 2193 511
rect 2256 502 2258 512
rect 2262 511 2263 515
rect 2267 511 2268 515
rect 2262 510 2268 511
rect 2270 515 2276 516
rect 2270 511 2271 515
rect 2275 514 2276 515
rect 2283 515 2289 516
rect 2283 514 2284 515
rect 2275 512 2284 514
rect 2275 511 2276 512
rect 2270 510 2276 511
rect 2283 511 2284 512
rect 2288 511 2289 515
rect 2283 510 2289 511
rect 2358 515 2364 516
rect 2358 511 2359 515
rect 2363 511 2364 515
rect 2358 510 2364 511
rect 2379 515 2388 516
rect 2379 511 2380 515
rect 2387 511 2388 515
rect 2379 510 2388 511
rect 2454 515 2460 516
rect 2454 511 2455 515
rect 2459 511 2460 515
rect 2454 510 2460 511
rect 2475 515 2481 516
rect 2475 511 2476 515
rect 2480 511 2481 515
rect 2502 512 2503 516
rect 2507 512 2508 516
rect 2502 511 2508 512
rect 2475 510 2481 511
rect 2477 506 2479 510
rect 2364 504 2479 506
rect 2364 502 2366 504
rect 1485 501 1553 502
rect 1485 500 1548 501
rect 1178 498 1184 499
rect 1387 499 1393 500
rect 851 497 857 498
rect 155 495 161 496
rect 155 491 156 495
rect 160 494 161 495
rect 238 495 244 496
rect 160 492 234 494
rect 160 491 161 492
rect 155 490 161 491
rect 232 486 234 492
rect 238 491 239 495
rect 243 494 244 495
rect 251 495 257 496
rect 251 494 252 495
rect 243 492 252 494
rect 243 491 244 492
rect 238 490 244 491
rect 251 491 252 492
rect 256 491 257 495
rect 251 490 257 491
rect 342 495 348 496
rect 342 491 343 495
rect 347 494 348 495
rect 371 495 377 496
rect 371 494 372 495
rect 347 492 372 494
rect 347 491 348 492
rect 342 490 348 491
rect 371 491 372 492
rect 376 491 377 495
rect 491 495 497 496
rect 491 494 492 495
rect 371 490 377 491
rect 388 492 492 494
rect 232 484 270 486
rect 268 482 270 484
rect 388 482 390 492
rect 491 491 492 492
rect 496 491 497 495
rect 491 490 497 491
rect 619 495 625 496
rect 619 491 620 495
rect 624 494 625 495
rect 739 495 748 496
rect 624 492 735 494
rect 624 491 625 492
rect 619 490 625 491
rect 733 486 735 492
rect 739 491 740 495
rect 747 491 748 495
rect 851 493 852 497
rect 856 493 857 497
rect 955 495 961 496
rect 955 494 956 495
rect 851 492 857 493
rect 868 492 956 494
rect 739 490 748 491
rect 733 484 758 486
rect 756 482 758 484
rect 868 482 870 492
rect 955 491 956 492
rect 960 491 961 495
rect 1059 495 1065 496
rect 1059 494 1060 495
rect 955 490 961 491
rect 972 492 1060 494
rect 972 482 974 492
rect 1059 491 1060 492
rect 1064 491 1065 495
rect 1059 490 1065 491
rect 1163 495 1169 496
rect 1163 491 1164 495
rect 1168 494 1169 495
rect 1243 495 1249 496
rect 1168 492 1222 494
rect 1168 491 1169 492
rect 1163 490 1169 491
rect 1220 486 1222 492
rect 1243 491 1244 495
rect 1248 494 1249 495
rect 1258 495 1264 496
rect 1258 494 1259 495
rect 1248 492 1259 494
rect 1248 491 1249 492
rect 1243 490 1249 491
rect 1258 491 1259 492
rect 1263 491 1264 495
rect 1387 495 1388 499
rect 1392 495 1393 499
rect 1387 494 1393 495
rect 1467 499 1476 500
rect 1467 495 1468 499
rect 1475 495 1476 499
rect 1547 497 1548 500
rect 1552 497 1553 501
rect 1653 501 1737 502
rect 1653 500 1732 501
rect 1547 496 1553 497
rect 1635 499 1641 500
rect 1467 494 1476 495
rect 1635 495 1636 499
rect 1640 498 1641 499
rect 1640 496 1722 498
rect 1731 497 1732 500
rect 1736 497 1737 501
rect 1749 501 1825 502
rect 1749 500 1820 501
rect 1731 496 1737 497
rect 1819 497 1820 500
rect 1824 497 1825 501
rect 1925 501 2001 502
rect 1925 500 1996 501
rect 1819 496 1825 497
rect 1907 499 1913 500
rect 1640 495 1641 496
rect 1635 494 1641 495
rect 1718 495 1724 496
rect 1258 490 1264 491
rect 1389 490 1391 494
rect 1550 491 1556 492
rect 1550 490 1551 491
rect 1389 488 1551 490
rect 1550 487 1551 488
rect 1555 487 1556 491
rect 1718 491 1719 495
rect 1723 491 1724 495
rect 1907 495 1908 499
rect 1912 498 1913 499
rect 1912 496 1958 498
rect 1995 497 1996 500
rect 2000 497 2001 501
rect 2068 501 2089 502
rect 2068 500 2084 501
rect 1995 496 2001 497
rect 2083 497 2084 500
rect 2088 497 2089 501
rect 2256 501 2273 502
rect 2256 500 2268 501
rect 2083 496 2089 497
rect 2158 499 2164 500
rect 1912 495 1913 496
rect 1907 494 1913 495
rect 1956 494 1958 496
rect 2054 495 2060 496
rect 2054 494 2055 495
rect 1956 492 2055 494
rect 1718 490 1724 491
rect 2054 491 2055 492
rect 2059 491 2060 495
rect 2158 495 2159 499
rect 2163 498 2164 499
rect 2171 499 2177 500
rect 2171 498 2172 499
rect 2163 496 2172 498
rect 2163 495 2164 496
rect 2158 494 2164 495
rect 2171 495 2172 496
rect 2176 495 2177 499
rect 2267 497 2268 500
rect 2272 497 2273 501
rect 2267 496 2273 497
rect 2363 501 2369 502
rect 2363 497 2364 501
rect 2368 497 2369 501
rect 2363 496 2369 497
rect 2459 499 2465 500
rect 2171 494 2177 495
rect 2459 495 2460 499
rect 2464 498 2465 499
rect 2478 499 2484 500
rect 2478 498 2479 499
rect 2464 496 2479 498
rect 2464 495 2465 496
rect 2459 494 2465 495
rect 2478 495 2479 496
rect 2483 495 2484 499
rect 2478 494 2484 495
rect 2054 490 2060 491
rect 1550 486 1556 487
rect 1220 484 1262 486
rect 1260 482 1262 484
rect 1390 483 1396 484
rect 1390 482 1391 483
rect 150 481 156 482
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 150 477 151 481
rect 155 477 156 481
rect 246 481 252 482
rect 150 476 156 477
rect 158 479 164 480
rect 110 475 116 476
rect 158 475 159 479
rect 163 478 164 479
rect 171 479 177 480
rect 171 478 172 479
rect 163 476 172 478
rect 163 475 164 476
rect 158 474 164 475
rect 171 475 172 476
rect 176 475 177 479
rect 246 477 247 481
rect 251 477 252 481
rect 246 476 252 477
rect 267 481 273 482
rect 267 477 268 481
rect 272 477 273 481
rect 267 476 273 477
rect 366 481 372 482
rect 366 477 367 481
rect 371 477 372 481
rect 366 476 372 477
rect 387 481 393 482
rect 387 477 388 481
rect 392 477 393 481
rect 387 476 393 477
rect 486 481 492 482
rect 486 477 487 481
rect 491 477 492 481
rect 614 481 620 482
rect 486 476 492 477
rect 494 479 500 480
rect 171 474 177 475
rect 494 475 495 479
rect 499 478 500 479
rect 507 479 513 480
rect 507 478 508 479
rect 499 476 508 478
rect 499 475 500 476
rect 494 474 500 475
rect 507 475 508 476
rect 512 475 513 479
rect 614 477 615 481
rect 619 477 620 481
rect 734 481 740 482
rect 614 476 620 477
rect 622 479 628 480
rect 507 474 513 475
rect 622 475 623 479
rect 627 478 628 479
rect 635 479 641 480
rect 635 478 636 479
rect 627 476 636 478
rect 627 475 628 476
rect 622 474 628 475
rect 635 475 636 476
rect 640 475 641 479
rect 734 477 735 481
rect 739 477 740 481
rect 734 476 740 477
rect 755 481 761 482
rect 755 477 756 481
rect 760 477 761 481
rect 755 476 761 477
rect 846 481 852 482
rect 846 477 847 481
rect 851 477 852 481
rect 846 476 852 477
rect 867 481 873 482
rect 867 477 868 481
rect 872 477 873 481
rect 867 476 873 477
rect 950 481 956 482
rect 950 477 951 481
rect 955 477 956 481
rect 950 476 956 477
rect 971 481 977 482
rect 971 477 972 481
rect 976 477 977 481
rect 971 476 977 477
rect 1054 481 1060 482
rect 1054 477 1055 481
rect 1059 477 1060 481
rect 1158 481 1164 482
rect 1054 476 1060 477
rect 1075 479 1084 480
rect 635 474 641 475
rect 1075 475 1076 479
rect 1083 475 1084 479
rect 1158 477 1159 481
rect 1163 477 1164 481
rect 1238 481 1244 482
rect 1158 476 1164 477
rect 1178 479 1185 480
rect 1075 474 1084 475
rect 1178 475 1179 479
rect 1184 475 1185 479
rect 1238 477 1239 481
rect 1243 477 1244 481
rect 1238 476 1244 477
rect 1259 481 1265 482
rect 1259 477 1260 481
rect 1264 477 1265 481
rect 1259 476 1265 477
rect 1286 480 1292 481
rect 1286 476 1287 480
rect 1291 476 1292 480
rect 1372 480 1391 482
rect 1372 478 1374 480
rect 1390 479 1391 480
rect 1395 479 1396 483
rect 2070 483 2076 484
rect 2070 482 2071 483
rect 1390 478 1396 479
rect 1820 480 2071 482
rect 1820 478 1822 480
rect 2070 479 2071 480
rect 2075 479 2076 483
rect 2350 483 2356 484
rect 2350 482 2351 483
rect 2070 478 2076 479
rect 2144 480 2351 482
rect 1286 475 1292 476
rect 1371 477 1377 478
rect 1178 474 1185 475
rect 1371 473 1372 477
rect 1376 473 1377 477
rect 1819 477 1825 478
rect 1435 475 1441 476
rect 1435 474 1436 475
rect 1371 472 1377 473
rect 1389 472 1436 474
rect 110 463 116 464
rect 110 459 111 463
rect 115 459 116 463
rect 1286 463 1292 464
rect 110 458 116 459
rect 134 460 140 461
rect 134 456 135 460
rect 139 456 140 460
rect 134 455 140 456
rect 230 460 236 461
rect 230 456 231 460
rect 235 456 236 460
rect 230 455 236 456
rect 350 460 356 461
rect 350 456 351 460
rect 355 456 356 460
rect 350 455 356 456
rect 470 460 476 461
rect 470 456 471 460
rect 475 456 476 460
rect 470 455 476 456
rect 598 460 604 461
rect 598 456 599 460
rect 603 456 604 460
rect 598 455 604 456
rect 718 460 724 461
rect 718 456 719 460
rect 723 456 724 460
rect 718 455 724 456
rect 830 460 836 461
rect 830 456 831 460
rect 835 456 836 460
rect 830 455 836 456
rect 934 460 940 461
rect 934 456 935 460
rect 939 456 940 460
rect 934 455 940 456
rect 1038 460 1044 461
rect 1038 456 1039 460
rect 1043 456 1044 460
rect 1038 455 1044 456
rect 1142 460 1148 461
rect 1142 456 1143 460
rect 1147 456 1148 460
rect 1142 455 1148 456
rect 1222 460 1228 461
rect 1222 456 1223 460
rect 1227 456 1228 460
rect 1286 459 1287 463
rect 1291 459 1292 463
rect 1389 462 1391 472
rect 1435 471 1436 472
rect 1440 471 1441 475
rect 1523 475 1529 476
rect 1523 474 1524 475
rect 1435 470 1441 471
rect 1452 472 1524 474
rect 1452 462 1454 472
rect 1523 471 1524 472
rect 1528 471 1529 475
rect 1523 470 1529 471
rect 1550 475 1556 476
rect 1550 471 1551 475
rect 1555 474 1556 475
rect 1619 475 1625 476
rect 1619 474 1620 475
rect 1555 472 1620 474
rect 1555 471 1556 472
rect 1550 470 1556 471
rect 1619 471 1620 472
rect 1624 471 1625 475
rect 1715 475 1721 476
rect 1715 474 1716 475
rect 1619 470 1625 471
rect 1668 472 1716 474
rect 1668 466 1670 472
rect 1715 471 1716 472
rect 1720 471 1721 475
rect 1819 473 1820 477
rect 1824 473 1825 477
rect 1819 472 1825 473
rect 1931 475 1937 476
rect 1715 470 1721 471
rect 1931 471 1932 475
rect 1936 471 1937 475
rect 1931 470 1937 471
rect 2059 475 2065 476
rect 2059 471 2060 475
rect 2064 474 2065 475
rect 2144 474 2146 480
rect 2350 479 2351 480
rect 2355 479 2356 483
rect 2350 478 2356 479
rect 2064 472 2146 474
rect 2150 475 2156 476
rect 2064 471 2065 472
rect 2059 470 2065 471
rect 2150 471 2151 475
rect 2155 474 2156 475
rect 2195 475 2201 476
rect 2195 474 2196 475
rect 2155 472 2196 474
rect 2155 471 2156 472
rect 2150 470 2156 471
rect 2195 471 2196 472
rect 2200 471 2201 475
rect 2339 475 2345 476
rect 2339 474 2340 475
rect 2195 470 2201 471
rect 2212 472 2340 474
rect 1933 466 1935 470
rect 1636 464 1670 466
rect 1837 464 1935 466
rect 1636 462 1638 464
rect 1837 462 1839 464
rect 2212 462 2214 472
rect 2339 471 2340 472
rect 2344 471 2345 475
rect 2339 470 2345 471
rect 2459 475 2468 476
rect 2459 471 2460 475
rect 2467 471 2468 475
rect 2459 470 2468 471
rect 1366 461 1372 462
rect 1286 458 1292 459
rect 1326 460 1332 461
rect 1222 455 1228 456
rect 1326 456 1327 460
rect 1331 456 1332 460
rect 1366 457 1367 461
rect 1371 457 1372 461
rect 1366 456 1372 457
rect 1387 461 1393 462
rect 1387 457 1388 461
rect 1392 457 1393 461
rect 1387 456 1393 457
rect 1430 461 1436 462
rect 1430 457 1431 461
rect 1435 457 1436 461
rect 1430 456 1436 457
rect 1451 461 1457 462
rect 1451 457 1452 461
rect 1456 457 1457 461
rect 1451 456 1457 457
rect 1518 461 1524 462
rect 1518 457 1519 461
rect 1523 457 1524 461
rect 1614 461 1620 462
rect 1518 456 1524 457
rect 1526 459 1532 460
rect 1326 455 1332 456
rect 1526 455 1527 459
rect 1531 458 1532 459
rect 1539 459 1545 460
rect 1539 458 1540 459
rect 1531 456 1540 458
rect 1531 455 1532 456
rect 1526 454 1532 455
rect 1539 455 1540 456
rect 1544 455 1545 459
rect 1614 457 1615 461
rect 1619 457 1620 461
rect 1614 456 1620 457
rect 1635 461 1641 462
rect 1635 457 1636 461
rect 1640 457 1641 461
rect 1635 456 1641 457
rect 1710 461 1716 462
rect 1710 457 1711 461
rect 1715 457 1716 461
rect 1814 461 1820 462
rect 1710 456 1716 457
rect 1718 459 1724 460
rect 1539 454 1545 455
rect 1718 455 1719 459
rect 1723 458 1724 459
rect 1731 459 1737 460
rect 1731 458 1732 459
rect 1723 456 1732 458
rect 1723 455 1724 456
rect 1718 454 1724 455
rect 1731 455 1732 456
rect 1736 455 1737 459
rect 1814 457 1815 461
rect 1819 457 1820 461
rect 1814 456 1820 457
rect 1835 461 1841 462
rect 1835 457 1836 461
rect 1840 457 1841 461
rect 1835 456 1841 457
rect 1926 461 1932 462
rect 1926 457 1927 461
rect 1931 457 1932 461
rect 2054 461 2060 462
rect 1926 456 1932 457
rect 1947 459 1953 460
rect 1731 454 1737 455
rect 1947 455 1948 459
rect 1952 458 1953 459
rect 2022 459 2028 460
rect 2022 458 2023 459
rect 1952 456 2023 458
rect 1952 455 1953 456
rect 1947 454 1953 455
rect 2022 455 2023 456
rect 2027 455 2028 459
rect 2054 457 2055 461
rect 2059 457 2060 461
rect 2190 461 2196 462
rect 2054 456 2060 457
rect 2070 459 2081 460
rect 2022 454 2028 455
rect 2070 455 2071 459
rect 2075 455 2076 459
rect 2080 455 2081 459
rect 2190 457 2191 461
rect 2195 457 2196 461
rect 2190 456 2196 457
rect 2211 461 2217 462
rect 2211 457 2212 461
rect 2216 457 2217 461
rect 2211 456 2217 457
rect 2334 461 2340 462
rect 2334 457 2335 461
rect 2339 457 2340 461
rect 2454 461 2460 462
rect 2334 456 2340 457
rect 2350 459 2361 460
rect 2070 454 2081 455
rect 2350 455 2351 459
rect 2355 455 2356 459
rect 2360 455 2361 459
rect 2454 457 2455 461
rect 2459 457 2460 461
rect 2502 460 2508 461
rect 2454 456 2460 457
rect 2470 459 2481 460
rect 2350 454 2361 455
rect 2470 455 2471 459
rect 2475 455 2476 459
rect 2480 455 2481 459
rect 2502 456 2503 460
rect 2507 456 2508 460
rect 2502 455 2508 456
rect 2470 454 2481 455
rect 134 444 140 445
rect 110 441 116 442
rect 110 437 111 441
rect 115 437 116 441
rect 134 440 135 444
rect 139 440 140 444
rect 134 439 140 440
rect 190 444 196 445
rect 190 440 191 444
rect 195 440 196 444
rect 190 439 196 440
rect 246 444 252 445
rect 246 440 247 444
rect 251 440 252 444
rect 246 439 252 440
rect 302 444 308 445
rect 302 440 303 444
rect 307 440 308 444
rect 302 439 308 440
rect 382 444 388 445
rect 382 440 383 444
rect 387 440 388 444
rect 382 439 388 440
rect 470 444 476 445
rect 470 440 471 444
rect 475 440 476 444
rect 470 439 476 440
rect 566 444 572 445
rect 566 440 567 444
rect 571 440 572 444
rect 566 439 572 440
rect 670 444 676 445
rect 670 440 671 444
rect 675 440 676 444
rect 670 439 676 440
rect 782 444 788 445
rect 782 440 783 444
rect 787 440 788 444
rect 782 439 788 440
rect 894 444 900 445
rect 894 440 895 444
rect 899 440 900 444
rect 894 439 900 440
rect 1006 444 1012 445
rect 1006 440 1007 444
rect 1011 440 1012 444
rect 1006 439 1012 440
rect 1126 444 1132 445
rect 1126 440 1127 444
rect 1131 440 1132 444
rect 1126 439 1132 440
rect 1222 444 1228 445
rect 1222 440 1223 444
rect 1227 440 1228 444
rect 1326 443 1332 444
rect 1222 439 1228 440
rect 1286 441 1292 442
rect 110 436 116 437
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1326 439 1327 443
rect 1331 439 1332 443
rect 2502 443 2508 444
rect 1326 438 1332 439
rect 1350 440 1356 441
rect 1286 436 1292 437
rect 1350 436 1351 440
rect 1355 436 1356 440
rect 1350 435 1356 436
rect 1414 440 1420 441
rect 1414 436 1415 440
rect 1419 436 1420 440
rect 1414 435 1420 436
rect 1502 440 1508 441
rect 1502 436 1503 440
rect 1507 436 1508 440
rect 1502 435 1508 436
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1694 440 1700 441
rect 1694 436 1695 440
rect 1699 436 1700 440
rect 1694 435 1700 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1910 440 1916 441
rect 1910 436 1911 440
rect 1915 436 1916 440
rect 1910 435 1916 436
rect 2038 440 2044 441
rect 2038 436 2039 440
rect 2043 436 2044 440
rect 2038 435 2044 436
rect 2174 440 2180 441
rect 2174 436 2175 440
rect 2179 436 2180 440
rect 2174 435 2180 436
rect 2318 440 2324 441
rect 2318 436 2319 440
rect 2323 436 2324 440
rect 2318 435 2324 436
rect 2438 440 2444 441
rect 2438 436 2439 440
rect 2443 436 2444 440
rect 2502 439 2503 443
rect 2507 439 2508 443
rect 2502 438 2508 439
rect 2438 435 2444 436
rect 110 424 116 425
rect 1286 424 1292 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 150 423 156 424
rect 150 419 151 423
rect 155 419 156 423
rect 150 418 156 419
rect 171 423 177 424
rect 171 419 172 423
rect 176 419 177 423
rect 171 418 177 419
rect 206 423 212 424
rect 206 419 207 423
rect 211 419 212 423
rect 206 418 212 419
rect 214 423 220 424
rect 214 419 215 423
rect 219 422 220 423
rect 227 423 233 424
rect 227 422 228 423
rect 219 420 228 422
rect 219 419 220 420
rect 214 418 220 419
rect 227 419 228 420
rect 232 419 233 423
rect 227 418 233 419
rect 262 423 268 424
rect 262 419 263 423
rect 267 419 268 423
rect 262 418 268 419
rect 283 423 289 424
rect 283 419 284 423
rect 288 422 289 423
rect 318 423 324 424
rect 288 420 306 422
rect 288 419 289 420
rect 283 418 289 419
rect 173 410 175 418
rect 304 410 306 420
rect 318 419 319 423
rect 323 419 324 423
rect 318 418 324 419
rect 339 423 348 424
rect 339 419 340 423
rect 347 419 348 423
rect 339 418 348 419
rect 398 423 404 424
rect 398 419 399 423
rect 403 419 404 423
rect 398 418 404 419
rect 414 423 425 424
rect 414 419 415 423
rect 419 419 420 423
rect 424 419 425 423
rect 414 418 425 419
rect 486 423 492 424
rect 486 419 487 423
rect 491 419 492 423
rect 507 423 513 424
rect 507 422 508 423
rect 486 418 492 419
rect 496 420 508 422
rect 496 414 498 420
rect 507 419 508 420
rect 512 419 513 423
rect 507 418 513 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 603 423 609 424
rect 603 419 604 423
rect 608 422 609 423
rect 686 423 692 424
rect 608 420 682 422
rect 608 419 609 420
rect 603 418 609 419
rect 404 412 498 414
rect 404 410 406 412
rect 680 410 682 420
rect 686 419 687 423
rect 691 419 692 423
rect 686 418 692 419
rect 707 423 713 424
rect 707 419 708 423
rect 712 422 713 423
rect 798 423 804 424
rect 712 420 794 422
rect 712 419 713 420
rect 707 418 713 419
rect 792 410 794 420
rect 798 419 799 423
rect 803 419 804 423
rect 798 418 804 419
rect 819 423 825 424
rect 819 419 820 423
rect 824 422 825 423
rect 910 423 916 424
rect 824 420 906 422
rect 824 419 825 420
rect 819 418 825 419
rect 904 410 906 420
rect 910 419 911 423
rect 915 419 916 423
rect 910 418 916 419
rect 918 423 924 424
rect 918 419 919 423
rect 923 422 924 423
rect 931 423 937 424
rect 931 422 932 423
rect 923 420 932 422
rect 923 419 924 420
rect 918 418 924 419
rect 931 419 932 420
rect 936 419 937 423
rect 931 418 937 419
rect 1022 423 1028 424
rect 1022 419 1023 423
rect 1027 419 1028 423
rect 1022 418 1028 419
rect 1043 423 1049 424
rect 1043 419 1044 423
rect 1048 422 1049 423
rect 1142 423 1148 424
rect 1048 420 1138 422
rect 1048 419 1049 420
rect 1043 418 1049 419
rect 1136 410 1138 420
rect 1142 419 1143 423
rect 1147 419 1148 423
rect 1142 418 1148 419
rect 1163 423 1169 424
rect 1163 419 1164 423
rect 1168 422 1169 423
rect 1238 423 1244 424
rect 1168 420 1234 422
rect 1168 419 1169 420
rect 1163 418 1169 419
rect 1232 410 1234 420
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1238 418 1244 419
rect 1258 423 1265 424
rect 1258 419 1259 423
rect 1264 419 1265 423
rect 1286 420 1287 424
rect 1291 420 1292 424
rect 1350 424 1356 425
rect 1286 419 1292 420
rect 1326 421 1332 422
rect 1258 418 1265 419
rect 1326 417 1327 421
rect 1331 417 1332 421
rect 1350 420 1351 424
rect 1355 420 1356 424
rect 1350 419 1356 420
rect 1422 424 1428 425
rect 1422 420 1423 424
rect 1427 420 1428 424
rect 1422 419 1428 420
rect 1510 424 1516 425
rect 1510 420 1511 424
rect 1515 420 1516 424
rect 1510 419 1516 420
rect 1598 424 1604 425
rect 1598 420 1599 424
rect 1603 420 1604 424
rect 1598 419 1604 420
rect 1678 424 1684 425
rect 1678 420 1679 424
rect 1683 420 1684 424
rect 1678 419 1684 420
rect 1774 424 1780 425
rect 1774 420 1775 424
rect 1779 420 1780 424
rect 1774 419 1780 420
rect 1886 424 1892 425
rect 1886 420 1887 424
rect 1891 420 1892 424
rect 1886 419 1892 420
rect 2014 424 2020 425
rect 2014 420 2015 424
rect 2019 420 2020 424
rect 2014 419 2020 420
rect 2158 424 2164 425
rect 2158 420 2159 424
rect 2163 420 2164 424
rect 2158 419 2164 420
rect 2310 424 2316 425
rect 2310 420 2311 424
rect 2315 420 2316 424
rect 2310 419 2316 420
rect 2438 424 2444 425
rect 2438 420 2439 424
rect 2443 420 2444 424
rect 2438 419 2444 420
rect 2502 421 2508 422
rect 1326 416 1332 417
rect 2502 417 2503 421
rect 2507 417 2508 421
rect 2502 416 2508 417
rect 173 409 217 410
rect 173 408 212 409
rect 155 407 164 408
rect 155 403 156 407
rect 163 403 164 407
rect 211 405 212 408
rect 216 405 217 409
rect 304 409 329 410
rect 304 408 324 409
rect 211 404 217 405
rect 267 407 273 408
rect 155 402 164 403
rect 267 403 268 407
rect 272 406 273 407
rect 272 404 321 406
rect 323 405 324 408
rect 328 405 329 409
rect 323 404 329 405
rect 403 409 409 410
rect 403 405 404 409
rect 408 405 409 409
rect 680 409 697 410
rect 680 408 692 409
rect 403 404 409 405
rect 491 407 497 408
rect 272 403 273 404
rect 267 402 273 403
rect 319 402 321 404
rect 414 403 420 404
rect 414 402 415 403
rect 319 400 415 402
rect 414 399 415 400
rect 419 399 420 403
rect 491 403 492 407
rect 496 406 497 407
rect 530 407 536 408
rect 530 406 531 407
rect 496 404 531 406
rect 496 403 497 404
rect 491 402 497 403
rect 530 403 531 404
rect 535 403 536 407
rect 530 402 536 403
rect 587 407 593 408
rect 587 403 588 407
rect 592 406 593 407
rect 622 407 628 408
rect 622 406 623 407
rect 592 404 623 406
rect 592 403 593 404
rect 587 402 593 403
rect 622 403 623 404
rect 627 403 628 407
rect 691 405 692 408
rect 696 405 697 409
rect 792 409 809 410
rect 792 408 804 409
rect 691 404 697 405
rect 803 405 804 408
rect 808 405 809 409
rect 904 409 921 410
rect 904 408 916 409
rect 803 404 809 405
rect 915 405 916 408
rect 920 405 921 409
rect 1136 409 1153 410
rect 1136 408 1148 409
rect 915 404 921 405
rect 990 407 996 408
rect 622 402 628 403
rect 990 403 991 407
rect 995 406 996 407
rect 1027 407 1033 408
rect 1027 406 1028 407
rect 995 404 1028 406
rect 995 403 996 404
rect 990 402 996 403
rect 1027 403 1028 404
rect 1032 403 1033 407
rect 1147 405 1148 408
rect 1152 405 1153 409
rect 1232 409 1249 410
rect 1232 408 1244 409
rect 1147 404 1153 405
rect 1243 405 1244 408
rect 1248 405 1249 409
rect 1243 404 1249 405
rect 1326 404 1332 405
rect 2502 404 2508 405
rect 1027 402 1033 403
rect 1326 400 1327 404
rect 1331 400 1332 404
rect 1326 399 1332 400
rect 1366 403 1372 404
rect 1366 399 1367 403
rect 1371 399 1372 403
rect 414 398 420 399
rect 1366 398 1372 399
rect 1374 403 1380 404
rect 1374 399 1375 403
rect 1379 402 1380 403
rect 1387 403 1393 404
rect 1387 402 1388 403
rect 1379 400 1388 402
rect 1379 399 1380 400
rect 1374 398 1380 399
rect 1387 399 1388 400
rect 1392 399 1393 403
rect 1387 398 1393 399
rect 1438 403 1444 404
rect 1438 399 1439 403
rect 1443 399 1444 403
rect 1438 398 1444 399
rect 1459 403 1465 404
rect 1459 399 1460 403
rect 1464 399 1465 403
rect 1459 398 1465 399
rect 1526 403 1532 404
rect 1526 399 1527 403
rect 1531 399 1532 403
rect 1526 398 1532 399
rect 1547 403 1556 404
rect 1547 399 1548 403
rect 1555 399 1556 403
rect 1547 398 1556 399
rect 1614 403 1620 404
rect 1614 399 1615 403
rect 1619 399 1620 403
rect 1635 403 1641 404
rect 1635 402 1636 403
rect 1614 398 1620 399
rect 1624 400 1636 402
rect 1461 394 1463 398
rect 1624 394 1626 400
rect 1635 399 1636 400
rect 1640 399 1641 403
rect 1635 398 1641 399
rect 1694 403 1700 404
rect 1694 399 1695 403
rect 1699 399 1700 403
rect 1694 398 1700 399
rect 1715 403 1721 404
rect 1715 399 1716 403
rect 1720 402 1721 403
rect 1790 403 1796 404
rect 1720 400 1786 402
rect 1720 399 1721 400
rect 1715 398 1721 399
rect 1372 392 1463 394
rect 1532 392 1626 394
rect 1372 390 1374 392
rect 1532 390 1534 392
rect 1784 390 1786 400
rect 1790 399 1791 403
rect 1795 399 1796 403
rect 1790 398 1796 399
rect 1811 403 1820 404
rect 1811 399 1812 403
rect 1819 399 1820 403
rect 1811 398 1820 399
rect 1902 403 1908 404
rect 1902 399 1903 403
rect 1907 399 1908 403
rect 1902 398 1908 399
rect 1923 403 1929 404
rect 1923 399 1924 403
rect 1928 399 1929 403
rect 1923 398 1929 399
rect 2030 403 2036 404
rect 2030 399 2031 403
rect 2035 399 2036 403
rect 2030 398 2036 399
rect 2051 403 2057 404
rect 2051 399 2052 403
rect 2056 402 2057 403
rect 2174 403 2180 404
rect 2056 400 2170 402
rect 2056 399 2057 400
rect 2051 398 2057 399
rect 1925 394 1927 398
rect 1812 392 1927 394
rect 1371 389 1377 390
rect 298 387 304 388
rect 298 386 299 387
rect 156 384 299 386
rect 156 382 158 384
rect 298 383 299 384
rect 303 383 304 387
rect 478 387 484 388
rect 478 386 479 387
rect 298 382 304 383
rect 364 384 479 386
rect 364 382 366 384
rect 478 383 479 384
rect 483 383 484 387
rect 842 387 848 388
rect 842 386 843 387
rect 478 382 484 383
rect 756 384 843 386
rect 756 382 758 384
rect 842 383 843 384
rect 847 383 848 387
rect 1371 385 1372 389
rect 1376 385 1377 389
rect 1531 389 1537 390
rect 1371 384 1377 385
rect 1443 387 1449 388
rect 842 382 848 383
rect 1443 383 1444 387
rect 1448 386 1449 387
rect 1518 387 1524 388
rect 1518 386 1519 387
rect 1448 384 1519 386
rect 1448 383 1449 384
rect 1443 382 1449 383
rect 1518 383 1519 384
rect 1523 383 1524 387
rect 1531 385 1532 389
rect 1536 385 1537 389
rect 1784 389 1801 390
rect 1784 388 1796 389
rect 1531 384 1537 385
rect 1619 387 1625 388
rect 1518 382 1524 383
rect 1619 383 1620 387
rect 1624 386 1625 387
rect 1699 387 1705 388
rect 1624 384 1694 386
rect 1624 383 1625 384
rect 1619 382 1625 383
rect 155 381 161 382
rect 155 377 156 381
rect 160 377 161 381
rect 363 381 369 382
rect 155 376 161 377
rect 211 379 220 380
rect 211 375 212 379
rect 219 375 220 379
rect 283 379 289 380
rect 283 378 284 379
rect 211 374 220 375
rect 232 376 284 378
rect 232 370 234 376
rect 283 375 284 376
rect 288 375 289 379
rect 363 377 364 381
rect 368 377 369 381
rect 755 381 761 382
rect 435 379 441 380
rect 435 378 436 379
rect 363 376 369 377
rect 380 376 436 378
rect 283 374 289 375
rect 228 368 234 370
rect 228 366 230 368
rect 380 366 382 376
rect 435 375 436 376
rect 440 375 441 379
rect 515 379 521 380
rect 515 378 516 379
rect 435 374 441 375
rect 476 376 516 378
rect 476 370 478 376
rect 515 375 516 376
rect 520 375 521 379
rect 515 374 521 375
rect 595 379 601 380
rect 595 375 596 379
rect 600 378 601 379
rect 675 379 681 380
rect 600 376 670 378
rect 600 375 601 376
rect 595 374 601 375
rect 452 368 478 370
rect 668 370 670 376
rect 675 375 676 379
rect 680 378 681 379
rect 680 376 750 378
rect 755 377 756 381
rect 760 377 761 381
rect 755 376 761 377
rect 827 379 833 380
rect 680 375 681 376
rect 675 374 681 375
rect 748 370 750 376
rect 827 375 828 379
rect 832 375 833 379
rect 827 374 833 375
rect 899 379 905 380
rect 899 375 900 379
rect 904 378 905 379
rect 918 379 924 380
rect 918 378 919 379
rect 904 376 919 378
rect 904 375 905 376
rect 899 374 905 375
rect 918 375 919 376
rect 923 375 924 379
rect 918 374 924 375
rect 971 379 977 380
rect 971 375 972 379
rect 976 378 977 379
rect 1043 379 1049 380
rect 976 376 1038 378
rect 976 375 977 376
rect 971 374 977 375
rect 829 370 831 374
rect 1036 370 1038 376
rect 1043 375 1044 379
rect 1048 378 1049 379
rect 1070 379 1076 380
rect 1048 376 1066 378
rect 1048 375 1049 376
rect 1043 374 1049 375
rect 1064 370 1066 376
rect 1070 375 1071 379
rect 1075 378 1076 379
rect 1115 379 1121 380
rect 1115 378 1116 379
rect 1075 376 1116 378
rect 1075 375 1076 376
rect 1070 374 1076 375
rect 1115 375 1116 376
rect 1120 375 1121 379
rect 1115 374 1121 375
rect 1187 379 1193 380
rect 1187 375 1188 379
rect 1192 378 1193 379
rect 1243 379 1249 380
rect 1192 376 1238 378
rect 1192 375 1193 376
rect 1187 374 1193 375
rect 1236 370 1238 376
rect 1243 375 1244 379
rect 1248 378 1249 379
rect 1374 379 1380 380
rect 1374 378 1375 379
rect 1248 376 1375 378
rect 1248 375 1249 376
rect 1243 374 1249 375
rect 1374 375 1375 376
rect 1379 375 1380 379
rect 1692 378 1694 384
rect 1699 383 1700 387
rect 1704 386 1705 387
rect 1704 384 1790 386
rect 1795 385 1796 388
rect 1800 385 1801 389
rect 1795 384 1801 385
rect 1704 383 1705 384
rect 1699 382 1705 383
rect 1788 382 1790 384
rect 1812 382 1814 392
rect 2168 390 2170 400
rect 2174 399 2175 403
rect 2179 399 2180 403
rect 2174 398 2180 399
rect 2195 403 2201 404
rect 2195 399 2196 403
rect 2200 399 2201 403
rect 2195 398 2201 399
rect 2326 403 2332 404
rect 2326 399 2327 403
rect 2331 399 2332 403
rect 2326 398 2332 399
rect 2334 403 2340 404
rect 2334 399 2335 403
rect 2339 402 2340 403
rect 2347 403 2353 404
rect 2347 402 2348 403
rect 2339 400 2348 402
rect 2339 399 2340 400
rect 2334 398 2340 399
rect 2347 399 2348 400
rect 2352 399 2353 403
rect 2347 398 2353 399
rect 2454 403 2460 404
rect 2454 399 2455 403
rect 2459 399 2460 403
rect 2454 398 2460 399
rect 2462 403 2468 404
rect 2462 399 2463 403
rect 2467 402 2468 403
rect 2475 403 2481 404
rect 2475 402 2476 403
rect 2467 400 2476 402
rect 2467 399 2468 400
rect 2462 398 2468 399
rect 2475 399 2476 400
rect 2480 399 2481 403
rect 2502 400 2503 404
rect 2507 400 2508 404
rect 2502 399 2508 400
rect 2475 398 2481 399
rect 2197 390 2199 398
rect 2168 389 2185 390
rect 2168 388 2180 389
rect 1907 387 1913 388
rect 1907 383 1908 387
rect 1912 386 1913 387
rect 2022 387 2028 388
rect 1912 384 2001 386
rect 1912 383 1913 384
rect 1907 382 1913 383
rect 1788 380 1814 382
rect 1754 379 1760 380
rect 1754 378 1755 379
rect 1692 376 1755 378
rect 1374 374 1380 375
rect 1754 375 1755 376
rect 1759 375 1760 379
rect 1999 378 2001 384
rect 2022 383 2023 387
rect 2027 386 2028 387
rect 2035 387 2041 388
rect 2035 386 2036 387
rect 2027 384 2036 386
rect 2027 383 2028 384
rect 2022 382 2028 383
rect 2035 383 2036 384
rect 2040 383 2041 387
rect 2179 385 2180 388
rect 2184 385 2185 389
rect 2197 389 2337 390
rect 2197 388 2332 389
rect 2179 384 2185 385
rect 2331 385 2332 388
rect 2336 385 2337 389
rect 2331 384 2337 385
rect 2459 387 2465 388
rect 2035 382 2041 383
rect 2459 383 2460 387
rect 2464 386 2465 387
rect 2470 387 2476 388
rect 2470 386 2471 387
rect 2464 384 2471 386
rect 2464 383 2465 384
rect 2459 382 2465 383
rect 2470 383 2471 384
rect 2475 383 2476 387
rect 2470 382 2476 383
rect 2334 379 2340 380
rect 2334 378 2335 379
rect 1999 376 2335 378
rect 1754 374 1760 375
rect 2334 375 2335 376
rect 2339 375 2340 379
rect 2334 374 2340 375
rect 668 368 694 370
rect 748 368 774 370
rect 829 368 918 370
rect 1036 368 1062 370
rect 1064 368 1135 370
rect 1236 368 1262 370
rect 452 366 454 368
rect 692 366 694 368
rect 772 366 774 368
rect 916 366 918 368
rect 1060 366 1062 368
rect 1133 366 1135 368
rect 1260 366 1262 368
rect 150 365 156 366
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 150 361 151 365
rect 155 361 156 365
rect 206 365 212 366
rect 150 360 156 361
rect 158 363 164 364
rect 110 359 116 360
rect 158 359 159 363
rect 163 362 164 363
rect 171 363 177 364
rect 171 362 172 363
rect 163 360 172 362
rect 163 359 164 360
rect 158 358 164 359
rect 171 359 172 360
rect 176 359 177 363
rect 206 361 207 365
rect 211 361 212 365
rect 206 360 212 361
rect 227 365 233 366
rect 227 361 228 365
rect 232 361 233 365
rect 227 360 233 361
rect 278 365 284 366
rect 278 361 279 365
rect 283 361 284 365
rect 358 365 364 366
rect 278 360 284 361
rect 298 363 305 364
rect 171 358 177 359
rect 298 359 299 363
rect 304 359 305 363
rect 358 361 359 365
rect 363 361 364 365
rect 358 360 364 361
rect 379 365 385 366
rect 379 361 380 365
rect 384 361 385 365
rect 379 360 385 361
rect 430 365 436 366
rect 430 361 431 365
rect 435 361 436 365
rect 430 360 436 361
rect 451 365 457 366
rect 451 361 452 365
rect 456 361 457 365
rect 451 360 457 361
rect 510 365 516 366
rect 510 361 511 365
rect 515 361 516 365
rect 590 365 596 366
rect 510 360 516 361
rect 530 363 537 364
rect 298 358 305 359
rect 530 359 531 363
rect 536 359 537 363
rect 590 361 591 365
rect 595 361 596 365
rect 670 365 676 366
rect 590 360 596 361
rect 611 363 617 364
rect 530 358 537 359
rect 611 359 612 363
rect 616 362 617 363
rect 638 363 644 364
rect 638 362 639 363
rect 616 360 639 362
rect 616 359 617 360
rect 611 358 617 359
rect 638 359 639 360
rect 643 359 644 363
rect 670 361 671 365
rect 675 361 676 365
rect 670 360 676 361
rect 691 365 697 366
rect 691 361 692 365
rect 696 361 697 365
rect 691 360 697 361
rect 750 365 756 366
rect 750 361 751 365
rect 755 361 756 365
rect 750 360 756 361
rect 771 365 777 366
rect 771 361 772 365
rect 776 361 777 365
rect 771 360 777 361
rect 822 365 828 366
rect 822 361 823 365
rect 827 361 828 365
rect 894 365 900 366
rect 822 360 828 361
rect 842 363 849 364
rect 638 358 644 359
rect 842 359 843 363
rect 848 359 849 363
rect 894 361 895 365
rect 899 361 900 365
rect 894 360 900 361
rect 915 365 921 366
rect 915 361 916 365
rect 920 361 921 365
rect 915 360 921 361
rect 966 365 972 366
rect 966 361 967 365
rect 971 361 972 365
rect 1038 365 1044 366
rect 966 360 972 361
rect 987 363 996 364
rect 842 358 849 359
rect 987 359 988 363
rect 995 359 996 363
rect 1038 361 1039 365
rect 1043 361 1044 365
rect 1038 360 1044 361
rect 1059 365 1065 366
rect 1059 361 1060 365
rect 1064 361 1065 365
rect 1059 360 1065 361
rect 1110 365 1116 366
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 1131 365 1137 366
rect 1131 361 1132 365
rect 1136 361 1137 365
rect 1131 360 1137 361
rect 1182 365 1188 366
rect 1182 361 1183 365
rect 1187 361 1188 365
rect 1238 365 1244 366
rect 1182 360 1188 361
rect 1203 363 1209 364
rect 987 358 996 359
rect 1203 359 1204 363
rect 1208 362 1209 363
rect 1230 363 1236 364
rect 1230 362 1231 363
rect 1208 360 1231 362
rect 1208 359 1209 360
rect 1203 358 1209 359
rect 1230 359 1231 360
rect 1235 359 1236 363
rect 1238 361 1239 365
rect 1243 361 1244 365
rect 1238 360 1244 361
rect 1259 365 1265 366
rect 1259 361 1260 365
rect 1264 361 1265 365
rect 1259 360 1265 361
rect 1286 364 1292 365
rect 1286 360 1287 364
rect 1291 360 1292 364
rect 1286 359 1292 360
rect 1670 363 1676 364
rect 1670 359 1671 363
rect 1675 362 1676 363
rect 1683 363 1689 364
rect 1683 362 1684 363
rect 1675 360 1684 362
rect 1675 359 1676 360
rect 1230 358 1236 359
rect 1670 358 1676 359
rect 1683 359 1684 360
rect 1688 359 1689 363
rect 1739 363 1745 364
rect 1739 362 1740 363
rect 1683 358 1689 359
rect 1716 360 1740 362
rect 1716 354 1718 360
rect 1739 359 1740 360
rect 1744 359 1745 363
rect 1739 358 1745 359
rect 1811 363 1820 364
rect 1811 359 1812 363
rect 1819 359 1820 363
rect 1907 363 1913 364
rect 1907 362 1908 363
rect 1811 358 1820 359
rect 1828 360 1908 362
rect 1700 352 1718 354
rect 1700 350 1702 352
rect 1828 350 1830 360
rect 1907 359 1908 360
rect 1912 359 1913 363
rect 2027 363 2033 364
rect 2027 362 2028 363
rect 1907 358 1913 359
rect 1999 360 2028 362
rect 1999 350 2001 360
rect 2027 359 2028 360
rect 2032 359 2033 363
rect 2163 363 2169 364
rect 2163 362 2164 363
rect 2027 358 2033 359
rect 2048 360 2164 362
rect 2048 350 2050 360
rect 2163 359 2164 360
rect 2168 359 2169 363
rect 2307 363 2313 364
rect 2307 362 2308 363
rect 2163 358 2169 359
rect 2180 360 2308 362
rect 2180 350 2182 360
rect 2307 359 2308 360
rect 2312 359 2313 363
rect 2307 358 2313 359
rect 2459 363 2468 364
rect 2459 359 2460 363
rect 2467 359 2468 363
rect 2459 358 2468 359
rect 1678 349 1684 350
rect 1326 348 1332 349
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 1286 347 1292 348
rect 110 342 116 343
rect 134 344 140 345
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 190 344 196 345
rect 190 340 191 344
rect 195 340 196 344
rect 190 339 196 340
rect 262 344 268 345
rect 262 340 263 344
rect 267 340 268 344
rect 262 339 268 340
rect 342 344 348 345
rect 342 340 343 344
rect 347 340 348 344
rect 342 339 348 340
rect 414 344 420 345
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 806 344 812 345
rect 806 340 807 344
rect 811 340 812 344
rect 806 339 812 340
rect 878 344 884 345
rect 878 340 879 344
rect 883 340 884 344
rect 878 339 884 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1022 344 1028 345
rect 1022 340 1023 344
rect 1027 340 1028 344
rect 1022 339 1028 340
rect 1094 344 1100 345
rect 1094 340 1095 344
rect 1099 340 1100 344
rect 1094 339 1100 340
rect 1166 344 1172 345
rect 1166 340 1167 344
rect 1171 340 1172 344
rect 1166 339 1172 340
rect 1222 344 1228 345
rect 1222 340 1223 344
rect 1227 340 1228 344
rect 1286 343 1287 347
rect 1291 343 1292 347
rect 1326 344 1327 348
rect 1331 344 1332 348
rect 1678 345 1679 349
rect 1683 345 1684 349
rect 1678 344 1684 345
rect 1699 349 1705 350
rect 1699 345 1700 349
rect 1704 345 1705 349
rect 1699 344 1705 345
rect 1734 349 1740 350
rect 1734 345 1735 349
rect 1739 345 1740 349
rect 1806 349 1812 350
rect 1734 344 1740 345
rect 1754 347 1761 348
rect 1326 343 1332 344
rect 1754 343 1755 347
rect 1760 343 1761 347
rect 1806 345 1807 349
rect 1811 345 1812 349
rect 1806 344 1812 345
rect 1827 349 1833 350
rect 1827 345 1828 349
rect 1832 345 1833 349
rect 1827 344 1833 345
rect 1902 349 1908 350
rect 1902 345 1903 349
rect 1907 345 1908 349
rect 1902 344 1908 345
rect 1923 349 2001 350
rect 1923 345 1924 349
rect 1928 348 2001 349
rect 2022 349 2028 350
rect 1928 345 1929 348
rect 1923 344 1929 345
rect 2022 345 2023 349
rect 2027 345 2028 349
rect 2022 344 2028 345
rect 2043 349 2050 350
rect 2043 345 2044 349
rect 2048 348 2050 349
rect 2158 349 2164 350
rect 2048 345 2049 348
rect 2043 344 2049 345
rect 2158 345 2159 349
rect 2163 345 2164 349
rect 2158 344 2164 345
rect 2179 349 2185 350
rect 2179 345 2180 349
rect 2184 345 2185 349
rect 2179 344 2185 345
rect 2302 349 2308 350
rect 2302 345 2303 349
rect 2307 345 2308 349
rect 2454 349 2460 350
rect 2302 344 2308 345
rect 2318 347 2329 348
rect 1286 342 1292 343
rect 1754 342 1761 343
rect 2318 343 2319 347
rect 2323 343 2324 347
rect 2328 343 2329 347
rect 2454 345 2455 349
rect 2459 345 2460 349
rect 2502 348 2508 349
rect 2454 344 2460 345
rect 2475 347 2484 348
rect 2318 342 2329 343
rect 2475 343 2476 347
rect 2483 343 2484 347
rect 2502 344 2503 348
rect 2507 344 2508 348
rect 2502 343 2508 344
rect 2475 342 2484 343
rect 1222 339 1228 340
rect 1326 331 1332 332
rect 1326 327 1327 331
rect 1331 327 1332 331
rect 2502 331 2508 332
rect 1326 326 1332 327
rect 1662 328 1668 329
rect 134 324 140 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 134 320 135 324
rect 139 320 140 324
rect 134 319 140 320
rect 198 324 204 325
rect 198 320 199 324
rect 203 320 204 324
rect 198 319 204 320
rect 286 324 292 325
rect 286 320 287 324
rect 291 320 292 324
rect 286 319 292 320
rect 374 324 380 325
rect 374 320 375 324
rect 379 320 380 324
rect 374 319 380 320
rect 454 324 460 325
rect 454 320 455 324
rect 459 320 460 324
rect 454 319 460 320
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 630 324 636 325
rect 630 320 631 324
rect 635 320 636 324
rect 630 319 636 320
rect 726 324 732 325
rect 726 320 727 324
rect 731 320 732 324
rect 726 319 732 320
rect 822 324 828 325
rect 822 320 823 324
rect 827 320 828 324
rect 822 319 828 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 1030 324 1036 325
rect 1030 320 1031 324
rect 1035 320 1036 324
rect 1030 319 1036 320
rect 1134 324 1140 325
rect 1134 320 1135 324
rect 1139 320 1140 324
rect 1134 319 1140 320
rect 1222 324 1228 325
rect 1222 320 1223 324
rect 1227 320 1228 324
rect 1662 324 1663 328
rect 1667 324 1668 328
rect 1662 323 1668 324
rect 1718 328 1724 329
rect 1718 324 1719 328
rect 1723 324 1724 328
rect 1718 323 1724 324
rect 1790 328 1796 329
rect 1790 324 1791 328
rect 1795 324 1796 328
rect 1790 323 1796 324
rect 1886 328 1892 329
rect 1886 324 1887 328
rect 1891 324 1892 328
rect 1886 323 1892 324
rect 2006 328 2012 329
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 2142 328 2148 329
rect 2142 324 2143 328
rect 2147 324 2148 328
rect 2142 323 2148 324
rect 2286 328 2292 329
rect 2286 324 2287 328
rect 2291 324 2292 328
rect 2286 323 2292 324
rect 2438 328 2444 329
rect 2438 324 2439 328
rect 2443 324 2444 328
rect 2502 327 2503 331
rect 2507 327 2508 331
rect 2502 326 2508 327
rect 2438 323 2444 324
rect 1222 319 1228 320
rect 1286 321 1292 322
rect 110 316 116 317
rect 1286 317 1287 321
rect 1291 317 1292 321
rect 1286 316 1292 317
rect 1350 316 1356 317
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1350 312 1351 316
rect 1355 312 1356 316
rect 1350 311 1356 312
rect 1430 316 1436 317
rect 1430 312 1431 316
rect 1435 312 1436 316
rect 1430 311 1436 312
rect 1526 316 1532 317
rect 1526 312 1527 316
rect 1531 312 1532 316
rect 1526 311 1532 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1710 316 1716 317
rect 1710 312 1711 316
rect 1715 312 1716 316
rect 1710 311 1716 312
rect 1806 316 1812 317
rect 1806 312 1807 316
rect 1811 312 1812 316
rect 1806 311 1812 312
rect 1910 316 1916 317
rect 1910 312 1911 316
rect 1915 312 1916 316
rect 1910 311 1916 312
rect 2022 316 2028 317
rect 2022 312 2023 316
rect 2027 312 2028 316
rect 2022 311 2028 312
rect 2150 316 2156 317
rect 2150 312 2151 316
rect 2155 312 2156 316
rect 2150 311 2156 312
rect 2286 316 2292 317
rect 2286 312 2287 316
rect 2291 312 2292 316
rect 2286 311 2292 312
rect 2422 316 2428 317
rect 2422 312 2423 316
rect 2427 312 2428 316
rect 2422 311 2428 312
rect 2502 313 2508 314
rect 1326 308 1332 309
rect 2502 309 2503 313
rect 2507 309 2508 313
rect 2502 308 2508 309
rect 110 304 116 305
rect 1286 304 1292 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 150 303 156 304
rect 150 299 151 303
rect 155 299 156 303
rect 150 298 156 299
rect 171 303 177 304
rect 171 299 172 303
rect 176 299 177 303
rect 171 298 177 299
rect 214 303 220 304
rect 214 299 215 303
rect 219 299 220 303
rect 214 298 220 299
rect 235 303 241 304
rect 235 299 236 303
rect 240 299 241 303
rect 235 298 241 299
rect 302 303 308 304
rect 302 299 303 303
rect 307 299 308 303
rect 302 298 308 299
rect 323 303 329 304
rect 323 299 324 303
rect 328 302 329 303
rect 334 303 340 304
rect 334 302 335 303
rect 328 300 335 302
rect 328 299 329 300
rect 323 298 329 299
rect 334 299 335 300
rect 339 299 340 303
rect 334 298 340 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 411 303 417 304
rect 411 299 412 303
rect 416 302 417 303
rect 470 303 476 304
rect 416 300 466 302
rect 416 299 417 300
rect 411 298 417 299
rect 173 290 175 298
rect 237 290 239 298
rect 464 290 466 300
rect 470 299 471 303
rect 475 299 476 303
rect 470 298 476 299
rect 478 303 484 304
rect 478 299 479 303
rect 483 302 484 303
rect 491 303 497 304
rect 491 302 492 303
rect 483 300 492 302
rect 483 299 484 300
rect 478 298 484 299
rect 491 299 492 300
rect 496 299 497 303
rect 491 298 497 299
rect 558 303 564 304
rect 558 299 559 303
rect 563 299 564 303
rect 579 303 585 304
rect 579 302 580 303
rect 558 298 564 299
rect 568 300 580 302
rect 568 294 570 300
rect 579 299 580 300
rect 584 299 585 303
rect 579 298 585 299
rect 646 303 652 304
rect 646 299 647 303
rect 651 299 652 303
rect 646 298 652 299
rect 667 303 673 304
rect 667 299 668 303
rect 672 302 673 303
rect 742 303 748 304
rect 672 300 738 302
rect 672 299 673 300
rect 667 298 673 299
rect 484 292 570 294
rect 173 289 225 290
rect 173 288 220 289
rect 155 287 164 288
rect 155 283 156 287
rect 163 283 164 287
rect 219 285 220 288
rect 224 285 225 289
rect 237 289 313 290
rect 237 288 308 289
rect 219 284 225 285
rect 307 285 308 288
rect 312 285 313 289
rect 464 289 481 290
rect 464 288 476 289
rect 307 284 313 285
rect 395 287 401 288
rect 155 282 164 283
rect 395 283 396 287
rect 400 286 401 287
rect 400 284 470 286
rect 475 285 476 288
rect 480 285 481 289
rect 475 284 481 285
rect 400 283 401 284
rect 395 282 401 283
rect 468 282 470 284
rect 484 282 486 292
rect 736 290 738 300
rect 742 299 743 303
rect 747 299 748 303
rect 742 298 748 299
rect 763 303 769 304
rect 763 299 764 303
rect 768 302 769 303
rect 838 303 844 304
rect 768 300 834 302
rect 768 299 769 300
rect 763 298 769 299
rect 832 290 834 300
rect 838 299 839 303
rect 843 299 844 303
rect 838 298 844 299
rect 859 303 865 304
rect 859 299 860 303
rect 864 302 865 303
rect 942 303 948 304
rect 864 300 934 302
rect 864 299 865 300
rect 859 298 865 299
rect 932 290 934 300
rect 942 299 943 303
rect 947 299 948 303
rect 942 298 948 299
rect 950 303 956 304
rect 950 299 951 303
rect 955 302 956 303
rect 963 303 969 304
rect 963 302 964 303
rect 955 300 964 302
rect 955 299 956 300
rect 950 298 956 299
rect 963 299 964 300
rect 968 299 969 303
rect 963 298 969 299
rect 1046 303 1052 304
rect 1046 299 1047 303
rect 1051 299 1052 303
rect 1046 298 1052 299
rect 1067 303 1076 304
rect 1067 299 1068 303
rect 1075 299 1076 303
rect 1067 298 1076 299
rect 1150 303 1156 304
rect 1150 299 1151 303
rect 1155 299 1156 303
rect 1171 303 1177 304
rect 1171 302 1172 303
rect 1150 298 1156 299
rect 1159 300 1172 302
rect 1159 294 1161 300
rect 1171 299 1172 300
rect 1176 299 1177 303
rect 1171 298 1177 299
rect 1238 303 1244 304
rect 1238 299 1239 303
rect 1243 299 1244 303
rect 1238 298 1244 299
rect 1259 303 1265 304
rect 1259 299 1260 303
rect 1264 302 1265 303
rect 1278 303 1284 304
rect 1278 302 1279 303
rect 1264 300 1279 302
rect 1264 299 1265 300
rect 1259 298 1265 299
rect 1278 299 1279 300
rect 1283 299 1284 303
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1278 298 1284 299
rect 1052 292 1161 294
rect 1326 296 1332 297
rect 2502 296 2508 297
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1052 290 1054 292
rect 1326 291 1332 292
rect 1366 295 1372 296
rect 1366 291 1367 295
rect 1371 291 1372 295
rect 1366 290 1372 291
rect 1387 295 1393 296
rect 1387 291 1388 295
rect 1392 291 1393 295
rect 1387 290 1393 291
rect 1446 295 1452 296
rect 1446 291 1447 295
rect 1451 291 1452 295
rect 1446 290 1452 291
rect 1467 295 1473 296
rect 1467 291 1468 295
rect 1472 294 1473 295
rect 1542 295 1548 296
rect 1472 292 1538 294
rect 1472 291 1473 292
rect 1467 290 1473 291
rect 736 289 753 290
rect 736 288 748 289
rect 542 287 548 288
rect 542 283 543 287
rect 547 286 548 287
rect 563 287 569 288
rect 563 286 564 287
rect 547 284 564 286
rect 547 283 548 284
rect 542 282 548 283
rect 563 283 564 284
rect 568 283 569 287
rect 563 282 569 283
rect 638 287 644 288
rect 638 283 639 287
rect 643 286 644 287
rect 651 287 657 288
rect 651 286 652 287
rect 643 284 652 286
rect 643 283 644 284
rect 638 282 644 283
rect 651 283 652 284
rect 656 283 657 287
rect 747 285 748 288
rect 752 285 753 289
rect 832 289 849 290
rect 832 288 844 289
rect 747 284 753 285
rect 843 285 844 288
rect 848 285 849 289
rect 932 289 953 290
rect 932 288 948 289
rect 843 284 849 285
rect 947 285 948 288
rect 952 285 953 289
rect 947 284 953 285
rect 1051 289 1057 290
rect 1051 285 1052 289
rect 1056 285 1057 289
rect 1051 284 1057 285
rect 1155 287 1161 288
rect 651 282 657 283
rect 1155 283 1156 287
rect 1160 286 1161 287
rect 1222 287 1228 288
rect 1222 286 1223 287
rect 1160 284 1223 286
rect 1160 283 1161 284
rect 1155 282 1161 283
rect 1222 283 1223 284
rect 1227 283 1228 287
rect 1222 282 1228 283
rect 1230 287 1236 288
rect 1230 283 1231 287
rect 1235 286 1236 287
rect 1243 287 1249 288
rect 1243 286 1244 287
rect 1235 284 1244 286
rect 1235 283 1236 284
rect 1230 282 1236 283
rect 1243 283 1244 284
rect 1248 283 1249 287
rect 1243 282 1249 283
rect 1389 282 1391 290
rect 1536 282 1538 292
rect 1542 291 1543 295
rect 1547 291 1548 295
rect 1542 290 1548 291
rect 1550 295 1556 296
rect 1550 291 1551 295
rect 1555 294 1556 295
rect 1563 295 1569 296
rect 1563 294 1564 295
rect 1555 292 1564 294
rect 1555 291 1556 292
rect 1550 290 1556 291
rect 1563 291 1564 292
rect 1568 291 1569 295
rect 1563 290 1569 291
rect 1638 295 1644 296
rect 1638 291 1639 295
rect 1643 291 1644 295
rect 1638 290 1644 291
rect 1659 295 1665 296
rect 1659 291 1660 295
rect 1664 294 1665 295
rect 1670 295 1676 296
rect 1670 294 1671 295
rect 1664 292 1671 294
rect 1664 291 1665 292
rect 1659 290 1665 291
rect 1670 291 1671 292
rect 1675 291 1676 295
rect 1670 290 1676 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1747 295 1753 296
rect 1747 291 1748 295
rect 1752 291 1753 295
rect 1747 290 1753 291
rect 1822 295 1828 296
rect 1822 291 1823 295
rect 1827 291 1828 295
rect 1822 290 1828 291
rect 1843 295 1849 296
rect 1843 291 1844 295
rect 1848 291 1849 295
rect 1843 290 1849 291
rect 1926 295 1932 296
rect 1926 291 1927 295
rect 1931 291 1932 295
rect 1926 290 1932 291
rect 1947 295 1953 296
rect 1947 291 1948 295
rect 1952 294 1953 295
rect 2038 295 2044 296
rect 1952 292 2001 294
rect 1952 291 1953 292
rect 1947 290 1953 291
rect 1749 286 1751 290
rect 1644 284 1751 286
rect 1845 286 1847 290
rect 1845 284 1935 286
rect 1644 282 1646 284
rect 1933 282 1935 284
rect 1999 282 2001 292
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2059 295 2065 296
rect 2059 291 2060 295
rect 2064 294 2065 295
rect 2166 295 2172 296
rect 2064 292 2158 294
rect 2064 291 2065 292
rect 2059 290 2065 291
rect 2156 282 2158 292
rect 2166 291 2167 295
rect 2171 291 2172 295
rect 2166 290 2172 291
rect 2187 295 2193 296
rect 2187 291 2188 295
rect 2192 294 2193 295
rect 2302 295 2308 296
rect 2192 292 2294 294
rect 2192 291 2193 292
rect 2187 290 2193 291
rect 2292 282 2294 292
rect 2302 291 2303 295
rect 2307 291 2308 295
rect 2302 290 2308 291
rect 2310 295 2316 296
rect 2310 291 2311 295
rect 2315 294 2316 295
rect 2323 295 2329 296
rect 2323 294 2324 295
rect 2315 292 2324 294
rect 2315 291 2316 292
rect 2310 290 2316 291
rect 2323 291 2324 292
rect 2328 291 2329 295
rect 2323 290 2329 291
rect 2438 295 2444 296
rect 2438 291 2439 295
rect 2443 291 2444 295
rect 2438 290 2444 291
rect 2459 295 2468 296
rect 2459 291 2460 295
rect 2467 291 2468 295
rect 2502 292 2503 296
rect 2507 292 2508 296
rect 2502 291 2508 292
rect 2459 290 2468 291
rect 468 280 486 282
rect 1389 281 1457 282
rect 1389 280 1452 281
rect 1278 279 1284 280
rect 1278 275 1279 279
rect 1283 278 1284 279
rect 1371 279 1377 280
rect 1371 278 1372 279
rect 1283 276 1372 278
rect 1283 275 1284 276
rect 1278 274 1284 275
rect 1371 275 1372 276
rect 1376 275 1377 279
rect 1451 277 1452 280
rect 1456 277 1457 281
rect 1536 281 1553 282
rect 1536 280 1548 281
rect 1451 276 1457 277
rect 1547 277 1548 280
rect 1552 277 1553 281
rect 1547 276 1553 277
rect 1643 281 1649 282
rect 1643 277 1644 281
rect 1648 277 1649 281
rect 1931 281 1937 282
rect 1643 276 1649 277
rect 1731 279 1737 280
rect 1371 274 1377 275
rect 1731 275 1732 279
rect 1736 278 1737 279
rect 1806 279 1812 280
rect 1806 278 1807 279
rect 1736 276 1807 278
rect 1736 275 1737 276
rect 1731 274 1737 275
rect 1806 275 1807 276
rect 1811 275 1812 279
rect 1806 274 1812 275
rect 1827 279 1833 280
rect 1827 275 1828 279
rect 1832 278 1833 279
rect 1832 276 1918 278
rect 1931 277 1932 281
rect 1936 277 1937 281
rect 1999 281 2049 282
rect 1999 280 2044 281
rect 1931 276 1937 277
rect 2043 277 2044 280
rect 2048 277 2049 281
rect 2156 281 2177 282
rect 2156 280 2172 281
rect 2043 276 2049 277
rect 2171 277 2172 280
rect 2176 277 2177 281
rect 2292 281 2313 282
rect 2292 280 2308 281
rect 2171 276 2177 277
rect 2307 277 2308 280
rect 2312 277 2313 281
rect 2307 276 2313 277
rect 2414 279 2420 280
rect 1832 275 1833 276
rect 1827 274 1833 275
rect 1916 274 1918 276
rect 2318 275 2324 276
rect 2318 274 2319 275
rect 1916 272 2319 274
rect 2318 271 2319 272
rect 2323 271 2324 275
rect 2414 275 2415 279
rect 2419 278 2420 279
rect 2443 279 2449 280
rect 2443 278 2444 279
rect 2419 276 2444 278
rect 2419 275 2420 276
rect 2414 274 2420 275
rect 2443 275 2444 276
rect 2448 275 2449 279
rect 2443 274 2449 275
rect 2318 270 2324 271
rect 346 267 352 268
rect 346 266 347 267
rect 156 264 347 266
rect 156 262 158 264
rect 346 263 347 264
rect 351 263 352 267
rect 634 267 640 268
rect 634 266 635 267
rect 346 262 352 263
rect 428 264 635 266
rect 428 262 430 264
rect 634 263 635 264
rect 639 263 640 267
rect 922 267 928 268
rect 922 266 923 267
rect 634 262 640 263
rect 716 264 923 266
rect 716 262 718 264
rect 922 263 923 264
rect 927 263 928 267
rect 922 262 928 263
rect 1550 263 1556 264
rect 1550 262 1551 263
rect 155 261 161 262
rect 155 257 156 261
rect 160 257 161 261
rect 427 261 433 262
rect 155 256 161 257
rect 235 259 241 260
rect 235 255 236 259
rect 240 255 241 259
rect 235 254 241 255
rect 331 259 340 260
rect 331 255 332 259
rect 339 255 340 259
rect 427 257 428 261
rect 432 257 433 261
rect 715 261 721 262
rect 523 259 529 260
rect 523 258 524 259
rect 427 256 433 257
rect 444 256 524 258
rect 331 254 340 255
rect 237 250 239 254
rect 172 248 239 250
rect 172 246 174 248
rect 444 246 446 256
rect 523 255 524 256
rect 528 255 529 259
rect 523 254 529 255
rect 619 259 625 260
rect 619 255 620 259
rect 624 258 625 259
rect 642 259 648 260
rect 642 258 643 259
rect 624 256 643 258
rect 624 255 625 256
rect 619 254 625 255
rect 642 255 643 256
rect 647 255 648 259
rect 715 257 716 261
rect 720 257 721 261
rect 1372 260 1551 262
rect 811 259 817 260
rect 811 258 812 259
rect 715 256 721 257
rect 776 256 812 258
rect 642 254 648 255
rect 776 250 778 256
rect 811 255 812 256
rect 816 255 817 259
rect 811 254 817 255
rect 907 259 913 260
rect 907 255 908 259
rect 912 258 913 259
rect 950 259 956 260
rect 950 258 951 259
rect 912 256 951 258
rect 912 255 913 256
rect 907 254 913 255
rect 950 255 951 256
rect 955 255 956 259
rect 950 254 956 255
rect 998 259 1004 260
rect 998 255 999 259
rect 1003 258 1004 259
rect 1011 259 1017 260
rect 1011 258 1012 259
rect 1003 256 1012 258
rect 1003 255 1004 256
rect 998 254 1004 255
rect 1011 255 1012 256
rect 1016 255 1017 259
rect 1115 259 1121 260
rect 1115 258 1116 259
rect 1011 254 1017 255
rect 1028 256 1116 258
rect 732 248 778 250
rect 732 246 734 248
rect 1028 246 1030 256
rect 1115 255 1116 256
rect 1120 255 1121 259
rect 1219 259 1225 260
rect 1219 258 1220 259
rect 1115 254 1121 255
rect 1132 256 1220 258
rect 1132 246 1134 256
rect 1219 255 1220 256
rect 1224 255 1225 259
rect 1372 258 1374 260
rect 1550 259 1551 260
rect 1555 259 1556 263
rect 1738 263 1744 264
rect 1738 262 1739 263
rect 1550 258 1556 259
rect 1636 260 1739 262
rect 1636 258 1638 260
rect 1738 259 1739 260
rect 1743 259 1744 263
rect 2310 263 2316 264
rect 2310 262 2311 263
rect 1738 258 1744 259
rect 1908 260 2311 262
rect 1908 258 1910 260
rect 2310 259 2311 260
rect 2315 259 2316 263
rect 2310 258 2316 259
rect 1219 254 1225 255
rect 1371 257 1377 258
rect 1371 253 1372 257
rect 1376 253 1377 257
rect 1635 257 1641 258
rect 1443 255 1449 256
rect 1443 254 1444 255
rect 1371 252 1377 253
rect 1388 252 1444 254
rect 150 245 156 246
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 150 241 151 245
rect 155 241 156 245
rect 150 240 156 241
rect 171 245 177 246
rect 171 241 172 245
rect 176 241 177 245
rect 171 240 177 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 326 245 332 246
rect 230 240 236 241
rect 251 243 257 244
rect 110 239 116 240
rect 251 239 252 243
rect 256 242 257 243
rect 262 243 268 244
rect 262 242 263 243
rect 256 240 263 242
rect 256 239 257 240
rect 251 238 257 239
rect 262 239 263 240
rect 267 239 268 243
rect 326 241 327 245
rect 331 241 332 245
rect 422 245 428 246
rect 326 240 332 241
rect 346 243 353 244
rect 262 238 268 239
rect 346 239 347 243
rect 352 239 353 243
rect 422 241 423 245
rect 427 241 428 245
rect 422 240 428 241
rect 443 245 449 246
rect 443 241 444 245
rect 448 241 449 245
rect 443 240 449 241
rect 518 245 524 246
rect 518 241 519 245
rect 523 241 524 245
rect 614 245 620 246
rect 518 240 524 241
rect 539 243 548 244
rect 346 238 353 239
rect 539 239 540 243
rect 547 239 548 243
rect 614 241 615 245
rect 619 241 620 245
rect 710 245 716 246
rect 614 240 620 241
rect 634 243 641 244
rect 539 238 548 239
rect 634 239 635 243
rect 640 239 641 243
rect 710 241 711 245
rect 715 241 716 245
rect 710 240 716 241
rect 731 245 737 246
rect 731 241 732 245
rect 736 241 737 245
rect 731 240 737 241
rect 806 245 812 246
rect 806 241 807 245
rect 811 241 812 245
rect 902 245 908 246
rect 806 240 812 241
rect 827 243 833 244
rect 634 238 641 239
rect 827 239 828 243
rect 832 242 833 243
rect 878 243 884 244
rect 878 242 879 243
rect 832 240 879 242
rect 832 239 833 240
rect 827 238 833 239
rect 878 239 879 240
rect 883 239 884 243
rect 902 241 903 245
rect 907 241 908 245
rect 1006 245 1012 246
rect 902 240 908 241
rect 922 243 929 244
rect 878 238 884 239
rect 922 239 923 243
rect 928 239 929 243
rect 1006 241 1007 245
rect 1011 241 1012 245
rect 1006 240 1012 241
rect 1027 245 1033 246
rect 1027 241 1028 245
rect 1032 241 1033 245
rect 1027 240 1033 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1131 245 1137 246
rect 1131 241 1132 245
rect 1136 241 1137 245
rect 1131 240 1137 241
rect 1214 245 1220 246
rect 1214 241 1215 245
rect 1219 241 1220 245
rect 1286 244 1292 245
rect 1214 240 1220 241
rect 1222 243 1228 244
rect 922 238 929 239
rect 1222 239 1223 243
rect 1227 242 1228 243
rect 1235 243 1241 244
rect 1235 242 1236 243
rect 1227 240 1236 242
rect 1227 239 1228 240
rect 1222 238 1228 239
rect 1235 239 1236 240
rect 1240 239 1241 243
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1388 242 1390 252
rect 1443 251 1444 252
rect 1448 251 1449 255
rect 1539 255 1545 256
rect 1539 254 1540 255
rect 1443 250 1449 251
rect 1519 252 1540 254
rect 1519 250 1521 252
rect 1539 251 1540 252
rect 1544 251 1545 255
rect 1635 253 1636 257
rect 1640 253 1641 257
rect 1907 257 1913 258
rect 1731 255 1737 256
rect 1731 254 1732 255
rect 1635 252 1641 253
rect 1652 252 1732 254
rect 1539 250 1545 251
rect 1460 248 1521 250
rect 1460 242 1462 248
rect 1652 242 1654 252
rect 1731 251 1732 252
rect 1736 251 1737 255
rect 1819 255 1825 256
rect 1819 254 1820 255
rect 1731 250 1737 251
rect 1748 252 1820 254
rect 1748 242 1750 252
rect 1819 251 1820 252
rect 1824 251 1825 255
rect 1907 253 1908 257
rect 1912 253 1913 257
rect 2003 255 2009 256
rect 2003 254 2004 255
rect 1907 252 1913 253
rect 1924 252 2004 254
rect 1819 250 1825 251
rect 1806 247 1812 248
rect 1806 243 1807 247
rect 1811 246 1812 247
rect 1811 244 1838 246
rect 1811 243 1812 244
rect 1806 242 1812 243
rect 1836 242 1838 244
rect 1924 242 1926 252
rect 2003 251 2004 252
rect 2008 251 2009 255
rect 2107 255 2113 256
rect 2107 254 2108 255
rect 2003 250 2009 251
rect 2020 252 2108 254
rect 2020 242 2022 252
rect 2107 251 2108 252
rect 2112 251 2113 255
rect 2219 255 2225 256
rect 2219 254 2220 255
rect 2107 250 2113 251
rect 2125 252 2220 254
rect 2125 242 2127 252
rect 2219 251 2220 252
rect 2224 251 2225 255
rect 2339 255 2345 256
rect 2339 254 2340 255
rect 2219 250 2225 251
rect 2236 252 2340 254
rect 2236 242 2238 252
rect 2339 251 2340 252
rect 2344 251 2345 255
rect 2339 250 2345 251
rect 2459 255 2468 256
rect 2459 251 2460 255
rect 2467 251 2468 255
rect 2459 250 2468 251
rect 1366 241 1372 242
rect 1286 239 1292 240
rect 1326 240 1332 241
rect 1235 238 1241 239
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1387 241 1393 242
rect 1387 237 1388 241
rect 1392 237 1393 241
rect 1387 236 1393 237
rect 1438 241 1444 242
rect 1438 237 1439 241
rect 1443 237 1444 241
rect 1438 236 1444 237
rect 1459 241 1465 242
rect 1459 237 1460 241
rect 1464 237 1465 241
rect 1459 236 1465 237
rect 1534 241 1540 242
rect 1534 237 1535 241
rect 1539 237 1540 241
rect 1630 241 1636 242
rect 1534 236 1540 237
rect 1555 239 1561 240
rect 1326 235 1332 236
rect 1555 235 1556 239
rect 1560 238 1561 239
rect 1606 239 1612 240
rect 1606 238 1607 239
rect 1560 236 1607 238
rect 1560 235 1561 236
rect 1555 234 1561 235
rect 1606 235 1607 236
rect 1611 235 1612 239
rect 1630 237 1631 241
rect 1635 237 1636 241
rect 1630 236 1636 237
rect 1651 241 1657 242
rect 1651 237 1652 241
rect 1656 237 1657 241
rect 1651 236 1657 237
rect 1726 241 1732 242
rect 1726 237 1727 241
rect 1731 237 1732 241
rect 1726 236 1732 237
rect 1747 241 1753 242
rect 1747 237 1748 241
rect 1752 237 1753 241
rect 1747 236 1753 237
rect 1814 241 1820 242
rect 1814 237 1815 241
rect 1819 237 1820 241
rect 1814 236 1820 237
rect 1835 241 1841 242
rect 1835 237 1836 241
rect 1840 237 1841 241
rect 1835 236 1841 237
rect 1902 241 1908 242
rect 1902 237 1903 241
rect 1907 237 1908 241
rect 1902 236 1908 237
rect 1923 241 1929 242
rect 1923 237 1924 241
rect 1928 237 1929 241
rect 1923 236 1929 237
rect 1998 241 2004 242
rect 1998 237 1999 241
rect 2003 237 2004 241
rect 1998 236 2004 237
rect 2019 241 2025 242
rect 2019 237 2020 241
rect 2024 237 2025 241
rect 2019 236 2025 237
rect 2102 241 2108 242
rect 2102 237 2103 241
rect 2107 237 2108 241
rect 2102 236 2108 237
rect 2123 241 2129 242
rect 2123 237 2124 241
rect 2128 237 2129 241
rect 2123 236 2129 237
rect 2214 241 2220 242
rect 2214 237 2215 241
rect 2219 237 2220 241
rect 2214 236 2220 237
rect 2235 241 2241 242
rect 2235 237 2236 241
rect 2240 237 2241 241
rect 2235 236 2241 237
rect 2334 241 2340 242
rect 2334 237 2335 241
rect 2339 237 2340 241
rect 2454 241 2460 242
rect 2334 236 2340 237
rect 2342 239 2348 240
rect 1606 234 1612 235
rect 2342 235 2343 239
rect 2347 238 2348 239
rect 2355 239 2361 240
rect 2355 238 2356 239
rect 2347 236 2356 238
rect 2347 235 2348 236
rect 2342 234 2348 235
rect 2355 235 2356 236
rect 2360 235 2361 239
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2502 240 2508 241
rect 2454 236 2460 237
rect 2470 239 2481 240
rect 2355 234 2361 235
rect 2470 235 2471 239
rect 2475 235 2476 239
rect 2480 235 2481 239
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 2502 235 2508 236
rect 2470 234 2481 235
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 1286 227 1292 228
rect 110 222 116 223
rect 134 224 140 225
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 214 224 220 225
rect 214 220 215 224
rect 219 220 220 224
rect 214 219 220 220
rect 310 224 316 225
rect 310 220 311 224
rect 315 220 316 224
rect 310 219 316 220
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 502 224 508 225
rect 502 220 503 224
rect 507 220 508 224
rect 502 219 508 220
rect 598 224 604 225
rect 598 220 599 224
rect 603 220 604 224
rect 598 219 604 220
rect 694 224 700 225
rect 694 220 695 224
rect 699 220 700 224
rect 694 219 700 220
rect 790 224 796 225
rect 790 220 791 224
rect 795 220 796 224
rect 790 219 796 220
rect 886 224 892 225
rect 886 220 887 224
rect 891 220 892 224
rect 886 219 892 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 1094 224 1100 225
rect 1094 220 1095 224
rect 1099 220 1100 224
rect 1094 219 1100 220
rect 1198 224 1204 225
rect 1198 220 1199 224
rect 1203 220 1204 224
rect 1286 223 1287 227
rect 1291 223 1292 227
rect 1286 222 1292 223
rect 1326 223 1332 224
rect 1198 219 1204 220
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 2502 223 2508 224
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1422 220 1428 221
rect 1422 216 1423 220
rect 1427 216 1428 220
rect 1422 215 1428 216
rect 1518 220 1524 221
rect 1518 216 1519 220
rect 1523 216 1524 220
rect 1518 215 1524 216
rect 1614 220 1620 221
rect 1614 216 1615 220
rect 1619 216 1620 220
rect 1614 215 1620 216
rect 1710 220 1716 221
rect 1710 216 1711 220
rect 1715 216 1716 220
rect 1710 215 1716 216
rect 1798 220 1804 221
rect 1798 216 1799 220
rect 1803 216 1804 220
rect 1798 215 1804 216
rect 1886 220 1892 221
rect 1886 216 1887 220
rect 1891 216 1892 220
rect 1886 215 1892 216
rect 1982 220 1988 221
rect 1982 216 1983 220
rect 1987 216 1988 220
rect 1982 215 1988 216
rect 2086 220 2092 221
rect 2086 216 2087 220
rect 2091 216 2092 220
rect 2086 215 2092 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2318 220 2324 221
rect 2318 216 2319 220
rect 2323 216 2324 220
rect 2318 215 2324 216
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2438 215 2444 216
rect 158 204 164 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 158 200 159 204
rect 163 200 164 204
rect 158 199 164 200
rect 238 204 244 205
rect 238 200 239 204
rect 243 200 244 204
rect 238 199 244 200
rect 326 204 332 205
rect 326 200 327 204
rect 331 200 332 204
rect 326 199 332 200
rect 414 204 420 205
rect 414 200 415 204
rect 419 200 420 204
rect 414 199 420 200
rect 510 204 516 205
rect 510 200 511 204
rect 515 200 516 204
rect 510 199 516 200
rect 606 204 612 205
rect 606 200 607 204
rect 611 200 612 204
rect 606 199 612 200
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 782 204 788 205
rect 782 200 783 204
rect 787 200 788 204
rect 782 199 788 200
rect 870 204 876 205
rect 870 200 871 204
rect 875 200 876 204
rect 870 199 876 200
rect 958 204 964 205
rect 958 200 959 204
rect 963 200 964 204
rect 958 199 964 200
rect 1046 204 1052 205
rect 1046 200 1047 204
rect 1051 200 1052 204
rect 1046 199 1052 200
rect 1134 204 1140 205
rect 1134 200 1135 204
rect 1139 200 1140 204
rect 1390 204 1396 205
rect 1134 199 1140 200
rect 1286 201 1292 202
rect 110 196 116 197
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1390 200 1391 204
rect 1395 200 1396 204
rect 1390 199 1396 200
rect 1494 204 1500 205
rect 1494 200 1495 204
rect 1499 200 1500 204
rect 1494 199 1500 200
rect 1598 204 1604 205
rect 1598 200 1599 204
rect 1603 200 1604 204
rect 1598 199 1604 200
rect 1710 204 1716 205
rect 1710 200 1711 204
rect 1715 200 1716 204
rect 1710 199 1716 200
rect 1814 204 1820 205
rect 1814 200 1815 204
rect 1819 200 1820 204
rect 1814 199 1820 200
rect 1918 204 1924 205
rect 1918 200 1919 204
rect 1923 200 1924 204
rect 1918 199 1924 200
rect 2014 204 2020 205
rect 2014 200 2015 204
rect 2019 200 2020 204
rect 2014 199 2020 200
rect 2110 204 2116 205
rect 2110 200 2111 204
rect 2115 200 2116 204
rect 2110 199 2116 200
rect 2198 204 2204 205
rect 2198 200 2199 204
rect 2203 200 2204 204
rect 2198 199 2204 200
rect 2286 204 2292 205
rect 2286 200 2287 204
rect 2291 200 2292 204
rect 2286 199 2292 200
rect 2374 204 2380 205
rect 2374 200 2375 204
rect 2379 200 2380 204
rect 2374 199 2380 200
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2502 201 2508 202
rect 1326 196 1332 197
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 110 184 116 185
rect 1286 184 1292 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 174 183 180 184
rect 174 179 175 183
rect 179 179 180 183
rect 174 178 180 179
rect 182 183 188 184
rect 182 179 183 183
rect 187 182 188 183
rect 195 183 201 184
rect 195 182 196 183
rect 187 180 196 182
rect 187 179 188 180
rect 182 178 188 179
rect 195 179 196 180
rect 200 179 201 183
rect 195 178 201 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 179 260 183
rect 254 178 260 179
rect 275 183 281 184
rect 275 179 276 183
rect 280 182 281 183
rect 342 183 348 184
rect 280 180 321 182
rect 280 179 281 180
rect 275 178 281 179
rect 319 170 321 180
rect 342 179 343 183
rect 347 179 348 183
rect 342 178 348 179
rect 350 183 356 184
rect 350 179 351 183
rect 355 182 356 183
rect 363 183 369 184
rect 363 182 364 183
rect 355 180 364 182
rect 355 179 356 180
rect 350 178 356 179
rect 363 179 364 180
rect 368 179 369 183
rect 363 178 369 179
rect 430 183 436 184
rect 430 179 431 183
rect 435 179 436 183
rect 430 178 436 179
rect 451 183 457 184
rect 451 179 452 183
rect 456 182 457 183
rect 526 183 532 184
rect 456 180 518 182
rect 456 179 457 180
rect 451 178 457 179
rect 516 170 518 180
rect 526 179 527 183
rect 531 179 532 183
rect 526 178 532 179
rect 547 183 553 184
rect 547 179 548 183
rect 552 182 553 183
rect 622 183 628 184
rect 552 180 614 182
rect 552 179 553 180
rect 547 178 553 179
rect 612 170 614 180
rect 622 179 623 183
rect 627 179 628 183
rect 622 178 628 179
rect 642 183 649 184
rect 642 179 643 183
rect 648 179 649 183
rect 642 178 649 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 718 183 724 184
rect 718 179 719 183
rect 723 182 724 183
rect 731 183 737 184
rect 731 182 732 183
rect 723 180 732 182
rect 723 179 724 180
rect 718 178 724 179
rect 731 179 732 180
rect 736 179 737 183
rect 731 178 737 179
rect 798 183 804 184
rect 798 179 799 183
rect 803 179 804 183
rect 798 178 804 179
rect 814 183 825 184
rect 814 179 815 183
rect 819 179 820 183
rect 824 179 825 183
rect 814 178 825 179
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 907 183 913 184
rect 907 179 908 183
rect 912 179 913 183
rect 907 178 913 179
rect 974 183 980 184
rect 974 179 975 183
rect 979 179 980 183
rect 974 178 980 179
rect 995 183 1004 184
rect 995 179 996 183
rect 1003 179 1004 183
rect 995 178 1004 179
rect 1062 183 1068 184
rect 1062 179 1063 183
rect 1067 179 1068 183
rect 1083 183 1089 184
rect 1083 182 1084 183
rect 1062 178 1068 179
rect 1072 180 1084 182
rect 909 174 911 178
rect 1072 174 1074 180
rect 1083 179 1084 180
rect 1088 179 1089 183
rect 1083 178 1089 179
rect 1150 183 1156 184
rect 1150 179 1151 183
rect 1155 179 1156 183
rect 1171 183 1177 184
rect 1171 182 1172 183
rect 1150 178 1156 179
rect 1159 180 1172 182
rect 1159 174 1161 180
rect 1171 179 1172 180
rect 1176 179 1177 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 2502 184 2508 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1406 183 1412 184
rect 1406 179 1407 183
rect 1411 179 1412 183
rect 1171 178 1177 179
rect 1406 178 1412 179
rect 1414 183 1420 184
rect 1414 179 1415 183
rect 1419 182 1420 183
rect 1427 183 1433 184
rect 1427 182 1428 183
rect 1419 180 1428 182
rect 1419 179 1420 180
rect 1414 178 1420 179
rect 1427 179 1428 180
rect 1432 179 1433 183
rect 1427 178 1433 179
rect 1510 183 1516 184
rect 1510 179 1511 183
rect 1515 179 1516 183
rect 1510 178 1516 179
rect 1526 183 1537 184
rect 1526 179 1527 183
rect 1531 179 1532 183
rect 1536 179 1537 183
rect 1526 178 1537 179
rect 1614 183 1620 184
rect 1614 179 1615 183
rect 1619 179 1620 183
rect 1614 178 1620 179
rect 1635 183 1641 184
rect 1635 179 1636 183
rect 1640 179 1641 183
rect 1635 178 1641 179
rect 1726 183 1732 184
rect 1726 179 1727 183
rect 1731 179 1732 183
rect 1726 178 1732 179
rect 1738 183 1744 184
rect 1738 179 1739 183
rect 1743 182 1744 183
rect 1747 183 1753 184
rect 1747 182 1748 183
rect 1743 180 1748 182
rect 1743 179 1744 180
rect 1738 178 1744 179
rect 1747 179 1748 180
rect 1752 179 1753 183
rect 1747 178 1753 179
rect 1830 183 1836 184
rect 1830 179 1831 183
rect 1835 179 1836 183
rect 1851 183 1857 184
rect 1851 182 1852 183
rect 1830 178 1836 179
rect 1840 180 1852 182
rect 1637 174 1639 178
rect 1840 174 1842 180
rect 1851 179 1852 180
rect 1856 179 1857 183
rect 1851 178 1857 179
rect 1934 183 1940 184
rect 1934 179 1935 183
rect 1939 179 1940 183
rect 1934 178 1940 179
rect 1955 183 1961 184
rect 1955 179 1956 183
rect 1960 182 1961 183
rect 2030 183 2036 184
rect 1960 180 2001 182
rect 1960 179 1961 180
rect 1955 178 1961 179
rect 804 172 911 174
rect 980 172 1074 174
rect 1076 172 1161 174
rect 1516 172 1639 174
rect 1733 172 1842 174
rect 804 170 806 172
rect 980 170 982 172
rect 1076 170 1078 172
rect 1516 170 1518 172
rect 1733 170 1735 172
rect 1999 170 2001 180
rect 2030 179 2031 183
rect 2035 179 2036 183
rect 2030 178 2036 179
rect 2051 183 2057 184
rect 2051 179 2052 183
rect 2056 182 2057 183
rect 2126 183 2132 184
rect 2056 180 2122 182
rect 2056 179 2057 180
rect 2051 178 2057 179
rect 2120 170 2122 180
rect 2126 179 2127 183
rect 2131 179 2132 183
rect 2126 178 2132 179
rect 2147 183 2153 184
rect 2147 179 2148 183
rect 2152 182 2153 183
rect 2214 183 2220 184
rect 2152 180 2186 182
rect 2152 179 2153 180
rect 2147 178 2153 179
rect 2184 170 2186 180
rect 2214 179 2215 183
rect 2219 179 2220 183
rect 2214 178 2220 179
rect 2230 183 2241 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2240 179 2241 183
rect 2230 178 2241 179
rect 2302 183 2308 184
rect 2302 179 2303 183
rect 2307 179 2308 183
rect 2302 178 2308 179
rect 2323 183 2329 184
rect 2323 179 2324 183
rect 2328 182 2329 183
rect 2390 183 2396 184
rect 2328 180 2366 182
rect 2328 179 2329 180
rect 2323 178 2329 179
rect 2364 170 2366 180
rect 2390 179 2391 183
rect 2395 179 2396 183
rect 2390 178 2396 179
rect 2411 183 2420 184
rect 2411 179 2412 183
rect 2419 179 2420 183
rect 2411 178 2420 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2454 178 2460 179
rect 2462 183 2468 184
rect 2462 179 2463 183
rect 2467 182 2468 183
rect 2475 183 2481 184
rect 2475 182 2476 183
rect 2467 180 2476 182
rect 2467 179 2468 180
rect 2462 178 2468 179
rect 2475 179 2476 180
rect 2480 179 2481 183
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2475 178 2481 179
rect 319 169 353 170
rect 319 168 348 169
rect 179 167 185 168
rect 179 163 180 167
rect 184 166 185 167
rect 259 167 268 168
rect 184 164 254 166
rect 184 163 185 164
rect 179 162 185 163
rect 252 158 254 164
rect 259 163 260 167
rect 267 163 268 167
rect 347 165 348 168
rect 352 165 353 169
rect 516 169 537 170
rect 516 168 532 169
rect 347 164 353 165
rect 435 167 441 168
rect 259 162 268 163
rect 435 163 436 167
rect 440 166 441 167
rect 440 164 527 166
rect 531 165 532 168
rect 536 165 537 169
rect 612 169 633 170
rect 612 168 628 169
rect 531 164 537 165
rect 627 165 628 168
rect 632 165 633 169
rect 803 169 809 170
rect 627 164 633 165
rect 715 167 721 168
rect 440 163 441 164
rect 435 162 441 163
rect 525 162 527 164
rect 642 163 648 164
rect 642 162 643 163
rect 525 160 643 162
rect 350 159 356 160
rect 350 158 351 159
rect 252 156 351 158
rect 350 155 351 156
rect 355 155 356 159
rect 642 159 643 160
rect 647 159 648 163
rect 715 163 716 167
rect 720 163 721 167
rect 803 165 804 169
rect 808 165 809 169
rect 979 169 985 170
rect 803 164 809 165
rect 878 167 884 168
rect 715 162 721 163
rect 814 163 820 164
rect 814 162 815 163
rect 717 160 815 162
rect 642 158 648 159
rect 814 159 815 160
rect 819 159 820 163
rect 878 163 879 167
rect 883 166 884 167
rect 891 167 897 168
rect 891 166 892 167
rect 883 164 892 166
rect 883 163 884 164
rect 878 162 884 163
rect 891 163 892 164
rect 896 163 897 167
rect 979 165 980 169
rect 984 165 985 169
rect 979 164 985 165
rect 1067 169 1078 170
rect 1067 165 1068 169
rect 1072 168 1078 169
rect 1515 169 1521 170
rect 1072 165 1073 168
rect 1067 164 1073 165
rect 1155 167 1161 168
rect 891 162 897 163
rect 1155 163 1156 167
rect 1160 166 1161 167
rect 1218 167 1224 168
rect 1218 166 1219 167
rect 1160 164 1219 166
rect 1160 163 1161 164
rect 1155 162 1161 163
rect 1218 163 1219 164
rect 1223 163 1224 167
rect 1218 162 1224 163
rect 1411 167 1417 168
rect 1411 163 1412 167
rect 1416 166 1417 167
rect 1416 164 1474 166
rect 1515 165 1516 169
rect 1520 165 1521 169
rect 1731 169 1737 170
rect 1515 164 1521 165
rect 1606 167 1612 168
rect 1416 163 1417 164
rect 1411 162 1417 163
rect 1472 162 1474 164
rect 1526 163 1532 164
rect 1526 162 1527 163
rect 1472 160 1527 162
rect 814 158 820 159
rect 1526 159 1527 160
rect 1531 159 1532 163
rect 1606 163 1607 167
rect 1611 166 1612 167
rect 1619 167 1625 168
rect 1619 166 1620 167
rect 1611 164 1620 166
rect 1611 163 1612 164
rect 1606 162 1612 163
rect 1619 163 1620 164
rect 1624 163 1625 167
rect 1731 165 1732 169
rect 1736 165 1737 169
rect 1999 169 2041 170
rect 1999 168 2036 169
rect 1731 164 1737 165
rect 1835 167 1844 168
rect 1619 162 1625 163
rect 1835 163 1836 167
rect 1843 163 1844 167
rect 1835 162 1844 163
rect 1939 167 1945 168
rect 1939 163 1940 167
rect 1944 166 1945 167
rect 1944 164 2001 166
rect 2035 165 2036 168
rect 2040 165 2041 169
rect 2120 169 2137 170
rect 2120 168 2132 169
rect 2035 164 2041 165
rect 2131 165 2132 168
rect 2136 165 2137 169
rect 2184 169 2225 170
rect 2184 168 2220 169
rect 2131 164 2137 165
rect 2219 165 2220 168
rect 2224 165 2225 169
rect 2364 169 2401 170
rect 2364 168 2396 169
rect 2219 164 2225 165
rect 2307 167 2313 168
rect 1944 163 1945 164
rect 1939 162 1945 163
rect 1526 158 1532 159
rect 1999 158 2001 164
rect 2307 163 2308 167
rect 2312 166 2313 167
rect 2354 167 2360 168
rect 2354 166 2355 167
rect 2312 164 2355 166
rect 2312 163 2313 164
rect 2307 162 2313 163
rect 2354 163 2355 164
rect 2359 163 2360 167
rect 2395 165 2396 168
rect 2400 165 2401 169
rect 2395 164 2401 165
rect 2459 167 2465 168
rect 2354 162 2360 163
rect 2459 163 2460 167
rect 2464 166 2465 167
rect 2470 167 2476 168
rect 2470 166 2471 167
rect 2464 164 2471 166
rect 2464 163 2465 164
rect 2459 162 2465 163
rect 2470 163 2471 164
rect 2475 163 2476 167
rect 2470 162 2476 163
rect 2342 159 2348 160
rect 2342 158 2343 159
rect 1999 156 2343 158
rect 350 154 356 155
rect 2342 155 2343 156
rect 2347 155 2348 159
rect 2342 154 2348 155
rect 182 135 188 136
rect 182 131 183 135
rect 187 131 188 135
rect 718 135 724 136
rect 718 134 719 135
rect 182 130 188 131
rect 692 132 719 134
rect 692 130 694 132
rect 718 131 719 132
rect 723 131 724 135
rect 718 130 724 131
rect 1414 135 1420 136
rect 1414 131 1415 135
rect 1419 131 1420 135
rect 2230 135 2236 136
rect 2230 134 2231 135
rect 1414 130 1420 131
rect 1876 132 2231 134
rect 1876 130 1878 132
rect 2230 131 2231 132
rect 2235 131 2236 135
rect 2230 130 2236 131
rect 155 129 186 130
rect 155 125 156 129
rect 160 128 186 129
rect 691 129 697 130
rect 160 125 161 128
rect 211 127 217 128
rect 211 126 212 127
rect 155 124 161 125
rect 172 124 212 126
rect 172 114 174 124
rect 211 123 212 124
rect 216 123 217 127
rect 267 127 273 128
rect 267 126 268 127
rect 211 122 217 123
rect 228 124 268 126
rect 228 114 230 124
rect 267 123 268 124
rect 272 123 273 127
rect 323 127 329 128
rect 323 126 324 127
rect 267 122 273 123
rect 319 124 324 126
rect 319 118 321 124
rect 323 123 324 124
rect 328 123 329 127
rect 379 127 385 128
rect 379 126 380 127
rect 323 122 329 123
rect 340 124 380 126
rect 284 116 321 118
rect 284 114 286 116
rect 340 114 342 124
rect 379 123 380 124
rect 384 123 385 127
rect 435 127 441 128
rect 435 126 436 127
rect 379 122 385 123
rect 396 124 436 126
rect 396 114 398 124
rect 435 123 436 124
rect 440 123 441 127
rect 491 127 497 128
rect 491 126 492 127
rect 435 122 441 123
rect 452 124 492 126
rect 452 114 454 124
rect 491 123 492 124
rect 496 123 497 127
rect 555 127 561 128
rect 555 126 556 127
rect 491 122 497 123
rect 508 124 556 126
rect 508 114 510 124
rect 555 123 556 124
rect 560 123 561 127
rect 627 127 633 128
rect 627 126 628 127
rect 555 122 561 123
rect 572 124 628 126
rect 572 114 574 124
rect 627 123 628 124
rect 632 123 633 127
rect 691 125 692 129
rect 696 125 697 129
rect 1371 129 1418 130
rect 755 127 761 128
rect 755 126 756 127
rect 691 124 697 125
rect 708 124 756 126
rect 627 122 633 123
rect 708 114 710 124
rect 755 123 756 124
rect 760 123 761 127
rect 819 127 825 128
rect 819 126 820 127
rect 755 122 761 123
rect 772 124 820 126
rect 772 114 774 124
rect 819 123 820 124
rect 824 123 825 127
rect 883 127 889 128
rect 883 126 884 127
rect 819 122 825 123
rect 836 124 884 126
rect 836 114 838 124
rect 883 123 884 124
rect 888 123 889 127
rect 947 127 953 128
rect 947 126 948 127
rect 883 122 889 123
rect 900 124 948 126
rect 900 114 902 124
rect 947 123 948 124
rect 952 123 953 127
rect 947 122 953 123
rect 1011 127 1017 128
rect 1011 123 1012 127
rect 1016 123 1017 127
rect 1075 127 1081 128
rect 1075 126 1076 127
rect 1011 122 1017 123
rect 1028 124 1076 126
rect 1013 118 1015 122
rect 964 116 1015 118
rect 964 114 966 116
rect 1028 114 1030 124
rect 1075 123 1076 124
rect 1080 123 1081 127
rect 1139 127 1145 128
rect 1139 126 1140 127
rect 1075 122 1081 123
rect 1092 124 1140 126
rect 1092 114 1094 124
rect 1139 123 1140 124
rect 1144 123 1145 127
rect 1203 127 1209 128
rect 1203 126 1204 127
rect 1139 122 1145 123
rect 1159 124 1204 126
rect 1159 114 1161 124
rect 1203 123 1204 124
rect 1208 123 1209 127
rect 1371 125 1372 129
rect 1376 128 1418 129
rect 1875 129 1881 130
rect 1376 125 1377 128
rect 1427 127 1433 128
rect 1427 126 1428 127
rect 1371 124 1377 125
rect 1388 124 1428 126
rect 1203 122 1209 123
rect 1388 114 1390 124
rect 1427 123 1428 124
rect 1432 123 1433 127
rect 1483 127 1489 128
rect 1483 126 1484 127
rect 1427 122 1433 123
rect 1445 124 1484 126
rect 1445 114 1447 124
rect 1483 123 1484 124
rect 1488 123 1489 127
rect 1483 122 1489 123
rect 1539 127 1545 128
rect 1539 123 1540 127
rect 1544 123 1545 127
rect 1595 127 1601 128
rect 1595 126 1596 127
rect 1539 122 1545 123
rect 1556 124 1596 126
rect 1541 118 1543 122
rect 1500 116 1543 118
rect 1500 114 1502 116
rect 1556 114 1558 124
rect 1595 123 1596 124
rect 1600 123 1601 127
rect 1651 127 1657 128
rect 1651 126 1652 127
rect 1595 122 1601 123
rect 1612 124 1652 126
rect 1612 114 1614 124
rect 1651 123 1652 124
rect 1656 123 1657 127
rect 1707 127 1713 128
rect 1707 126 1708 127
rect 1651 122 1657 123
rect 1668 124 1708 126
rect 1668 114 1670 124
rect 1707 123 1708 124
rect 1712 123 1713 127
rect 1763 127 1769 128
rect 1763 126 1764 127
rect 1707 122 1713 123
rect 1724 124 1764 126
rect 1724 114 1726 124
rect 1763 123 1764 124
rect 1768 123 1769 127
rect 1763 122 1769 123
rect 1819 127 1825 128
rect 1819 123 1820 127
rect 1824 123 1825 127
rect 1875 125 1876 129
rect 1880 125 1881 129
rect 1875 124 1881 125
rect 1931 127 1937 128
rect 1819 122 1825 123
rect 1931 123 1932 127
rect 1936 123 1937 127
rect 1987 127 1993 128
rect 1987 126 1988 127
rect 1931 122 1937 123
rect 1948 124 1988 126
rect 1821 118 1823 122
rect 1933 118 1935 122
rect 1780 116 1823 118
rect 1892 116 1935 118
rect 1780 114 1782 116
rect 1892 114 1894 116
rect 1948 114 1950 124
rect 1987 123 1988 124
rect 1992 123 1993 127
rect 1987 122 1993 123
rect 2043 127 2049 128
rect 2043 123 2044 127
rect 2048 123 2049 127
rect 2099 127 2105 128
rect 2099 126 2100 127
rect 2043 122 2049 123
rect 2060 124 2100 126
rect 2045 118 2047 122
rect 2005 116 2047 118
rect 2005 114 2007 116
rect 2060 114 2062 124
rect 2099 123 2100 124
rect 2104 123 2105 127
rect 2163 127 2169 128
rect 2163 126 2164 127
rect 2099 122 2105 123
rect 2116 124 2164 126
rect 2116 114 2118 124
rect 2163 123 2164 124
rect 2168 123 2169 127
rect 2227 127 2233 128
rect 2227 126 2228 127
rect 2163 122 2169 123
rect 2180 124 2228 126
rect 2180 114 2182 124
rect 2227 123 2228 124
rect 2232 123 2233 127
rect 2291 127 2297 128
rect 2291 126 2292 127
rect 2227 122 2233 123
rect 2244 124 2292 126
rect 2244 114 2246 124
rect 2291 123 2292 124
rect 2296 123 2297 127
rect 2347 127 2353 128
rect 2347 126 2348 127
rect 2291 122 2297 123
rect 2309 124 2348 126
rect 2309 114 2311 124
rect 2347 123 2348 124
rect 2352 123 2353 127
rect 2347 122 2353 123
rect 2403 127 2409 128
rect 2403 123 2404 127
rect 2408 126 2409 127
rect 2459 127 2468 128
rect 2408 124 2454 126
rect 2408 123 2409 124
rect 2403 122 2409 123
rect 2452 118 2454 124
rect 2459 123 2460 127
rect 2467 123 2468 127
rect 2459 122 2468 123
rect 2452 116 2478 118
rect 2476 114 2478 116
rect 150 113 156 114
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 150 109 151 113
rect 155 109 156 113
rect 150 108 156 109
rect 171 113 177 114
rect 171 109 172 113
rect 176 109 177 113
rect 171 108 177 109
rect 206 113 212 114
rect 206 109 207 113
rect 211 109 212 113
rect 206 108 212 109
rect 227 113 233 114
rect 227 109 228 113
rect 232 109 233 113
rect 227 108 233 109
rect 262 113 268 114
rect 262 109 263 113
rect 267 109 268 113
rect 262 108 268 109
rect 283 113 289 114
rect 283 109 284 113
rect 288 109 289 113
rect 283 108 289 109
rect 318 113 324 114
rect 318 109 319 113
rect 323 109 324 113
rect 318 108 324 109
rect 339 113 345 114
rect 339 109 340 113
rect 344 109 345 113
rect 339 108 345 109
rect 374 113 380 114
rect 374 109 375 113
rect 379 109 380 113
rect 374 108 380 109
rect 395 113 401 114
rect 395 109 396 113
rect 400 109 401 113
rect 395 108 401 109
rect 430 113 436 114
rect 430 109 431 113
rect 435 109 436 113
rect 430 108 436 109
rect 451 113 457 114
rect 451 109 452 113
rect 456 109 457 113
rect 451 108 457 109
rect 486 113 492 114
rect 486 109 487 113
rect 491 109 492 113
rect 486 108 492 109
rect 507 113 513 114
rect 507 109 508 113
rect 512 109 513 113
rect 507 108 513 109
rect 550 113 556 114
rect 550 109 551 113
rect 555 109 556 113
rect 550 108 556 109
rect 571 113 577 114
rect 571 109 572 113
rect 576 109 577 113
rect 571 108 577 109
rect 622 113 628 114
rect 622 109 623 113
rect 627 109 628 113
rect 686 113 692 114
rect 622 108 628 109
rect 642 111 649 112
rect 110 107 116 108
rect 642 107 643 111
rect 648 107 649 111
rect 686 109 687 113
rect 691 109 692 113
rect 686 108 692 109
rect 707 113 713 114
rect 707 109 708 113
rect 712 109 713 113
rect 707 108 713 109
rect 750 113 756 114
rect 750 109 751 113
rect 755 109 756 113
rect 750 108 756 109
rect 771 113 777 114
rect 771 109 772 113
rect 776 109 777 113
rect 771 108 777 109
rect 814 113 820 114
rect 814 109 815 113
rect 819 109 820 113
rect 814 108 820 109
rect 835 113 841 114
rect 835 109 836 113
rect 840 109 841 113
rect 835 108 841 109
rect 878 113 884 114
rect 878 109 879 113
rect 883 109 884 113
rect 878 108 884 109
rect 899 113 905 114
rect 899 109 900 113
rect 904 109 905 113
rect 899 108 905 109
rect 942 113 948 114
rect 942 109 943 113
rect 947 109 948 113
rect 942 108 948 109
rect 963 113 969 114
rect 963 109 964 113
rect 968 109 969 113
rect 963 108 969 109
rect 1006 113 1012 114
rect 1006 109 1007 113
rect 1011 109 1012 113
rect 1006 108 1012 109
rect 1027 113 1033 114
rect 1027 109 1028 113
rect 1032 109 1033 113
rect 1027 108 1033 109
rect 1070 113 1076 114
rect 1070 109 1071 113
rect 1075 109 1076 113
rect 1070 108 1076 109
rect 1091 113 1097 114
rect 1091 109 1092 113
rect 1096 109 1097 113
rect 1091 108 1097 109
rect 1134 113 1140 114
rect 1134 109 1135 113
rect 1139 109 1140 113
rect 1134 108 1140 109
rect 1155 113 1161 114
rect 1155 109 1156 113
rect 1160 109 1161 113
rect 1155 108 1161 109
rect 1198 113 1204 114
rect 1366 113 1372 114
rect 1198 109 1199 113
rect 1203 109 1204 113
rect 1286 112 1292 113
rect 1198 108 1204 109
rect 1218 111 1225 112
rect 642 106 649 107
rect 1218 107 1219 111
rect 1224 107 1225 111
rect 1286 108 1287 112
rect 1291 108 1292 112
rect 1286 107 1292 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1387 113 1393 114
rect 1387 109 1388 113
rect 1392 109 1393 113
rect 1387 108 1393 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1443 113 1449 114
rect 1443 109 1444 113
rect 1448 109 1449 113
rect 1443 108 1449 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1499 113 1505 114
rect 1499 109 1500 113
rect 1504 109 1505 113
rect 1499 108 1505 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1555 113 1561 114
rect 1555 109 1556 113
rect 1560 109 1561 113
rect 1555 108 1561 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1611 113 1617 114
rect 1611 109 1612 113
rect 1616 109 1617 113
rect 1611 108 1617 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1667 113 1673 114
rect 1667 109 1668 113
rect 1672 109 1673 113
rect 1667 108 1673 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1723 113 1729 114
rect 1723 109 1724 113
rect 1728 109 1729 113
rect 1723 108 1729 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1779 113 1785 114
rect 1779 109 1780 113
rect 1784 109 1785 113
rect 1779 108 1785 109
rect 1814 113 1820 114
rect 1814 109 1815 113
rect 1819 109 1820 113
rect 1870 113 1876 114
rect 1814 108 1820 109
rect 1835 111 1844 112
rect 1326 107 1332 108
rect 1835 107 1836 111
rect 1843 107 1844 111
rect 1870 109 1871 113
rect 1875 109 1876 113
rect 1870 108 1876 109
rect 1891 113 1897 114
rect 1891 109 1892 113
rect 1896 109 1897 113
rect 1891 108 1897 109
rect 1926 113 1932 114
rect 1926 109 1927 113
rect 1931 109 1932 113
rect 1926 108 1932 109
rect 1947 113 1953 114
rect 1947 109 1948 113
rect 1952 109 1953 113
rect 1947 108 1953 109
rect 1982 113 1988 114
rect 1982 109 1983 113
rect 1987 109 1988 113
rect 1982 108 1988 109
rect 2003 113 2009 114
rect 2003 109 2004 113
rect 2008 109 2009 113
rect 2003 108 2009 109
rect 2038 113 2044 114
rect 2038 109 2039 113
rect 2043 109 2044 113
rect 2038 108 2044 109
rect 2059 113 2065 114
rect 2059 109 2060 113
rect 2064 109 2065 113
rect 2059 108 2065 109
rect 2094 113 2100 114
rect 2094 109 2095 113
rect 2099 109 2100 113
rect 2094 108 2100 109
rect 2115 113 2121 114
rect 2115 109 2116 113
rect 2120 109 2121 113
rect 2115 108 2121 109
rect 2158 113 2164 114
rect 2158 109 2159 113
rect 2163 109 2164 113
rect 2158 108 2164 109
rect 2179 113 2185 114
rect 2179 109 2180 113
rect 2184 109 2185 113
rect 2179 108 2185 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2243 113 2249 114
rect 2243 109 2244 113
rect 2248 109 2249 113
rect 2243 108 2249 109
rect 2286 113 2292 114
rect 2286 109 2287 113
rect 2291 109 2292 113
rect 2286 108 2292 109
rect 2307 113 2313 114
rect 2307 109 2308 113
rect 2312 109 2313 113
rect 2307 108 2313 109
rect 2342 113 2348 114
rect 2342 109 2343 113
rect 2347 109 2348 113
rect 2398 113 2404 114
rect 2342 108 2348 109
rect 2354 111 2360 112
rect 1218 106 1225 107
rect 1835 106 1844 107
rect 2354 107 2355 111
rect 2359 110 2360 111
rect 2363 111 2369 112
rect 2363 110 2364 111
rect 2359 108 2364 110
rect 2359 107 2360 108
rect 2354 106 2360 107
rect 2363 107 2364 108
rect 2368 107 2369 111
rect 2398 109 2399 113
rect 2403 109 2404 113
rect 2398 108 2404 109
rect 2454 113 2460 114
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2475 113 2481 114
rect 2475 109 2476 113
rect 2480 109 2481 113
rect 2475 108 2481 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 2502 107 2508 108
rect 2363 106 2369 107
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1286 95 1292 96
rect 110 90 116 91
rect 134 92 140 93
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 246 92 252 93
rect 246 88 247 92
rect 251 88 252 92
rect 246 87 252 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 358 92 364 93
rect 358 88 359 92
rect 363 88 364 92
rect 358 87 364 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 606 92 612 93
rect 606 88 607 92
rect 611 88 612 92
rect 606 87 612 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 798 92 804 93
rect 798 88 799 92
rect 803 88 804 92
rect 798 87 804 88
rect 862 92 868 93
rect 862 88 863 92
rect 867 88 868 92
rect 862 87 868 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1054 92 1060 93
rect 1054 88 1055 92
rect 1059 88 1060 92
rect 1054 87 1060 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1182 92 1188 93
rect 1182 88 1183 92
rect 1187 88 1188 92
rect 1286 91 1287 95
rect 1291 91 1292 95
rect 1286 90 1292 91
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1182 87 1188 88
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1798 92 1804 93
rect 1798 88 1799 92
rect 1803 88 1804 92
rect 1798 87 1804 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1910 92 1916 93
rect 1910 88 1911 92
rect 1915 88 1916 92
rect 1910 87 1916 88
rect 1966 92 1972 93
rect 1966 88 1967 92
rect 1971 88 1972 92
rect 1966 87 1972 88
rect 2022 92 2028 93
rect 2022 88 2023 92
rect 2027 88 2028 92
rect 2022 87 2028 88
rect 2078 92 2084 93
rect 2078 88 2079 92
rect 2083 88 2084 92
rect 2078 87 2084 88
rect 2142 92 2148 93
rect 2142 88 2143 92
rect 2147 88 2148 92
rect 2142 87 2148 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2270 92 2276 93
rect 2270 88 2271 92
rect 2275 88 2276 92
rect 2270 87 2276 88
rect 2326 92 2332 93
rect 2326 88 2327 92
rect 2331 88 2332 92
rect 2326 87 2332 88
rect 2382 92 2388 93
rect 2382 88 2383 92
rect 2387 88 2388 92
rect 2382 87 2388 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
<< m3c >>
rect 111 2552 115 2556
rect 719 2553 723 2557
rect 775 2553 779 2557
rect 831 2553 835 2557
rect 887 2553 891 2557
rect 943 2553 947 2557
rect 951 2551 955 2555
rect 1287 2552 1291 2556
rect 1711 2551 1715 2555
rect 111 2535 115 2539
rect 703 2532 707 2536
rect 759 2532 763 2536
rect 815 2532 819 2536
rect 871 2532 875 2536
rect 927 2532 931 2536
rect 1287 2535 1291 2539
rect 1327 2528 1331 2532
rect 1399 2529 1403 2533
rect 1455 2529 1459 2533
rect 1511 2529 1515 2533
rect 1567 2529 1571 2533
rect 1623 2529 1627 2533
rect 1679 2529 1683 2533
rect 1735 2529 1739 2533
rect 1791 2529 1795 2533
rect 1847 2529 1851 2533
rect 1903 2529 1907 2533
rect 1959 2529 1963 2533
rect 2015 2529 2019 2533
rect 2071 2529 2075 2533
rect 2127 2529 2131 2533
rect 2183 2529 2187 2533
rect 2191 2527 2195 2531
rect 2503 2528 2507 2532
rect 111 2517 115 2521
rect 167 2520 171 2524
rect 223 2520 227 2524
rect 279 2520 283 2524
rect 343 2520 347 2524
rect 407 2520 411 2524
rect 479 2520 483 2524
rect 559 2520 563 2524
rect 639 2520 643 2524
rect 719 2520 723 2524
rect 799 2520 803 2524
rect 879 2520 883 2524
rect 959 2520 963 2524
rect 1039 2520 1043 2524
rect 1287 2517 1291 2521
rect 1327 2511 1331 2515
rect 1383 2508 1387 2512
rect 1439 2508 1443 2512
rect 1495 2508 1499 2512
rect 1551 2508 1555 2512
rect 1607 2508 1611 2512
rect 1663 2508 1667 2512
rect 1719 2508 1723 2512
rect 1775 2508 1779 2512
rect 1831 2508 1835 2512
rect 1887 2508 1891 2512
rect 1943 2508 1947 2512
rect 1999 2508 2003 2512
rect 2055 2508 2059 2512
rect 2111 2508 2115 2512
rect 2167 2508 2171 2512
rect 2503 2511 2507 2515
rect 111 2500 115 2504
rect 183 2499 187 2503
rect 239 2499 243 2503
rect 255 2499 259 2503
rect 295 2499 299 2503
rect 359 2499 363 2503
rect 423 2499 427 2503
rect 495 2499 499 2503
rect 575 2499 579 2503
rect 591 2499 595 2503
rect 655 2499 659 2503
rect 735 2499 739 2503
rect 815 2499 819 2503
rect 895 2499 899 2503
rect 975 2499 979 2503
rect 1055 2499 1059 2503
rect 1071 2499 1075 2503
rect 1287 2500 1291 2504
rect 1799 2495 1803 2499
rect 2191 2495 2195 2499
rect 591 2479 595 2483
rect 623 2483 627 2487
rect 1327 2485 1331 2489
rect 1351 2488 1355 2492
rect 1423 2488 1427 2492
rect 1511 2488 1515 2492
rect 1599 2488 1603 2492
rect 1687 2488 1691 2492
rect 1775 2488 1779 2492
rect 1863 2488 1867 2492
rect 1951 2488 1955 2492
rect 2039 2488 2043 2492
rect 2127 2488 2131 2492
rect 2503 2485 2507 2489
rect 951 2479 955 2483
rect 435 2471 439 2475
rect 715 2471 719 2475
rect 1071 2471 1075 2475
rect 255 2463 256 2467
rect 256 2463 259 2467
rect 763 2463 767 2467
rect 1327 2468 1331 2472
rect 1367 2467 1371 2471
rect 1439 2467 1443 2471
rect 1527 2467 1531 2471
rect 1615 2467 1619 2471
rect 1703 2467 1707 2471
rect 1711 2467 1715 2471
rect 1791 2467 1795 2471
rect 1879 2467 1883 2471
rect 1967 2467 1971 2471
rect 2055 2467 2059 2471
rect 2143 2467 2147 2471
rect 2151 2467 2155 2471
rect 2503 2468 2507 2472
rect 111 2448 115 2452
rect 183 2449 187 2453
rect 191 2447 195 2451
rect 247 2449 251 2453
rect 327 2449 331 2453
rect 415 2449 419 2453
rect 435 2447 436 2451
rect 436 2447 439 2451
rect 503 2449 507 2453
rect 599 2449 603 2453
rect 623 2447 624 2451
rect 624 2447 627 2451
rect 695 2449 699 2453
rect 715 2447 716 2451
rect 716 2447 719 2451
rect 791 2449 795 2453
rect 879 2449 883 2453
rect 967 2449 971 2453
rect 1063 2449 1067 2453
rect 1159 2449 1163 2453
rect 1183 2447 1184 2451
rect 1184 2447 1187 2451
rect 1287 2448 1291 2452
rect 1659 2447 1663 2451
rect 1799 2451 1800 2455
rect 1800 2451 1803 2455
rect 111 2431 115 2435
rect 167 2428 171 2432
rect 231 2428 235 2432
rect 311 2428 315 2432
rect 399 2428 403 2432
rect 487 2428 491 2432
rect 583 2428 587 2432
rect 679 2428 683 2432
rect 775 2428 779 2432
rect 863 2428 867 2432
rect 951 2428 955 2432
rect 1047 2428 1051 2432
rect 1143 2428 1147 2432
rect 1287 2431 1291 2435
rect 1375 2423 1376 2427
rect 1376 2423 1379 2427
rect 111 2409 115 2413
rect 151 2412 155 2416
rect 231 2412 235 2416
rect 319 2412 323 2416
rect 415 2412 419 2416
rect 519 2412 523 2416
rect 623 2412 627 2416
rect 727 2412 731 2416
rect 831 2412 835 2416
rect 935 2412 939 2416
rect 1039 2412 1043 2416
rect 1151 2412 1155 2416
rect 2151 2423 2155 2427
rect 1287 2409 1291 2413
rect 1327 2408 1331 2412
rect 1367 2409 1371 2413
rect 1439 2409 1443 2413
rect 1543 2409 1547 2413
rect 1639 2409 1643 2413
rect 1659 2407 1660 2411
rect 1660 2407 1663 2411
rect 1735 2409 1739 2413
rect 1759 2407 1760 2411
rect 1760 2407 1763 2411
rect 1823 2409 1827 2413
rect 1911 2409 1915 2413
rect 2007 2409 2011 2413
rect 2103 2409 2107 2413
rect 2503 2408 2507 2412
rect 111 2392 115 2396
rect 167 2391 171 2395
rect 247 2391 251 2395
rect 335 2391 339 2395
rect 431 2391 435 2395
rect 439 2391 443 2395
rect 535 2391 539 2395
rect 639 2391 643 2395
rect 743 2391 747 2395
rect 763 2391 764 2395
rect 764 2391 767 2395
rect 847 2391 851 2395
rect 951 2391 955 2395
rect 1055 2391 1059 2395
rect 1167 2391 1171 2395
rect 1175 2391 1179 2395
rect 1287 2392 1291 2396
rect 1327 2391 1331 2395
rect 1351 2388 1355 2392
rect 1423 2388 1427 2392
rect 1527 2388 1531 2392
rect 1623 2388 1627 2392
rect 1719 2388 1723 2392
rect 1807 2388 1811 2392
rect 1895 2388 1899 2392
rect 1991 2388 1995 2392
rect 2087 2388 2091 2392
rect 2503 2391 2507 2395
rect 191 2375 195 2379
rect 631 2371 635 2375
rect 1183 2371 1187 2375
rect 439 2363 443 2367
rect 1147 2363 1151 2367
rect 1327 2365 1331 2369
rect 1351 2368 1355 2372
rect 1407 2368 1411 2372
rect 1495 2368 1499 2372
rect 1583 2368 1587 2372
rect 1671 2368 1675 2372
rect 1751 2368 1755 2372
rect 1831 2368 1835 2372
rect 1919 2368 1923 2372
rect 2007 2368 2011 2372
rect 2095 2368 2099 2372
rect 2503 2365 2507 2369
rect 771 2355 775 2359
rect 1175 2355 1179 2359
rect 1327 2348 1331 2352
rect 1367 2347 1371 2351
rect 1375 2347 1379 2351
rect 1423 2347 1427 2351
rect 111 2340 115 2344
rect 175 2341 179 2345
rect 279 2341 283 2345
rect 391 2341 395 2345
rect 503 2341 507 2345
rect 511 2339 515 2343
rect 623 2341 627 2345
rect 631 2339 635 2343
rect 743 2341 747 2345
rect 871 2341 875 2345
rect 999 2341 1003 2345
rect 1015 2339 1019 2343
rect 1127 2341 1131 2345
rect 1147 2339 1148 2343
rect 1148 2339 1151 2343
rect 1287 2340 1291 2344
rect 1511 2347 1515 2351
rect 1599 2347 1603 2351
rect 1687 2347 1691 2351
rect 1695 2347 1699 2351
rect 1767 2347 1771 2351
rect 1847 2347 1851 2351
rect 1935 2347 1939 2351
rect 2023 2347 2027 2351
rect 2111 2347 2115 2351
rect 2119 2347 2123 2351
rect 2503 2348 2507 2352
rect 111 2323 115 2327
rect 159 2320 163 2324
rect 263 2320 267 2324
rect 375 2320 379 2324
rect 487 2320 491 2324
rect 607 2320 611 2324
rect 727 2320 731 2324
rect 855 2320 859 2324
rect 983 2320 987 2324
rect 1111 2320 1115 2324
rect 1287 2323 1291 2327
rect 1567 2331 1571 2335
rect 1759 2331 1763 2335
rect 1695 2323 1699 2327
rect 1659 2315 1663 2319
rect 2119 2315 2123 2319
rect 111 2301 115 2305
rect 207 2304 211 2308
rect 287 2304 291 2308
rect 375 2304 379 2308
rect 471 2304 475 2308
rect 559 2304 563 2308
rect 647 2304 651 2308
rect 735 2304 739 2308
rect 815 2304 819 2308
rect 903 2304 907 2308
rect 991 2304 995 2308
rect 1079 2304 1083 2308
rect 1287 2301 1291 2305
rect 1823 2307 1827 2311
rect 1327 2292 1331 2296
rect 1367 2293 1371 2297
rect 1455 2293 1459 2297
rect 1543 2293 1547 2297
rect 1567 2291 1568 2295
rect 1568 2291 1571 2295
rect 1639 2293 1643 2297
rect 1659 2291 1660 2295
rect 1660 2291 1663 2295
rect 1735 2293 1739 2297
rect 1831 2293 1835 2297
rect 1927 2293 1931 2297
rect 2015 2293 2019 2297
rect 2111 2293 2115 2297
rect 2207 2293 2211 2297
rect 2223 2291 2227 2295
rect 2503 2292 2507 2296
rect 111 2284 115 2288
rect 223 2283 227 2287
rect 303 2283 307 2287
rect 391 2283 395 2287
rect 487 2283 491 2287
rect 495 2283 499 2287
rect 575 2283 579 2287
rect 663 2283 667 2287
rect 751 2283 755 2287
rect 771 2283 772 2287
rect 772 2283 775 2287
rect 831 2283 835 2287
rect 919 2283 923 2287
rect 975 2283 979 2287
rect 1007 2283 1011 2287
rect 1095 2283 1099 2287
rect 1103 2283 1107 2287
rect 1287 2284 1291 2288
rect 1327 2275 1331 2279
rect 511 2263 515 2267
rect 583 2267 584 2271
rect 584 2267 587 2271
rect 1015 2267 1016 2271
rect 1016 2267 1019 2271
rect 1351 2272 1355 2276
rect 1439 2272 1443 2276
rect 1527 2272 1531 2276
rect 1623 2272 1627 2276
rect 1719 2272 1723 2276
rect 1815 2272 1819 2276
rect 1911 2272 1915 2276
rect 1823 2267 1827 2271
rect 1999 2272 2003 2276
rect 2095 2272 2099 2276
rect 2191 2272 2195 2276
rect 2503 2275 2507 2279
rect 1875 2267 1879 2271
rect 1103 2259 1107 2263
rect 1327 2257 1331 2261
rect 1455 2260 1459 2264
rect 1543 2260 1547 2264
rect 1639 2260 1643 2264
rect 1735 2260 1739 2264
rect 1839 2260 1843 2264
rect 1935 2260 1939 2264
rect 2031 2260 2035 2264
rect 2119 2260 2123 2264
rect 2215 2260 2219 2264
rect 2311 2260 2315 2264
rect 2503 2257 2507 2261
rect 495 2251 499 2255
rect 1131 2251 1135 2255
rect 975 2243 979 2247
rect 1327 2240 1331 2244
rect 1471 2239 1475 2243
rect 111 2228 115 2232
rect 263 2229 267 2233
rect 319 2229 323 2233
rect 383 2229 387 2233
rect 447 2229 451 2233
rect 503 2229 507 2233
rect 511 2227 515 2231
rect 559 2229 563 2233
rect 583 2227 584 2231
rect 584 2227 587 2231
rect 615 2229 619 2233
rect 671 2229 675 2233
rect 727 2229 731 2233
rect 791 2229 795 2233
rect 855 2229 859 2233
rect 919 2229 923 2233
rect 983 2229 987 2233
rect 1047 2229 1051 2233
rect 1111 2229 1115 2233
rect 1131 2227 1132 2231
rect 1132 2227 1135 2231
rect 1287 2228 1291 2232
rect 1559 2239 1563 2243
rect 1655 2239 1659 2243
rect 1751 2239 1755 2243
rect 1855 2239 1859 2243
rect 1875 2239 1876 2243
rect 1876 2239 1879 2243
rect 1951 2239 1955 2243
rect 2047 2239 2051 2243
rect 2135 2239 2139 2243
rect 2231 2239 2235 2243
rect 2327 2239 2331 2243
rect 2335 2239 2339 2243
rect 2503 2240 2507 2244
rect 1587 2219 1591 2223
rect 2223 2219 2227 2223
rect 111 2211 115 2215
rect 247 2208 251 2212
rect 303 2208 307 2212
rect 367 2208 371 2212
rect 431 2208 435 2212
rect 487 2208 491 2212
rect 543 2208 547 2212
rect 599 2208 603 2212
rect 655 2208 659 2212
rect 711 2208 715 2212
rect 775 2208 779 2212
rect 839 2208 843 2212
rect 903 2208 907 2212
rect 967 2208 971 2212
rect 1031 2208 1035 2212
rect 1095 2208 1099 2212
rect 1287 2211 1291 2215
rect 1891 2207 1895 2211
rect 2335 2207 2339 2211
rect 359 2199 363 2203
rect 511 2199 515 2203
rect 111 2189 115 2193
rect 335 2192 339 2196
rect 391 2192 395 2196
rect 447 2192 451 2196
rect 503 2192 507 2196
rect 559 2192 563 2196
rect 1827 2199 1831 2203
rect 1287 2189 1291 2193
rect 1327 2184 1331 2188
rect 1567 2185 1571 2189
rect 1587 2183 1588 2187
rect 1588 2183 1591 2187
rect 1623 2185 1627 2189
rect 1679 2185 1683 2189
rect 1743 2185 1747 2189
rect 1807 2185 1811 2189
rect 1871 2185 1875 2189
rect 1891 2183 1892 2187
rect 1892 2183 1895 2187
rect 1927 2185 1931 2189
rect 1983 2185 1987 2189
rect 2039 2185 2043 2189
rect 2095 2185 2099 2189
rect 2159 2185 2163 2189
rect 2223 2185 2227 2189
rect 2287 2185 2291 2189
rect 2343 2185 2347 2189
rect 2399 2185 2403 2189
rect 2455 2185 2459 2189
rect 2471 2183 2475 2187
rect 2503 2184 2507 2188
rect 111 2172 115 2176
rect 351 2171 355 2175
rect 407 2171 411 2175
rect 463 2171 467 2175
rect 519 2171 523 2175
rect 575 2171 579 2175
rect 583 2171 587 2175
rect 1287 2172 1291 2176
rect 1327 2167 1331 2171
rect 1551 2164 1555 2168
rect 1607 2164 1611 2168
rect 1663 2164 1667 2168
rect 1727 2164 1731 2168
rect 1791 2164 1795 2168
rect 1855 2164 1859 2168
rect 1911 2164 1915 2168
rect 1967 2164 1971 2168
rect 2023 2164 2027 2168
rect 2079 2164 2083 2168
rect 2143 2164 2147 2168
rect 2207 2164 2211 2168
rect 2271 2164 2275 2168
rect 2327 2164 2331 2168
rect 2383 2164 2387 2168
rect 2439 2164 2443 2168
rect 2503 2167 2507 2171
rect 359 2155 360 2159
rect 360 2155 363 2159
rect 583 2143 587 2147
rect 1127 2143 1131 2147
rect 1327 2137 1331 2141
rect 1663 2140 1667 2144
rect 1719 2140 1723 2144
rect 1791 2140 1795 2144
rect 1871 2140 1875 2144
rect 1967 2140 1971 2144
rect 2079 2140 2083 2144
rect 2199 2140 2203 2144
rect 2327 2140 2331 2144
rect 2439 2140 2443 2144
rect 2503 2137 2507 2141
rect 111 2120 115 2124
rect 415 2121 419 2125
rect 511 2121 515 2125
rect 607 2121 611 2125
rect 711 2121 715 2125
rect 815 2121 819 2125
rect 823 2119 827 2123
rect 927 2121 931 2125
rect 1039 2121 1043 2125
rect 1151 2121 1155 2125
rect 1239 2121 1243 2125
rect 1255 2119 1259 2123
rect 1287 2120 1291 2124
rect 1327 2120 1331 2124
rect 1679 2119 1683 2123
rect 1735 2119 1739 2123
rect 1807 2119 1811 2123
rect 1827 2119 1828 2123
rect 1828 2119 1831 2123
rect 1887 2119 1891 2123
rect 1983 2119 1987 2123
rect 1991 2119 1995 2123
rect 2095 2119 2099 2123
rect 2215 2119 2219 2123
rect 2343 2119 2347 2123
rect 111 2103 115 2107
rect 399 2100 403 2104
rect 495 2100 499 2104
rect 591 2100 595 2104
rect 695 2100 699 2104
rect 799 2100 803 2104
rect 911 2100 915 2104
rect 1023 2100 1027 2104
rect 1135 2100 1139 2104
rect 1223 2100 1227 2104
rect 1287 2103 1291 2107
rect 2455 2119 2459 2123
rect 2463 2119 2467 2123
rect 2503 2120 2507 2124
rect 2335 2103 2339 2107
rect 1991 2095 1995 2099
rect 2471 2099 2475 2103
rect 111 2085 115 2089
rect 375 2088 379 2092
rect 447 2088 451 2092
rect 519 2088 523 2092
rect 599 2088 603 2092
rect 679 2088 683 2092
rect 759 2088 763 2092
rect 831 2088 835 2092
rect 903 2088 907 2092
rect 967 2088 971 2092
rect 1031 2088 1035 2092
rect 1103 2088 1107 2092
rect 1167 2088 1171 2092
rect 1223 2088 1227 2092
rect 1287 2085 1291 2089
rect 1859 2079 1863 2083
rect 111 2068 115 2072
rect 391 2067 395 2071
rect 455 2067 459 2071
rect 463 2067 467 2071
rect 479 2067 483 2071
rect 535 2067 539 2071
rect 615 2067 619 2071
rect 631 2067 635 2071
rect 695 2067 699 2071
rect 775 2067 779 2071
rect 823 2059 827 2063
rect 847 2067 851 2071
rect 919 2067 923 2071
rect 983 2067 987 2071
rect 1047 2067 1051 2071
rect 1119 2067 1123 2071
rect 1127 2067 1131 2071
rect 1183 2067 1187 2071
rect 1239 2067 1243 2071
rect 1287 2068 1291 2072
rect 2463 2071 2464 2075
rect 2464 2071 2467 2075
rect 479 2047 483 2051
rect 631 2047 635 2051
rect 1083 2047 1087 2051
rect 1327 2056 1331 2060
rect 1367 2057 1371 2061
rect 1423 2057 1427 2061
rect 1503 2057 1507 2061
rect 1591 2057 1595 2061
rect 1679 2057 1683 2061
rect 1687 2055 1691 2059
rect 1783 2057 1787 2061
rect 1895 2057 1899 2061
rect 2023 2057 2027 2061
rect 2167 2057 2171 2061
rect 2319 2057 2323 2061
rect 2335 2055 2339 2059
rect 2455 2057 2459 2061
rect 2471 2055 2475 2059
rect 2503 2056 2507 2060
rect 1255 2047 1259 2051
rect 659 2035 663 2039
rect 1327 2039 1331 2043
rect 1351 2036 1355 2040
rect 1407 2036 1411 2040
rect 1487 2036 1491 2040
rect 1575 2036 1579 2040
rect 1663 2036 1667 2040
rect 1767 2036 1771 2040
rect 1879 2036 1883 2040
rect 2007 2036 2011 2040
rect 2151 2036 2155 2040
rect 2303 2036 2307 2040
rect 2439 2036 2443 2040
rect 2503 2039 2507 2043
rect 455 2027 459 2031
rect 727 2027 728 2031
rect 728 2027 731 2031
rect 1327 2021 1331 2025
rect 1351 2024 1355 2028
rect 1423 2024 1427 2028
rect 1519 2024 1523 2028
rect 1615 2024 1619 2028
rect 1719 2024 1723 2028
rect 1823 2024 1827 2028
rect 1935 2024 1939 2028
rect 2055 2024 2059 2028
rect 2183 2024 2187 2028
rect 2319 2024 2323 2028
rect 2439 2024 2443 2028
rect 2503 2021 2507 2025
rect 111 2012 115 2016
rect 295 2013 299 2017
rect 375 2013 379 2017
rect 407 2011 411 2015
rect 463 2013 467 2017
rect 551 2013 555 2017
rect 639 2013 643 2017
rect 659 2011 660 2015
rect 660 2011 663 2015
rect 719 2013 723 2017
rect 799 2013 803 2017
rect 887 2013 891 2017
rect 975 2013 979 2017
rect 1063 2013 1067 2017
rect 1083 2011 1084 2015
rect 1084 2011 1087 2015
rect 1287 2012 1291 2016
rect 1327 2004 1331 2008
rect 1367 2003 1371 2007
rect 111 1995 115 1999
rect 279 1992 283 1996
rect 359 1992 363 1996
rect 447 1992 451 1996
rect 535 1992 539 1996
rect 623 1992 627 1996
rect 703 1992 707 1996
rect 783 1992 787 1996
rect 871 1992 875 1996
rect 959 1992 963 1996
rect 1047 1992 1051 1996
rect 1287 1995 1291 1999
rect 1439 2003 1443 2007
rect 1535 2003 1539 2007
rect 1631 2003 1635 2007
rect 1735 2003 1739 2007
rect 1743 2003 1747 2007
rect 1839 2003 1843 2007
rect 1859 2003 1860 2007
rect 1860 2003 1863 2007
rect 1951 2003 1955 2007
rect 1967 2003 1971 2007
rect 2071 2003 2075 2007
rect 2199 2003 2203 2007
rect 2115 1995 2119 1999
rect 2311 1995 2315 1999
rect 2335 2003 2339 2007
rect 2343 2003 2347 2007
rect 2455 2003 2459 2007
rect 2463 2003 2467 2007
rect 2503 2004 2507 2008
rect 1687 1983 1691 1987
rect 1967 1983 1971 1987
rect 2175 1987 2179 1991
rect 2471 1987 2475 1991
rect 111 1973 115 1977
rect 135 1976 139 1980
rect 207 1976 211 1980
rect 287 1976 291 1980
rect 383 1976 387 1980
rect 487 1976 491 1980
rect 591 1976 595 1980
rect 695 1976 699 1980
rect 799 1976 803 1980
rect 903 1976 907 1980
rect 1015 1976 1019 1980
rect 2343 1979 2347 1983
rect 1287 1973 1291 1977
rect 1743 1971 1747 1975
rect 2115 1971 2119 1975
rect 111 1956 115 1960
rect 151 1955 155 1959
rect 223 1955 227 1959
rect 303 1955 307 1959
rect 367 1955 371 1959
rect 399 1955 403 1959
rect 503 1955 507 1959
rect 607 1955 611 1959
rect 615 1955 619 1959
rect 711 1955 715 1959
rect 727 1955 731 1959
rect 815 1955 819 1959
rect 919 1955 923 1959
rect 1031 1955 1035 1959
rect 1039 1955 1043 1959
rect 1287 1956 1291 1960
rect 2247 1963 2251 1967
rect 2463 1963 2464 1967
rect 2464 1963 2467 1967
rect 2311 1955 2315 1959
rect 1327 1948 1331 1952
rect 1455 1949 1459 1953
rect 1543 1949 1547 1953
rect 1639 1949 1643 1953
rect 1735 1949 1739 1953
rect 1839 1949 1843 1953
rect 1847 1947 1851 1951
rect 1943 1949 1947 1953
rect 2047 1949 2051 1953
rect 2151 1949 2155 1953
rect 2175 1947 2176 1951
rect 2176 1947 2179 1951
rect 2255 1949 2259 1953
rect 2367 1949 2371 1953
rect 2455 1949 2459 1953
rect 2463 1947 2467 1951
rect 2503 1948 2507 1952
rect 407 1939 408 1943
rect 408 1939 411 1943
rect 615 1931 619 1935
rect 887 1939 891 1943
rect 1039 1931 1043 1935
rect 1327 1931 1331 1935
rect 1439 1928 1443 1932
rect 1527 1928 1531 1932
rect 1623 1928 1627 1932
rect 1719 1928 1723 1932
rect 1823 1928 1827 1932
rect 1927 1928 1931 1932
rect 2031 1928 2035 1932
rect 2135 1928 2139 1932
rect 2239 1928 2243 1932
rect 2351 1928 2355 1932
rect 2439 1928 2443 1932
rect 2503 1931 2507 1935
rect 703 1919 707 1923
rect 367 1911 371 1915
rect 1075 1911 1079 1915
rect 1327 1909 1331 1913
rect 1527 1912 1531 1916
rect 1615 1912 1619 1916
rect 1711 1912 1715 1916
rect 1815 1912 1819 1916
rect 1919 1912 1923 1916
rect 2015 1912 2019 1916
rect 2111 1912 2115 1916
rect 2199 1912 2203 1916
rect 2287 1912 2291 1916
rect 2375 1912 2379 1916
rect 2439 1912 2443 1916
rect 2503 1909 2507 1913
rect 111 1896 115 1900
rect 151 1897 155 1901
rect 199 1895 203 1899
rect 239 1897 243 1901
rect 375 1897 379 1901
rect 527 1897 531 1901
rect 687 1897 691 1901
rect 703 1895 707 1899
rect 863 1897 867 1901
rect 887 1895 888 1899
rect 888 1895 891 1899
rect 1039 1897 1043 1901
rect 1287 1896 1291 1900
rect 1327 1892 1331 1896
rect 1543 1891 1547 1895
rect 1631 1891 1635 1895
rect 1727 1891 1731 1895
rect 111 1879 115 1883
rect 135 1876 139 1880
rect 223 1876 227 1880
rect 359 1876 363 1880
rect 511 1876 515 1880
rect 671 1876 675 1880
rect 847 1876 851 1880
rect 1023 1876 1027 1880
rect 1287 1879 1291 1883
rect 1831 1891 1835 1895
rect 1935 1891 1939 1895
rect 1975 1891 1979 1895
rect 2031 1891 2035 1895
rect 2127 1891 2131 1895
rect 2215 1891 2219 1895
rect 2247 1891 2251 1895
rect 2303 1891 2307 1895
rect 2319 1891 2323 1895
rect 2391 1891 2395 1895
rect 2455 1891 2459 1895
rect 2487 1891 2491 1895
rect 2503 1892 2507 1896
rect 1847 1871 1851 1875
rect 2319 1871 2323 1875
rect 2463 1875 2464 1879
rect 2464 1875 2467 1879
rect 111 1861 115 1865
rect 135 1864 139 1868
rect 191 1864 195 1868
rect 263 1864 267 1868
rect 335 1864 339 1868
rect 407 1864 411 1868
rect 479 1864 483 1868
rect 551 1864 555 1868
rect 615 1864 619 1868
rect 679 1864 683 1868
rect 743 1864 747 1868
rect 815 1864 819 1868
rect 887 1864 891 1868
rect 959 1864 963 1868
rect 1039 1864 1043 1868
rect 1287 1861 1291 1865
rect 1803 1863 1807 1867
rect 2475 1867 2479 1871
rect 111 1844 115 1848
rect 151 1843 155 1847
rect 159 1843 163 1847
rect 207 1843 211 1847
rect 279 1843 283 1847
rect 351 1843 355 1847
rect 359 1843 363 1847
rect 423 1843 427 1847
rect 495 1843 499 1847
rect 567 1843 571 1847
rect 631 1843 635 1847
rect 695 1843 699 1847
rect 759 1843 763 1847
rect 831 1843 835 1847
rect 903 1843 907 1847
rect 975 1843 979 1847
rect 983 1843 987 1847
rect 1055 1843 1059 1847
rect 1075 1843 1076 1847
rect 1076 1843 1079 1847
rect 1287 1844 1291 1848
rect 1975 1855 1979 1859
rect 2167 1855 2171 1859
rect 1327 1840 1331 1844
rect 1535 1841 1539 1845
rect 1607 1841 1611 1845
rect 1687 1841 1691 1845
rect 1695 1839 1699 1843
rect 1783 1841 1787 1845
rect 1803 1839 1804 1843
rect 1804 1839 1807 1843
rect 1879 1841 1883 1845
rect 1983 1841 1987 1845
rect 2079 1841 2083 1845
rect 2175 1841 2179 1845
rect 2271 1841 2275 1845
rect 2367 1841 2371 1845
rect 2455 1841 2459 1845
rect 2475 1839 2476 1843
rect 2476 1839 2479 1843
rect 2503 1840 2507 1844
rect 199 1827 203 1831
rect 459 1827 463 1831
rect 1063 1827 1064 1831
rect 1064 1827 1067 1831
rect 359 1819 363 1823
rect 1327 1823 1331 1827
rect 1519 1820 1523 1824
rect 1591 1820 1595 1824
rect 1671 1820 1675 1824
rect 1767 1820 1771 1824
rect 1863 1820 1867 1824
rect 1967 1820 1971 1824
rect 2063 1820 2067 1824
rect 2159 1820 2163 1824
rect 2255 1820 2259 1824
rect 2351 1820 2355 1824
rect 2439 1820 2443 1824
rect 2503 1823 2507 1827
rect 651 1807 655 1811
rect 983 1807 987 1811
rect 159 1799 160 1803
rect 160 1799 163 1803
rect 499 1799 503 1803
rect 1139 1799 1143 1803
rect 1327 1801 1331 1805
rect 1463 1804 1467 1808
rect 1559 1804 1563 1808
rect 1663 1804 1667 1808
rect 1767 1804 1771 1808
rect 1879 1804 1883 1808
rect 1983 1804 1987 1808
rect 2087 1804 2091 1808
rect 2183 1804 2187 1808
rect 2271 1804 2275 1808
rect 2367 1804 2371 1808
rect 2439 1804 2443 1808
rect 2503 1801 2507 1805
rect 111 1784 115 1788
rect 151 1785 155 1789
rect 231 1785 235 1789
rect 335 1785 339 1789
rect 359 1783 360 1787
rect 360 1783 363 1787
rect 439 1785 443 1789
rect 459 1783 460 1787
rect 460 1783 463 1787
rect 535 1785 539 1789
rect 631 1785 635 1789
rect 651 1783 652 1787
rect 652 1783 655 1787
rect 719 1785 723 1789
rect 799 1785 803 1789
rect 879 1785 883 1789
rect 959 1785 963 1789
rect 999 1783 1003 1787
rect 1039 1785 1043 1789
rect 1063 1783 1064 1787
rect 1064 1783 1067 1787
rect 1119 1785 1123 1789
rect 1287 1784 1291 1788
rect 1327 1784 1331 1788
rect 1479 1783 1483 1787
rect 1559 1783 1563 1787
rect 1575 1783 1579 1787
rect 1679 1783 1683 1787
rect 1783 1783 1787 1787
rect 1895 1783 1899 1787
rect 1903 1783 1907 1787
rect 1999 1783 2003 1787
rect 2103 1783 2107 1787
rect 2199 1783 2203 1787
rect 2287 1783 2291 1787
rect 2383 1783 2387 1787
rect 2403 1783 2404 1787
rect 2404 1783 2407 1787
rect 2455 1783 2459 1787
rect 2463 1783 2467 1787
rect 2503 1784 2507 1788
rect 111 1767 115 1771
rect 135 1764 139 1768
rect 215 1764 219 1768
rect 319 1764 323 1768
rect 423 1764 427 1768
rect 519 1764 523 1768
rect 615 1764 619 1768
rect 703 1764 707 1768
rect 783 1764 787 1768
rect 863 1764 867 1768
rect 943 1764 947 1768
rect 1023 1764 1027 1768
rect 1103 1764 1107 1768
rect 1287 1767 1291 1771
rect 1695 1767 1699 1771
rect 1903 1759 1907 1763
rect 2371 1763 2375 1767
rect 2487 1767 2491 1771
rect 111 1745 115 1749
rect 135 1748 139 1752
rect 239 1748 243 1752
rect 351 1748 355 1752
rect 463 1748 467 1752
rect 575 1748 579 1752
rect 679 1748 683 1752
rect 783 1748 787 1752
rect 887 1748 891 1752
rect 991 1748 995 1752
rect 1103 1748 1107 1752
rect 1795 1751 1799 1755
rect 2343 1751 2347 1755
rect 1287 1745 1291 1749
rect 1559 1743 1563 1747
rect 2463 1743 2464 1747
rect 2464 1743 2467 1747
rect 111 1728 115 1732
rect 151 1727 155 1731
rect 183 1727 187 1731
rect 255 1727 259 1731
rect 367 1727 371 1731
rect 479 1727 483 1731
rect 499 1727 500 1731
rect 500 1727 503 1731
rect 591 1727 595 1731
rect 695 1727 699 1731
rect 735 1727 739 1731
rect 799 1727 803 1731
rect 903 1727 907 1731
rect 919 1727 923 1731
rect 1007 1727 1011 1731
rect 1119 1727 1123 1731
rect 1139 1727 1140 1731
rect 1140 1727 1143 1731
rect 1287 1728 1291 1732
rect 1327 1728 1331 1732
rect 1375 1729 1379 1733
rect 1439 1727 1443 1731
rect 1471 1729 1475 1733
rect 1567 1729 1571 1733
rect 1671 1729 1675 1733
rect 1775 1729 1779 1733
rect 1795 1727 1796 1731
rect 1796 1727 1799 1731
rect 1887 1729 1891 1733
rect 1999 1729 2003 1733
rect 2111 1729 2115 1733
rect 2231 1729 2235 1733
rect 2351 1729 2355 1733
rect 2371 1727 2372 1731
rect 2372 1727 2375 1731
rect 2455 1729 2459 1733
rect 2471 1727 2475 1731
rect 2503 1728 2507 1732
rect 359 1711 363 1715
rect 659 1711 663 1715
rect 919 1707 923 1711
rect 999 1711 1003 1715
rect 1195 1711 1199 1715
rect 1327 1711 1331 1715
rect 1359 1708 1363 1712
rect 1455 1708 1459 1712
rect 1551 1708 1555 1712
rect 1655 1708 1659 1712
rect 1759 1708 1763 1712
rect 1871 1708 1875 1712
rect 1983 1708 1987 1712
rect 2095 1708 2099 1712
rect 2215 1708 2219 1712
rect 2335 1708 2339 1712
rect 2439 1708 2443 1712
rect 2503 1711 2507 1715
rect 1327 1693 1331 1697
rect 1351 1696 1355 1700
rect 1431 1696 1435 1700
rect 1535 1696 1539 1700
rect 1647 1696 1651 1700
rect 1759 1696 1763 1700
rect 1879 1696 1883 1700
rect 2015 1696 2019 1700
rect 2159 1696 2163 1700
rect 2311 1696 2315 1700
rect 2439 1696 2443 1700
rect 2503 1693 2507 1697
rect 183 1687 187 1691
rect 447 1687 448 1691
rect 448 1687 451 1691
rect 735 1687 739 1691
rect 1091 1687 1095 1691
rect 111 1672 115 1676
rect 191 1673 195 1677
rect 271 1673 275 1677
rect 351 1673 355 1677
rect 359 1671 363 1675
rect 439 1673 443 1677
rect 535 1673 539 1677
rect 639 1673 643 1677
rect 659 1671 660 1675
rect 660 1671 663 1675
rect 743 1673 747 1677
rect 847 1673 851 1677
rect 951 1673 955 1677
rect 967 1671 971 1675
rect 1063 1673 1067 1677
rect 1175 1673 1179 1677
rect 1195 1671 1196 1675
rect 1196 1671 1199 1675
rect 1287 1672 1291 1676
rect 1327 1676 1331 1680
rect 1367 1675 1371 1679
rect 1375 1675 1379 1679
rect 1447 1675 1451 1679
rect 1551 1675 1555 1679
rect 1663 1675 1667 1679
rect 1671 1675 1675 1679
rect 1775 1675 1779 1679
rect 1895 1675 1899 1679
rect 2031 1675 2035 1679
rect 2175 1675 2179 1679
rect 2327 1675 2331 1679
rect 2343 1675 2347 1679
rect 2455 1675 2459 1679
rect 2463 1675 2467 1679
rect 2503 1676 2507 1680
rect 111 1655 115 1659
rect 175 1652 179 1656
rect 255 1652 259 1656
rect 335 1652 339 1656
rect 423 1652 427 1656
rect 519 1652 523 1656
rect 623 1652 627 1656
rect 727 1652 731 1656
rect 831 1652 835 1656
rect 935 1652 939 1656
rect 1047 1652 1051 1656
rect 1159 1652 1163 1656
rect 1287 1655 1291 1659
rect 1383 1659 1387 1663
rect 1439 1659 1443 1663
rect 2347 1655 2351 1659
rect 2471 1659 2475 1663
rect 111 1637 115 1641
rect 215 1640 219 1644
rect 271 1640 275 1644
rect 335 1640 339 1644
rect 407 1640 411 1644
rect 479 1640 483 1644
rect 559 1640 563 1644
rect 647 1640 651 1644
rect 743 1640 747 1644
rect 839 1640 843 1644
rect 943 1640 947 1644
rect 1055 1640 1059 1644
rect 1175 1640 1179 1644
rect 1287 1637 1291 1641
rect 2139 1639 2143 1643
rect 1375 1631 1376 1635
rect 1376 1631 1379 1635
rect 111 1620 115 1624
rect 231 1619 235 1623
rect 287 1619 291 1623
rect 295 1619 299 1623
rect 351 1619 355 1623
rect 423 1619 427 1623
rect 447 1619 448 1623
rect 448 1619 451 1623
rect 495 1619 499 1623
rect 575 1619 579 1623
rect 663 1619 667 1623
rect 359 1603 360 1607
rect 360 1603 363 1607
rect 759 1619 763 1623
rect 807 1619 811 1623
rect 855 1619 859 1623
rect 871 1619 875 1623
rect 959 1619 963 1623
rect 1071 1619 1075 1623
rect 1091 1619 1092 1623
rect 1092 1619 1095 1623
rect 1191 1619 1195 1623
rect 1287 1620 1291 1624
rect 2463 1631 2464 1635
rect 2464 1631 2467 1635
rect 1327 1616 1331 1620
rect 1367 1617 1371 1621
rect 1431 1617 1435 1621
rect 1519 1617 1523 1621
rect 1535 1615 1539 1619
rect 1599 1617 1603 1621
rect 1679 1617 1683 1621
rect 1751 1617 1755 1621
rect 1839 1617 1843 1621
rect 1935 1617 1939 1621
rect 2055 1617 2059 1621
rect 2183 1617 2187 1621
rect 2327 1617 2331 1621
rect 2347 1615 2348 1619
rect 2348 1615 2351 1619
rect 2455 1617 2459 1621
rect 2463 1615 2467 1619
rect 2503 1616 2507 1620
rect 527 1603 531 1607
rect 871 1599 875 1603
rect 967 1603 968 1607
rect 968 1603 971 1607
rect 1211 1603 1215 1607
rect 1327 1599 1331 1603
rect 1351 1596 1355 1600
rect 1415 1596 1419 1600
rect 1503 1596 1507 1600
rect 1583 1596 1587 1600
rect 1663 1596 1667 1600
rect 1735 1596 1739 1600
rect 1823 1596 1827 1600
rect 1919 1596 1923 1600
rect 2039 1596 2043 1600
rect 2167 1596 2171 1600
rect 2311 1596 2315 1600
rect 2439 1596 2443 1600
rect 2503 1599 2507 1603
rect 295 1583 296 1587
rect 296 1583 299 1587
rect 619 1583 623 1587
rect 807 1583 811 1587
rect 991 1583 995 1587
rect 1327 1577 1331 1581
rect 1351 1580 1355 1584
rect 1423 1580 1427 1584
rect 1527 1580 1531 1584
rect 1647 1580 1651 1584
rect 1783 1580 1787 1584
rect 1935 1580 1939 1584
rect 2103 1580 2107 1584
rect 2279 1580 2283 1584
rect 2439 1580 2443 1584
rect 2503 1577 2507 1581
rect 111 1568 115 1572
rect 287 1569 291 1573
rect 351 1569 355 1573
rect 423 1569 427 1573
rect 503 1569 507 1573
rect 527 1567 528 1571
rect 528 1567 531 1571
rect 599 1569 603 1573
rect 703 1569 707 1573
rect 743 1567 747 1571
rect 815 1569 819 1573
rect 935 1569 939 1573
rect 955 1567 956 1571
rect 956 1567 959 1571
rect 1063 1569 1067 1573
rect 1191 1569 1195 1573
rect 1211 1567 1212 1571
rect 1212 1567 1215 1571
rect 1287 1568 1291 1572
rect 1327 1560 1331 1564
rect 1367 1559 1371 1563
rect 1375 1559 1379 1563
rect 1439 1559 1443 1563
rect 111 1551 115 1555
rect 271 1548 275 1552
rect 335 1548 339 1552
rect 407 1548 411 1552
rect 487 1548 491 1552
rect 583 1548 587 1552
rect 687 1548 691 1552
rect 799 1548 803 1552
rect 919 1548 923 1552
rect 1047 1548 1051 1552
rect 1175 1548 1179 1552
rect 1287 1551 1291 1555
rect 1543 1559 1547 1563
rect 1663 1559 1667 1563
rect 1799 1559 1803 1563
rect 1951 1559 1955 1563
rect 2119 1559 2123 1563
rect 2139 1559 2140 1563
rect 2140 1559 2143 1563
rect 2295 1559 2299 1563
rect 2311 1559 2315 1563
rect 2455 1559 2459 1563
rect 2471 1559 2475 1563
rect 2503 1560 2507 1564
rect 1535 1543 1539 1547
rect 1875 1539 1879 1543
rect 2271 1543 2275 1547
rect 2311 1539 2315 1543
rect 2463 1543 2464 1547
rect 2464 1543 2467 1547
rect 111 1525 115 1529
rect 471 1528 475 1532
rect 551 1528 555 1532
rect 639 1528 643 1532
rect 735 1528 739 1532
rect 839 1528 843 1532
rect 951 1528 955 1532
rect 1063 1528 1067 1532
rect 1175 1528 1179 1532
rect 2363 1531 2367 1535
rect 1287 1525 1291 1529
rect 1375 1523 1376 1527
rect 1376 1523 1379 1527
rect 1655 1523 1656 1527
rect 1656 1523 1659 1527
rect 1471 1515 1475 1519
rect 2351 1523 2352 1527
rect 2352 1523 2355 1527
rect 2471 1523 2475 1527
rect 111 1508 115 1512
rect 487 1507 491 1511
rect 567 1507 571 1511
rect 655 1507 659 1511
rect 663 1507 667 1511
rect 751 1507 755 1511
rect 855 1507 859 1511
rect 871 1507 875 1511
rect 967 1507 971 1511
rect 991 1507 992 1511
rect 992 1507 995 1511
rect 1079 1507 1083 1511
rect 1095 1507 1099 1511
rect 1191 1507 1195 1511
rect 1287 1508 1291 1512
rect 1327 1508 1331 1512
rect 1367 1509 1371 1513
rect 1439 1509 1443 1513
rect 1543 1509 1547 1513
rect 1647 1509 1651 1513
rect 1751 1509 1755 1513
rect 1855 1509 1859 1513
rect 1875 1507 1876 1511
rect 1876 1507 1879 1511
rect 1959 1509 1963 1513
rect 2055 1509 2059 1513
rect 2143 1507 2147 1511
rect 2151 1509 2155 1513
rect 2247 1509 2251 1513
rect 2271 1507 2272 1511
rect 2272 1507 2275 1511
rect 2343 1509 2347 1513
rect 2363 1507 2364 1511
rect 2364 1507 2367 1511
rect 2439 1509 2443 1513
rect 2463 1507 2464 1511
rect 2464 1507 2467 1511
rect 2503 1508 2507 1512
rect 743 1491 747 1495
rect 871 1487 875 1491
rect 1095 1487 1099 1491
rect 1199 1491 1200 1495
rect 1200 1491 1203 1495
rect 1327 1491 1331 1495
rect 1351 1488 1355 1492
rect 1423 1488 1427 1492
rect 1527 1488 1531 1492
rect 1631 1488 1635 1492
rect 1735 1488 1739 1492
rect 1839 1488 1843 1492
rect 1943 1488 1947 1492
rect 2039 1488 2043 1492
rect 2135 1488 2139 1492
rect 2231 1488 2235 1492
rect 2327 1488 2331 1492
rect 2423 1488 2427 1492
rect 2503 1491 2507 1495
rect 663 1471 664 1475
rect 664 1471 667 1475
rect 771 1475 775 1479
rect 1123 1479 1127 1483
rect 1327 1469 1331 1473
rect 1351 1472 1355 1476
rect 1423 1472 1427 1476
rect 1519 1472 1523 1476
rect 1615 1472 1619 1476
rect 1711 1472 1715 1476
rect 1815 1472 1819 1476
rect 1927 1472 1931 1476
rect 2047 1472 2051 1476
rect 2175 1472 2179 1476
rect 2303 1472 2307 1476
rect 2439 1472 2443 1476
rect 2503 1469 2507 1473
rect 111 1456 115 1460
rect 375 1457 379 1461
rect 463 1457 467 1461
rect 559 1457 563 1461
rect 623 1455 627 1459
rect 655 1457 659 1461
rect 751 1457 755 1461
rect 771 1455 772 1459
rect 772 1455 775 1459
rect 855 1457 859 1461
rect 959 1457 963 1461
rect 1063 1457 1067 1461
rect 1167 1457 1171 1461
rect 1199 1455 1203 1459
rect 1287 1456 1291 1460
rect 1327 1452 1331 1456
rect 1367 1451 1371 1455
rect 1415 1451 1419 1455
rect 1439 1451 1443 1455
rect 1535 1451 1539 1455
rect 1631 1451 1635 1455
rect 1655 1451 1656 1455
rect 1656 1451 1659 1455
rect 1727 1451 1731 1455
rect 111 1439 115 1443
rect 359 1436 363 1440
rect 447 1436 451 1440
rect 543 1436 547 1440
rect 639 1436 643 1440
rect 735 1436 739 1440
rect 839 1436 843 1440
rect 943 1436 947 1440
rect 1047 1436 1051 1440
rect 1151 1436 1155 1440
rect 1287 1439 1291 1443
rect 1831 1451 1835 1455
rect 1839 1451 1843 1455
rect 1943 1451 1947 1455
rect 1959 1451 1963 1455
rect 2063 1451 2067 1455
rect 2191 1451 2195 1455
rect 2319 1451 2323 1455
rect 2351 1451 2355 1455
rect 2455 1451 2459 1455
rect 2471 1451 2475 1455
rect 2503 1452 2507 1456
rect 1471 1435 1475 1439
rect 1703 1435 1707 1439
rect 1959 1431 1963 1435
rect 2143 1435 2147 1439
rect 2255 1435 2259 1439
rect 2463 1435 2464 1439
rect 2464 1435 2467 1439
rect 111 1421 115 1425
rect 231 1424 235 1428
rect 319 1424 323 1428
rect 415 1424 419 1428
rect 511 1424 515 1428
rect 615 1424 619 1428
rect 711 1424 715 1428
rect 807 1424 811 1428
rect 895 1424 899 1428
rect 991 1424 995 1428
rect 1087 1424 1091 1428
rect 1287 1421 1291 1425
rect 1603 1419 1607 1423
rect 1839 1419 1843 1423
rect 111 1404 115 1408
rect 247 1403 251 1407
rect 335 1403 339 1407
rect 431 1403 435 1407
rect 503 1403 507 1407
rect 527 1403 531 1407
rect 543 1403 547 1407
rect 631 1403 635 1407
rect 727 1403 731 1407
rect 823 1403 827 1407
rect 911 1403 915 1407
rect 1007 1403 1011 1407
rect 1103 1403 1107 1407
rect 1123 1403 1124 1407
rect 1124 1403 1127 1407
rect 1287 1404 1291 1408
rect 1415 1411 1419 1415
rect 2359 1411 2360 1415
rect 2360 1411 2363 1415
rect 2471 1411 2475 1415
rect 1327 1396 1331 1400
rect 1367 1397 1371 1401
rect 1375 1395 1379 1399
rect 1423 1397 1427 1401
rect 1503 1397 1507 1401
rect 1591 1397 1595 1401
rect 1679 1397 1683 1401
rect 1703 1395 1704 1399
rect 1704 1395 1707 1399
rect 1775 1397 1779 1401
rect 1879 1397 1883 1401
rect 1991 1397 1995 1401
rect 2111 1397 2115 1401
rect 2119 1395 2123 1399
rect 2231 1397 2235 1401
rect 2255 1395 2256 1399
rect 2256 1395 2259 1399
rect 2351 1397 2355 1401
rect 2455 1397 2459 1401
rect 2463 1395 2467 1399
rect 2503 1396 2507 1400
rect 543 1383 547 1387
rect 623 1387 627 1391
rect 1023 1383 1027 1387
rect 903 1375 907 1379
rect 1327 1379 1331 1383
rect 1351 1376 1355 1380
rect 1407 1376 1411 1380
rect 1487 1376 1491 1380
rect 1575 1376 1579 1380
rect 1663 1376 1667 1380
rect 1759 1376 1763 1380
rect 1863 1376 1867 1380
rect 1975 1376 1979 1380
rect 2095 1376 2099 1380
rect 2215 1376 2219 1380
rect 2335 1376 2339 1380
rect 2439 1376 2443 1380
rect 2503 1379 2507 1383
rect 503 1367 507 1371
rect 111 1352 115 1356
rect 151 1353 155 1357
rect 159 1351 163 1355
rect 215 1353 219 1357
rect 311 1353 315 1357
rect 407 1353 411 1357
rect 511 1353 515 1357
rect 607 1353 611 1357
rect 703 1353 707 1357
rect 799 1353 803 1357
rect 895 1353 899 1357
rect 1327 1357 1331 1361
rect 1351 1360 1355 1364
rect 1407 1360 1411 1364
rect 1479 1360 1483 1364
rect 1567 1360 1571 1364
rect 1655 1360 1659 1364
rect 1751 1360 1755 1364
rect 1855 1360 1859 1364
rect 1967 1360 1971 1364
rect 2079 1360 2083 1364
rect 2199 1360 2203 1364
rect 2327 1360 2331 1364
rect 2439 1360 2443 1364
rect 999 1353 1003 1357
rect 2503 1357 2507 1361
rect 1023 1351 1024 1355
rect 1024 1351 1027 1355
rect 1287 1352 1291 1356
rect 1327 1340 1331 1344
rect 111 1335 115 1339
rect 1367 1339 1371 1343
rect 135 1332 139 1336
rect 199 1332 203 1336
rect 295 1332 299 1336
rect 391 1332 395 1336
rect 495 1332 499 1336
rect 591 1332 595 1336
rect 687 1332 691 1336
rect 783 1332 787 1336
rect 879 1332 883 1336
rect 983 1332 987 1336
rect 1287 1335 1291 1339
rect 1423 1339 1427 1343
rect 1495 1339 1499 1343
rect 1527 1339 1531 1343
rect 1583 1339 1587 1343
rect 1603 1339 1604 1343
rect 1604 1339 1607 1343
rect 1671 1339 1675 1343
rect 1767 1339 1771 1343
rect 1871 1339 1875 1343
rect 111 1317 115 1321
rect 135 1320 139 1324
rect 215 1320 219 1324
rect 319 1320 323 1324
rect 415 1320 419 1324
rect 511 1320 515 1324
rect 599 1320 603 1324
rect 687 1320 691 1324
rect 783 1320 787 1324
rect 879 1320 883 1324
rect 1375 1323 1376 1327
rect 1376 1323 1379 1327
rect 1983 1339 1987 1343
rect 2095 1339 2099 1343
rect 2215 1339 2219 1343
rect 2223 1339 2227 1343
rect 2343 1339 2347 1343
rect 2359 1339 2363 1343
rect 2455 1339 2459 1343
rect 2471 1339 2475 1343
rect 2503 1340 2507 1344
rect 1743 1323 1747 1327
rect 1287 1317 1291 1321
rect 2119 1319 2123 1323
rect 2351 1323 2352 1327
rect 2352 1323 2355 1327
rect 2463 1323 2464 1327
rect 2464 1323 2467 1327
rect 111 1300 115 1304
rect 151 1299 155 1303
rect 231 1299 235 1303
rect 335 1299 339 1303
rect 431 1299 435 1303
rect 447 1299 451 1303
rect 527 1299 531 1303
rect 615 1299 619 1303
rect 703 1299 707 1303
rect 799 1299 803 1303
rect 895 1299 899 1303
rect 903 1299 907 1303
rect 1287 1300 1291 1304
rect 1843 1303 1847 1307
rect 2223 1303 2227 1307
rect 2471 1303 2475 1307
rect 159 1283 160 1287
rect 160 1283 163 1287
rect 1247 1287 1251 1291
rect 1527 1295 1528 1299
rect 1528 1295 1531 1299
rect 1851 1295 1855 1299
rect 2411 1287 2415 1291
rect 1115 1279 1119 1283
rect 1327 1280 1331 1284
rect 1367 1281 1371 1285
rect 1423 1281 1427 1285
rect 1519 1281 1523 1285
rect 1615 1281 1619 1285
rect 1719 1281 1723 1285
rect 1743 1279 1744 1283
rect 1744 1279 1747 1283
rect 1823 1281 1827 1285
rect 1843 1279 1844 1283
rect 1844 1279 1847 1283
rect 1919 1281 1923 1285
rect 2015 1281 2019 1285
rect 2103 1281 2107 1285
rect 2183 1281 2187 1285
rect 2255 1281 2259 1285
rect 2263 1279 2267 1283
rect 2327 1281 2331 1285
rect 2351 1279 2352 1283
rect 2352 1279 2355 1283
rect 2399 1281 2403 1285
rect 2455 1281 2459 1285
rect 2463 1279 2467 1283
rect 2503 1280 2507 1284
rect 447 1271 451 1275
rect 655 1263 659 1267
rect 1247 1263 1248 1267
rect 1248 1263 1251 1267
rect 1327 1263 1331 1267
rect 1351 1260 1355 1264
rect 1407 1260 1411 1264
rect 1503 1260 1507 1264
rect 1599 1260 1603 1264
rect 1703 1260 1707 1264
rect 1807 1260 1811 1264
rect 1903 1260 1907 1264
rect 1999 1260 2003 1264
rect 2087 1260 2091 1264
rect 2167 1260 2171 1264
rect 2239 1260 2243 1264
rect 2311 1260 2315 1264
rect 2383 1260 2387 1264
rect 2439 1260 2443 1264
rect 2503 1263 2507 1267
rect 111 1248 115 1252
rect 191 1249 195 1253
rect 247 1249 251 1253
rect 303 1249 307 1253
rect 367 1249 371 1253
rect 439 1249 443 1253
rect 527 1249 531 1253
rect 551 1247 552 1251
rect 552 1247 555 1251
rect 639 1249 643 1253
rect 775 1249 779 1253
rect 927 1249 931 1253
rect 1095 1249 1099 1253
rect 1115 1247 1116 1251
rect 1116 1247 1119 1251
rect 1239 1249 1243 1253
rect 1279 1247 1283 1251
rect 1287 1248 1291 1252
rect 111 1231 115 1235
rect 175 1228 179 1232
rect 231 1228 235 1232
rect 287 1228 291 1232
rect 351 1228 355 1232
rect 423 1228 427 1232
rect 511 1228 515 1232
rect 623 1228 627 1232
rect 759 1228 763 1232
rect 911 1228 915 1232
rect 1079 1228 1083 1232
rect 1223 1228 1227 1232
rect 1287 1231 1291 1235
rect 1327 1229 1331 1233
rect 1351 1232 1355 1236
rect 1447 1232 1451 1236
rect 1575 1232 1579 1236
rect 1695 1232 1699 1236
rect 1815 1232 1819 1236
rect 1927 1232 1931 1236
rect 2031 1232 2035 1236
rect 2127 1232 2131 1236
rect 2215 1232 2219 1236
rect 2295 1232 2299 1236
rect 2375 1232 2379 1236
rect 2439 1232 2443 1236
rect 2503 1229 2507 1233
rect 111 1213 115 1217
rect 351 1216 355 1220
rect 407 1216 411 1220
rect 463 1216 467 1220
rect 519 1216 523 1220
rect 575 1216 579 1220
rect 631 1216 635 1220
rect 687 1216 691 1220
rect 743 1216 747 1220
rect 799 1216 803 1220
rect 855 1216 859 1220
rect 911 1216 915 1220
rect 1287 1213 1291 1217
rect 1327 1212 1331 1216
rect 1367 1211 1371 1215
rect 1463 1211 1467 1215
rect 1479 1211 1483 1215
rect 1591 1211 1595 1215
rect 1279 1203 1283 1207
rect 1711 1211 1715 1215
rect 1831 1211 1835 1215
rect 1851 1211 1852 1215
rect 1852 1211 1855 1215
rect 1943 1211 1947 1215
rect 2047 1211 2051 1215
rect 2143 1211 2147 1215
rect 2231 1211 2235 1215
rect 2311 1211 2315 1215
rect 2375 1211 2379 1215
rect 2391 1211 2395 1215
rect 2411 1211 2412 1215
rect 2412 1211 2415 1215
rect 2455 1211 2459 1215
rect 2471 1211 2475 1215
rect 2503 1212 2507 1216
rect 111 1196 115 1200
rect 367 1195 371 1199
rect 423 1195 427 1199
rect 479 1195 483 1199
rect 535 1195 539 1199
rect 591 1195 595 1199
rect 639 1195 643 1199
rect 647 1195 651 1199
rect 655 1195 659 1199
rect 703 1195 707 1199
rect 759 1195 763 1199
rect 775 1195 779 1199
rect 815 1195 819 1199
rect 871 1195 875 1199
rect 887 1195 891 1199
rect 927 1195 931 1199
rect 1287 1196 1291 1200
rect 1755 1191 1759 1195
rect 1951 1195 1952 1199
rect 1952 1195 1955 1199
rect 2435 1195 2439 1199
rect 2463 1195 2464 1199
rect 2464 1195 2467 1199
rect 551 1175 555 1179
rect 775 1175 779 1179
rect 887 1175 891 1179
rect 895 1179 899 1183
rect 1479 1183 1483 1187
rect 2211 1183 2215 1187
rect 723 1163 727 1167
rect 1003 1163 1007 1167
rect 1855 1175 1859 1179
rect 2375 1175 2379 1179
rect 2479 1175 2483 1179
rect 2435 1167 2439 1171
rect 639 1155 643 1159
rect 1327 1160 1331 1164
rect 1367 1161 1371 1165
rect 1471 1161 1475 1165
rect 1599 1161 1603 1165
rect 887 1155 891 1159
rect 1607 1159 1611 1163
rect 1735 1161 1739 1165
rect 1755 1159 1756 1163
rect 1756 1159 1759 1163
rect 1863 1161 1867 1165
rect 1983 1161 1987 1165
rect 2087 1161 2091 1165
rect 2167 1159 2171 1163
rect 2191 1161 2195 1165
rect 2211 1159 2212 1163
rect 2212 1159 2215 1163
rect 2287 1161 2291 1165
rect 2383 1161 2387 1165
rect 2455 1161 2459 1165
rect 2503 1160 2507 1164
rect 111 1140 115 1144
rect 423 1141 427 1145
rect 479 1141 483 1145
rect 535 1141 539 1145
rect 583 1139 587 1143
rect 591 1141 595 1145
rect 647 1141 651 1145
rect 703 1141 707 1145
rect 723 1139 724 1143
rect 724 1139 727 1143
rect 759 1141 763 1145
rect 815 1141 819 1145
rect 871 1141 875 1145
rect 895 1139 896 1143
rect 896 1139 899 1143
rect 927 1141 931 1145
rect 983 1141 987 1145
rect 1003 1139 1004 1143
rect 1004 1139 1007 1143
rect 1287 1140 1291 1144
rect 1327 1143 1331 1147
rect 1351 1140 1355 1144
rect 1455 1140 1459 1144
rect 1583 1140 1587 1144
rect 1719 1140 1723 1144
rect 1847 1140 1851 1144
rect 1967 1140 1971 1144
rect 2071 1140 2075 1144
rect 2175 1140 2179 1144
rect 2271 1140 2275 1144
rect 2367 1140 2371 1144
rect 2439 1140 2443 1144
rect 2503 1143 2507 1147
rect 111 1123 115 1127
rect 407 1120 411 1124
rect 463 1120 467 1124
rect 519 1120 523 1124
rect 575 1120 579 1124
rect 631 1120 635 1124
rect 687 1120 691 1124
rect 743 1120 747 1124
rect 799 1120 803 1124
rect 855 1120 859 1124
rect 911 1120 915 1124
rect 967 1120 971 1124
rect 1287 1123 1291 1127
rect 1327 1121 1331 1125
rect 1367 1124 1371 1128
rect 1447 1124 1451 1128
rect 1535 1124 1539 1128
rect 1631 1124 1635 1128
rect 1719 1124 1723 1128
rect 1807 1124 1811 1128
rect 1895 1124 1899 1128
rect 1983 1124 1987 1128
rect 2071 1124 2075 1128
rect 2159 1124 2163 1128
rect 2255 1124 2259 1128
rect 2359 1124 2363 1128
rect 2439 1124 2443 1128
rect 2503 1121 2507 1125
rect 111 1101 115 1105
rect 223 1104 227 1108
rect 311 1104 315 1108
rect 399 1104 403 1108
rect 495 1104 499 1108
rect 591 1104 595 1108
rect 679 1104 683 1108
rect 767 1104 771 1108
rect 847 1104 851 1108
rect 927 1104 931 1108
rect 1015 1104 1019 1108
rect 1103 1104 1107 1108
rect 1287 1101 1291 1105
rect 1327 1104 1331 1108
rect 1383 1103 1387 1107
rect 1423 1103 1427 1107
rect 1463 1103 1467 1107
rect 1479 1103 1483 1107
rect 1551 1103 1555 1107
rect 1647 1103 1651 1107
rect 1735 1103 1739 1107
rect 1823 1103 1827 1107
rect 1855 1103 1859 1107
rect 1911 1103 1915 1107
rect 1999 1103 2003 1107
rect 2087 1103 2091 1107
rect 2119 1103 2123 1107
rect 2175 1103 2179 1107
rect 2271 1103 2275 1107
rect 2375 1103 2379 1107
rect 2383 1103 2387 1107
rect 2455 1103 2459 1107
rect 2463 1103 2467 1107
rect 2503 1104 2507 1108
rect 111 1084 115 1088
rect 239 1083 243 1087
rect 327 1083 331 1087
rect 415 1083 419 1087
rect 423 1083 427 1087
rect 511 1083 515 1087
rect 527 1083 531 1087
rect 607 1083 611 1087
rect 695 1083 699 1087
rect 783 1083 787 1087
rect 863 1083 867 1087
rect 887 1083 888 1087
rect 888 1083 891 1087
rect 943 1083 947 1087
rect 1031 1083 1035 1087
rect 527 1063 531 1067
rect 583 1067 587 1071
rect 1119 1083 1123 1087
rect 1127 1083 1131 1087
rect 1287 1084 1291 1088
rect 1479 1083 1483 1087
rect 1607 1087 1611 1091
rect 1787 1083 1791 1087
rect 1959 1087 1963 1091
rect 2167 1087 2171 1091
rect 2471 1087 2475 1091
rect 1007 1067 1011 1071
rect 2367 1067 2371 1071
rect 1127 1059 1131 1063
rect 1423 1059 1427 1063
rect 675 1051 679 1055
rect 799 1051 803 1055
rect 1711 1059 1712 1063
rect 1712 1059 1715 1063
rect 2119 1059 2120 1063
rect 2120 1059 2123 1063
rect 2463 1059 2464 1063
rect 2464 1059 2467 1063
rect 423 1043 424 1047
rect 424 1043 427 1047
rect 775 1043 776 1047
rect 776 1043 779 1047
rect 1327 1044 1331 1048
rect 1431 1045 1435 1049
rect 1495 1045 1499 1049
rect 1567 1045 1571 1049
rect 1639 1045 1643 1049
rect 1647 1043 1651 1047
rect 1703 1045 1707 1049
rect 1767 1045 1771 1049
rect 1787 1043 1788 1047
rect 1788 1043 1791 1047
rect 1839 1045 1843 1049
rect 1919 1045 1923 1049
rect 2007 1045 2011 1049
rect 2015 1043 2019 1047
rect 2111 1045 2115 1049
rect 2231 1045 2235 1049
rect 2351 1045 2355 1049
rect 2367 1043 2371 1047
rect 2455 1045 2459 1049
rect 2463 1043 2467 1047
rect 2503 1044 2507 1048
rect 111 1028 115 1032
rect 151 1029 155 1033
rect 207 1029 211 1033
rect 303 1029 307 1033
rect 335 1027 339 1031
rect 415 1029 419 1033
rect 535 1029 539 1033
rect 655 1029 659 1033
rect 675 1027 676 1031
rect 676 1027 679 1031
rect 767 1029 771 1033
rect 879 1029 883 1033
rect 983 1029 987 1033
rect 1007 1027 1008 1031
rect 1008 1027 1011 1031
rect 1095 1029 1099 1033
rect 1207 1029 1211 1033
rect 1227 1027 1228 1031
rect 1228 1027 1231 1031
rect 1287 1028 1291 1032
rect 1327 1027 1331 1031
rect 1415 1024 1419 1028
rect 1479 1024 1483 1028
rect 1551 1024 1555 1028
rect 1623 1024 1627 1028
rect 1687 1024 1691 1028
rect 1751 1024 1755 1028
rect 1823 1024 1827 1028
rect 1903 1024 1907 1028
rect 1991 1024 1995 1028
rect 2095 1024 2099 1028
rect 2215 1024 2219 1028
rect 2335 1024 2339 1028
rect 2439 1024 2443 1028
rect 2503 1027 2507 1031
rect 111 1011 115 1015
rect 135 1008 139 1012
rect 191 1008 195 1012
rect 287 1008 291 1012
rect 399 1008 403 1012
rect 519 1008 523 1012
rect 639 1008 643 1012
rect 751 1008 755 1012
rect 863 1008 867 1012
rect 967 1008 971 1012
rect 1079 1008 1083 1012
rect 1191 1008 1195 1012
rect 1287 1011 1291 1015
rect 1327 1001 1331 1005
rect 1511 1004 1515 1008
rect 1567 1004 1571 1008
rect 1623 1004 1627 1008
rect 1679 1004 1683 1008
rect 1735 1004 1739 1008
rect 1807 1004 1811 1008
rect 1887 1004 1891 1008
rect 1983 1004 1987 1008
rect 2095 1004 2099 1008
rect 2215 1004 2219 1008
rect 2335 1004 2339 1008
rect 2439 1004 2443 1008
rect 2503 1001 2507 1005
rect 111 989 115 993
rect 135 992 139 996
rect 215 992 219 996
rect 327 992 331 996
rect 439 992 443 996
rect 551 992 555 996
rect 663 992 667 996
rect 759 992 763 996
rect 847 992 851 996
rect 935 992 939 996
rect 1015 992 1019 996
rect 1087 992 1091 996
rect 1167 992 1171 996
rect 1223 992 1227 996
rect 1287 989 1291 993
rect 1327 984 1331 988
rect 1527 983 1531 987
rect 1535 983 1539 987
rect 1583 983 1587 987
rect 1599 983 1603 987
rect 1639 983 1643 987
rect 1695 983 1699 987
rect 1711 983 1715 987
rect 1751 983 1755 987
rect 1783 983 1787 987
rect 1823 983 1827 987
rect 1903 983 1907 987
rect 1999 983 2003 987
rect 2111 983 2115 987
rect 111 972 115 976
rect 151 971 155 975
rect 159 971 163 975
rect 231 971 235 975
rect 343 971 347 975
rect 455 971 459 975
rect 567 971 571 975
rect 575 971 579 975
rect 679 971 683 975
rect 775 971 779 975
rect 799 971 800 975
rect 800 971 803 975
rect 863 971 867 975
rect 919 971 923 975
rect 951 971 955 975
rect 1031 971 1035 975
rect 1047 971 1051 975
rect 1103 971 1107 975
rect 1183 971 1187 975
rect 335 955 339 959
rect 1239 971 1243 975
rect 1247 971 1251 975
rect 1287 972 1291 976
rect 1599 963 1603 967
rect 1647 967 1648 971
rect 1648 967 1651 971
rect 1655 967 1659 971
rect 2007 973 2011 975
rect 2007 971 2008 973
rect 2008 971 2011 973
rect 2231 983 2235 987
rect 2247 983 2251 987
rect 2351 983 2355 987
rect 2431 983 2435 987
rect 2455 983 2459 987
rect 2479 983 2480 987
rect 2480 983 2483 987
rect 2503 984 2507 988
rect 2247 963 2251 967
rect 2447 967 2451 971
rect 2463 967 2464 971
rect 2464 967 2467 971
rect 855 955 859 959
rect 575 947 579 951
rect 1047 951 1051 955
rect 1191 955 1192 959
rect 1192 955 1195 959
rect 767 943 771 947
rect 1247 947 1251 951
rect 159 935 160 939
rect 160 935 163 939
rect 535 935 539 939
rect 431 927 435 931
rect 919 935 923 939
rect 1247 935 1248 939
rect 1248 935 1251 939
rect 1263 935 1267 939
rect 1535 939 1539 943
rect 111 920 115 924
rect 151 921 155 925
rect 207 921 211 925
rect 295 921 299 925
rect 399 921 403 925
rect 511 921 515 925
rect 535 919 536 923
rect 536 919 539 923
rect 623 921 627 925
rect 735 921 739 925
rect 831 921 835 925
rect 855 919 856 923
rect 856 919 859 923
rect 927 921 931 925
rect 1015 921 1019 925
rect 1095 921 1099 925
rect 1119 919 1120 923
rect 1120 919 1123 923
rect 1175 921 1179 925
rect 1191 919 1195 923
rect 1239 921 1243 925
rect 1263 919 1264 923
rect 1264 919 1267 923
rect 1287 920 1291 924
rect 1723 931 1727 935
rect 1783 931 1787 935
rect 2407 931 2411 935
rect 1327 916 1331 920
rect 1367 917 1371 921
rect 1439 917 1443 921
rect 1527 917 1531 921
rect 1567 915 1571 919
rect 1615 917 1619 921
rect 1655 915 1659 919
rect 1695 917 1699 921
rect 1791 917 1795 921
rect 1895 917 1899 921
rect 2015 917 2019 921
rect 2151 917 2155 921
rect 2295 917 2299 921
rect 2303 915 2307 919
rect 2439 917 2443 921
rect 2447 915 2451 919
rect 2503 916 2507 920
rect 111 903 115 907
rect 135 900 139 904
rect 191 900 195 904
rect 279 900 283 904
rect 383 900 387 904
rect 495 900 499 904
rect 607 900 611 904
rect 719 900 723 904
rect 815 900 819 904
rect 911 900 915 904
rect 999 900 1003 904
rect 1079 900 1083 904
rect 1159 900 1163 904
rect 1223 900 1227 904
rect 1287 903 1291 907
rect 1327 899 1331 903
rect 1351 896 1355 900
rect 1423 896 1427 900
rect 1511 896 1515 900
rect 1599 896 1603 900
rect 1679 896 1683 900
rect 1775 896 1779 900
rect 1879 896 1883 900
rect 1999 896 2003 900
rect 2135 896 2139 900
rect 2279 896 2283 900
rect 2423 896 2427 900
rect 2503 899 2507 903
rect 111 881 115 885
rect 247 884 251 888
rect 343 884 347 888
rect 439 884 443 888
rect 543 884 547 888
rect 647 884 651 888
rect 743 884 747 888
rect 839 884 843 888
rect 927 884 931 888
rect 1007 884 1011 888
rect 1087 884 1091 888
rect 1167 884 1171 888
rect 1223 884 1227 888
rect 1287 881 1291 885
rect 1327 873 1331 877
rect 1487 876 1491 880
rect 1559 876 1563 880
rect 1623 876 1627 880
rect 1687 876 1691 880
rect 1751 876 1755 880
rect 1815 876 1819 880
rect 1887 876 1891 880
rect 1975 876 1979 880
rect 2079 876 2083 880
rect 2199 876 2203 880
rect 2319 876 2323 880
rect 2439 876 2443 880
rect 2503 873 2507 877
rect 111 864 115 868
rect 263 863 267 867
rect 359 863 363 867
rect 455 863 459 867
rect 559 863 563 867
rect 663 863 667 867
rect 671 863 675 867
rect 759 863 763 867
rect 767 863 771 867
rect 855 863 859 867
rect 943 863 947 867
rect 1023 863 1027 867
rect 1103 863 1107 867
rect 1183 863 1187 867
rect 1239 863 1243 867
rect 1247 863 1251 867
rect 1287 864 1291 868
rect 1327 856 1331 860
rect 1503 855 1507 859
rect 1519 855 1523 859
rect 1575 855 1579 859
rect 431 843 435 847
rect 1119 843 1123 847
rect 1639 855 1643 859
rect 1647 855 1651 859
rect 1703 855 1707 859
rect 1723 855 1724 859
rect 1724 855 1727 859
rect 1767 855 1771 859
rect 1831 855 1835 859
rect 1903 855 1907 859
rect 1991 855 1995 859
rect 2095 855 2099 859
rect 2215 855 2219 859
rect 2335 855 2339 859
rect 2343 855 2347 859
rect 2455 855 2459 859
rect 2463 855 2467 859
rect 2503 856 2507 860
rect 403 831 407 835
rect 1091 835 1095 839
rect 1567 839 1571 843
rect 1819 839 1823 843
rect 1839 839 1840 843
rect 1840 839 1843 843
rect 2431 839 2435 843
rect 1647 831 1651 835
rect 671 823 675 827
rect 763 823 767 827
rect 1519 819 1523 823
rect 1723 819 1727 823
rect 2343 819 2347 823
rect 111 808 115 812
rect 239 809 243 813
rect 303 809 307 813
rect 351 807 355 811
rect 383 809 387 813
rect 403 807 404 811
rect 404 807 407 811
rect 463 809 467 813
rect 551 809 555 813
rect 639 809 643 813
rect 727 809 731 813
rect 807 809 811 813
rect 895 809 899 813
rect 983 809 987 813
rect 1071 809 1075 813
rect 1091 807 1092 811
rect 1092 807 1095 811
rect 1287 808 1291 812
rect 1819 803 1823 807
rect 2391 811 2392 815
rect 2392 811 2395 815
rect 2463 811 2464 815
rect 2464 811 2467 815
rect 1327 796 1331 800
rect 1439 797 1443 801
rect 1511 797 1515 801
rect 1591 797 1595 801
rect 111 791 115 795
rect 1599 795 1603 799
rect 223 788 227 792
rect 287 788 291 792
rect 367 788 371 792
rect 447 788 451 792
rect 535 788 539 792
rect 623 788 627 792
rect 711 788 715 792
rect 791 788 795 792
rect 879 788 883 792
rect 967 788 971 792
rect 1055 788 1059 792
rect 1287 791 1291 795
rect 1671 797 1675 801
rect 1759 797 1763 801
rect 1847 797 1851 801
rect 1935 797 1939 801
rect 2023 797 2027 801
rect 2111 797 2115 801
rect 2199 797 2203 801
rect 2287 797 2291 801
rect 2295 795 2299 799
rect 2383 797 2387 801
rect 2407 795 2408 799
rect 2408 795 2411 799
rect 2455 797 2459 801
rect 2471 795 2475 799
rect 2503 796 2507 800
rect 763 779 767 783
rect 1011 779 1015 783
rect 1327 779 1331 783
rect 111 769 115 773
rect 151 772 155 776
rect 247 772 251 776
rect 343 772 347 776
rect 439 772 443 776
rect 527 772 531 776
rect 607 772 611 776
rect 679 772 683 776
rect 751 772 755 776
rect 823 772 827 776
rect 895 772 899 776
rect 975 772 979 776
rect 1423 776 1427 780
rect 1495 776 1499 780
rect 1575 776 1579 780
rect 1655 776 1659 780
rect 1743 776 1747 780
rect 1831 776 1835 780
rect 1919 776 1923 780
rect 2007 776 2011 780
rect 2095 776 2099 780
rect 2183 776 2187 780
rect 2271 776 2275 780
rect 2367 776 2371 780
rect 2439 776 2443 780
rect 2503 779 2507 783
rect 1287 769 1291 773
rect 1327 757 1331 761
rect 1351 760 1355 764
rect 1447 760 1451 764
rect 1567 760 1571 764
rect 1687 760 1691 764
rect 1807 760 1811 764
rect 1927 760 1931 764
rect 2039 760 2043 764
rect 2143 760 2147 764
rect 2247 760 2251 764
rect 2351 760 2355 764
rect 2439 760 2443 764
rect 2503 757 2507 761
rect 111 752 115 756
rect 167 751 171 755
rect 183 751 187 755
rect 263 751 267 755
rect 279 751 283 755
rect 359 751 363 755
rect 455 751 459 755
rect 543 751 547 755
rect 567 751 568 755
rect 568 751 571 755
rect 623 751 627 755
rect 695 751 699 755
rect 767 751 771 755
rect 839 751 843 755
rect 911 751 915 755
rect 991 751 995 755
rect 1011 751 1012 755
rect 1012 751 1015 755
rect 1287 752 1291 756
rect 279 731 283 735
rect 351 735 355 739
rect 375 735 379 739
rect 1327 740 1331 744
rect 1367 739 1371 743
rect 1375 739 1379 743
rect 1463 739 1467 743
rect 1583 739 1587 743
rect 931 731 935 735
rect 1703 739 1707 743
rect 1723 739 1724 743
rect 1724 739 1727 743
rect 1823 739 1827 743
rect 1943 739 1947 743
rect 2055 739 2059 743
rect 2159 739 2163 743
rect 2263 739 2267 743
rect 2271 739 2275 743
rect 2367 739 2371 743
rect 2391 739 2392 743
rect 2392 739 2395 743
rect 2455 739 2459 743
rect 2463 739 2467 743
rect 2503 740 2507 744
rect 595 719 599 723
rect 1599 723 1603 727
rect 1883 723 1887 727
rect 2295 719 2299 723
rect 2411 723 2415 727
rect 2471 723 2475 727
rect 183 711 184 715
rect 184 711 187 715
rect 311 711 315 715
rect 567 711 571 715
rect 631 711 635 715
rect 111 696 115 700
rect 175 697 179 701
rect 223 695 227 699
rect 263 697 267 701
rect 343 697 347 701
rect 375 695 379 699
rect 423 697 427 701
rect 503 697 507 701
rect 535 695 539 699
rect 575 697 579 701
rect 595 695 596 699
rect 596 695 599 699
rect 639 697 643 701
rect 703 697 707 701
rect 767 697 771 701
rect 839 697 843 701
rect 911 697 915 701
rect 931 695 932 699
rect 932 695 935 699
rect 1287 696 1291 700
rect 1375 699 1376 703
rect 1376 699 1379 703
rect 1759 699 1760 703
rect 1760 699 1763 703
rect 1975 699 1976 703
rect 1976 699 1979 703
rect 2275 699 2279 703
rect 2463 699 2464 703
rect 2464 699 2467 703
rect 1327 684 1331 688
rect 1367 685 1371 689
rect 1431 685 1435 689
rect 1535 685 1539 689
rect 1639 685 1643 689
rect 111 679 115 683
rect 1655 683 1659 687
rect 1751 685 1755 689
rect 1863 685 1867 689
rect 159 676 163 680
rect 247 676 251 680
rect 327 676 331 680
rect 407 676 411 680
rect 487 676 491 680
rect 559 676 563 680
rect 623 676 627 680
rect 687 676 691 680
rect 751 676 755 680
rect 823 676 827 680
rect 895 676 899 680
rect 1287 679 1291 683
rect 1883 683 1884 687
rect 1884 683 1887 687
rect 1967 685 1971 689
rect 2063 685 2067 689
rect 2151 685 2155 689
rect 2231 685 2235 689
rect 2247 683 2251 687
rect 2311 685 2315 689
rect 2391 685 2395 689
rect 2411 683 2412 687
rect 2412 683 2415 687
rect 2455 685 2459 689
rect 2471 683 2475 687
rect 2503 684 2507 688
rect 111 661 115 665
rect 215 664 219 668
rect 295 664 299 668
rect 375 664 379 668
rect 455 664 459 668
rect 527 664 531 668
rect 591 664 595 668
rect 655 664 659 668
rect 719 664 723 668
rect 783 664 787 668
rect 847 664 851 668
rect 919 664 923 668
rect 1327 667 1331 671
rect 1287 661 1291 665
rect 1351 664 1355 668
rect 1415 664 1419 668
rect 1519 664 1523 668
rect 1623 664 1627 668
rect 1735 664 1739 668
rect 1847 664 1851 668
rect 1951 664 1955 668
rect 2047 664 2051 668
rect 2135 664 2139 668
rect 2215 664 2219 668
rect 2295 664 2299 668
rect 2375 664 2379 668
rect 2439 664 2443 668
rect 2503 667 2507 671
rect 111 644 115 648
rect 231 643 235 647
rect 295 643 299 647
rect 311 643 315 647
rect 319 643 323 647
rect 391 643 395 647
rect 471 643 475 647
rect 495 643 496 647
rect 496 643 499 647
rect 543 643 547 647
rect 607 643 611 647
rect 631 643 632 647
rect 632 643 635 647
rect 671 643 675 647
rect 735 643 739 647
rect 751 643 755 647
rect 799 643 803 647
rect 863 643 867 647
rect 935 643 939 647
rect 943 643 947 647
rect 1287 644 1291 648
rect 1327 641 1331 645
rect 1479 644 1483 648
rect 1559 644 1563 648
rect 1647 644 1651 648
rect 1735 644 1739 648
rect 1831 644 1835 648
rect 1919 644 1923 648
rect 2007 644 2011 648
rect 2087 644 2091 648
rect 2167 644 2171 648
rect 2239 644 2243 648
rect 2311 644 2315 648
rect 2383 644 2387 648
rect 2439 644 2443 648
rect 2503 641 2507 645
rect 223 627 227 631
rect 427 627 431 631
rect 535 627 539 631
rect 751 623 755 627
rect 871 627 872 631
rect 872 627 875 631
rect 1327 624 1331 628
rect 1495 623 1499 627
rect 943 619 947 623
rect 295 603 299 607
rect 415 603 416 607
rect 416 603 419 607
rect 495 603 499 607
rect 1107 611 1111 615
rect 1575 623 1579 627
rect 1663 623 1667 627
rect 1679 623 1683 627
rect 1751 623 1755 627
rect 1759 623 1763 627
rect 1847 623 1851 627
rect 1863 623 1867 627
rect 1935 623 1939 627
rect 2023 623 2027 627
rect 2103 623 2107 627
rect 2175 623 2179 627
rect 2183 623 2187 627
rect 2255 623 2259 627
rect 2275 623 2276 627
rect 2276 623 2279 627
rect 2327 623 2331 627
rect 2343 623 2347 627
rect 2399 623 2403 627
rect 2455 623 2459 627
rect 2463 623 2467 627
rect 2503 624 2507 628
rect 1015 603 1016 607
rect 1016 603 1019 607
rect 1655 603 1659 607
rect 1863 603 1867 607
rect 1903 607 1907 611
rect 2247 607 2251 611
rect 2343 603 2347 607
rect 2407 607 2408 611
rect 2408 607 2411 611
rect 2471 607 2475 611
rect 111 588 115 592
rect 207 589 211 593
rect 215 587 219 591
rect 303 589 307 593
rect 407 589 411 593
rect 427 587 428 591
rect 428 587 431 591
rect 503 589 507 593
rect 599 589 603 593
rect 623 587 624 591
rect 624 587 627 591
rect 687 589 691 593
rect 767 589 771 593
rect 847 589 851 593
rect 871 587 872 591
rect 872 587 875 591
rect 927 589 931 593
rect 1007 589 1011 593
rect 1087 589 1091 593
rect 1107 587 1108 591
rect 1108 587 1111 591
rect 1287 588 1291 592
rect 2299 591 2303 595
rect 1679 583 1680 587
rect 1680 583 1683 587
rect 1835 583 1839 587
rect 2175 583 2179 587
rect 111 571 115 575
rect 191 568 195 572
rect 287 568 291 572
rect 391 568 395 572
rect 487 568 491 572
rect 583 568 587 572
rect 671 568 675 572
rect 751 568 755 572
rect 831 568 835 572
rect 911 568 915 572
rect 991 568 995 572
rect 1071 568 1075 572
rect 1287 571 1291 575
rect 2383 583 2384 587
rect 2384 583 2387 587
rect 2463 583 2464 587
rect 2464 583 2467 587
rect 1327 568 1331 572
rect 1455 569 1459 573
rect 1471 567 1475 571
rect 1559 569 1563 573
rect 1671 569 1675 573
rect 1775 569 1779 573
rect 1879 569 1883 573
rect 1903 567 1904 571
rect 1904 567 1907 571
rect 1983 569 1987 573
rect 2087 569 2091 573
rect 2159 567 2163 571
rect 2183 569 2187 573
rect 2279 569 2283 573
rect 2299 567 2300 571
rect 2300 567 2303 571
rect 2375 569 2379 573
rect 2407 567 2411 571
rect 2455 569 2459 573
rect 2463 567 2467 571
rect 2503 568 2507 572
rect 111 549 115 553
rect 175 552 179 556
rect 271 552 275 556
rect 375 552 379 556
rect 487 552 491 556
rect 591 552 595 556
rect 695 552 699 556
rect 791 552 795 556
rect 879 552 883 556
rect 967 552 971 556
rect 1055 552 1059 556
rect 1151 552 1155 556
rect 1287 549 1291 553
rect 1327 551 1331 555
rect 1439 548 1443 552
rect 1543 548 1547 552
rect 1655 548 1659 552
rect 1759 548 1763 552
rect 1863 548 1867 552
rect 1967 548 1971 552
rect 2071 548 2075 552
rect 2167 548 2171 552
rect 2263 548 2267 552
rect 2359 548 2363 552
rect 2439 548 2443 552
rect 2503 551 2507 555
rect 111 532 115 536
rect 191 531 195 535
rect 239 531 243 535
rect 287 531 291 535
rect 391 531 395 535
rect 415 531 416 535
rect 416 531 419 535
rect 503 531 507 535
rect 607 531 611 535
rect 711 531 715 535
rect 743 531 747 535
rect 807 531 811 535
rect 895 531 899 535
rect 983 531 987 535
rect 1015 531 1019 535
rect 1071 531 1075 535
rect 1167 531 1171 535
rect 1175 531 1179 535
rect 1287 532 1291 536
rect 1327 529 1331 533
rect 1367 532 1371 536
rect 1447 532 1451 536
rect 1527 532 1531 536
rect 1615 532 1619 536
rect 1711 532 1715 536
rect 1799 532 1803 536
rect 1887 532 1891 536
rect 1975 532 1979 536
rect 2063 532 2067 536
rect 2151 532 2155 536
rect 2247 532 2251 536
rect 2343 532 2347 536
rect 2439 532 2443 536
rect 2503 529 2507 533
rect 215 515 219 519
rect 495 511 499 515
rect 623 511 627 515
rect 1079 515 1080 519
rect 1080 515 1083 519
rect 1327 512 1331 516
rect 1383 511 1387 515
rect 1175 507 1179 511
rect 1391 511 1395 515
rect 1463 511 1467 515
rect 1543 511 1547 515
rect 1551 511 1555 515
rect 1631 511 1635 515
rect 1727 511 1731 515
rect 1815 511 1819 515
rect 1835 511 1836 515
rect 1836 511 1839 515
rect 1903 511 1907 515
rect 1991 511 1995 515
rect 1179 499 1183 503
rect 2079 511 2083 515
rect 2151 511 2155 515
rect 2167 511 2171 515
rect 2263 511 2267 515
rect 2271 511 2275 515
rect 2359 511 2363 515
rect 2383 511 2384 515
rect 2384 511 2387 515
rect 2455 511 2459 515
rect 2503 512 2507 516
rect 239 491 243 495
rect 343 491 347 495
rect 743 491 744 495
rect 744 491 747 495
rect 1259 491 1263 495
rect 1471 495 1472 499
rect 1472 495 1475 499
rect 1551 487 1555 491
rect 1719 491 1723 495
rect 2055 491 2059 495
rect 2159 495 2163 499
rect 2479 495 2483 499
rect 111 476 115 480
rect 151 477 155 481
rect 159 475 163 479
rect 247 477 251 481
rect 367 477 371 481
rect 487 477 491 481
rect 495 475 499 479
rect 615 477 619 481
rect 623 475 627 479
rect 735 477 739 481
rect 847 477 851 481
rect 951 477 955 481
rect 1055 477 1059 481
rect 1079 475 1080 479
rect 1080 475 1083 479
rect 1159 477 1163 481
rect 1179 475 1180 479
rect 1180 475 1183 479
rect 1239 477 1243 481
rect 1287 476 1291 480
rect 1391 479 1395 483
rect 2071 479 2075 483
rect 111 459 115 463
rect 135 456 139 460
rect 231 456 235 460
rect 351 456 355 460
rect 471 456 475 460
rect 599 456 603 460
rect 719 456 723 460
rect 831 456 835 460
rect 935 456 939 460
rect 1039 456 1043 460
rect 1143 456 1147 460
rect 1223 456 1227 460
rect 1287 459 1291 463
rect 1551 471 1555 475
rect 2351 479 2355 483
rect 2151 471 2155 475
rect 2463 471 2464 475
rect 2464 471 2467 475
rect 1327 456 1331 460
rect 1367 457 1371 461
rect 1431 457 1435 461
rect 1519 457 1523 461
rect 1527 455 1531 459
rect 1615 457 1619 461
rect 1711 457 1715 461
rect 1719 455 1723 459
rect 1815 457 1819 461
rect 1927 457 1931 461
rect 2023 455 2027 459
rect 2055 457 2059 461
rect 2071 455 2075 459
rect 2191 457 2195 461
rect 2335 457 2339 461
rect 2351 455 2355 459
rect 2455 457 2459 461
rect 2471 455 2475 459
rect 2503 456 2507 460
rect 111 437 115 441
rect 135 440 139 444
rect 191 440 195 444
rect 247 440 251 444
rect 303 440 307 444
rect 383 440 387 444
rect 471 440 475 444
rect 567 440 571 444
rect 671 440 675 444
rect 783 440 787 444
rect 895 440 899 444
rect 1007 440 1011 444
rect 1127 440 1131 444
rect 1223 440 1227 444
rect 1287 437 1291 441
rect 1327 439 1331 443
rect 1351 436 1355 440
rect 1415 436 1419 440
rect 1503 436 1507 440
rect 1599 436 1603 440
rect 1695 436 1699 440
rect 1799 436 1803 440
rect 1911 436 1915 440
rect 2039 436 2043 440
rect 2175 436 2179 440
rect 2319 436 2323 440
rect 2439 436 2443 440
rect 2503 439 2507 443
rect 111 420 115 424
rect 151 419 155 423
rect 207 419 211 423
rect 215 419 219 423
rect 263 419 267 423
rect 319 419 323 423
rect 343 419 344 423
rect 344 419 347 423
rect 399 419 403 423
rect 415 419 419 423
rect 487 419 491 423
rect 583 419 587 423
rect 687 419 691 423
rect 799 419 803 423
rect 911 419 915 423
rect 919 419 923 423
rect 1023 419 1027 423
rect 1143 419 1147 423
rect 1239 419 1243 423
rect 1259 419 1260 423
rect 1260 419 1263 423
rect 1287 420 1291 424
rect 1327 417 1331 421
rect 1351 420 1355 424
rect 1423 420 1427 424
rect 1511 420 1515 424
rect 1599 420 1603 424
rect 1679 420 1683 424
rect 1775 420 1779 424
rect 1887 420 1891 424
rect 2015 420 2019 424
rect 2159 420 2163 424
rect 2311 420 2315 424
rect 2439 420 2443 424
rect 2503 417 2507 421
rect 159 403 160 407
rect 160 403 163 407
rect 415 399 419 403
rect 531 403 535 407
rect 623 403 627 407
rect 991 403 995 407
rect 1327 400 1331 404
rect 1367 399 1371 403
rect 1375 399 1379 403
rect 1439 399 1443 403
rect 1527 399 1531 403
rect 1551 399 1552 403
rect 1552 399 1555 403
rect 1615 399 1619 403
rect 1695 399 1699 403
rect 1791 399 1795 403
rect 1815 399 1816 403
rect 1816 399 1819 403
rect 1903 399 1907 403
rect 2031 399 2035 403
rect 299 383 303 387
rect 479 383 483 387
rect 843 383 847 387
rect 1519 383 1523 387
rect 215 375 216 379
rect 216 375 219 379
rect 919 375 923 379
rect 1071 375 1075 379
rect 1375 375 1379 379
rect 2175 399 2179 403
rect 2327 399 2331 403
rect 2335 399 2339 403
rect 2455 399 2459 403
rect 2463 399 2467 403
rect 2503 400 2507 404
rect 1755 375 1759 379
rect 2023 383 2027 387
rect 2471 383 2475 387
rect 2335 375 2339 379
rect 111 360 115 364
rect 151 361 155 365
rect 159 359 163 363
rect 207 361 211 365
rect 279 361 283 365
rect 299 359 300 363
rect 300 359 303 363
rect 359 361 363 365
rect 431 361 435 365
rect 511 361 515 365
rect 531 359 532 363
rect 532 359 535 363
rect 591 361 595 365
rect 639 359 643 363
rect 671 361 675 365
rect 751 361 755 365
rect 823 361 827 365
rect 843 359 844 363
rect 844 359 847 363
rect 895 361 899 365
rect 967 361 971 365
rect 991 359 992 363
rect 992 359 995 363
rect 1039 361 1043 365
rect 1111 361 1115 365
rect 1183 361 1187 365
rect 1231 359 1235 363
rect 1239 361 1243 365
rect 1287 360 1291 364
rect 1671 359 1675 363
rect 1815 359 1816 363
rect 1816 359 1819 363
rect 2463 359 2464 363
rect 2464 359 2467 363
rect 111 343 115 347
rect 135 340 139 344
rect 191 340 195 344
rect 263 340 267 344
rect 343 340 347 344
rect 415 340 419 344
rect 495 340 499 344
rect 575 340 579 344
rect 655 340 659 344
rect 735 340 739 344
rect 807 340 811 344
rect 879 340 883 344
rect 951 340 955 344
rect 1023 340 1027 344
rect 1095 340 1099 344
rect 1167 340 1171 344
rect 1223 340 1227 344
rect 1287 343 1291 347
rect 1327 344 1331 348
rect 1679 345 1683 349
rect 1735 345 1739 349
rect 1755 343 1756 347
rect 1756 343 1759 347
rect 1807 345 1811 349
rect 1903 345 1907 349
rect 2023 345 2027 349
rect 2159 345 2163 349
rect 2303 345 2307 349
rect 2319 343 2323 347
rect 2455 345 2459 349
rect 2479 343 2480 347
rect 2480 343 2483 347
rect 2503 344 2507 348
rect 1327 327 1331 331
rect 111 317 115 321
rect 135 320 139 324
rect 199 320 203 324
rect 287 320 291 324
rect 375 320 379 324
rect 455 320 459 324
rect 543 320 547 324
rect 631 320 635 324
rect 727 320 731 324
rect 823 320 827 324
rect 927 320 931 324
rect 1031 320 1035 324
rect 1135 320 1139 324
rect 1223 320 1227 324
rect 1663 324 1667 328
rect 1719 324 1723 328
rect 1791 324 1795 328
rect 1887 324 1891 328
rect 2007 324 2011 328
rect 2143 324 2147 328
rect 2287 324 2291 328
rect 2439 324 2443 328
rect 2503 327 2507 331
rect 1287 317 1291 321
rect 1327 309 1331 313
rect 1351 312 1355 316
rect 1431 312 1435 316
rect 1527 312 1531 316
rect 1623 312 1627 316
rect 1711 312 1715 316
rect 1807 312 1811 316
rect 1911 312 1915 316
rect 2023 312 2027 316
rect 2151 312 2155 316
rect 2287 312 2291 316
rect 2423 312 2427 316
rect 2503 309 2507 313
rect 111 300 115 304
rect 151 299 155 303
rect 215 299 219 303
rect 303 299 307 303
rect 335 299 339 303
rect 391 299 395 303
rect 471 299 475 303
rect 479 299 483 303
rect 559 299 563 303
rect 647 299 651 303
rect 159 283 160 287
rect 160 283 163 287
rect 743 299 747 303
rect 839 299 843 303
rect 943 299 947 303
rect 951 299 955 303
rect 1047 299 1051 303
rect 1071 299 1072 303
rect 1072 299 1075 303
rect 1151 299 1155 303
rect 1239 299 1243 303
rect 1279 299 1283 303
rect 1287 300 1291 304
rect 1327 292 1331 296
rect 1367 291 1371 295
rect 1447 291 1451 295
rect 543 283 547 287
rect 639 283 643 287
rect 1223 283 1227 287
rect 1231 283 1235 287
rect 1543 291 1547 295
rect 1551 291 1555 295
rect 1639 291 1643 295
rect 1671 291 1675 295
rect 1727 291 1731 295
rect 1823 291 1827 295
rect 1927 291 1931 295
rect 2039 291 2043 295
rect 2167 291 2171 295
rect 2303 291 2307 295
rect 2311 291 2315 295
rect 2439 291 2443 295
rect 2463 291 2464 295
rect 2464 291 2467 295
rect 2503 292 2507 296
rect 1279 275 1283 279
rect 1807 275 1811 279
rect 2319 271 2323 275
rect 2415 275 2419 279
rect 347 263 351 267
rect 635 263 639 267
rect 923 263 927 267
rect 335 255 336 259
rect 336 255 339 259
rect 643 255 647 259
rect 951 255 955 259
rect 999 255 1003 259
rect 1551 259 1555 263
rect 1739 259 1743 263
rect 2311 259 2315 263
rect 111 240 115 244
rect 151 241 155 245
rect 231 241 235 245
rect 263 239 267 243
rect 327 241 331 245
rect 347 239 348 243
rect 348 239 351 243
rect 423 241 427 245
rect 519 241 523 245
rect 543 239 544 243
rect 544 239 547 243
rect 615 241 619 245
rect 635 239 636 243
rect 636 239 639 243
rect 711 241 715 245
rect 807 241 811 245
rect 879 239 883 243
rect 903 241 907 245
rect 923 239 924 243
rect 924 239 927 243
rect 1007 241 1011 245
rect 1111 241 1115 245
rect 1215 241 1219 245
rect 1223 239 1227 243
rect 1287 240 1291 244
rect 1807 243 1811 247
rect 2463 251 2464 255
rect 2464 251 2467 255
rect 1327 236 1331 240
rect 1367 237 1371 241
rect 1439 237 1443 241
rect 1535 237 1539 241
rect 1607 235 1611 239
rect 1631 237 1635 241
rect 1727 237 1731 241
rect 1815 237 1819 241
rect 1903 237 1907 241
rect 1999 237 2003 241
rect 2103 237 2107 241
rect 2215 237 2219 241
rect 2335 237 2339 241
rect 2343 235 2347 239
rect 2455 237 2459 241
rect 2471 235 2475 239
rect 2503 236 2507 240
rect 111 223 115 227
rect 135 220 139 224
rect 215 220 219 224
rect 311 220 315 224
rect 407 220 411 224
rect 503 220 507 224
rect 599 220 603 224
rect 695 220 699 224
rect 791 220 795 224
rect 887 220 891 224
rect 991 220 995 224
rect 1095 220 1099 224
rect 1199 220 1203 224
rect 1287 223 1291 227
rect 1327 219 1331 223
rect 1351 216 1355 220
rect 1423 216 1427 220
rect 1519 216 1523 220
rect 1615 216 1619 220
rect 1711 216 1715 220
rect 1799 216 1803 220
rect 1887 216 1891 220
rect 1983 216 1987 220
rect 2087 216 2091 220
rect 2199 216 2203 220
rect 2319 216 2323 220
rect 2439 216 2443 220
rect 2503 219 2507 223
rect 111 197 115 201
rect 159 200 163 204
rect 239 200 243 204
rect 327 200 331 204
rect 415 200 419 204
rect 511 200 515 204
rect 607 200 611 204
rect 695 200 699 204
rect 783 200 787 204
rect 871 200 875 204
rect 959 200 963 204
rect 1047 200 1051 204
rect 1135 200 1139 204
rect 1287 197 1291 201
rect 1327 197 1331 201
rect 1391 200 1395 204
rect 1495 200 1499 204
rect 1599 200 1603 204
rect 1711 200 1715 204
rect 1815 200 1819 204
rect 1919 200 1923 204
rect 2015 200 2019 204
rect 2111 200 2115 204
rect 2199 200 2203 204
rect 2287 200 2291 204
rect 2375 200 2379 204
rect 2439 200 2443 204
rect 2503 197 2507 201
rect 111 180 115 184
rect 175 179 179 183
rect 183 179 187 183
rect 255 179 259 183
rect 343 179 347 183
rect 351 179 355 183
rect 431 179 435 183
rect 527 179 531 183
rect 623 179 627 183
rect 643 179 644 183
rect 644 179 647 183
rect 711 179 715 183
rect 719 179 723 183
rect 799 179 803 183
rect 815 179 819 183
rect 887 179 891 183
rect 975 179 979 183
rect 999 179 1000 183
rect 1000 179 1003 183
rect 1063 179 1067 183
rect 1151 179 1155 183
rect 1287 180 1291 184
rect 1327 180 1331 184
rect 1407 179 1411 183
rect 1415 179 1419 183
rect 1511 179 1515 183
rect 1527 179 1531 183
rect 1615 179 1619 183
rect 1727 179 1731 183
rect 1739 179 1743 183
rect 1831 179 1835 183
rect 1935 179 1939 183
rect 2031 179 2035 183
rect 2127 179 2131 183
rect 2215 179 2219 183
rect 2231 179 2235 183
rect 2303 179 2307 183
rect 2391 179 2395 183
rect 2415 179 2416 183
rect 2416 179 2419 183
rect 2455 179 2459 183
rect 2463 179 2467 183
rect 2503 180 2507 184
rect 263 163 264 167
rect 264 163 267 167
rect 351 155 355 159
rect 643 159 647 163
rect 815 159 819 163
rect 879 163 883 167
rect 1219 163 1223 167
rect 1527 159 1531 163
rect 1607 163 1611 167
rect 1839 163 1840 167
rect 1840 163 1843 167
rect 2355 163 2359 167
rect 2471 163 2475 167
rect 2343 155 2347 159
rect 183 131 187 135
rect 719 131 723 135
rect 1415 131 1419 135
rect 2231 131 2235 135
rect 2463 123 2464 127
rect 2464 123 2467 127
rect 111 108 115 112
rect 151 109 155 113
rect 207 109 211 113
rect 263 109 267 113
rect 319 109 323 113
rect 375 109 379 113
rect 431 109 435 113
rect 487 109 491 113
rect 551 109 555 113
rect 623 109 627 113
rect 643 107 644 111
rect 644 107 647 111
rect 687 109 691 113
rect 751 109 755 113
rect 815 109 819 113
rect 879 109 883 113
rect 943 109 947 113
rect 1007 109 1011 113
rect 1071 109 1075 113
rect 1135 109 1139 113
rect 1199 109 1203 113
rect 1219 107 1220 111
rect 1220 107 1223 111
rect 1287 108 1291 112
rect 1327 108 1331 112
rect 1367 109 1371 113
rect 1423 109 1427 113
rect 1479 109 1483 113
rect 1535 109 1539 113
rect 1591 109 1595 113
rect 1647 109 1651 113
rect 1703 109 1707 113
rect 1759 109 1763 113
rect 1815 109 1819 113
rect 1839 107 1840 111
rect 1840 107 1843 111
rect 1871 109 1875 113
rect 1927 109 1931 113
rect 1983 109 1987 113
rect 2039 109 2043 113
rect 2095 109 2099 113
rect 2159 109 2163 113
rect 2223 109 2227 113
rect 2287 109 2291 113
rect 2343 109 2347 113
rect 2355 107 2359 111
rect 2399 109 2403 113
rect 2455 109 2459 113
rect 2503 108 2507 112
rect 111 91 115 95
rect 135 88 139 92
rect 191 88 195 92
rect 247 88 251 92
rect 303 88 307 92
rect 359 88 363 92
rect 415 88 419 92
rect 471 88 475 92
rect 535 88 539 92
rect 607 88 611 92
rect 671 88 675 92
rect 735 88 739 92
rect 799 88 803 92
rect 863 88 867 92
rect 927 88 931 92
rect 991 88 995 92
rect 1055 88 1059 92
rect 1119 88 1123 92
rect 1183 88 1187 92
rect 1287 91 1291 95
rect 1327 91 1331 95
rect 1351 88 1355 92
rect 1407 88 1411 92
rect 1463 88 1467 92
rect 1519 88 1523 92
rect 1575 88 1579 92
rect 1631 88 1635 92
rect 1687 88 1691 92
rect 1743 88 1747 92
rect 1799 88 1803 92
rect 1855 88 1859 92
rect 1911 88 1915 92
rect 1967 88 1971 92
rect 2023 88 2027 92
rect 2079 88 2083 92
rect 2143 88 2147 92
rect 2207 88 2211 92
rect 2271 88 2275 92
rect 2327 88 2331 92
rect 2383 88 2387 92
rect 2439 88 2443 92
rect 2503 91 2507 95
<< m3 >>
rect 111 2582 115 2583
rect 111 2577 115 2578
rect 719 2582 723 2583
rect 719 2577 723 2578
rect 775 2582 779 2583
rect 775 2577 779 2578
rect 831 2582 835 2583
rect 831 2577 835 2578
rect 887 2582 891 2583
rect 887 2577 891 2578
rect 943 2582 947 2583
rect 943 2577 947 2578
rect 1287 2582 1291 2583
rect 1287 2577 1291 2578
rect 112 2557 114 2577
rect 720 2558 722 2577
rect 776 2558 778 2577
rect 832 2558 834 2577
rect 888 2558 890 2577
rect 944 2558 946 2577
rect 718 2557 724 2558
rect 110 2556 116 2557
rect 110 2552 111 2556
rect 115 2552 116 2556
rect 718 2553 719 2557
rect 723 2553 724 2557
rect 718 2552 724 2553
rect 774 2557 780 2558
rect 774 2553 775 2557
rect 779 2553 780 2557
rect 774 2552 780 2553
rect 830 2557 836 2558
rect 830 2553 831 2557
rect 835 2553 836 2557
rect 830 2552 836 2553
rect 886 2557 892 2558
rect 886 2553 887 2557
rect 891 2553 892 2557
rect 886 2552 892 2553
rect 942 2557 948 2558
rect 1288 2557 1290 2577
rect 1327 2558 1331 2559
rect 942 2553 943 2557
rect 947 2553 948 2557
rect 1286 2556 1292 2557
rect 942 2552 948 2553
rect 950 2555 956 2556
rect 110 2551 116 2552
rect 950 2551 951 2555
rect 955 2551 956 2555
rect 1286 2552 1287 2556
rect 1291 2552 1292 2556
rect 1327 2553 1331 2554
rect 1399 2558 1403 2559
rect 1399 2553 1403 2554
rect 1455 2558 1459 2559
rect 1455 2553 1459 2554
rect 1511 2558 1515 2559
rect 1511 2553 1515 2554
rect 1567 2558 1571 2559
rect 1567 2553 1571 2554
rect 1623 2558 1627 2559
rect 1623 2553 1627 2554
rect 1679 2558 1683 2559
rect 1735 2558 1739 2559
rect 1679 2553 1683 2554
rect 1710 2555 1716 2556
rect 1286 2551 1292 2552
rect 950 2550 956 2551
rect 110 2539 116 2540
rect 110 2535 111 2539
rect 115 2535 116 2539
rect 110 2534 116 2535
rect 702 2536 708 2537
rect 112 2531 114 2534
rect 702 2532 703 2536
rect 707 2532 708 2536
rect 702 2531 708 2532
rect 758 2536 764 2537
rect 758 2532 759 2536
rect 763 2532 764 2536
rect 758 2531 764 2532
rect 814 2536 820 2537
rect 814 2532 815 2536
rect 819 2532 820 2536
rect 814 2531 820 2532
rect 870 2536 876 2537
rect 870 2532 871 2536
rect 875 2532 876 2536
rect 870 2531 876 2532
rect 926 2536 932 2537
rect 926 2532 927 2536
rect 931 2532 932 2536
rect 926 2531 932 2532
rect 111 2530 115 2531
rect 111 2525 115 2526
rect 167 2530 171 2531
rect 167 2525 171 2526
rect 223 2530 227 2531
rect 223 2525 227 2526
rect 279 2530 283 2531
rect 279 2525 283 2526
rect 343 2530 347 2531
rect 343 2525 347 2526
rect 407 2530 411 2531
rect 407 2525 411 2526
rect 479 2530 483 2531
rect 479 2525 483 2526
rect 559 2530 563 2531
rect 559 2525 563 2526
rect 639 2530 643 2531
rect 639 2525 643 2526
rect 703 2530 707 2531
rect 703 2525 707 2526
rect 719 2530 723 2531
rect 719 2525 723 2526
rect 759 2530 763 2531
rect 759 2525 763 2526
rect 799 2530 803 2531
rect 799 2525 803 2526
rect 815 2530 819 2531
rect 815 2525 819 2526
rect 871 2530 875 2531
rect 871 2525 875 2526
rect 879 2530 883 2531
rect 879 2525 883 2526
rect 927 2530 931 2531
rect 927 2525 931 2526
rect 112 2522 114 2525
rect 166 2524 172 2525
rect 110 2521 116 2522
rect 110 2517 111 2521
rect 115 2517 116 2521
rect 166 2520 167 2524
rect 171 2520 172 2524
rect 166 2519 172 2520
rect 222 2524 228 2525
rect 222 2520 223 2524
rect 227 2520 228 2524
rect 222 2519 228 2520
rect 278 2524 284 2525
rect 278 2520 279 2524
rect 283 2520 284 2524
rect 278 2519 284 2520
rect 342 2524 348 2525
rect 342 2520 343 2524
rect 347 2520 348 2524
rect 342 2519 348 2520
rect 406 2524 412 2525
rect 406 2520 407 2524
rect 411 2520 412 2524
rect 406 2519 412 2520
rect 478 2524 484 2525
rect 478 2520 479 2524
rect 483 2520 484 2524
rect 478 2519 484 2520
rect 558 2524 564 2525
rect 558 2520 559 2524
rect 563 2520 564 2524
rect 558 2519 564 2520
rect 638 2524 644 2525
rect 638 2520 639 2524
rect 643 2520 644 2524
rect 638 2519 644 2520
rect 718 2524 724 2525
rect 718 2520 719 2524
rect 723 2520 724 2524
rect 718 2519 724 2520
rect 798 2524 804 2525
rect 798 2520 799 2524
rect 803 2520 804 2524
rect 798 2519 804 2520
rect 878 2524 884 2525
rect 878 2520 879 2524
rect 883 2520 884 2524
rect 878 2519 884 2520
rect 110 2516 116 2517
rect 110 2504 116 2505
rect 110 2500 111 2504
rect 115 2500 116 2504
rect 110 2499 116 2500
rect 182 2503 188 2504
rect 182 2499 183 2503
rect 187 2499 188 2503
rect 112 2479 114 2499
rect 182 2498 188 2499
rect 238 2503 244 2504
rect 238 2499 239 2503
rect 243 2499 244 2503
rect 238 2498 244 2499
rect 254 2503 260 2504
rect 254 2499 255 2503
rect 259 2499 260 2503
rect 254 2498 260 2499
rect 294 2503 300 2504
rect 294 2499 295 2503
rect 299 2499 300 2503
rect 294 2498 300 2499
rect 358 2503 364 2504
rect 358 2499 359 2503
rect 363 2499 364 2503
rect 358 2498 364 2499
rect 422 2503 428 2504
rect 422 2499 423 2503
rect 427 2499 428 2503
rect 422 2498 428 2499
rect 494 2503 500 2504
rect 494 2499 495 2503
rect 499 2499 500 2503
rect 494 2498 500 2499
rect 574 2503 580 2504
rect 574 2499 575 2503
rect 579 2499 580 2503
rect 574 2498 580 2499
rect 590 2503 596 2504
rect 590 2499 591 2503
rect 595 2499 596 2503
rect 590 2498 596 2499
rect 654 2503 660 2504
rect 654 2499 655 2503
rect 659 2499 660 2503
rect 654 2498 660 2499
rect 734 2503 740 2504
rect 734 2499 735 2503
rect 739 2499 740 2503
rect 734 2498 740 2499
rect 814 2503 820 2504
rect 814 2499 815 2503
rect 819 2499 820 2503
rect 814 2498 820 2499
rect 894 2503 900 2504
rect 894 2499 895 2503
rect 899 2499 900 2503
rect 894 2498 900 2499
rect 184 2479 186 2498
rect 240 2479 242 2498
rect 111 2478 115 2479
rect 111 2473 115 2474
rect 183 2478 187 2479
rect 183 2473 187 2474
rect 239 2478 243 2479
rect 239 2473 243 2474
rect 247 2478 251 2479
rect 247 2473 251 2474
rect 112 2453 114 2473
rect 184 2454 186 2473
rect 248 2454 250 2473
rect 256 2468 258 2498
rect 296 2479 298 2498
rect 360 2479 362 2498
rect 424 2479 426 2498
rect 496 2479 498 2498
rect 576 2479 578 2498
rect 592 2484 594 2498
rect 622 2487 628 2488
rect 590 2483 596 2484
rect 590 2479 591 2483
rect 595 2479 596 2483
rect 622 2483 623 2487
rect 627 2483 628 2487
rect 622 2482 628 2483
rect 295 2478 299 2479
rect 295 2473 299 2474
rect 327 2478 331 2479
rect 327 2473 331 2474
rect 359 2478 363 2479
rect 359 2473 363 2474
rect 415 2478 419 2479
rect 415 2473 419 2474
rect 423 2478 427 2479
rect 495 2478 499 2479
rect 423 2473 427 2474
rect 434 2475 440 2476
rect 254 2467 260 2468
rect 254 2463 255 2467
rect 259 2463 260 2467
rect 254 2462 260 2463
rect 328 2454 330 2473
rect 416 2454 418 2473
rect 434 2471 435 2475
rect 439 2471 440 2475
rect 495 2473 499 2474
rect 503 2478 507 2479
rect 503 2473 507 2474
rect 575 2478 579 2479
rect 590 2478 596 2479
rect 599 2478 603 2479
rect 575 2473 579 2474
rect 599 2473 603 2474
rect 434 2470 440 2471
rect 182 2453 188 2454
rect 110 2452 116 2453
rect 110 2448 111 2452
rect 115 2448 116 2452
rect 182 2449 183 2453
rect 187 2449 188 2453
rect 246 2453 252 2454
rect 182 2448 188 2449
rect 190 2451 196 2452
rect 110 2447 116 2448
rect 190 2447 191 2451
rect 195 2447 196 2451
rect 246 2449 247 2453
rect 251 2449 252 2453
rect 246 2448 252 2449
rect 326 2453 332 2454
rect 326 2449 327 2453
rect 331 2449 332 2453
rect 326 2448 332 2449
rect 414 2453 420 2454
rect 414 2449 415 2453
rect 419 2449 420 2453
rect 436 2452 438 2470
rect 504 2454 506 2473
rect 600 2454 602 2473
rect 502 2453 508 2454
rect 414 2448 420 2449
rect 434 2451 440 2452
rect 190 2446 196 2447
rect 434 2447 435 2451
rect 439 2447 440 2451
rect 502 2449 503 2453
rect 507 2449 508 2453
rect 502 2448 508 2449
rect 598 2453 604 2454
rect 598 2449 599 2453
rect 603 2449 604 2453
rect 624 2452 626 2482
rect 656 2479 658 2498
rect 736 2479 738 2498
rect 816 2479 818 2498
rect 896 2479 898 2498
rect 952 2484 954 2550
rect 1286 2539 1292 2540
rect 1286 2535 1287 2539
rect 1291 2535 1292 2539
rect 1286 2534 1292 2535
rect 1288 2531 1290 2534
rect 1328 2533 1330 2553
rect 1400 2534 1402 2553
rect 1456 2534 1458 2553
rect 1512 2534 1514 2553
rect 1568 2534 1570 2553
rect 1624 2534 1626 2553
rect 1680 2534 1682 2553
rect 1710 2551 1711 2555
rect 1715 2551 1716 2555
rect 1735 2553 1739 2554
rect 1791 2558 1795 2559
rect 1791 2553 1795 2554
rect 1847 2558 1851 2559
rect 1847 2553 1851 2554
rect 1903 2558 1907 2559
rect 1903 2553 1907 2554
rect 1959 2558 1963 2559
rect 1959 2553 1963 2554
rect 2015 2558 2019 2559
rect 2015 2553 2019 2554
rect 2071 2558 2075 2559
rect 2071 2553 2075 2554
rect 2127 2558 2131 2559
rect 2127 2553 2131 2554
rect 2183 2558 2187 2559
rect 2183 2553 2187 2554
rect 2503 2558 2507 2559
rect 2503 2553 2507 2554
rect 1710 2550 1716 2551
rect 1398 2533 1404 2534
rect 1326 2532 1332 2533
rect 959 2530 963 2531
rect 959 2525 963 2526
rect 1039 2530 1043 2531
rect 1039 2525 1043 2526
rect 1287 2530 1291 2531
rect 1326 2528 1327 2532
rect 1331 2528 1332 2532
rect 1398 2529 1399 2533
rect 1403 2529 1404 2533
rect 1398 2528 1404 2529
rect 1454 2533 1460 2534
rect 1454 2529 1455 2533
rect 1459 2529 1460 2533
rect 1454 2528 1460 2529
rect 1510 2533 1516 2534
rect 1510 2529 1511 2533
rect 1515 2529 1516 2533
rect 1510 2528 1516 2529
rect 1566 2533 1572 2534
rect 1566 2529 1567 2533
rect 1571 2529 1572 2533
rect 1566 2528 1572 2529
rect 1622 2533 1628 2534
rect 1622 2529 1623 2533
rect 1627 2529 1628 2533
rect 1622 2528 1628 2529
rect 1678 2533 1684 2534
rect 1678 2529 1679 2533
rect 1683 2529 1684 2533
rect 1678 2528 1684 2529
rect 1326 2527 1332 2528
rect 1287 2525 1291 2526
rect 958 2524 964 2525
rect 958 2520 959 2524
rect 963 2520 964 2524
rect 958 2519 964 2520
rect 1038 2524 1044 2525
rect 1038 2520 1039 2524
rect 1043 2520 1044 2524
rect 1288 2522 1290 2525
rect 1038 2519 1044 2520
rect 1286 2521 1292 2522
rect 1286 2517 1287 2521
rect 1291 2517 1292 2521
rect 1286 2516 1292 2517
rect 1326 2515 1332 2516
rect 1326 2511 1327 2515
rect 1331 2511 1332 2515
rect 1326 2510 1332 2511
rect 1382 2512 1388 2513
rect 1286 2504 1292 2505
rect 974 2503 980 2504
rect 974 2499 975 2503
rect 979 2499 980 2503
rect 974 2498 980 2499
rect 1054 2503 1060 2504
rect 1054 2499 1055 2503
rect 1059 2499 1060 2503
rect 1054 2498 1060 2499
rect 1070 2503 1076 2504
rect 1070 2499 1071 2503
rect 1075 2499 1076 2503
rect 1286 2500 1287 2504
rect 1291 2500 1292 2504
rect 1286 2499 1292 2500
rect 1328 2499 1330 2510
rect 1382 2508 1383 2512
rect 1387 2508 1388 2512
rect 1382 2507 1388 2508
rect 1438 2512 1444 2513
rect 1438 2508 1439 2512
rect 1443 2508 1444 2512
rect 1438 2507 1444 2508
rect 1494 2512 1500 2513
rect 1494 2508 1495 2512
rect 1499 2508 1500 2512
rect 1494 2507 1500 2508
rect 1550 2512 1556 2513
rect 1550 2508 1551 2512
rect 1555 2508 1556 2512
rect 1550 2507 1556 2508
rect 1606 2512 1612 2513
rect 1606 2508 1607 2512
rect 1611 2508 1612 2512
rect 1606 2507 1612 2508
rect 1662 2512 1668 2513
rect 1662 2508 1663 2512
rect 1667 2508 1668 2512
rect 1662 2507 1668 2508
rect 1384 2499 1386 2507
rect 1440 2499 1442 2507
rect 1496 2499 1498 2507
rect 1552 2499 1554 2507
rect 1608 2499 1610 2507
rect 1664 2499 1666 2507
rect 1070 2498 1076 2499
rect 950 2483 956 2484
rect 950 2479 951 2483
rect 955 2479 956 2483
rect 976 2479 978 2498
rect 1056 2479 1058 2498
rect 655 2478 659 2479
rect 655 2473 659 2474
rect 695 2478 699 2479
rect 735 2478 739 2479
rect 695 2473 699 2474
rect 714 2475 720 2476
rect 696 2454 698 2473
rect 714 2471 715 2475
rect 719 2471 720 2475
rect 735 2473 739 2474
rect 791 2478 795 2479
rect 791 2473 795 2474
rect 815 2478 819 2479
rect 815 2473 819 2474
rect 879 2478 883 2479
rect 879 2473 883 2474
rect 895 2478 899 2479
rect 950 2478 956 2479
rect 967 2478 971 2479
rect 895 2473 899 2474
rect 967 2473 971 2474
rect 975 2478 979 2479
rect 975 2473 979 2474
rect 1055 2478 1059 2479
rect 1055 2473 1059 2474
rect 1063 2478 1067 2479
rect 1072 2476 1074 2498
rect 1288 2479 1290 2499
rect 1327 2498 1331 2499
rect 1327 2493 1331 2494
rect 1351 2498 1355 2499
rect 1351 2493 1355 2494
rect 1383 2498 1387 2499
rect 1383 2493 1387 2494
rect 1423 2498 1427 2499
rect 1423 2493 1427 2494
rect 1439 2498 1443 2499
rect 1439 2493 1443 2494
rect 1495 2498 1499 2499
rect 1495 2493 1499 2494
rect 1511 2498 1515 2499
rect 1511 2493 1515 2494
rect 1551 2498 1555 2499
rect 1551 2493 1555 2494
rect 1599 2498 1603 2499
rect 1599 2493 1603 2494
rect 1607 2498 1611 2499
rect 1607 2493 1611 2494
rect 1663 2498 1667 2499
rect 1663 2493 1667 2494
rect 1687 2498 1691 2499
rect 1687 2493 1691 2494
rect 1328 2490 1330 2493
rect 1350 2492 1356 2493
rect 1326 2489 1332 2490
rect 1326 2485 1327 2489
rect 1331 2485 1332 2489
rect 1350 2488 1351 2492
rect 1355 2488 1356 2492
rect 1350 2487 1356 2488
rect 1422 2492 1428 2493
rect 1422 2488 1423 2492
rect 1427 2488 1428 2492
rect 1422 2487 1428 2488
rect 1510 2492 1516 2493
rect 1510 2488 1511 2492
rect 1515 2488 1516 2492
rect 1510 2487 1516 2488
rect 1598 2492 1604 2493
rect 1598 2488 1599 2492
rect 1603 2488 1604 2492
rect 1598 2487 1604 2488
rect 1686 2492 1692 2493
rect 1686 2488 1687 2492
rect 1691 2488 1692 2492
rect 1686 2487 1692 2488
rect 1326 2484 1332 2485
rect 1159 2478 1163 2479
rect 1063 2473 1067 2474
rect 1070 2475 1076 2476
rect 714 2470 720 2471
rect 694 2453 700 2454
rect 598 2448 604 2449
rect 622 2451 628 2452
rect 434 2446 440 2447
rect 622 2447 623 2451
rect 627 2447 628 2451
rect 694 2449 695 2453
rect 699 2449 700 2453
rect 716 2452 718 2470
rect 762 2467 768 2468
rect 762 2463 763 2467
rect 767 2463 768 2467
rect 762 2462 768 2463
rect 694 2448 700 2449
rect 714 2451 720 2452
rect 622 2446 628 2447
rect 714 2447 715 2451
rect 719 2447 720 2451
rect 714 2446 720 2447
rect 110 2435 116 2436
rect 110 2431 111 2435
rect 115 2431 116 2435
rect 110 2430 116 2431
rect 166 2432 172 2433
rect 112 2423 114 2430
rect 166 2428 167 2432
rect 171 2428 172 2432
rect 166 2427 172 2428
rect 168 2423 170 2427
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 151 2422 155 2423
rect 151 2417 155 2418
rect 167 2422 171 2423
rect 167 2417 171 2418
rect 112 2414 114 2417
rect 150 2416 156 2417
rect 110 2413 116 2414
rect 110 2409 111 2413
rect 115 2409 116 2413
rect 150 2412 151 2416
rect 155 2412 156 2416
rect 150 2411 156 2412
rect 110 2408 116 2409
rect 110 2396 116 2397
rect 110 2392 111 2396
rect 115 2392 116 2396
rect 110 2391 116 2392
rect 166 2395 172 2396
rect 166 2391 167 2395
rect 171 2391 172 2395
rect 112 2371 114 2391
rect 166 2390 172 2391
rect 168 2371 170 2390
rect 192 2380 194 2446
rect 230 2432 236 2433
rect 230 2428 231 2432
rect 235 2428 236 2432
rect 230 2427 236 2428
rect 310 2432 316 2433
rect 310 2428 311 2432
rect 315 2428 316 2432
rect 310 2427 316 2428
rect 398 2432 404 2433
rect 398 2428 399 2432
rect 403 2428 404 2432
rect 398 2427 404 2428
rect 486 2432 492 2433
rect 486 2428 487 2432
rect 491 2428 492 2432
rect 486 2427 492 2428
rect 582 2432 588 2433
rect 582 2428 583 2432
rect 587 2428 588 2432
rect 582 2427 588 2428
rect 678 2432 684 2433
rect 678 2428 679 2432
rect 683 2428 684 2432
rect 678 2427 684 2428
rect 232 2423 234 2427
rect 312 2423 314 2427
rect 400 2423 402 2427
rect 488 2423 490 2427
rect 584 2423 586 2427
rect 680 2423 682 2427
rect 231 2422 235 2423
rect 231 2417 235 2418
rect 311 2422 315 2423
rect 311 2417 315 2418
rect 319 2422 323 2423
rect 319 2417 323 2418
rect 399 2422 403 2423
rect 399 2417 403 2418
rect 415 2422 419 2423
rect 415 2417 419 2418
rect 487 2422 491 2423
rect 487 2417 491 2418
rect 519 2422 523 2423
rect 519 2417 523 2418
rect 583 2422 587 2423
rect 583 2417 587 2418
rect 623 2422 627 2423
rect 623 2417 627 2418
rect 679 2422 683 2423
rect 679 2417 683 2418
rect 727 2422 731 2423
rect 727 2417 731 2418
rect 230 2416 236 2417
rect 230 2412 231 2416
rect 235 2412 236 2416
rect 230 2411 236 2412
rect 318 2416 324 2417
rect 318 2412 319 2416
rect 323 2412 324 2416
rect 318 2411 324 2412
rect 414 2416 420 2417
rect 414 2412 415 2416
rect 419 2412 420 2416
rect 414 2411 420 2412
rect 518 2416 524 2417
rect 518 2412 519 2416
rect 523 2412 524 2416
rect 518 2411 524 2412
rect 622 2416 628 2417
rect 622 2412 623 2416
rect 627 2412 628 2416
rect 622 2411 628 2412
rect 726 2416 732 2417
rect 726 2412 727 2416
rect 731 2412 732 2416
rect 726 2411 732 2412
rect 764 2396 766 2462
rect 792 2454 794 2473
rect 880 2454 882 2473
rect 968 2454 970 2473
rect 1064 2454 1066 2473
rect 1070 2471 1071 2475
rect 1075 2471 1076 2475
rect 1159 2473 1163 2474
rect 1287 2478 1291 2479
rect 1287 2473 1291 2474
rect 1070 2470 1076 2471
rect 1160 2454 1162 2473
rect 790 2453 796 2454
rect 790 2449 791 2453
rect 795 2449 796 2453
rect 790 2448 796 2449
rect 878 2453 884 2454
rect 878 2449 879 2453
rect 883 2449 884 2453
rect 878 2448 884 2449
rect 966 2453 972 2454
rect 966 2449 967 2453
rect 971 2449 972 2453
rect 966 2448 972 2449
rect 1062 2453 1068 2454
rect 1062 2449 1063 2453
rect 1067 2449 1068 2453
rect 1062 2448 1068 2449
rect 1158 2453 1164 2454
rect 1288 2453 1290 2473
rect 1326 2472 1332 2473
rect 1712 2472 1714 2550
rect 1736 2534 1738 2553
rect 1792 2534 1794 2553
rect 1848 2534 1850 2553
rect 1904 2534 1906 2553
rect 1960 2534 1962 2553
rect 2016 2534 2018 2553
rect 2072 2534 2074 2553
rect 2128 2534 2130 2553
rect 2184 2534 2186 2553
rect 1734 2533 1740 2534
rect 1734 2529 1735 2533
rect 1739 2529 1740 2533
rect 1734 2528 1740 2529
rect 1790 2533 1796 2534
rect 1790 2529 1791 2533
rect 1795 2529 1796 2533
rect 1790 2528 1796 2529
rect 1846 2533 1852 2534
rect 1846 2529 1847 2533
rect 1851 2529 1852 2533
rect 1846 2528 1852 2529
rect 1902 2533 1908 2534
rect 1902 2529 1903 2533
rect 1907 2529 1908 2533
rect 1902 2528 1908 2529
rect 1958 2533 1964 2534
rect 1958 2529 1959 2533
rect 1963 2529 1964 2533
rect 1958 2528 1964 2529
rect 2014 2533 2020 2534
rect 2014 2529 2015 2533
rect 2019 2529 2020 2533
rect 2014 2528 2020 2529
rect 2070 2533 2076 2534
rect 2070 2529 2071 2533
rect 2075 2529 2076 2533
rect 2070 2528 2076 2529
rect 2126 2533 2132 2534
rect 2126 2529 2127 2533
rect 2131 2529 2132 2533
rect 2126 2528 2132 2529
rect 2182 2533 2188 2534
rect 2504 2533 2506 2553
rect 2182 2529 2183 2533
rect 2187 2529 2188 2533
rect 2502 2532 2508 2533
rect 2182 2528 2188 2529
rect 2190 2531 2196 2532
rect 2190 2527 2191 2531
rect 2195 2527 2196 2531
rect 2502 2528 2503 2532
rect 2507 2528 2508 2532
rect 2502 2527 2508 2528
rect 2190 2526 2196 2527
rect 1718 2512 1724 2513
rect 1718 2508 1719 2512
rect 1723 2508 1724 2512
rect 1718 2507 1724 2508
rect 1774 2512 1780 2513
rect 1774 2508 1775 2512
rect 1779 2508 1780 2512
rect 1774 2507 1780 2508
rect 1830 2512 1836 2513
rect 1830 2508 1831 2512
rect 1835 2508 1836 2512
rect 1830 2507 1836 2508
rect 1886 2512 1892 2513
rect 1886 2508 1887 2512
rect 1891 2508 1892 2512
rect 1886 2507 1892 2508
rect 1942 2512 1948 2513
rect 1942 2508 1943 2512
rect 1947 2508 1948 2512
rect 1942 2507 1948 2508
rect 1998 2512 2004 2513
rect 1998 2508 1999 2512
rect 2003 2508 2004 2512
rect 1998 2507 2004 2508
rect 2054 2512 2060 2513
rect 2054 2508 2055 2512
rect 2059 2508 2060 2512
rect 2054 2507 2060 2508
rect 2110 2512 2116 2513
rect 2110 2508 2111 2512
rect 2115 2508 2116 2512
rect 2110 2507 2116 2508
rect 2166 2512 2172 2513
rect 2166 2508 2167 2512
rect 2171 2508 2172 2512
rect 2166 2507 2172 2508
rect 1720 2499 1722 2507
rect 1776 2499 1778 2507
rect 1798 2499 1804 2500
rect 1832 2499 1834 2507
rect 1888 2499 1890 2507
rect 1944 2499 1946 2507
rect 2000 2499 2002 2507
rect 2056 2499 2058 2507
rect 2112 2499 2114 2507
rect 2168 2499 2170 2507
rect 2192 2500 2194 2526
rect 2502 2515 2508 2516
rect 2502 2511 2503 2515
rect 2507 2511 2508 2515
rect 2502 2510 2508 2511
rect 2190 2499 2196 2500
rect 2504 2499 2506 2510
rect 1719 2498 1723 2499
rect 1719 2493 1723 2494
rect 1775 2498 1779 2499
rect 1798 2495 1799 2499
rect 1803 2495 1804 2499
rect 1798 2494 1804 2495
rect 1831 2498 1835 2499
rect 1775 2493 1779 2494
rect 1774 2492 1780 2493
rect 1774 2488 1775 2492
rect 1779 2488 1780 2492
rect 1774 2487 1780 2488
rect 1326 2468 1327 2472
rect 1331 2468 1332 2472
rect 1326 2467 1332 2468
rect 1366 2471 1372 2472
rect 1366 2467 1367 2471
rect 1371 2467 1372 2471
rect 1158 2449 1159 2453
rect 1163 2449 1164 2453
rect 1286 2452 1292 2453
rect 1158 2448 1164 2449
rect 1182 2451 1188 2452
rect 1182 2447 1183 2451
rect 1187 2447 1188 2451
rect 1286 2448 1287 2452
rect 1291 2448 1292 2452
rect 1286 2447 1292 2448
rect 1182 2446 1188 2447
rect 774 2432 780 2433
rect 774 2428 775 2432
rect 779 2428 780 2432
rect 774 2427 780 2428
rect 862 2432 868 2433
rect 862 2428 863 2432
rect 867 2428 868 2432
rect 862 2427 868 2428
rect 950 2432 956 2433
rect 950 2428 951 2432
rect 955 2428 956 2432
rect 950 2427 956 2428
rect 1046 2432 1052 2433
rect 1046 2428 1047 2432
rect 1051 2428 1052 2432
rect 1046 2427 1052 2428
rect 1142 2432 1148 2433
rect 1142 2428 1143 2432
rect 1147 2428 1148 2432
rect 1142 2427 1148 2428
rect 776 2423 778 2427
rect 864 2423 866 2427
rect 952 2423 954 2427
rect 1048 2423 1050 2427
rect 1144 2423 1146 2427
rect 775 2422 779 2423
rect 775 2417 779 2418
rect 831 2422 835 2423
rect 831 2417 835 2418
rect 863 2422 867 2423
rect 863 2417 867 2418
rect 935 2422 939 2423
rect 935 2417 939 2418
rect 951 2422 955 2423
rect 951 2417 955 2418
rect 1039 2422 1043 2423
rect 1039 2417 1043 2418
rect 1047 2422 1051 2423
rect 1047 2417 1051 2418
rect 1143 2422 1147 2423
rect 1143 2417 1147 2418
rect 1151 2422 1155 2423
rect 1151 2417 1155 2418
rect 830 2416 836 2417
rect 830 2412 831 2416
rect 835 2412 836 2416
rect 830 2411 836 2412
rect 934 2416 940 2417
rect 934 2412 935 2416
rect 939 2412 940 2416
rect 934 2411 940 2412
rect 1038 2416 1044 2417
rect 1038 2412 1039 2416
rect 1043 2412 1044 2416
rect 1038 2411 1044 2412
rect 1150 2416 1156 2417
rect 1150 2412 1151 2416
rect 1155 2412 1156 2416
rect 1150 2411 1156 2412
rect 246 2395 252 2396
rect 246 2391 247 2395
rect 251 2391 252 2395
rect 246 2390 252 2391
rect 334 2395 340 2396
rect 334 2391 335 2395
rect 339 2391 340 2395
rect 334 2390 340 2391
rect 430 2395 436 2396
rect 430 2391 431 2395
rect 435 2391 436 2395
rect 430 2390 436 2391
rect 438 2395 444 2396
rect 438 2391 439 2395
rect 443 2391 444 2395
rect 438 2390 444 2391
rect 534 2395 540 2396
rect 534 2391 535 2395
rect 539 2391 540 2395
rect 534 2390 540 2391
rect 638 2395 644 2396
rect 638 2391 639 2395
rect 643 2391 644 2395
rect 638 2390 644 2391
rect 742 2395 748 2396
rect 742 2391 743 2395
rect 747 2391 748 2395
rect 742 2390 748 2391
rect 762 2395 768 2396
rect 762 2391 763 2395
rect 767 2391 768 2395
rect 762 2390 768 2391
rect 846 2395 852 2396
rect 846 2391 847 2395
rect 851 2391 852 2395
rect 846 2390 852 2391
rect 950 2395 956 2396
rect 950 2391 951 2395
rect 955 2391 956 2395
rect 950 2390 956 2391
rect 1054 2395 1060 2396
rect 1054 2391 1055 2395
rect 1059 2391 1060 2395
rect 1054 2390 1060 2391
rect 1166 2395 1172 2396
rect 1166 2391 1167 2395
rect 1171 2391 1172 2395
rect 1166 2390 1172 2391
rect 1174 2395 1180 2396
rect 1174 2391 1175 2395
rect 1179 2391 1180 2395
rect 1174 2390 1180 2391
rect 190 2379 196 2380
rect 190 2375 191 2379
rect 195 2375 196 2379
rect 190 2374 196 2375
rect 248 2371 250 2390
rect 336 2371 338 2390
rect 432 2371 434 2390
rect 111 2370 115 2371
rect 111 2365 115 2366
rect 167 2370 171 2371
rect 167 2365 171 2366
rect 175 2370 179 2371
rect 175 2365 179 2366
rect 247 2370 251 2371
rect 247 2365 251 2366
rect 279 2370 283 2371
rect 279 2365 283 2366
rect 335 2370 339 2371
rect 335 2365 339 2366
rect 391 2370 395 2371
rect 391 2365 395 2366
rect 431 2370 435 2371
rect 440 2368 442 2390
rect 536 2371 538 2390
rect 630 2375 636 2376
rect 630 2371 631 2375
rect 635 2371 636 2375
rect 640 2371 642 2390
rect 744 2371 746 2390
rect 848 2371 850 2390
rect 952 2371 954 2390
rect 1056 2371 1058 2390
rect 1168 2371 1170 2390
rect 503 2370 507 2371
rect 431 2365 435 2366
rect 438 2367 444 2368
rect 112 2345 114 2365
rect 176 2346 178 2365
rect 280 2346 282 2365
rect 392 2346 394 2365
rect 438 2363 439 2367
rect 443 2363 444 2367
rect 503 2365 507 2366
rect 535 2370 539 2371
rect 535 2365 539 2366
rect 623 2370 627 2371
rect 630 2370 636 2371
rect 639 2370 643 2371
rect 623 2365 627 2366
rect 438 2362 444 2363
rect 504 2346 506 2365
rect 624 2346 626 2365
rect 174 2345 180 2346
rect 110 2344 116 2345
rect 110 2340 111 2344
rect 115 2340 116 2344
rect 174 2341 175 2345
rect 179 2341 180 2345
rect 174 2340 180 2341
rect 278 2345 284 2346
rect 278 2341 279 2345
rect 283 2341 284 2345
rect 278 2340 284 2341
rect 390 2345 396 2346
rect 390 2341 391 2345
rect 395 2341 396 2345
rect 390 2340 396 2341
rect 502 2345 508 2346
rect 502 2341 503 2345
rect 507 2341 508 2345
rect 622 2345 628 2346
rect 502 2340 508 2341
rect 510 2343 516 2344
rect 110 2339 116 2340
rect 510 2339 511 2343
rect 515 2339 516 2343
rect 622 2341 623 2345
rect 627 2341 628 2345
rect 632 2344 634 2370
rect 639 2365 643 2366
rect 743 2370 747 2371
rect 743 2365 747 2366
rect 847 2370 851 2371
rect 847 2365 851 2366
rect 871 2370 875 2371
rect 871 2365 875 2366
rect 951 2370 955 2371
rect 951 2365 955 2366
rect 999 2370 1003 2371
rect 999 2365 1003 2366
rect 1055 2370 1059 2371
rect 1055 2365 1059 2366
rect 1127 2370 1131 2371
rect 1167 2370 1171 2371
rect 1127 2365 1131 2366
rect 1146 2367 1152 2368
rect 744 2346 746 2365
rect 770 2359 776 2360
rect 770 2355 771 2359
rect 775 2355 776 2359
rect 770 2354 776 2355
rect 742 2345 748 2346
rect 622 2340 628 2341
rect 630 2343 636 2344
rect 510 2338 516 2339
rect 630 2339 631 2343
rect 635 2339 636 2343
rect 742 2341 743 2345
rect 747 2341 748 2345
rect 742 2340 748 2341
rect 630 2338 636 2339
rect 110 2327 116 2328
rect 110 2323 111 2327
rect 115 2323 116 2327
rect 110 2322 116 2323
rect 158 2324 164 2325
rect 112 2315 114 2322
rect 158 2320 159 2324
rect 163 2320 164 2324
rect 158 2319 164 2320
rect 262 2324 268 2325
rect 262 2320 263 2324
rect 267 2320 268 2324
rect 262 2319 268 2320
rect 374 2324 380 2325
rect 374 2320 375 2324
rect 379 2320 380 2324
rect 374 2319 380 2320
rect 486 2324 492 2325
rect 486 2320 487 2324
rect 491 2320 492 2324
rect 486 2319 492 2320
rect 160 2315 162 2319
rect 264 2315 266 2319
rect 376 2315 378 2319
rect 488 2315 490 2319
rect 111 2314 115 2315
rect 111 2309 115 2310
rect 159 2314 163 2315
rect 159 2309 163 2310
rect 207 2314 211 2315
rect 207 2309 211 2310
rect 263 2314 267 2315
rect 263 2309 267 2310
rect 287 2314 291 2315
rect 287 2309 291 2310
rect 375 2314 379 2315
rect 375 2309 379 2310
rect 471 2314 475 2315
rect 471 2309 475 2310
rect 487 2314 491 2315
rect 487 2309 491 2310
rect 112 2306 114 2309
rect 206 2308 212 2309
rect 110 2305 116 2306
rect 110 2301 111 2305
rect 115 2301 116 2305
rect 206 2304 207 2308
rect 211 2304 212 2308
rect 206 2303 212 2304
rect 286 2308 292 2309
rect 286 2304 287 2308
rect 291 2304 292 2308
rect 286 2303 292 2304
rect 374 2308 380 2309
rect 374 2304 375 2308
rect 379 2304 380 2308
rect 374 2303 380 2304
rect 470 2308 476 2309
rect 470 2304 471 2308
rect 475 2304 476 2308
rect 470 2303 476 2304
rect 110 2300 116 2301
rect 110 2288 116 2289
rect 110 2284 111 2288
rect 115 2284 116 2288
rect 110 2283 116 2284
rect 222 2287 228 2288
rect 222 2283 223 2287
rect 227 2283 228 2287
rect 112 2259 114 2283
rect 222 2282 228 2283
rect 302 2287 308 2288
rect 302 2283 303 2287
rect 307 2283 308 2287
rect 302 2282 308 2283
rect 390 2287 396 2288
rect 390 2283 391 2287
rect 395 2283 396 2287
rect 390 2282 396 2283
rect 486 2287 492 2288
rect 486 2283 487 2287
rect 491 2283 492 2287
rect 486 2282 492 2283
rect 494 2287 500 2288
rect 494 2283 495 2287
rect 499 2283 500 2287
rect 494 2282 500 2283
rect 224 2259 226 2282
rect 304 2259 306 2282
rect 392 2259 394 2282
rect 488 2259 490 2282
rect 111 2258 115 2259
rect 111 2253 115 2254
rect 223 2258 227 2259
rect 223 2253 227 2254
rect 263 2258 267 2259
rect 263 2253 267 2254
rect 303 2258 307 2259
rect 303 2253 307 2254
rect 319 2258 323 2259
rect 319 2253 323 2254
rect 383 2258 387 2259
rect 383 2253 387 2254
rect 391 2258 395 2259
rect 391 2253 395 2254
rect 447 2258 451 2259
rect 447 2253 451 2254
rect 487 2258 491 2259
rect 496 2256 498 2282
rect 512 2268 514 2338
rect 606 2324 612 2325
rect 606 2320 607 2324
rect 611 2320 612 2324
rect 606 2319 612 2320
rect 726 2324 732 2325
rect 726 2320 727 2324
rect 731 2320 732 2324
rect 726 2319 732 2320
rect 608 2315 610 2319
rect 728 2315 730 2319
rect 559 2314 563 2315
rect 559 2309 563 2310
rect 607 2314 611 2315
rect 607 2309 611 2310
rect 647 2314 651 2315
rect 647 2309 651 2310
rect 727 2314 731 2315
rect 727 2309 731 2310
rect 735 2314 739 2315
rect 735 2309 739 2310
rect 558 2308 564 2309
rect 558 2304 559 2308
rect 563 2304 564 2308
rect 558 2303 564 2304
rect 646 2308 652 2309
rect 646 2304 647 2308
rect 651 2304 652 2308
rect 646 2303 652 2304
rect 734 2308 740 2309
rect 734 2304 735 2308
rect 739 2304 740 2308
rect 734 2303 740 2304
rect 772 2288 774 2354
rect 872 2346 874 2365
rect 1000 2346 1002 2365
rect 1128 2346 1130 2365
rect 1146 2363 1147 2367
rect 1151 2363 1152 2367
rect 1167 2365 1171 2366
rect 1146 2362 1152 2363
rect 870 2345 876 2346
rect 870 2341 871 2345
rect 875 2341 876 2345
rect 870 2340 876 2341
rect 998 2345 1004 2346
rect 998 2341 999 2345
rect 1003 2341 1004 2345
rect 1126 2345 1132 2346
rect 998 2340 1004 2341
rect 1014 2343 1020 2344
rect 1014 2339 1015 2343
rect 1019 2339 1020 2343
rect 1126 2341 1127 2345
rect 1131 2341 1132 2345
rect 1148 2344 1150 2362
rect 1176 2360 1178 2390
rect 1184 2376 1186 2446
rect 1328 2439 1330 2467
rect 1366 2466 1372 2467
rect 1438 2471 1444 2472
rect 1438 2467 1439 2471
rect 1443 2467 1444 2471
rect 1438 2466 1444 2467
rect 1526 2471 1532 2472
rect 1526 2467 1527 2471
rect 1531 2467 1532 2471
rect 1526 2466 1532 2467
rect 1614 2471 1620 2472
rect 1614 2467 1615 2471
rect 1619 2467 1620 2471
rect 1614 2466 1620 2467
rect 1702 2471 1708 2472
rect 1702 2467 1703 2471
rect 1707 2467 1708 2471
rect 1702 2466 1708 2467
rect 1710 2471 1716 2472
rect 1710 2467 1711 2471
rect 1715 2467 1716 2471
rect 1710 2466 1716 2467
rect 1790 2471 1796 2472
rect 1790 2467 1791 2471
rect 1795 2467 1796 2471
rect 1790 2466 1796 2467
rect 1368 2439 1370 2466
rect 1440 2439 1442 2466
rect 1528 2439 1530 2466
rect 1616 2439 1618 2466
rect 1658 2451 1664 2452
rect 1658 2447 1659 2451
rect 1663 2447 1664 2451
rect 1658 2446 1664 2447
rect 1327 2438 1331 2439
rect 1286 2435 1292 2436
rect 1286 2431 1287 2435
rect 1291 2431 1292 2435
rect 1327 2433 1331 2434
rect 1367 2438 1371 2439
rect 1367 2433 1371 2434
rect 1439 2438 1443 2439
rect 1439 2433 1443 2434
rect 1527 2438 1531 2439
rect 1527 2433 1531 2434
rect 1543 2438 1547 2439
rect 1543 2433 1547 2434
rect 1615 2438 1619 2439
rect 1615 2433 1619 2434
rect 1639 2438 1643 2439
rect 1639 2433 1643 2434
rect 1286 2430 1292 2431
rect 1288 2423 1290 2430
rect 1287 2422 1291 2423
rect 1287 2417 1291 2418
rect 1288 2414 1290 2417
rect 1286 2413 1292 2414
rect 1328 2413 1330 2433
rect 1368 2414 1370 2433
rect 1374 2427 1380 2428
rect 1374 2423 1375 2427
rect 1379 2423 1380 2427
rect 1374 2422 1380 2423
rect 1366 2413 1372 2414
rect 1286 2409 1287 2413
rect 1291 2409 1292 2413
rect 1286 2408 1292 2409
rect 1326 2412 1332 2413
rect 1326 2408 1327 2412
rect 1331 2408 1332 2412
rect 1366 2409 1367 2413
rect 1371 2409 1372 2413
rect 1366 2408 1372 2409
rect 1326 2407 1332 2408
rect 1286 2396 1292 2397
rect 1286 2392 1287 2396
rect 1291 2392 1292 2396
rect 1286 2391 1292 2392
rect 1326 2395 1332 2396
rect 1326 2391 1327 2395
rect 1331 2391 1332 2395
rect 1182 2375 1188 2376
rect 1182 2371 1183 2375
rect 1187 2371 1188 2375
rect 1288 2371 1290 2391
rect 1326 2390 1332 2391
rect 1350 2392 1356 2393
rect 1328 2379 1330 2390
rect 1350 2388 1351 2392
rect 1355 2388 1356 2392
rect 1350 2387 1356 2388
rect 1352 2379 1354 2387
rect 1327 2378 1331 2379
rect 1327 2373 1331 2374
rect 1351 2378 1355 2379
rect 1351 2373 1355 2374
rect 1182 2370 1188 2371
rect 1287 2370 1291 2371
rect 1328 2370 1330 2373
rect 1350 2372 1356 2373
rect 1287 2365 1291 2366
rect 1326 2369 1332 2370
rect 1326 2365 1327 2369
rect 1331 2365 1332 2369
rect 1350 2368 1351 2372
rect 1355 2368 1356 2372
rect 1350 2367 1356 2368
rect 1174 2359 1180 2360
rect 1174 2355 1175 2359
rect 1179 2355 1180 2359
rect 1174 2354 1180 2355
rect 1288 2345 1290 2365
rect 1326 2364 1332 2365
rect 1326 2352 1332 2353
rect 1376 2352 1378 2422
rect 1440 2414 1442 2433
rect 1544 2414 1546 2433
rect 1640 2414 1642 2433
rect 1438 2413 1444 2414
rect 1438 2409 1439 2413
rect 1443 2409 1444 2413
rect 1438 2408 1444 2409
rect 1542 2413 1548 2414
rect 1542 2409 1543 2413
rect 1547 2409 1548 2413
rect 1542 2408 1548 2409
rect 1638 2413 1644 2414
rect 1638 2409 1639 2413
rect 1643 2409 1644 2413
rect 1660 2412 1662 2446
rect 1704 2439 1706 2466
rect 1792 2439 1794 2466
rect 1800 2456 1802 2494
rect 1831 2493 1835 2494
rect 1863 2498 1867 2499
rect 1863 2493 1867 2494
rect 1887 2498 1891 2499
rect 1887 2493 1891 2494
rect 1943 2498 1947 2499
rect 1943 2493 1947 2494
rect 1951 2498 1955 2499
rect 1951 2493 1955 2494
rect 1999 2498 2003 2499
rect 1999 2493 2003 2494
rect 2039 2498 2043 2499
rect 2039 2493 2043 2494
rect 2055 2498 2059 2499
rect 2055 2493 2059 2494
rect 2111 2498 2115 2499
rect 2111 2493 2115 2494
rect 2127 2498 2131 2499
rect 2127 2493 2131 2494
rect 2167 2498 2171 2499
rect 2190 2495 2191 2499
rect 2195 2495 2196 2499
rect 2190 2494 2196 2495
rect 2503 2498 2507 2499
rect 2167 2493 2171 2494
rect 2503 2493 2507 2494
rect 1862 2492 1868 2493
rect 1862 2488 1863 2492
rect 1867 2488 1868 2492
rect 1862 2487 1868 2488
rect 1950 2492 1956 2493
rect 1950 2488 1951 2492
rect 1955 2488 1956 2492
rect 1950 2487 1956 2488
rect 2038 2492 2044 2493
rect 2038 2488 2039 2492
rect 2043 2488 2044 2492
rect 2038 2487 2044 2488
rect 2126 2492 2132 2493
rect 2126 2488 2127 2492
rect 2131 2488 2132 2492
rect 2504 2490 2506 2493
rect 2126 2487 2132 2488
rect 2502 2489 2508 2490
rect 2502 2485 2503 2489
rect 2507 2485 2508 2489
rect 2502 2484 2508 2485
rect 2502 2472 2508 2473
rect 1878 2471 1884 2472
rect 1878 2467 1879 2471
rect 1883 2467 1884 2471
rect 1878 2466 1884 2467
rect 1966 2471 1972 2472
rect 1966 2467 1967 2471
rect 1971 2467 1972 2471
rect 1966 2466 1972 2467
rect 2054 2471 2060 2472
rect 2054 2467 2055 2471
rect 2059 2467 2060 2471
rect 2054 2466 2060 2467
rect 2142 2471 2148 2472
rect 2142 2467 2143 2471
rect 2147 2467 2148 2471
rect 2142 2466 2148 2467
rect 2150 2471 2156 2472
rect 2150 2467 2151 2471
rect 2155 2467 2156 2471
rect 2502 2468 2503 2472
rect 2507 2468 2508 2472
rect 2502 2467 2508 2468
rect 2150 2466 2156 2467
rect 1798 2455 1804 2456
rect 1798 2451 1799 2455
rect 1803 2451 1804 2455
rect 1798 2450 1804 2451
rect 1880 2439 1882 2466
rect 1968 2439 1970 2466
rect 2056 2439 2058 2466
rect 2144 2439 2146 2466
rect 1703 2438 1707 2439
rect 1703 2433 1707 2434
rect 1735 2438 1739 2439
rect 1735 2433 1739 2434
rect 1791 2438 1795 2439
rect 1791 2433 1795 2434
rect 1823 2438 1827 2439
rect 1823 2433 1827 2434
rect 1879 2438 1883 2439
rect 1879 2433 1883 2434
rect 1911 2438 1915 2439
rect 1911 2433 1915 2434
rect 1967 2438 1971 2439
rect 1967 2433 1971 2434
rect 2007 2438 2011 2439
rect 2007 2433 2011 2434
rect 2055 2438 2059 2439
rect 2055 2433 2059 2434
rect 2103 2438 2107 2439
rect 2103 2433 2107 2434
rect 2143 2438 2147 2439
rect 2143 2433 2147 2434
rect 1736 2414 1738 2433
rect 1824 2414 1826 2433
rect 1912 2414 1914 2433
rect 2008 2414 2010 2433
rect 2104 2414 2106 2433
rect 2152 2428 2154 2466
rect 2504 2439 2506 2467
rect 2503 2438 2507 2439
rect 2503 2433 2507 2434
rect 2150 2427 2156 2428
rect 2150 2423 2151 2427
rect 2155 2423 2156 2427
rect 2150 2422 2156 2423
rect 1734 2413 1740 2414
rect 1638 2408 1644 2409
rect 1658 2411 1664 2412
rect 1658 2407 1659 2411
rect 1663 2407 1664 2411
rect 1734 2409 1735 2413
rect 1739 2409 1740 2413
rect 1822 2413 1828 2414
rect 1734 2408 1740 2409
rect 1758 2411 1764 2412
rect 1658 2406 1664 2407
rect 1758 2407 1759 2411
rect 1763 2407 1764 2411
rect 1822 2409 1823 2413
rect 1827 2409 1828 2413
rect 1822 2408 1828 2409
rect 1910 2413 1916 2414
rect 1910 2409 1911 2413
rect 1915 2409 1916 2413
rect 1910 2408 1916 2409
rect 2006 2413 2012 2414
rect 2006 2409 2007 2413
rect 2011 2409 2012 2413
rect 2006 2408 2012 2409
rect 2102 2413 2108 2414
rect 2504 2413 2506 2433
rect 2102 2409 2103 2413
rect 2107 2409 2108 2413
rect 2102 2408 2108 2409
rect 2502 2412 2508 2413
rect 2502 2408 2503 2412
rect 2507 2408 2508 2412
rect 2502 2407 2508 2408
rect 1758 2406 1764 2407
rect 1422 2392 1428 2393
rect 1422 2388 1423 2392
rect 1427 2388 1428 2392
rect 1422 2387 1428 2388
rect 1526 2392 1532 2393
rect 1526 2388 1527 2392
rect 1531 2388 1532 2392
rect 1526 2387 1532 2388
rect 1622 2392 1628 2393
rect 1622 2388 1623 2392
rect 1627 2388 1628 2392
rect 1622 2387 1628 2388
rect 1718 2392 1724 2393
rect 1718 2388 1719 2392
rect 1723 2388 1724 2392
rect 1718 2387 1724 2388
rect 1424 2379 1426 2387
rect 1528 2379 1530 2387
rect 1624 2379 1626 2387
rect 1720 2379 1722 2387
rect 1407 2378 1411 2379
rect 1407 2373 1411 2374
rect 1423 2378 1427 2379
rect 1423 2373 1427 2374
rect 1495 2378 1499 2379
rect 1495 2373 1499 2374
rect 1527 2378 1531 2379
rect 1527 2373 1531 2374
rect 1583 2378 1587 2379
rect 1583 2373 1587 2374
rect 1623 2378 1627 2379
rect 1623 2373 1627 2374
rect 1671 2378 1675 2379
rect 1671 2373 1675 2374
rect 1719 2378 1723 2379
rect 1719 2373 1723 2374
rect 1751 2378 1755 2379
rect 1751 2373 1755 2374
rect 1406 2372 1412 2373
rect 1406 2368 1407 2372
rect 1411 2368 1412 2372
rect 1406 2367 1412 2368
rect 1494 2372 1500 2373
rect 1494 2368 1495 2372
rect 1499 2368 1500 2372
rect 1494 2367 1500 2368
rect 1582 2372 1588 2373
rect 1582 2368 1583 2372
rect 1587 2368 1588 2372
rect 1582 2367 1588 2368
rect 1670 2372 1676 2373
rect 1670 2368 1671 2372
rect 1675 2368 1676 2372
rect 1670 2367 1676 2368
rect 1750 2372 1756 2373
rect 1750 2368 1751 2372
rect 1755 2368 1756 2372
rect 1750 2367 1756 2368
rect 1326 2348 1327 2352
rect 1331 2348 1332 2352
rect 1326 2347 1332 2348
rect 1366 2351 1372 2352
rect 1366 2347 1367 2351
rect 1371 2347 1372 2351
rect 1286 2344 1292 2345
rect 1126 2340 1132 2341
rect 1146 2343 1152 2344
rect 1014 2338 1020 2339
rect 1146 2339 1147 2343
rect 1151 2339 1152 2343
rect 1286 2340 1287 2344
rect 1291 2340 1292 2344
rect 1286 2339 1292 2340
rect 1146 2338 1152 2339
rect 854 2324 860 2325
rect 854 2320 855 2324
rect 859 2320 860 2324
rect 854 2319 860 2320
rect 982 2324 988 2325
rect 982 2320 983 2324
rect 987 2320 988 2324
rect 982 2319 988 2320
rect 856 2315 858 2319
rect 984 2315 986 2319
rect 815 2314 819 2315
rect 815 2309 819 2310
rect 855 2314 859 2315
rect 855 2309 859 2310
rect 903 2314 907 2315
rect 903 2309 907 2310
rect 983 2314 987 2315
rect 983 2309 987 2310
rect 991 2314 995 2315
rect 991 2309 995 2310
rect 814 2308 820 2309
rect 814 2304 815 2308
rect 819 2304 820 2308
rect 814 2303 820 2304
rect 902 2308 908 2309
rect 902 2304 903 2308
rect 907 2304 908 2308
rect 902 2303 908 2304
rect 990 2308 996 2309
rect 990 2304 991 2308
rect 995 2304 996 2308
rect 990 2303 996 2304
rect 574 2287 580 2288
rect 574 2283 575 2287
rect 579 2283 580 2287
rect 574 2282 580 2283
rect 662 2287 668 2288
rect 662 2283 663 2287
rect 667 2283 668 2287
rect 662 2282 668 2283
rect 750 2287 756 2288
rect 750 2283 751 2287
rect 755 2283 756 2287
rect 750 2282 756 2283
rect 770 2287 776 2288
rect 770 2283 771 2287
rect 775 2283 776 2287
rect 770 2282 776 2283
rect 830 2287 836 2288
rect 830 2283 831 2287
rect 835 2283 836 2287
rect 830 2282 836 2283
rect 918 2287 924 2288
rect 918 2283 919 2287
rect 923 2283 924 2287
rect 918 2282 924 2283
rect 974 2287 980 2288
rect 974 2283 975 2287
rect 979 2283 980 2287
rect 974 2282 980 2283
rect 1006 2287 1012 2288
rect 1006 2283 1007 2287
rect 1011 2283 1012 2287
rect 1006 2282 1012 2283
rect 510 2267 516 2268
rect 510 2263 511 2267
rect 515 2263 516 2267
rect 510 2262 516 2263
rect 576 2259 578 2282
rect 582 2271 588 2272
rect 582 2267 583 2271
rect 587 2267 588 2271
rect 582 2266 588 2267
rect 503 2258 507 2259
rect 487 2253 491 2254
rect 494 2255 500 2256
rect 112 2233 114 2253
rect 264 2234 266 2253
rect 320 2234 322 2253
rect 384 2234 386 2253
rect 448 2234 450 2253
rect 494 2251 495 2255
rect 499 2251 500 2255
rect 503 2253 507 2254
rect 559 2258 563 2259
rect 559 2253 563 2254
rect 575 2258 579 2259
rect 575 2253 579 2254
rect 494 2250 500 2251
rect 504 2234 506 2253
rect 560 2234 562 2253
rect 262 2233 268 2234
rect 110 2232 116 2233
rect 110 2228 111 2232
rect 115 2228 116 2232
rect 262 2229 263 2233
rect 267 2229 268 2233
rect 262 2228 268 2229
rect 318 2233 324 2234
rect 318 2229 319 2233
rect 323 2229 324 2233
rect 318 2228 324 2229
rect 382 2233 388 2234
rect 382 2229 383 2233
rect 387 2229 388 2233
rect 382 2228 388 2229
rect 446 2233 452 2234
rect 446 2229 447 2233
rect 451 2229 452 2233
rect 446 2228 452 2229
rect 502 2233 508 2234
rect 502 2229 503 2233
rect 507 2229 508 2233
rect 558 2233 564 2234
rect 502 2228 508 2229
rect 510 2231 516 2232
rect 110 2227 116 2228
rect 510 2227 511 2231
rect 515 2227 516 2231
rect 558 2229 559 2233
rect 563 2229 564 2233
rect 584 2232 586 2266
rect 664 2259 666 2282
rect 752 2259 754 2282
rect 832 2259 834 2282
rect 920 2259 922 2282
rect 615 2258 619 2259
rect 615 2253 619 2254
rect 663 2258 667 2259
rect 663 2253 667 2254
rect 671 2258 675 2259
rect 671 2253 675 2254
rect 727 2258 731 2259
rect 727 2253 731 2254
rect 751 2258 755 2259
rect 751 2253 755 2254
rect 791 2258 795 2259
rect 791 2253 795 2254
rect 831 2258 835 2259
rect 831 2253 835 2254
rect 855 2258 859 2259
rect 855 2253 859 2254
rect 919 2258 923 2259
rect 919 2253 923 2254
rect 616 2234 618 2253
rect 672 2234 674 2253
rect 728 2234 730 2253
rect 792 2234 794 2253
rect 856 2234 858 2253
rect 920 2234 922 2253
rect 976 2248 978 2282
rect 1008 2259 1010 2282
rect 1016 2272 1018 2338
rect 1286 2327 1292 2328
rect 1110 2324 1116 2325
rect 1110 2320 1111 2324
rect 1115 2320 1116 2324
rect 1286 2323 1287 2327
rect 1291 2323 1292 2327
rect 1328 2323 1330 2347
rect 1366 2346 1372 2347
rect 1374 2351 1380 2352
rect 1374 2347 1375 2351
rect 1379 2347 1380 2351
rect 1374 2346 1380 2347
rect 1422 2351 1428 2352
rect 1422 2347 1423 2351
rect 1427 2347 1428 2351
rect 1422 2346 1428 2347
rect 1510 2351 1516 2352
rect 1510 2347 1511 2351
rect 1515 2347 1516 2351
rect 1510 2346 1516 2347
rect 1598 2351 1604 2352
rect 1598 2347 1599 2351
rect 1603 2347 1604 2351
rect 1598 2346 1604 2347
rect 1686 2351 1692 2352
rect 1686 2347 1687 2351
rect 1691 2347 1692 2351
rect 1686 2346 1692 2347
rect 1694 2351 1700 2352
rect 1694 2347 1695 2351
rect 1699 2347 1700 2351
rect 1694 2346 1700 2347
rect 1368 2323 1370 2346
rect 1424 2323 1426 2346
rect 1512 2323 1514 2346
rect 1566 2335 1572 2336
rect 1566 2331 1567 2335
rect 1571 2331 1572 2335
rect 1566 2330 1572 2331
rect 1286 2322 1292 2323
rect 1327 2322 1331 2323
rect 1110 2319 1116 2320
rect 1112 2315 1114 2319
rect 1288 2315 1290 2322
rect 1327 2317 1331 2318
rect 1367 2322 1371 2323
rect 1367 2317 1371 2318
rect 1423 2322 1427 2323
rect 1423 2317 1427 2318
rect 1455 2322 1459 2323
rect 1455 2317 1459 2318
rect 1511 2322 1515 2323
rect 1511 2317 1515 2318
rect 1543 2322 1547 2323
rect 1543 2317 1547 2318
rect 1079 2314 1083 2315
rect 1079 2309 1083 2310
rect 1111 2314 1115 2315
rect 1111 2309 1115 2310
rect 1287 2314 1291 2315
rect 1287 2309 1291 2310
rect 1078 2308 1084 2309
rect 1078 2304 1079 2308
rect 1083 2304 1084 2308
rect 1288 2306 1290 2309
rect 1078 2303 1084 2304
rect 1286 2305 1292 2306
rect 1286 2301 1287 2305
rect 1291 2301 1292 2305
rect 1286 2300 1292 2301
rect 1328 2297 1330 2317
rect 1368 2298 1370 2317
rect 1456 2298 1458 2317
rect 1544 2298 1546 2317
rect 1366 2297 1372 2298
rect 1326 2296 1332 2297
rect 1326 2292 1327 2296
rect 1331 2292 1332 2296
rect 1366 2293 1367 2297
rect 1371 2293 1372 2297
rect 1366 2292 1372 2293
rect 1454 2297 1460 2298
rect 1454 2293 1455 2297
rect 1459 2293 1460 2297
rect 1454 2292 1460 2293
rect 1542 2297 1548 2298
rect 1542 2293 1543 2297
rect 1547 2293 1548 2297
rect 1568 2296 1570 2330
rect 1600 2323 1602 2346
rect 1688 2323 1690 2346
rect 1696 2328 1698 2346
rect 1760 2336 1762 2406
rect 2502 2395 2508 2396
rect 1806 2392 1812 2393
rect 1806 2388 1807 2392
rect 1811 2388 1812 2392
rect 1806 2387 1812 2388
rect 1894 2392 1900 2393
rect 1894 2388 1895 2392
rect 1899 2388 1900 2392
rect 1894 2387 1900 2388
rect 1990 2392 1996 2393
rect 1990 2388 1991 2392
rect 1995 2388 1996 2392
rect 1990 2387 1996 2388
rect 2086 2392 2092 2393
rect 2086 2388 2087 2392
rect 2091 2388 2092 2392
rect 2502 2391 2503 2395
rect 2507 2391 2508 2395
rect 2502 2390 2508 2391
rect 2086 2387 2092 2388
rect 1808 2379 1810 2387
rect 1896 2379 1898 2387
rect 1992 2379 1994 2387
rect 2088 2379 2090 2387
rect 2504 2379 2506 2390
rect 1807 2378 1811 2379
rect 1807 2373 1811 2374
rect 1831 2378 1835 2379
rect 1831 2373 1835 2374
rect 1895 2378 1899 2379
rect 1895 2373 1899 2374
rect 1919 2378 1923 2379
rect 1919 2373 1923 2374
rect 1991 2378 1995 2379
rect 1991 2373 1995 2374
rect 2007 2378 2011 2379
rect 2007 2373 2011 2374
rect 2087 2378 2091 2379
rect 2087 2373 2091 2374
rect 2095 2378 2099 2379
rect 2095 2373 2099 2374
rect 2503 2378 2507 2379
rect 2503 2373 2507 2374
rect 1830 2372 1836 2373
rect 1830 2368 1831 2372
rect 1835 2368 1836 2372
rect 1830 2367 1836 2368
rect 1918 2372 1924 2373
rect 1918 2368 1919 2372
rect 1923 2368 1924 2372
rect 1918 2367 1924 2368
rect 2006 2372 2012 2373
rect 2006 2368 2007 2372
rect 2011 2368 2012 2372
rect 2006 2367 2012 2368
rect 2094 2372 2100 2373
rect 2094 2368 2095 2372
rect 2099 2368 2100 2372
rect 2504 2370 2506 2373
rect 2094 2367 2100 2368
rect 2502 2369 2508 2370
rect 2502 2365 2503 2369
rect 2507 2365 2508 2369
rect 2502 2364 2508 2365
rect 2502 2352 2508 2353
rect 1766 2351 1772 2352
rect 1766 2347 1767 2351
rect 1771 2347 1772 2351
rect 1766 2346 1772 2347
rect 1846 2351 1852 2352
rect 1846 2347 1847 2351
rect 1851 2347 1852 2351
rect 1846 2346 1852 2347
rect 1934 2351 1940 2352
rect 1934 2347 1935 2351
rect 1939 2347 1940 2351
rect 1934 2346 1940 2347
rect 2022 2351 2028 2352
rect 2022 2347 2023 2351
rect 2027 2347 2028 2351
rect 2022 2346 2028 2347
rect 2110 2351 2116 2352
rect 2110 2347 2111 2351
rect 2115 2347 2116 2351
rect 2110 2346 2116 2347
rect 2118 2351 2124 2352
rect 2118 2347 2119 2351
rect 2123 2347 2124 2351
rect 2502 2348 2503 2352
rect 2507 2348 2508 2352
rect 2502 2347 2508 2348
rect 2118 2346 2124 2347
rect 1758 2335 1764 2336
rect 1758 2331 1759 2335
rect 1763 2331 1764 2335
rect 1758 2330 1764 2331
rect 1694 2327 1700 2328
rect 1694 2323 1695 2327
rect 1699 2323 1700 2327
rect 1768 2323 1770 2346
rect 1848 2323 1850 2346
rect 1936 2323 1938 2346
rect 2024 2323 2026 2346
rect 2112 2323 2114 2346
rect 1599 2322 1603 2323
rect 1599 2317 1603 2318
rect 1639 2322 1643 2323
rect 1687 2322 1691 2323
rect 1694 2322 1700 2323
rect 1735 2322 1739 2323
rect 1639 2317 1643 2318
rect 1658 2319 1664 2320
rect 1640 2298 1642 2317
rect 1658 2315 1659 2319
rect 1663 2315 1664 2319
rect 1687 2317 1691 2318
rect 1735 2317 1739 2318
rect 1767 2322 1771 2323
rect 1767 2317 1771 2318
rect 1831 2322 1835 2323
rect 1831 2317 1835 2318
rect 1847 2322 1851 2323
rect 1847 2317 1851 2318
rect 1927 2322 1931 2323
rect 1927 2317 1931 2318
rect 1935 2322 1939 2323
rect 1935 2317 1939 2318
rect 2015 2322 2019 2323
rect 2015 2317 2019 2318
rect 2023 2322 2027 2323
rect 2023 2317 2027 2318
rect 2111 2322 2115 2323
rect 2120 2320 2122 2346
rect 2504 2323 2506 2347
rect 2207 2322 2211 2323
rect 2111 2317 2115 2318
rect 2118 2319 2124 2320
rect 1658 2314 1664 2315
rect 1638 2297 1644 2298
rect 1542 2292 1548 2293
rect 1566 2295 1572 2296
rect 1326 2291 1332 2292
rect 1566 2291 1567 2295
rect 1571 2291 1572 2295
rect 1638 2293 1639 2297
rect 1643 2293 1644 2297
rect 1660 2296 1662 2314
rect 1736 2298 1738 2317
rect 1822 2311 1828 2312
rect 1822 2307 1823 2311
rect 1827 2307 1828 2311
rect 1822 2306 1828 2307
rect 1734 2297 1740 2298
rect 1638 2292 1644 2293
rect 1658 2295 1664 2296
rect 1566 2290 1572 2291
rect 1658 2291 1659 2295
rect 1663 2291 1664 2295
rect 1734 2293 1735 2297
rect 1739 2293 1740 2297
rect 1734 2292 1740 2293
rect 1658 2290 1664 2291
rect 1286 2288 1292 2289
rect 1094 2287 1100 2288
rect 1094 2283 1095 2287
rect 1099 2283 1100 2287
rect 1094 2282 1100 2283
rect 1102 2287 1108 2288
rect 1102 2283 1103 2287
rect 1107 2283 1108 2287
rect 1286 2284 1287 2288
rect 1291 2284 1292 2288
rect 1286 2283 1292 2284
rect 1102 2282 1108 2283
rect 1014 2271 1020 2272
rect 1014 2267 1015 2271
rect 1019 2267 1020 2271
rect 1014 2266 1020 2267
rect 1096 2259 1098 2282
rect 1104 2264 1106 2282
rect 1102 2263 1108 2264
rect 1102 2259 1103 2263
rect 1107 2259 1108 2263
rect 1288 2259 1290 2283
rect 1326 2279 1332 2280
rect 1326 2275 1327 2279
rect 1331 2275 1332 2279
rect 1326 2274 1332 2275
rect 1350 2276 1356 2277
rect 1328 2271 1330 2274
rect 1350 2272 1351 2276
rect 1355 2272 1356 2276
rect 1350 2271 1356 2272
rect 1438 2276 1444 2277
rect 1438 2272 1439 2276
rect 1443 2272 1444 2276
rect 1438 2271 1444 2272
rect 1526 2276 1532 2277
rect 1526 2272 1527 2276
rect 1531 2272 1532 2276
rect 1526 2271 1532 2272
rect 1622 2276 1628 2277
rect 1622 2272 1623 2276
rect 1627 2272 1628 2276
rect 1622 2271 1628 2272
rect 1718 2276 1724 2277
rect 1718 2272 1719 2276
rect 1723 2272 1724 2276
rect 1718 2271 1724 2272
rect 1814 2276 1820 2277
rect 1814 2272 1815 2276
rect 1819 2272 1820 2276
rect 1824 2272 1826 2306
rect 1832 2298 1834 2317
rect 1928 2298 1930 2317
rect 2016 2298 2018 2317
rect 2112 2298 2114 2317
rect 2118 2315 2119 2319
rect 2123 2315 2124 2319
rect 2207 2317 2211 2318
rect 2503 2322 2507 2323
rect 2503 2317 2507 2318
rect 2118 2314 2124 2315
rect 2208 2298 2210 2317
rect 1830 2297 1836 2298
rect 1830 2293 1831 2297
rect 1835 2293 1836 2297
rect 1830 2292 1836 2293
rect 1926 2297 1932 2298
rect 1926 2293 1927 2297
rect 1931 2293 1932 2297
rect 1926 2292 1932 2293
rect 2014 2297 2020 2298
rect 2014 2293 2015 2297
rect 2019 2293 2020 2297
rect 2014 2292 2020 2293
rect 2110 2297 2116 2298
rect 2110 2293 2111 2297
rect 2115 2293 2116 2297
rect 2110 2292 2116 2293
rect 2206 2297 2212 2298
rect 2504 2297 2506 2317
rect 2206 2293 2207 2297
rect 2211 2293 2212 2297
rect 2502 2296 2508 2297
rect 2206 2292 2212 2293
rect 2222 2295 2228 2296
rect 2222 2291 2223 2295
rect 2227 2291 2228 2295
rect 2502 2292 2503 2296
rect 2507 2292 2508 2296
rect 2502 2291 2508 2292
rect 2222 2290 2228 2291
rect 1910 2276 1916 2277
rect 1910 2272 1911 2276
rect 1915 2272 1916 2276
rect 1814 2271 1820 2272
rect 1822 2271 1828 2272
rect 1874 2271 1880 2272
rect 1910 2271 1916 2272
rect 1998 2276 2004 2277
rect 1998 2272 1999 2276
rect 2003 2272 2004 2276
rect 1998 2271 2004 2272
rect 2094 2276 2100 2277
rect 2094 2272 2095 2276
rect 2099 2272 2100 2276
rect 2094 2271 2100 2272
rect 2190 2276 2196 2277
rect 2190 2272 2191 2276
rect 2195 2272 2196 2276
rect 2190 2271 2196 2272
rect 1327 2270 1331 2271
rect 1327 2265 1331 2266
rect 1351 2270 1355 2271
rect 1351 2265 1355 2266
rect 1439 2270 1443 2271
rect 1439 2265 1443 2266
rect 1455 2270 1459 2271
rect 1455 2265 1459 2266
rect 1527 2270 1531 2271
rect 1527 2265 1531 2266
rect 1543 2270 1547 2271
rect 1543 2265 1547 2266
rect 1623 2270 1627 2271
rect 1623 2265 1627 2266
rect 1639 2270 1643 2271
rect 1639 2265 1643 2266
rect 1719 2270 1723 2271
rect 1719 2265 1723 2266
rect 1735 2270 1739 2271
rect 1735 2265 1739 2266
rect 1815 2270 1819 2271
rect 1822 2267 1823 2271
rect 1827 2267 1828 2271
rect 1822 2266 1828 2267
rect 1839 2270 1843 2271
rect 1874 2267 1875 2271
rect 1879 2267 1880 2271
rect 1874 2266 1880 2267
rect 1911 2270 1915 2271
rect 1815 2265 1819 2266
rect 1839 2265 1843 2266
rect 1328 2262 1330 2265
rect 1454 2264 1460 2265
rect 1326 2261 1332 2262
rect 983 2258 987 2259
rect 983 2253 987 2254
rect 1007 2258 1011 2259
rect 1007 2253 1011 2254
rect 1047 2258 1051 2259
rect 1047 2253 1051 2254
rect 1095 2258 1099 2259
rect 1102 2258 1108 2259
rect 1111 2258 1115 2259
rect 1095 2253 1099 2254
rect 1287 2258 1291 2259
rect 1111 2253 1115 2254
rect 1130 2255 1136 2256
rect 974 2247 980 2248
rect 974 2243 975 2247
rect 979 2243 980 2247
rect 974 2242 980 2243
rect 984 2234 986 2253
rect 1048 2234 1050 2253
rect 1112 2234 1114 2253
rect 1130 2251 1131 2255
rect 1135 2251 1136 2255
rect 1326 2257 1327 2261
rect 1331 2257 1332 2261
rect 1454 2260 1455 2264
rect 1459 2260 1460 2264
rect 1454 2259 1460 2260
rect 1542 2264 1548 2265
rect 1542 2260 1543 2264
rect 1547 2260 1548 2264
rect 1542 2259 1548 2260
rect 1638 2264 1644 2265
rect 1638 2260 1639 2264
rect 1643 2260 1644 2264
rect 1638 2259 1644 2260
rect 1734 2264 1740 2265
rect 1734 2260 1735 2264
rect 1739 2260 1740 2264
rect 1734 2259 1740 2260
rect 1838 2264 1844 2265
rect 1838 2260 1839 2264
rect 1843 2260 1844 2264
rect 1838 2259 1844 2260
rect 1326 2256 1332 2257
rect 1287 2253 1291 2254
rect 1130 2250 1136 2251
rect 614 2233 620 2234
rect 558 2228 564 2229
rect 582 2231 588 2232
rect 510 2226 516 2227
rect 582 2227 583 2231
rect 587 2227 588 2231
rect 614 2229 615 2233
rect 619 2229 620 2233
rect 614 2228 620 2229
rect 670 2233 676 2234
rect 670 2229 671 2233
rect 675 2229 676 2233
rect 670 2228 676 2229
rect 726 2233 732 2234
rect 726 2229 727 2233
rect 731 2229 732 2233
rect 726 2228 732 2229
rect 790 2233 796 2234
rect 790 2229 791 2233
rect 795 2229 796 2233
rect 790 2228 796 2229
rect 854 2233 860 2234
rect 854 2229 855 2233
rect 859 2229 860 2233
rect 854 2228 860 2229
rect 918 2233 924 2234
rect 918 2229 919 2233
rect 923 2229 924 2233
rect 918 2228 924 2229
rect 982 2233 988 2234
rect 982 2229 983 2233
rect 987 2229 988 2233
rect 982 2228 988 2229
rect 1046 2233 1052 2234
rect 1046 2229 1047 2233
rect 1051 2229 1052 2233
rect 1046 2228 1052 2229
rect 1110 2233 1116 2234
rect 1110 2229 1111 2233
rect 1115 2229 1116 2233
rect 1132 2232 1134 2250
rect 1288 2233 1290 2253
rect 1326 2244 1332 2245
rect 1876 2244 1878 2266
rect 1911 2265 1915 2266
rect 1935 2270 1939 2271
rect 1935 2265 1939 2266
rect 1999 2270 2003 2271
rect 1999 2265 2003 2266
rect 2031 2270 2035 2271
rect 2031 2265 2035 2266
rect 2095 2270 2099 2271
rect 2095 2265 2099 2266
rect 2119 2270 2123 2271
rect 2119 2265 2123 2266
rect 2191 2270 2195 2271
rect 2191 2265 2195 2266
rect 2215 2270 2219 2271
rect 2215 2265 2219 2266
rect 1934 2264 1940 2265
rect 1934 2260 1935 2264
rect 1939 2260 1940 2264
rect 1934 2259 1940 2260
rect 2030 2264 2036 2265
rect 2030 2260 2031 2264
rect 2035 2260 2036 2264
rect 2030 2259 2036 2260
rect 2118 2264 2124 2265
rect 2118 2260 2119 2264
rect 2123 2260 2124 2264
rect 2118 2259 2124 2260
rect 2214 2264 2220 2265
rect 2214 2260 2215 2264
rect 2219 2260 2220 2264
rect 2214 2259 2220 2260
rect 1326 2240 1327 2244
rect 1331 2240 1332 2244
rect 1326 2239 1332 2240
rect 1470 2243 1476 2244
rect 1470 2239 1471 2243
rect 1475 2239 1476 2243
rect 1286 2232 1292 2233
rect 1110 2228 1116 2229
rect 1130 2231 1136 2232
rect 582 2226 588 2227
rect 1130 2227 1131 2231
rect 1135 2227 1136 2231
rect 1286 2228 1287 2232
rect 1291 2228 1292 2232
rect 1286 2227 1292 2228
rect 1130 2226 1136 2227
rect 110 2215 116 2216
rect 110 2211 111 2215
rect 115 2211 116 2215
rect 110 2210 116 2211
rect 246 2212 252 2213
rect 112 2203 114 2210
rect 246 2208 247 2212
rect 251 2208 252 2212
rect 246 2207 252 2208
rect 302 2212 308 2213
rect 302 2208 303 2212
rect 307 2208 308 2212
rect 302 2207 308 2208
rect 366 2212 372 2213
rect 366 2208 367 2212
rect 371 2208 372 2212
rect 366 2207 372 2208
rect 430 2212 436 2213
rect 430 2208 431 2212
rect 435 2208 436 2212
rect 430 2207 436 2208
rect 486 2212 492 2213
rect 486 2208 487 2212
rect 491 2208 492 2212
rect 486 2207 492 2208
rect 248 2203 250 2207
rect 304 2203 306 2207
rect 358 2203 364 2204
rect 368 2203 370 2207
rect 432 2203 434 2207
rect 488 2203 490 2207
rect 512 2204 514 2226
rect 1286 2215 1292 2216
rect 1328 2215 1330 2239
rect 1470 2238 1476 2239
rect 1558 2243 1564 2244
rect 1558 2239 1559 2243
rect 1563 2239 1564 2243
rect 1558 2238 1564 2239
rect 1654 2243 1660 2244
rect 1654 2239 1655 2243
rect 1659 2239 1660 2243
rect 1654 2238 1660 2239
rect 1750 2243 1756 2244
rect 1750 2239 1751 2243
rect 1755 2239 1756 2243
rect 1750 2238 1756 2239
rect 1854 2243 1860 2244
rect 1854 2239 1855 2243
rect 1859 2239 1860 2243
rect 1854 2238 1860 2239
rect 1874 2243 1880 2244
rect 1874 2239 1875 2243
rect 1879 2239 1880 2243
rect 1874 2238 1880 2239
rect 1950 2243 1956 2244
rect 1950 2239 1951 2243
rect 1955 2239 1956 2243
rect 1950 2238 1956 2239
rect 2046 2243 2052 2244
rect 2046 2239 2047 2243
rect 2051 2239 2052 2243
rect 2046 2238 2052 2239
rect 2134 2243 2140 2244
rect 2134 2239 2135 2243
rect 2139 2239 2140 2243
rect 2134 2238 2140 2239
rect 1472 2215 1474 2238
rect 1560 2215 1562 2238
rect 1586 2223 1592 2224
rect 1586 2219 1587 2223
rect 1591 2219 1592 2223
rect 1586 2218 1592 2219
rect 542 2212 548 2213
rect 542 2208 543 2212
rect 547 2208 548 2212
rect 542 2207 548 2208
rect 598 2212 604 2213
rect 598 2208 599 2212
rect 603 2208 604 2212
rect 598 2207 604 2208
rect 654 2212 660 2213
rect 654 2208 655 2212
rect 659 2208 660 2212
rect 654 2207 660 2208
rect 710 2212 716 2213
rect 710 2208 711 2212
rect 715 2208 716 2212
rect 710 2207 716 2208
rect 774 2212 780 2213
rect 774 2208 775 2212
rect 779 2208 780 2212
rect 774 2207 780 2208
rect 838 2212 844 2213
rect 838 2208 839 2212
rect 843 2208 844 2212
rect 838 2207 844 2208
rect 902 2212 908 2213
rect 902 2208 903 2212
rect 907 2208 908 2212
rect 902 2207 908 2208
rect 966 2212 972 2213
rect 966 2208 967 2212
rect 971 2208 972 2212
rect 966 2207 972 2208
rect 1030 2212 1036 2213
rect 1030 2208 1031 2212
rect 1035 2208 1036 2212
rect 1030 2207 1036 2208
rect 1094 2212 1100 2213
rect 1094 2208 1095 2212
rect 1099 2208 1100 2212
rect 1286 2211 1287 2215
rect 1291 2211 1292 2215
rect 1286 2210 1292 2211
rect 1327 2214 1331 2215
rect 1094 2207 1100 2208
rect 510 2203 516 2204
rect 544 2203 546 2207
rect 600 2203 602 2207
rect 656 2203 658 2207
rect 712 2203 714 2207
rect 776 2203 778 2207
rect 840 2203 842 2207
rect 904 2203 906 2207
rect 968 2203 970 2207
rect 1032 2203 1034 2207
rect 1096 2203 1098 2207
rect 1288 2203 1290 2210
rect 1327 2209 1331 2210
rect 1471 2214 1475 2215
rect 1471 2209 1475 2210
rect 1559 2214 1563 2215
rect 1559 2209 1563 2210
rect 1567 2214 1571 2215
rect 1567 2209 1571 2210
rect 111 2202 115 2203
rect 111 2197 115 2198
rect 247 2202 251 2203
rect 247 2197 251 2198
rect 303 2202 307 2203
rect 303 2197 307 2198
rect 335 2202 339 2203
rect 358 2199 359 2203
rect 363 2199 364 2203
rect 358 2198 364 2199
rect 367 2202 371 2203
rect 335 2197 339 2198
rect 112 2194 114 2197
rect 334 2196 340 2197
rect 110 2193 116 2194
rect 110 2189 111 2193
rect 115 2189 116 2193
rect 334 2192 335 2196
rect 339 2192 340 2196
rect 334 2191 340 2192
rect 110 2188 116 2189
rect 110 2176 116 2177
rect 110 2172 111 2176
rect 115 2172 116 2176
rect 110 2171 116 2172
rect 350 2175 356 2176
rect 350 2171 351 2175
rect 355 2171 356 2175
rect 112 2151 114 2171
rect 350 2170 356 2171
rect 352 2151 354 2170
rect 360 2160 362 2198
rect 367 2197 371 2198
rect 391 2202 395 2203
rect 391 2197 395 2198
rect 431 2202 435 2203
rect 431 2197 435 2198
rect 447 2202 451 2203
rect 447 2197 451 2198
rect 487 2202 491 2203
rect 487 2197 491 2198
rect 503 2202 507 2203
rect 510 2199 511 2203
rect 515 2199 516 2203
rect 510 2198 516 2199
rect 543 2202 547 2203
rect 503 2197 507 2198
rect 543 2197 547 2198
rect 559 2202 563 2203
rect 559 2197 563 2198
rect 599 2202 603 2203
rect 599 2197 603 2198
rect 655 2202 659 2203
rect 655 2197 659 2198
rect 711 2202 715 2203
rect 711 2197 715 2198
rect 775 2202 779 2203
rect 775 2197 779 2198
rect 839 2202 843 2203
rect 839 2197 843 2198
rect 903 2202 907 2203
rect 903 2197 907 2198
rect 967 2202 971 2203
rect 967 2197 971 2198
rect 1031 2202 1035 2203
rect 1031 2197 1035 2198
rect 1095 2202 1099 2203
rect 1095 2197 1099 2198
rect 1287 2202 1291 2203
rect 1287 2197 1291 2198
rect 390 2196 396 2197
rect 390 2192 391 2196
rect 395 2192 396 2196
rect 390 2191 396 2192
rect 446 2196 452 2197
rect 446 2192 447 2196
rect 451 2192 452 2196
rect 446 2191 452 2192
rect 502 2196 508 2197
rect 502 2192 503 2196
rect 507 2192 508 2196
rect 502 2191 508 2192
rect 558 2196 564 2197
rect 558 2192 559 2196
rect 563 2192 564 2196
rect 1288 2194 1290 2197
rect 558 2191 564 2192
rect 1286 2193 1292 2194
rect 1286 2189 1287 2193
rect 1291 2189 1292 2193
rect 1328 2189 1330 2209
rect 1568 2190 1570 2209
rect 1566 2189 1572 2190
rect 1286 2188 1292 2189
rect 1326 2188 1332 2189
rect 1326 2184 1327 2188
rect 1331 2184 1332 2188
rect 1566 2185 1567 2189
rect 1571 2185 1572 2189
rect 1588 2188 1590 2218
rect 1656 2215 1658 2238
rect 1752 2215 1754 2238
rect 1856 2215 1858 2238
rect 1952 2215 1954 2238
rect 2048 2215 2050 2238
rect 2136 2215 2138 2238
rect 2224 2224 2226 2290
rect 2502 2279 2508 2280
rect 2502 2275 2503 2279
rect 2507 2275 2508 2279
rect 2502 2274 2508 2275
rect 2504 2271 2506 2274
rect 2311 2270 2315 2271
rect 2311 2265 2315 2266
rect 2503 2270 2507 2271
rect 2503 2265 2507 2266
rect 2310 2264 2316 2265
rect 2310 2260 2311 2264
rect 2315 2260 2316 2264
rect 2504 2262 2506 2265
rect 2310 2259 2316 2260
rect 2502 2261 2508 2262
rect 2502 2257 2503 2261
rect 2507 2257 2508 2261
rect 2502 2256 2508 2257
rect 2502 2244 2508 2245
rect 2230 2243 2236 2244
rect 2230 2239 2231 2243
rect 2235 2239 2236 2243
rect 2230 2238 2236 2239
rect 2326 2243 2332 2244
rect 2326 2239 2327 2243
rect 2331 2239 2332 2243
rect 2326 2238 2332 2239
rect 2334 2243 2340 2244
rect 2334 2239 2335 2243
rect 2339 2239 2340 2243
rect 2502 2240 2503 2244
rect 2507 2240 2508 2244
rect 2502 2239 2508 2240
rect 2334 2238 2340 2239
rect 2222 2223 2228 2224
rect 2222 2219 2223 2223
rect 2227 2219 2228 2223
rect 2222 2218 2228 2219
rect 2232 2215 2234 2238
rect 2328 2215 2330 2238
rect 1623 2214 1627 2215
rect 1623 2209 1627 2210
rect 1655 2214 1659 2215
rect 1655 2209 1659 2210
rect 1679 2214 1683 2215
rect 1679 2209 1683 2210
rect 1743 2214 1747 2215
rect 1743 2209 1747 2210
rect 1751 2214 1755 2215
rect 1751 2209 1755 2210
rect 1807 2214 1811 2215
rect 1807 2209 1811 2210
rect 1855 2214 1859 2215
rect 1855 2209 1859 2210
rect 1871 2214 1875 2215
rect 1927 2214 1931 2215
rect 1871 2209 1875 2210
rect 1890 2211 1896 2212
rect 1624 2190 1626 2209
rect 1680 2190 1682 2209
rect 1744 2190 1746 2209
rect 1808 2190 1810 2209
rect 1826 2203 1832 2204
rect 1826 2199 1827 2203
rect 1831 2199 1832 2203
rect 1826 2198 1832 2199
rect 1622 2189 1628 2190
rect 1566 2184 1572 2185
rect 1586 2187 1592 2188
rect 1326 2183 1332 2184
rect 1586 2183 1587 2187
rect 1591 2183 1592 2187
rect 1622 2185 1623 2189
rect 1627 2185 1628 2189
rect 1622 2184 1628 2185
rect 1678 2189 1684 2190
rect 1678 2185 1679 2189
rect 1683 2185 1684 2189
rect 1678 2184 1684 2185
rect 1742 2189 1748 2190
rect 1742 2185 1743 2189
rect 1747 2185 1748 2189
rect 1742 2184 1748 2185
rect 1806 2189 1812 2190
rect 1806 2185 1807 2189
rect 1811 2185 1812 2189
rect 1806 2184 1812 2185
rect 1586 2182 1592 2183
rect 1286 2176 1292 2177
rect 406 2175 412 2176
rect 406 2171 407 2175
rect 411 2171 412 2175
rect 406 2170 412 2171
rect 462 2175 468 2176
rect 462 2171 463 2175
rect 467 2171 468 2175
rect 462 2170 468 2171
rect 518 2175 524 2176
rect 518 2171 519 2175
rect 523 2171 524 2175
rect 518 2170 524 2171
rect 574 2175 580 2176
rect 574 2171 575 2175
rect 579 2171 580 2175
rect 574 2170 580 2171
rect 582 2175 588 2176
rect 582 2171 583 2175
rect 587 2171 588 2175
rect 1286 2172 1287 2176
rect 1291 2172 1292 2176
rect 1286 2171 1292 2172
rect 1326 2171 1332 2172
rect 582 2170 588 2171
rect 358 2159 364 2160
rect 358 2155 359 2159
rect 363 2155 364 2159
rect 358 2154 364 2155
rect 408 2151 410 2170
rect 464 2151 466 2170
rect 520 2151 522 2170
rect 576 2151 578 2170
rect 111 2150 115 2151
rect 111 2145 115 2146
rect 351 2150 355 2151
rect 351 2145 355 2146
rect 407 2150 411 2151
rect 407 2145 411 2146
rect 415 2150 419 2151
rect 415 2145 419 2146
rect 463 2150 467 2151
rect 463 2145 467 2146
rect 511 2150 515 2151
rect 511 2145 515 2146
rect 519 2150 523 2151
rect 519 2145 523 2146
rect 575 2150 579 2151
rect 584 2148 586 2170
rect 1288 2151 1290 2171
rect 1326 2167 1327 2171
rect 1331 2167 1332 2171
rect 1326 2166 1332 2167
rect 1550 2168 1556 2169
rect 1328 2151 1330 2166
rect 1550 2164 1551 2168
rect 1555 2164 1556 2168
rect 1550 2163 1556 2164
rect 1606 2168 1612 2169
rect 1606 2164 1607 2168
rect 1611 2164 1612 2168
rect 1606 2163 1612 2164
rect 1662 2168 1668 2169
rect 1662 2164 1663 2168
rect 1667 2164 1668 2168
rect 1662 2163 1668 2164
rect 1726 2168 1732 2169
rect 1726 2164 1727 2168
rect 1731 2164 1732 2168
rect 1726 2163 1732 2164
rect 1790 2168 1796 2169
rect 1790 2164 1791 2168
rect 1795 2164 1796 2168
rect 1790 2163 1796 2164
rect 1552 2151 1554 2163
rect 1608 2151 1610 2163
rect 1664 2151 1666 2163
rect 1728 2151 1730 2163
rect 1792 2151 1794 2163
rect 607 2150 611 2151
rect 575 2145 579 2146
rect 582 2147 588 2148
rect 112 2125 114 2145
rect 416 2126 418 2145
rect 512 2126 514 2145
rect 582 2143 583 2147
rect 587 2143 588 2147
rect 607 2145 611 2146
rect 711 2150 715 2151
rect 711 2145 715 2146
rect 815 2150 819 2151
rect 815 2145 819 2146
rect 927 2150 931 2151
rect 927 2145 931 2146
rect 1039 2150 1043 2151
rect 1151 2150 1155 2151
rect 1039 2145 1043 2146
rect 1126 2147 1132 2148
rect 582 2142 588 2143
rect 608 2126 610 2145
rect 712 2126 714 2145
rect 816 2126 818 2145
rect 928 2126 930 2145
rect 1040 2126 1042 2145
rect 1126 2143 1127 2147
rect 1131 2143 1132 2147
rect 1151 2145 1155 2146
rect 1239 2150 1243 2151
rect 1239 2145 1243 2146
rect 1287 2150 1291 2151
rect 1287 2145 1291 2146
rect 1327 2150 1331 2151
rect 1327 2145 1331 2146
rect 1551 2150 1555 2151
rect 1551 2145 1555 2146
rect 1607 2150 1611 2151
rect 1607 2145 1611 2146
rect 1663 2150 1667 2151
rect 1663 2145 1667 2146
rect 1719 2150 1723 2151
rect 1719 2145 1723 2146
rect 1727 2150 1731 2151
rect 1727 2145 1731 2146
rect 1791 2150 1795 2151
rect 1791 2145 1795 2146
rect 1126 2142 1132 2143
rect 414 2125 420 2126
rect 110 2124 116 2125
rect 110 2120 111 2124
rect 115 2120 116 2124
rect 414 2121 415 2125
rect 419 2121 420 2125
rect 414 2120 420 2121
rect 510 2125 516 2126
rect 510 2121 511 2125
rect 515 2121 516 2125
rect 510 2120 516 2121
rect 606 2125 612 2126
rect 606 2121 607 2125
rect 611 2121 612 2125
rect 606 2120 612 2121
rect 710 2125 716 2126
rect 710 2121 711 2125
rect 715 2121 716 2125
rect 710 2120 716 2121
rect 814 2125 820 2126
rect 814 2121 815 2125
rect 819 2121 820 2125
rect 926 2125 932 2126
rect 814 2120 820 2121
rect 822 2123 828 2124
rect 110 2119 116 2120
rect 822 2119 823 2123
rect 827 2119 828 2123
rect 926 2121 927 2125
rect 931 2121 932 2125
rect 926 2120 932 2121
rect 1038 2125 1044 2126
rect 1038 2121 1039 2125
rect 1043 2121 1044 2125
rect 1038 2120 1044 2121
rect 822 2118 828 2119
rect 110 2107 116 2108
rect 110 2103 111 2107
rect 115 2103 116 2107
rect 110 2102 116 2103
rect 398 2104 404 2105
rect 112 2099 114 2102
rect 398 2100 399 2104
rect 403 2100 404 2104
rect 398 2099 404 2100
rect 494 2104 500 2105
rect 494 2100 495 2104
rect 499 2100 500 2104
rect 494 2099 500 2100
rect 590 2104 596 2105
rect 590 2100 591 2104
rect 595 2100 596 2104
rect 590 2099 596 2100
rect 694 2104 700 2105
rect 694 2100 695 2104
rect 699 2100 700 2104
rect 694 2099 700 2100
rect 798 2104 804 2105
rect 798 2100 799 2104
rect 803 2100 804 2104
rect 798 2099 804 2100
rect 111 2098 115 2099
rect 111 2093 115 2094
rect 375 2098 379 2099
rect 375 2093 379 2094
rect 399 2098 403 2099
rect 399 2093 403 2094
rect 447 2098 451 2099
rect 447 2093 451 2094
rect 495 2098 499 2099
rect 495 2093 499 2094
rect 519 2098 523 2099
rect 519 2093 523 2094
rect 591 2098 595 2099
rect 591 2093 595 2094
rect 599 2098 603 2099
rect 599 2093 603 2094
rect 679 2098 683 2099
rect 679 2093 683 2094
rect 695 2098 699 2099
rect 695 2093 699 2094
rect 759 2098 763 2099
rect 759 2093 763 2094
rect 799 2098 803 2099
rect 799 2093 803 2094
rect 112 2090 114 2093
rect 374 2092 380 2093
rect 110 2089 116 2090
rect 110 2085 111 2089
rect 115 2085 116 2089
rect 374 2088 375 2092
rect 379 2088 380 2092
rect 374 2087 380 2088
rect 446 2092 452 2093
rect 446 2088 447 2092
rect 451 2088 452 2092
rect 446 2087 452 2088
rect 518 2092 524 2093
rect 518 2088 519 2092
rect 523 2088 524 2092
rect 518 2087 524 2088
rect 598 2092 604 2093
rect 598 2088 599 2092
rect 603 2088 604 2092
rect 598 2087 604 2088
rect 678 2092 684 2093
rect 678 2088 679 2092
rect 683 2088 684 2092
rect 678 2087 684 2088
rect 758 2092 764 2093
rect 758 2088 759 2092
rect 763 2088 764 2092
rect 758 2087 764 2088
rect 110 2084 116 2085
rect 110 2072 116 2073
rect 110 2068 111 2072
rect 115 2068 116 2072
rect 110 2067 116 2068
rect 390 2071 396 2072
rect 390 2067 391 2071
rect 395 2067 396 2071
rect 112 2043 114 2067
rect 390 2066 396 2067
rect 454 2071 460 2072
rect 454 2067 455 2071
rect 459 2067 460 2071
rect 454 2066 460 2067
rect 462 2071 468 2072
rect 462 2067 463 2071
rect 467 2067 468 2071
rect 462 2066 468 2067
rect 478 2071 484 2072
rect 478 2067 479 2071
rect 483 2067 484 2071
rect 478 2066 484 2067
rect 534 2071 540 2072
rect 534 2067 535 2071
rect 539 2067 540 2071
rect 534 2066 540 2067
rect 614 2071 620 2072
rect 614 2067 615 2071
rect 619 2067 620 2071
rect 614 2066 620 2067
rect 630 2071 636 2072
rect 630 2067 631 2071
rect 635 2067 636 2071
rect 630 2066 636 2067
rect 694 2071 700 2072
rect 694 2067 695 2071
rect 699 2067 700 2071
rect 694 2066 700 2067
rect 774 2071 780 2072
rect 774 2067 775 2071
rect 779 2067 780 2071
rect 774 2066 780 2067
rect 392 2043 394 2066
rect 111 2042 115 2043
rect 111 2037 115 2038
rect 295 2042 299 2043
rect 295 2037 299 2038
rect 375 2042 379 2043
rect 375 2037 379 2038
rect 391 2042 395 2043
rect 391 2037 395 2038
rect 112 2017 114 2037
rect 296 2018 298 2037
rect 376 2018 378 2037
rect 456 2032 458 2066
rect 464 2043 466 2066
rect 480 2052 482 2066
rect 478 2051 484 2052
rect 478 2047 479 2051
rect 483 2047 484 2051
rect 478 2046 484 2047
rect 536 2043 538 2066
rect 616 2043 618 2066
rect 632 2052 634 2066
rect 630 2051 636 2052
rect 630 2047 631 2051
rect 635 2047 636 2051
rect 630 2046 636 2047
rect 696 2043 698 2066
rect 776 2043 778 2066
rect 824 2064 826 2118
rect 910 2104 916 2105
rect 910 2100 911 2104
rect 915 2100 916 2104
rect 910 2099 916 2100
rect 1022 2104 1028 2105
rect 1022 2100 1023 2104
rect 1027 2100 1028 2104
rect 1022 2099 1028 2100
rect 831 2098 835 2099
rect 831 2093 835 2094
rect 903 2098 907 2099
rect 903 2093 907 2094
rect 911 2098 915 2099
rect 911 2093 915 2094
rect 967 2098 971 2099
rect 967 2093 971 2094
rect 1023 2098 1027 2099
rect 1023 2093 1027 2094
rect 1031 2098 1035 2099
rect 1031 2093 1035 2094
rect 1103 2098 1107 2099
rect 1103 2093 1107 2094
rect 830 2092 836 2093
rect 830 2088 831 2092
rect 835 2088 836 2092
rect 830 2087 836 2088
rect 902 2092 908 2093
rect 902 2088 903 2092
rect 907 2088 908 2092
rect 902 2087 908 2088
rect 966 2092 972 2093
rect 966 2088 967 2092
rect 971 2088 972 2092
rect 966 2087 972 2088
rect 1030 2092 1036 2093
rect 1030 2088 1031 2092
rect 1035 2088 1036 2092
rect 1030 2087 1036 2088
rect 1102 2092 1108 2093
rect 1102 2088 1103 2092
rect 1107 2088 1108 2092
rect 1102 2087 1108 2088
rect 1128 2072 1130 2142
rect 1152 2126 1154 2145
rect 1240 2126 1242 2145
rect 1150 2125 1156 2126
rect 1150 2121 1151 2125
rect 1155 2121 1156 2125
rect 1150 2120 1156 2121
rect 1238 2125 1244 2126
rect 1288 2125 1290 2145
rect 1328 2142 1330 2145
rect 1662 2144 1668 2145
rect 1326 2141 1332 2142
rect 1326 2137 1327 2141
rect 1331 2137 1332 2141
rect 1662 2140 1663 2144
rect 1667 2140 1668 2144
rect 1662 2139 1668 2140
rect 1718 2144 1724 2145
rect 1718 2140 1719 2144
rect 1723 2140 1724 2144
rect 1718 2139 1724 2140
rect 1790 2144 1796 2145
rect 1790 2140 1791 2144
rect 1795 2140 1796 2144
rect 1790 2139 1796 2140
rect 1326 2136 1332 2137
rect 1238 2121 1239 2125
rect 1243 2121 1244 2125
rect 1286 2124 1292 2125
rect 1238 2120 1244 2121
rect 1254 2123 1260 2124
rect 1254 2119 1255 2123
rect 1259 2119 1260 2123
rect 1286 2120 1287 2124
rect 1291 2120 1292 2124
rect 1286 2119 1292 2120
rect 1326 2124 1332 2125
rect 1828 2124 1830 2198
rect 1872 2190 1874 2209
rect 1890 2207 1891 2211
rect 1895 2207 1896 2211
rect 1927 2209 1931 2210
rect 1951 2214 1955 2215
rect 1951 2209 1955 2210
rect 1983 2214 1987 2215
rect 1983 2209 1987 2210
rect 2039 2214 2043 2215
rect 2039 2209 2043 2210
rect 2047 2214 2051 2215
rect 2047 2209 2051 2210
rect 2095 2214 2099 2215
rect 2095 2209 2099 2210
rect 2135 2214 2139 2215
rect 2135 2209 2139 2210
rect 2159 2214 2163 2215
rect 2159 2209 2163 2210
rect 2223 2214 2227 2215
rect 2223 2209 2227 2210
rect 2231 2214 2235 2215
rect 2231 2209 2235 2210
rect 2287 2214 2291 2215
rect 2287 2209 2291 2210
rect 2327 2214 2331 2215
rect 2336 2212 2338 2238
rect 2504 2215 2506 2239
rect 2343 2214 2347 2215
rect 2327 2209 2331 2210
rect 2334 2211 2340 2212
rect 1890 2206 1896 2207
rect 1870 2189 1876 2190
rect 1870 2185 1871 2189
rect 1875 2185 1876 2189
rect 1892 2188 1894 2206
rect 1928 2190 1930 2209
rect 1984 2190 1986 2209
rect 2040 2190 2042 2209
rect 2096 2190 2098 2209
rect 2160 2190 2162 2209
rect 2224 2190 2226 2209
rect 2288 2190 2290 2209
rect 2334 2207 2335 2211
rect 2339 2207 2340 2211
rect 2343 2209 2347 2210
rect 2399 2214 2403 2215
rect 2399 2209 2403 2210
rect 2455 2214 2459 2215
rect 2455 2209 2459 2210
rect 2503 2214 2507 2215
rect 2503 2209 2507 2210
rect 2334 2206 2340 2207
rect 2344 2190 2346 2209
rect 2400 2190 2402 2209
rect 2456 2190 2458 2209
rect 1926 2189 1932 2190
rect 1870 2184 1876 2185
rect 1890 2187 1896 2188
rect 1890 2183 1891 2187
rect 1895 2183 1896 2187
rect 1926 2185 1927 2189
rect 1931 2185 1932 2189
rect 1926 2184 1932 2185
rect 1982 2189 1988 2190
rect 1982 2185 1983 2189
rect 1987 2185 1988 2189
rect 1982 2184 1988 2185
rect 2038 2189 2044 2190
rect 2038 2185 2039 2189
rect 2043 2185 2044 2189
rect 2038 2184 2044 2185
rect 2094 2189 2100 2190
rect 2094 2185 2095 2189
rect 2099 2185 2100 2189
rect 2094 2184 2100 2185
rect 2158 2189 2164 2190
rect 2158 2185 2159 2189
rect 2163 2185 2164 2189
rect 2158 2184 2164 2185
rect 2222 2189 2228 2190
rect 2222 2185 2223 2189
rect 2227 2185 2228 2189
rect 2222 2184 2228 2185
rect 2286 2189 2292 2190
rect 2286 2185 2287 2189
rect 2291 2185 2292 2189
rect 2286 2184 2292 2185
rect 2342 2189 2348 2190
rect 2342 2185 2343 2189
rect 2347 2185 2348 2189
rect 2342 2184 2348 2185
rect 2398 2189 2404 2190
rect 2398 2185 2399 2189
rect 2403 2185 2404 2189
rect 2398 2184 2404 2185
rect 2454 2189 2460 2190
rect 2504 2189 2506 2209
rect 2454 2185 2455 2189
rect 2459 2185 2460 2189
rect 2502 2188 2508 2189
rect 2454 2184 2460 2185
rect 2470 2187 2476 2188
rect 1890 2182 1896 2183
rect 2470 2183 2471 2187
rect 2475 2183 2476 2187
rect 2502 2184 2503 2188
rect 2507 2184 2508 2188
rect 2502 2183 2508 2184
rect 2470 2182 2476 2183
rect 1854 2168 1860 2169
rect 1854 2164 1855 2168
rect 1859 2164 1860 2168
rect 1854 2163 1860 2164
rect 1910 2168 1916 2169
rect 1910 2164 1911 2168
rect 1915 2164 1916 2168
rect 1910 2163 1916 2164
rect 1966 2168 1972 2169
rect 1966 2164 1967 2168
rect 1971 2164 1972 2168
rect 1966 2163 1972 2164
rect 2022 2168 2028 2169
rect 2022 2164 2023 2168
rect 2027 2164 2028 2168
rect 2022 2163 2028 2164
rect 2078 2168 2084 2169
rect 2078 2164 2079 2168
rect 2083 2164 2084 2168
rect 2078 2163 2084 2164
rect 2142 2168 2148 2169
rect 2142 2164 2143 2168
rect 2147 2164 2148 2168
rect 2142 2163 2148 2164
rect 2206 2168 2212 2169
rect 2206 2164 2207 2168
rect 2211 2164 2212 2168
rect 2206 2163 2212 2164
rect 2270 2168 2276 2169
rect 2270 2164 2271 2168
rect 2275 2164 2276 2168
rect 2270 2163 2276 2164
rect 2326 2168 2332 2169
rect 2326 2164 2327 2168
rect 2331 2164 2332 2168
rect 2326 2163 2332 2164
rect 2382 2168 2388 2169
rect 2382 2164 2383 2168
rect 2387 2164 2388 2168
rect 2382 2163 2388 2164
rect 2438 2168 2444 2169
rect 2438 2164 2439 2168
rect 2443 2164 2444 2168
rect 2438 2163 2444 2164
rect 1856 2151 1858 2163
rect 1912 2151 1914 2163
rect 1968 2151 1970 2163
rect 2024 2151 2026 2163
rect 2080 2151 2082 2163
rect 2144 2151 2146 2163
rect 2208 2151 2210 2163
rect 2272 2151 2274 2163
rect 2328 2151 2330 2163
rect 2384 2151 2386 2163
rect 2440 2151 2442 2163
rect 1855 2150 1859 2151
rect 1855 2145 1859 2146
rect 1871 2150 1875 2151
rect 1871 2145 1875 2146
rect 1911 2150 1915 2151
rect 1911 2145 1915 2146
rect 1967 2150 1971 2151
rect 1967 2145 1971 2146
rect 2023 2150 2027 2151
rect 2023 2145 2027 2146
rect 2079 2150 2083 2151
rect 2079 2145 2083 2146
rect 2143 2150 2147 2151
rect 2143 2145 2147 2146
rect 2199 2150 2203 2151
rect 2199 2145 2203 2146
rect 2207 2150 2211 2151
rect 2207 2145 2211 2146
rect 2271 2150 2275 2151
rect 2271 2145 2275 2146
rect 2327 2150 2331 2151
rect 2327 2145 2331 2146
rect 2383 2150 2387 2151
rect 2383 2145 2387 2146
rect 2439 2150 2443 2151
rect 2439 2145 2443 2146
rect 1870 2144 1876 2145
rect 1870 2140 1871 2144
rect 1875 2140 1876 2144
rect 1870 2139 1876 2140
rect 1966 2144 1972 2145
rect 1966 2140 1967 2144
rect 1971 2140 1972 2144
rect 1966 2139 1972 2140
rect 2078 2144 2084 2145
rect 2078 2140 2079 2144
rect 2083 2140 2084 2144
rect 2078 2139 2084 2140
rect 2198 2144 2204 2145
rect 2198 2140 2199 2144
rect 2203 2140 2204 2144
rect 2198 2139 2204 2140
rect 2326 2144 2332 2145
rect 2326 2140 2327 2144
rect 2331 2140 2332 2144
rect 2326 2139 2332 2140
rect 2438 2144 2444 2145
rect 2438 2140 2439 2144
rect 2443 2140 2444 2144
rect 2438 2139 2444 2140
rect 1326 2120 1327 2124
rect 1331 2120 1332 2124
rect 1326 2119 1332 2120
rect 1678 2123 1684 2124
rect 1678 2119 1679 2123
rect 1683 2119 1684 2123
rect 1254 2118 1260 2119
rect 1134 2104 1140 2105
rect 1134 2100 1135 2104
rect 1139 2100 1140 2104
rect 1134 2099 1140 2100
rect 1222 2104 1228 2105
rect 1222 2100 1223 2104
rect 1227 2100 1228 2104
rect 1222 2099 1228 2100
rect 1135 2098 1139 2099
rect 1135 2093 1139 2094
rect 1167 2098 1171 2099
rect 1167 2093 1171 2094
rect 1223 2098 1227 2099
rect 1223 2093 1227 2094
rect 1166 2092 1172 2093
rect 1166 2088 1167 2092
rect 1171 2088 1172 2092
rect 1166 2087 1172 2088
rect 1222 2092 1228 2093
rect 1222 2088 1223 2092
rect 1227 2088 1228 2092
rect 1222 2087 1228 2088
rect 846 2071 852 2072
rect 846 2067 847 2071
rect 851 2067 852 2071
rect 846 2066 852 2067
rect 918 2071 924 2072
rect 918 2067 919 2071
rect 923 2067 924 2071
rect 918 2066 924 2067
rect 982 2071 988 2072
rect 982 2067 983 2071
rect 987 2067 988 2071
rect 982 2066 988 2067
rect 1046 2071 1052 2072
rect 1046 2067 1047 2071
rect 1051 2067 1052 2071
rect 1046 2066 1052 2067
rect 1118 2071 1124 2072
rect 1118 2067 1119 2071
rect 1123 2067 1124 2071
rect 1118 2066 1124 2067
rect 1126 2071 1132 2072
rect 1126 2067 1127 2071
rect 1131 2067 1132 2071
rect 1126 2066 1132 2067
rect 1182 2071 1188 2072
rect 1182 2067 1183 2071
rect 1187 2067 1188 2071
rect 1182 2066 1188 2067
rect 1238 2071 1244 2072
rect 1238 2067 1239 2071
rect 1243 2067 1244 2071
rect 1238 2066 1244 2067
rect 822 2063 828 2064
rect 822 2059 823 2063
rect 827 2059 828 2063
rect 822 2058 828 2059
rect 848 2043 850 2066
rect 920 2043 922 2066
rect 984 2043 986 2066
rect 1048 2043 1050 2066
rect 1082 2051 1088 2052
rect 1082 2047 1083 2051
rect 1087 2047 1088 2051
rect 1082 2046 1088 2047
rect 463 2042 467 2043
rect 463 2037 467 2038
rect 535 2042 539 2043
rect 535 2037 539 2038
rect 551 2042 555 2043
rect 551 2037 555 2038
rect 615 2042 619 2043
rect 615 2037 619 2038
rect 639 2042 643 2043
rect 695 2042 699 2043
rect 639 2037 643 2038
rect 658 2039 664 2040
rect 454 2031 460 2032
rect 454 2027 455 2031
rect 459 2027 460 2031
rect 454 2026 460 2027
rect 464 2018 466 2037
rect 552 2018 554 2037
rect 640 2018 642 2037
rect 658 2035 659 2039
rect 663 2035 664 2039
rect 695 2037 699 2038
rect 719 2042 723 2043
rect 719 2037 723 2038
rect 775 2042 779 2043
rect 775 2037 779 2038
rect 799 2042 803 2043
rect 799 2037 803 2038
rect 847 2042 851 2043
rect 847 2037 851 2038
rect 887 2042 891 2043
rect 887 2037 891 2038
rect 919 2042 923 2043
rect 919 2037 923 2038
rect 975 2042 979 2043
rect 975 2037 979 2038
rect 983 2042 987 2043
rect 983 2037 987 2038
rect 1047 2042 1051 2043
rect 1047 2037 1051 2038
rect 1063 2042 1067 2043
rect 1063 2037 1067 2038
rect 658 2034 664 2035
rect 294 2017 300 2018
rect 110 2016 116 2017
rect 110 2012 111 2016
rect 115 2012 116 2016
rect 294 2013 295 2017
rect 299 2013 300 2017
rect 294 2012 300 2013
rect 374 2017 380 2018
rect 374 2013 375 2017
rect 379 2013 380 2017
rect 462 2017 468 2018
rect 374 2012 380 2013
rect 406 2015 412 2016
rect 110 2011 116 2012
rect 406 2011 407 2015
rect 411 2011 412 2015
rect 462 2013 463 2017
rect 467 2013 468 2017
rect 462 2012 468 2013
rect 550 2017 556 2018
rect 550 2013 551 2017
rect 555 2013 556 2017
rect 550 2012 556 2013
rect 638 2017 644 2018
rect 638 2013 639 2017
rect 643 2013 644 2017
rect 660 2016 662 2034
rect 720 2018 722 2037
rect 726 2031 732 2032
rect 726 2027 727 2031
rect 731 2027 732 2031
rect 726 2026 732 2027
rect 718 2017 724 2018
rect 638 2012 644 2013
rect 658 2015 664 2016
rect 406 2010 412 2011
rect 658 2011 659 2015
rect 663 2011 664 2015
rect 718 2013 719 2017
rect 723 2013 724 2017
rect 718 2012 724 2013
rect 658 2010 664 2011
rect 110 1999 116 2000
rect 110 1995 111 1999
rect 115 1995 116 1999
rect 110 1994 116 1995
rect 278 1996 284 1997
rect 112 1987 114 1994
rect 278 1992 279 1996
rect 283 1992 284 1996
rect 278 1991 284 1992
rect 358 1996 364 1997
rect 358 1992 359 1996
rect 363 1992 364 1996
rect 358 1991 364 1992
rect 280 1987 282 1991
rect 360 1987 362 1991
rect 111 1986 115 1987
rect 111 1981 115 1982
rect 135 1986 139 1987
rect 135 1981 139 1982
rect 207 1986 211 1987
rect 207 1981 211 1982
rect 279 1986 283 1987
rect 279 1981 283 1982
rect 287 1986 291 1987
rect 287 1981 291 1982
rect 359 1986 363 1987
rect 359 1981 363 1982
rect 383 1986 387 1987
rect 383 1981 387 1982
rect 112 1978 114 1981
rect 134 1980 140 1981
rect 110 1977 116 1978
rect 110 1973 111 1977
rect 115 1973 116 1977
rect 134 1976 135 1980
rect 139 1976 140 1980
rect 134 1975 140 1976
rect 206 1980 212 1981
rect 206 1976 207 1980
rect 211 1976 212 1980
rect 206 1975 212 1976
rect 286 1980 292 1981
rect 286 1976 287 1980
rect 291 1976 292 1980
rect 286 1975 292 1976
rect 382 1980 388 1981
rect 382 1976 383 1980
rect 387 1976 388 1980
rect 382 1975 388 1976
rect 110 1972 116 1973
rect 110 1960 116 1961
rect 110 1956 111 1960
rect 115 1956 116 1960
rect 110 1955 116 1956
rect 150 1959 156 1960
rect 150 1955 151 1959
rect 155 1955 156 1959
rect 112 1927 114 1955
rect 150 1954 156 1955
rect 222 1959 228 1960
rect 222 1955 223 1959
rect 227 1955 228 1959
rect 222 1954 228 1955
rect 302 1959 308 1960
rect 302 1955 303 1959
rect 307 1955 308 1959
rect 302 1954 308 1955
rect 366 1959 372 1960
rect 366 1955 367 1959
rect 371 1955 372 1959
rect 366 1954 372 1955
rect 398 1959 404 1960
rect 398 1955 399 1959
rect 403 1955 404 1959
rect 398 1954 404 1955
rect 152 1927 154 1954
rect 224 1927 226 1954
rect 304 1927 306 1954
rect 111 1926 115 1927
rect 111 1921 115 1922
rect 151 1926 155 1927
rect 151 1921 155 1922
rect 223 1926 227 1927
rect 223 1921 227 1922
rect 239 1926 243 1927
rect 239 1921 243 1922
rect 303 1926 307 1927
rect 303 1921 307 1922
rect 112 1901 114 1921
rect 152 1902 154 1921
rect 240 1902 242 1921
rect 368 1916 370 1954
rect 400 1927 402 1954
rect 408 1944 410 2010
rect 446 1996 452 1997
rect 446 1992 447 1996
rect 451 1992 452 1996
rect 446 1991 452 1992
rect 534 1996 540 1997
rect 534 1992 535 1996
rect 539 1992 540 1996
rect 534 1991 540 1992
rect 622 1996 628 1997
rect 622 1992 623 1996
rect 627 1992 628 1996
rect 622 1991 628 1992
rect 702 1996 708 1997
rect 702 1992 703 1996
rect 707 1992 708 1996
rect 702 1991 708 1992
rect 448 1987 450 1991
rect 536 1987 538 1991
rect 624 1987 626 1991
rect 704 1987 706 1991
rect 447 1986 451 1987
rect 447 1981 451 1982
rect 487 1986 491 1987
rect 487 1981 491 1982
rect 535 1986 539 1987
rect 535 1981 539 1982
rect 591 1986 595 1987
rect 591 1981 595 1982
rect 623 1986 627 1987
rect 623 1981 627 1982
rect 695 1986 699 1987
rect 695 1981 699 1982
rect 703 1986 707 1987
rect 703 1981 707 1982
rect 486 1980 492 1981
rect 486 1976 487 1980
rect 491 1976 492 1980
rect 486 1975 492 1976
rect 590 1980 596 1981
rect 590 1976 591 1980
rect 595 1976 596 1980
rect 590 1975 596 1976
rect 694 1980 700 1981
rect 694 1976 695 1980
rect 699 1976 700 1980
rect 694 1975 700 1976
rect 728 1960 730 2026
rect 800 2018 802 2037
rect 888 2018 890 2037
rect 976 2018 978 2037
rect 1064 2018 1066 2037
rect 798 2017 804 2018
rect 798 2013 799 2017
rect 803 2013 804 2017
rect 798 2012 804 2013
rect 886 2017 892 2018
rect 886 2013 887 2017
rect 891 2013 892 2017
rect 886 2012 892 2013
rect 974 2017 980 2018
rect 974 2013 975 2017
rect 979 2013 980 2017
rect 974 2012 980 2013
rect 1062 2017 1068 2018
rect 1062 2013 1063 2017
rect 1067 2013 1068 2017
rect 1084 2016 1086 2046
rect 1120 2043 1122 2066
rect 1184 2043 1186 2066
rect 1240 2043 1242 2066
rect 1256 2052 1258 2118
rect 1286 2107 1292 2108
rect 1286 2103 1287 2107
rect 1291 2103 1292 2107
rect 1286 2102 1292 2103
rect 1288 2099 1290 2102
rect 1287 2098 1291 2099
rect 1287 2093 1291 2094
rect 1288 2090 1290 2093
rect 1286 2089 1292 2090
rect 1286 2085 1287 2089
rect 1291 2085 1292 2089
rect 1328 2087 1330 2119
rect 1678 2118 1684 2119
rect 1734 2123 1740 2124
rect 1734 2119 1735 2123
rect 1739 2119 1740 2123
rect 1734 2118 1740 2119
rect 1806 2123 1812 2124
rect 1806 2119 1807 2123
rect 1811 2119 1812 2123
rect 1806 2118 1812 2119
rect 1826 2123 1832 2124
rect 1826 2119 1827 2123
rect 1831 2119 1832 2123
rect 1826 2118 1832 2119
rect 1886 2123 1892 2124
rect 1886 2119 1887 2123
rect 1891 2119 1892 2123
rect 1886 2118 1892 2119
rect 1982 2123 1988 2124
rect 1982 2119 1983 2123
rect 1987 2119 1988 2123
rect 1982 2118 1988 2119
rect 1990 2123 1996 2124
rect 1990 2119 1991 2123
rect 1995 2119 1996 2123
rect 1990 2118 1996 2119
rect 2094 2123 2100 2124
rect 2094 2119 2095 2123
rect 2099 2119 2100 2123
rect 2094 2118 2100 2119
rect 2214 2123 2220 2124
rect 2214 2119 2215 2123
rect 2219 2119 2220 2123
rect 2214 2118 2220 2119
rect 2342 2123 2348 2124
rect 2342 2119 2343 2123
rect 2347 2119 2348 2123
rect 2342 2118 2348 2119
rect 2454 2123 2460 2124
rect 2454 2119 2455 2123
rect 2459 2119 2460 2123
rect 2454 2118 2460 2119
rect 2462 2123 2468 2124
rect 2462 2119 2463 2123
rect 2467 2119 2468 2123
rect 2462 2118 2468 2119
rect 1680 2087 1682 2118
rect 1736 2087 1738 2118
rect 1808 2087 1810 2118
rect 1888 2087 1890 2118
rect 1984 2087 1986 2118
rect 1992 2100 1994 2118
rect 1990 2099 1996 2100
rect 1990 2095 1991 2099
rect 1995 2095 1996 2099
rect 1990 2094 1996 2095
rect 2096 2087 2098 2118
rect 2216 2087 2218 2118
rect 2334 2107 2340 2108
rect 2334 2103 2335 2107
rect 2339 2103 2340 2107
rect 2334 2102 2340 2103
rect 1286 2084 1292 2085
rect 1327 2086 1331 2087
rect 1327 2081 1331 2082
rect 1367 2086 1371 2087
rect 1367 2081 1371 2082
rect 1423 2086 1427 2087
rect 1423 2081 1427 2082
rect 1503 2086 1507 2087
rect 1503 2081 1507 2082
rect 1591 2086 1595 2087
rect 1591 2081 1595 2082
rect 1679 2086 1683 2087
rect 1679 2081 1683 2082
rect 1735 2086 1739 2087
rect 1735 2081 1739 2082
rect 1783 2086 1787 2087
rect 1783 2081 1787 2082
rect 1807 2086 1811 2087
rect 1887 2086 1891 2087
rect 1807 2081 1811 2082
rect 1858 2083 1864 2084
rect 1286 2072 1292 2073
rect 1286 2068 1287 2072
rect 1291 2068 1292 2072
rect 1286 2067 1292 2068
rect 1254 2051 1260 2052
rect 1254 2047 1255 2051
rect 1259 2047 1260 2051
rect 1254 2046 1260 2047
rect 1288 2043 1290 2067
rect 1328 2061 1330 2081
rect 1368 2062 1370 2081
rect 1424 2062 1426 2081
rect 1504 2062 1506 2081
rect 1592 2062 1594 2081
rect 1680 2062 1682 2081
rect 1784 2062 1786 2081
rect 1858 2079 1859 2083
rect 1863 2079 1864 2083
rect 1887 2081 1891 2082
rect 1895 2086 1899 2087
rect 1895 2081 1899 2082
rect 1983 2086 1987 2087
rect 1983 2081 1987 2082
rect 2023 2086 2027 2087
rect 2023 2081 2027 2082
rect 2095 2086 2099 2087
rect 2095 2081 2099 2082
rect 2167 2086 2171 2087
rect 2167 2081 2171 2082
rect 2215 2086 2219 2087
rect 2215 2081 2219 2082
rect 2319 2086 2323 2087
rect 2319 2081 2323 2082
rect 1858 2078 1864 2079
rect 1366 2061 1372 2062
rect 1326 2060 1332 2061
rect 1326 2056 1327 2060
rect 1331 2056 1332 2060
rect 1366 2057 1367 2061
rect 1371 2057 1372 2061
rect 1366 2056 1372 2057
rect 1422 2061 1428 2062
rect 1422 2057 1423 2061
rect 1427 2057 1428 2061
rect 1422 2056 1428 2057
rect 1502 2061 1508 2062
rect 1502 2057 1503 2061
rect 1507 2057 1508 2061
rect 1502 2056 1508 2057
rect 1590 2061 1596 2062
rect 1590 2057 1591 2061
rect 1595 2057 1596 2061
rect 1590 2056 1596 2057
rect 1678 2061 1684 2062
rect 1678 2057 1679 2061
rect 1683 2057 1684 2061
rect 1782 2061 1788 2062
rect 1678 2056 1684 2057
rect 1686 2059 1692 2060
rect 1326 2055 1332 2056
rect 1686 2055 1687 2059
rect 1691 2055 1692 2059
rect 1782 2057 1783 2061
rect 1787 2057 1788 2061
rect 1782 2056 1788 2057
rect 1686 2054 1692 2055
rect 1326 2043 1332 2044
rect 1119 2042 1123 2043
rect 1119 2037 1123 2038
rect 1183 2042 1187 2043
rect 1183 2037 1187 2038
rect 1239 2042 1243 2043
rect 1239 2037 1243 2038
rect 1287 2042 1291 2043
rect 1326 2039 1327 2043
rect 1331 2039 1332 2043
rect 1326 2038 1332 2039
rect 1350 2040 1356 2041
rect 1287 2037 1291 2038
rect 1288 2017 1290 2037
rect 1328 2035 1330 2038
rect 1350 2036 1351 2040
rect 1355 2036 1356 2040
rect 1350 2035 1356 2036
rect 1406 2040 1412 2041
rect 1406 2036 1407 2040
rect 1411 2036 1412 2040
rect 1406 2035 1412 2036
rect 1486 2040 1492 2041
rect 1486 2036 1487 2040
rect 1491 2036 1492 2040
rect 1486 2035 1492 2036
rect 1574 2040 1580 2041
rect 1574 2036 1575 2040
rect 1579 2036 1580 2040
rect 1574 2035 1580 2036
rect 1662 2040 1668 2041
rect 1662 2036 1663 2040
rect 1667 2036 1668 2040
rect 1662 2035 1668 2036
rect 1327 2034 1331 2035
rect 1327 2029 1331 2030
rect 1351 2034 1355 2035
rect 1351 2029 1355 2030
rect 1407 2034 1411 2035
rect 1407 2029 1411 2030
rect 1423 2034 1427 2035
rect 1423 2029 1427 2030
rect 1487 2034 1491 2035
rect 1487 2029 1491 2030
rect 1519 2034 1523 2035
rect 1519 2029 1523 2030
rect 1575 2034 1579 2035
rect 1575 2029 1579 2030
rect 1615 2034 1619 2035
rect 1615 2029 1619 2030
rect 1663 2034 1667 2035
rect 1663 2029 1667 2030
rect 1328 2026 1330 2029
rect 1350 2028 1356 2029
rect 1326 2025 1332 2026
rect 1326 2021 1327 2025
rect 1331 2021 1332 2025
rect 1350 2024 1351 2028
rect 1355 2024 1356 2028
rect 1350 2023 1356 2024
rect 1422 2028 1428 2029
rect 1422 2024 1423 2028
rect 1427 2024 1428 2028
rect 1422 2023 1428 2024
rect 1518 2028 1524 2029
rect 1518 2024 1519 2028
rect 1523 2024 1524 2028
rect 1518 2023 1524 2024
rect 1614 2028 1620 2029
rect 1614 2024 1615 2028
rect 1619 2024 1620 2028
rect 1614 2023 1620 2024
rect 1326 2020 1332 2021
rect 1286 2016 1292 2017
rect 1062 2012 1068 2013
rect 1082 2015 1088 2016
rect 1082 2011 1083 2015
rect 1087 2011 1088 2015
rect 1286 2012 1287 2016
rect 1291 2012 1292 2016
rect 1286 2011 1292 2012
rect 1082 2010 1088 2011
rect 1326 2008 1332 2009
rect 1326 2004 1327 2008
rect 1331 2004 1332 2008
rect 1326 2003 1332 2004
rect 1366 2007 1372 2008
rect 1366 2003 1367 2007
rect 1371 2003 1372 2007
rect 1286 1999 1292 2000
rect 782 1996 788 1997
rect 782 1992 783 1996
rect 787 1992 788 1996
rect 782 1991 788 1992
rect 870 1996 876 1997
rect 870 1992 871 1996
rect 875 1992 876 1996
rect 870 1991 876 1992
rect 958 1996 964 1997
rect 958 1992 959 1996
rect 963 1992 964 1996
rect 958 1991 964 1992
rect 1046 1996 1052 1997
rect 1046 1992 1047 1996
rect 1051 1992 1052 1996
rect 1286 1995 1287 1999
rect 1291 1995 1292 1999
rect 1286 1994 1292 1995
rect 1046 1991 1052 1992
rect 784 1987 786 1991
rect 872 1987 874 1991
rect 960 1987 962 1991
rect 1048 1987 1050 1991
rect 1288 1987 1290 1994
rect 783 1986 787 1987
rect 783 1981 787 1982
rect 799 1986 803 1987
rect 799 1981 803 1982
rect 871 1986 875 1987
rect 871 1981 875 1982
rect 903 1986 907 1987
rect 903 1981 907 1982
rect 959 1986 963 1987
rect 959 1981 963 1982
rect 1015 1986 1019 1987
rect 1015 1981 1019 1982
rect 1047 1986 1051 1987
rect 1047 1981 1051 1982
rect 1287 1986 1291 1987
rect 1287 1981 1291 1982
rect 798 1980 804 1981
rect 798 1976 799 1980
rect 803 1976 804 1980
rect 798 1975 804 1976
rect 902 1980 908 1981
rect 902 1976 903 1980
rect 907 1976 908 1980
rect 902 1975 908 1976
rect 1014 1980 1020 1981
rect 1014 1976 1015 1980
rect 1019 1976 1020 1980
rect 1288 1978 1290 1981
rect 1328 1979 1330 2003
rect 1366 2002 1372 2003
rect 1438 2007 1444 2008
rect 1438 2003 1439 2007
rect 1443 2003 1444 2007
rect 1438 2002 1444 2003
rect 1534 2007 1540 2008
rect 1534 2003 1535 2007
rect 1539 2003 1540 2007
rect 1534 2002 1540 2003
rect 1630 2007 1636 2008
rect 1630 2003 1631 2007
rect 1635 2003 1636 2007
rect 1630 2002 1636 2003
rect 1368 1979 1370 2002
rect 1440 1979 1442 2002
rect 1536 1979 1538 2002
rect 1632 1979 1634 2002
rect 1688 1988 1690 2054
rect 1766 2040 1772 2041
rect 1766 2036 1767 2040
rect 1771 2036 1772 2040
rect 1766 2035 1772 2036
rect 1719 2034 1723 2035
rect 1719 2029 1723 2030
rect 1767 2034 1771 2035
rect 1767 2029 1771 2030
rect 1823 2034 1827 2035
rect 1823 2029 1827 2030
rect 1718 2028 1724 2029
rect 1718 2024 1719 2028
rect 1723 2024 1724 2028
rect 1718 2023 1724 2024
rect 1822 2028 1828 2029
rect 1822 2024 1823 2028
rect 1827 2024 1828 2028
rect 1822 2023 1828 2024
rect 1860 2008 1862 2078
rect 1896 2062 1898 2081
rect 2024 2062 2026 2081
rect 2168 2062 2170 2081
rect 2320 2062 2322 2081
rect 1894 2061 1900 2062
rect 1894 2057 1895 2061
rect 1899 2057 1900 2061
rect 1894 2056 1900 2057
rect 2022 2061 2028 2062
rect 2022 2057 2023 2061
rect 2027 2057 2028 2061
rect 2022 2056 2028 2057
rect 2166 2061 2172 2062
rect 2166 2057 2167 2061
rect 2171 2057 2172 2061
rect 2166 2056 2172 2057
rect 2318 2061 2324 2062
rect 2318 2057 2319 2061
rect 2323 2057 2324 2061
rect 2336 2060 2338 2102
rect 2344 2087 2346 2118
rect 2456 2087 2458 2118
rect 2343 2086 2347 2087
rect 2343 2081 2347 2082
rect 2455 2086 2459 2087
rect 2455 2081 2459 2082
rect 2456 2062 2458 2081
rect 2464 2076 2466 2118
rect 2472 2104 2474 2182
rect 2502 2171 2508 2172
rect 2502 2167 2503 2171
rect 2507 2167 2508 2171
rect 2502 2166 2508 2167
rect 2504 2151 2506 2166
rect 2503 2150 2507 2151
rect 2503 2145 2507 2146
rect 2504 2142 2506 2145
rect 2502 2141 2508 2142
rect 2502 2137 2503 2141
rect 2507 2137 2508 2141
rect 2502 2136 2508 2137
rect 2502 2124 2508 2125
rect 2502 2120 2503 2124
rect 2507 2120 2508 2124
rect 2502 2119 2508 2120
rect 2470 2103 2476 2104
rect 2470 2099 2471 2103
rect 2475 2099 2476 2103
rect 2470 2098 2476 2099
rect 2504 2087 2506 2119
rect 2503 2086 2507 2087
rect 2503 2081 2507 2082
rect 2462 2075 2468 2076
rect 2462 2071 2463 2075
rect 2467 2071 2468 2075
rect 2462 2070 2468 2071
rect 2454 2061 2460 2062
rect 2504 2061 2506 2081
rect 2318 2056 2324 2057
rect 2334 2059 2340 2060
rect 2334 2055 2335 2059
rect 2339 2055 2340 2059
rect 2454 2057 2455 2061
rect 2459 2057 2460 2061
rect 2502 2060 2508 2061
rect 2454 2056 2460 2057
rect 2470 2059 2476 2060
rect 2334 2054 2340 2055
rect 2470 2055 2471 2059
rect 2475 2055 2476 2059
rect 2502 2056 2503 2060
rect 2507 2056 2508 2060
rect 2502 2055 2508 2056
rect 2470 2054 2476 2055
rect 1878 2040 1884 2041
rect 1878 2036 1879 2040
rect 1883 2036 1884 2040
rect 1878 2035 1884 2036
rect 2006 2040 2012 2041
rect 2006 2036 2007 2040
rect 2011 2036 2012 2040
rect 2006 2035 2012 2036
rect 2150 2040 2156 2041
rect 2150 2036 2151 2040
rect 2155 2036 2156 2040
rect 2150 2035 2156 2036
rect 2302 2040 2308 2041
rect 2302 2036 2303 2040
rect 2307 2036 2308 2040
rect 2302 2035 2308 2036
rect 2438 2040 2444 2041
rect 2438 2036 2439 2040
rect 2443 2036 2444 2040
rect 2438 2035 2444 2036
rect 1879 2034 1883 2035
rect 1879 2029 1883 2030
rect 1935 2034 1939 2035
rect 1935 2029 1939 2030
rect 2007 2034 2011 2035
rect 2007 2029 2011 2030
rect 2055 2034 2059 2035
rect 2055 2029 2059 2030
rect 2151 2034 2155 2035
rect 2151 2029 2155 2030
rect 2183 2034 2187 2035
rect 2183 2029 2187 2030
rect 2303 2034 2307 2035
rect 2303 2029 2307 2030
rect 2319 2034 2323 2035
rect 2319 2029 2323 2030
rect 2439 2034 2443 2035
rect 2439 2029 2443 2030
rect 1934 2028 1940 2029
rect 1934 2024 1935 2028
rect 1939 2024 1940 2028
rect 1934 2023 1940 2024
rect 2054 2028 2060 2029
rect 2054 2024 2055 2028
rect 2059 2024 2060 2028
rect 2054 2023 2060 2024
rect 2182 2028 2188 2029
rect 2182 2024 2183 2028
rect 2187 2024 2188 2028
rect 2182 2023 2188 2024
rect 2318 2028 2324 2029
rect 2318 2024 2319 2028
rect 2323 2024 2324 2028
rect 2318 2023 2324 2024
rect 2438 2028 2444 2029
rect 2438 2024 2439 2028
rect 2443 2024 2444 2028
rect 2438 2023 2444 2024
rect 1734 2007 1740 2008
rect 1734 2003 1735 2007
rect 1739 2003 1740 2007
rect 1734 2002 1740 2003
rect 1742 2007 1748 2008
rect 1742 2003 1743 2007
rect 1747 2003 1748 2007
rect 1742 2002 1748 2003
rect 1838 2007 1844 2008
rect 1838 2003 1839 2007
rect 1843 2003 1844 2007
rect 1838 2002 1844 2003
rect 1858 2007 1864 2008
rect 1858 2003 1859 2007
rect 1863 2003 1864 2007
rect 1858 2002 1864 2003
rect 1950 2007 1956 2008
rect 1950 2003 1951 2007
rect 1955 2003 1956 2007
rect 1950 2002 1956 2003
rect 1966 2007 1972 2008
rect 1966 2003 1967 2007
rect 1971 2003 1972 2007
rect 1966 2002 1972 2003
rect 2070 2007 2076 2008
rect 2070 2003 2071 2007
rect 2075 2003 2076 2007
rect 2070 2002 2076 2003
rect 2198 2007 2204 2008
rect 2198 2003 2199 2007
rect 2203 2003 2204 2007
rect 2198 2002 2204 2003
rect 2334 2007 2340 2008
rect 2334 2003 2335 2007
rect 2339 2003 2340 2007
rect 2334 2002 2340 2003
rect 2342 2007 2348 2008
rect 2342 2003 2343 2007
rect 2347 2003 2348 2007
rect 2342 2002 2348 2003
rect 2454 2007 2460 2008
rect 2454 2003 2455 2007
rect 2459 2003 2460 2007
rect 2454 2002 2460 2003
rect 2462 2007 2468 2008
rect 2462 2003 2463 2007
rect 2467 2003 2468 2007
rect 2462 2002 2468 2003
rect 1686 1987 1692 1988
rect 1686 1983 1687 1987
rect 1691 1983 1692 1987
rect 1686 1982 1692 1983
rect 1736 1979 1738 2002
rect 1327 1978 1331 1979
rect 1014 1975 1020 1976
rect 1286 1977 1292 1978
rect 1286 1973 1287 1977
rect 1291 1973 1292 1977
rect 1327 1973 1331 1974
rect 1367 1978 1371 1979
rect 1367 1973 1371 1974
rect 1439 1978 1443 1979
rect 1439 1973 1443 1974
rect 1455 1978 1459 1979
rect 1455 1973 1459 1974
rect 1535 1978 1539 1979
rect 1535 1973 1539 1974
rect 1543 1978 1547 1979
rect 1543 1973 1547 1974
rect 1631 1978 1635 1979
rect 1631 1973 1635 1974
rect 1639 1978 1643 1979
rect 1639 1973 1643 1974
rect 1735 1978 1739 1979
rect 1744 1976 1746 2002
rect 1840 1979 1842 2002
rect 1952 1979 1954 2002
rect 1968 1988 1970 2002
rect 1966 1987 1972 1988
rect 1966 1983 1967 1987
rect 1971 1983 1972 1987
rect 1966 1982 1972 1983
rect 2072 1979 2074 2002
rect 2114 1999 2120 2000
rect 2114 1995 2115 1999
rect 2119 1995 2120 1999
rect 2114 1994 2120 1995
rect 1839 1978 1843 1979
rect 1735 1973 1739 1974
rect 1742 1975 1748 1976
rect 1286 1972 1292 1973
rect 1286 1960 1292 1961
rect 502 1959 508 1960
rect 502 1955 503 1959
rect 507 1955 508 1959
rect 502 1954 508 1955
rect 606 1959 612 1960
rect 606 1955 607 1959
rect 611 1955 612 1959
rect 606 1954 612 1955
rect 614 1959 620 1960
rect 614 1955 615 1959
rect 619 1955 620 1959
rect 614 1954 620 1955
rect 710 1959 716 1960
rect 710 1955 711 1959
rect 715 1955 716 1959
rect 710 1954 716 1955
rect 726 1959 732 1960
rect 726 1955 727 1959
rect 731 1955 732 1959
rect 726 1954 732 1955
rect 814 1959 820 1960
rect 814 1955 815 1959
rect 819 1955 820 1959
rect 814 1954 820 1955
rect 918 1959 924 1960
rect 918 1955 919 1959
rect 923 1955 924 1959
rect 918 1954 924 1955
rect 1030 1959 1036 1960
rect 1030 1955 1031 1959
rect 1035 1955 1036 1959
rect 1030 1954 1036 1955
rect 1038 1959 1044 1960
rect 1038 1955 1039 1959
rect 1043 1955 1044 1959
rect 1286 1956 1287 1960
rect 1291 1956 1292 1960
rect 1286 1955 1292 1956
rect 1038 1954 1044 1955
rect 406 1943 412 1944
rect 406 1939 407 1943
rect 411 1939 412 1943
rect 406 1938 412 1939
rect 504 1927 506 1954
rect 608 1927 610 1954
rect 616 1936 618 1954
rect 614 1935 620 1936
rect 614 1931 615 1935
rect 619 1931 620 1935
rect 614 1930 620 1931
rect 712 1927 714 1954
rect 816 1927 818 1954
rect 886 1943 892 1944
rect 886 1939 887 1943
rect 891 1939 892 1943
rect 886 1938 892 1939
rect 375 1926 379 1927
rect 375 1921 379 1922
rect 399 1926 403 1927
rect 399 1921 403 1922
rect 503 1926 507 1927
rect 503 1921 507 1922
rect 527 1926 531 1927
rect 527 1921 531 1922
rect 607 1926 611 1927
rect 607 1921 611 1922
rect 687 1926 691 1927
rect 711 1926 715 1927
rect 687 1921 691 1922
rect 702 1923 708 1924
rect 366 1915 372 1916
rect 366 1911 367 1915
rect 371 1911 372 1915
rect 366 1910 372 1911
rect 376 1902 378 1921
rect 528 1902 530 1921
rect 688 1902 690 1921
rect 702 1919 703 1923
rect 707 1919 708 1923
rect 711 1921 715 1922
rect 815 1926 819 1927
rect 815 1921 819 1922
rect 863 1926 867 1927
rect 863 1921 867 1922
rect 702 1918 708 1919
rect 150 1901 156 1902
rect 110 1900 116 1901
rect 110 1896 111 1900
rect 115 1896 116 1900
rect 150 1897 151 1901
rect 155 1897 156 1901
rect 238 1901 244 1902
rect 150 1896 156 1897
rect 198 1899 204 1900
rect 110 1895 116 1896
rect 198 1895 199 1899
rect 203 1895 204 1899
rect 238 1897 239 1901
rect 243 1897 244 1901
rect 238 1896 244 1897
rect 374 1901 380 1902
rect 374 1897 375 1901
rect 379 1897 380 1901
rect 374 1896 380 1897
rect 526 1901 532 1902
rect 526 1897 527 1901
rect 531 1897 532 1901
rect 526 1896 532 1897
rect 686 1901 692 1902
rect 686 1897 687 1901
rect 691 1897 692 1901
rect 704 1900 706 1918
rect 864 1902 866 1921
rect 862 1901 868 1902
rect 686 1896 692 1897
rect 702 1899 708 1900
rect 198 1894 204 1895
rect 702 1895 703 1899
rect 707 1895 708 1899
rect 862 1897 863 1901
rect 867 1897 868 1901
rect 888 1900 890 1938
rect 920 1927 922 1954
rect 1032 1927 1034 1954
rect 1040 1936 1042 1954
rect 1038 1935 1044 1936
rect 1038 1931 1039 1935
rect 1043 1931 1044 1935
rect 1038 1930 1044 1931
rect 1288 1927 1290 1955
rect 1328 1953 1330 1973
rect 1456 1954 1458 1973
rect 1544 1954 1546 1973
rect 1640 1954 1642 1973
rect 1736 1954 1738 1973
rect 1742 1971 1743 1975
rect 1747 1971 1748 1975
rect 1839 1973 1843 1974
rect 1943 1978 1947 1979
rect 1943 1973 1947 1974
rect 1951 1978 1955 1979
rect 1951 1973 1955 1974
rect 2047 1978 2051 1979
rect 2047 1973 2051 1974
rect 2071 1978 2075 1979
rect 2116 1976 2118 1994
rect 2174 1991 2180 1992
rect 2174 1987 2175 1991
rect 2179 1987 2180 1991
rect 2174 1986 2180 1987
rect 2151 1978 2155 1979
rect 2071 1973 2075 1974
rect 2114 1975 2120 1976
rect 1742 1970 1748 1971
rect 1840 1954 1842 1973
rect 1944 1954 1946 1973
rect 2048 1954 2050 1973
rect 2114 1971 2115 1975
rect 2119 1971 2120 1975
rect 2151 1973 2155 1974
rect 2114 1970 2120 1971
rect 2152 1954 2154 1973
rect 1454 1953 1460 1954
rect 1326 1952 1332 1953
rect 1326 1948 1327 1952
rect 1331 1948 1332 1952
rect 1454 1949 1455 1953
rect 1459 1949 1460 1953
rect 1454 1948 1460 1949
rect 1542 1953 1548 1954
rect 1542 1949 1543 1953
rect 1547 1949 1548 1953
rect 1542 1948 1548 1949
rect 1638 1953 1644 1954
rect 1638 1949 1639 1953
rect 1643 1949 1644 1953
rect 1638 1948 1644 1949
rect 1734 1953 1740 1954
rect 1734 1949 1735 1953
rect 1739 1949 1740 1953
rect 1734 1948 1740 1949
rect 1838 1953 1844 1954
rect 1838 1949 1839 1953
rect 1843 1949 1844 1953
rect 1942 1953 1948 1954
rect 1838 1948 1844 1949
rect 1846 1951 1852 1952
rect 1326 1947 1332 1948
rect 1846 1947 1847 1951
rect 1851 1947 1852 1951
rect 1942 1949 1943 1953
rect 1947 1949 1948 1953
rect 1942 1948 1948 1949
rect 2046 1953 2052 1954
rect 2046 1949 2047 1953
rect 2051 1949 2052 1953
rect 2046 1948 2052 1949
rect 2150 1953 2156 1954
rect 2150 1949 2151 1953
rect 2155 1949 2156 1953
rect 2176 1952 2178 1986
rect 2200 1979 2202 2002
rect 2310 1999 2316 2000
rect 2310 1995 2311 1999
rect 2315 1995 2316 1999
rect 2310 1994 2316 1995
rect 2199 1978 2203 1979
rect 2199 1973 2203 1974
rect 2255 1978 2259 1979
rect 2255 1973 2259 1974
rect 2246 1967 2252 1968
rect 2246 1963 2247 1967
rect 2251 1963 2252 1967
rect 2246 1962 2252 1963
rect 2150 1948 2156 1949
rect 2174 1951 2180 1952
rect 1846 1946 1852 1947
rect 2174 1947 2175 1951
rect 2179 1947 2180 1951
rect 2174 1946 2180 1947
rect 1326 1935 1332 1936
rect 1326 1931 1327 1935
rect 1331 1931 1332 1935
rect 1326 1930 1332 1931
rect 1438 1932 1444 1933
rect 919 1926 923 1927
rect 919 1921 923 1922
rect 1031 1926 1035 1927
rect 1031 1921 1035 1922
rect 1039 1926 1043 1927
rect 1039 1921 1043 1922
rect 1287 1926 1291 1927
rect 1328 1923 1330 1930
rect 1438 1928 1439 1932
rect 1443 1928 1444 1932
rect 1438 1927 1444 1928
rect 1526 1932 1532 1933
rect 1526 1928 1527 1932
rect 1531 1928 1532 1932
rect 1526 1927 1532 1928
rect 1622 1932 1628 1933
rect 1622 1928 1623 1932
rect 1627 1928 1628 1932
rect 1622 1927 1628 1928
rect 1718 1932 1724 1933
rect 1718 1928 1719 1932
rect 1723 1928 1724 1932
rect 1718 1927 1724 1928
rect 1822 1932 1828 1933
rect 1822 1928 1823 1932
rect 1827 1928 1828 1932
rect 1822 1927 1828 1928
rect 1440 1923 1442 1927
rect 1528 1923 1530 1927
rect 1624 1923 1626 1927
rect 1720 1923 1722 1927
rect 1824 1923 1826 1927
rect 1287 1921 1291 1922
rect 1327 1922 1331 1923
rect 1040 1902 1042 1921
rect 1074 1915 1080 1916
rect 1074 1911 1075 1915
rect 1079 1911 1080 1915
rect 1074 1910 1080 1911
rect 1038 1901 1044 1902
rect 862 1896 868 1897
rect 886 1899 892 1900
rect 702 1894 708 1895
rect 886 1895 887 1899
rect 891 1895 892 1899
rect 1038 1897 1039 1901
rect 1043 1897 1044 1901
rect 1038 1896 1044 1897
rect 886 1894 892 1895
rect 110 1883 116 1884
rect 110 1879 111 1883
rect 115 1879 116 1883
rect 110 1878 116 1879
rect 134 1880 140 1881
rect 112 1875 114 1878
rect 134 1876 135 1880
rect 139 1876 140 1880
rect 134 1875 140 1876
rect 111 1874 115 1875
rect 111 1869 115 1870
rect 135 1874 139 1875
rect 135 1869 139 1870
rect 191 1874 195 1875
rect 191 1869 195 1870
rect 112 1866 114 1869
rect 134 1868 140 1869
rect 110 1865 116 1866
rect 110 1861 111 1865
rect 115 1861 116 1865
rect 134 1864 135 1868
rect 139 1864 140 1868
rect 134 1863 140 1864
rect 190 1868 196 1869
rect 190 1864 191 1868
rect 195 1864 196 1868
rect 190 1863 196 1864
rect 110 1860 116 1861
rect 110 1848 116 1849
rect 110 1844 111 1848
rect 115 1844 116 1848
rect 110 1843 116 1844
rect 150 1847 156 1848
rect 150 1843 151 1847
rect 155 1843 156 1847
rect 112 1815 114 1843
rect 150 1842 156 1843
rect 158 1847 164 1848
rect 158 1843 159 1847
rect 163 1843 164 1847
rect 158 1842 164 1843
rect 152 1815 154 1842
rect 111 1814 115 1815
rect 111 1809 115 1810
rect 151 1814 155 1815
rect 151 1809 155 1810
rect 112 1789 114 1809
rect 152 1790 154 1809
rect 160 1804 162 1842
rect 200 1832 202 1894
rect 222 1880 228 1881
rect 222 1876 223 1880
rect 227 1876 228 1880
rect 222 1875 228 1876
rect 358 1880 364 1881
rect 358 1876 359 1880
rect 363 1876 364 1880
rect 358 1875 364 1876
rect 510 1880 516 1881
rect 510 1876 511 1880
rect 515 1876 516 1880
rect 510 1875 516 1876
rect 670 1880 676 1881
rect 670 1876 671 1880
rect 675 1876 676 1880
rect 670 1875 676 1876
rect 846 1880 852 1881
rect 846 1876 847 1880
rect 851 1876 852 1880
rect 846 1875 852 1876
rect 1022 1880 1028 1881
rect 1022 1876 1023 1880
rect 1027 1876 1028 1880
rect 1022 1875 1028 1876
rect 223 1874 227 1875
rect 223 1869 227 1870
rect 263 1874 267 1875
rect 263 1869 267 1870
rect 335 1874 339 1875
rect 335 1869 339 1870
rect 359 1874 363 1875
rect 359 1869 363 1870
rect 407 1874 411 1875
rect 407 1869 411 1870
rect 479 1874 483 1875
rect 479 1869 483 1870
rect 511 1874 515 1875
rect 511 1869 515 1870
rect 551 1874 555 1875
rect 551 1869 555 1870
rect 615 1874 619 1875
rect 615 1869 619 1870
rect 671 1874 675 1875
rect 671 1869 675 1870
rect 679 1874 683 1875
rect 679 1869 683 1870
rect 743 1874 747 1875
rect 743 1869 747 1870
rect 815 1874 819 1875
rect 815 1869 819 1870
rect 847 1874 851 1875
rect 847 1869 851 1870
rect 887 1874 891 1875
rect 887 1869 891 1870
rect 959 1874 963 1875
rect 959 1869 963 1870
rect 1023 1874 1027 1875
rect 1023 1869 1027 1870
rect 1039 1874 1043 1875
rect 1039 1869 1043 1870
rect 262 1868 268 1869
rect 262 1864 263 1868
rect 267 1864 268 1868
rect 262 1863 268 1864
rect 334 1868 340 1869
rect 334 1864 335 1868
rect 339 1864 340 1868
rect 334 1863 340 1864
rect 406 1868 412 1869
rect 406 1864 407 1868
rect 411 1864 412 1868
rect 406 1863 412 1864
rect 478 1868 484 1869
rect 478 1864 479 1868
rect 483 1864 484 1868
rect 478 1863 484 1864
rect 550 1868 556 1869
rect 550 1864 551 1868
rect 555 1864 556 1868
rect 550 1863 556 1864
rect 614 1868 620 1869
rect 614 1864 615 1868
rect 619 1864 620 1868
rect 614 1863 620 1864
rect 678 1868 684 1869
rect 678 1864 679 1868
rect 683 1864 684 1868
rect 678 1863 684 1864
rect 742 1868 748 1869
rect 742 1864 743 1868
rect 747 1864 748 1868
rect 742 1863 748 1864
rect 814 1868 820 1869
rect 814 1864 815 1868
rect 819 1864 820 1868
rect 814 1863 820 1864
rect 886 1868 892 1869
rect 886 1864 887 1868
rect 891 1864 892 1868
rect 886 1863 892 1864
rect 958 1868 964 1869
rect 958 1864 959 1868
rect 963 1864 964 1868
rect 958 1863 964 1864
rect 1038 1868 1044 1869
rect 1038 1864 1039 1868
rect 1043 1864 1044 1868
rect 1038 1863 1044 1864
rect 1076 1848 1078 1910
rect 1288 1901 1290 1921
rect 1327 1917 1331 1918
rect 1439 1922 1443 1923
rect 1439 1917 1443 1918
rect 1527 1922 1531 1923
rect 1527 1917 1531 1918
rect 1615 1922 1619 1923
rect 1615 1917 1619 1918
rect 1623 1922 1627 1923
rect 1623 1917 1627 1918
rect 1711 1922 1715 1923
rect 1711 1917 1715 1918
rect 1719 1922 1723 1923
rect 1719 1917 1723 1918
rect 1815 1922 1819 1923
rect 1815 1917 1819 1918
rect 1823 1922 1827 1923
rect 1823 1917 1827 1918
rect 1328 1914 1330 1917
rect 1526 1916 1532 1917
rect 1326 1913 1332 1914
rect 1326 1909 1327 1913
rect 1331 1909 1332 1913
rect 1526 1912 1527 1916
rect 1531 1912 1532 1916
rect 1526 1911 1532 1912
rect 1614 1916 1620 1917
rect 1614 1912 1615 1916
rect 1619 1912 1620 1916
rect 1614 1911 1620 1912
rect 1710 1916 1716 1917
rect 1710 1912 1711 1916
rect 1715 1912 1716 1916
rect 1710 1911 1716 1912
rect 1814 1916 1820 1917
rect 1814 1912 1815 1916
rect 1819 1912 1820 1916
rect 1814 1911 1820 1912
rect 1326 1908 1332 1909
rect 1286 1900 1292 1901
rect 1286 1896 1287 1900
rect 1291 1896 1292 1900
rect 1286 1895 1292 1896
rect 1326 1896 1332 1897
rect 1326 1892 1327 1896
rect 1331 1892 1332 1896
rect 1326 1891 1332 1892
rect 1542 1895 1548 1896
rect 1542 1891 1543 1895
rect 1547 1891 1548 1895
rect 1286 1883 1292 1884
rect 1286 1879 1287 1883
rect 1291 1879 1292 1883
rect 1286 1878 1292 1879
rect 1288 1875 1290 1878
rect 1287 1874 1291 1875
rect 1328 1871 1330 1891
rect 1542 1890 1548 1891
rect 1630 1895 1636 1896
rect 1630 1891 1631 1895
rect 1635 1891 1636 1895
rect 1630 1890 1636 1891
rect 1726 1895 1732 1896
rect 1726 1891 1727 1895
rect 1731 1891 1732 1895
rect 1726 1890 1732 1891
rect 1830 1895 1836 1896
rect 1830 1891 1831 1895
rect 1835 1891 1836 1895
rect 1830 1890 1836 1891
rect 1544 1871 1546 1890
rect 1632 1871 1634 1890
rect 1728 1871 1730 1890
rect 1832 1871 1834 1890
rect 1848 1876 1850 1946
rect 1926 1932 1932 1933
rect 1926 1928 1927 1932
rect 1931 1928 1932 1932
rect 1926 1927 1932 1928
rect 2030 1932 2036 1933
rect 2030 1928 2031 1932
rect 2035 1928 2036 1932
rect 2030 1927 2036 1928
rect 2134 1932 2140 1933
rect 2134 1928 2135 1932
rect 2139 1928 2140 1932
rect 2134 1927 2140 1928
rect 2238 1932 2244 1933
rect 2238 1928 2239 1932
rect 2243 1928 2244 1932
rect 2238 1927 2244 1928
rect 1928 1923 1930 1927
rect 2032 1923 2034 1927
rect 2136 1923 2138 1927
rect 2240 1923 2242 1927
rect 1919 1922 1923 1923
rect 1919 1917 1923 1918
rect 1927 1922 1931 1923
rect 1927 1917 1931 1918
rect 2015 1922 2019 1923
rect 2015 1917 2019 1918
rect 2031 1922 2035 1923
rect 2031 1917 2035 1918
rect 2111 1922 2115 1923
rect 2111 1917 2115 1918
rect 2135 1922 2139 1923
rect 2135 1917 2139 1918
rect 2199 1922 2203 1923
rect 2199 1917 2203 1918
rect 2239 1922 2243 1923
rect 2239 1917 2243 1918
rect 1918 1916 1924 1917
rect 1918 1912 1919 1916
rect 1923 1912 1924 1916
rect 1918 1911 1924 1912
rect 2014 1916 2020 1917
rect 2014 1912 2015 1916
rect 2019 1912 2020 1916
rect 2014 1911 2020 1912
rect 2110 1916 2116 1917
rect 2110 1912 2111 1916
rect 2115 1912 2116 1916
rect 2110 1911 2116 1912
rect 2198 1916 2204 1917
rect 2198 1912 2199 1916
rect 2203 1912 2204 1916
rect 2198 1911 2204 1912
rect 2248 1896 2250 1962
rect 2256 1954 2258 1973
rect 2312 1960 2314 1994
rect 2336 1979 2338 2002
rect 2344 1984 2346 2002
rect 2342 1983 2348 1984
rect 2342 1979 2343 1983
rect 2347 1979 2348 1983
rect 2456 1979 2458 2002
rect 2335 1978 2339 1979
rect 2342 1978 2348 1979
rect 2367 1978 2371 1979
rect 2335 1973 2339 1974
rect 2367 1973 2371 1974
rect 2455 1978 2459 1979
rect 2455 1973 2459 1974
rect 2310 1959 2316 1960
rect 2310 1955 2311 1959
rect 2315 1955 2316 1959
rect 2310 1954 2316 1955
rect 2368 1954 2370 1973
rect 2456 1954 2458 1973
rect 2464 1968 2466 2002
rect 2472 1992 2474 2054
rect 2502 2043 2508 2044
rect 2502 2039 2503 2043
rect 2507 2039 2508 2043
rect 2502 2038 2508 2039
rect 2504 2035 2506 2038
rect 2503 2034 2507 2035
rect 2503 2029 2507 2030
rect 2504 2026 2506 2029
rect 2502 2025 2508 2026
rect 2502 2021 2503 2025
rect 2507 2021 2508 2025
rect 2502 2020 2508 2021
rect 2502 2008 2508 2009
rect 2502 2004 2503 2008
rect 2507 2004 2508 2008
rect 2502 2003 2508 2004
rect 2470 1991 2476 1992
rect 2470 1987 2471 1991
rect 2475 1987 2476 1991
rect 2470 1986 2476 1987
rect 2504 1979 2506 2003
rect 2503 1978 2507 1979
rect 2503 1973 2507 1974
rect 2462 1967 2468 1968
rect 2462 1963 2463 1967
rect 2467 1963 2468 1967
rect 2462 1962 2468 1963
rect 2254 1953 2260 1954
rect 2254 1949 2255 1953
rect 2259 1949 2260 1953
rect 2254 1948 2260 1949
rect 2366 1953 2372 1954
rect 2366 1949 2367 1953
rect 2371 1949 2372 1953
rect 2366 1948 2372 1949
rect 2454 1953 2460 1954
rect 2504 1953 2506 1973
rect 2454 1949 2455 1953
rect 2459 1949 2460 1953
rect 2502 1952 2508 1953
rect 2454 1948 2460 1949
rect 2462 1951 2468 1952
rect 2462 1947 2463 1951
rect 2467 1947 2468 1951
rect 2502 1948 2503 1952
rect 2507 1948 2508 1952
rect 2502 1947 2508 1948
rect 2462 1946 2468 1947
rect 2350 1932 2356 1933
rect 2350 1928 2351 1932
rect 2355 1928 2356 1932
rect 2350 1927 2356 1928
rect 2438 1932 2444 1933
rect 2438 1928 2439 1932
rect 2443 1928 2444 1932
rect 2438 1927 2444 1928
rect 2352 1923 2354 1927
rect 2440 1923 2442 1927
rect 2287 1922 2291 1923
rect 2287 1917 2291 1918
rect 2351 1922 2355 1923
rect 2351 1917 2355 1918
rect 2375 1922 2379 1923
rect 2375 1917 2379 1918
rect 2439 1922 2443 1923
rect 2439 1917 2443 1918
rect 2286 1916 2292 1917
rect 2286 1912 2287 1916
rect 2291 1912 2292 1916
rect 2286 1911 2292 1912
rect 2374 1916 2380 1917
rect 2374 1912 2375 1916
rect 2379 1912 2380 1916
rect 2374 1911 2380 1912
rect 2438 1916 2444 1917
rect 2438 1912 2439 1916
rect 2443 1912 2444 1916
rect 2438 1911 2444 1912
rect 1934 1895 1940 1896
rect 1934 1891 1935 1895
rect 1939 1891 1940 1895
rect 1934 1890 1940 1891
rect 1974 1895 1980 1896
rect 1974 1891 1975 1895
rect 1979 1891 1980 1895
rect 1974 1890 1980 1891
rect 2030 1895 2036 1896
rect 2030 1891 2031 1895
rect 2035 1891 2036 1895
rect 2030 1890 2036 1891
rect 2126 1895 2132 1896
rect 2126 1891 2127 1895
rect 2131 1891 2132 1895
rect 2126 1890 2132 1891
rect 2214 1895 2220 1896
rect 2214 1891 2215 1895
rect 2219 1891 2220 1895
rect 2214 1890 2220 1891
rect 2246 1895 2252 1896
rect 2246 1891 2247 1895
rect 2251 1891 2252 1895
rect 2246 1890 2252 1891
rect 2302 1895 2308 1896
rect 2302 1891 2303 1895
rect 2307 1891 2308 1895
rect 2302 1890 2308 1891
rect 2318 1895 2324 1896
rect 2318 1891 2319 1895
rect 2323 1891 2324 1895
rect 2318 1890 2324 1891
rect 2390 1895 2396 1896
rect 2390 1891 2391 1895
rect 2395 1891 2396 1895
rect 2390 1890 2396 1891
rect 2454 1895 2460 1896
rect 2454 1891 2455 1895
rect 2459 1891 2460 1895
rect 2454 1890 2460 1891
rect 1846 1875 1852 1876
rect 1846 1871 1847 1875
rect 1851 1871 1852 1875
rect 1936 1871 1938 1890
rect 1287 1869 1291 1870
rect 1327 1870 1331 1871
rect 1288 1866 1290 1869
rect 1286 1865 1292 1866
rect 1327 1865 1331 1866
rect 1535 1870 1539 1871
rect 1535 1865 1539 1866
rect 1543 1870 1547 1871
rect 1543 1865 1547 1866
rect 1607 1870 1611 1871
rect 1607 1865 1611 1866
rect 1631 1870 1635 1871
rect 1631 1865 1635 1866
rect 1687 1870 1691 1871
rect 1687 1865 1691 1866
rect 1727 1870 1731 1871
rect 1727 1865 1731 1866
rect 1783 1870 1787 1871
rect 1831 1870 1835 1871
rect 1846 1870 1852 1871
rect 1879 1870 1883 1871
rect 1783 1865 1787 1866
rect 1802 1867 1808 1868
rect 1286 1861 1287 1865
rect 1291 1861 1292 1865
rect 1286 1860 1292 1861
rect 1286 1848 1292 1849
rect 206 1847 212 1848
rect 206 1843 207 1847
rect 211 1843 212 1847
rect 206 1842 212 1843
rect 278 1847 284 1848
rect 278 1843 279 1847
rect 283 1843 284 1847
rect 278 1842 284 1843
rect 350 1847 356 1848
rect 350 1843 351 1847
rect 355 1843 356 1847
rect 350 1842 356 1843
rect 358 1847 364 1848
rect 358 1843 359 1847
rect 363 1843 364 1847
rect 358 1842 364 1843
rect 422 1847 428 1848
rect 422 1843 423 1847
rect 427 1843 428 1847
rect 422 1842 428 1843
rect 494 1847 500 1848
rect 494 1843 495 1847
rect 499 1843 500 1847
rect 494 1842 500 1843
rect 566 1847 572 1848
rect 566 1843 567 1847
rect 571 1843 572 1847
rect 566 1842 572 1843
rect 630 1847 636 1848
rect 630 1843 631 1847
rect 635 1843 636 1847
rect 630 1842 636 1843
rect 694 1847 700 1848
rect 694 1843 695 1847
rect 699 1843 700 1847
rect 694 1842 700 1843
rect 758 1847 764 1848
rect 758 1843 759 1847
rect 763 1843 764 1847
rect 758 1842 764 1843
rect 830 1847 836 1848
rect 830 1843 831 1847
rect 835 1843 836 1847
rect 830 1842 836 1843
rect 902 1847 908 1848
rect 902 1843 903 1847
rect 907 1843 908 1847
rect 902 1842 908 1843
rect 974 1847 980 1848
rect 974 1843 975 1847
rect 979 1843 980 1847
rect 974 1842 980 1843
rect 982 1847 988 1848
rect 982 1843 983 1847
rect 987 1843 988 1847
rect 982 1842 988 1843
rect 1054 1847 1060 1848
rect 1054 1843 1055 1847
rect 1059 1843 1060 1847
rect 1054 1842 1060 1843
rect 1074 1847 1080 1848
rect 1074 1843 1075 1847
rect 1079 1843 1080 1847
rect 1286 1844 1287 1848
rect 1291 1844 1292 1848
rect 1328 1845 1330 1865
rect 1536 1846 1538 1865
rect 1608 1846 1610 1865
rect 1688 1846 1690 1865
rect 1784 1846 1786 1865
rect 1802 1863 1803 1867
rect 1807 1863 1808 1867
rect 1831 1865 1835 1866
rect 1879 1865 1883 1866
rect 1935 1870 1939 1871
rect 1935 1865 1939 1866
rect 1802 1862 1808 1863
rect 1534 1845 1540 1846
rect 1286 1843 1292 1844
rect 1326 1844 1332 1845
rect 1074 1842 1080 1843
rect 198 1831 204 1832
rect 198 1827 199 1831
rect 203 1827 204 1831
rect 198 1826 204 1827
rect 208 1815 210 1842
rect 280 1815 282 1842
rect 352 1815 354 1842
rect 360 1824 362 1842
rect 358 1823 364 1824
rect 358 1819 359 1823
rect 363 1819 364 1823
rect 358 1818 364 1819
rect 424 1815 426 1842
rect 458 1831 464 1832
rect 458 1827 459 1831
rect 463 1827 464 1831
rect 458 1826 464 1827
rect 207 1814 211 1815
rect 207 1809 211 1810
rect 231 1814 235 1815
rect 231 1809 235 1810
rect 279 1814 283 1815
rect 279 1809 283 1810
rect 335 1814 339 1815
rect 335 1809 339 1810
rect 351 1814 355 1815
rect 351 1809 355 1810
rect 423 1814 427 1815
rect 423 1809 427 1810
rect 439 1814 443 1815
rect 439 1809 443 1810
rect 158 1803 164 1804
rect 158 1799 159 1803
rect 163 1799 164 1803
rect 158 1798 164 1799
rect 232 1790 234 1809
rect 336 1790 338 1809
rect 440 1790 442 1809
rect 150 1789 156 1790
rect 110 1788 116 1789
rect 110 1784 111 1788
rect 115 1784 116 1788
rect 150 1785 151 1789
rect 155 1785 156 1789
rect 150 1784 156 1785
rect 230 1789 236 1790
rect 230 1785 231 1789
rect 235 1785 236 1789
rect 230 1784 236 1785
rect 334 1789 340 1790
rect 334 1785 335 1789
rect 339 1785 340 1789
rect 438 1789 444 1790
rect 334 1784 340 1785
rect 358 1787 364 1788
rect 110 1783 116 1784
rect 358 1783 359 1787
rect 363 1783 364 1787
rect 438 1785 439 1789
rect 443 1785 444 1789
rect 460 1788 462 1826
rect 496 1815 498 1842
rect 568 1815 570 1842
rect 632 1815 634 1842
rect 696 1815 698 1842
rect 760 1815 762 1842
rect 832 1815 834 1842
rect 904 1815 906 1842
rect 976 1815 978 1842
rect 495 1814 499 1815
rect 495 1809 499 1810
rect 535 1814 539 1815
rect 535 1809 539 1810
rect 567 1814 571 1815
rect 567 1809 571 1810
rect 631 1814 635 1815
rect 695 1814 699 1815
rect 631 1809 635 1810
rect 650 1811 656 1812
rect 498 1803 504 1804
rect 498 1799 499 1803
rect 503 1799 504 1803
rect 498 1798 504 1799
rect 438 1784 444 1785
rect 458 1787 464 1788
rect 358 1782 364 1783
rect 458 1783 459 1787
rect 463 1783 464 1787
rect 458 1782 464 1783
rect 110 1771 116 1772
rect 110 1767 111 1771
rect 115 1767 116 1771
rect 110 1766 116 1767
rect 134 1768 140 1769
rect 112 1759 114 1766
rect 134 1764 135 1768
rect 139 1764 140 1768
rect 134 1763 140 1764
rect 214 1768 220 1769
rect 214 1764 215 1768
rect 219 1764 220 1768
rect 214 1763 220 1764
rect 318 1768 324 1769
rect 318 1764 319 1768
rect 323 1764 324 1768
rect 318 1763 324 1764
rect 136 1759 138 1763
rect 216 1759 218 1763
rect 320 1759 322 1763
rect 111 1758 115 1759
rect 111 1753 115 1754
rect 135 1758 139 1759
rect 135 1753 139 1754
rect 215 1758 219 1759
rect 215 1753 219 1754
rect 239 1758 243 1759
rect 239 1753 243 1754
rect 319 1758 323 1759
rect 319 1753 323 1754
rect 351 1758 355 1759
rect 351 1753 355 1754
rect 112 1750 114 1753
rect 134 1752 140 1753
rect 110 1749 116 1750
rect 110 1745 111 1749
rect 115 1745 116 1749
rect 134 1748 135 1752
rect 139 1748 140 1752
rect 134 1747 140 1748
rect 238 1752 244 1753
rect 238 1748 239 1752
rect 243 1748 244 1752
rect 238 1747 244 1748
rect 350 1752 356 1753
rect 350 1748 351 1752
rect 355 1748 356 1752
rect 350 1747 356 1748
rect 110 1744 116 1745
rect 110 1732 116 1733
rect 110 1728 111 1732
rect 115 1728 116 1732
rect 110 1727 116 1728
rect 150 1731 156 1732
rect 150 1727 151 1731
rect 155 1727 156 1731
rect 112 1703 114 1727
rect 150 1726 156 1727
rect 182 1731 188 1732
rect 182 1727 183 1731
rect 187 1727 188 1731
rect 182 1726 188 1727
rect 254 1731 260 1732
rect 254 1727 255 1731
rect 259 1727 260 1731
rect 254 1726 260 1727
rect 152 1703 154 1726
rect 111 1702 115 1703
rect 111 1697 115 1698
rect 151 1702 155 1703
rect 151 1697 155 1698
rect 112 1677 114 1697
rect 184 1692 186 1726
rect 256 1703 258 1726
rect 360 1716 362 1782
rect 422 1768 428 1769
rect 422 1764 423 1768
rect 427 1764 428 1768
rect 422 1763 428 1764
rect 424 1759 426 1763
rect 423 1758 427 1759
rect 423 1753 427 1754
rect 463 1758 467 1759
rect 463 1753 467 1754
rect 462 1752 468 1753
rect 462 1748 463 1752
rect 467 1748 468 1752
rect 462 1747 468 1748
rect 500 1732 502 1798
rect 536 1790 538 1809
rect 632 1790 634 1809
rect 650 1807 651 1811
rect 655 1807 656 1811
rect 695 1809 699 1810
rect 719 1814 723 1815
rect 719 1809 723 1810
rect 759 1814 763 1815
rect 759 1809 763 1810
rect 799 1814 803 1815
rect 799 1809 803 1810
rect 831 1814 835 1815
rect 831 1809 835 1810
rect 879 1814 883 1815
rect 879 1809 883 1810
rect 903 1814 907 1815
rect 903 1809 907 1810
rect 959 1814 963 1815
rect 959 1809 963 1810
rect 975 1814 979 1815
rect 984 1812 986 1842
rect 1056 1815 1058 1842
rect 1062 1831 1068 1832
rect 1062 1827 1063 1831
rect 1067 1827 1068 1831
rect 1062 1826 1068 1827
rect 1039 1814 1043 1815
rect 975 1809 979 1810
rect 982 1811 988 1812
rect 650 1806 656 1807
rect 534 1789 540 1790
rect 534 1785 535 1789
rect 539 1785 540 1789
rect 534 1784 540 1785
rect 630 1789 636 1790
rect 630 1785 631 1789
rect 635 1785 636 1789
rect 652 1788 654 1806
rect 720 1790 722 1809
rect 800 1790 802 1809
rect 880 1790 882 1809
rect 960 1790 962 1809
rect 982 1807 983 1811
rect 987 1807 988 1811
rect 1039 1809 1043 1810
rect 1055 1814 1059 1815
rect 1055 1809 1059 1810
rect 982 1806 988 1807
rect 1040 1790 1042 1809
rect 718 1789 724 1790
rect 630 1784 636 1785
rect 650 1787 656 1788
rect 650 1783 651 1787
rect 655 1783 656 1787
rect 718 1785 719 1789
rect 723 1785 724 1789
rect 718 1784 724 1785
rect 798 1789 804 1790
rect 798 1785 799 1789
rect 803 1785 804 1789
rect 798 1784 804 1785
rect 878 1789 884 1790
rect 878 1785 879 1789
rect 883 1785 884 1789
rect 878 1784 884 1785
rect 958 1789 964 1790
rect 958 1785 959 1789
rect 963 1785 964 1789
rect 1038 1789 1044 1790
rect 958 1784 964 1785
rect 998 1787 1004 1788
rect 650 1782 656 1783
rect 998 1783 999 1787
rect 1003 1783 1004 1787
rect 1038 1785 1039 1789
rect 1043 1785 1044 1789
rect 1064 1788 1066 1826
rect 1288 1815 1290 1843
rect 1326 1840 1327 1844
rect 1331 1840 1332 1844
rect 1534 1841 1535 1845
rect 1539 1841 1540 1845
rect 1534 1840 1540 1841
rect 1606 1845 1612 1846
rect 1606 1841 1607 1845
rect 1611 1841 1612 1845
rect 1606 1840 1612 1841
rect 1686 1845 1692 1846
rect 1686 1841 1687 1845
rect 1691 1841 1692 1845
rect 1782 1845 1788 1846
rect 1686 1840 1692 1841
rect 1694 1843 1700 1844
rect 1326 1839 1332 1840
rect 1694 1839 1695 1843
rect 1699 1839 1700 1843
rect 1782 1841 1783 1845
rect 1787 1841 1788 1845
rect 1804 1844 1806 1862
rect 1880 1846 1882 1865
rect 1976 1860 1978 1890
rect 2032 1871 2034 1890
rect 2128 1871 2130 1890
rect 2216 1871 2218 1890
rect 2304 1871 2306 1890
rect 2320 1876 2322 1890
rect 2318 1875 2324 1876
rect 2318 1871 2319 1875
rect 2323 1871 2324 1875
rect 2392 1871 2394 1890
rect 2456 1871 2458 1890
rect 2464 1880 2466 1946
rect 2502 1935 2508 1936
rect 2502 1931 2503 1935
rect 2507 1931 2508 1935
rect 2502 1930 2508 1931
rect 2504 1923 2506 1930
rect 2503 1922 2507 1923
rect 2503 1917 2507 1918
rect 2504 1914 2506 1917
rect 2502 1913 2508 1914
rect 2502 1909 2503 1913
rect 2507 1909 2508 1913
rect 2502 1908 2508 1909
rect 2502 1896 2508 1897
rect 2486 1895 2492 1896
rect 2486 1891 2487 1895
rect 2491 1891 2492 1895
rect 2502 1892 2503 1896
rect 2507 1892 2508 1896
rect 2502 1891 2508 1892
rect 2486 1890 2492 1891
rect 2462 1879 2468 1880
rect 2462 1875 2463 1879
rect 2467 1875 2468 1879
rect 2462 1874 2468 1875
rect 2474 1871 2480 1872
rect 1983 1870 1987 1871
rect 1983 1865 1987 1866
rect 2031 1870 2035 1871
rect 2031 1865 2035 1866
rect 2079 1870 2083 1871
rect 2079 1865 2083 1866
rect 2127 1870 2131 1871
rect 2127 1865 2131 1866
rect 2175 1870 2179 1871
rect 2175 1865 2179 1866
rect 2215 1870 2219 1871
rect 2215 1865 2219 1866
rect 2271 1870 2275 1871
rect 2271 1865 2275 1866
rect 2303 1870 2307 1871
rect 2318 1870 2324 1871
rect 2367 1870 2371 1871
rect 2303 1865 2307 1866
rect 2367 1865 2371 1866
rect 2391 1870 2395 1871
rect 2391 1865 2395 1866
rect 2455 1870 2459 1871
rect 2474 1867 2475 1871
rect 2479 1867 2480 1871
rect 2474 1866 2480 1867
rect 2455 1865 2459 1866
rect 1974 1859 1980 1860
rect 1974 1855 1975 1859
rect 1979 1855 1980 1859
rect 1974 1854 1980 1855
rect 1984 1846 1986 1865
rect 2080 1846 2082 1865
rect 2166 1859 2172 1860
rect 2166 1855 2167 1859
rect 2171 1855 2172 1859
rect 2166 1854 2172 1855
rect 1878 1845 1884 1846
rect 1782 1840 1788 1841
rect 1802 1843 1808 1844
rect 1694 1838 1700 1839
rect 1802 1839 1803 1843
rect 1807 1839 1808 1843
rect 1878 1841 1879 1845
rect 1883 1841 1884 1845
rect 1878 1840 1884 1841
rect 1982 1845 1988 1846
rect 1982 1841 1983 1845
rect 1987 1841 1988 1845
rect 1982 1840 1988 1841
rect 2078 1845 2084 1846
rect 2078 1841 2079 1845
rect 2083 1841 2084 1845
rect 2078 1840 2084 1841
rect 1802 1838 1808 1839
rect 1326 1827 1332 1828
rect 1326 1823 1327 1827
rect 1331 1823 1332 1827
rect 1326 1822 1332 1823
rect 1518 1824 1524 1825
rect 1328 1815 1330 1822
rect 1518 1820 1519 1824
rect 1523 1820 1524 1824
rect 1518 1819 1524 1820
rect 1590 1824 1596 1825
rect 1590 1820 1591 1824
rect 1595 1820 1596 1824
rect 1590 1819 1596 1820
rect 1670 1824 1676 1825
rect 1670 1820 1671 1824
rect 1675 1820 1676 1824
rect 1670 1819 1676 1820
rect 1520 1815 1522 1819
rect 1592 1815 1594 1819
rect 1672 1815 1674 1819
rect 1119 1814 1123 1815
rect 1119 1809 1123 1810
rect 1287 1814 1291 1815
rect 1287 1809 1291 1810
rect 1327 1814 1331 1815
rect 1327 1809 1331 1810
rect 1463 1814 1467 1815
rect 1463 1809 1467 1810
rect 1519 1814 1523 1815
rect 1519 1809 1523 1810
rect 1559 1814 1563 1815
rect 1559 1809 1563 1810
rect 1591 1814 1595 1815
rect 1591 1809 1595 1810
rect 1663 1814 1667 1815
rect 1663 1809 1667 1810
rect 1671 1814 1675 1815
rect 1671 1809 1675 1810
rect 1120 1790 1122 1809
rect 1138 1803 1144 1804
rect 1138 1799 1139 1803
rect 1143 1799 1144 1803
rect 1138 1798 1144 1799
rect 1118 1789 1124 1790
rect 1038 1784 1044 1785
rect 1062 1787 1068 1788
rect 998 1782 1004 1783
rect 1062 1783 1063 1787
rect 1067 1783 1068 1787
rect 1118 1785 1119 1789
rect 1123 1785 1124 1789
rect 1118 1784 1124 1785
rect 1062 1782 1068 1783
rect 518 1768 524 1769
rect 518 1764 519 1768
rect 523 1764 524 1768
rect 518 1763 524 1764
rect 614 1768 620 1769
rect 614 1764 615 1768
rect 619 1764 620 1768
rect 614 1763 620 1764
rect 702 1768 708 1769
rect 702 1764 703 1768
rect 707 1764 708 1768
rect 702 1763 708 1764
rect 782 1768 788 1769
rect 782 1764 783 1768
rect 787 1764 788 1768
rect 782 1763 788 1764
rect 862 1768 868 1769
rect 862 1764 863 1768
rect 867 1764 868 1768
rect 862 1763 868 1764
rect 942 1768 948 1769
rect 942 1764 943 1768
rect 947 1764 948 1768
rect 942 1763 948 1764
rect 520 1759 522 1763
rect 616 1759 618 1763
rect 704 1759 706 1763
rect 784 1759 786 1763
rect 864 1759 866 1763
rect 944 1759 946 1763
rect 519 1758 523 1759
rect 519 1753 523 1754
rect 575 1758 579 1759
rect 575 1753 579 1754
rect 615 1758 619 1759
rect 615 1753 619 1754
rect 679 1758 683 1759
rect 679 1753 683 1754
rect 703 1758 707 1759
rect 703 1753 707 1754
rect 783 1758 787 1759
rect 783 1753 787 1754
rect 863 1758 867 1759
rect 863 1753 867 1754
rect 887 1758 891 1759
rect 887 1753 891 1754
rect 943 1758 947 1759
rect 943 1753 947 1754
rect 991 1758 995 1759
rect 991 1753 995 1754
rect 574 1752 580 1753
rect 574 1748 575 1752
rect 579 1748 580 1752
rect 574 1747 580 1748
rect 678 1752 684 1753
rect 678 1748 679 1752
rect 683 1748 684 1752
rect 678 1747 684 1748
rect 782 1752 788 1753
rect 782 1748 783 1752
rect 787 1748 788 1752
rect 782 1747 788 1748
rect 886 1752 892 1753
rect 886 1748 887 1752
rect 891 1748 892 1752
rect 886 1747 892 1748
rect 990 1752 996 1753
rect 990 1748 991 1752
rect 995 1748 996 1752
rect 990 1747 996 1748
rect 366 1731 372 1732
rect 366 1727 367 1731
rect 371 1727 372 1731
rect 366 1726 372 1727
rect 478 1731 484 1732
rect 478 1727 479 1731
rect 483 1727 484 1731
rect 478 1726 484 1727
rect 498 1731 504 1732
rect 498 1727 499 1731
rect 503 1727 504 1731
rect 498 1726 504 1727
rect 590 1731 596 1732
rect 590 1727 591 1731
rect 595 1727 596 1731
rect 590 1726 596 1727
rect 694 1731 700 1732
rect 694 1727 695 1731
rect 699 1727 700 1731
rect 694 1726 700 1727
rect 734 1731 740 1732
rect 734 1727 735 1731
rect 739 1727 740 1731
rect 734 1726 740 1727
rect 798 1731 804 1732
rect 798 1727 799 1731
rect 803 1727 804 1731
rect 798 1726 804 1727
rect 902 1731 908 1732
rect 902 1727 903 1731
rect 907 1727 908 1731
rect 902 1726 908 1727
rect 918 1731 924 1732
rect 918 1727 919 1731
rect 923 1727 924 1731
rect 918 1726 924 1727
rect 358 1715 364 1716
rect 358 1711 359 1715
rect 363 1711 364 1715
rect 358 1710 364 1711
rect 368 1703 370 1726
rect 480 1703 482 1726
rect 592 1703 594 1726
rect 658 1715 664 1716
rect 658 1711 659 1715
rect 663 1711 664 1715
rect 658 1710 664 1711
rect 191 1702 195 1703
rect 191 1697 195 1698
rect 255 1702 259 1703
rect 255 1697 259 1698
rect 271 1702 275 1703
rect 271 1697 275 1698
rect 351 1702 355 1703
rect 351 1697 355 1698
rect 367 1702 371 1703
rect 367 1697 371 1698
rect 439 1702 443 1703
rect 439 1697 443 1698
rect 479 1702 483 1703
rect 479 1697 483 1698
rect 535 1702 539 1703
rect 535 1697 539 1698
rect 591 1702 595 1703
rect 591 1697 595 1698
rect 639 1702 643 1703
rect 639 1697 643 1698
rect 182 1691 188 1692
rect 182 1687 183 1691
rect 187 1687 188 1691
rect 182 1686 188 1687
rect 192 1678 194 1697
rect 272 1678 274 1697
rect 352 1678 354 1697
rect 440 1678 442 1697
rect 446 1691 452 1692
rect 446 1687 447 1691
rect 451 1687 452 1691
rect 446 1686 452 1687
rect 190 1677 196 1678
rect 110 1676 116 1677
rect 110 1672 111 1676
rect 115 1672 116 1676
rect 190 1673 191 1677
rect 195 1673 196 1677
rect 190 1672 196 1673
rect 270 1677 276 1678
rect 270 1673 271 1677
rect 275 1673 276 1677
rect 270 1672 276 1673
rect 350 1677 356 1678
rect 350 1673 351 1677
rect 355 1673 356 1677
rect 438 1677 444 1678
rect 350 1672 356 1673
rect 358 1675 364 1676
rect 110 1671 116 1672
rect 358 1671 359 1675
rect 363 1671 364 1675
rect 438 1673 439 1677
rect 443 1673 444 1677
rect 438 1672 444 1673
rect 358 1670 364 1671
rect 110 1659 116 1660
rect 110 1655 111 1659
rect 115 1655 116 1659
rect 110 1654 116 1655
rect 174 1656 180 1657
rect 112 1651 114 1654
rect 174 1652 175 1656
rect 179 1652 180 1656
rect 174 1651 180 1652
rect 254 1656 260 1657
rect 254 1652 255 1656
rect 259 1652 260 1656
rect 254 1651 260 1652
rect 334 1656 340 1657
rect 334 1652 335 1656
rect 339 1652 340 1656
rect 334 1651 340 1652
rect 111 1650 115 1651
rect 111 1645 115 1646
rect 175 1650 179 1651
rect 175 1645 179 1646
rect 215 1650 219 1651
rect 215 1645 219 1646
rect 255 1650 259 1651
rect 255 1645 259 1646
rect 271 1650 275 1651
rect 271 1645 275 1646
rect 335 1650 339 1651
rect 335 1645 339 1646
rect 112 1642 114 1645
rect 214 1644 220 1645
rect 110 1641 116 1642
rect 110 1637 111 1641
rect 115 1637 116 1641
rect 214 1640 215 1644
rect 219 1640 220 1644
rect 214 1639 220 1640
rect 270 1644 276 1645
rect 270 1640 271 1644
rect 275 1640 276 1644
rect 270 1639 276 1640
rect 334 1644 340 1645
rect 334 1640 335 1644
rect 339 1640 340 1644
rect 334 1639 340 1640
rect 110 1636 116 1637
rect 110 1624 116 1625
rect 110 1620 111 1624
rect 115 1620 116 1624
rect 110 1619 116 1620
rect 230 1623 236 1624
rect 230 1619 231 1623
rect 235 1619 236 1623
rect 112 1599 114 1619
rect 230 1618 236 1619
rect 286 1623 292 1624
rect 286 1619 287 1623
rect 291 1619 292 1623
rect 286 1618 292 1619
rect 294 1623 300 1624
rect 294 1619 295 1623
rect 299 1619 300 1623
rect 294 1618 300 1619
rect 350 1623 356 1624
rect 350 1619 351 1623
rect 355 1619 356 1623
rect 350 1618 356 1619
rect 232 1599 234 1618
rect 288 1599 290 1618
rect 111 1598 115 1599
rect 111 1593 115 1594
rect 231 1598 235 1599
rect 231 1593 235 1594
rect 287 1598 291 1599
rect 287 1593 291 1594
rect 112 1573 114 1593
rect 288 1574 290 1593
rect 296 1588 298 1618
rect 352 1599 354 1618
rect 360 1608 362 1670
rect 422 1656 428 1657
rect 422 1652 423 1656
rect 427 1652 428 1656
rect 422 1651 428 1652
rect 407 1650 411 1651
rect 407 1645 411 1646
rect 423 1650 427 1651
rect 423 1645 427 1646
rect 406 1644 412 1645
rect 406 1640 407 1644
rect 411 1640 412 1644
rect 406 1639 412 1640
rect 448 1624 450 1686
rect 536 1678 538 1697
rect 640 1678 642 1697
rect 534 1677 540 1678
rect 534 1673 535 1677
rect 539 1673 540 1677
rect 534 1672 540 1673
rect 638 1677 644 1678
rect 638 1673 639 1677
rect 643 1673 644 1677
rect 660 1676 662 1710
rect 696 1703 698 1726
rect 695 1702 699 1703
rect 695 1697 699 1698
rect 736 1692 738 1726
rect 800 1703 802 1726
rect 904 1703 906 1726
rect 920 1712 922 1726
rect 1000 1716 1002 1782
rect 1022 1768 1028 1769
rect 1022 1764 1023 1768
rect 1027 1764 1028 1768
rect 1022 1763 1028 1764
rect 1102 1768 1108 1769
rect 1102 1764 1103 1768
rect 1107 1764 1108 1768
rect 1102 1763 1108 1764
rect 1024 1759 1026 1763
rect 1104 1759 1106 1763
rect 1023 1758 1027 1759
rect 1023 1753 1027 1754
rect 1103 1758 1107 1759
rect 1103 1753 1107 1754
rect 1102 1752 1108 1753
rect 1102 1748 1103 1752
rect 1107 1748 1108 1752
rect 1102 1747 1108 1748
rect 1140 1732 1142 1798
rect 1288 1789 1290 1809
rect 1328 1806 1330 1809
rect 1462 1808 1468 1809
rect 1326 1805 1332 1806
rect 1326 1801 1327 1805
rect 1331 1801 1332 1805
rect 1462 1804 1463 1808
rect 1467 1804 1468 1808
rect 1462 1803 1468 1804
rect 1558 1808 1564 1809
rect 1558 1804 1559 1808
rect 1563 1804 1564 1808
rect 1558 1803 1564 1804
rect 1662 1808 1668 1809
rect 1662 1804 1663 1808
rect 1667 1804 1668 1808
rect 1662 1803 1668 1804
rect 1326 1800 1332 1801
rect 1286 1788 1292 1789
rect 1286 1784 1287 1788
rect 1291 1784 1292 1788
rect 1286 1783 1292 1784
rect 1326 1788 1332 1789
rect 1326 1784 1327 1788
rect 1331 1784 1332 1788
rect 1326 1783 1332 1784
rect 1478 1787 1484 1788
rect 1478 1783 1479 1787
rect 1483 1783 1484 1787
rect 1286 1771 1292 1772
rect 1286 1767 1287 1771
rect 1291 1767 1292 1771
rect 1286 1766 1292 1767
rect 1288 1759 1290 1766
rect 1328 1759 1330 1783
rect 1478 1782 1484 1783
rect 1558 1787 1564 1788
rect 1558 1783 1559 1787
rect 1563 1783 1564 1787
rect 1558 1782 1564 1783
rect 1574 1787 1580 1788
rect 1574 1783 1575 1787
rect 1579 1783 1580 1787
rect 1574 1782 1580 1783
rect 1678 1787 1684 1788
rect 1678 1783 1679 1787
rect 1683 1783 1684 1787
rect 1678 1782 1684 1783
rect 1480 1759 1482 1782
rect 1287 1758 1291 1759
rect 1287 1753 1291 1754
rect 1327 1758 1331 1759
rect 1327 1753 1331 1754
rect 1375 1758 1379 1759
rect 1375 1753 1379 1754
rect 1471 1758 1475 1759
rect 1471 1753 1475 1754
rect 1479 1758 1483 1759
rect 1479 1753 1483 1754
rect 1288 1750 1290 1753
rect 1286 1749 1292 1750
rect 1286 1745 1287 1749
rect 1291 1745 1292 1749
rect 1286 1744 1292 1745
rect 1328 1733 1330 1753
rect 1376 1734 1378 1753
rect 1472 1734 1474 1753
rect 1560 1748 1562 1782
rect 1576 1759 1578 1782
rect 1680 1759 1682 1782
rect 1696 1772 1698 1838
rect 1766 1824 1772 1825
rect 1766 1820 1767 1824
rect 1771 1820 1772 1824
rect 1766 1819 1772 1820
rect 1862 1824 1868 1825
rect 1862 1820 1863 1824
rect 1867 1820 1868 1824
rect 1862 1819 1868 1820
rect 1966 1824 1972 1825
rect 1966 1820 1967 1824
rect 1971 1820 1972 1824
rect 1966 1819 1972 1820
rect 2062 1824 2068 1825
rect 2062 1820 2063 1824
rect 2067 1820 2068 1824
rect 2062 1819 2068 1820
rect 2158 1824 2164 1825
rect 2158 1820 2159 1824
rect 2163 1820 2164 1824
rect 2158 1819 2164 1820
rect 1768 1815 1770 1819
rect 1864 1815 1866 1819
rect 1968 1815 1970 1819
rect 2064 1815 2066 1819
rect 2160 1815 2162 1819
rect 1767 1814 1771 1815
rect 1767 1809 1771 1810
rect 1863 1814 1867 1815
rect 1863 1809 1867 1810
rect 1879 1814 1883 1815
rect 1879 1809 1883 1810
rect 1967 1814 1971 1815
rect 1967 1809 1971 1810
rect 1983 1814 1987 1815
rect 1983 1809 1987 1810
rect 2063 1814 2067 1815
rect 2063 1809 2067 1810
rect 2087 1814 2091 1815
rect 2087 1809 2091 1810
rect 2159 1814 2163 1815
rect 2159 1809 2163 1810
rect 1766 1808 1772 1809
rect 1766 1804 1767 1808
rect 1771 1804 1772 1808
rect 1766 1803 1772 1804
rect 1878 1808 1884 1809
rect 1878 1804 1879 1808
rect 1883 1804 1884 1808
rect 1878 1803 1884 1804
rect 1982 1808 1988 1809
rect 1982 1804 1983 1808
rect 1987 1804 1988 1808
rect 1982 1803 1988 1804
rect 2086 1808 2092 1809
rect 2086 1804 2087 1808
rect 2091 1804 2092 1808
rect 2086 1803 2092 1804
rect 2168 1797 2170 1854
rect 2176 1846 2178 1865
rect 2272 1846 2274 1865
rect 2368 1846 2370 1865
rect 2456 1846 2458 1865
rect 2174 1845 2180 1846
rect 2174 1841 2175 1845
rect 2179 1841 2180 1845
rect 2174 1840 2180 1841
rect 2270 1845 2276 1846
rect 2270 1841 2271 1845
rect 2275 1841 2276 1845
rect 2270 1840 2276 1841
rect 2366 1845 2372 1846
rect 2366 1841 2367 1845
rect 2371 1841 2372 1845
rect 2366 1840 2372 1841
rect 2454 1845 2460 1846
rect 2454 1841 2455 1845
rect 2459 1841 2460 1845
rect 2476 1844 2478 1866
rect 2454 1840 2460 1841
rect 2474 1843 2480 1844
rect 2474 1839 2475 1843
rect 2479 1839 2480 1843
rect 2474 1838 2480 1839
rect 2254 1824 2260 1825
rect 2254 1820 2255 1824
rect 2259 1820 2260 1824
rect 2254 1819 2260 1820
rect 2350 1824 2356 1825
rect 2350 1820 2351 1824
rect 2355 1820 2356 1824
rect 2350 1819 2356 1820
rect 2438 1824 2444 1825
rect 2438 1820 2439 1824
rect 2443 1820 2444 1824
rect 2438 1819 2444 1820
rect 2256 1815 2258 1819
rect 2352 1815 2354 1819
rect 2440 1815 2442 1819
rect 2183 1814 2187 1815
rect 2183 1809 2187 1810
rect 2255 1814 2259 1815
rect 2255 1809 2259 1810
rect 2271 1814 2275 1815
rect 2271 1809 2275 1810
rect 2351 1814 2355 1815
rect 2351 1809 2355 1810
rect 2367 1814 2371 1815
rect 2367 1809 2371 1810
rect 2439 1814 2443 1815
rect 2439 1809 2443 1810
rect 2182 1808 2188 1809
rect 2182 1804 2183 1808
rect 2187 1804 2188 1808
rect 2182 1803 2188 1804
rect 2270 1808 2276 1809
rect 2270 1804 2271 1808
rect 2275 1804 2276 1808
rect 2270 1803 2276 1804
rect 2366 1808 2372 1809
rect 2366 1804 2367 1808
rect 2371 1804 2372 1808
rect 2366 1803 2372 1804
rect 2438 1808 2444 1809
rect 2438 1804 2439 1808
rect 2443 1804 2444 1808
rect 2438 1803 2444 1804
rect 2167 1796 2171 1797
rect 2167 1791 2171 1792
rect 2403 1796 2407 1797
rect 2403 1791 2407 1792
rect 2404 1788 2406 1791
rect 1782 1787 1788 1788
rect 1782 1783 1783 1787
rect 1787 1783 1788 1787
rect 1782 1782 1788 1783
rect 1894 1787 1900 1788
rect 1894 1783 1895 1787
rect 1899 1783 1900 1787
rect 1894 1782 1900 1783
rect 1902 1787 1908 1788
rect 1902 1783 1903 1787
rect 1907 1783 1908 1787
rect 1902 1782 1908 1783
rect 1998 1787 2004 1788
rect 1998 1783 1999 1787
rect 2003 1783 2004 1787
rect 1998 1782 2004 1783
rect 2102 1787 2108 1788
rect 2102 1783 2103 1787
rect 2107 1783 2108 1787
rect 2102 1782 2108 1783
rect 2198 1787 2204 1788
rect 2198 1783 2199 1787
rect 2203 1783 2204 1787
rect 2198 1782 2204 1783
rect 2286 1787 2292 1788
rect 2286 1783 2287 1787
rect 2291 1783 2292 1787
rect 2286 1782 2292 1783
rect 2382 1787 2388 1788
rect 2382 1783 2383 1787
rect 2387 1783 2388 1787
rect 2382 1782 2388 1783
rect 2402 1787 2408 1788
rect 2402 1783 2403 1787
rect 2407 1783 2408 1787
rect 2402 1782 2408 1783
rect 2454 1787 2460 1788
rect 2454 1783 2455 1787
rect 2459 1783 2460 1787
rect 2454 1782 2460 1783
rect 2462 1787 2468 1788
rect 2462 1783 2463 1787
rect 2467 1783 2468 1787
rect 2462 1782 2468 1783
rect 1694 1771 1700 1772
rect 1694 1767 1695 1771
rect 1699 1767 1700 1771
rect 1694 1766 1700 1767
rect 1784 1759 1786 1782
rect 1896 1759 1898 1782
rect 1904 1764 1906 1782
rect 1902 1763 1908 1764
rect 1902 1759 1903 1763
rect 1907 1759 1908 1763
rect 2000 1759 2002 1782
rect 2104 1759 2106 1782
rect 2200 1759 2202 1782
rect 2288 1759 2290 1782
rect 2370 1767 2376 1768
rect 2370 1763 2371 1767
rect 2375 1763 2376 1767
rect 2370 1762 2376 1763
rect 1567 1758 1571 1759
rect 1567 1753 1571 1754
rect 1575 1758 1579 1759
rect 1575 1753 1579 1754
rect 1671 1758 1675 1759
rect 1671 1753 1675 1754
rect 1679 1758 1683 1759
rect 1679 1753 1683 1754
rect 1775 1758 1779 1759
rect 1775 1753 1779 1754
rect 1783 1758 1787 1759
rect 1887 1758 1891 1759
rect 1783 1753 1787 1754
rect 1794 1755 1800 1756
rect 1558 1747 1564 1748
rect 1558 1743 1559 1747
rect 1563 1743 1564 1747
rect 1558 1742 1564 1743
rect 1568 1734 1570 1753
rect 1672 1734 1674 1753
rect 1776 1734 1778 1753
rect 1794 1751 1795 1755
rect 1799 1751 1800 1755
rect 1887 1753 1891 1754
rect 1895 1758 1899 1759
rect 1902 1758 1908 1759
rect 1999 1758 2003 1759
rect 1895 1753 1899 1754
rect 1999 1753 2003 1754
rect 2103 1758 2107 1759
rect 2103 1753 2107 1754
rect 2111 1758 2115 1759
rect 2111 1753 2115 1754
rect 2199 1758 2203 1759
rect 2199 1753 2203 1754
rect 2231 1758 2235 1759
rect 2231 1753 2235 1754
rect 2287 1758 2291 1759
rect 2351 1758 2355 1759
rect 2287 1753 2291 1754
rect 2342 1755 2348 1756
rect 1794 1750 1800 1751
rect 1374 1733 1380 1734
rect 1286 1732 1292 1733
rect 1006 1731 1012 1732
rect 1006 1727 1007 1731
rect 1011 1727 1012 1731
rect 1006 1726 1012 1727
rect 1118 1731 1124 1732
rect 1118 1727 1119 1731
rect 1123 1727 1124 1731
rect 1118 1726 1124 1727
rect 1138 1731 1144 1732
rect 1138 1727 1139 1731
rect 1143 1727 1144 1731
rect 1286 1728 1287 1732
rect 1291 1728 1292 1732
rect 1286 1727 1292 1728
rect 1326 1732 1332 1733
rect 1326 1728 1327 1732
rect 1331 1728 1332 1732
rect 1374 1729 1375 1733
rect 1379 1729 1380 1733
rect 1470 1733 1476 1734
rect 1374 1728 1380 1729
rect 1438 1731 1444 1732
rect 1326 1727 1332 1728
rect 1438 1727 1439 1731
rect 1443 1727 1444 1731
rect 1470 1729 1471 1733
rect 1475 1729 1476 1733
rect 1470 1728 1476 1729
rect 1566 1733 1572 1734
rect 1566 1729 1567 1733
rect 1571 1729 1572 1733
rect 1566 1728 1572 1729
rect 1670 1733 1676 1734
rect 1670 1729 1671 1733
rect 1675 1729 1676 1733
rect 1670 1728 1676 1729
rect 1774 1733 1780 1734
rect 1774 1729 1775 1733
rect 1779 1729 1780 1733
rect 1796 1732 1798 1750
rect 1888 1734 1890 1753
rect 2000 1734 2002 1753
rect 2112 1734 2114 1753
rect 2232 1734 2234 1753
rect 2342 1751 2343 1755
rect 2347 1751 2348 1755
rect 2351 1753 2355 1754
rect 2342 1750 2348 1751
rect 1886 1733 1892 1734
rect 1774 1728 1780 1729
rect 1794 1731 1800 1732
rect 1138 1726 1144 1727
rect 998 1715 1004 1716
rect 918 1711 924 1712
rect 918 1707 919 1711
rect 923 1707 924 1711
rect 998 1711 999 1715
rect 1003 1711 1004 1715
rect 998 1710 1004 1711
rect 918 1706 924 1707
rect 1008 1703 1010 1726
rect 1120 1703 1122 1726
rect 1194 1715 1200 1716
rect 1194 1711 1195 1715
rect 1199 1711 1200 1715
rect 1194 1710 1200 1711
rect 743 1702 747 1703
rect 743 1697 747 1698
rect 799 1702 803 1703
rect 799 1697 803 1698
rect 847 1702 851 1703
rect 847 1697 851 1698
rect 903 1702 907 1703
rect 903 1697 907 1698
rect 951 1702 955 1703
rect 951 1697 955 1698
rect 1007 1702 1011 1703
rect 1007 1697 1011 1698
rect 1063 1702 1067 1703
rect 1063 1697 1067 1698
rect 1119 1702 1123 1703
rect 1119 1697 1123 1698
rect 1175 1702 1179 1703
rect 1175 1697 1179 1698
rect 734 1691 740 1692
rect 734 1687 735 1691
rect 739 1687 740 1691
rect 734 1686 740 1687
rect 744 1678 746 1697
rect 848 1678 850 1697
rect 952 1678 954 1697
rect 1064 1678 1066 1697
rect 1090 1691 1096 1692
rect 1090 1687 1091 1691
rect 1095 1687 1096 1691
rect 1090 1686 1096 1687
rect 742 1677 748 1678
rect 638 1672 644 1673
rect 658 1675 664 1676
rect 658 1671 659 1675
rect 663 1671 664 1675
rect 742 1673 743 1677
rect 747 1673 748 1677
rect 742 1672 748 1673
rect 846 1677 852 1678
rect 846 1673 847 1677
rect 851 1673 852 1677
rect 846 1672 852 1673
rect 950 1677 956 1678
rect 950 1673 951 1677
rect 955 1673 956 1677
rect 1062 1677 1068 1678
rect 950 1672 956 1673
rect 966 1675 972 1676
rect 658 1670 664 1671
rect 966 1671 967 1675
rect 971 1671 972 1675
rect 1062 1673 1063 1677
rect 1067 1673 1068 1677
rect 1062 1672 1068 1673
rect 966 1670 972 1671
rect 518 1656 524 1657
rect 518 1652 519 1656
rect 523 1652 524 1656
rect 518 1651 524 1652
rect 622 1656 628 1657
rect 622 1652 623 1656
rect 627 1652 628 1656
rect 622 1651 628 1652
rect 726 1656 732 1657
rect 726 1652 727 1656
rect 731 1652 732 1656
rect 726 1651 732 1652
rect 830 1656 836 1657
rect 830 1652 831 1656
rect 835 1652 836 1656
rect 830 1651 836 1652
rect 934 1656 940 1657
rect 934 1652 935 1656
rect 939 1652 940 1656
rect 934 1651 940 1652
rect 479 1650 483 1651
rect 479 1645 483 1646
rect 519 1650 523 1651
rect 519 1645 523 1646
rect 559 1650 563 1651
rect 559 1645 563 1646
rect 623 1650 627 1651
rect 623 1645 627 1646
rect 647 1650 651 1651
rect 647 1645 651 1646
rect 727 1650 731 1651
rect 727 1645 731 1646
rect 743 1650 747 1651
rect 743 1645 747 1646
rect 831 1650 835 1651
rect 831 1645 835 1646
rect 839 1650 843 1651
rect 839 1645 843 1646
rect 935 1650 939 1651
rect 935 1645 939 1646
rect 943 1650 947 1651
rect 943 1645 947 1646
rect 478 1644 484 1645
rect 478 1640 479 1644
rect 483 1640 484 1644
rect 478 1639 484 1640
rect 558 1644 564 1645
rect 558 1640 559 1644
rect 563 1640 564 1644
rect 558 1639 564 1640
rect 646 1644 652 1645
rect 646 1640 647 1644
rect 651 1640 652 1644
rect 646 1639 652 1640
rect 742 1644 748 1645
rect 742 1640 743 1644
rect 747 1640 748 1644
rect 742 1639 748 1640
rect 838 1644 844 1645
rect 838 1640 839 1644
rect 843 1640 844 1644
rect 838 1639 844 1640
rect 942 1644 948 1645
rect 942 1640 943 1644
rect 947 1640 948 1644
rect 942 1639 948 1640
rect 422 1623 428 1624
rect 422 1619 423 1623
rect 427 1619 428 1623
rect 422 1618 428 1619
rect 446 1623 452 1624
rect 446 1619 447 1623
rect 451 1619 452 1623
rect 446 1618 452 1619
rect 494 1623 500 1624
rect 494 1619 495 1623
rect 499 1619 500 1623
rect 494 1618 500 1619
rect 574 1623 580 1624
rect 574 1619 575 1623
rect 579 1619 580 1623
rect 574 1618 580 1619
rect 662 1623 668 1624
rect 662 1619 663 1623
rect 667 1619 668 1623
rect 662 1618 668 1619
rect 758 1623 764 1624
rect 758 1619 759 1623
rect 763 1619 764 1623
rect 758 1618 764 1619
rect 806 1623 812 1624
rect 806 1619 807 1623
rect 811 1619 812 1623
rect 806 1618 812 1619
rect 854 1623 860 1624
rect 854 1619 855 1623
rect 859 1619 860 1623
rect 854 1618 860 1619
rect 870 1623 876 1624
rect 870 1619 871 1623
rect 875 1619 876 1623
rect 870 1618 876 1619
rect 958 1623 964 1624
rect 958 1619 959 1623
rect 963 1619 964 1623
rect 958 1618 964 1619
rect 358 1607 364 1608
rect 358 1603 359 1607
rect 363 1603 364 1607
rect 358 1602 364 1603
rect 424 1599 426 1618
rect 496 1599 498 1618
rect 526 1607 532 1608
rect 526 1603 527 1607
rect 531 1603 532 1607
rect 526 1602 532 1603
rect 351 1598 355 1599
rect 351 1593 355 1594
rect 423 1598 427 1599
rect 423 1593 427 1594
rect 495 1598 499 1599
rect 495 1593 499 1594
rect 503 1598 507 1599
rect 503 1593 507 1594
rect 294 1587 300 1588
rect 294 1583 295 1587
rect 299 1583 300 1587
rect 294 1582 300 1583
rect 352 1574 354 1593
rect 424 1574 426 1593
rect 504 1574 506 1593
rect 286 1573 292 1574
rect 110 1572 116 1573
rect 110 1568 111 1572
rect 115 1568 116 1572
rect 286 1569 287 1573
rect 291 1569 292 1573
rect 286 1568 292 1569
rect 350 1573 356 1574
rect 350 1569 351 1573
rect 355 1569 356 1573
rect 350 1568 356 1569
rect 422 1573 428 1574
rect 422 1569 423 1573
rect 427 1569 428 1573
rect 422 1568 428 1569
rect 502 1573 508 1574
rect 502 1569 503 1573
rect 507 1569 508 1573
rect 528 1572 530 1602
rect 576 1599 578 1618
rect 664 1599 666 1618
rect 760 1599 762 1618
rect 575 1598 579 1599
rect 575 1593 579 1594
rect 599 1598 603 1599
rect 599 1593 603 1594
rect 663 1598 667 1599
rect 663 1593 667 1594
rect 703 1598 707 1599
rect 703 1593 707 1594
rect 759 1598 763 1599
rect 759 1593 763 1594
rect 600 1574 602 1593
rect 618 1587 624 1588
rect 618 1583 619 1587
rect 623 1583 624 1587
rect 618 1582 624 1583
rect 598 1573 604 1574
rect 620 1573 622 1582
rect 704 1574 706 1593
rect 808 1588 810 1618
rect 856 1599 858 1618
rect 872 1604 874 1618
rect 870 1603 876 1604
rect 870 1599 871 1603
rect 875 1599 876 1603
rect 960 1599 962 1618
rect 968 1608 970 1670
rect 1046 1656 1052 1657
rect 1046 1652 1047 1656
rect 1051 1652 1052 1656
rect 1046 1651 1052 1652
rect 1047 1650 1051 1651
rect 1047 1645 1051 1646
rect 1055 1650 1059 1651
rect 1055 1645 1059 1646
rect 1054 1644 1060 1645
rect 1054 1640 1055 1644
rect 1059 1640 1060 1644
rect 1054 1639 1060 1640
rect 1092 1624 1094 1686
rect 1176 1678 1178 1697
rect 1174 1677 1180 1678
rect 1174 1673 1175 1677
rect 1179 1673 1180 1677
rect 1196 1676 1198 1710
rect 1288 1703 1290 1727
rect 1438 1726 1444 1727
rect 1794 1727 1795 1731
rect 1799 1727 1800 1731
rect 1886 1729 1887 1733
rect 1891 1729 1892 1733
rect 1886 1728 1892 1729
rect 1998 1733 2004 1734
rect 1998 1729 1999 1733
rect 2003 1729 2004 1733
rect 1998 1728 2004 1729
rect 2110 1733 2116 1734
rect 2110 1729 2111 1733
rect 2115 1729 2116 1733
rect 2110 1728 2116 1729
rect 2230 1733 2236 1734
rect 2230 1729 2231 1733
rect 2235 1729 2236 1733
rect 2230 1728 2236 1729
rect 1794 1726 1800 1727
rect 1326 1715 1332 1716
rect 1326 1711 1327 1715
rect 1331 1711 1332 1715
rect 1326 1710 1332 1711
rect 1358 1712 1364 1713
rect 1328 1707 1330 1710
rect 1358 1708 1359 1712
rect 1363 1708 1364 1712
rect 1358 1707 1364 1708
rect 1327 1706 1331 1707
rect 1287 1702 1291 1703
rect 1327 1701 1331 1702
rect 1351 1706 1355 1707
rect 1351 1701 1355 1702
rect 1359 1706 1363 1707
rect 1359 1701 1363 1702
rect 1431 1706 1435 1707
rect 1431 1701 1435 1702
rect 1328 1698 1330 1701
rect 1350 1700 1356 1701
rect 1287 1697 1291 1698
rect 1326 1697 1332 1698
rect 1288 1677 1290 1697
rect 1326 1693 1327 1697
rect 1331 1693 1332 1697
rect 1350 1696 1351 1700
rect 1355 1696 1356 1700
rect 1350 1695 1356 1696
rect 1430 1700 1436 1701
rect 1430 1696 1431 1700
rect 1435 1696 1436 1700
rect 1430 1695 1436 1696
rect 1326 1692 1332 1693
rect 1326 1680 1332 1681
rect 1286 1676 1292 1677
rect 1174 1672 1180 1673
rect 1194 1675 1200 1676
rect 1194 1671 1195 1675
rect 1199 1671 1200 1675
rect 1286 1672 1287 1676
rect 1291 1672 1292 1676
rect 1326 1676 1327 1680
rect 1331 1676 1332 1680
rect 1326 1675 1332 1676
rect 1366 1679 1372 1680
rect 1366 1675 1367 1679
rect 1371 1675 1372 1679
rect 1286 1671 1292 1672
rect 1194 1670 1200 1671
rect 1286 1659 1292 1660
rect 1158 1656 1164 1657
rect 1158 1652 1159 1656
rect 1163 1652 1164 1656
rect 1286 1655 1287 1659
rect 1291 1655 1292 1659
rect 1286 1654 1292 1655
rect 1158 1651 1164 1652
rect 1288 1651 1290 1654
rect 1159 1650 1163 1651
rect 1159 1645 1163 1646
rect 1175 1650 1179 1651
rect 1175 1645 1179 1646
rect 1287 1650 1291 1651
rect 1328 1647 1330 1675
rect 1366 1674 1372 1675
rect 1374 1679 1380 1680
rect 1374 1675 1375 1679
rect 1379 1675 1380 1679
rect 1374 1674 1380 1675
rect 1368 1647 1370 1674
rect 1287 1645 1291 1646
rect 1327 1646 1331 1647
rect 1174 1644 1180 1645
rect 1174 1640 1175 1644
rect 1179 1640 1180 1644
rect 1288 1642 1290 1645
rect 1174 1639 1180 1640
rect 1286 1641 1292 1642
rect 1327 1641 1331 1642
rect 1367 1646 1371 1647
rect 1367 1641 1371 1642
rect 1286 1637 1287 1641
rect 1291 1637 1292 1641
rect 1286 1636 1292 1637
rect 1286 1624 1292 1625
rect 1070 1623 1076 1624
rect 1070 1619 1071 1623
rect 1075 1619 1076 1623
rect 1070 1618 1076 1619
rect 1090 1623 1096 1624
rect 1090 1619 1091 1623
rect 1095 1619 1096 1623
rect 1090 1618 1096 1619
rect 1190 1623 1196 1624
rect 1190 1619 1191 1623
rect 1195 1619 1196 1623
rect 1286 1620 1287 1624
rect 1291 1620 1292 1624
rect 1328 1621 1330 1641
rect 1368 1622 1370 1641
rect 1376 1636 1378 1674
rect 1383 1668 1387 1669
rect 1440 1664 1442 1726
rect 1454 1712 1460 1713
rect 1454 1708 1455 1712
rect 1459 1708 1460 1712
rect 1454 1707 1460 1708
rect 1550 1712 1556 1713
rect 1550 1708 1551 1712
rect 1555 1708 1556 1712
rect 1550 1707 1556 1708
rect 1654 1712 1660 1713
rect 1654 1708 1655 1712
rect 1659 1708 1660 1712
rect 1654 1707 1660 1708
rect 1758 1712 1764 1713
rect 1758 1708 1759 1712
rect 1763 1708 1764 1712
rect 1758 1707 1764 1708
rect 1870 1712 1876 1713
rect 1870 1708 1871 1712
rect 1875 1708 1876 1712
rect 1870 1707 1876 1708
rect 1982 1712 1988 1713
rect 1982 1708 1983 1712
rect 1987 1708 1988 1712
rect 1982 1707 1988 1708
rect 2094 1712 2100 1713
rect 2094 1708 2095 1712
rect 2099 1708 2100 1712
rect 2094 1707 2100 1708
rect 2214 1712 2220 1713
rect 2214 1708 2215 1712
rect 2219 1708 2220 1712
rect 2214 1707 2220 1708
rect 2334 1712 2340 1713
rect 2334 1708 2335 1712
rect 2339 1708 2340 1712
rect 2334 1707 2340 1708
rect 1455 1706 1459 1707
rect 1455 1701 1459 1702
rect 1535 1706 1539 1707
rect 1535 1701 1539 1702
rect 1551 1706 1555 1707
rect 1551 1701 1555 1702
rect 1647 1706 1651 1707
rect 1647 1701 1651 1702
rect 1655 1706 1659 1707
rect 1655 1701 1659 1702
rect 1759 1706 1763 1707
rect 1759 1701 1763 1702
rect 1871 1706 1875 1707
rect 1871 1701 1875 1702
rect 1879 1706 1883 1707
rect 1879 1701 1883 1702
rect 1983 1706 1987 1707
rect 1983 1701 1987 1702
rect 2015 1706 2019 1707
rect 2015 1701 2019 1702
rect 2095 1706 2099 1707
rect 2095 1701 2099 1702
rect 2159 1706 2163 1707
rect 2159 1701 2163 1702
rect 2215 1706 2219 1707
rect 2215 1701 2219 1702
rect 2311 1706 2315 1707
rect 2311 1701 2315 1702
rect 2335 1706 2339 1707
rect 2335 1701 2339 1702
rect 1534 1700 1540 1701
rect 1534 1696 1535 1700
rect 1539 1696 1540 1700
rect 1534 1695 1540 1696
rect 1646 1700 1652 1701
rect 1646 1696 1647 1700
rect 1651 1696 1652 1700
rect 1646 1695 1652 1696
rect 1758 1700 1764 1701
rect 1758 1696 1759 1700
rect 1763 1696 1764 1700
rect 1758 1695 1764 1696
rect 1878 1700 1884 1701
rect 1878 1696 1879 1700
rect 1883 1696 1884 1700
rect 1878 1695 1884 1696
rect 2014 1700 2020 1701
rect 2014 1696 2015 1700
rect 2019 1696 2020 1700
rect 2014 1695 2020 1696
rect 2158 1700 2164 1701
rect 2158 1696 2159 1700
rect 2163 1696 2164 1700
rect 2158 1695 2164 1696
rect 2310 1700 2316 1701
rect 2310 1696 2311 1700
rect 2315 1696 2316 1700
rect 2310 1695 2316 1696
rect 2344 1680 2346 1750
rect 2352 1734 2354 1753
rect 2350 1733 2356 1734
rect 2350 1729 2351 1733
rect 2355 1729 2356 1733
rect 2372 1732 2374 1762
rect 2384 1759 2386 1782
rect 2456 1759 2458 1782
rect 2383 1758 2387 1759
rect 2383 1753 2387 1754
rect 2455 1758 2459 1759
rect 2455 1753 2459 1754
rect 2456 1734 2458 1753
rect 2464 1748 2466 1782
rect 2488 1772 2490 1890
rect 2504 1871 2506 1891
rect 2503 1870 2507 1871
rect 2503 1865 2507 1866
rect 2504 1845 2506 1865
rect 2502 1844 2508 1845
rect 2502 1840 2503 1844
rect 2507 1840 2508 1844
rect 2502 1839 2508 1840
rect 2502 1827 2508 1828
rect 2502 1823 2503 1827
rect 2507 1823 2508 1827
rect 2502 1822 2508 1823
rect 2504 1815 2506 1822
rect 2503 1814 2507 1815
rect 2503 1809 2507 1810
rect 2504 1806 2506 1809
rect 2502 1805 2508 1806
rect 2502 1801 2503 1805
rect 2507 1801 2508 1805
rect 2502 1800 2508 1801
rect 2502 1788 2508 1789
rect 2502 1784 2503 1788
rect 2507 1784 2508 1788
rect 2502 1783 2508 1784
rect 2486 1771 2492 1772
rect 2486 1767 2487 1771
rect 2491 1767 2492 1771
rect 2486 1766 2492 1767
rect 2504 1759 2506 1783
rect 2503 1758 2507 1759
rect 2503 1753 2507 1754
rect 2462 1747 2468 1748
rect 2462 1743 2463 1747
rect 2467 1743 2468 1747
rect 2462 1742 2468 1743
rect 2454 1733 2460 1734
rect 2504 1733 2506 1753
rect 2350 1728 2356 1729
rect 2370 1731 2376 1732
rect 2370 1727 2371 1731
rect 2375 1727 2376 1731
rect 2454 1729 2455 1733
rect 2459 1729 2460 1733
rect 2502 1732 2508 1733
rect 2454 1728 2460 1729
rect 2470 1731 2476 1732
rect 2370 1726 2376 1727
rect 2470 1727 2471 1731
rect 2475 1727 2476 1731
rect 2502 1728 2503 1732
rect 2507 1728 2508 1732
rect 2502 1727 2508 1728
rect 2470 1726 2476 1727
rect 2438 1712 2444 1713
rect 2438 1708 2439 1712
rect 2443 1708 2444 1712
rect 2438 1707 2444 1708
rect 2439 1706 2443 1707
rect 2439 1701 2443 1702
rect 2438 1700 2444 1701
rect 2438 1696 2439 1700
rect 2443 1696 2444 1700
rect 2438 1695 2444 1696
rect 1446 1679 1452 1680
rect 1446 1675 1447 1679
rect 1451 1675 1452 1679
rect 1446 1674 1452 1675
rect 1550 1679 1556 1680
rect 1550 1675 1551 1679
rect 1555 1675 1556 1679
rect 1550 1674 1556 1675
rect 1662 1679 1668 1680
rect 1662 1675 1663 1679
rect 1667 1675 1668 1679
rect 1662 1674 1668 1675
rect 1670 1679 1676 1680
rect 1670 1675 1671 1679
rect 1675 1675 1676 1679
rect 1670 1674 1676 1675
rect 1774 1679 1780 1680
rect 1774 1675 1775 1679
rect 1779 1675 1780 1679
rect 1774 1674 1780 1675
rect 1894 1679 1900 1680
rect 1894 1675 1895 1679
rect 1899 1675 1900 1679
rect 1894 1674 1900 1675
rect 2030 1679 2036 1680
rect 2030 1675 2031 1679
rect 2035 1675 2036 1679
rect 2030 1674 2036 1675
rect 2174 1679 2180 1680
rect 2174 1675 2175 1679
rect 2179 1675 2180 1679
rect 2174 1674 2180 1675
rect 2326 1679 2332 1680
rect 2326 1675 2327 1679
rect 2331 1675 2332 1679
rect 2326 1674 2332 1675
rect 2342 1679 2348 1680
rect 2342 1675 2343 1679
rect 2347 1675 2348 1679
rect 2342 1674 2348 1675
rect 2454 1679 2460 1680
rect 2454 1675 2455 1679
rect 2459 1675 2460 1679
rect 2454 1674 2460 1675
rect 2462 1679 2468 1680
rect 2462 1675 2463 1679
rect 2467 1675 2468 1679
rect 2462 1674 2468 1675
rect 1382 1663 1388 1664
rect 1382 1659 1383 1663
rect 1387 1659 1388 1663
rect 1382 1658 1388 1659
rect 1438 1663 1444 1664
rect 1438 1659 1439 1663
rect 1443 1659 1444 1663
rect 1438 1658 1444 1659
rect 1448 1647 1450 1674
rect 1552 1647 1554 1674
rect 1664 1647 1666 1674
rect 1672 1669 1674 1674
rect 1671 1668 1675 1669
rect 1671 1663 1675 1664
rect 1776 1647 1778 1674
rect 1896 1647 1898 1674
rect 2032 1647 2034 1674
rect 2176 1647 2178 1674
rect 2328 1647 2330 1674
rect 2346 1659 2352 1660
rect 2346 1655 2347 1659
rect 2351 1655 2352 1659
rect 2346 1654 2352 1655
rect 1431 1646 1435 1647
rect 1431 1641 1435 1642
rect 1447 1646 1451 1647
rect 1447 1641 1451 1642
rect 1519 1646 1523 1647
rect 1519 1641 1523 1642
rect 1551 1646 1555 1647
rect 1551 1641 1555 1642
rect 1599 1646 1603 1647
rect 1599 1641 1603 1642
rect 1663 1646 1667 1647
rect 1663 1641 1667 1642
rect 1679 1646 1683 1647
rect 1679 1641 1683 1642
rect 1751 1646 1755 1647
rect 1751 1641 1755 1642
rect 1775 1646 1779 1647
rect 1775 1641 1779 1642
rect 1839 1646 1843 1647
rect 1839 1641 1843 1642
rect 1895 1646 1899 1647
rect 1895 1641 1899 1642
rect 1935 1646 1939 1647
rect 1935 1641 1939 1642
rect 2031 1646 2035 1647
rect 2031 1641 2035 1642
rect 2055 1646 2059 1647
rect 2175 1646 2179 1647
rect 2055 1641 2059 1642
rect 2138 1643 2144 1644
rect 1374 1635 1380 1636
rect 1374 1631 1375 1635
rect 1379 1631 1380 1635
rect 1374 1630 1380 1631
rect 1432 1622 1434 1641
rect 1520 1622 1522 1641
rect 1600 1622 1602 1641
rect 1680 1622 1682 1641
rect 1752 1622 1754 1641
rect 1840 1622 1842 1641
rect 1936 1622 1938 1641
rect 2056 1622 2058 1641
rect 2138 1639 2139 1643
rect 2143 1639 2144 1643
rect 2175 1641 2179 1642
rect 2183 1646 2187 1647
rect 2183 1641 2187 1642
rect 2327 1646 2331 1647
rect 2327 1641 2331 1642
rect 2138 1638 2144 1639
rect 1366 1621 1372 1622
rect 1286 1619 1292 1620
rect 1326 1620 1332 1621
rect 1190 1618 1196 1619
rect 966 1607 972 1608
rect 966 1603 967 1607
rect 971 1603 972 1607
rect 966 1602 972 1603
rect 1072 1599 1074 1618
rect 1192 1599 1194 1618
rect 1210 1607 1216 1608
rect 1210 1603 1211 1607
rect 1215 1603 1216 1607
rect 1210 1602 1216 1603
rect 815 1598 819 1599
rect 815 1593 819 1594
rect 855 1598 859 1599
rect 870 1598 876 1599
rect 935 1598 939 1599
rect 855 1593 859 1594
rect 935 1593 939 1594
rect 959 1598 963 1599
rect 959 1593 963 1594
rect 1063 1598 1067 1599
rect 1063 1593 1067 1594
rect 1071 1598 1075 1599
rect 1071 1593 1075 1594
rect 1191 1598 1195 1599
rect 1191 1593 1195 1594
rect 806 1587 812 1588
rect 806 1583 807 1587
rect 811 1583 812 1587
rect 806 1582 812 1583
rect 816 1574 818 1593
rect 936 1574 938 1593
rect 990 1587 996 1588
rect 990 1583 991 1587
rect 995 1583 996 1587
rect 990 1582 996 1583
rect 702 1573 708 1574
rect 502 1568 508 1569
rect 526 1571 532 1572
rect 110 1567 116 1568
rect 526 1567 527 1571
rect 531 1567 532 1571
rect 598 1569 599 1573
rect 603 1569 604 1573
rect 598 1568 604 1569
rect 619 1572 623 1573
rect 702 1569 703 1573
rect 707 1569 708 1573
rect 814 1573 820 1574
rect 702 1568 708 1569
rect 742 1571 748 1572
rect 619 1567 623 1568
rect 742 1567 743 1571
rect 747 1567 748 1571
rect 814 1569 815 1573
rect 819 1569 820 1573
rect 814 1568 820 1569
rect 934 1573 940 1574
rect 934 1569 935 1573
rect 939 1569 940 1573
rect 955 1572 959 1573
rect 934 1568 940 1569
rect 526 1566 532 1567
rect 742 1566 748 1567
rect 954 1567 955 1572
rect 959 1567 960 1572
rect 954 1566 960 1567
rect 110 1555 116 1556
rect 110 1551 111 1555
rect 115 1551 116 1555
rect 110 1550 116 1551
rect 270 1552 276 1553
rect 112 1539 114 1550
rect 270 1548 271 1552
rect 275 1548 276 1552
rect 270 1547 276 1548
rect 334 1552 340 1553
rect 334 1548 335 1552
rect 339 1548 340 1552
rect 334 1547 340 1548
rect 406 1552 412 1553
rect 406 1548 407 1552
rect 411 1548 412 1552
rect 406 1547 412 1548
rect 486 1552 492 1553
rect 486 1548 487 1552
rect 491 1548 492 1552
rect 486 1547 492 1548
rect 582 1552 588 1553
rect 582 1548 583 1552
rect 587 1548 588 1552
rect 582 1547 588 1548
rect 686 1552 692 1553
rect 686 1548 687 1552
rect 691 1548 692 1552
rect 686 1547 692 1548
rect 272 1539 274 1547
rect 336 1539 338 1547
rect 408 1539 410 1547
rect 488 1539 490 1547
rect 584 1539 586 1547
rect 688 1539 690 1547
rect 111 1538 115 1539
rect 111 1533 115 1534
rect 271 1538 275 1539
rect 271 1533 275 1534
rect 335 1538 339 1539
rect 335 1533 339 1534
rect 407 1538 411 1539
rect 407 1533 411 1534
rect 471 1538 475 1539
rect 471 1533 475 1534
rect 487 1538 491 1539
rect 487 1533 491 1534
rect 551 1538 555 1539
rect 551 1533 555 1534
rect 583 1538 587 1539
rect 583 1533 587 1534
rect 639 1538 643 1539
rect 639 1533 643 1534
rect 687 1538 691 1539
rect 687 1533 691 1534
rect 735 1538 739 1539
rect 735 1533 739 1534
rect 112 1530 114 1533
rect 470 1532 476 1533
rect 110 1529 116 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 470 1528 471 1532
rect 475 1528 476 1532
rect 470 1527 476 1528
rect 550 1532 556 1533
rect 550 1528 551 1532
rect 555 1528 556 1532
rect 550 1527 556 1528
rect 638 1532 644 1533
rect 638 1528 639 1532
rect 643 1528 644 1532
rect 638 1527 644 1528
rect 734 1532 740 1533
rect 734 1528 735 1532
rect 739 1528 740 1532
rect 734 1527 740 1528
rect 110 1524 116 1525
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 110 1507 116 1508
rect 486 1511 492 1512
rect 486 1507 487 1511
rect 491 1507 492 1511
rect 112 1487 114 1507
rect 486 1506 492 1507
rect 566 1511 572 1512
rect 566 1507 567 1511
rect 571 1507 572 1511
rect 566 1506 572 1507
rect 654 1511 660 1512
rect 654 1507 655 1511
rect 659 1507 660 1511
rect 654 1506 660 1507
rect 662 1511 668 1512
rect 662 1507 663 1511
rect 667 1507 668 1511
rect 662 1506 668 1507
rect 488 1487 490 1506
rect 568 1487 570 1506
rect 656 1487 658 1506
rect 111 1486 115 1487
rect 111 1481 115 1482
rect 375 1486 379 1487
rect 375 1481 379 1482
rect 463 1486 467 1487
rect 463 1481 467 1482
rect 487 1486 491 1487
rect 487 1481 491 1482
rect 559 1486 563 1487
rect 559 1481 563 1482
rect 567 1486 571 1487
rect 567 1481 571 1482
rect 655 1486 659 1487
rect 655 1481 659 1482
rect 112 1461 114 1481
rect 376 1462 378 1481
rect 464 1462 466 1481
rect 560 1462 562 1481
rect 656 1462 658 1481
rect 664 1476 666 1506
rect 744 1496 746 1566
rect 798 1552 804 1553
rect 798 1548 799 1552
rect 803 1548 804 1552
rect 798 1547 804 1548
rect 918 1552 924 1553
rect 918 1548 919 1552
rect 923 1548 924 1552
rect 918 1547 924 1548
rect 800 1539 802 1547
rect 920 1539 922 1547
rect 799 1538 803 1539
rect 799 1533 803 1534
rect 839 1538 843 1539
rect 839 1533 843 1534
rect 919 1538 923 1539
rect 919 1533 923 1534
rect 951 1538 955 1539
rect 951 1533 955 1534
rect 838 1532 844 1533
rect 838 1528 839 1532
rect 843 1528 844 1532
rect 838 1527 844 1528
rect 950 1532 956 1533
rect 950 1528 951 1532
rect 955 1528 956 1532
rect 950 1527 956 1528
rect 992 1512 994 1582
rect 1064 1574 1066 1593
rect 1192 1574 1194 1593
rect 1062 1573 1068 1574
rect 1062 1569 1063 1573
rect 1067 1569 1068 1573
rect 1062 1568 1068 1569
rect 1190 1573 1196 1574
rect 1190 1569 1191 1573
rect 1195 1569 1196 1573
rect 1212 1572 1214 1602
rect 1288 1599 1290 1619
rect 1326 1616 1327 1620
rect 1331 1616 1332 1620
rect 1366 1617 1367 1621
rect 1371 1617 1372 1621
rect 1366 1616 1372 1617
rect 1430 1621 1436 1622
rect 1430 1617 1431 1621
rect 1435 1617 1436 1621
rect 1430 1616 1436 1617
rect 1518 1621 1524 1622
rect 1518 1617 1519 1621
rect 1523 1617 1524 1621
rect 1598 1621 1604 1622
rect 1518 1616 1524 1617
rect 1534 1619 1540 1620
rect 1326 1615 1332 1616
rect 1534 1615 1535 1619
rect 1539 1615 1540 1619
rect 1598 1617 1599 1621
rect 1603 1617 1604 1621
rect 1598 1616 1604 1617
rect 1678 1621 1684 1622
rect 1678 1617 1679 1621
rect 1683 1617 1684 1621
rect 1678 1616 1684 1617
rect 1750 1621 1756 1622
rect 1750 1617 1751 1621
rect 1755 1617 1756 1621
rect 1750 1616 1756 1617
rect 1838 1621 1844 1622
rect 1838 1617 1839 1621
rect 1843 1617 1844 1621
rect 1838 1616 1844 1617
rect 1934 1621 1940 1622
rect 1934 1617 1935 1621
rect 1939 1617 1940 1621
rect 1934 1616 1940 1617
rect 2054 1621 2060 1622
rect 2054 1617 2055 1621
rect 2059 1617 2060 1621
rect 2054 1616 2060 1617
rect 1534 1614 1540 1615
rect 1326 1603 1332 1604
rect 1326 1599 1327 1603
rect 1331 1599 1332 1603
rect 1287 1598 1291 1599
rect 1326 1598 1332 1599
rect 1350 1600 1356 1601
rect 1287 1593 1291 1594
rect 1288 1573 1290 1593
rect 1328 1591 1330 1598
rect 1350 1596 1351 1600
rect 1355 1596 1356 1600
rect 1350 1595 1356 1596
rect 1414 1600 1420 1601
rect 1414 1596 1415 1600
rect 1419 1596 1420 1600
rect 1414 1595 1420 1596
rect 1502 1600 1508 1601
rect 1502 1596 1503 1600
rect 1507 1596 1508 1600
rect 1502 1595 1508 1596
rect 1352 1591 1354 1595
rect 1416 1591 1418 1595
rect 1504 1591 1506 1595
rect 1327 1590 1331 1591
rect 1327 1585 1331 1586
rect 1351 1590 1355 1591
rect 1351 1585 1355 1586
rect 1415 1590 1419 1591
rect 1415 1585 1419 1586
rect 1423 1590 1427 1591
rect 1423 1585 1427 1586
rect 1503 1590 1507 1591
rect 1503 1585 1507 1586
rect 1527 1590 1531 1591
rect 1527 1585 1531 1586
rect 1328 1582 1330 1585
rect 1350 1584 1356 1585
rect 1326 1581 1332 1582
rect 1326 1577 1327 1581
rect 1331 1577 1332 1581
rect 1350 1580 1351 1584
rect 1355 1580 1356 1584
rect 1350 1579 1356 1580
rect 1422 1584 1428 1585
rect 1422 1580 1423 1584
rect 1427 1580 1428 1584
rect 1422 1579 1428 1580
rect 1526 1584 1532 1585
rect 1526 1580 1527 1584
rect 1531 1580 1532 1584
rect 1526 1579 1532 1580
rect 1326 1576 1332 1577
rect 1286 1572 1292 1573
rect 1190 1568 1196 1569
rect 1210 1571 1216 1572
rect 1210 1567 1211 1571
rect 1215 1567 1216 1571
rect 1286 1568 1287 1572
rect 1291 1568 1292 1572
rect 1286 1567 1292 1568
rect 1210 1566 1216 1567
rect 1326 1564 1332 1565
rect 1326 1560 1327 1564
rect 1331 1560 1332 1564
rect 1326 1559 1332 1560
rect 1366 1563 1372 1564
rect 1366 1559 1367 1563
rect 1371 1559 1372 1563
rect 1286 1555 1292 1556
rect 1046 1552 1052 1553
rect 1046 1548 1047 1552
rect 1051 1548 1052 1552
rect 1046 1547 1052 1548
rect 1174 1552 1180 1553
rect 1174 1548 1175 1552
rect 1179 1548 1180 1552
rect 1286 1551 1287 1555
rect 1291 1551 1292 1555
rect 1286 1550 1292 1551
rect 1174 1547 1180 1548
rect 1048 1539 1050 1547
rect 1176 1539 1178 1547
rect 1288 1539 1290 1550
rect 1328 1539 1330 1559
rect 1366 1558 1372 1559
rect 1374 1563 1380 1564
rect 1374 1559 1375 1563
rect 1379 1559 1380 1563
rect 1374 1558 1380 1559
rect 1438 1563 1444 1564
rect 1438 1559 1439 1563
rect 1443 1559 1444 1563
rect 1438 1558 1444 1559
rect 1368 1539 1370 1558
rect 1047 1538 1051 1539
rect 1047 1533 1051 1534
rect 1063 1538 1067 1539
rect 1063 1533 1067 1534
rect 1175 1538 1179 1539
rect 1175 1533 1179 1534
rect 1287 1538 1291 1539
rect 1287 1533 1291 1534
rect 1327 1538 1331 1539
rect 1327 1533 1331 1534
rect 1367 1538 1371 1539
rect 1367 1533 1371 1534
rect 1062 1532 1068 1533
rect 1062 1528 1063 1532
rect 1067 1528 1068 1532
rect 1062 1527 1068 1528
rect 1174 1532 1180 1533
rect 1174 1528 1175 1532
rect 1179 1528 1180 1532
rect 1288 1530 1290 1533
rect 1174 1527 1180 1528
rect 1286 1529 1292 1530
rect 1286 1525 1287 1529
rect 1291 1525 1292 1529
rect 1286 1524 1292 1525
rect 1328 1513 1330 1533
rect 1368 1514 1370 1533
rect 1376 1528 1378 1558
rect 1440 1539 1442 1558
rect 1536 1548 1538 1614
rect 1582 1600 1588 1601
rect 1582 1596 1583 1600
rect 1587 1596 1588 1600
rect 1582 1595 1588 1596
rect 1662 1600 1668 1601
rect 1662 1596 1663 1600
rect 1667 1596 1668 1600
rect 1662 1595 1668 1596
rect 1734 1600 1740 1601
rect 1734 1596 1735 1600
rect 1739 1596 1740 1600
rect 1734 1595 1740 1596
rect 1822 1600 1828 1601
rect 1822 1596 1823 1600
rect 1827 1596 1828 1600
rect 1822 1595 1828 1596
rect 1918 1600 1924 1601
rect 1918 1596 1919 1600
rect 1923 1596 1924 1600
rect 1918 1595 1924 1596
rect 2038 1600 2044 1601
rect 2038 1596 2039 1600
rect 2043 1596 2044 1600
rect 2038 1595 2044 1596
rect 1584 1591 1586 1595
rect 1664 1591 1666 1595
rect 1736 1591 1738 1595
rect 1824 1591 1826 1595
rect 1920 1591 1922 1595
rect 2040 1591 2042 1595
rect 1583 1590 1587 1591
rect 1583 1585 1587 1586
rect 1647 1590 1651 1591
rect 1647 1585 1651 1586
rect 1663 1590 1667 1591
rect 1663 1585 1667 1586
rect 1735 1590 1739 1591
rect 1735 1585 1739 1586
rect 1783 1590 1787 1591
rect 1783 1585 1787 1586
rect 1823 1590 1827 1591
rect 1823 1585 1827 1586
rect 1919 1590 1923 1591
rect 1919 1585 1923 1586
rect 1935 1590 1939 1591
rect 1935 1585 1939 1586
rect 2039 1590 2043 1591
rect 2039 1585 2043 1586
rect 2103 1590 2107 1591
rect 2103 1585 2107 1586
rect 1646 1584 1652 1585
rect 1646 1580 1647 1584
rect 1651 1580 1652 1584
rect 1646 1579 1652 1580
rect 1782 1584 1788 1585
rect 1782 1580 1783 1584
rect 1787 1580 1788 1584
rect 1782 1579 1788 1580
rect 1934 1584 1940 1585
rect 1934 1580 1935 1584
rect 1939 1580 1940 1584
rect 1934 1579 1940 1580
rect 2102 1584 2108 1585
rect 2102 1580 2103 1584
rect 2107 1580 2108 1584
rect 2102 1579 2108 1580
rect 2140 1564 2142 1638
rect 2184 1622 2186 1641
rect 2328 1622 2330 1641
rect 2182 1621 2188 1622
rect 2182 1617 2183 1621
rect 2187 1617 2188 1621
rect 2182 1616 2188 1617
rect 2326 1621 2332 1622
rect 2326 1617 2327 1621
rect 2331 1617 2332 1621
rect 2348 1620 2350 1654
rect 2456 1647 2458 1674
rect 2455 1646 2459 1647
rect 2455 1641 2459 1642
rect 2456 1622 2458 1641
rect 2464 1636 2466 1674
rect 2472 1664 2474 1726
rect 2502 1715 2508 1716
rect 2502 1711 2503 1715
rect 2507 1711 2508 1715
rect 2502 1710 2508 1711
rect 2504 1707 2506 1710
rect 2503 1706 2507 1707
rect 2503 1701 2507 1702
rect 2504 1698 2506 1701
rect 2502 1697 2508 1698
rect 2502 1693 2503 1697
rect 2507 1693 2508 1697
rect 2502 1692 2508 1693
rect 2502 1680 2508 1681
rect 2502 1676 2503 1680
rect 2507 1676 2508 1680
rect 2502 1675 2508 1676
rect 2470 1663 2476 1664
rect 2470 1659 2471 1663
rect 2475 1659 2476 1663
rect 2470 1658 2476 1659
rect 2504 1647 2506 1675
rect 2503 1646 2507 1647
rect 2503 1641 2507 1642
rect 2462 1635 2468 1636
rect 2462 1631 2463 1635
rect 2467 1631 2468 1635
rect 2462 1630 2468 1631
rect 2454 1621 2460 1622
rect 2504 1621 2506 1641
rect 2326 1616 2332 1617
rect 2346 1619 2352 1620
rect 2346 1615 2347 1619
rect 2351 1615 2352 1619
rect 2454 1617 2455 1621
rect 2459 1617 2460 1621
rect 2502 1620 2508 1621
rect 2454 1616 2460 1617
rect 2462 1619 2468 1620
rect 2346 1614 2352 1615
rect 2462 1615 2463 1619
rect 2467 1615 2468 1619
rect 2502 1616 2503 1620
rect 2507 1616 2508 1620
rect 2502 1615 2508 1616
rect 2462 1614 2468 1615
rect 2166 1600 2172 1601
rect 2166 1596 2167 1600
rect 2171 1596 2172 1600
rect 2166 1595 2172 1596
rect 2310 1600 2316 1601
rect 2310 1596 2311 1600
rect 2315 1596 2316 1600
rect 2310 1595 2316 1596
rect 2438 1600 2444 1601
rect 2438 1596 2439 1600
rect 2443 1596 2444 1600
rect 2438 1595 2444 1596
rect 2168 1591 2170 1595
rect 2312 1591 2314 1595
rect 2440 1591 2442 1595
rect 2167 1590 2171 1591
rect 2167 1585 2171 1586
rect 2279 1590 2283 1591
rect 2279 1585 2283 1586
rect 2311 1590 2315 1591
rect 2311 1585 2315 1586
rect 2439 1590 2443 1591
rect 2439 1585 2443 1586
rect 2278 1584 2284 1585
rect 2278 1580 2279 1584
rect 2283 1580 2284 1584
rect 2278 1579 2284 1580
rect 2438 1584 2444 1585
rect 2438 1580 2439 1584
rect 2443 1580 2444 1584
rect 2438 1579 2444 1580
rect 1542 1563 1548 1564
rect 1542 1559 1543 1563
rect 1547 1559 1548 1563
rect 1542 1558 1548 1559
rect 1662 1563 1668 1564
rect 1662 1559 1663 1563
rect 1667 1559 1668 1563
rect 1662 1558 1668 1559
rect 1798 1563 1804 1564
rect 1798 1559 1799 1563
rect 1803 1559 1804 1563
rect 1798 1558 1804 1559
rect 1950 1563 1956 1564
rect 1950 1559 1951 1563
rect 1955 1559 1956 1563
rect 1950 1558 1956 1559
rect 2118 1563 2124 1564
rect 2118 1559 2119 1563
rect 2123 1559 2124 1563
rect 2118 1558 2124 1559
rect 2138 1563 2144 1564
rect 2138 1559 2139 1563
rect 2143 1559 2144 1563
rect 2138 1558 2144 1559
rect 2294 1563 2300 1564
rect 2294 1559 2295 1563
rect 2299 1559 2300 1563
rect 2294 1558 2300 1559
rect 2310 1563 2316 1564
rect 2310 1559 2311 1563
rect 2315 1559 2316 1563
rect 2310 1558 2316 1559
rect 2454 1563 2460 1564
rect 2454 1559 2455 1563
rect 2459 1559 2460 1563
rect 2454 1558 2460 1559
rect 1534 1547 1540 1548
rect 1534 1543 1535 1547
rect 1539 1543 1540 1547
rect 1534 1542 1540 1543
rect 1544 1539 1546 1558
rect 1664 1539 1666 1558
rect 1800 1539 1802 1558
rect 1874 1543 1880 1544
rect 1874 1539 1875 1543
rect 1879 1539 1880 1543
rect 1952 1539 1954 1558
rect 2120 1539 2122 1558
rect 2270 1547 2276 1548
rect 2270 1543 2271 1547
rect 2275 1543 2276 1547
rect 2270 1542 2276 1543
rect 1439 1538 1443 1539
rect 1439 1533 1443 1534
rect 1543 1538 1547 1539
rect 1543 1533 1547 1534
rect 1647 1538 1651 1539
rect 1647 1533 1651 1534
rect 1663 1538 1667 1539
rect 1663 1533 1667 1534
rect 1751 1538 1755 1539
rect 1751 1533 1755 1534
rect 1799 1538 1803 1539
rect 1799 1533 1803 1534
rect 1855 1538 1859 1539
rect 1874 1538 1880 1539
rect 1951 1538 1955 1539
rect 1855 1533 1859 1534
rect 1374 1527 1380 1528
rect 1374 1523 1375 1527
rect 1379 1523 1380 1527
rect 1374 1522 1380 1523
rect 1440 1514 1442 1533
rect 1470 1519 1476 1520
rect 1470 1515 1471 1519
rect 1475 1515 1476 1519
rect 1470 1514 1476 1515
rect 1544 1514 1546 1533
rect 1648 1514 1650 1533
rect 1654 1527 1660 1528
rect 1654 1523 1655 1527
rect 1659 1523 1660 1527
rect 1654 1522 1660 1523
rect 1366 1513 1372 1514
rect 1286 1512 1292 1513
rect 750 1511 756 1512
rect 750 1507 751 1511
rect 755 1507 756 1511
rect 750 1506 756 1507
rect 854 1511 860 1512
rect 854 1507 855 1511
rect 859 1507 860 1511
rect 854 1506 860 1507
rect 870 1511 876 1512
rect 870 1507 871 1511
rect 875 1507 876 1511
rect 870 1506 876 1507
rect 966 1511 972 1512
rect 966 1507 967 1511
rect 971 1507 972 1511
rect 966 1506 972 1507
rect 990 1511 996 1512
rect 990 1507 991 1511
rect 995 1507 996 1511
rect 990 1506 996 1507
rect 1078 1511 1084 1512
rect 1078 1507 1079 1511
rect 1083 1507 1084 1511
rect 1078 1506 1084 1507
rect 1094 1511 1100 1512
rect 1094 1507 1095 1511
rect 1099 1507 1100 1511
rect 1094 1506 1100 1507
rect 1190 1511 1196 1512
rect 1190 1507 1191 1511
rect 1195 1507 1196 1511
rect 1286 1508 1287 1512
rect 1291 1508 1292 1512
rect 1286 1507 1292 1508
rect 1326 1512 1332 1513
rect 1326 1508 1327 1512
rect 1331 1508 1332 1512
rect 1366 1509 1367 1513
rect 1371 1509 1372 1513
rect 1366 1508 1372 1509
rect 1438 1513 1444 1514
rect 1438 1509 1439 1513
rect 1443 1509 1444 1513
rect 1438 1508 1444 1509
rect 1326 1507 1332 1508
rect 1190 1506 1196 1507
rect 742 1495 748 1496
rect 742 1491 743 1495
rect 747 1491 748 1495
rect 742 1490 748 1491
rect 752 1487 754 1506
rect 856 1487 858 1506
rect 872 1492 874 1506
rect 870 1491 876 1492
rect 870 1487 871 1491
rect 875 1487 876 1491
rect 968 1487 970 1506
rect 1080 1487 1082 1506
rect 1096 1492 1098 1506
rect 1094 1491 1100 1492
rect 1094 1487 1095 1491
rect 1099 1487 1100 1491
rect 1192 1487 1194 1506
rect 1198 1495 1204 1496
rect 1198 1491 1199 1495
rect 1203 1491 1204 1495
rect 1198 1490 1204 1491
rect 751 1486 755 1487
rect 751 1481 755 1482
rect 855 1486 859 1487
rect 870 1486 876 1487
rect 959 1486 963 1487
rect 855 1481 859 1482
rect 959 1481 963 1482
rect 967 1486 971 1487
rect 967 1481 971 1482
rect 1063 1486 1067 1487
rect 1063 1481 1067 1482
rect 1079 1486 1083 1487
rect 1094 1486 1100 1487
rect 1167 1486 1171 1487
rect 1079 1481 1083 1482
rect 1122 1483 1128 1484
rect 662 1475 668 1476
rect 662 1471 663 1475
rect 667 1471 668 1475
rect 662 1470 668 1471
rect 752 1462 754 1481
rect 770 1479 776 1480
rect 770 1475 771 1479
rect 775 1475 776 1479
rect 770 1474 776 1475
rect 374 1461 380 1462
rect 110 1460 116 1461
rect 110 1456 111 1460
rect 115 1456 116 1460
rect 374 1457 375 1461
rect 379 1457 380 1461
rect 374 1456 380 1457
rect 462 1461 468 1462
rect 462 1457 463 1461
rect 467 1457 468 1461
rect 462 1456 468 1457
rect 558 1461 564 1462
rect 558 1457 559 1461
rect 563 1457 564 1461
rect 654 1461 660 1462
rect 558 1456 564 1457
rect 622 1459 628 1460
rect 110 1455 116 1456
rect 622 1455 623 1459
rect 627 1455 628 1459
rect 654 1457 655 1461
rect 659 1457 660 1461
rect 654 1456 660 1457
rect 750 1461 756 1462
rect 750 1457 751 1461
rect 755 1457 756 1461
rect 772 1460 774 1474
rect 856 1462 858 1481
rect 960 1462 962 1481
rect 1064 1462 1066 1481
rect 1122 1479 1123 1483
rect 1127 1479 1128 1483
rect 1167 1481 1171 1482
rect 1191 1486 1195 1487
rect 1191 1481 1195 1482
rect 1122 1478 1128 1479
rect 854 1461 860 1462
rect 750 1456 756 1457
rect 770 1459 776 1460
rect 622 1454 628 1455
rect 770 1455 771 1459
rect 775 1455 776 1459
rect 854 1457 855 1461
rect 859 1457 860 1461
rect 854 1456 860 1457
rect 958 1461 964 1462
rect 958 1457 959 1461
rect 963 1457 964 1461
rect 958 1456 964 1457
rect 1062 1461 1068 1462
rect 1062 1457 1063 1461
rect 1067 1457 1068 1461
rect 1062 1456 1068 1457
rect 770 1454 776 1455
rect 110 1443 116 1444
rect 110 1439 111 1443
rect 115 1439 116 1443
rect 110 1438 116 1439
rect 358 1440 364 1441
rect 112 1435 114 1438
rect 358 1436 359 1440
rect 363 1436 364 1440
rect 358 1435 364 1436
rect 446 1440 452 1441
rect 446 1436 447 1440
rect 451 1436 452 1440
rect 446 1435 452 1436
rect 542 1440 548 1441
rect 542 1436 543 1440
rect 547 1436 548 1440
rect 542 1435 548 1436
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 231 1434 235 1435
rect 231 1429 235 1430
rect 319 1434 323 1435
rect 319 1429 323 1430
rect 359 1434 363 1435
rect 359 1429 363 1430
rect 415 1434 419 1435
rect 415 1429 419 1430
rect 447 1434 451 1435
rect 447 1429 451 1430
rect 511 1434 515 1435
rect 511 1429 515 1430
rect 543 1434 547 1435
rect 543 1429 547 1430
rect 615 1434 619 1435
rect 615 1429 619 1430
rect 112 1426 114 1429
rect 230 1428 236 1429
rect 110 1425 116 1426
rect 110 1421 111 1425
rect 115 1421 116 1425
rect 230 1424 231 1428
rect 235 1424 236 1428
rect 230 1423 236 1424
rect 318 1428 324 1429
rect 318 1424 319 1428
rect 323 1424 324 1428
rect 318 1423 324 1424
rect 414 1428 420 1429
rect 414 1424 415 1428
rect 419 1424 420 1428
rect 414 1423 420 1424
rect 510 1428 516 1429
rect 510 1424 511 1428
rect 515 1424 516 1428
rect 510 1423 516 1424
rect 614 1428 620 1429
rect 614 1424 615 1428
rect 619 1424 620 1428
rect 614 1423 620 1424
rect 110 1420 116 1421
rect 110 1408 116 1409
rect 110 1404 111 1408
rect 115 1404 116 1408
rect 110 1403 116 1404
rect 246 1407 252 1408
rect 246 1403 247 1407
rect 251 1403 252 1407
rect 112 1383 114 1403
rect 246 1402 252 1403
rect 334 1407 340 1408
rect 334 1403 335 1407
rect 339 1403 340 1407
rect 334 1402 340 1403
rect 430 1407 436 1408
rect 430 1403 431 1407
rect 435 1403 436 1407
rect 430 1402 436 1403
rect 502 1407 508 1408
rect 502 1403 503 1407
rect 507 1403 508 1407
rect 502 1402 508 1403
rect 526 1407 532 1408
rect 526 1403 527 1407
rect 531 1403 532 1407
rect 526 1402 532 1403
rect 542 1407 548 1408
rect 542 1403 543 1407
rect 547 1403 548 1407
rect 542 1402 548 1403
rect 248 1383 250 1402
rect 336 1383 338 1402
rect 432 1383 434 1402
rect 111 1382 115 1383
rect 111 1377 115 1378
rect 151 1382 155 1383
rect 151 1377 155 1378
rect 215 1382 219 1383
rect 215 1377 219 1378
rect 247 1382 251 1383
rect 247 1377 251 1378
rect 311 1382 315 1383
rect 311 1377 315 1378
rect 335 1382 339 1383
rect 335 1377 339 1378
rect 407 1382 411 1383
rect 407 1377 411 1378
rect 431 1382 435 1383
rect 431 1377 435 1378
rect 112 1357 114 1377
rect 152 1358 154 1377
rect 216 1358 218 1377
rect 312 1358 314 1377
rect 408 1358 410 1377
rect 504 1372 506 1402
rect 528 1383 530 1402
rect 544 1388 546 1402
rect 624 1392 626 1454
rect 638 1440 644 1441
rect 638 1436 639 1440
rect 643 1436 644 1440
rect 638 1435 644 1436
rect 734 1440 740 1441
rect 734 1436 735 1440
rect 739 1436 740 1440
rect 734 1435 740 1436
rect 838 1440 844 1441
rect 838 1436 839 1440
rect 843 1436 844 1440
rect 838 1435 844 1436
rect 942 1440 948 1441
rect 942 1436 943 1440
rect 947 1436 948 1440
rect 942 1435 948 1436
rect 1046 1440 1052 1441
rect 1046 1436 1047 1440
rect 1051 1436 1052 1440
rect 1046 1435 1052 1436
rect 639 1434 643 1435
rect 639 1429 643 1430
rect 711 1434 715 1435
rect 711 1429 715 1430
rect 735 1434 739 1435
rect 735 1429 739 1430
rect 807 1434 811 1435
rect 807 1429 811 1430
rect 839 1434 843 1435
rect 839 1429 843 1430
rect 895 1434 899 1435
rect 895 1429 899 1430
rect 943 1434 947 1435
rect 943 1429 947 1430
rect 991 1434 995 1435
rect 991 1429 995 1430
rect 1047 1434 1051 1435
rect 1047 1429 1051 1430
rect 1087 1434 1091 1435
rect 1087 1429 1091 1430
rect 710 1428 716 1429
rect 710 1424 711 1428
rect 715 1424 716 1428
rect 710 1423 716 1424
rect 806 1428 812 1429
rect 806 1424 807 1428
rect 811 1424 812 1428
rect 806 1423 812 1424
rect 894 1428 900 1429
rect 894 1424 895 1428
rect 899 1424 900 1428
rect 894 1423 900 1424
rect 990 1428 996 1429
rect 990 1424 991 1428
rect 995 1424 996 1428
rect 990 1423 996 1424
rect 1086 1428 1092 1429
rect 1086 1424 1087 1428
rect 1091 1424 1092 1428
rect 1086 1423 1092 1424
rect 1124 1408 1126 1478
rect 1168 1462 1170 1481
rect 1166 1461 1172 1462
rect 1166 1457 1167 1461
rect 1171 1457 1172 1461
rect 1200 1460 1202 1490
rect 1288 1487 1290 1507
rect 1326 1495 1332 1496
rect 1326 1491 1327 1495
rect 1331 1491 1332 1495
rect 1326 1490 1332 1491
rect 1350 1492 1356 1493
rect 1287 1486 1291 1487
rect 1328 1483 1330 1490
rect 1350 1488 1351 1492
rect 1355 1488 1356 1492
rect 1350 1487 1356 1488
rect 1422 1492 1428 1493
rect 1422 1488 1423 1492
rect 1427 1488 1428 1492
rect 1422 1487 1428 1488
rect 1352 1483 1354 1487
rect 1424 1483 1426 1487
rect 1287 1481 1291 1482
rect 1327 1482 1331 1483
rect 1288 1461 1290 1481
rect 1327 1477 1331 1478
rect 1351 1482 1355 1483
rect 1351 1477 1355 1478
rect 1423 1482 1427 1483
rect 1423 1477 1427 1478
rect 1328 1474 1330 1477
rect 1350 1476 1356 1477
rect 1326 1473 1332 1474
rect 1326 1469 1327 1473
rect 1331 1469 1332 1473
rect 1350 1472 1351 1476
rect 1355 1472 1356 1476
rect 1350 1471 1356 1472
rect 1422 1476 1428 1477
rect 1422 1472 1423 1476
rect 1427 1472 1428 1476
rect 1422 1471 1428 1472
rect 1326 1468 1332 1469
rect 1286 1460 1292 1461
rect 1166 1456 1172 1457
rect 1198 1459 1204 1460
rect 1198 1455 1199 1459
rect 1203 1455 1204 1459
rect 1286 1456 1287 1460
rect 1291 1456 1292 1460
rect 1286 1455 1292 1456
rect 1326 1456 1332 1457
rect 1198 1454 1204 1455
rect 1326 1452 1327 1456
rect 1331 1452 1332 1456
rect 1326 1451 1332 1452
rect 1366 1455 1372 1456
rect 1366 1451 1367 1455
rect 1371 1451 1372 1455
rect 1286 1443 1292 1444
rect 1150 1440 1156 1441
rect 1150 1436 1151 1440
rect 1155 1436 1156 1440
rect 1286 1439 1287 1443
rect 1291 1439 1292 1443
rect 1286 1438 1292 1439
rect 1150 1435 1156 1436
rect 1288 1435 1290 1438
rect 1151 1434 1155 1435
rect 1151 1429 1155 1430
rect 1287 1434 1291 1435
rect 1287 1429 1291 1430
rect 1288 1426 1290 1429
rect 1328 1427 1330 1451
rect 1366 1450 1372 1451
rect 1414 1455 1420 1456
rect 1414 1451 1415 1455
rect 1419 1451 1420 1455
rect 1414 1450 1420 1451
rect 1438 1455 1444 1456
rect 1438 1451 1439 1455
rect 1443 1451 1444 1455
rect 1438 1450 1444 1451
rect 1368 1427 1370 1450
rect 1327 1426 1331 1427
rect 1286 1425 1292 1426
rect 1286 1421 1287 1425
rect 1291 1421 1292 1425
rect 1327 1421 1331 1422
rect 1367 1426 1371 1427
rect 1367 1421 1371 1422
rect 1286 1420 1292 1421
rect 1286 1408 1292 1409
rect 630 1407 636 1408
rect 630 1403 631 1407
rect 635 1403 636 1407
rect 630 1402 636 1403
rect 726 1407 732 1408
rect 726 1403 727 1407
rect 731 1403 732 1407
rect 726 1402 732 1403
rect 822 1407 828 1408
rect 822 1403 823 1407
rect 827 1403 828 1407
rect 822 1402 828 1403
rect 910 1407 916 1408
rect 910 1403 911 1407
rect 915 1403 916 1407
rect 910 1402 916 1403
rect 1006 1407 1012 1408
rect 1006 1403 1007 1407
rect 1011 1403 1012 1407
rect 1006 1402 1012 1403
rect 1102 1407 1108 1408
rect 1102 1403 1103 1407
rect 1107 1403 1108 1407
rect 1102 1402 1108 1403
rect 1122 1407 1128 1408
rect 1122 1403 1123 1407
rect 1127 1403 1128 1407
rect 1286 1404 1287 1408
rect 1291 1404 1292 1408
rect 1286 1403 1292 1404
rect 1122 1402 1128 1403
rect 622 1391 628 1392
rect 542 1387 548 1388
rect 542 1383 543 1387
rect 547 1383 548 1387
rect 622 1387 623 1391
rect 627 1387 628 1391
rect 622 1386 628 1387
rect 632 1383 634 1402
rect 728 1383 730 1402
rect 824 1383 826 1402
rect 912 1383 914 1402
rect 1008 1383 1010 1402
rect 1022 1387 1028 1388
rect 1022 1383 1023 1387
rect 1027 1383 1028 1387
rect 1104 1383 1106 1402
rect 1288 1383 1290 1403
rect 1328 1401 1330 1421
rect 1368 1402 1370 1421
rect 1416 1416 1418 1450
rect 1440 1427 1442 1450
rect 1472 1440 1474 1514
rect 1542 1513 1548 1514
rect 1542 1509 1543 1513
rect 1547 1509 1548 1513
rect 1542 1508 1548 1509
rect 1646 1513 1652 1514
rect 1646 1509 1647 1513
rect 1651 1509 1652 1513
rect 1646 1508 1652 1509
rect 1526 1492 1532 1493
rect 1526 1488 1527 1492
rect 1531 1488 1532 1492
rect 1526 1487 1532 1488
rect 1630 1492 1636 1493
rect 1630 1488 1631 1492
rect 1635 1488 1636 1492
rect 1630 1487 1636 1488
rect 1528 1483 1530 1487
rect 1632 1483 1634 1487
rect 1519 1482 1523 1483
rect 1519 1477 1523 1478
rect 1527 1482 1531 1483
rect 1527 1477 1531 1478
rect 1615 1482 1619 1483
rect 1615 1477 1619 1478
rect 1631 1482 1635 1483
rect 1631 1477 1635 1478
rect 1518 1476 1524 1477
rect 1518 1472 1519 1476
rect 1523 1472 1524 1476
rect 1518 1471 1524 1472
rect 1614 1476 1620 1477
rect 1614 1472 1615 1476
rect 1619 1472 1620 1476
rect 1614 1471 1620 1472
rect 1656 1456 1658 1522
rect 1752 1514 1754 1533
rect 1856 1514 1858 1533
rect 1750 1513 1756 1514
rect 1750 1509 1751 1513
rect 1755 1509 1756 1513
rect 1750 1508 1756 1509
rect 1854 1513 1860 1514
rect 1854 1509 1855 1513
rect 1859 1509 1860 1513
rect 1876 1512 1878 1538
rect 1951 1533 1955 1534
rect 1959 1538 1963 1539
rect 1959 1533 1963 1534
rect 2055 1538 2059 1539
rect 2055 1533 2059 1534
rect 2119 1538 2123 1539
rect 2119 1533 2123 1534
rect 2151 1538 2155 1539
rect 2151 1533 2155 1534
rect 2247 1538 2251 1539
rect 2247 1533 2251 1534
rect 1960 1514 1962 1533
rect 2056 1514 2058 1533
rect 2152 1514 2154 1533
rect 2248 1514 2250 1533
rect 1958 1513 1964 1514
rect 1854 1508 1860 1509
rect 1874 1511 1880 1512
rect 1874 1507 1875 1511
rect 1879 1507 1880 1511
rect 1958 1509 1959 1513
rect 1963 1509 1964 1513
rect 1958 1508 1964 1509
rect 2054 1513 2060 1514
rect 2054 1509 2055 1513
rect 2059 1509 2060 1513
rect 2150 1513 2156 1514
rect 2054 1508 2060 1509
rect 2142 1511 2148 1512
rect 1874 1506 1880 1507
rect 2142 1507 2143 1511
rect 2147 1507 2148 1511
rect 2150 1509 2151 1513
rect 2155 1509 2156 1513
rect 2150 1508 2156 1509
rect 2246 1513 2252 1514
rect 2246 1509 2247 1513
rect 2251 1509 2252 1513
rect 2272 1512 2274 1542
rect 2296 1539 2298 1558
rect 2312 1544 2314 1558
rect 2310 1543 2316 1544
rect 2310 1539 2311 1543
rect 2315 1539 2316 1543
rect 2456 1539 2458 1558
rect 2464 1548 2466 1614
rect 2502 1603 2508 1604
rect 2502 1599 2503 1603
rect 2507 1599 2508 1603
rect 2502 1598 2508 1599
rect 2504 1591 2506 1598
rect 2503 1590 2507 1591
rect 2503 1585 2507 1586
rect 2504 1582 2506 1585
rect 2502 1581 2508 1582
rect 2502 1577 2503 1581
rect 2507 1577 2508 1581
rect 2502 1576 2508 1577
rect 2502 1564 2508 1565
rect 2470 1563 2476 1564
rect 2470 1559 2471 1563
rect 2475 1559 2476 1563
rect 2502 1560 2503 1564
rect 2507 1560 2508 1564
rect 2502 1559 2508 1560
rect 2470 1558 2476 1559
rect 2462 1547 2468 1548
rect 2462 1543 2463 1547
rect 2467 1543 2468 1547
rect 2462 1542 2468 1543
rect 2295 1538 2299 1539
rect 2310 1538 2316 1539
rect 2343 1538 2347 1539
rect 2295 1533 2299 1534
rect 2439 1538 2443 1539
rect 2343 1533 2347 1534
rect 2362 1535 2368 1536
rect 2344 1514 2346 1533
rect 2362 1531 2363 1535
rect 2367 1531 2368 1535
rect 2439 1533 2443 1534
rect 2455 1538 2459 1539
rect 2455 1533 2459 1534
rect 2362 1530 2368 1531
rect 2350 1527 2356 1528
rect 2350 1523 2351 1527
rect 2355 1523 2356 1527
rect 2350 1522 2356 1523
rect 2342 1513 2348 1514
rect 2246 1508 2252 1509
rect 2270 1511 2276 1512
rect 2142 1506 2148 1507
rect 2270 1507 2271 1511
rect 2275 1507 2276 1511
rect 2342 1509 2343 1513
rect 2347 1509 2348 1513
rect 2342 1508 2348 1509
rect 2270 1506 2276 1507
rect 1734 1492 1740 1493
rect 1734 1488 1735 1492
rect 1739 1488 1740 1492
rect 1734 1487 1740 1488
rect 1838 1492 1844 1493
rect 1838 1488 1839 1492
rect 1843 1488 1844 1492
rect 1838 1487 1844 1488
rect 1942 1492 1948 1493
rect 1942 1488 1943 1492
rect 1947 1488 1948 1492
rect 1942 1487 1948 1488
rect 2038 1492 2044 1493
rect 2038 1488 2039 1492
rect 2043 1488 2044 1492
rect 2038 1487 2044 1488
rect 2134 1492 2140 1493
rect 2134 1488 2135 1492
rect 2139 1488 2140 1492
rect 2134 1487 2140 1488
rect 1736 1483 1738 1487
rect 1840 1483 1842 1487
rect 1944 1483 1946 1487
rect 2040 1483 2042 1487
rect 2136 1483 2138 1487
rect 1711 1482 1715 1483
rect 1711 1477 1715 1478
rect 1735 1482 1739 1483
rect 1735 1477 1739 1478
rect 1815 1482 1819 1483
rect 1815 1477 1819 1478
rect 1839 1482 1843 1483
rect 1839 1477 1843 1478
rect 1927 1482 1931 1483
rect 1927 1477 1931 1478
rect 1943 1482 1947 1483
rect 1943 1477 1947 1478
rect 2039 1482 2043 1483
rect 2039 1477 2043 1478
rect 2047 1482 2051 1483
rect 2047 1477 2051 1478
rect 2135 1482 2139 1483
rect 2135 1477 2139 1478
rect 1710 1476 1716 1477
rect 1710 1472 1711 1476
rect 1715 1472 1716 1476
rect 1710 1471 1716 1472
rect 1814 1476 1820 1477
rect 1814 1472 1815 1476
rect 1819 1472 1820 1476
rect 1814 1471 1820 1472
rect 1926 1476 1932 1477
rect 1926 1472 1927 1476
rect 1931 1472 1932 1476
rect 1926 1471 1932 1472
rect 2046 1476 2052 1477
rect 2046 1472 2047 1476
rect 2051 1472 2052 1476
rect 2046 1471 2052 1472
rect 1534 1455 1540 1456
rect 1534 1451 1535 1455
rect 1539 1451 1540 1455
rect 1534 1450 1540 1451
rect 1630 1455 1636 1456
rect 1630 1451 1631 1455
rect 1635 1451 1636 1455
rect 1630 1450 1636 1451
rect 1654 1455 1660 1456
rect 1654 1451 1655 1455
rect 1659 1451 1660 1455
rect 1654 1450 1660 1451
rect 1726 1455 1732 1456
rect 1726 1451 1727 1455
rect 1731 1451 1732 1455
rect 1726 1450 1732 1451
rect 1830 1455 1836 1456
rect 1830 1451 1831 1455
rect 1835 1451 1836 1455
rect 1830 1450 1836 1451
rect 1838 1455 1844 1456
rect 1838 1451 1839 1455
rect 1843 1451 1844 1455
rect 1838 1450 1844 1451
rect 1942 1455 1948 1456
rect 1942 1451 1943 1455
rect 1947 1451 1948 1455
rect 1942 1450 1948 1451
rect 1958 1455 1964 1456
rect 1958 1451 1959 1455
rect 1963 1451 1964 1455
rect 1958 1450 1964 1451
rect 2062 1455 2068 1456
rect 2062 1451 2063 1455
rect 2067 1451 2068 1455
rect 2062 1450 2068 1451
rect 1470 1439 1476 1440
rect 1470 1435 1471 1439
rect 1475 1435 1476 1439
rect 1470 1434 1476 1435
rect 1536 1427 1538 1450
rect 1632 1427 1634 1450
rect 1702 1439 1708 1440
rect 1702 1435 1703 1439
rect 1707 1435 1708 1439
rect 1702 1434 1708 1435
rect 1423 1426 1427 1427
rect 1423 1421 1427 1422
rect 1439 1426 1443 1427
rect 1439 1421 1443 1422
rect 1503 1426 1507 1427
rect 1503 1421 1507 1422
rect 1535 1426 1539 1427
rect 1535 1421 1539 1422
rect 1591 1426 1595 1427
rect 1631 1426 1635 1427
rect 1591 1421 1595 1422
rect 1602 1423 1608 1424
rect 1414 1415 1420 1416
rect 1414 1411 1415 1415
rect 1419 1411 1420 1415
rect 1414 1410 1420 1411
rect 1424 1402 1426 1421
rect 1504 1402 1506 1421
rect 1592 1402 1594 1421
rect 1602 1419 1603 1423
rect 1607 1419 1608 1423
rect 1631 1421 1635 1422
rect 1679 1426 1683 1427
rect 1679 1421 1683 1422
rect 1602 1418 1608 1419
rect 1366 1401 1372 1402
rect 1326 1400 1332 1401
rect 1326 1396 1327 1400
rect 1331 1396 1332 1400
rect 1366 1397 1367 1401
rect 1371 1397 1372 1401
rect 1422 1401 1428 1402
rect 1366 1396 1372 1397
rect 1374 1399 1380 1400
rect 1326 1395 1332 1396
rect 1374 1395 1375 1399
rect 1379 1395 1380 1399
rect 1422 1397 1423 1401
rect 1427 1397 1428 1401
rect 1422 1396 1428 1397
rect 1502 1401 1508 1402
rect 1502 1397 1503 1401
rect 1507 1397 1508 1401
rect 1502 1396 1508 1397
rect 1590 1401 1596 1402
rect 1590 1397 1591 1401
rect 1595 1397 1596 1401
rect 1590 1396 1596 1397
rect 1374 1394 1380 1395
rect 1326 1383 1332 1384
rect 511 1382 515 1383
rect 511 1377 515 1378
rect 527 1382 531 1383
rect 542 1382 548 1383
rect 607 1382 611 1383
rect 527 1377 531 1378
rect 607 1377 611 1378
rect 631 1382 635 1383
rect 631 1377 635 1378
rect 703 1382 707 1383
rect 703 1377 707 1378
rect 727 1382 731 1383
rect 727 1377 731 1378
rect 799 1382 803 1383
rect 799 1377 803 1378
rect 823 1382 827 1383
rect 823 1377 827 1378
rect 895 1382 899 1383
rect 911 1382 915 1383
rect 895 1377 899 1378
rect 902 1379 908 1380
rect 502 1371 508 1372
rect 502 1367 503 1371
rect 507 1367 508 1371
rect 502 1366 508 1367
rect 512 1358 514 1377
rect 608 1358 610 1377
rect 704 1358 706 1377
rect 800 1358 802 1377
rect 896 1358 898 1377
rect 902 1375 903 1379
rect 907 1375 908 1379
rect 911 1377 915 1378
rect 999 1382 1003 1383
rect 999 1377 1003 1378
rect 1007 1382 1011 1383
rect 1022 1382 1028 1383
rect 1103 1382 1107 1383
rect 1007 1377 1011 1378
rect 902 1374 908 1375
rect 150 1357 156 1358
rect 110 1356 116 1357
rect 110 1352 111 1356
rect 115 1352 116 1356
rect 150 1353 151 1357
rect 155 1353 156 1357
rect 214 1357 220 1358
rect 150 1352 156 1353
rect 158 1355 164 1356
rect 110 1351 116 1352
rect 158 1351 159 1355
rect 163 1351 164 1355
rect 214 1353 215 1357
rect 219 1353 220 1357
rect 214 1352 220 1353
rect 310 1357 316 1358
rect 310 1353 311 1357
rect 315 1353 316 1357
rect 310 1352 316 1353
rect 406 1357 412 1358
rect 406 1353 407 1357
rect 411 1353 412 1357
rect 406 1352 412 1353
rect 510 1357 516 1358
rect 510 1353 511 1357
rect 515 1353 516 1357
rect 510 1352 516 1353
rect 606 1357 612 1358
rect 606 1353 607 1357
rect 611 1353 612 1357
rect 606 1352 612 1353
rect 702 1357 708 1358
rect 702 1353 703 1357
rect 707 1353 708 1357
rect 702 1352 708 1353
rect 798 1357 804 1358
rect 798 1353 799 1357
rect 803 1353 804 1357
rect 798 1352 804 1353
rect 894 1357 900 1358
rect 894 1353 895 1357
rect 899 1353 900 1357
rect 894 1352 900 1353
rect 158 1350 164 1351
rect 110 1339 116 1340
rect 110 1335 111 1339
rect 115 1335 116 1339
rect 110 1334 116 1335
rect 134 1336 140 1337
rect 112 1331 114 1334
rect 134 1332 135 1336
rect 139 1332 140 1336
rect 134 1331 140 1332
rect 111 1330 115 1331
rect 111 1325 115 1326
rect 135 1330 139 1331
rect 135 1325 139 1326
rect 112 1322 114 1325
rect 134 1324 140 1325
rect 110 1321 116 1322
rect 110 1317 111 1321
rect 115 1317 116 1321
rect 134 1320 135 1324
rect 139 1320 140 1324
rect 134 1319 140 1320
rect 110 1316 116 1317
rect 110 1304 116 1305
rect 110 1300 111 1304
rect 115 1300 116 1304
rect 110 1299 116 1300
rect 150 1303 156 1304
rect 150 1299 151 1303
rect 155 1299 156 1303
rect 112 1279 114 1299
rect 150 1298 156 1299
rect 152 1279 154 1298
rect 160 1288 162 1350
rect 198 1336 204 1337
rect 198 1332 199 1336
rect 203 1332 204 1336
rect 198 1331 204 1332
rect 294 1336 300 1337
rect 294 1332 295 1336
rect 299 1332 300 1336
rect 294 1331 300 1332
rect 390 1336 396 1337
rect 390 1332 391 1336
rect 395 1332 396 1336
rect 390 1331 396 1332
rect 494 1336 500 1337
rect 494 1332 495 1336
rect 499 1332 500 1336
rect 494 1331 500 1332
rect 590 1336 596 1337
rect 590 1332 591 1336
rect 595 1332 596 1336
rect 590 1331 596 1332
rect 686 1336 692 1337
rect 686 1332 687 1336
rect 691 1332 692 1336
rect 686 1331 692 1332
rect 782 1336 788 1337
rect 782 1332 783 1336
rect 787 1332 788 1336
rect 782 1331 788 1332
rect 878 1336 884 1337
rect 878 1332 879 1336
rect 883 1332 884 1336
rect 878 1331 884 1332
rect 199 1330 203 1331
rect 199 1325 203 1326
rect 215 1330 219 1331
rect 215 1325 219 1326
rect 295 1330 299 1331
rect 295 1325 299 1326
rect 319 1330 323 1331
rect 319 1325 323 1326
rect 391 1330 395 1331
rect 391 1325 395 1326
rect 415 1330 419 1331
rect 415 1325 419 1326
rect 495 1330 499 1331
rect 495 1325 499 1326
rect 511 1330 515 1331
rect 511 1325 515 1326
rect 591 1330 595 1331
rect 591 1325 595 1326
rect 599 1330 603 1331
rect 599 1325 603 1326
rect 687 1330 691 1331
rect 687 1325 691 1326
rect 783 1330 787 1331
rect 783 1325 787 1326
rect 879 1330 883 1331
rect 879 1325 883 1326
rect 214 1324 220 1325
rect 214 1320 215 1324
rect 219 1320 220 1324
rect 214 1319 220 1320
rect 318 1324 324 1325
rect 318 1320 319 1324
rect 323 1320 324 1324
rect 318 1319 324 1320
rect 414 1324 420 1325
rect 414 1320 415 1324
rect 419 1320 420 1324
rect 414 1319 420 1320
rect 510 1324 516 1325
rect 510 1320 511 1324
rect 515 1320 516 1324
rect 510 1319 516 1320
rect 598 1324 604 1325
rect 598 1320 599 1324
rect 603 1320 604 1324
rect 598 1319 604 1320
rect 686 1324 692 1325
rect 686 1320 687 1324
rect 691 1320 692 1324
rect 686 1319 692 1320
rect 782 1324 788 1325
rect 782 1320 783 1324
rect 787 1320 788 1324
rect 782 1319 788 1320
rect 878 1324 884 1325
rect 878 1320 879 1324
rect 883 1320 884 1324
rect 878 1319 884 1320
rect 904 1304 906 1374
rect 1000 1358 1002 1377
rect 998 1357 1004 1358
rect 998 1353 999 1357
rect 1003 1353 1004 1357
rect 1024 1356 1026 1382
rect 1103 1377 1107 1378
rect 1287 1382 1291 1383
rect 1326 1379 1327 1383
rect 1331 1379 1332 1383
rect 1326 1378 1332 1379
rect 1350 1380 1356 1381
rect 1287 1377 1291 1378
rect 1288 1357 1290 1377
rect 1328 1371 1330 1378
rect 1350 1376 1351 1380
rect 1355 1376 1356 1380
rect 1350 1375 1356 1376
rect 1352 1371 1354 1375
rect 1327 1370 1331 1371
rect 1327 1365 1331 1366
rect 1351 1370 1355 1371
rect 1351 1365 1355 1366
rect 1328 1362 1330 1365
rect 1350 1364 1356 1365
rect 1326 1361 1332 1362
rect 1326 1357 1327 1361
rect 1331 1357 1332 1361
rect 1350 1360 1351 1364
rect 1355 1360 1356 1364
rect 1350 1359 1356 1360
rect 1286 1356 1292 1357
rect 1326 1356 1332 1357
rect 998 1352 1004 1353
rect 1022 1355 1028 1356
rect 1022 1351 1023 1355
rect 1027 1351 1028 1355
rect 1286 1352 1287 1356
rect 1291 1352 1292 1356
rect 1286 1351 1292 1352
rect 1022 1350 1028 1351
rect 1326 1344 1332 1345
rect 1326 1340 1327 1344
rect 1331 1340 1332 1344
rect 1286 1339 1292 1340
rect 1326 1339 1332 1340
rect 1366 1343 1372 1344
rect 1366 1339 1367 1343
rect 1371 1339 1372 1343
rect 982 1336 988 1337
rect 982 1332 983 1336
rect 987 1332 988 1336
rect 1286 1335 1287 1339
rect 1291 1335 1292 1339
rect 1286 1334 1292 1335
rect 982 1331 988 1332
rect 1288 1331 1290 1334
rect 983 1330 987 1331
rect 983 1325 987 1326
rect 1287 1330 1291 1331
rect 1287 1325 1291 1326
rect 1288 1322 1290 1325
rect 1286 1321 1292 1322
rect 1286 1317 1287 1321
rect 1291 1317 1292 1321
rect 1286 1316 1292 1317
rect 1328 1311 1330 1339
rect 1366 1338 1372 1339
rect 1368 1311 1370 1338
rect 1376 1328 1378 1394
rect 1406 1380 1412 1381
rect 1406 1376 1407 1380
rect 1411 1376 1412 1380
rect 1406 1375 1412 1376
rect 1486 1380 1492 1381
rect 1486 1376 1487 1380
rect 1491 1376 1492 1380
rect 1486 1375 1492 1376
rect 1574 1380 1580 1381
rect 1574 1376 1575 1380
rect 1579 1376 1580 1380
rect 1574 1375 1580 1376
rect 1408 1371 1410 1375
rect 1488 1371 1490 1375
rect 1576 1371 1578 1375
rect 1407 1370 1411 1371
rect 1407 1365 1411 1366
rect 1479 1370 1483 1371
rect 1479 1365 1483 1366
rect 1487 1370 1491 1371
rect 1487 1365 1491 1366
rect 1567 1370 1571 1371
rect 1567 1365 1571 1366
rect 1575 1370 1579 1371
rect 1575 1365 1579 1366
rect 1406 1364 1412 1365
rect 1406 1360 1407 1364
rect 1411 1360 1412 1364
rect 1406 1359 1412 1360
rect 1478 1364 1484 1365
rect 1478 1360 1479 1364
rect 1483 1360 1484 1364
rect 1478 1359 1484 1360
rect 1566 1364 1572 1365
rect 1566 1360 1567 1364
rect 1571 1360 1572 1364
rect 1566 1359 1572 1360
rect 1604 1344 1606 1418
rect 1680 1402 1682 1421
rect 1678 1401 1684 1402
rect 1678 1397 1679 1401
rect 1683 1397 1684 1401
rect 1704 1400 1706 1434
rect 1728 1427 1730 1450
rect 1832 1427 1834 1450
rect 1727 1426 1731 1427
rect 1727 1421 1731 1422
rect 1775 1426 1779 1427
rect 1775 1421 1779 1422
rect 1831 1426 1835 1427
rect 1840 1424 1842 1450
rect 1944 1427 1946 1450
rect 1960 1436 1962 1450
rect 1958 1435 1964 1436
rect 1958 1431 1959 1435
rect 1963 1431 1964 1435
rect 1958 1430 1964 1431
rect 2064 1427 2066 1450
rect 2144 1440 2146 1506
rect 2230 1492 2236 1493
rect 2230 1488 2231 1492
rect 2235 1488 2236 1492
rect 2230 1487 2236 1488
rect 2326 1492 2332 1493
rect 2326 1488 2327 1492
rect 2331 1488 2332 1492
rect 2326 1487 2332 1488
rect 2232 1483 2234 1487
rect 2328 1483 2330 1487
rect 2175 1482 2179 1483
rect 2175 1477 2179 1478
rect 2231 1482 2235 1483
rect 2231 1477 2235 1478
rect 2303 1482 2307 1483
rect 2303 1477 2307 1478
rect 2327 1482 2331 1483
rect 2327 1477 2331 1478
rect 2174 1476 2180 1477
rect 2174 1472 2175 1476
rect 2179 1472 2180 1476
rect 2174 1471 2180 1472
rect 2302 1476 2308 1477
rect 2302 1472 2303 1476
rect 2307 1472 2308 1476
rect 2302 1471 2308 1472
rect 2352 1456 2354 1522
rect 2364 1512 2366 1530
rect 2440 1514 2442 1533
rect 2472 1528 2474 1558
rect 2504 1539 2506 1559
rect 2503 1538 2507 1539
rect 2503 1533 2507 1534
rect 2470 1527 2476 1528
rect 2470 1523 2471 1527
rect 2475 1523 2476 1527
rect 2470 1522 2476 1523
rect 2438 1513 2444 1514
rect 2504 1513 2506 1533
rect 2362 1511 2368 1512
rect 2362 1507 2363 1511
rect 2367 1507 2368 1511
rect 2438 1509 2439 1513
rect 2443 1509 2444 1513
rect 2502 1512 2508 1513
rect 2438 1508 2444 1509
rect 2462 1511 2468 1512
rect 2362 1506 2368 1507
rect 2462 1507 2463 1511
rect 2467 1507 2468 1511
rect 2502 1508 2503 1512
rect 2507 1508 2508 1512
rect 2502 1507 2508 1508
rect 2462 1506 2468 1507
rect 2422 1492 2428 1493
rect 2422 1488 2423 1492
rect 2427 1488 2428 1492
rect 2422 1487 2428 1488
rect 2424 1483 2426 1487
rect 2423 1482 2427 1483
rect 2423 1477 2427 1478
rect 2439 1482 2443 1483
rect 2439 1477 2443 1478
rect 2438 1476 2444 1477
rect 2438 1472 2439 1476
rect 2443 1472 2444 1476
rect 2438 1471 2444 1472
rect 2190 1455 2196 1456
rect 2190 1451 2191 1455
rect 2195 1451 2196 1455
rect 2190 1450 2196 1451
rect 2318 1455 2324 1456
rect 2318 1451 2319 1455
rect 2323 1451 2324 1455
rect 2318 1450 2324 1451
rect 2350 1455 2356 1456
rect 2350 1451 2351 1455
rect 2355 1451 2356 1455
rect 2350 1450 2356 1451
rect 2454 1455 2460 1456
rect 2454 1451 2455 1455
rect 2459 1451 2460 1455
rect 2454 1450 2460 1451
rect 2142 1439 2148 1440
rect 2142 1435 2143 1439
rect 2147 1435 2148 1439
rect 2142 1434 2148 1435
rect 2192 1427 2194 1450
rect 2254 1439 2260 1440
rect 2254 1435 2255 1439
rect 2259 1435 2260 1439
rect 2254 1434 2260 1435
rect 1879 1426 1883 1427
rect 1831 1421 1835 1422
rect 1838 1423 1844 1424
rect 1776 1402 1778 1421
rect 1838 1419 1839 1423
rect 1843 1419 1844 1423
rect 1879 1421 1883 1422
rect 1943 1426 1947 1427
rect 1943 1421 1947 1422
rect 1991 1426 1995 1427
rect 1991 1421 1995 1422
rect 2063 1426 2067 1427
rect 2063 1421 2067 1422
rect 2111 1426 2115 1427
rect 2111 1421 2115 1422
rect 2191 1426 2195 1427
rect 2191 1421 2195 1422
rect 2231 1426 2235 1427
rect 2231 1421 2235 1422
rect 1838 1418 1844 1419
rect 1880 1402 1882 1421
rect 1992 1402 1994 1421
rect 2112 1402 2114 1421
rect 2232 1402 2234 1421
rect 1774 1401 1780 1402
rect 1678 1396 1684 1397
rect 1702 1399 1708 1400
rect 1702 1395 1703 1399
rect 1707 1395 1708 1399
rect 1774 1397 1775 1401
rect 1779 1397 1780 1401
rect 1774 1396 1780 1397
rect 1878 1401 1884 1402
rect 1878 1397 1879 1401
rect 1883 1397 1884 1401
rect 1878 1396 1884 1397
rect 1990 1401 1996 1402
rect 1990 1397 1991 1401
rect 1995 1397 1996 1401
rect 1990 1396 1996 1397
rect 2110 1401 2116 1402
rect 2110 1397 2111 1401
rect 2115 1397 2116 1401
rect 2230 1401 2236 1402
rect 2110 1396 2116 1397
rect 2118 1399 2124 1400
rect 1702 1394 1708 1395
rect 2118 1395 2119 1399
rect 2123 1395 2124 1399
rect 2230 1397 2231 1401
rect 2235 1397 2236 1401
rect 2256 1400 2258 1434
rect 2320 1427 2322 1450
rect 2456 1427 2458 1450
rect 2464 1440 2466 1506
rect 2502 1495 2508 1496
rect 2502 1491 2503 1495
rect 2507 1491 2508 1495
rect 2502 1490 2508 1491
rect 2504 1483 2506 1490
rect 2503 1482 2507 1483
rect 2503 1477 2507 1478
rect 2504 1474 2506 1477
rect 2502 1473 2508 1474
rect 2502 1469 2503 1473
rect 2507 1469 2508 1473
rect 2502 1468 2508 1469
rect 2502 1456 2508 1457
rect 2470 1455 2476 1456
rect 2470 1451 2471 1455
rect 2475 1451 2476 1455
rect 2502 1452 2503 1456
rect 2507 1452 2508 1456
rect 2502 1451 2508 1452
rect 2470 1450 2476 1451
rect 2462 1439 2468 1440
rect 2462 1435 2463 1439
rect 2467 1435 2468 1439
rect 2462 1434 2468 1435
rect 2319 1426 2323 1427
rect 2319 1421 2323 1422
rect 2351 1426 2355 1427
rect 2351 1421 2355 1422
rect 2455 1426 2459 1427
rect 2455 1421 2459 1422
rect 2352 1402 2354 1421
rect 2358 1415 2364 1416
rect 2358 1411 2359 1415
rect 2363 1411 2364 1415
rect 2358 1410 2364 1411
rect 2350 1401 2356 1402
rect 2230 1396 2236 1397
rect 2254 1399 2260 1400
rect 2118 1394 2124 1395
rect 2254 1395 2255 1399
rect 2259 1395 2260 1399
rect 2350 1397 2351 1401
rect 2355 1397 2356 1401
rect 2350 1396 2356 1397
rect 2254 1394 2260 1395
rect 1662 1380 1668 1381
rect 1662 1376 1663 1380
rect 1667 1376 1668 1380
rect 1662 1375 1668 1376
rect 1758 1380 1764 1381
rect 1758 1376 1759 1380
rect 1763 1376 1764 1380
rect 1758 1375 1764 1376
rect 1862 1380 1868 1381
rect 1862 1376 1863 1380
rect 1867 1376 1868 1380
rect 1862 1375 1868 1376
rect 1974 1380 1980 1381
rect 1974 1376 1975 1380
rect 1979 1376 1980 1380
rect 1974 1375 1980 1376
rect 2094 1380 2100 1381
rect 2094 1376 2095 1380
rect 2099 1376 2100 1380
rect 2094 1375 2100 1376
rect 1664 1371 1666 1375
rect 1760 1371 1762 1375
rect 1864 1371 1866 1375
rect 1976 1371 1978 1375
rect 2096 1371 2098 1375
rect 1655 1370 1659 1371
rect 1655 1365 1659 1366
rect 1663 1370 1667 1371
rect 1663 1365 1667 1366
rect 1751 1370 1755 1371
rect 1751 1365 1755 1366
rect 1759 1370 1763 1371
rect 1759 1365 1763 1366
rect 1855 1370 1859 1371
rect 1855 1365 1859 1366
rect 1863 1370 1867 1371
rect 1863 1365 1867 1366
rect 1967 1370 1971 1371
rect 1967 1365 1971 1366
rect 1975 1370 1979 1371
rect 1975 1365 1979 1366
rect 2079 1370 2083 1371
rect 2079 1365 2083 1366
rect 2095 1370 2099 1371
rect 2095 1365 2099 1366
rect 1654 1364 1660 1365
rect 1654 1360 1655 1364
rect 1659 1360 1660 1364
rect 1654 1359 1660 1360
rect 1750 1364 1756 1365
rect 1750 1360 1751 1364
rect 1755 1360 1756 1364
rect 1750 1359 1756 1360
rect 1854 1364 1860 1365
rect 1854 1360 1855 1364
rect 1859 1360 1860 1364
rect 1854 1359 1860 1360
rect 1966 1364 1972 1365
rect 1966 1360 1967 1364
rect 1971 1360 1972 1364
rect 1966 1359 1972 1360
rect 2078 1364 2084 1365
rect 2078 1360 2079 1364
rect 2083 1360 2084 1364
rect 2078 1359 2084 1360
rect 1422 1343 1428 1344
rect 1422 1339 1423 1343
rect 1427 1339 1428 1343
rect 1422 1338 1428 1339
rect 1494 1343 1500 1344
rect 1494 1339 1495 1343
rect 1499 1339 1500 1343
rect 1494 1338 1500 1339
rect 1526 1343 1532 1344
rect 1526 1339 1527 1343
rect 1531 1339 1532 1343
rect 1526 1338 1532 1339
rect 1582 1343 1588 1344
rect 1582 1339 1583 1343
rect 1587 1339 1588 1343
rect 1582 1338 1588 1339
rect 1602 1343 1608 1344
rect 1602 1339 1603 1343
rect 1607 1339 1608 1343
rect 1602 1338 1608 1339
rect 1670 1343 1676 1344
rect 1670 1339 1671 1343
rect 1675 1339 1676 1343
rect 1670 1338 1676 1339
rect 1766 1343 1772 1344
rect 1766 1339 1767 1343
rect 1771 1339 1772 1343
rect 1766 1338 1772 1339
rect 1870 1343 1876 1344
rect 1870 1339 1871 1343
rect 1875 1339 1876 1343
rect 1870 1338 1876 1339
rect 1982 1343 1988 1344
rect 1982 1339 1983 1343
rect 1987 1339 1988 1343
rect 1982 1338 1988 1339
rect 2094 1343 2100 1344
rect 2094 1339 2095 1343
rect 2099 1339 2100 1343
rect 2094 1338 2100 1339
rect 1374 1327 1380 1328
rect 1374 1323 1375 1327
rect 1379 1323 1380 1327
rect 1374 1322 1380 1323
rect 1424 1311 1426 1338
rect 1496 1311 1498 1338
rect 1327 1310 1331 1311
rect 1327 1305 1331 1306
rect 1367 1310 1371 1311
rect 1367 1305 1371 1306
rect 1423 1310 1427 1311
rect 1423 1305 1427 1306
rect 1495 1310 1499 1311
rect 1495 1305 1499 1306
rect 1519 1310 1523 1311
rect 1519 1305 1523 1306
rect 1286 1304 1292 1305
rect 230 1303 236 1304
rect 230 1299 231 1303
rect 235 1299 236 1303
rect 230 1298 236 1299
rect 334 1303 340 1304
rect 334 1299 335 1303
rect 339 1299 340 1303
rect 334 1298 340 1299
rect 430 1303 436 1304
rect 430 1299 431 1303
rect 435 1299 436 1303
rect 430 1298 436 1299
rect 446 1303 452 1304
rect 446 1299 447 1303
rect 451 1299 452 1303
rect 446 1298 452 1299
rect 526 1303 532 1304
rect 526 1299 527 1303
rect 531 1299 532 1303
rect 526 1298 532 1299
rect 614 1303 620 1304
rect 614 1299 615 1303
rect 619 1299 620 1303
rect 614 1298 620 1299
rect 702 1303 708 1304
rect 702 1299 703 1303
rect 707 1299 708 1303
rect 702 1298 708 1299
rect 798 1303 804 1304
rect 798 1299 799 1303
rect 803 1299 804 1303
rect 798 1298 804 1299
rect 894 1303 900 1304
rect 894 1299 895 1303
rect 899 1299 900 1303
rect 894 1298 900 1299
rect 902 1303 908 1304
rect 902 1299 903 1303
rect 907 1299 908 1303
rect 1286 1300 1287 1304
rect 1291 1300 1292 1304
rect 1286 1299 1292 1300
rect 902 1298 908 1299
rect 158 1287 164 1288
rect 158 1283 159 1287
rect 163 1283 164 1287
rect 158 1282 164 1283
rect 232 1279 234 1298
rect 336 1279 338 1298
rect 432 1279 434 1298
rect 111 1278 115 1279
rect 111 1273 115 1274
rect 151 1278 155 1279
rect 151 1273 155 1274
rect 191 1278 195 1279
rect 191 1273 195 1274
rect 231 1278 235 1279
rect 231 1273 235 1274
rect 247 1278 251 1279
rect 247 1273 251 1274
rect 303 1278 307 1279
rect 303 1273 307 1274
rect 335 1278 339 1279
rect 335 1273 339 1274
rect 367 1278 371 1279
rect 367 1273 371 1274
rect 431 1278 435 1279
rect 431 1273 435 1274
rect 439 1278 443 1279
rect 448 1276 450 1298
rect 528 1279 530 1298
rect 616 1279 618 1298
rect 704 1279 706 1298
rect 800 1279 802 1298
rect 896 1279 898 1298
rect 1246 1291 1252 1292
rect 1246 1287 1247 1291
rect 1251 1287 1252 1291
rect 1246 1286 1252 1287
rect 1114 1283 1120 1284
rect 1114 1279 1115 1283
rect 1119 1279 1120 1283
rect 527 1278 531 1279
rect 439 1273 443 1274
rect 446 1275 452 1276
rect 112 1253 114 1273
rect 192 1254 194 1273
rect 248 1254 250 1273
rect 304 1254 306 1273
rect 368 1254 370 1273
rect 440 1254 442 1273
rect 446 1271 447 1275
rect 451 1271 452 1275
rect 527 1273 531 1274
rect 615 1278 619 1279
rect 615 1273 619 1274
rect 639 1278 643 1279
rect 639 1273 643 1274
rect 703 1278 707 1279
rect 703 1273 707 1274
rect 775 1278 779 1279
rect 775 1273 779 1274
rect 799 1278 803 1279
rect 799 1273 803 1274
rect 895 1278 899 1279
rect 895 1273 899 1274
rect 927 1278 931 1279
rect 927 1273 931 1274
rect 1095 1278 1099 1279
rect 1114 1278 1120 1279
rect 1239 1278 1243 1279
rect 1095 1273 1099 1274
rect 446 1270 452 1271
rect 528 1254 530 1273
rect 640 1254 642 1273
rect 654 1267 660 1268
rect 654 1263 655 1267
rect 659 1263 660 1267
rect 654 1262 660 1263
rect 190 1253 196 1254
rect 110 1252 116 1253
rect 110 1248 111 1252
rect 115 1248 116 1252
rect 190 1249 191 1253
rect 195 1249 196 1253
rect 190 1248 196 1249
rect 246 1253 252 1254
rect 246 1249 247 1253
rect 251 1249 252 1253
rect 246 1248 252 1249
rect 302 1253 308 1254
rect 302 1249 303 1253
rect 307 1249 308 1253
rect 302 1248 308 1249
rect 366 1253 372 1254
rect 366 1249 367 1253
rect 371 1249 372 1253
rect 366 1248 372 1249
rect 438 1253 444 1254
rect 438 1249 439 1253
rect 443 1249 444 1253
rect 438 1248 444 1249
rect 526 1253 532 1254
rect 526 1249 527 1253
rect 531 1249 532 1253
rect 638 1253 644 1254
rect 526 1248 532 1249
rect 550 1251 556 1252
rect 110 1247 116 1248
rect 550 1247 551 1251
rect 555 1247 556 1251
rect 638 1249 639 1253
rect 643 1249 644 1253
rect 638 1248 644 1249
rect 550 1246 556 1247
rect 110 1235 116 1236
rect 110 1231 111 1235
rect 115 1231 116 1235
rect 110 1230 116 1231
rect 174 1232 180 1233
rect 112 1227 114 1230
rect 174 1228 175 1232
rect 179 1228 180 1232
rect 174 1227 180 1228
rect 230 1232 236 1233
rect 230 1228 231 1232
rect 235 1228 236 1232
rect 230 1227 236 1228
rect 286 1232 292 1233
rect 286 1228 287 1232
rect 291 1228 292 1232
rect 286 1227 292 1228
rect 350 1232 356 1233
rect 350 1228 351 1232
rect 355 1228 356 1232
rect 350 1227 356 1228
rect 422 1232 428 1233
rect 422 1228 423 1232
rect 427 1228 428 1232
rect 422 1227 428 1228
rect 510 1232 516 1233
rect 510 1228 511 1232
rect 515 1228 516 1232
rect 510 1227 516 1228
rect 111 1226 115 1227
rect 111 1221 115 1222
rect 175 1226 179 1227
rect 175 1221 179 1222
rect 231 1226 235 1227
rect 231 1221 235 1222
rect 287 1226 291 1227
rect 287 1221 291 1222
rect 351 1226 355 1227
rect 351 1221 355 1222
rect 407 1226 411 1227
rect 407 1221 411 1222
rect 423 1226 427 1227
rect 423 1221 427 1222
rect 463 1226 467 1227
rect 463 1221 467 1222
rect 511 1226 515 1227
rect 511 1221 515 1222
rect 519 1226 523 1227
rect 519 1221 523 1222
rect 112 1218 114 1221
rect 350 1220 356 1221
rect 110 1217 116 1218
rect 110 1213 111 1217
rect 115 1213 116 1217
rect 350 1216 351 1220
rect 355 1216 356 1220
rect 350 1215 356 1216
rect 406 1220 412 1221
rect 406 1216 407 1220
rect 411 1216 412 1220
rect 406 1215 412 1216
rect 462 1220 468 1221
rect 462 1216 463 1220
rect 467 1216 468 1220
rect 462 1215 468 1216
rect 518 1220 524 1221
rect 518 1216 519 1220
rect 523 1216 524 1220
rect 518 1215 524 1216
rect 110 1212 116 1213
rect 110 1200 116 1201
rect 110 1196 111 1200
rect 115 1196 116 1200
rect 110 1195 116 1196
rect 366 1199 372 1200
rect 366 1195 367 1199
rect 371 1195 372 1199
rect 112 1171 114 1195
rect 366 1194 372 1195
rect 422 1199 428 1200
rect 422 1195 423 1199
rect 427 1195 428 1199
rect 422 1194 428 1195
rect 478 1199 484 1200
rect 478 1195 479 1199
rect 483 1195 484 1199
rect 478 1194 484 1195
rect 534 1199 540 1200
rect 534 1195 535 1199
rect 539 1195 540 1199
rect 534 1194 540 1195
rect 368 1171 370 1194
rect 424 1171 426 1194
rect 480 1171 482 1194
rect 536 1171 538 1194
rect 552 1180 554 1246
rect 622 1232 628 1233
rect 622 1228 623 1232
rect 627 1228 628 1232
rect 622 1227 628 1228
rect 575 1226 579 1227
rect 575 1221 579 1222
rect 623 1226 627 1227
rect 623 1221 627 1222
rect 631 1226 635 1227
rect 631 1221 635 1222
rect 574 1220 580 1221
rect 574 1216 575 1220
rect 579 1216 580 1220
rect 574 1215 580 1216
rect 630 1220 636 1221
rect 630 1216 631 1220
rect 635 1216 636 1220
rect 630 1215 636 1216
rect 656 1200 658 1262
rect 776 1254 778 1273
rect 928 1254 930 1273
rect 1096 1254 1098 1273
rect 774 1253 780 1254
rect 774 1249 775 1253
rect 779 1249 780 1253
rect 774 1248 780 1249
rect 926 1253 932 1254
rect 926 1249 927 1253
rect 931 1249 932 1253
rect 926 1248 932 1249
rect 1094 1253 1100 1254
rect 1094 1249 1095 1253
rect 1099 1249 1100 1253
rect 1116 1252 1118 1278
rect 1239 1273 1243 1274
rect 1240 1254 1242 1273
rect 1248 1268 1250 1286
rect 1288 1279 1290 1299
rect 1328 1285 1330 1305
rect 1368 1286 1370 1305
rect 1424 1286 1426 1305
rect 1520 1286 1522 1305
rect 1528 1300 1530 1338
rect 1584 1311 1586 1338
rect 1672 1311 1674 1338
rect 1742 1327 1748 1328
rect 1742 1323 1743 1327
rect 1747 1323 1748 1327
rect 1742 1322 1748 1323
rect 1583 1310 1587 1311
rect 1583 1305 1587 1306
rect 1615 1310 1619 1311
rect 1615 1305 1619 1306
rect 1671 1310 1675 1311
rect 1671 1305 1675 1306
rect 1719 1310 1723 1311
rect 1719 1305 1723 1306
rect 1526 1299 1532 1300
rect 1526 1295 1527 1299
rect 1531 1295 1532 1299
rect 1526 1294 1532 1295
rect 1616 1286 1618 1305
rect 1720 1286 1722 1305
rect 1366 1285 1372 1286
rect 1326 1284 1332 1285
rect 1326 1280 1327 1284
rect 1331 1280 1332 1284
rect 1366 1281 1367 1285
rect 1371 1281 1372 1285
rect 1366 1280 1372 1281
rect 1422 1285 1428 1286
rect 1422 1281 1423 1285
rect 1427 1281 1428 1285
rect 1422 1280 1428 1281
rect 1518 1285 1524 1286
rect 1518 1281 1519 1285
rect 1523 1281 1524 1285
rect 1518 1280 1524 1281
rect 1614 1285 1620 1286
rect 1614 1281 1615 1285
rect 1619 1281 1620 1285
rect 1614 1280 1620 1281
rect 1718 1285 1724 1286
rect 1718 1281 1719 1285
rect 1723 1281 1724 1285
rect 1744 1284 1746 1322
rect 1768 1311 1770 1338
rect 1872 1311 1874 1338
rect 1984 1311 1986 1338
rect 2096 1311 2098 1338
rect 2120 1324 2122 1394
rect 2214 1380 2220 1381
rect 2214 1376 2215 1380
rect 2219 1376 2220 1380
rect 2214 1375 2220 1376
rect 2334 1380 2340 1381
rect 2334 1376 2335 1380
rect 2339 1376 2340 1380
rect 2334 1375 2340 1376
rect 2216 1371 2218 1375
rect 2336 1371 2338 1375
rect 2199 1370 2203 1371
rect 2199 1365 2203 1366
rect 2215 1370 2219 1371
rect 2215 1365 2219 1366
rect 2327 1370 2331 1371
rect 2327 1365 2331 1366
rect 2335 1370 2339 1371
rect 2335 1365 2339 1366
rect 2198 1364 2204 1365
rect 2198 1360 2199 1364
rect 2203 1360 2204 1364
rect 2198 1359 2204 1360
rect 2326 1364 2332 1365
rect 2326 1360 2327 1364
rect 2331 1360 2332 1364
rect 2326 1359 2332 1360
rect 2360 1344 2362 1410
rect 2456 1402 2458 1421
rect 2472 1416 2474 1450
rect 2504 1427 2506 1451
rect 2503 1426 2507 1427
rect 2503 1421 2507 1422
rect 2470 1415 2476 1416
rect 2470 1411 2471 1415
rect 2475 1411 2476 1415
rect 2470 1410 2476 1411
rect 2454 1401 2460 1402
rect 2504 1401 2506 1421
rect 2454 1397 2455 1401
rect 2459 1397 2460 1401
rect 2502 1400 2508 1401
rect 2454 1396 2460 1397
rect 2462 1399 2468 1400
rect 2462 1395 2463 1399
rect 2467 1395 2468 1399
rect 2502 1396 2503 1400
rect 2507 1396 2508 1400
rect 2502 1395 2508 1396
rect 2462 1394 2468 1395
rect 2438 1380 2444 1381
rect 2438 1376 2439 1380
rect 2443 1376 2444 1380
rect 2438 1375 2444 1376
rect 2440 1371 2442 1375
rect 2439 1370 2443 1371
rect 2439 1365 2443 1366
rect 2438 1364 2444 1365
rect 2438 1360 2439 1364
rect 2443 1360 2444 1364
rect 2438 1359 2444 1360
rect 2214 1343 2220 1344
rect 2214 1339 2215 1343
rect 2219 1339 2220 1343
rect 2214 1338 2220 1339
rect 2222 1343 2228 1344
rect 2222 1339 2223 1343
rect 2227 1339 2228 1343
rect 2222 1338 2228 1339
rect 2342 1343 2348 1344
rect 2342 1339 2343 1343
rect 2347 1339 2348 1343
rect 2342 1338 2348 1339
rect 2358 1343 2364 1344
rect 2358 1339 2359 1343
rect 2363 1339 2364 1343
rect 2358 1338 2364 1339
rect 2454 1343 2460 1344
rect 2454 1339 2455 1343
rect 2459 1339 2460 1343
rect 2454 1338 2460 1339
rect 2118 1323 2124 1324
rect 2118 1319 2119 1323
rect 2123 1319 2124 1323
rect 2118 1318 2124 1319
rect 2216 1311 2218 1338
rect 1767 1310 1771 1311
rect 1767 1305 1771 1306
rect 1823 1310 1827 1311
rect 1871 1310 1875 1311
rect 1823 1305 1827 1306
rect 1842 1307 1848 1308
rect 1824 1286 1826 1305
rect 1842 1303 1843 1307
rect 1847 1303 1848 1307
rect 1871 1305 1875 1306
rect 1919 1310 1923 1311
rect 1919 1305 1923 1306
rect 1983 1310 1987 1311
rect 1983 1305 1987 1306
rect 2015 1310 2019 1311
rect 2015 1305 2019 1306
rect 2095 1310 2099 1311
rect 2095 1305 2099 1306
rect 2103 1310 2107 1311
rect 2103 1305 2107 1306
rect 2183 1310 2187 1311
rect 2183 1305 2187 1306
rect 2215 1310 2219 1311
rect 2224 1308 2226 1338
rect 2344 1311 2346 1338
rect 2350 1327 2356 1328
rect 2350 1323 2351 1327
rect 2355 1323 2356 1327
rect 2350 1322 2356 1323
rect 2255 1310 2259 1311
rect 2215 1305 2219 1306
rect 2222 1307 2228 1308
rect 1842 1302 1848 1303
rect 1822 1285 1828 1286
rect 1718 1280 1724 1281
rect 1742 1283 1748 1284
rect 1326 1279 1332 1280
rect 1742 1279 1743 1283
rect 1747 1279 1748 1283
rect 1822 1281 1823 1285
rect 1827 1281 1828 1285
rect 1844 1284 1846 1302
rect 1850 1299 1856 1300
rect 1850 1295 1851 1299
rect 1855 1295 1856 1299
rect 1850 1294 1856 1295
rect 1822 1280 1828 1281
rect 1842 1283 1848 1284
rect 1287 1278 1291 1279
rect 1742 1278 1748 1279
rect 1842 1279 1843 1283
rect 1847 1279 1848 1283
rect 1842 1278 1848 1279
rect 1287 1273 1291 1274
rect 1246 1267 1252 1268
rect 1246 1263 1247 1267
rect 1251 1263 1252 1267
rect 1246 1262 1252 1263
rect 1238 1253 1244 1254
rect 1288 1253 1290 1273
rect 1326 1267 1332 1268
rect 1326 1263 1327 1267
rect 1331 1263 1332 1267
rect 1326 1262 1332 1263
rect 1350 1264 1356 1265
rect 1094 1248 1100 1249
rect 1114 1251 1120 1252
rect 1114 1247 1115 1251
rect 1119 1247 1120 1251
rect 1238 1249 1239 1253
rect 1243 1249 1244 1253
rect 1286 1252 1292 1253
rect 1238 1248 1244 1249
rect 1278 1251 1284 1252
rect 1114 1246 1120 1247
rect 1278 1247 1279 1251
rect 1283 1247 1284 1251
rect 1286 1248 1287 1252
rect 1291 1248 1292 1252
rect 1286 1247 1292 1248
rect 1278 1246 1284 1247
rect 758 1232 764 1233
rect 758 1228 759 1232
rect 763 1228 764 1232
rect 758 1227 764 1228
rect 910 1232 916 1233
rect 910 1228 911 1232
rect 915 1228 916 1232
rect 910 1227 916 1228
rect 1078 1232 1084 1233
rect 1078 1228 1079 1232
rect 1083 1228 1084 1232
rect 1078 1227 1084 1228
rect 1222 1232 1228 1233
rect 1222 1228 1223 1232
rect 1227 1228 1228 1232
rect 1222 1227 1228 1228
rect 687 1226 691 1227
rect 687 1221 691 1222
rect 743 1226 747 1227
rect 743 1221 747 1222
rect 759 1226 763 1227
rect 759 1221 763 1222
rect 799 1226 803 1227
rect 799 1221 803 1222
rect 855 1226 859 1227
rect 855 1221 859 1222
rect 911 1226 915 1227
rect 911 1221 915 1222
rect 1079 1226 1083 1227
rect 1079 1221 1083 1222
rect 1223 1226 1227 1227
rect 1223 1221 1227 1222
rect 686 1220 692 1221
rect 686 1216 687 1220
rect 691 1216 692 1220
rect 686 1215 692 1216
rect 742 1220 748 1221
rect 742 1216 743 1220
rect 747 1216 748 1220
rect 742 1215 748 1216
rect 798 1220 804 1221
rect 798 1216 799 1220
rect 803 1216 804 1220
rect 798 1215 804 1216
rect 854 1220 860 1221
rect 854 1216 855 1220
rect 859 1216 860 1220
rect 854 1215 860 1216
rect 910 1220 916 1221
rect 910 1216 911 1220
rect 915 1216 916 1220
rect 910 1215 916 1216
rect 1280 1208 1282 1246
rect 1328 1243 1330 1262
rect 1350 1260 1351 1264
rect 1355 1260 1356 1264
rect 1350 1259 1356 1260
rect 1406 1264 1412 1265
rect 1406 1260 1407 1264
rect 1411 1260 1412 1264
rect 1406 1259 1412 1260
rect 1502 1264 1508 1265
rect 1502 1260 1503 1264
rect 1507 1260 1508 1264
rect 1502 1259 1508 1260
rect 1598 1264 1604 1265
rect 1598 1260 1599 1264
rect 1603 1260 1604 1264
rect 1598 1259 1604 1260
rect 1702 1264 1708 1265
rect 1702 1260 1703 1264
rect 1707 1260 1708 1264
rect 1702 1259 1708 1260
rect 1806 1264 1812 1265
rect 1806 1260 1807 1264
rect 1811 1260 1812 1264
rect 1806 1259 1812 1260
rect 1352 1243 1354 1259
rect 1408 1243 1410 1259
rect 1504 1243 1506 1259
rect 1600 1243 1602 1259
rect 1704 1243 1706 1259
rect 1808 1243 1810 1259
rect 1327 1242 1331 1243
rect 1327 1237 1331 1238
rect 1351 1242 1355 1243
rect 1351 1237 1355 1238
rect 1407 1242 1411 1243
rect 1407 1237 1411 1238
rect 1447 1242 1451 1243
rect 1447 1237 1451 1238
rect 1503 1242 1507 1243
rect 1503 1237 1507 1238
rect 1575 1242 1579 1243
rect 1575 1237 1579 1238
rect 1599 1242 1603 1243
rect 1599 1237 1603 1238
rect 1695 1242 1699 1243
rect 1695 1237 1699 1238
rect 1703 1242 1707 1243
rect 1703 1237 1707 1238
rect 1807 1242 1811 1243
rect 1807 1237 1811 1238
rect 1815 1242 1819 1243
rect 1815 1237 1819 1238
rect 1286 1235 1292 1236
rect 1286 1231 1287 1235
rect 1291 1231 1292 1235
rect 1328 1234 1330 1237
rect 1350 1236 1356 1237
rect 1286 1230 1292 1231
rect 1326 1233 1332 1234
rect 1288 1227 1290 1230
rect 1326 1229 1327 1233
rect 1331 1229 1332 1233
rect 1350 1232 1351 1236
rect 1355 1232 1356 1236
rect 1350 1231 1356 1232
rect 1446 1236 1452 1237
rect 1446 1232 1447 1236
rect 1451 1232 1452 1236
rect 1446 1231 1452 1232
rect 1574 1236 1580 1237
rect 1574 1232 1575 1236
rect 1579 1232 1580 1236
rect 1574 1231 1580 1232
rect 1694 1236 1700 1237
rect 1694 1232 1695 1236
rect 1699 1232 1700 1236
rect 1694 1231 1700 1232
rect 1814 1236 1820 1237
rect 1814 1232 1815 1236
rect 1819 1232 1820 1236
rect 1814 1231 1820 1232
rect 1326 1228 1332 1229
rect 1287 1226 1291 1227
rect 1287 1221 1291 1222
rect 1288 1218 1290 1221
rect 1286 1217 1292 1218
rect 1286 1213 1287 1217
rect 1291 1213 1292 1217
rect 1286 1212 1292 1213
rect 1326 1216 1332 1217
rect 1852 1216 1854 1294
rect 1920 1286 1922 1305
rect 2016 1286 2018 1305
rect 2104 1286 2106 1305
rect 2184 1286 2186 1305
rect 2222 1303 2223 1307
rect 2227 1303 2228 1307
rect 2255 1305 2259 1306
rect 2327 1310 2331 1311
rect 2327 1305 2331 1306
rect 2343 1310 2347 1311
rect 2343 1305 2347 1306
rect 2222 1302 2228 1303
rect 2256 1286 2258 1305
rect 2328 1286 2330 1305
rect 1918 1285 1924 1286
rect 1918 1281 1919 1285
rect 1923 1281 1924 1285
rect 1918 1280 1924 1281
rect 2014 1285 2020 1286
rect 2014 1281 2015 1285
rect 2019 1281 2020 1285
rect 2014 1280 2020 1281
rect 2102 1285 2108 1286
rect 2102 1281 2103 1285
rect 2107 1281 2108 1285
rect 2102 1280 2108 1281
rect 2182 1285 2188 1286
rect 2182 1281 2183 1285
rect 2187 1281 2188 1285
rect 2182 1280 2188 1281
rect 2254 1285 2260 1286
rect 2254 1281 2255 1285
rect 2259 1281 2260 1285
rect 2326 1285 2332 1286
rect 2254 1280 2260 1281
rect 2262 1283 2268 1284
rect 2262 1279 2263 1283
rect 2267 1279 2268 1283
rect 2326 1281 2327 1285
rect 2331 1281 2332 1285
rect 2352 1284 2354 1322
rect 2456 1311 2458 1338
rect 2464 1328 2466 1394
rect 2502 1383 2508 1384
rect 2502 1379 2503 1383
rect 2507 1379 2508 1383
rect 2502 1378 2508 1379
rect 2504 1371 2506 1378
rect 2503 1370 2507 1371
rect 2503 1365 2507 1366
rect 2504 1362 2506 1365
rect 2502 1361 2508 1362
rect 2502 1357 2503 1361
rect 2507 1357 2508 1361
rect 2502 1356 2508 1357
rect 2502 1344 2508 1345
rect 2470 1343 2476 1344
rect 2470 1339 2471 1343
rect 2475 1339 2476 1343
rect 2502 1340 2503 1344
rect 2507 1340 2508 1344
rect 2502 1339 2508 1340
rect 2470 1338 2476 1339
rect 2462 1327 2468 1328
rect 2462 1323 2463 1327
rect 2467 1323 2468 1327
rect 2462 1322 2468 1323
rect 2399 1310 2403 1311
rect 2399 1305 2403 1306
rect 2455 1310 2459 1311
rect 2472 1308 2474 1338
rect 2504 1311 2506 1339
rect 2503 1310 2507 1311
rect 2455 1305 2459 1306
rect 2470 1307 2476 1308
rect 2400 1286 2402 1305
rect 2410 1291 2416 1292
rect 2410 1287 2411 1291
rect 2415 1287 2416 1291
rect 2410 1286 2416 1287
rect 2456 1286 2458 1305
rect 2470 1303 2471 1307
rect 2475 1303 2476 1307
rect 2503 1305 2507 1306
rect 2470 1302 2476 1303
rect 2398 1285 2404 1286
rect 2326 1280 2332 1281
rect 2350 1283 2356 1284
rect 2262 1278 2268 1279
rect 2350 1279 2351 1283
rect 2355 1279 2356 1283
rect 2398 1281 2399 1285
rect 2403 1281 2404 1285
rect 2398 1280 2404 1281
rect 2350 1278 2356 1279
rect 1902 1264 1908 1265
rect 1902 1260 1903 1264
rect 1907 1260 1908 1264
rect 1902 1259 1908 1260
rect 1998 1264 2004 1265
rect 1998 1260 1999 1264
rect 2003 1260 2004 1264
rect 1998 1259 2004 1260
rect 2086 1264 2092 1265
rect 2086 1260 2087 1264
rect 2091 1260 2092 1264
rect 2086 1259 2092 1260
rect 2166 1264 2172 1265
rect 2166 1260 2167 1264
rect 2171 1260 2172 1264
rect 2166 1259 2172 1260
rect 2238 1264 2244 1265
rect 2238 1260 2239 1264
rect 2243 1260 2244 1264
rect 2238 1259 2244 1260
rect 1904 1243 1906 1259
rect 2000 1243 2002 1259
rect 2088 1243 2090 1259
rect 2168 1243 2170 1259
rect 2240 1243 2242 1259
rect 1903 1242 1907 1243
rect 1903 1237 1907 1238
rect 1927 1242 1931 1243
rect 1927 1237 1931 1238
rect 1999 1242 2003 1243
rect 1999 1237 2003 1238
rect 2031 1242 2035 1243
rect 2031 1237 2035 1238
rect 2087 1242 2091 1243
rect 2087 1237 2091 1238
rect 2127 1242 2131 1243
rect 2127 1237 2131 1238
rect 2167 1242 2171 1243
rect 2167 1237 2171 1238
rect 2215 1242 2219 1243
rect 2215 1237 2219 1238
rect 2239 1242 2243 1243
rect 2239 1237 2243 1238
rect 1926 1236 1932 1237
rect 1926 1232 1927 1236
rect 1931 1232 1932 1236
rect 1926 1231 1932 1232
rect 2030 1236 2036 1237
rect 2030 1232 2031 1236
rect 2035 1232 2036 1236
rect 2030 1231 2036 1232
rect 2126 1236 2132 1237
rect 2126 1232 2127 1236
rect 2131 1232 2132 1236
rect 2126 1231 2132 1232
rect 2214 1236 2220 1237
rect 2214 1232 2215 1236
rect 2219 1232 2220 1236
rect 2214 1231 2220 1232
rect 1326 1212 1327 1216
rect 1331 1212 1332 1216
rect 1326 1211 1332 1212
rect 1366 1215 1372 1216
rect 1366 1211 1367 1215
rect 1371 1211 1372 1215
rect 1278 1207 1284 1208
rect 1278 1203 1279 1207
rect 1283 1203 1284 1207
rect 1278 1202 1284 1203
rect 1286 1200 1292 1201
rect 590 1199 596 1200
rect 590 1195 591 1199
rect 595 1195 596 1199
rect 590 1194 596 1195
rect 638 1199 644 1200
rect 638 1195 639 1199
rect 643 1195 644 1199
rect 638 1194 644 1195
rect 646 1199 652 1200
rect 646 1195 647 1199
rect 651 1195 652 1199
rect 646 1194 652 1195
rect 654 1199 660 1200
rect 654 1195 655 1199
rect 659 1195 660 1199
rect 654 1194 660 1195
rect 702 1199 708 1200
rect 702 1195 703 1199
rect 707 1195 708 1199
rect 702 1194 708 1195
rect 758 1199 764 1200
rect 758 1195 759 1199
rect 763 1195 764 1199
rect 758 1194 764 1195
rect 774 1199 780 1200
rect 774 1195 775 1199
rect 779 1195 780 1199
rect 774 1194 780 1195
rect 814 1199 820 1200
rect 814 1195 815 1199
rect 819 1195 820 1199
rect 814 1194 820 1195
rect 870 1199 876 1200
rect 870 1195 871 1199
rect 875 1195 876 1199
rect 870 1194 876 1195
rect 886 1199 892 1200
rect 886 1195 887 1199
rect 891 1195 892 1199
rect 886 1194 892 1195
rect 926 1199 932 1200
rect 926 1195 927 1199
rect 931 1195 932 1199
rect 1286 1196 1287 1200
rect 1291 1196 1292 1200
rect 1286 1195 1292 1196
rect 926 1194 932 1195
rect 550 1179 556 1180
rect 550 1175 551 1179
rect 555 1175 556 1179
rect 550 1174 556 1175
rect 592 1171 594 1194
rect 111 1170 115 1171
rect 111 1165 115 1166
rect 367 1170 371 1171
rect 367 1165 371 1166
rect 423 1170 427 1171
rect 423 1165 427 1166
rect 479 1170 483 1171
rect 479 1165 483 1166
rect 535 1170 539 1171
rect 535 1165 539 1166
rect 591 1170 595 1171
rect 591 1165 595 1166
rect 112 1145 114 1165
rect 424 1146 426 1165
rect 480 1146 482 1165
rect 536 1146 538 1165
rect 592 1146 594 1165
rect 640 1160 642 1194
rect 648 1171 650 1194
rect 704 1171 706 1194
rect 760 1171 762 1194
rect 776 1180 778 1194
rect 774 1179 780 1180
rect 774 1175 775 1179
rect 779 1175 780 1179
rect 774 1174 780 1175
rect 816 1171 818 1194
rect 872 1171 874 1194
rect 888 1180 890 1194
rect 894 1183 900 1184
rect 886 1179 892 1180
rect 886 1175 887 1179
rect 891 1175 892 1179
rect 894 1179 895 1183
rect 899 1179 900 1183
rect 894 1178 900 1179
rect 886 1174 892 1175
rect 647 1170 651 1171
rect 647 1165 651 1166
rect 703 1170 707 1171
rect 759 1170 763 1171
rect 703 1165 707 1166
rect 722 1167 728 1168
rect 638 1159 644 1160
rect 638 1155 639 1159
rect 643 1155 644 1159
rect 638 1154 644 1155
rect 648 1146 650 1165
rect 704 1146 706 1165
rect 722 1163 723 1167
rect 727 1163 728 1167
rect 759 1165 763 1166
rect 815 1170 819 1171
rect 815 1165 819 1166
rect 871 1170 875 1171
rect 871 1165 875 1166
rect 722 1162 728 1163
rect 422 1145 428 1146
rect 110 1144 116 1145
rect 110 1140 111 1144
rect 115 1140 116 1144
rect 422 1141 423 1145
rect 427 1141 428 1145
rect 422 1140 428 1141
rect 478 1145 484 1146
rect 478 1141 479 1145
rect 483 1141 484 1145
rect 478 1140 484 1141
rect 534 1145 540 1146
rect 534 1141 535 1145
rect 539 1141 540 1145
rect 590 1145 596 1146
rect 534 1140 540 1141
rect 582 1143 588 1144
rect 110 1139 116 1140
rect 582 1139 583 1143
rect 587 1139 588 1143
rect 590 1141 591 1145
rect 595 1141 596 1145
rect 590 1140 596 1141
rect 646 1145 652 1146
rect 646 1141 647 1145
rect 651 1141 652 1145
rect 646 1140 652 1141
rect 702 1145 708 1146
rect 702 1141 703 1145
rect 707 1141 708 1145
rect 724 1144 726 1162
rect 760 1146 762 1165
rect 816 1146 818 1165
rect 872 1146 874 1165
rect 886 1159 892 1160
rect 886 1155 887 1159
rect 891 1155 892 1159
rect 886 1154 892 1155
rect 758 1145 764 1146
rect 702 1140 708 1141
rect 722 1143 728 1144
rect 582 1138 588 1139
rect 722 1139 723 1143
rect 727 1139 728 1143
rect 758 1141 759 1145
rect 763 1141 764 1145
rect 758 1140 764 1141
rect 814 1145 820 1146
rect 814 1141 815 1145
rect 819 1141 820 1145
rect 814 1140 820 1141
rect 870 1145 876 1146
rect 870 1141 871 1145
rect 875 1141 876 1145
rect 870 1140 876 1141
rect 722 1138 728 1139
rect 110 1127 116 1128
rect 110 1123 111 1127
rect 115 1123 116 1127
rect 110 1122 116 1123
rect 406 1124 412 1125
rect 112 1115 114 1122
rect 406 1120 407 1124
rect 411 1120 412 1124
rect 406 1119 412 1120
rect 462 1124 468 1125
rect 462 1120 463 1124
rect 467 1120 468 1124
rect 462 1119 468 1120
rect 518 1124 524 1125
rect 518 1120 519 1124
rect 523 1120 524 1124
rect 518 1119 524 1120
rect 574 1124 580 1125
rect 574 1120 575 1124
rect 579 1120 580 1124
rect 574 1119 580 1120
rect 408 1115 410 1119
rect 464 1115 466 1119
rect 520 1115 522 1119
rect 576 1115 578 1119
rect 111 1114 115 1115
rect 111 1109 115 1110
rect 223 1114 227 1115
rect 223 1109 227 1110
rect 311 1114 315 1115
rect 311 1109 315 1110
rect 399 1114 403 1115
rect 399 1109 403 1110
rect 407 1114 411 1115
rect 407 1109 411 1110
rect 463 1114 467 1115
rect 463 1109 467 1110
rect 495 1114 499 1115
rect 495 1109 499 1110
rect 519 1114 523 1115
rect 519 1109 523 1110
rect 575 1114 579 1115
rect 575 1109 579 1110
rect 112 1106 114 1109
rect 222 1108 228 1109
rect 110 1105 116 1106
rect 110 1101 111 1105
rect 115 1101 116 1105
rect 222 1104 223 1108
rect 227 1104 228 1108
rect 222 1103 228 1104
rect 310 1108 316 1109
rect 310 1104 311 1108
rect 315 1104 316 1108
rect 310 1103 316 1104
rect 398 1108 404 1109
rect 398 1104 399 1108
rect 403 1104 404 1108
rect 398 1103 404 1104
rect 494 1108 500 1109
rect 494 1104 495 1108
rect 499 1104 500 1108
rect 494 1103 500 1104
rect 110 1100 116 1101
rect 110 1088 116 1089
rect 110 1084 111 1088
rect 115 1084 116 1088
rect 110 1083 116 1084
rect 238 1087 244 1088
rect 238 1083 239 1087
rect 243 1083 244 1087
rect 112 1059 114 1083
rect 238 1082 244 1083
rect 326 1087 332 1088
rect 326 1083 327 1087
rect 331 1083 332 1087
rect 326 1082 332 1083
rect 414 1087 420 1088
rect 414 1083 415 1087
rect 419 1083 420 1087
rect 414 1082 420 1083
rect 422 1087 428 1088
rect 422 1083 423 1087
rect 427 1083 428 1087
rect 422 1082 428 1083
rect 510 1087 516 1088
rect 510 1083 511 1087
rect 515 1083 516 1087
rect 510 1082 516 1083
rect 526 1087 532 1088
rect 526 1083 527 1087
rect 531 1083 532 1087
rect 526 1082 532 1083
rect 240 1059 242 1082
rect 328 1059 330 1082
rect 416 1059 418 1082
rect 111 1058 115 1059
rect 111 1053 115 1054
rect 151 1058 155 1059
rect 151 1053 155 1054
rect 207 1058 211 1059
rect 207 1053 211 1054
rect 239 1058 243 1059
rect 239 1053 243 1054
rect 303 1058 307 1059
rect 303 1053 307 1054
rect 327 1058 331 1059
rect 327 1053 331 1054
rect 415 1058 419 1059
rect 415 1053 419 1054
rect 112 1033 114 1053
rect 152 1034 154 1053
rect 208 1034 210 1053
rect 304 1034 306 1053
rect 416 1034 418 1053
rect 424 1048 426 1082
rect 512 1059 514 1082
rect 528 1068 530 1082
rect 584 1072 586 1138
rect 630 1124 636 1125
rect 630 1120 631 1124
rect 635 1120 636 1124
rect 630 1119 636 1120
rect 686 1124 692 1125
rect 686 1120 687 1124
rect 691 1120 692 1124
rect 686 1119 692 1120
rect 742 1124 748 1125
rect 742 1120 743 1124
rect 747 1120 748 1124
rect 742 1119 748 1120
rect 798 1124 804 1125
rect 798 1120 799 1124
rect 803 1120 804 1124
rect 798 1119 804 1120
rect 854 1124 860 1125
rect 854 1120 855 1124
rect 859 1120 860 1124
rect 854 1119 860 1120
rect 632 1115 634 1119
rect 688 1115 690 1119
rect 744 1115 746 1119
rect 800 1115 802 1119
rect 856 1115 858 1119
rect 591 1114 595 1115
rect 591 1109 595 1110
rect 631 1114 635 1115
rect 631 1109 635 1110
rect 679 1114 683 1115
rect 679 1109 683 1110
rect 687 1114 691 1115
rect 687 1109 691 1110
rect 743 1114 747 1115
rect 743 1109 747 1110
rect 767 1114 771 1115
rect 767 1109 771 1110
rect 799 1114 803 1115
rect 799 1109 803 1110
rect 847 1114 851 1115
rect 847 1109 851 1110
rect 855 1114 859 1115
rect 855 1109 859 1110
rect 590 1108 596 1109
rect 590 1104 591 1108
rect 595 1104 596 1108
rect 590 1103 596 1104
rect 678 1108 684 1109
rect 678 1104 679 1108
rect 683 1104 684 1108
rect 678 1103 684 1104
rect 766 1108 772 1109
rect 766 1104 767 1108
rect 771 1104 772 1108
rect 766 1103 772 1104
rect 846 1108 852 1109
rect 846 1104 847 1108
rect 851 1104 852 1108
rect 846 1103 852 1104
rect 888 1088 890 1154
rect 896 1144 898 1178
rect 928 1171 930 1194
rect 1288 1171 1290 1195
rect 1328 1191 1330 1211
rect 1366 1210 1372 1211
rect 1462 1215 1468 1216
rect 1462 1211 1463 1215
rect 1467 1211 1468 1215
rect 1462 1210 1468 1211
rect 1478 1215 1484 1216
rect 1478 1211 1479 1215
rect 1483 1211 1484 1215
rect 1478 1210 1484 1211
rect 1590 1215 1596 1216
rect 1590 1211 1591 1215
rect 1595 1211 1596 1215
rect 1590 1210 1596 1211
rect 1710 1215 1716 1216
rect 1710 1211 1711 1215
rect 1715 1211 1716 1215
rect 1710 1210 1716 1211
rect 1830 1215 1836 1216
rect 1830 1211 1831 1215
rect 1835 1211 1836 1215
rect 1830 1210 1836 1211
rect 1850 1215 1856 1216
rect 1850 1211 1851 1215
rect 1855 1211 1856 1215
rect 1850 1210 1856 1211
rect 1942 1215 1948 1216
rect 1942 1211 1943 1215
rect 1947 1211 1948 1215
rect 1942 1210 1948 1211
rect 2046 1215 2052 1216
rect 2046 1211 2047 1215
rect 2051 1211 2052 1215
rect 2046 1210 2052 1211
rect 2142 1215 2148 1216
rect 2142 1211 2143 1215
rect 2147 1211 2148 1215
rect 2142 1210 2148 1211
rect 2230 1215 2236 1216
rect 2230 1211 2231 1215
rect 2235 1211 2236 1215
rect 2230 1210 2236 1211
rect 1368 1191 1370 1210
rect 1464 1191 1466 1210
rect 1327 1190 1331 1191
rect 1327 1185 1331 1186
rect 1367 1190 1371 1191
rect 1367 1185 1371 1186
rect 1463 1190 1467 1191
rect 1463 1185 1467 1186
rect 1471 1190 1475 1191
rect 1480 1188 1482 1210
rect 1592 1191 1594 1210
rect 1712 1191 1714 1210
rect 1754 1195 1760 1196
rect 1754 1191 1755 1195
rect 1759 1191 1760 1195
rect 1832 1191 1834 1210
rect 1944 1191 1946 1210
rect 1951 1204 1955 1205
rect 1950 1199 1956 1200
rect 1950 1195 1951 1199
rect 1955 1195 1956 1199
rect 1950 1194 1956 1195
rect 2048 1191 2050 1210
rect 2144 1191 2146 1210
rect 2232 1191 2234 1210
rect 2264 1205 2266 1278
rect 2310 1264 2316 1265
rect 2310 1260 2311 1264
rect 2315 1260 2316 1264
rect 2310 1259 2316 1260
rect 2382 1264 2388 1265
rect 2382 1260 2383 1264
rect 2387 1260 2388 1264
rect 2382 1259 2388 1260
rect 2312 1243 2314 1259
rect 2384 1243 2386 1259
rect 2295 1242 2299 1243
rect 2295 1237 2299 1238
rect 2311 1242 2315 1243
rect 2311 1237 2315 1238
rect 2375 1242 2379 1243
rect 2375 1237 2379 1238
rect 2383 1242 2387 1243
rect 2383 1237 2387 1238
rect 2294 1236 2300 1237
rect 2294 1232 2295 1236
rect 2299 1232 2300 1236
rect 2294 1231 2300 1232
rect 2374 1236 2380 1237
rect 2374 1232 2375 1236
rect 2379 1232 2380 1236
rect 2374 1231 2380 1232
rect 2412 1216 2414 1286
rect 2454 1285 2460 1286
rect 2504 1285 2506 1305
rect 2454 1281 2455 1285
rect 2459 1281 2460 1285
rect 2502 1284 2508 1285
rect 2454 1280 2460 1281
rect 2462 1283 2468 1284
rect 2462 1279 2463 1283
rect 2467 1279 2468 1283
rect 2502 1280 2503 1284
rect 2507 1280 2508 1284
rect 2502 1279 2508 1280
rect 2462 1278 2468 1279
rect 2438 1264 2444 1265
rect 2438 1260 2439 1264
rect 2443 1260 2444 1264
rect 2438 1259 2444 1260
rect 2440 1243 2442 1259
rect 2439 1242 2443 1243
rect 2439 1237 2443 1238
rect 2438 1236 2444 1237
rect 2438 1232 2439 1236
rect 2443 1232 2444 1236
rect 2438 1231 2444 1232
rect 2310 1215 2316 1216
rect 2310 1211 2311 1215
rect 2315 1211 2316 1215
rect 2310 1210 2316 1211
rect 2374 1215 2380 1216
rect 2374 1211 2375 1215
rect 2379 1211 2380 1215
rect 2374 1210 2380 1211
rect 2390 1215 2396 1216
rect 2390 1211 2391 1215
rect 2395 1211 2396 1215
rect 2390 1210 2396 1211
rect 2410 1215 2416 1216
rect 2410 1211 2411 1215
rect 2415 1211 2416 1215
rect 2410 1210 2416 1211
rect 2454 1215 2460 1216
rect 2454 1211 2455 1215
rect 2459 1211 2460 1215
rect 2454 1210 2460 1211
rect 2263 1204 2267 1205
rect 2263 1199 2267 1200
rect 2312 1191 2314 1210
rect 1591 1190 1595 1191
rect 1471 1185 1475 1186
rect 1478 1187 1484 1188
rect 927 1170 931 1171
rect 927 1165 931 1166
rect 983 1170 987 1171
rect 1287 1170 1291 1171
rect 983 1165 987 1166
rect 1002 1167 1008 1168
rect 928 1146 930 1165
rect 984 1146 986 1165
rect 1002 1163 1003 1167
rect 1007 1163 1008 1167
rect 1287 1165 1291 1166
rect 1328 1165 1330 1185
rect 1368 1166 1370 1185
rect 1472 1166 1474 1185
rect 1478 1183 1479 1187
rect 1483 1183 1484 1187
rect 1591 1185 1595 1186
rect 1599 1190 1603 1191
rect 1599 1185 1603 1186
rect 1711 1190 1715 1191
rect 1711 1185 1715 1186
rect 1735 1190 1739 1191
rect 1754 1190 1760 1191
rect 1831 1190 1835 1191
rect 1735 1185 1739 1186
rect 1478 1182 1484 1183
rect 1600 1166 1602 1185
rect 1736 1166 1738 1185
rect 1366 1165 1372 1166
rect 1002 1162 1008 1163
rect 926 1145 932 1146
rect 894 1143 900 1144
rect 894 1139 895 1143
rect 899 1139 900 1143
rect 926 1141 927 1145
rect 931 1141 932 1145
rect 926 1140 932 1141
rect 982 1145 988 1146
rect 982 1141 983 1145
rect 987 1141 988 1145
rect 1004 1144 1006 1162
rect 1288 1145 1290 1165
rect 1326 1164 1332 1165
rect 1326 1160 1327 1164
rect 1331 1160 1332 1164
rect 1366 1161 1367 1165
rect 1371 1161 1372 1165
rect 1366 1160 1372 1161
rect 1470 1165 1476 1166
rect 1470 1161 1471 1165
rect 1475 1161 1476 1165
rect 1470 1160 1476 1161
rect 1598 1165 1604 1166
rect 1598 1161 1599 1165
rect 1603 1161 1604 1165
rect 1734 1165 1740 1166
rect 1598 1160 1604 1161
rect 1606 1163 1612 1164
rect 1326 1159 1332 1160
rect 1606 1159 1607 1163
rect 1611 1159 1612 1163
rect 1734 1161 1735 1165
rect 1739 1161 1740 1165
rect 1756 1164 1758 1190
rect 1831 1185 1835 1186
rect 1863 1190 1867 1191
rect 1863 1185 1867 1186
rect 1943 1190 1947 1191
rect 1943 1185 1947 1186
rect 1983 1190 1987 1191
rect 1983 1185 1987 1186
rect 2047 1190 2051 1191
rect 2047 1185 2051 1186
rect 2087 1190 2091 1191
rect 2087 1185 2091 1186
rect 2143 1190 2147 1191
rect 2143 1185 2147 1186
rect 2191 1190 2195 1191
rect 2231 1190 2235 1191
rect 2191 1185 2195 1186
rect 2210 1187 2216 1188
rect 1854 1179 1860 1180
rect 1854 1175 1855 1179
rect 1859 1175 1860 1179
rect 1854 1174 1860 1175
rect 1734 1160 1740 1161
rect 1754 1163 1760 1164
rect 1606 1158 1612 1159
rect 1754 1159 1755 1163
rect 1759 1159 1760 1163
rect 1754 1158 1760 1159
rect 1326 1147 1332 1148
rect 1286 1144 1292 1145
rect 982 1140 988 1141
rect 1002 1143 1008 1144
rect 894 1138 900 1139
rect 1002 1139 1003 1143
rect 1007 1139 1008 1143
rect 1286 1140 1287 1144
rect 1291 1140 1292 1144
rect 1326 1143 1327 1147
rect 1331 1143 1332 1147
rect 1326 1142 1332 1143
rect 1350 1144 1356 1145
rect 1286 1139 1292 1140
rect 1002 1138 1008 1139
rect 1328 1135 1330 1142
rect 1350 1140 1351 1144
rect 1355 1140 1356 1144
rect 1350 1139 1356 1140
rect 1454 1144 1460 1145
rect 1454 1140 1455 1144
rect 1459 1140 1460 1144
rect 1454 1139 1460 1140
rect 1582 1144 1588 1145
rect 1582 1140 1583 1144
rect 1587 1140 1588 1144
rect 1582 1139 1588 1140
rect 1352 1135 1354 1139
rect 1456 1135 1458 1139
rect 1584 1135 1586 1139
rect 1327 1134 1331 1135
rect 1327 1129 1331 1130
rect 1351 1134 1355 1135
rect 1351 1129 1355 1130
rect 1367 1134 1371 1135
rect 1367 1129 1371 1130
rect 1447 1134 1451 1135
rect 1447 1129 1451 1130
rect 1455 1134 1459 1135
rect 1455 1129 1459 1130
rect 1535 1134 1539 1135
rect 1535 1129 1539 1130
rect 1583 1134 1587 1135
rect 1583 1129 1587 1130
rect 1286 1127 1292 1128
rect 910 1124 916 1125
rect 910 1120 911 1124
rect 915 1120 916 1124
rect 910 1119 916 1120
rect 966 1124 972 1125
rect 966 1120 967 1124
rect 971 1120 972 1124
rect 1286 1123 1287 1127
rect 1291 1123 1292 1127
rect 1328 1126 1330 1129
rect 1366 1128 1372 1129
rect 1286 1122 1292 1123
rect 1326 1125 1332 1126
rect 966 1119 972 1120
rect 912 1115 914 1119
rect 968 1115 970 1119
rect 1288 1115 1290 1122
rect 1326 1121 1327 1125
rect 1331 1121 1332 1125
rect 1366 1124 1367 1128
rect 1371 1124 1372 1128
rect 1366 1123 1372 1124
rect 1446 1128 1452 1129
rect 1446 1124 1447 1128
rect 1451 1124 1452 1128
rect 1446 1123 1452 1124
rect 1534 1128 1540 1129
rect 1534 1124 1535 1128
rect 1539 1124 1540 1128
rect 1534 1123 1540 1124
rect 1326 1120 1332 1121
rect 911 1114 915 1115
rect 911 1109 915 1110
rect 927 1114 931 1115
rect 927 1109 931 1110
rect 967 1114 971 1115
rect 967 1109 971 1110
rect 1015 1114 1019 1115
rect 1015 1109 1019 1110
rect 1103 1114 1107 1115
rect 1103 1109 1107 1110
rect 1287 1114 1291 1115
rect 1287 1109 1291 1110
rect 926 1108 932 1109
rect 926 1104 927 1108
rect 931 1104 932 1108
rect 926 1103 932 1104
rect 1014 1108 1020 1109
rect 1014 1104 1015 1108
rect 1019 1104 1020 1108
rect 1014 1103 1020 1104
rect 1102 1108 1108 1109
rect 1102 1104 1103 1108
rect 1107 1104 1108 1108
rect 1288 1106 1290 1109
rect 1326 1108 1332 1109
rect 1102 1103 1108 1104
rect 1286 1105 1292 1106
rect 1286 1101 1287 1105
rect 1291 1101 1292 1105
rect 1326 1104 1327 1108
rect 1331 1104 1332 1108
rect 1326 1103 1332 1104
rect 1382 1107 1388 1108
rect 1382 1103 1383 1107
rect 1387 1103 1388 1107
rect 1286 1100 1292 1101
rect 1286 1088 1292 1089
rect 606 1087 612 1088
rect 606 1083 607 1087
rect 611 1083 612 1087
rect 606 1082 612 1083
rect 694 1087 700 1088
rect 694 1083 695 1087
rect 699 1083 700 1087
rect 694 1082 700 1083
rect 782 1087 788 1088
rect 782 1083 783 1087
rect 787 1083 788 1087
rect 782 1082 788 1083
rect 862 1087 868 1088
rect 862 1083 863 1087
rect 867 1083 868 1087
rect 862 1082 868 1083
rect 886 1087 892 1088
rect 886 1083 887 1087
rect 891 1083 892 1087
rect 886 1082 892 1083
rect 942 1087 948 1088
rect 942 1083 943 1087
rect 947 1083 948 1087
rect 942 1082 948 1083
rect 1030 1087 1036 1088
rect 1030 1083 1031 1087
rect 1035 1083 1036 1087
rect 1030 1082 1036 1083
rect 1118 1087 1124 1088
rect 1118 1083 1119 1087
rect 1123 1083 1124 1087
rect 1118 1082 1124 1083
rect 1126 1087 1132 1088
rect 1126 1083 1127 1087
rect 1131 1083 1132 1087
rect 1286 1084 1287 1088
rect 1291 1084 1292 1088
rect 1286 1083 1292 1084
rect 1126 1082 1132 1083
rect 582 1071 588 1072
rect 526 1067 532 1068
rect 526 1063 527 1067
rect 531 1063 532 1067
rect 582 1067 583 1071
rect 587 1067 588 1071
rect 582 1066 588 1067
rect 526 1062 532 1063
rect 608 1059 610 1082
rect 696 1059 698 1082
rect 784 1059 786 1082
rect 864 1059 866 1082
rect 944 1059 946 1082
rect 1006 1071 1012 1072
rect 1006 1067 1007 1071
rect 1011 1067 1012 1071
rect 1006 1066 1012 1067
rect 511 1058 515 1059
rect 511 1053 515 1054
rect 535 1058 539 1059
rect 535 1053 539 1054
rect 607 1058 611 1059
rect 607 1053 611 1054
rect 655 1058 659 1059
rect 695 1058 699 1059
rect 655 1053 659 1054
rect 674 1055 680 1056
rect 422 1047 428 1048
rect 422 1043 423 1047
rect 427 1043 428 1047
rect 422 1042 428 1043
rect 536 1034 538 1053
rect 656 1034 658 1053
rect 674 1051 675 1055
rect 679 1051 680 1055
rect 695 1053 699 1054
rect 767 1058 771 1059
rect 767 1053 771 1054
rect 783 1058 787 1059
rect 863 1058 867 1059
rect 783 1053 787 1054
rect 798 1055 804 1056
rect 674 1050 680 1051
rect 150 1033 156 1034
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 150 1029 151 1033
rect 155 1029 156 1033
rect 150 1028 156 1029
rect 206 1033 212 1034
rect 206 1029 207 1033
rect 211 1029 212 1033
rect 206 1028 212 1029
rect 302 1033 308 1034
rect 302 1029 303 1033
rect 307 1029 308 1033
rect 414 1033 420 1034
rect 302 1028 308 1029
rect 334 1031 340 1032
rect 110 1027 116 1028
rect 334 1027 335 1031
rect 339 1027 340 1031
rect 414 1029 415 1033
rect 419 1029 420 1033
rect 414 1028 420 1029
rect 534 1033 540 1034
rect 534 1029 535 1033
rect 539 1029 540 1033
rect 534 1028 540 1029
rect 654 1033 660 1034
rect 654 1029 655 1033
rect 659 1029 660 1033
rect 676 1032 678 1050
rect 768 1034 770 1053
rect 798 1051 799 1055
rect 803 1051 804 1055
rect 863 1053 867 1054
rect 879 1058 883 1059
rect 879 1053 883 1054
rect 943 1058 947 1059
rect 943 1053 947 1054
rect 983 1058 987 1059
rect 983 1053 987 1054
rect 798 1050 804 1051
rect 774 1047 780 1048
rect 774 1043 775 1047
rect 779 1043 780 1047
rect 774 1042 780 1043
rect 776 1037 778 1042
rect 775 1036 779 1037
rect 766 1033 772 1034
rect 654 1028 660 1029
rect 674 1031 680 1032
rect 334 1026 340 1027
rect 674 1027 675 1031
rect 679 1027 680 1031
rect 766 1029 767 1033
rect 771 1029 772 1033
rect 775 1031 779 1032
rect 766 1028 772 1029
rect 674 1026 680 1027
rect 110 1015 116 1016
rect 110 1011 111 1015
rect 115 1011 116 1015
rect 110 1010 116 1011
rect 134 1012 140 1013
rect 112 1003 114 1010
rect 134 1008 135 1012
rect 139 1008 140 1012
rect 134 1007 140 1008
rect 190 1012 196 1013
rect 190 1008 191 1012
rect 195 1008 196 1012
rect 190 1007 196 1008
rect 286 1012 292 1013
rect 286 1008 287 1012
rect 291 1008 292 1012
rect 286 1007 292 1008
rect 136 1003 138 1007
rect 192 1003 194 1007
rect 288 1003 290 1007
rect 111 1002 115 1003
rect 111 997 115 998
rect 135 1002 139 1003
rect 135 997 139 998
rect 191 1002 195 1003
rect 191 997 195 998
rect 215 1002 219 1003
rect 215 997 219 998
rect 287 1002 291 1003
rect 287 997 291 998
rect 327 1002 331 1003
rect 327 997 331 998
rect 112 994 114 997
rect 134 996 140 997
rect 110 993 116 994
rect 110 989 111 993
rect 115 989 116 993
rect 134 992 135 996
rect 139 992 140 996
rect 134 991 140 992
rect 214 996 220 997
rect 214 992 215 996
rect 219 992 220 996
rect 214 991 220 992
rect 326 996 332 997
rect 326 992 327 996
rect 331 992 332 996
rect 326 991 332 992
rect 110 988 116 989
rect 110 976 116 977
rect 110 972 111 976
rect 115 972 116 976
rect 110 971 116 972
rect 150 975 156 976
rect 150 971 151 975
rect 155 971 156 975
rect 112 951 114 971
rect 150 970 156 971
rect 158 975 164 976
rect 158 971 159 975
rect 163 971 164 975
rect 158 970 164 971
rect 230 975 236 976
rect 230 971 231 975
rect 235 971 236 975
rect 230 970 236 971
rect 152 951 154 970
rect 111 950 115 951
rect 111 945 115 946
rect 151 950 155 951
rect 151 945 155 946
rect 112 925 114 945
rect 152 926 154 945
rect 160 940 162 970
rect 232 951 234 970
rect 336 960 338 1026
rect 398 1012 404 1013
rect 398 1008 399 1012
rect 403 1008 404 1012
rect 398 1007 404 1008
rect 518 1012 524 1013
rect 518 1008 519 1012
rect 523 1008 524 1012
rect 518 1007 524 1008
rect 638 1012 644 1013
rect 638 1008 639 1012
rect 643 1008 644 1012
rect 638 1007 644 1008
rect 750 1012 756 1013
rect 750 1008 751 1012
rect 755 1008 756 1012
rect 750 1007 756 1008
rect 400 1003 402 1007
rect 520 1003 522 1007
rect 640 1003 642 1007
rect 752 1003 754 1007
rect 399 1002 403 1003
rect 399 997 403 998
rect 439 1002 443 1003
rect 439 997 443 998
rect 519 1002 523 1003
rect 519 997 523 998
rect 551 1002 555 1003
rect 551 997 555 998
rect 639 1002 643 1003
rect 639 997 643 998
rect 663 1002 667 1003
rect 663 997 667 998
rect 751 1002 755 1003
rect 751 997 755 998
rect 759 1002 763 1003
rect 759 997 763 998
rect 438 996 444 997
rect 438 992 439 996
rect 443 992 444 996
rect 438 991 444 992
rect 550 996 556 997
rect 550 992 551 996
rect 555 992 556 996
rect 550 991 556 992
rect 662 996 668 997
rect 662 992 663 996
rect 667 992 668 996
rect 662 991 668 992
rect 758 996 764 997
rect 758 992 759 996
rect 763 992 764 996
rect 758 991 764 992
rect 800 976 802 1050
rect 880 1034 882 1053
rect 984 1034 986 1053
rect 878 1033 884 1034
rect 878 1029 879 1033
rect 883 1029 884 1033
rect 878 1028 884 1029
rect 982 1033 988 1034
rect 982 1029 983 1033
rect 987 1029 988 1033
rect 1008 1032 1010 1066
rect 1032 1059 1034 1082
rect 1120 1059 1122 1082
rect 1128 1064 1130 1082
rect 1126 1063 1132 1064
rect 1126 1059 1127 1063
rect 1131 1059 1132 1063
rect 1288 1059 1290 1083
rect 1328 1075 1330 1103
rect 1382 1102 1388 1103
rect 1422 1107 1428 1108
rect 1422 1103 1423 1107
rect 1427 1103 1428 1107
rect 1422 1102 1428 1103
rect 1462 1107 1468 1108
rect 1462 1103 1463 1107
rect 1467 1103 1468 1107
rect 1462 1102 1468 1103
rect 1478 1107 1484 1108
rect 1478 1103 1479 1107
rect 1483 1103 1484 1107
rect 1478 1102 1484 1103
rect 1550 1107 1556 1108
rect 1550 1103 1551 1107
rect 1555 1103 1556 1107
rect 1550 1102 1556 1103
rect 1384 1075 1386 1102
rect 1327 1074 1331 1075
rect 1327 1069 1331 1070
rect 1383 1074 1387 1075
rect 1383 1069 1387 1070
rect 1031 1058 1035 1059
rect 1031 1053 1035 1054
rect 1095 1058 1099 1059
rect 1095 1053 1099 1054
rect 1119 1058 1123 1059
rect 1126 1058 1132 1059
rect 1207 1058 1211 1059
rect 1119 1053 1123 1054
rect 1207 1053 1211 1054
rect 1287 1058 1291 1059
rect 1287 1053 1291 1054
rect 1096 1034 1098 1053
rect 1208 1034 1210 1053
rect 1227 1036 1231 1037
rect 1094 1033 1100 1034
rect 982 1028 988 1029
rect 1006 1031 1012 1032
rect 1006 1027 1007 1031
rect 1011 1027 1012 1031
rect 1094 1029 1095 1033
rect 1099 1029 1100 1033
rect 1094 1028 1100 1029
rect 1206 1033 1212 1034
rect 1206 1029 1207 1033
rect 1211 1029 1212 1033
rect 1288 1033 1290 1053
rect 1328 1049 1330 1069
rect 1424 1064 1426 1102
rect 1464 1075 1466 1102
rect 1480 1088 1482 1102
rect 1478 1087 1484 1088
rect 1478 1083 1479 1087
rect 1483 1083 1484 1087
rect 1478 1082 1484 1083
rect 1552 1075 1554 1102
rect 1608 1092 1610 1158
rect 1718 1144 1724 1145
rect 1718 1140 1719 1144
rect 1723 1140 1724 1144
rect 1718 1139 1724 1140
rect 1846 1144 1852 1145
rect 1846 1140 1847 1144
rect 1851 1140 1852 1144
rect 1846 1139 1852 1140
rect 1720 1135 1722 1139
rect 1848 1135 1850 1139
rect 1631 1134 1635 1135
rect 1631 1129 1635 1130
rect 1719 1134 1723 1135
rect 1719 1129 1723 1130
rect 1807 1134 1811 1135
rect 1807 1129 1811 1130
rect 1847 1134 1851 1135
rect 1847 1129 1851 1130
rect 1630 1128 1636 1129
rect 1630 1124 1631 1128
rect 1635 1124 1636 1128
rect 1630 1123 1636 1124
rect 1718 1128 1724 1129
rect 1718 1124 1719 1128
rect 1723 1124 1724 1128
rect 1718 1123 1724 1124
rect 1806 1128 1812 1129
rect 1806 1124 1807 1128
rect 1811 1124 1812 1128
rect 1806 1123 1812 1124
rect 1856 1108 1858 1174
rect 1864 1166 1866 1185
rect 1984 1166 1986 1185
rect 2088 1166 2090 1185
rect 2192 1166 2194 1185
rect 2210 1183 2211 1187
rect 2215 1183 2216 1187
rect 2231 1185 2235 1186
rect 2287 1190 2291 1191
rect 2287 1185 2291 1186
rect 2311 1190 2315 1191
rect 2311 1185 2315 1186
rect 2210 1182 2216 1183
rect 1862 1165 1868 1166
rect 1862 1161 1863 1165
rect 1867 1161 1868 1165
rect 1862 1160 1868 1161
rect 1982 1165 1988 1166
rect 1982 1161 1983 1165
rect 1987 1161 1988 1165
rect 1982 1160 1988 1161
rect 2086 1165 2092 1166
rect 2086 1161 2087 1165
rect 2091 1161 2092 1165
rect 2190 1165 2196 1166
rect 2086 1160 2092 1161
rect 2166 1163 2172 1164
rect 2166 1159 2167 1163
rect 2171 1159 2172 1163
rect 2190 1161 2191 1165
rect 2195 1161 2196 1165
rect 2212 1164 2214 1182
rect 2288 1166 2290 1185
rect 2376 1180 2378 1210
rect 2392 1191 2394 1210
rect 2434 1199 2440 1200
rect 2434 1195 2435 1199
rect 2439 1195 2440 1199
rect 2434 1194 2440 1195
rect 2383 1190 2387 1191
rect 2383 1185 2387 1186
rect 2391 1190 2395 1191
rect 2391 1185 2395 1186
rect 2374 1179 2380 1180
rect 2374 1175 2375 1179
rect 2379 1175 2380 1179
rect 2374 1174 2380 1175
rect 2384 1166 2386 1185
rect 2436 1172 2438 1194
rect 2456 1191 2458 1210
rect 2464 1200 2466 1278
rect 2502 1267 2508 1268
rect 2502 1263 2503 1267
rect 2507 1263 2508 1267
rect 2502 1262 2508 1263
rect 2504 1243 2506 1262
rect 2503 1242 2507 1243
rect 2503 1237 2507 1238
rect 2504 1234 2506 1237
rect 2502 1233 2508 1234
rect 2502 1229 2503 1233
rect 2507 1229 2508 1233
rect 2502 1228 2508 1229
rect 2502 1216 2508 1217
rect 2470 1215 2476 1216
rect 2470 1211 2471 1215
rect 2475 1211 2476 1215
rect 2502 1212 2503 1216
rect 2507 1212 2508 1216
rect 2502 1211 2508 1212
rect 2470 1210 2476 1211
rect 2462 1199 2468 1200
rect 2462 1195 2463 1199
rect 2467 1195 2468 1199
rect 2462 1194 2468 1195
rect 2455 1190 2459 1191
rect 2455 1185 2459 1186
rect 2434 1171 2440 1172
rect 2434 1167 2435 1171
rect 2439 1167 2440 1171
rect 2434 1166 2440 1167
rect 2456 1166 2458 1185
rect 2286 1165 2292 1166
rect 2190 1160 2196 1161
rect 2210 1163 2216 1164
rect 2166 1158 2172 1159
rect 2210 1159 2211 1163
rect 2215 1159 2216 1163
rect 2286 1161 2287 1165
rect 2291 1161 2292 1165
rect 2286 1160 2292 1161
rect 2382 1165 2388 1166
rect 2382 1161 2383 1165
rect 2387 1161 2388 1165
rect 2382 1160 2388 1161
rect 2454 1165 2460 1166
rect 2454 1161 2455 1165
rect 2459 1161 2460 1165
rect 2454 1160 2460 1161
rect 2210 1158 2216 1159
rect 1966 1144 1972 1145
rect 1966 1140 1967 1144
rect 1971 1140 1972 1144
rect 1966 1139 1972 1140
rect 2070 1144 2076 1145
rect 2070 1140 2071 1144
rect 2075 1140 2076 1144
rect 2070 1139 2076 1140
rect 1968 1135 1970 1139
rect 2072 1135 2074 1139
rect 1895 1134 1899 1135
rect 1895 1129 1899 1130
rect 1967 1134 1971 1135
rect 1967 1129 1971 1130
rect 1983 1134 1987 1135
rect 1983 1129 1987 1130
rect 2071 1134 2075 1135
rect 2071 1129 2075 1130
rect 2159 1134 2163 1135
rect 2159 1129 2163 1130
rect 1894 1128 1900 1129
rect 1894 1124 1895 1128
rect 1899 1124 1900 1128
rect 1894 1123 1900 1124
rect 1982 1128 1988 1129
rect 1982 1124 1983 1128
rect 1987 1124 1988 1128
rect 1982 1123 1988 1124
rect 2070 1128 2076 1129
rect 2070 1124 2071 1128
rect 2075 1124 2076 1128
rect 2070 1123 2076 1124
rect 2158 1128 2164 1129
rect 2158 1124 2159 1128
rect 2163 1124 2164 1128
rect 2158 1123 2164 1124
rect 1646 1107 1652 1108
rect 1646 1103 1647 1107
rect 1651 1103 1652 1107
rect 1646 1102 1652 1103
rect 1734 1107 1740 1108
rect 1734 1103 1735 1107
rect 1739 1103 1740 1107
rect 1734 1102 1740 1103
rect 1822 1107 1828 1108
rect 1822 1103 1823 1107
rect 1827 1103 1828 1107
rect 1822 1102 1828 1103
rect 1854 1107 1860 1108
rect 1854 1103 1855 1107
rect 1859 1103 1860 1107
rect 1854 1102 1860 1103
rect 1910 1107 1916 1108
rect 1910 1103 1911 1107
rect 1915 1103 1916 1107
rect 1910 1102 1916 1103
rect 1998 1107 2004 1108
rect 1998 1103 1999 1107
rect 2003 1103 2004 1107
rect 1998 1102 2004 1103
rect 2086 1107 2092 1108
rect 2086 1103 2087 1107
rect 2091 1103 2092 1107
rect 2086 1102 2092 1103
rect 2118 1107 2124 1108
rect 2118 1103 2119 1107
rect 2123 1103 2124 1107
rect 2118 1102 2124 1103
rect 1606 1091 1612 1092
rect 1606 1087 1607 1091
rect 1611 1087 1612 1091
rect 1606 1086 1612 1087
rect 1648 1075 1650 1102
rect 1736 1075 1738 1102
rect 1786 1087 1792 1088
rect 1786 1083 1787 1087
rect 1791 1083 1792 1087
rect 1786 1082 1792 1083
rect 1431 1074 1435 1075
rect 1431 1069 1435 1070
rect 1463 1074 1467 1075
rect 1463 1069 1467 1070
rect 1495 1074 1499 1075
rect 1495 1069 1499 1070
rect 1551 1074 1555 1075
rect 1551 1069 1555 1070
rect 1567 1074 1571 1075
rect 1567 1069 1571 1070
rect 1639 1074 1643 1075
rect 1639 1069 1643 1070
rect 1647 1074 1651 1075
rect 1647 1069 1651 1070
rect 1703 1074 1707 1075
rect 1703 1069 1707 1070
rect 1735 1074 1739 1075
rect 1735 1069 1739 1070
rect 1767 1074 1771 1075
rect 1767 1069 1771 1070
rect 1422 1063 1428 1064
rect 1422 1059 1423 1063
rect 1427 1059 1428 1063
rect 1422 1058 1428 1059
rect 1432 1050 1434 1069
rect 1496 1050 1498 1069
rect 1568 1050 1570 1069
rect 1640 1050 1642 1069
rect 1704 1050 1706 1069
rect 1710 1063 1716 1064
rect 1710 1059 1711 1063
rect 1715 1059 1716 1063
rect 1710 1058 1716 1059
rect 1430 1049 1436 1050
rect 1326 1048 1332 1049
rect 1326 1044 1327 1048
rect 1331 1044 1332 1048
rect 1430 1045 1431 1049
rect 1435 1045 1436 1049
rect 1430 1044 1436 1045
rect 1494 1049 1500 1050
rect 1494 1045 1495 1049
rect 1499 1045 1500 1049
rect 1494 1044 1500 1045
rect 1566 1049 1572 1050
rect 1566 1045 1567 1049
rect 1571 1045 1572 1049
rect 1566 1044 1572 1045
rect 1638 1049 1644 1050
rect 1638 1045 1639 1049
rect 1643 1045 1644 1049
rect 1702 1049 1708 1050
rect 1638 1044 1644 1045
rect 1646 1047 1652 1048
rect 1326 1043 1332 1044
rect 1646 1043 1647 1047
rect 1651 1043 1652 1047
rect 1702 1045 1703 1049
rect 1707 1045 1708 1049
rect 1702 1044 1708 1045
rect 1646 1042 1652 1043
rect 1286 1032 1292 1033
rect 1206 1028 1212 1029
rect 1226 1031 1232 1032
rect 1006 1026 1012 1027
rect 1226 1027 1227 1031
rect 1231 1027 1232 1031
rect 1286 1028 1287 1032
rect 1291 1028 1292 1032
rect 1286 1027 1292 1028
rect 1326 1031 1332 1032
rect 1326 1027 1327 1031
rect 1331 1027 1332 1031
rect 1226 1026 1232 1027
rect 1326 1026 1332 1027
rect 1414 1028 1420 1029
rect 1286 1015 1292 1016
rect 1328 1015 1330 1026
rect 1414 1024 1415 1028
rect 1419 1024 1420 1028
rect 1414 1023 1420 1024
rect 1478 1028 1484 1029
rect 1478 1024 1479 1028
rect 1483 1024 1484 1028
rect 1478 1023 1484 1024
rect 1550 1028 1556 1029
rect 1550 1024 1551 1028
rect 1555 1024 1556 1028
rect 1550 1023 1556 1024
rect 1622 1028 1628 1029
rect 1622 1024 1623 1028
rect 1627 1024 1628 1028
rect 1622 1023 1628 1024
rect 1416 1015 1418 1023
rect 1480 1015 1482 1023
rect 1552 1015 1554 1023
rect 1624 1015 1626 1023
rect 862 1012 868 1013
rect 862 1008 863 1012
rect 867 1008 868 1012
rect 862 1007 868 1008
rect 966 1012 972 1013
rect 966 1008 967 1012
rect 971 1008 972 1012
rect 966 1007 972 1008
rect 1078 1012 1084 1013
rect 1078 1008 1079 1012
rect 1083 1008 1084 1012
rect 1078 1007 1084 1008
rect 1190 1012 1196 1013
rect 1190 1008 1191 1012
rect 1195 1008 1196 1012
rect 1286 1011 1287 1015
rect 1291 1011 1292 1015
rect 1286 1010 1292 1011
rect 1327 1014 1331 1015
rect 1190 1007 1196 1008
rect 864 1003 866 1007
rect 968 1003 970 1007
rect 1080 1003 1082 1007
rect 1192 1003 1194 1007
rect 1288 1003 1290 1010
rect 1327 1009 1331 1010
rect 1415 1014 1419 1015
rect 1415 1009 1419 1010
rect 1479 1014 1483 1015
rect 1479 1009 1483 1010
rect 1511 1014 1515 1015
rect 1511 1009 1515 1010
rect 1551 1014 1555 1015
rect 1551 1009 1555 1010
rect 1567 1014 1571 1015
rect 1567 1009 1571 1010
rect 1623 1014 1627 1015
rect 1623 1009 1627 1010
rect 1328 1006 1330 1009
rect 1510 1008 1516 1009
rect 1326 1005 1332 1006
rect 847 1002 851 1003
rect 847 997 851 998
rect 863 1002 867 1003
rect 863 997 867 998
rect 935 1002 939 1003
rect 935 997 939 998
rect 967 1002 971 1003
rect 967 997 971 998
rect 1015 1002 1019 1003
rect 1015 997 1019 998
rect 1079 1002 1083 1003
rect 1079 997 1083 998
rect 1087 1002 1091 1003
rect 1087 997 1091 998
rect 1167 1002 1171 1003
rect 1167 997 1171 998
rect 1191 1002 1195 1003
rect 1191 997 1195 998
rect 1223 1002 1227 1003
rect 1223 997 1227 998
rect 1287 1002 1291 1003
rect 1326 1001 1327 1005
rect 1331 1001 1332 1005
rect 1510 1004 1511 1008
rect 1515 1004 1516 1008
rect 1510 1003 1516 1004
rect 1566 1008 1572 1009
rect 1566 1004 1567 1008
rect 1571 1004 1572 1008
rect 1566 1003 1572 1004
rect 1622 1008 1628 1009
rect 1622 1004 1623 1008
rect 1627 1004 1628 1008
rect 1622 1003 1628 1004
rect 1326 1000 1332 1001
rect 1287 997 1291 998
rect 846 996 852 997
rect 846 992 847 996
rect 851 992 852 996
rect 846 991 852 992
rect 934 996 940 997
rect 934 992 935 996
rect 939 992 940 996
rect 934 991 940 992
rect 1014 996 1020 997
rect 1014 992 1015 996
rect 1019 992 1020 996
rect 1014 991 1020 992
rect 1086 996 1092 997
rect 1086 992 1087 996
rect 1091 992 1092 996
rect 1086 991 1092 992
rect 1166 996 1172 997
rect 1166 992 1167 996
rect 1171 992 1172 996
rect 1166 991 1172 992
rect 1222 996 1228 997
rect 1222 992 1223 996
rect 1227 992 1228 996
rect 1288 994 1290 997
rect 1222 991 1228 992
rect 1286 993 1292 994
rect 1286 989 1287 993
rect 1291 989 1292 993
rect 1286 988 1292 989
rect 1326 988 1332 989
rect 1326 984 1327 988
rect 1331 984 1332 988
rect 1326 983 1332 984
rect 1526 987 1532 988
rect 1526 983 1527 987
rect 1531 983 1532 987
rect 1286 976 1292 977
rect 342 975 348 976
rect 342 971 343 975
rect 347 971 348 975
rect 342 970 348 971
rect 454 975 460 976
rect 454 971 455 975
rect 459 971 460 975
rect 454 970 460 971
rect 566 975 572 976
rect 566 971 567 975
rect 571 971 572 975
rect 566 970 572 971
rect 574 975 580 976
rect 574 971 575 975
rect 579 971 580 975
rect 574 970 580 971
rect 678 975 684 976
rect 678 971 679 975
rect 683 971 684 975
rect 678 970 684 971
rect 774 975 780 976
rect 774 971 775 975
rect 779 971 780 975
rect 774 970 780 971
rect 798 975 804 976
rect 798 971 799 975
rect 803 971 804 975
rect 798 970 804 971
rect 862 975 868 976
rect 862 971 863 975
rect 867 971 868 975
rect 862 970 868 971
rect 918 975 924 976
rect 918 971 919 975
rect 923 971 924 975
rect 918 970 924 971
rect 950 975 956 976
rect 950 971 951 975
rect 955 971 956 975
rect 950 970 956 971
rect 1030 975 1036 976
rect 1030 971 1031 975
rect 1035 971 1036 975
rect 1030 970 1036 971
rect 1046 975 1052 976
rect 1046 971 1047 975
rect 1051 971 1052 975
rect 1046 970 1052 971
rect 1102 975 1108 976
rect 1102 971 1103 975
rect 1107 971 1108 975
rect 1102 970 1108 971
rect 1182 975 1188 976
rect 1182 971 1183 975
rect 1187 971 1188 975
rect 1182 970 1188 971
rect 1238 975 1244 976
rect 1238 971 1239 975
rect 1243 971 1244 975
rect 1238 970 1244 971
rect 1246 975 1252 976
rect 1246 971 1247 975
rect 1251 971 1252 975
rect 1286 972 1287 976
rect 1291 972 1292 976
rect 1286 971 1292 972
rect 1246 970 1252 971
rect 334 959 340 960
rect 334 955 335 959
rect 339 955 340 959
rect 334 954 340 955
rect 344 951 346 970
rect 456 951 458 970
rect 568 951 570 970
rect 576 952 578 970
rect 574 951 580 952
rect 680 951 682 970
rect 776 951 778 970
rect 854 959 860 960
rect 854 955 855 959
rect 859 955 860 959
rect 854 954 860 955
rect 207 950 211 951
rect 207 945 211 946
rect 231 950 235 951
rect 231 945 235 946
rect 295 950 299 951
rect 295 945 299 946
rect 343 950 347 951
rect 343 945 347 946
rect 399 950 403 951
rect 399 945 403 946
rect 455 950 459 951
rect 455 945 459 946
rect 511 950 515 951
rect 511 945 515 946
rect 567 950 571 951
rect 574 947 575 951
rect 579 947 580 951
rect 574 946 580 947
rect 623 950 627 951
rect 567 945 571 946
rect 623 945 627 946
rect 679 950 683 951
rect 679 945 683 946
rect 735 950 739 951
rect 775 950 779 951
rect 735 945 739 946
rect 766 947 772 948
rect 158 939 164 940
rect 158 935 159 939
rect 163 935 164 939
rect 158 934 164 935
rect 208 926 210 945
rect 296 926 298 945
rect 400 926 402 945
rect 430 931 436 932
rect 430 927 431 931
rect 435 927 436 931
rect 430 926 436 927
rect 512 926 514 945
rect 534 939 540 940
rect 534 935 535 939
rect 539 935 540 939
rect 534 934 540 935
rect 150 925 156 926
rect 110 924 116 925
rect 110 920 111 924
rect 115 920 116 924
rect 150 921 151 925
rect 155 921 156 925
rect 150 920 156 921
rect 206 925 212 926
rect 206 921 207 925
rect 211 921 212 925
rect 206 920 212 921
rect 294 925 300 926
rect 294 921 295 925
rect 299 921 300 925
rect 294 920 300 921
rect 398 925 404 926
rect 398 921 399 925
rect 403 921 404 925
rect 398 920 404 921
rect 110 919 116 920
rect 110 907 116 908
rect 110 903 111 907
rect 115 903 116 907
rect 110 902 116 903
rect 134 904 140 905
rect 112 895 114 902
rect 134 900 135 904
rect 139 900 140 904
rect 134 899 140 900
rect 190 904 196 905
rect 190 900 191 904
rect 195 900 196 904
rect 190 899 196 900
rect 278 904 284 905
rect 278 900 279 904
rect 283 900 284 904
rect 278 899 284 900
rect 382 904 388 905
rect 382 900 383 904
rect 387 900 388 904
rect 382 899 388 900
rect 136 895 138 899
rect 192 895 194 899
rect 280 895 282 899
rect 384 895 386 899
rect 111 894 115 895
rect 111 889 115 890
rect 135 894 139 895
rect 135 889 139 890
rect 191 894 195 895
rect 191 889 195 890
rect 247 894 251 895
rect 247 889 251 890
rect 279 894 283 895
rect 279 889 283 890
rect 343 894 347 895
rect 343 889 347 890
rect 383 894 387 895
rect 383 889 387 890
rect 112 886 114 889
rect 246 888 252 889
rect 110 885 116 886
rect 110 881 111 885
rect 115 881 116 885
rect 246 884 247 888
rect 251 884 252 888
rect 246 883 252 884
rect 342 888 348 889
rect 342 884 343 888
rect 347 884 348 888
rect 342 883 348 884
rect 110 880 116 881
rect 110 868 116 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 262 867 268 868
rect 262 863 263 867
rect 267 863 268 867
rect 112 839 114 863
rect 262 862 268 863
rect 358 867 364 868
rect 358 863 359 867
rect 363 863 364 867
rect 358 862 364 863
rect 264 839 266 862
rect 360 839 362 862
rect 432 848 434 926
rect 510 925 516 926
rect 510 921 511 925
rect 515 921 516 925
rect 536 924 538 934
rect 624 926 626 945
rect 736 926 738 945
rect 766 943 767 947
rect 771 943 772 947
rect 775 945 779 946
rect 831 950 835 951
rect 831 945 835 946
rect 766 942 772 943
rect 622 925 628 926
rect 510 920 516 921
rect 534 923 540 924
rect 534 919 535 923
rect 539 919 540 923
rect 622 921 623 925
rect 627 921 628 925
rect 622 920 628 921
rect 734 925 740 926
rect 734 921 735 925
rect 739 921 740 925
rect 734 920 740 921
rect 534 918 540 919
rect 494 904 500 905
rect 494 900 495 904
rect 499 900 500 904
rect 494 899 500 900
rect 606 904 612 905
rect 606 900 607 904
rect 611 900 612 904
rect 606 899 612 900
rect 718 904 724 905
rect 718 900 719 904
rect 723 900 724 904
rect 718 899 724 900
rect 496 895 498 899
rect 608 895 610 899
rect 720 895 722 899
rect 439 894 443 895
rect 439 889 443 890
rect 495 894 499 895
rect 495 889 499 890
rect 543 894 547 895
rect 543 889 547 890
rect 607 894 611 895
rect 607 889 611 890
rect 647 894 651 895
rect 647 889 651 890
rect 719 894 723 895
rect 719 889 723 890
rect 743 894 747 895
rect 743 889 747 890
rect 438 888 444 889
rect 438 884 439 888
rect 443 884 444 888
rect 438 883 444 884
rect 542 888 548 889
rect 542 884 543 888
rect 547 884 548 888
rect 542 883 548 884
rect 646 888 652 889
rect 646 884 647 888
rect 651 884 652 888
rect 646 883 652 884
rect 742 888 748 889
rect 742 884 743 888
rect 747 884 748 888
rect 742 883 748 884
rect 768 868 770 942
rect 832 926 834 945
rect 830 925 836 926
rect 830 921 831 925
rect 835 921 836 925
rect 856 924 858 954
rect 864 951 866 970
rect 863 950 867 951
rect 863 945 867 946
rect 920 940 922 970
rect 952 951 954 970
rect 1032 951 1034 970
rect 1048 956 1050 970
rect 1046 955 1052 956
rect 1046 951 1047 955
rect 1051 951 1052 955
rect 1104 951 1106 970
rect 1184 951 1186 970
rect 1190 959 1196 960
rect 1190 955 1191 959
rect 1195 955 1196 959
rect 1190 954 1196 955
rect 927 950 931 951
rect 927 945 931 946
rect 951 950 955 951
rect 951 945 955 946
rect 1015 950 1019 951
rect 1015 945 1019 946
rect 1031 950 1035 951
rect 1046 950 1052 951
rect 1095 950 1099 951
rect 1031 945 1035 946
rect 1095 945 1099 946
rect 1103 950 1107 951
rect 1103 945 1107 946
rect 1175 950 1179 951
rect 1175 945 1179 946
rect 1183 950 1187 951
rect 1183 945 1187 946
rect 918 939 924 940
rect 918 935 919 939
rect 923 935 924 939
rect 918 934 924 935
rect 928 926 930 945
rect 1016 926 1018 945
rect 1096 926 1098 945
rect 1176 926 1178 945
rect 926 925 932 926
rect 830 920 836 921
rect 854 923 860 924
rect 854 919 855 923
rect 859 919 860 923
rect 926 921 927 925
rect 931 921 932 925
rect 926 920 932 921
rect 1014 925 1020 926
rect 1014 921 1015 925
rect 1019 921 1020 925
rect 1014 920 1020 921
rect 1094 925 1100 926
rect 1094 921 1095 925
rect 1099 921 1100 925
rect 1174 925 1180 926
rect 1094 920 1100 921
rect 1118 923 1124 924
rect 854 918 860 919
rect 1118 919 1119 923
rect 1123 919 1124 923
rect 1174 921 1175 925
rect 1179 921 1180 925
rect 1192 924 1194 954
rect 1240 951 1242 970
rect 1248 952 1250 970
rect 1246 951 1252 952
rect 1288 951 1290 971
rect 1239 950 1243 951
rect 1246 947 1247 951
rect 1251 947 1252 951
rect 1246 946 1252 947
rect 1287 950 1291 951
rect 1328 947 1330 983
rect 1526 982 1532 983
rect 1534 987 1540 988
rect 1534 983 1535 987
rect 1539 983 1540 987
rect 1534 982 1540 983
rect 1582 987 1588 988
rect 1582 983 1583 987
rect 1587 983 1588 987
rect 1582 982 1588 983
rect 1598 987 1604 988
rect 1598 983 1599 987
rect 1603 983 1604 987
rect 1598 982 1604 983
rect 1638 987 1644 988
rect 1638 983 1639 987
rect 1643 983 1644 987
rect 1638 982 1644 983
rect 1528 947 1530 982
rect 1239 945 1243 946
rect 1287 945 1291 946
rect 1327 946 1331 947
rect 1240 926 1242 945
rect 1246 939 1252 940
rect 1246 935 1247 939
rect 1251 935 1252 939
rect 1246 934 1252 935
rect 1262 939 1268 940
rect 1262 935 1263 939
rect 1267 935 1268 939
rect 1262 934 1268 935
rect 1238 925 1244 926
rect 1174 920 1180 921
rect 1190 923 1196 924
rect 1118 918 1124 919
rect 1190 919 1191 923
rect 1195 919 1196 923
rect 1238 921 1239 925
rect 1243 921 1244 925
rect 1238 920 1244 921
rect 1190 918 1196 919
rect 814 904 820 905
rect 814 900 815 904
rect 819 900 820 904
rect 814 899 820 900
rect 910 904 916 905
rect 910 900 911 904
rect 915 900 916 904
rect 910 899 916 900
rect 998 904 1004 905
rect 998 900 999 904
rect 1003 900 1004 904
rect 998 899 1004 900
rect 1078 904 1084 905
rect 1078 900 1079 904
rect 1083 900 1084 904
rect 1078 899 1084 900
rect 816 895 818 899
rect 912 895 914 899
rect 1000 895 1002 899
rect 1080 895 1082 899
rect 815 894 819 895
rect 815 889 819 890
rect 839 894 843 895
rect 839 889 843 890
rect 911 894 915 895
rect 911 889 915 890
rect 927 894 931 895
rect 927 889 931 890
rect 999 894 1003 895
rect 999 889 1003 890
rect 1007 894 1011 895
rect 1007 889 1011 890
rect 1079 894 1083 895
rect 1079 889 1083 890
rect 1087 894 1091 895
rect 1087 889 1091 890
rect 838 888 844 889
rect 838 884 839 888
rect 843 884 844 888
rect 838 883 844 884
rect 926 888 932 889
rect 926 884 927 888
rect 931 884 932 888
rect 926 883 932 884
rect 1006 888 1012 889
rect 1006 884 1007 888
rect 1011 884 1012 888
rect 1006 883 1012 884
rect 1086 888 1092 889
rect 1086 884 1087 888
rect 1091 884 1092 888
rect 1086 883 1092 884
rect 454 867 460 868
rect 454 863 455 867
rect 459 863 460 867
rect 454 862 460 863
rect 558 867 564 868
rect 558 863 559 867
rect 563 863 564 867
rect 558 862 564 863
rect 662 867 668 868
rect 662 863 663 867
rect 667 863 668 867
rect 662 862 668 863
rect 670 867 676 868
rect 670 863 671 867
rect 675 863 676 867
rect 670 862 676 863
rect 758 867 764 868
rect 758 863 759 867
rect 763 863 764 867
rect 758 862 764 863
rect 766 867 772 868
rect 766 863 767 867
rect 771 863 772 867
rect 766 862 772 863
rect 854 867 860 868
rect 854 863 855 867
rect 859 863 860 867
rect 854 862 860 863
rect 942 867 948 868
rect 942 863 943 867
rect 947 863 948 867
rect 942 862 948 863
rect 1022 867 1028 868
rect 1022 863 1023 867
rect 1027 863 1028 867
rect 1022 862 1028 863
rect 1102 867 1108 868
rect 1102 863 1103 867
rect 1107 863 1108 867
rect 1102 862 1108 863
rect 430 847 436 848
rect 430 843 431 847
rect 435 843 436 847
rect 430 842 436 843
rect 456 839 458 862
rect 560 839 562 862
rect 664 839 666 862
rect 111 838 115 839
rect 111 833 115 834
rect 239 838 243 839
rect 239 833 243 834
rect 263 838 267 839
rect 263 833 267 834
rect 303 838 307 839
rect 303 833 307 834
rect 359 838 363 839
rect 359 833 363 834
rect 383 838 387 839
rect 455 838 459 839
rect 383 833 387 834
rect 402 835 408 836
rect 112 813 114 833
rect 240 814 242 833
rect 304 814 306 833
rect 384 814 386 833
rect 402 831 403 835
rect 407 831 408 835
rect 455 833 459 834
rect 463 838 467 839
rect 463 833 467 834
rect 551 838 555 839
rect 551 833 555 834
rect 559 838 563 839
rect 559 833 563 834
rect 639 838 643 839
rect 639 833 643 834
rect 663 838 667 839
rect 663 833 667 834
rect 402 830 408 831
rect 238 813 244 814
rect 110 812 116 813
rect 110 808 111 812
rect 115 808 116 812
rect 238 809 239 813
rect 243 809 244 813
rect 238 808 244 809
rect 302 813 308 814
rect 302 809 303 813
rect 307 809 308 813
rect 382 813 388 814
rect 302 808 308 809
rect 350 811 356 812
rect 110 807 116 808
rect 350 807 351 811
rect 355 807 356 811
rect 382 809 383 813
rect 387 809 388 813
rect 404 812 406 830
rect 464 814 466 833
rect 552 814 554 833
rect 640 814 642 833
rect 672 828 674 862
rect 760 839 762 862
rect 856 839 858 862
rect 944 839 946 862
rect 1024 839 1026 862
rect 1090 839 1096 840
rect 1104 839 1106 862
rect 1120 848 1122 918
rect 1158 904 1164 905
rect 1158 900 1159 904
rect 1163 900 1164 904
rect 1158 899 1164 900
rect 1222 904 1228 905
rect 1222 900 1223 904
rect 1227 900 1228 904
rect 1222 899 1228 900
rect 1160 895 1162 899
rect 1224 895 1226 899
rect 1159 894 1163 895
rect 1159 889 1163 890
rect 1167 894 1171 895
rect 1167 889 1171 890
rect 1223 894 1227 895
rect 1223 889 1227 890
rect 1166 888 1172 889
rect 1166 884 1167 888
rect 1171 884 1172 888
rect 1166 883 1172 884
rect 1222 888 1228 889
rect 1222 884 1223 888
rect 1227 884 1228 888
rect 1222 883 1228 884
rect 1248 868 1250 934
rect 1264 924 1266 934
rect 1288 925 1290 945
rect 1327 941 1331 942
rect 1367 946 1371 947
rect 1367 941 1371 942
rect 1439 946 1443 947
rect 1439 941 1443 942
rect 1527 946 1531 947
rect 1536 944 1538 982
rect 1584 947 1586 982
rect 1600 968 1602 982
rect 1598 967 1604 968
rect 1598 963 1599 967
rect 1603 963 1604 967
rect 1598 962 1604 963
rect 1640 947 1642 982
rect 1648 972 1650 1042
rect 1686 1028 1692 1029
rect 1686 1024 1687 1028
rect 1691 1024 1692 1028
rect 1686 1023 1692 1024
rect 1688 1015 1690 1023
rect 1679 1014 1683 1015
rect 1679 1009 1683 1010
rect 1687 1014 1691 1015
rect 1687 1009 1691 1010
rect 1678 1008 1684 1009
rect 1678 1004 1679 1008
rect 1683 1004 1684 1008
rect 1678 1003 1684 1004
rect 1712 988 1714 1058
rect 1768 1050 1770 1069
rect 1766 1049 1772 1050
rect 1766 1045 1767 1049
rect 1771 1045 1772 1049
rect 1788 1048 1790 1082
rect 1824 1075 1826 1102
rect 1912 1075 1914 1102
rect 1959 1092 1963 1093
rect 1958 1087 1959 1092
rect 1963 1087 1964 1092
rect 1958 1086 1964 1087
rect 2000 1075 2002 1102
rect 2088 1075 2090 1102
rect 1823 1074 1827 1075
rect 1823 1069 1827 1070
rect 1839 1074 1843 1075
rect 1839 1069 1843 1070
rect 1911 1074 1915 1075
rect 1911 1069 1915 1070
rect 1919 1074 1923 1075
rect 1919 1069 1923 1070
rect 1999 1074 2003 1075
rect 1999 1069 2003 1070
rect 2007 1074 2011 1075
rect 2007 1069 2011 1070
rect 2087 1074 2091 1075
rect 2087 1069 2091 1070
rect 2111 1074 2115 1075
rect 2111 1069 2115 1070
rect 1840 1050 1842 1069
rect 1920 1050 1922 1069
rect 2008 1050 2010 1069
rect 2112 1050 2114 1069
rect 2120 1064 2122 1102
rect 2168 1092 2170 1158
rect 2174 1144 2180 1145
rect 2174 1140 2175 1144
rect 2179 1140 2180 1144
rect 2174 1139 2180 1140
rect 2270 1144 2276 1145
rect 2270 1140 2271 1144
rect 2275 1140 2276 1144
rect 2270 1139 2276 1140
rect 2366 1144 2372 1145
rect 2366 1140 2367 1144
rect 2371 1140 2372 1144
rect 2366 1139 2372 1140
rect 2438 1144 2444 1145
rect 2438 1140 2439 1144
rect 2443 1140 2444 1144
rect 2438 1139 2444 1140
rect 2176 1135 2178 1139
rect 2272 1135 2274 1139
rect 2368 1135 2370 1139
rect 2440 1135 2442 1139
rect 2175 1134 2179 1135
rect 2175 1129 2179 1130
rect 2255 1134 2259 1135
rect 2255 1129 2259 1130
rect 2271 1134 2275 1135
rect 2271 1129 2275 1130
rect 2359 1134 2363 1135
rect 2359 1129 2363 1130
rect 2367 1134 2371 1135
rect 2367 1129 2371 1130
rect 2439 1134 2443 1135
rect 2439 1129 2443 1130
rect 2254 1128 2260 1129
rect 2254 1124 2255 1128
rect 2259 1124 2260 1128
rect 2254 1123 2260 1124
rect 2358 1128 2364 1129
rect 2358 1124 2359 1128
rect 2363 1124 2364 1128
rect 2358 1123 2364 1124
rect 2438 1128 2444 1129
rect 2438 1124 2439 1128
rect 2443 1124 2444 1128
rect 2438 1123 2444 1124
rect 2174 1107 2180 1108
rect 2174 1103 2175 1107
rect 2179 1103 2180 1107
rect 2174 1102 2180 1103
rect 2270 1107 2276 1108
rect 2270 1103 2271 1107
rect 2275 1103 2276 1107
rect 2270 1102 2276 1103
rect 2374 1107 2380 1108
rect 2374 1103 2375 1107
rect 2379 1103 2380 1107
rect 2374 1102 2380 1103
rect 2382 1107 2388 1108
rect 2382 1103 2383 1107
rect 2387 1103 2388 1107
rect 2382 1102 2388 1103
rect 2454 1107 2460 1108
rect 2454 1103 2455 1107
rect 2459 1103 2460 1107
rect 2454 1102 2460 1103
rect 2462 1107 2468 1108
rect 2462 1103 2463 1107
rect 2467 1103 2468 1107
rect 2462 1102 2468 1103
rect 2166 1091 2172 1092
rect 2166 1087 2167 1091
rect 2171 1087 2172 1091
rect 2166 1086 2172 1087
rect 2176 1075 2178 1102
rect 2272 1075 2274 1102
rect 2376 1075 2378 1102
rect 2384 1093 2386 1102
rect 2383 1092 2387 1093
rect 2383 1087 2387 1088
rect 2456 1075 2458 1102
rect 2175 1074 2179 1075
rect 2175 1069 2179 1070
rect 2231 1074 2235 1075
rect 2231 1069 2235 1070
rect 2271 1074 2275 1075
rect 2271 1069 2275 1070
rect 2351 1074 2355 1075
rect 2375 1074 2379 1075
rect 2351 1069 2355 1070
rect 2366 1071 2372 1072
rect 2118 1063 2124 1064
rect 2118 1059 2119 1063
rect 2123 1059 2124 1063
rect 2118 1058 2124 1059
rect 2232 1050 2234 1069
rect 2352 1050 2354 1069
rect 2366 1067 2367 1071
rect 2371 1067 2372 1071
rect 2375 1069 2379 1070
rect 2455 1074 2459 1075
rect 2455 1069 2459 1070
rect 2366 1066 2372 1067
rect 1838 1049 1844 1050
rect 1766 1044 1772 1045
rect 1786 1047 1792 1048
rect 1786 1043 1787 1047
rect 1791 1043 1792 1047
rect 1838 1045 1839 1049
rect 1843 1045 1844 1049
rect 1838 1044 1844 1045
rect 1918 1049 1924 1050
rect 1918 1045 1919 1049
rect 1923 1045 1924 1049
rect 1918 1044 1924 1045
rect 2006 1049 2012 1050
rect 2006 1045 2007 1049
rect 2011 1045 2012 1049
rect 2110 1049 2116 1050
rect 2006 1044 2012 1045
rect 2014 1047 2020 1048
rect 1786 1042 1792 1043
rect 2014 1043 2015 1047
rect 2019 1043 2020 1047
rect 2110 1045 2111 1049
rect 2115 1045 2116 1049
rect 2110 1044 2116 1045
rect 2230 1049 2236 1050
rect 2230 1045 2231 1049
rect 2235 1045 2236 1049
rect 2230 1044 2236 1045
rect 2350 1049 2356 1050
rect 2350 1045 2351 1049
rect 2355 1045 2356 1049
rect 2368 1048 2370 1066
rect 2456 1050 2458 1069
rect 2464 1064 2466 1102
rect 2472 1092 2474 1210
rect 2504 1191 2506 1211
rect 2503 1190 2507 1191
rect 2503 1185 2507 1186
rect 2478 1179 2484 1180
rect 2478 1175 2479 1179
rect 2483 1175 2484 1179
rect 2478 1174 2484 1175
rect 2470 1091 2476 1092
rect 2470 1087 2471 1091
rect 2475 1087 2476 1091
rect 2470 1086 2476 1087
rect 2462 1063 2468 1064
rect 2462 1059 2463 1063
rect 2467 1059 2468 1063
rect 2462 1058 2468 1059
rect 2454 1049 2460 1050
rect 2350 1044 2356 1045
rect 2366 1047 2372 1048
rect 2014 1042 2020 1043
rect 2366 1043 2367 1047
rect 2371 1043 2372 1047
rect 2454 1045 2455 1049
rect 2459 1045 2460 1049
rect 2454 1044 2460 1045
rect 2462 1047 2468 1048
rect 2366 1042 2372 1043
rect 2462 1043 2463 1047
rect 2467 1043 2468 1047
rect 2462 1042 2468 1043
rect 1750 1028 1756 1029
rect 1750 1024 1751 1028
rect 1755 1024 1756 1028
rect 1750 1023 1756 1024
rect 1822 1028 1828 1029
rect 1822 1024 1823 1028
rect 1827 1024 1828 1028
rect 1822 1023 1828 1024
rect 1902 1028 1908 1029
rect 1902 1024 1903 1028
rect 1907 1024 1908 1028
rect 1902 1023 1908 1024
rect 1990 1028 1996 1029
rect 1990 1024 1991 1028
rect 1995 1024 1996 1028
rect 1990 1023 1996 1024
rect 1752 1015 1754 1023
rect 1824 1015 1826 1023
rect 1904 1015 1906 1023
rect 1992 1015 1994 1023
rect 1735 1014 1739 1015
rect 1735 1009 1739 1010
rect 1751 1014 1755 1015
rect 1751 1009 1755 1010
rect 1807 1014 1811 1015
rect 1807 1009 1811 1010
rect 1823 1014 1827 1015
rect 1823 1009 1827 1010
rect 1887 1014 1891 1015
rect 1887 1009 1891 1010
rect 1903 1014 1907 1015
rect 1903 1009 1907 1010
rect 1983 1014 1987 1015
rect 1983 1009 1987 1010
rect 1991 1014 1995 1015
rect 1991 1009 1995 1010
rect 1734 1008 1740 1009
rect 1734 1004 1735 1008
rect 1739 1004 1740 1008
rect 1734 1003 1740 1004
rect 1806 1008 1812 1009
rect 1806 1004 1807 1008
rect 1811 1004 1812 1008
rect 1806 1003 1812 1004
rect 1886 1008 1892 1009
rect 1886 1004 1887 1008
rect 1891 1004 1892 1008
rect 1886 1003 1892 1004
rect 1982 1008 1988 1009
rect 1982 1004 1983 1008
rect 1987 1004 1988 1008
rect 1982 1003 1988 1004
rect 1694 987 1700 988
rect 1694 983 1695 987
rect 1699 983 1700 987
rect 1694 982 1700 983
rect 1710 987 1716 988
rect 1710 983 1711 987
rect 1715 983 1716 987
rect 1710 982 1716 983
rect 1750 987 1756 988
rect 1750 983 1751 987
rect 1755 983 1756 987
rect 1750 982 1756 983
rect 1782 987 1788 988
rect 1782 983 1783 987
rect 1787 983 1788 987
rect 1782 982 1788 983
rect 1822 987 1828 988
rect 1822 983 1823 987
rect 1827 983 1828 987
rect 1822 982 1828 983
rect 1902 987 1908 988
rect 1902 983 1903 987
rect 1907 983 1908 987
rect 1902 982 1908 983
rect 1998 987 2004 988
rect 2016 987 2018 1042
rect 2094 1028 2100 1029
rect 2094 1024 2095 1028
rect 2099 1024 2100 1028
rect 2094 1023 2100 1024
rect 2214 1028 2220 1029
rect 2214 1024 2215 1028
rect 2219 1024 2220 1028
rect 2214 1023 2220 1024
rect 2334 1028 2340 1029
rect 2334 1024 2335 1028
rect 2339 1024 2340 1028
rect 2334 1023 2340 1024
rect 2438 1028 2444 1029
rect 2438 1024 2439 1028
rect 2443 1024 2444 1028
rect 2438 1023 2444 1024
rect 2096 1015 2098 1023
rect 2216 1015 2218 1023
rect 2336 1015 2338 1023
rect 2440 1015 2442 1023
rect 2095 1014 2099 1015
rect 2095 1009 2099 1010
rect 2215 1014 2219 1015
rect 2215 1009 2219 1010
rect 2335 1014 2339 1015
rect 2335 1009 2339 1010
rect 2439 1014 2443 1015
rect 2439 1009 2443 1010
rect 2094 1008 2100 1009
rect 2094 1004 2095 1008
rect 2099 1004 2100 1008
rect 2094 1003 2100 1004
rect 2214 1008 2220 1009
rect 2214 1004 2215 1008
rect 2219 1004 2220 1008
rect 2214 1003 2220 1004
rect 2334 1008 2340 1009
rect 2334 1004 2335 1008
rect 2339 1004 2340 1008
rect 2334 1003 2340 1004
rect 2438 1008 2444 1009
rect 2438 1004 2439 1008
rect 2443 1004 2444 1008
rect 2438 1003 2444 1004
rect 1998 983 1999 987
rect 2003 983 2004 987
rect 1998 982 2004 983
rect 2008 985 2018 987
rect 2110 987 2116 988
rect 1646 971 1652 972
rect 1646 967 1647 971
rect 1651 967 1652 971
rect 1646 966 1652 967
rect 1654 971 1660 972
rect 1654 967 1655 971
rect 1659 967 1660 971
rect 1654 966 1660 967
rect 1583 946 1587 947
rect 1527 941 1531 942
rect 1534 943 1540 944
rect 1286 924 1292 925
rect 1262 923 1268 924
rect 1262 919 1263 923
rect 1267 919 1268 923
rect 1286 920 1287 924
rect 1291 920 1292 924
rect 1328 921 1330 941
rect 1368 922 1370 941
rect 1440 922 1442 941
rect 1528 922 1530 941
rect 1534 939 1535 943
rect 1539 939 1540 943
rect 1583 941 1587 942
rect 1615 946 1619 947
rect 1615 941 1619 942
rect 1639 946 1643 947
rect 1639 941 1643 942
rect 1534 938 1540 939
rect 1616 922 1618 941
rect 1366 921 1372 922
rect 1286 919 1292 920
rect 1326 920 1332 921
rect 1262 918 1268 919
rect 1326 916 1327 920
rect 1331 916 1332 920
rect 1366 917 1367 921
rect 1371 917 1372 921
rect 1366 916 1372 917
rect 1438 921 1444 922
rect 1438 917 1439 921
rect 1443 917 1444 921
rect 1438 916 1444 917
rect 1526 921 1532 922
rect 1526 917 1527 921
rect 1531 917 1532 921
rect 1614 921 1620 922
rect 1526 916 1532 917
rect 1566 919 1572 920
rect 1326 915 1332 916
rect 1566 915 1567 919
rect 1571 915 1572 919
rect 1614 917 1615 921
rect 1619 917 1620 921
rect 1656 920 1658 966
rect 1696 947 1698 982
rect 1752 947 1754 982
rect 1695 946 1699 947
rect 1695 941 1699 942
rect 1751 946 1755 947
rect 1751 941 1755 942
rect 1696 922 1698 941
rect 1784 936 1786 982
rect 1824 947 1826 982
rect 1904 947 1906 982
rect 2000 947 2002 982
rect 2008 976 2010 985
rect 2110 983 2111 987
rect 2115 983 2116 987
rect 2110 982 2116 983
rect 2230 987 2236 988
rect 2230 983 2231 987
rect 2235 983 2236 987
rect 2230 982 2236 983
rect 2246 987 2252 988
rect 2246 983 2247 987
rect 2251 983 2252 987
rect 2246 982 2252 983
rect 2350 987 2356 988
rect 2350 983 2351 987
rect 2355 983 2356 987
rect 2350 982 2356 983
rect 2430 987 2436 988
rect 2430 983 2431 987
rect 2435 983 2436 987
rect 2430 982 2436 983
rect 2454 987 2460 988
rect 2454 983 2455 987
rect 2459 983 2460 987
rect 2454 982 2460 983
rect 2006 975 2012 976
rect 2006 971 2007 975
rect 2011 971 2012 975
rect 2006 970 2012 971
rect 2112 947 2114 982
rect 2232 947 2234 982
rect 2248 968 2250 982
rect 2246 967 2252 968
rect 2246 963 2247 967
rect 2251 963 2252 967
rect 2246 962 2252 963
rect 2352 947 2354 982
rect 1791 946 1795 947
rect 1791 941 1795 942
rect 1823 946 1827 947
rect 1823 941 1827 942
rect 1895 946 1899 947
rect 1895 941 1899 942
rect 1903 946 1907 947
rect 1903 941 1907 942
rect 1999 946 2003 947
rect 1999 941 2003 942
rect 2015 946 2019 947
rect 2015 941 2019 942
rect 2111 946 2115 947
rect 2111 941 2115 942
rect 2151 946 2155 947
rect 2151 941 2155 942
rect 2231 946 2235 947
rect 2231 941 2235 942
rect 2295 946 2299 947
rect 2295 941 2299 942
rect 2351 946 2355 947
rect 2351 941 2355 942
rect 1722 935 1728 936
rect 1722 931 1723 935
rect 1727 931 1728 935
rect 1722 930 1728 931
rect 1782 935 1788 936
rect 1782 931 1783 935
rect 1787 931 1788 935
rect 1782 930 1788 931
rect 1694 921 1700 922
rect 1614 916 1620 917
rect 1654 919 1660 920
rect 1566 914 1572 915
rect 1654 915 1655 919
rect 1659 915 1660 919
rect 1694 917 1695 921
rect 1699 917 1700 921
rect 1694 916 1700 917
rect 1654 914 1660 915
rect 1286 907 1292 908
rect 1286 903 1287 907
rect 1291 903 1292 907
rect 1286 902 1292 903
rect 1326 903 1332 904
rect 1288 895 1290 902
rect 1326 899 1327 903
rect 1331 899 1332 903
rect 1326 898 1332 899
rect 1350 900 1356 901
rect 1287 894 1291 895
rect 1287 889 1291 890
rect 1288 886 1290 889
rect 1328 887 1330 898
rect 1350 896 1351 900
rect 1355 896 1356 900
rect 1350 895 1356 896
rect 1422 900 1428 901
rect 1422 896 1423 900
rect 1427 896 1428 900
rect 1422 895 1428 896
rect 1510 900 1516 901
rect 1510 896 1511 900
rect 1515 896 1516 900
rect 1510 895 1516 896
rect 1352 887 1354 895
rect 1424 887 1426 895
rect 1512 887 1514 895
rect 1327 886 1331 887
rect 1286 885 1292 886
rect 1286 881 1287 885
rect 1291 881 1292 885
rect 1327 881 1331 882
rect 1351 886 1355 887
rect 1351 881 1355 882
rect 1423 886 1427 887
rect 1423 881 1427 882
rect 1487 886 1491 887
rect 1487 881 1491 882
rect 1511 886 1515 887
rect 1511 881 1515 882
rect 1559 886 1563 887
rect 1559 881 1563 882
rect 1286 880 1292 881
rect 1328 878 1330 881
rect 1486 880 1492 881
rect 1326 877 1332 878
rect 1326 873 1327 877
rect 1331 873 1332 877
rect 1486 876 1487 880
rect 1491 876 1492 880
rect 1486 875 1492 876
rect 1558 880 1564 881
rect 1558 876 1559 880
rect 1563 876 1564 880
rect 1558 875 1564 876
rect 1326 872 1332 873
rect 1286 868 1292 869
rect 1182 867 1188 868
rect 1182 863 1183 867
rect 1187 863 1188 867
rect 1182 862 1188 863
rect 1238 867 1244 868
rect 1238 863 1239 867
rect 1243 863 1244 867
rect 1238 862 1244 863
rect 1246 867 1252 868
rect 1246 863 1247 867
rect 1251 863 1252 867
rect 1286 864 1287 868
rect 1291 864 1292 868
rect 1286 863 1292 864
rect 1246 862 1252 863
rect 1118 847 1124 848
rect 1118 843 1119 847
rect 1123 843 1124 847
rect 1118 842 1124 843
rect 1184 839 1186 862
rect 1240 839 1242 862
rect 1288 839 1290 863
rect 1326 860 1332 861
rect 1326 856 1327 860
rect 1331 856 1332 860
rect 1326 855 1332 856
rect 1502 859 1508 860
rect 1502 855 1503 859
rect 1507 855 1508 859
rect 727 838 731 839
rect 727 833 731 834
rect 759 838 763 839
rect 759 833 763 834
rect 807 838 811 839
rect 807 833 811 834
rect 855 838 859 839
rect 855 833 859 834
rect 895 838 899 839
rect 895 833 899 834
rect 943 838 947 839
rect 943 833 947 834
rect 983 838 987 839
rect 983 833 987 834
rect 1023 838 1027 839
rect 1023 833 1027 834
rect 1071 838 1075 839
rect 1090 835 1091 839
rect 1095 835 1096 839
rect 1090 834 1096 835
rect 1103 838 1107 839
rect 1071 833 1075 834
rect 670 827 676 828
rect 670 823 671 827
rect 675 823 676 827
rect 670 822 676 823
rect 728 814 730 833
rect 762 827 768 828
rect 762 823 763 827
rect 767 823 768 827
rect 762 822 768 823
rect 462 813 468 814
rect 382 808 388 809
rect 402 811 408 812
rect 350 806 356 807
rect 402 807 403 811
rect 407 807 408 811
rect 462 809 463 813
rect 467 809 468 813
rect 462 808 468 809
rect 550 813 556 814
rect 550 809 551 813
rect 555 809 556 813
rect 550 808 556 809
rect 638 813 644 814
rect 638 809 639 813
rect 643 809 644 813
rect 638 808 644 809
rect 726 813 732 814
rect 726 809 727 813
rect 731 809 732 813
rect 726 808 732 809
rect 402 806 408 807
rect 110 795 116 796
rect 110 791 111 795
rect 115 791 116 795
rect 110 790 116 791
rect 222 792 228 793
rect 112 783 114 790
rect 222 788 223 792
rect 227 788 228 792
rect 222 787 228 788
rect 286 792 292 793
rect 286 788 287 792
rect 291 788 292 792
rect 286 787 292 788
rect 224 783 226 787
rect 288 783 290 787
rect 111 782 115 783
rect 111 777 115 778
rect 151 782 155 783
rect 151 777 155 778
rect 223 782 227 783
rect 223 777 227 778
rect 247 782 251 783
rect 247 777 251 778
rect 287 782 291 783
rect 287 777 291 778
rect 343 782 347 783
rect 343 777 347 778
rect 112 774 114 777
rect 150 776 156 777
rect 110 773 116 774
rect 110 769 111 773
rect 115 769 116 773
rect 150 772 151 776
rect 155 772 156 776
rect 150 771 156 772
rect 246 776 252 777
rect 246 772 247 776
rect 251 772 252 776
rect 246 771 252 772
rect 342 776 348 777
rect 342 772 343 776
rect 347 772 348 776
rect 342 771 348 772
rect 110 768 116 769
rect 110 756 116 757
rect 110 752 111 756
rect 115 752 116 756
rect 110 751 116 752
rect 166 755 172 756
rect 166 751 167 755
rect 171 751 172 755
rect 112 727 114 751
rect 166 750 172 751
rect 182 755 188 756
rect 182 751 183 755
rect 187 751 188 755
rect 182 750 188 751
rect 262 755 268 756
rect 262 751 263 755
rect 267 751 268 755
rect 262 750 268 751
rect 278 755 284 756
rect 278 751 279 755
rect 283 751 284 755
rect 278 750 284 751
rect 168 727 170 750
rect 111 726 115 727
rect 111 721 115 722
rect 167 726 171 727
rect 167 721 171 722
rect 175 726 179 727
rect 175 721 179 722
rect 112 701 114 721
rect 176 702 178 721
rect 184 716 186 750
rect 264 727 266 750
rect 280 736 282 750
rect 352 740 354 806
rect 366 792 372 793
rect 366 788 367 792
rect 371 788 372 792
rect 366 787 372 788
rect 446 792 452 793
rect 446 788 447 792
rect 451 788 452 792
rect 446 787 452 788
rect 534 792 540 793
rect 534 788 535 792
rect 539 788 540 792
rect 534 787 540 788
rect 622 792 628 793
rect 622 788 623 792
rect 627 788 628 792
rect 622 787 628 788
rect 710 792 716 793
rect 710 788 711 792
rect 715 788 716 792
rect 710 787 716 788
rect 368 783 370 787
rect 448 783 450 787
rect 536 783 538 787
rect 624 783 626 787
rect 712 783 714 787
rect 764 784 766 822
rect 808 814 810 833
rect 896 814 898 833
rect 984 814 986 833
rect 1072 814 1074 833
rect 806 813 812 814
rect 806 809 807 813
rect 811 809 812 813
rect 806 808 812 809
rect 894 813 900 814
rect 894 809 895 813
rect 899 809 900 813
rect 894 808 900 809
rect 982 813 988 814
rect 982 809 983 813
rect 987 809 988 813
rect 982 808 988 809
rect 1070 813 1076 814
rect 1070 809 1071 813
rect 1075 809 1076 813
rect 1092 812 1094 834
rect 1103 833 1107 834
rect 1183 838 1187 839
rect 1183 833 1187 834
rect 1239 838 1243 839
rect 1239 833 1243 834
rect 1287 838 1291 839
rect 1287 833 1291 834
rect 1288 813 1290 833
rect 1328 827 1330 855
rect 1502 854 1508 855
rect 1518 859 1524 860
rect 1518 855 1519 859
rect 1523 855 1524 859
rect 1518 854 1524 855
rect 1504 827 1506 854
rect 1327 826 1331 827
rect 1327 821 1331 822
rect 1439 826 1443 827
rect 1439 821 1443 822
rect 1503 826 1507 827
rect 1503 821 1507 822
rect 1511 826 1515 827
rect 1520 824 1522 854
rect 1568 844 1570 914
rect 1598 900 1604 901
rect 1598 896 1599 900
rect 1603 896 1604 900
rect 1598 895 1604 896
rect 1678 900 1684 901
rect 1678 896 1679 900
rect 1683 896 1684 900
rect 1678 895 1684 896
rect 1600 887 1602 895
rect 1680 887 1682 895
rect 1599 886 1603 887
rect 1599 881 1603 882
rect 1623 886 1627 887
rect 1623 881 1627 882
rect 1679 886 1683 887
rect 1679 881 1683 882
rect 1687 886 1691 887
rect 1687 881 1691 882
rect 1622 880 1628 881
rect 1622 876 1623 880
rect 1627 876 1628 880
rect 1622 875 1628 876
rect 1686 880 1692 881
rect 1686 876 1687 880
rect 1691 876 1692 880
rect 1686 875 1692 876
rect 1724 860 1726 930
rect 1792 922 1794 941
rect 1896 922 1898 941
rect 2016 922 2018 941
rect 2152 922 2154 941
rect 2296 922 2298 941
rect 2406 935 2412 936
rect 2406 931 2407 935
rect 2411 931 2412 935
rect 2406 930 2412 931
rect 1790 921 1796 922
rect 1790 917 1791 921
rect 1795 917 1796 921
rect 1790 916 1796 917
rect 1894 921 1900 922
rect 1894 917 1895 921
rect 1899 917 1900 921
rect 1894 916 1900 917
rect 2014 921 2020 922
rect 2014 917 2015 921
rect 2019 917 2020 921
rect 2014 916 2020 917
rect 2150 921 2156 922
rect 2150 917 2151 921
rect 2155 917 2156 921
rect 2150 916 2156 917
rect 2294 921 2300 922
rect 2294 917 2295 921
rect 2299 917 2300 921
rect 2294 916 2300 917
rect 2302 919 2308 920
rect 2302 915 2303 919
rect 2307 915 2308 919
rect 2302 914 2308 915
rect 1774 900 1780 901
rect 1774 896 1775 900
rect 1779 896 1780 900
rect 1774 895 1780 896
rect 1878 900 1884 901
rect 1878 896 1879 900
rect 1883 896 1884 900
rect 1878 895 1884 896
rect 1998 900 2004 901
rect 1998 896 1999 900
rect 2003 896 2004 900
rect 1998 895 2004 896
rect 2134 900 2140 901
rect 2134 896 2135 900
rect 2139 896 2140 900
rect 2134 895 2140 896
rect 2278 900 2284 901
rect 2278 896 2279 900
rect 2283 896 2284 900
rect 2278 895 2284 896
rect 1776 887 1778 895
rect 1880 887 1882 895
rect 2000 887 2002 895
rect 2136 887 2138 895
rect 2280 887 2282 895
rect 1751 886 1755 887
rect 1751 881 1755 882
rect 1775 886 1779 887
rect 1775 881 1779 882
rect 1815 886 1819 887
rect 1815 881 1819 882
rect 1879 886 1883 887
rect 1879 881 1883 882
rect 1887 886 1891 887
rect 1887 881 1891 882
rect 1975 886 1979 887
rect 1975 881 1979 882
rect 1999 886 2003 887
rect 1999 881 2003 882
rect 2079 886 2083 887
rect 2079 881 2083 882
rect 2135 886 2139 887
rect 2135 881 2139 882
rect 2199 886 2203 887
rect 2199 881 2203 882
rect 2279 886 2283 887
rect 2279 881 2283 882
rect 1750 880 1756 881
rect 1750 876 1751 880
rect 1755 876 1756 880
rect 1750 875 1756 876
rect 1814 880 1820 881
rect 1814 876 1815 880
rect 1819 876 1820 880
rect 1814 875 1820 876
rect 1886 880 1892 881
rect 1886 876 1887 880
rect 1891 876 1892 880
rect 1886 875 1892 876
rect 1974 880 1980 881
rect 1974 876 1975 880
rect 1979 876 1980 880
rect 1974 875 1980 876
rect 2078 880 2084 881
rect 2078 876 2079 880
rect 2083 876 2084 880
rect 2078 875 2084 876
rect 2198 880 2204 881
rect 2198 876 2199 880
rect 2203 876 2204 880
rect 2198 875 2204 876
rect 1574 859 1580 860
rect 1574 855 1575 859
rect 1579 855 1580 859
rect 1574 854 1580 855
rect 1638 859 1644 860
rect 1638 855 1639 859
rect 1643 855 1644 859
rect 1638 854 1644 855
rect 1646 859 1652 860
rect 1646 855 1647 859
rect 1651 855 1652 859
rect 1646 854 1652 855
rect 1702 859 1708 860
rect 1702 855 1703 859
rect 1707 855 1708 859
rect 1702 854 1708 855
rect 1722 859 1728 860
rect 1722 855 1723 859
rect 1727 855 1728 859
rect 1722 854 1728 855
rect 1766 859 1772 860
rect 1766 855 1767 859
rect 1771 855 1772 859
rect 1766 854 1772 855
rect 1830 859 1836 860
rect 1830 855 1831 859
rect 1835 855 1836 859
rect 1830 854 1836 855
rect 1902 859 1908 860
rect 1902 855 1903 859
rect 1907 855 1908 859
rect 1902 854 1908 855
rect 1990 859 1996 860
rect 1990 855 1991 859
rect 1995 855 1996 859
rect 1990 854 1996 855
rect 2094 859 2100 860
rect 2094 855 2095 859
rect 2099 855 2100 859
rect 2094 854 2100 855
rect 2214 859 2220 860
rect 2214 855 2215 859
rect 2219 855 2220 859
rect 2214 854 2220 855
rect 1566 843 1572 844
rect 1566 839 1567 843
rect 1571 839 1572 843
rect 1566 838 1572 839
rect 1576 827 1578 854
rect 1640 827 1642 854
rect 1648 836 1650 854
rect 1646 835 1652 836
rect 1646 831 1647 835
rect 1651 831 1652 835
rect 1646 830 1652 831
rect 1704 827 1706 854
rect 1768 827 1770 854
rect 1818 843 1824 844
rect 1818 839 1819 843
rect 1823 839 1824 843
rect 1818 838 1824 839
rect 1575 826 1579 827
rect 1511 821 1515 822
rect 1518 823 1524 824
rect 1286 812 1292 813
rect 1070 808 1076 809
rect 1090 811 1096 812
rect 1090 807 1091 811
rect 1095 807 1096 811
rect 1286 808 1287 812
rect 1291 808 1292 812
rect 1286 807 1292 808
rect 1090 806 1096 807
rect 1328 801 1330 821
rect 1440 802 1442 821
rect 1512 802 1514 821
rect 1518 819 1519 823
rect 1523 819 1524 823
rect 1575 821 1579 822
rect 1591 826 1595 827
rect 1591 821 1595 822
rect 1639 826 1643 827
rect 1639 821 1643 822
rect 1671 826 1675 827
rect 1671 821 1675 822
rect 1703 826 1707 827
rect 1759 826 1763 827
rect 1703 821 1707 822
rect 1722 823 1728 824
rect 1518 818 1524 819
rect 1592 802 1594 821
rect 1672 802 1674 821
rect 1722 819 1723 823
rect 1727 819 1728 823
rect 1759 821 1763 822
rect 1767 826 1771 827
rect 1767 821 1771 822
rect 1722 818 1728 819
rect 1438 801 1444 802
rect 1326 800 1332 801
rect 1326 796 1327 800
rect 1331 796 1332 800
rect 1438 797 1439 801
rect 1443 797 1444 801
rect 1438 796 1444 797
rect 1510 801 1516 802
rect 1510 797 1511 801
rect 1515 797 1516 801
rect 1510 796 1516 797
rect 1590 801 1596 802
rect 1590 797 1591 801
rect 1595 797 1596 801
rect 1670 801 1676 802
rect 1590 796 1596 797
rect 1598 799 1604 800
rect 1286 795 1292 796
rect 1326 795 1332 796
rect 1598 795 1599 799
rect 1603 795 1604 799
rect 1670 797 1671 801
rect 1675 797 1676 801
rect 1670 796 1676 797
rect 790 792 796 793
rect 790 788 791 792
rect 795 788 796 792
rect 790 787 796 788
rect 878 792 884 793
rect 878 788 879 792
rect 883 788 884 792
rect 878 787 884 788
rect 966 792 972 793
rect 966 788 967 792
rect 971 788 972 792
rect 966 787 972 788
rect 1054 792 1060 793
rect 1054 788 1055 792
rect 1059 788 1060 792
rect 1286 791 1287 795
rect 1291 791 1292 795
rect 1598 794 1604 795
rect 1286 790 1292 791
rect 1054 787 1060 788
rect 762 783 768 784
rect 792 783 794 787
rect 880 783 882 787
rect 968 783 970 787
rect 1010 783 1016 784
rect 1056 783 1058 787
rect 1288 783 1290 790
rect 1326 783 1332 784
rect 367 782 371 783
rect 367 777 371 778
rect 439 782 443 783
rect 439 777 443 778
rect 447 782 451 783
rect 447 777 451 778
rect 527 782 531 783
rect 527 777 531 778
rect 535 782 539 783
rect 535 777 539 778
rect 607 782 611 783
rect 607 777 611 778
rect 623 782 627 783
rect 623 777 627 778
rect 679 782 683 783
rect 679 777 683 778
rect 711 782 715 783
rect 711 777 715 778
rect 751 782 755 783
rect 762 779 763 783
rect 767 779 768 783
rect 762 778 768 779
rect 791 782 795 783
rect 751 777 755 778
rect 791 777 795 778
rect 823 782 827 783
rect 823 777 827 778
rect 879 782 883 783
rect 879 777 883 778
rect 895 782 899 783
rect 895 777 899 778
rect 967 782 971 783
rect 967 777 971 778
rect 975 782 979 783
rect 1010 779 1011 783
rect 1015 779 1016 783
rect 1010 778 1016 779
rect 1055 782 1059 783
rect 975 777 979 778
rect 438 776 444 777
rect 438 772 439 776
rect 443 772 444 776
rect 438 771 444 772
rect 526 776 532 777
rect 526 772 527 776
rect 531 772 532 776
rect 526 771 532 772
rect 606 776 612 777
rect 606 772 607 776
rect 611 772 612 776
rect 606 771 612 772
rect 678 776 684 777
rect 678 772 679 776
rect 683 772 684 776
rect 678 771 684 772
rect 750 776 756 777
rect 750 772 751 776
rect 755 772 756 776
rect 750 771 756 772
rect 822 776 828 777
rect 822 772 823 776
rect 827 772 828 776
rect 822 771 828 772
rect 894 776 900 777
rect 894 772 895 776
rect 899 772 900 776
rect 894 771 900 772
rect 974 776 980 777
rect 974 772 975 776
rect 979 772 980 776
rect 974 771 980 772
rect 1012 756 1014 778
rect 1055 777 1059 778
rect 1287 782 1291 783
rect 1326 779 1327 783
rect 1331 779 1332 783
rect 1326 778 1332 779
rect 1422 780 1428 781
rect 1287 777 1291 778
rect 1288 774 1290 777
rect 1286 773 1292 774
rect 1286 769 1287 773
rect 1291 769 1292 773
rect 1328 771 1330 778
rect 1422 776 1423 780
rect 1427 776 1428 780
rect 1422 775 1428 776
rect 1494 780 1500 781
rect 1494 776 1495 780
rect 1499 776 1500 780
rect 1494 775 1500 776
rect 1574 780 1580 781
rect 1574 776 1575 780
rect 1579 776 1580 780
rect 1574 775 1580 776
rect 1424 771 1426 775
rect 1496 771 1498 775
rect 1576 771 1578 775
rect 1286 768 1292 769
rect 1327 770 1331 771
rect 1327 765 1331 766
rect 1351 770 1355 771
rect 1351 765 1355 766
rect 1423 770 1427 771
rect 1423 765 1427 766
rect 1447 770 1451 771
rect 1447 765 1451 766
rect 1495 770 1499 771
rect 1495 765 1499 766
rect 1567 770 1571 771
rect 1567 765 1571 766
rect 1575 770 1579 771
rect 1575 765 1579 766
rect 1328 762 1330 765
rect 1350 764 1356 765
rect 1326 761 1332 762
rect 1326 757 1327 761
rect 1331 757 1332 761
rect 1350 760 1351 764
rect 1355 760 1356 764
rect 1350 759 1356 760
rect 1446 764 1452 765
rect 1446 760 1447 764
rect 1451 760 1452 764
rect 1446 759 1452 760
rect 1566 764 1572 765
rect 1566 760 1567 764
rect 1571 760 1572 764
rect 1566 759 1572 760
rect 1286 756 1292 757
rect 1326 756 1332 757
rect 358 755 364 756
rect 358 751 359 755
rect 363 751 364 755
rect 358 750 364 751
rect 454 755 460 756
rect 454 751 455 755
rect 459 751 460 755
rect 454 750 460 751
rect 542 755 548 756
rect 542 751 543 755
rect 547 751 548 755
rect 542 750 548 751
rect 566 755 572 756
rect 566 751 567 755
rect 571 751 572 755
rect 566 750 572 751
rect 622 755 628 756
rect 622 751 623 755
rect 627 751 628 755
rect 622 750 628 751
rect 694 755 700 756
rect 694 751 695 755
rect 699 751 700 755
rect 694 750 700 751
rect 766 755 772 756
rect 766 751 767 755
rect 771 751 772 755
rect 766 750 772 751
rect 838 755 844 756
rect 838 751 839 755
rect 843 751 844 755
rect 838 750 844 751
rect 910 755 916 756
rect 910 751 911 755
rect 915 751 916 755
rect 910 750 916 751
rect 990 755 996 756
rect 990 751 991 755
rect 995 751 996 755
rect 990 750 996 751
rect 1010 755 1016 756
rect 1010 751 1011 755
rect 1015 751 1016 755
rect 1286 752 1287 756
rect 1291 752 1292 756
rect 1286 751 1292 752
rect 1010 750 1016 751
rect 350 739 356 740
rect 278 735 284 736
rect 278 731 279 735
rect 283 731 284 735
rect 350 735 351 739
rect 355 735 356 739
rect 350 734 356 735
rect 278 730 284 731
rect 360 727 362 750
rect 374 739 380 740
rect 374 735 375 739
rect 379 735 380 739
rect 374 734 380 735
rect 263 726 267 727
rect 263 721 267 722
rect 343 726 347 727
rect 343 721 347 722
rect 359 726 363 727
rect 359 721 363 722
rect 182 715 188 716
rect 182 711 183 715
rect 187 711 188 715
rect 182 710 188 711
rect 264 702 266 721
rect 310 715 316 716
rect 310 711 311 715
rect 315 711 316 715
rect 310 710 316 711
rect 174 701 180 702
rect 110 700 116 701
rect 110 696 111 700
rect 115 696 116 700
rect 174 697 175 701
rect 179 697 180 701
rect 262 701 268 702
rect 174 696 180 697
rect 222 699 228 700
rect 110 695 116 696
rect 222 695 223 699
rect 227 695 228 699
rect 262 697 263 701
rect 267 697 268 701
rect 262 696 268 697
rect 222 694 228 695
rect 110 683 116 684
rect 110 679 111 683
rect 115 679 116 683
rect 110 678 116 679
rect 158 680 164 681
rect 112 675 114 678
rect 158 676 159 680
rect 163 676 164 680
rect 158 675 164 676
rect 111 674 115 675
rect 111 669 115 670
rect 159 674 163 675
rect 159 669 163 670
rect 215 674 219 675
rect 215 669 219 670
rect 112 666 114 669
rect 214 668 220 669
rect 110 665 116 666
rect 110 661 111 665
rect 115 661 116 665
rect 214 664 215 668
rect 219 664 220 668
rect 214 663 220 664
rect 110 660 116 661
rect 110 648 116 649
rect 110 644 111 648
rect 115 644 116 648
rect 110 643 116 644
rect 112 619 114 643
rect 224 632 226 694
rect 246 680 252 681
rect 246 676 247 680
rect 251 676 252 680
rect 246 675 252 676
rect 247 674 251 675
rect 247 669 251 670
rect 295 674 299 675
rect 295 669 299 670
rect 294 668 300 669
rect 294 664 295 668
rect 299 664 300 668
rect 294 663 300 664
rect 312 659 314 710
rect 344 702 346 721
rect 342 701 348 702
rect 342 697 343 701
rect 347 697 348 701
rect 376 700 378 734
rect 456 727 458 750
rect 544 727 546 750
rect 423 726 427 727
rect 423 721 427 722
rect 455 726 459 727
rect 455 721 459 722
rect 503 726 507 727
rect 503 721 507 722
rect 543 726 547 727
rect 543 721 547 722
rect 424 702 426 721
rect 504 702 506 721
rect 568 716 570 750
rect 624 727 626 750
rect 696 727 698 750
rect 768 727 770 750
rect 840 727 842 750
rect 912 727 914 750
rect 930 735 936 736
rect 930 731 931 735
rect 935 731 936 735
rect 930 730 936 731
rect 575 726 579 727
rect 623 726 627 727
rect 575 721 579 722
rect 594 723 600 724
rect 566 715 572 716
rect 566 711 567 715
rect 571 711 572 715
rect 566 710 572 711
rect 576 702 578 721
rect 594 719 595 723
rect 599 719 600 723
rect 623 721 627 722
rect 639 726 643 727
rect 639 721 643 722
rect 695 726 699 727
rect 695 721 699 722
rect 703 726 707 727
rect 703 721 707 722
rect 767 726 771 727
rect 767 721 771 722
rect 839 726 843 727
rect 839 721 843 722
rect 911 726 915 727
rect 911 721 915 722
rect 594 718 600 719
rect 422 701 428 702
rect 342 696 348 697
rect 374 699 380 700
rect 374 695 375 699
rect 379 695 380 699
rect 422 697 423 701
rect 427 697 428 701
rect 422 696 428 697
rect 502 701 508 702
rect 502 697 503 701
rect 507 697 508 701
rect 574 701 580 702
rect 502 696 508 697
rect 534 699 540 700
rect 374 694 380 695
rect 534 695 535 699
rect 539 695 540 699
rect 574 697 575 701
rect 579 697 580 701
rect 596 700 598 718
rect 630 715 636 716
rect 630 711 631 715
rect 635 711 636 715
rect 630 710 636 711
rect 574 696 580 697
rect 594 699 600 700
rect 534 694 540 695
rect 594 695 595 699
rect 599 695 600 699
rect 594 694 600 695
rect 326 680 332 681
rect 326 676 327 680
rect 331 676 332 680
rect 326 675 332 676
rect 406 680 412 681
rect 406 676 407 680
rect 411 676 412 680
rect 406 675 412 676
rect 486 680 492 681
rect 486 676 487 680
rect 491 676 492 680
rect 486 675 492 676
rect 327 674 331 675
rect 327 669 331 670
rect 375 674 379 675
rect 375 669 379 670
rect 407 674 411 675
rect 407 669 411 670
rect 455 674 459 675
rect 455 669 459 670
rect 487 674 491 675
rect 487 669 491 670
rect 527 674 531 675
rect 527 669 531 670
rect 374 668 380 669
rect 374 664 375 668
rect 379 664 380 668
rect 374 663 380 664
rect 454 668 460 669
rect 454 664 455 668
rect 459 664 460 668
rect 454 663 460 664
rect 526 668 532 669
rect 526 664 527 668
rect 531 664 532 668
rect 526 663 532 664
rect 312 657 322 659
rect 320 648 322 657
rect 230 647 236 648
rect 230 643 231 647
rect 235 643 236 647
rect 230 642 236 643
rect 294 647 300 648
rect 294 643 295 647
rect 299 643 300 647
rect 294 642 300 643
rect 310 647 316 648
rect 310 643 311 647
rect 315 643 316 647
rect 310 642 316 643
rect 318 647 324 648
rect 318 643 319 647
rect 323 643 324 647
rect 318 642 324 643
rect 390 647 396 648
rect 390 643 391 647
rect 395 643 396 647
rect 390 642 396 643
rect 470 647 476 648
rect 470 643 471 647
rect 475 643 476 647
rect 470 642 476 643
rect 494 647 500 648
rect 494 643 495 647
rect 499 643 500 647
rect 494 642 500 643
rect 222 631 228 632
rect 222 627 223 631
rect 227 627 228 631
rect 222 626 228 627
rect 232 619 234 642
rect 111 618 115 619
rect 111 613 115 614
rect 207 618 211 619
rect 207 613 211 614
rect 231 618 235 619
rect 231 613 235 614
rect 112 593 114 613
rect 208 594 210 613
rect 296 608 298 642
rect 312 619 314 642
rect 392 619 394 642
rect 426 631 432 632
rect 426 627 427 631
rect 431 627 432 631
rect 426 626 432 627
rect 303 618 307 619
rect 303 613 307 614
rect 311 618 315 619
rect 311 613 315 614
rect 391 618 395 619
rect 391 613 395 614
rect 407 618 411 619
rect 407 613 411 614
rect 294 607 300 608
rect 294 603 295 607
rect 299 603 300 607
rect 294 602 300 603
rect 304 594 306 613
rect 408 594 410 613
rect 414 607 420 608
rect 414 603 415 607
rect 419 603 420 607
rect 414 602 420 603
rect 206 593 212 594
rect 110 592 116 593
rect 110 588 111 592
rect 115 588 116 592
rect 206 589 207 593
rect 211 589 212 593
rect 302 593 308 594
rect 206 588 212 589
rect 214 591 220 592
rect 110 587 116 588
rect 214 587 215 591
rect 219 587 220 591
rect 302 589 303 593
rect 307 589 308 593
rect 302 588 308 589
rect 406 593 412 594
rect 406 589 407 593
rect 411 589 412 593
rect 406 588 412 589
rect 214 586 220 587
rect 110 575 116 576
rect 110 571 111 575
rect 115 571 116 575
rect 110 570 116 571
rect 190 572 196 573
rect 112 563 114 570
rect 190 568 191 572
rect 195 568 196 572
rect 190 567 196 568
rect 192 563 194 567
rect 111 562 115 563
rect 111 557 115 558
rect 175 562 179 563
rect 175 557 179 558
rect 191 562 195 563
rect 191 557 195 558
rect 112 554 114 557
rect 174 556 180 557
rect 110 553 116 554
rect 110 549 111 553
rect 115 549 116 553
rect 174 552 175 556
rect 179 552 180 556
rect 174 551 180 552
rect 110 548 116 549
rect 110 536 116 537
rect 110 532 111 536
rect 115 532 116 536
rect 110 531 116 532
rect 190 535 196 536
rect 190 531 191 535
rect 195 531 196 535
rect 112 507 114 531
rect 190 530 196 531
rect 192 507 194 530
rect 216 520 218 586
rect 286 572 292 573
rect 286 568 287 572
rect 291 568 292 572
rect 286 567 292 568
rect 390 572 396 573
rect 390 568 391 572
rect 395 568 396 572
rect 390 567 396 568
rect 288 563 290 567
rect 392 563 394 567
rect 271 562 275 563
rect 271 557 275 558
rect 287 562 291 563
rect 287 557 291 558
rect 375 562 379 563
rect 375 557 379 558
rect 391 562 395 563
rect 391 557 395 558
rect 270 556 276 557
rect 270 552 271 556
rect 275 552 276 556
rect 270 551 276 552
rect 374 556 380 557
rect 374 552 375 556
rect 379 552 380 556
rect 374 551 380 552
rect 416 536 418 602
rect 428 592 430 626
rect 472 619 474 642
rect 471 618 475 619
rect 471 613 475 614
rect 496 608 498 642
rect 536 632 538 694
rect 558 680 564 681
rect 558 676 559 680
rect 563 676 564 680
rect 558 675 564 676
rect 622 680 628 681
rect 622 676 623 680
rect 627 676 628 680
rect 622 675 628 676
rect 559 674 563 675
rect 559 669 563 670
rect 591 674 595 675
rect 591 669 595 670
rect 623 674 627 675
rect 623 669 627 670
rect 590 668 596 669
rect 590 664 591 668
rect 595 664 596 668
rect 590 663 596 664
rect 632 648 634 710
rect 640 702 642 721
rect 704 702 706 721
rect 768 702 770 721
rect 840 702 842 721
rect 912 702 914 721
rect 638 701 644 702
rect 638 697 639 701
rect 643 697 644 701
rect 638 696 644 697
rect 702 701 708 702
rect 702 697 703 701
rect 707 697 708 701
rect 702 696 708 697
rect 766 701 772 702
rect 766 697 767 701
rect 771 697 772 701
rect 766 696 772 697
rect 838 701 844 702
rect 838 697 839 701
rect 843 697 844 701
rect 838 696 844 697
rect 910 701 916 702
rect 910 697 911 701
rect 915 697 916 701
rect 932 700 934 730
rect 992 727 994 750
rect 1288 727 1290 751
rect 1326 744 1332 745
rect 1326 740 1327 744
rect 1331 740 1332 744
rect 1326 739 1332 740
rect 1366 743 1372 744
rect 1366 739 1367 743
rect 1371 739 1372 743
rect 991 726 995 727
rect 991 721 995 722
rect 1287 726 1291 727
rect 1287 721 1291 722
rect 1288 701 1290 721
rect 1328 715 1330 739
rect 1366 738 1372 739
rect 1374 743 1380 744
rect 1374 739 1375 743
rect 1379 739 1380 743
rect 1374 738 1380 739
rect 1462 743 1468 744
rect 1462 739 1463 743
rect 1467 739 1468 743
rect 1462 738 1468 739
rect 1582 743 1588 744
rect 1582 739 1583 743
rect 1587 739 1588 743
rect 1582 738 1588 739
rect 1368 715 1370 738
rect 1327 714 1331 715
rect 1327 709 1331 710
rect 1367 714 1371 715
rect 1367 709 1371 710
rect 1286 700 1292 701
rect 910 696 916 697
rect 930 699 936 700
rect 930 695 931 699
rect 935 695 936 699
rect 1286 696 1287 700
rect 1291 696 1292 700
rect 1286 695 1292 696
rect 930 694 936 695
rect 1328 689 1330 709
rect 1368 690 1370 709
rect 1376 704 1378 738
rect 1464 715 1466 738
rect 1584 715 1586 738
rect 1600 728 1602 794
rect 1654 780 1660 781
rect 1654 776 1655 780
rect 1659 776 1660 780
rect 1654 775 1660 776
rect 1656 771 1658 775
rect 1655 770 1659 771
rect 1655 765 1659 766
rect 1687 770 1691 771
rect 1687 765 1691 766
rect 1686 764 1692 765
rect 1686 760 1687 764
rect 1691 760 1692 764
rect 1686 759 1692 760
rect 1724 744 1726 818
rect 1760 802 1762 821
rect 1820 808 1822 838
rect 1832 827 1834 854
rect 1839 852 1843 853
rect 1839 847 1843 848
rect 1840 844 1842 847
rect 1838 843 1844 844
rect 1838 839 1839 843
rect 1843 839 1844 843
rect 1838 838 1844 839
rect 1904 827 1906 854
rect 1992 827 1994 854
rect 2096 827 2098 854
rect 2216 827 2218 854
rect 2304 853 2306 914
rect 2319 886 2323 887
rect 2319 881 2323 882
rect 2318 880 2324 881
rect 2318 876 2319 880
rect 2323 876 2324 880
rect 2318 875 2324 876
rect 2334 859 2340 860
rect 2334 855 2335 859
rect 2339 855 2340 859
rect 2334 854 2340 855
rect 2342 859 2348 860
rect 2342 855 2343 859
rect 2347 855 2348 859
rect 2342 854 2348 855
rect 2303 852 2307 853
rect 2303 847 2307 848
rect 2336 827 2338 854
rect 1831 826 1835 827
rect 1831 821 1835 822
rect 1847 826 1851 827
rect 1847 821 1851 822
rect 1903 826 1907 827
rect 1903 821 1907 822
rect 1935 826 1939 827
rect 1935 821 1939 822
rect 1991 826 1995 827
rect 1991 821 1995 822
rect 2023 826 2027 827
rect 2023 821 2027 822
rect 2095 826 2099 827
rect 2095 821 2099 822
rect 2111 826 2115 827
rect 2111 821 2115 822
rect 2199 826 2203 827
rect 2199 821 2203 822
rect 2215 826 2219 827
rect 2215 821 2219 822
rect 2287 826 2291 827
rect 2287 821 2291 822
rect 2335 826 2339 827
rect 2344 824 2346 854
rect 2383 826 2387 827
rect 2335 821 2339 822
rect 2342 823 2348 824
rect 1818 807 1824 808
rect 1818 803 1819 807
rect 1823 803 1824 807
rect 1818 802 1824 803
rect 1848 802 1850 821
rect 1936 802 1938 821
rect 2024 802 2026 821
rect 2112 802 2114 821
rect 2200 802 2202 821
rect 2288 802 2290 821
rect 2342 819 2343 823
rect 2347 819 2348 823
rect 2383 821 2387 822
rect 2342 818 2348 819
rect 2384 802 2386 821
rect 2390 815 2396 816
rect 2390 811 2391 815
rect 2395 811 2396 815
rect 2390 810 2396 811
rect 1758 801 1764 802
rect 1758 797 1759 801
rect 1763 797 1764 801
rect 1758 796 1764 797
rect 1846 801 1852 802
rect 1846 797 1847 801
rect 1851 797 1852 801
rect 1846 796 1852 797
rect 1934 801 1940 802
rect 1934 797 1935 801
rect 1939 797 1940 801
rect 1934 796 1940 797
rect 2022 801 2028 802
rect 2022 797 2023 801
rect 2027 797 2028 801
rect 2022 796 2028 797
rect 2110 801 2116 802
rect 2110 797 2111 801
rect 2115 797 2116 801
rect 2110 796 2116 797
rect 2198 801 2204 802
rect 2198 797 2199 801
rect 2203 797 2204 801
rect 2198 796 2204 797
rect 2286 801 2292 802
rect 2286 797 2287 801
rect 2291 797 2292 801
rect 2382 801 2388 802
rect 2286 796 2292 797
rect 2294 799 2300 800
rect 2294 795 2295 799
rect 2299 795 2300 799
rect 2382 797 2383 801
rect 2387 797 2388 801
rect 2382 796 2388 797
rect 2294 794 2300 795
rect 1742 780 1748 781
rect 1742 776 1743 780
rect 1747 776 1748 780
rect 1742 775 1748 776
rect 1830 780 1836 781
rect 1830 776 1831 780
rect 1835 776 1836 780
rect 1830 775 1836 776
rect 1918 780 1924 781
rect 1918 776 1919 780
rect 1923 776 1924 780
rect 1918 775 1924 776
rect 2006 780 2012 781
rect 2006 776 2007 780
rect 2011 776 2012 780
rect 2006 775 2012 776
rect 2094 780 2100 781
rect 2094 776 2095 780
rect 2099 776 2100 780
rect 2094 775 2100 776
rect 2182 780 2188 781
rect 2182 776 2183 780
rect 2187 776 2188 780
rect 2182 775 2188 776
rect 2270 780 2276 781
rect 2270 776 2271 780
rect 2275 776 2276 780
rect 2270 775 2276 776
rect 1744 771 1746 775
rect 1832 771 1834 775
rect 1920 771 1922 775
rect 2008 771 2010 775
rect 2096 771 2098 775
rect 2184 771 2186 775
rect 2272 771 2274 775
rect 1743 770 1747 771
rect 1743 765 1747 766
rect 1807 770 1811 771
rect 1807 765 1811 766
rect 1831 770 1835 771
rect 1831 765 1835 766
rect 1919 770 1923 771
rect 1919 765 1923 766
rect 1927 770 1931 771
rect 1927 765 1931 766
rect 2007 770 2011 771
rect 2007 765 2011 766
rect 2039 770 2043 771
rect 2039 765 2043 766
rect 2095 770 2099 771
rect 2095 765 2099 766
rect 2143 770 2147 771
rect 2143 765 2147 766
rect 2183 770 2187 771
rect 2183 765 2187 766
rect 2247 770 2251 771
rect 2247 765 2251 766
rect 2271 770 2275 771
rect 2271 765 2275 766
rect 1806 764 1812 765
rect 1806 760 1807 764
rect 1811 760 1812 764
rect 1806 759 1812 760
rect 1926 764 1932 765
rect 1926 760 1927 764
rect 1931 760 1932 764
rect 1926 759 1932 760
rect 2038 764 2044 765
rect 2038 760 2039 764
rect 2043 760 2044 764
rect 2038 759 2044 760
rect 2142 764 2148 765
rect 2142 760 2143 764
rect 2147 760 2148 764
rect 2142 759 2148 760
rect 2246 764 2252 765
rect 2246 760 2247 764
rect 2251 760 2252 764
rect 2246 759 2252 760
rect 1702 743 1708 744
rect 1702 739 1703 743
rect 1707 739 1708 743
rect 1702 738 1708 739
rect 1722 743 1728 744
rect 1722 739 1723 743
rect 1727 739 1728 743
rect 1722 738 1728 739
rect 1822 743 1828 744
rect 1822 739 1823 743
rect 1827 739 1828 743
rect 1822 738 1828 739
rect 1942 743 1948 744
rect 1942 739 1943 743
rect 1947 739 1948 743
rect 1942 738 1948 739
rect 2054 743 2060 744
rect 2054 739 2055 743
rect 2059 739 2060 743
rect 2054 738 2060 739
rect 2158 743 2164 744
rect 2158 739 2159 743
rect 2163 739 2164 743
rect 2158 738 2164 739
rect 2262 743 2268 744
rect 2262 739 2263 743
rect 2267 739 2268 743
rect 2262 738 2268 739
rect 2270 743 2276 744
rect 2270 739 2271 743
rect 2275 739 2276 743
rect 2270 738 2276 739
rect 1598 727 1604 728
rect 1598 723 1599 727
rect 1603 723 1604 727
rect 1598 722 1604 723
rect 1704 715 1706 738
rect 1824 715 1826 738
rect 1882 727 1888 728
rect 1882 723 1883 727
rect 1887 723 1888 727
rect 1882 722 1888 723
rect 1431 714 1435 715
rect 1431 709 1435 710
rect 1463 714 1467 715
rect 1463 709 1467 710
rect 1535 714 1539 715
rect 1535 709 1539 710
rect 1583 714 1587 715
rect 1583 709 1587 710
rect 1639 714 1643 715
rect 1639 709 1643 710
rect 1703 714 1707 715
rect 1703 709 1707 710
rect 1751 714 1755 715
rect 1751 709 1755 710
rect 1823 714 1827 715
rect 1823 709 1827 710
rect 1863 714 1867 715
rect 1863 709 1867 710
rect 1374 703 1380 704
rect 1374 699 1375 703
rect 1379 699 1380 703
rect 1374 698 1380 699
rect 1432 690 1434 709
rect 1536 690 1538 709
rect 1640 690 1642 709
rect 1752 690 1754 709
rect 1758 703 1764 704
rect 1758 699 1759 703
rect 1763 699 1764 703
rect 1758 698 1764 699
rect 1366 689 1372 690
rect 1326 688 1332 689
rect 1326 684 1327 688
rect 1331 684 1332 688
rect 1366 685 1367 689
rect 1371 685 1372 689
rect 1366 684 1372 685
rect 1430 689 1436 690
rect 1430 685 1431 689
rect 1435 685 1436 689
rect 1430 684 1436 685
rect 1534 689 1540 690
rect 1534 685 1535 689
rect 1539 685 1540 689
rect 1534 684 1540 685
rect 1638 689 1644 690
rect 1638 685 1639 689
rect 1643 685 1644 689
rect 1750 689 1756 690
rect 1638 684 1644 685
rect 1654 687 1660 688
rect 1286 683 1292 684
rect 1326 683 1332 684
rect 1654 683 1655 687
rect 1659 683 1660 687
rect 1750 685 1751 689
rect 1755 685 1756 689
rect 1750 684 1756 685
rect 686 680 692 681
rect 686 676 687 680
rect 691 676 692 680
rect 686 675 692 676
rect 750 680 756 681
rect 750 676 751 680
rect 755 676 756 680
rect 750 675 756 676
rect 822 680 828 681
rect 822 676 823 680
rect 827 676 828 680
rect 822 675 828 676
rect 894 680 900 681
rect 894 676 895 680
rect 899 676 900 680
rect 1286 679 1287 683
rect 1291 679 1292 683
rect 1654 682 1660 683
rect 1286 678 1292 679
rect 894 675 900 676
rect 1288 675 1290 678
rect 655 674 659 675
rect 655 669 659 670
rect 687 674 691 675
rect 687 669 691 670
rect 719 674 723 675
rect 719 669 723 670
rect 751 674 755 675
rect 751 669 755 670
rect 783 674 787 675
rect 783 669 787 670
rect 823 674 827 675
rect 823 669 827 670
rect 847 674 851 675
rect 847 669 851 670
rect 895 674 899 675
rect 895 669 899 670
rect 919 674 923 675
rect 919 669 923 670
rect 1287 674 1291 675
rect 1287 669 1291 670
rect 1326 671 1332 672
rect 654 668 660 669
rect 654 664 655 668
rect 659 664 660 668
rect 654 663 660 664
rect 718 668 724 669
rect 718 664 719 668
rect 723 664 724 668
rect 718 663 724 664
rect 782 668 788 669
rect 782 664 783 668
rect 787 664 788 668
rect 782 663 788 664
rect 846 668 852 669
rect 846 664 847 668
rect 851 664 852 668
rect 846 663 852 664
rect 918 668 924 669
rect 918 664 919 668
rect 923 664 924 668
rect 1288 666 1290 669
rect 1326 667 1327 671
rect 1331 667 1332 671
rect 1326 666 1332 667
rect 1350 668 1356 669
rect 918 663 924 664
rect 1286 665 1292 666
rect 1286 661 1287 665
rect 1291 661 1292 665
rect 1286 660 1292 661
rect 1328 655 1330 666
rect 1350 664 1351 668
rect 1355 664 1356 668
rect 1350 663 1356 664
rect 1414 668 1420 669
rect 1414 664 1415 668
rect 1419 664 1420 668
rect 1414 663 1420 664
rect 1518 668 1524 669
rect 1518 664 1519 668
rect 1523 664 1524 668
rect 1518 663 1524 664
rect 1622 668 1628 669
rect 1622 664 1623 668
rect 1627 664 1628 668
rect 1622 663 1628 664
rect 1352 655 1354 663
rect 1416 655 1418 663
rect 1520 655 1522 663
rect 1624 655 1626 663
rect 1327 654 1331 655
rect 1327 649 1331 650
rect 1351 654 1355 655
rect 1351 649 1355 650
rect 1415 654 1419 655
rect 1415 649 1419 650
rect 1479 654 1483 655
rect 1479 649 1483 650
rect 1519 654 1523 655
rect 1519 649 1523 650
rect 1559 654 1563 655
rect 1559 649 1563 650
rect 1623 654 1627 655
rect 1623 649 1627 650
rect 1647 654 1651 655
rect 1647 649 1651 650
rect 1286 648 1292 649
rect 542 647 548 648
rect 542 643 543 647
rect 547 643 548 647
rect 542 642 548 643
rect 606 647 612 648
rect 606 643 607 647
rect 611 643 612 647
rect 606 642 612 643
rect 630 647 636 648
rect 630 643 631 647
rect 635 643 636 647
rect 630 642 636 643
rect 670 647 676 648
rect 670 643 671 647
rect 675 643 676 647
rect 670 642 676 643
rect 734 647 740 648
rect 734 643 735 647
rect 739 643 740 647
rect 734 642 740 643
rect 750 647 756 648
rect 750 643 751 647
rect 755 643 756 647
rect 750 642 756 643
rect 798 647 804 648
rect 798 643 799 647
rect 803 643 804 647
rect 798 642 804 643
rect 862 647 868 648
rect 862 643 863 647
rect 867 643 868 647
rect 862 642 868 643
rect 934 647 940 648
rect 934 643 935 647
rect 939 643 940 647
rect 934 642 940 643
rect 942 647 948 648
rect 942 643 943 647
rect 947 643 948 647
rect 1286 644 1287 648
rect 1291 644 1292 648
rect 1328 646 1330 649
rect 1478 648 1484 649
rect 1286 643 1292 644
rect 1326 645 1332 646
rect 942 642 948 643
rect 534 631 540 632
rect 534 627 535 631
rect 539 627 540 631
rect 534 626 540 627
rect 544 619 546 642
rect 608 619 610 642
rect 672 619 674 642
rect 736 619 738 642
rect 752 628 754 642
rect 750 627 756 628
rect 750 623 751 627
rect 755 623 756 627
rect 750 622 756 623
rect 800 619 802 642
rect 864 619 866 642
rect 870 631 876 632
rect 870 627 871 631
rect 875 627 876 631
rect 870 626 876 627
rect 503 618 507 619
rect 503 613 507 614
rect 543 618 547 619
rect 543 613 547 614
rect 599 618 603 619
rect 599 613 603 614
rect 607 618 611 619
rect 607 613 611 614
rect 671 618 675 619
rect 671 613 675 614
rect 687 618 691 619
rect 687 613 691 614
rect 735 618 739 619
rect 735 613 739 614
rect 767 618 771 619
rect 767 613 771 614
rect 799 618 803 619
rect 799 613 803 614
rect 847 618 851 619
rect 847 613 851 614
rect 863 618 867 619
rect 863 613 867 614
rect 494 607 500 608
rect 494 603 495 607
rect 499 603 500 607
rect 494 602 500 603
rect 504 594 506 613
rect 600 594 602 613
rect 688 594 690 613
rect 768 594 770 613
rect 848 594 850 613
rect 502 593 508 594
rect 426 591 432 592
rect 426 587 427 591
rect 431 587 432 591
rect 502 589 503 593
rect 507 589 508 593
rect 502 588 508 589
rect 598 593 604 594
rect 598 589 599 593
rect 603 589 604 593
rect 686 593 692 594
rect 598 588 604 589
rect 622 591 628 592
rect 426 586 432 587
rect 622 587 623 591
rect 627 587 628 591
rect 686 589 687 593
rect 691 589 692 593
rect 686 588 692 589
rect 766 593 772 594
rect 766 589 767 593
rect 771 589 772 593
rect 766 588 772 589
rect 846 593 852 594
rect 846 589 847 593
rect 851 589 852 593
rect 872 592 874 626
rect 936 619 938 642
rect 944 624 946 642
rect 942 623 948 624
rect 942 619 943 623
rect 947 619 948 623
rect 1288 619 1290 643
rect 1326 641 1327 645
rect 1331 641 1332 645
rect 1478 644 1479 648
rect 1483 644 1484 648
rect 1478 643 1484 644
rect 1558 648 1564 649
rect 1558 644 1559 648
rect 1563 644 1564 648
rect 1558 643 1564 644
rect 1646 648 1652 649
rect 1646 644 1647 648
rect 1651 644 1652 648
rect 1646 643 1652 644
rect 1326 640 1332 641
rect 1326 628 1332 629
rect 1326 624 1327 628
rect 1331 624 1332 628
rect 1326 623 1332 624
rect 1494 627 1500 628
rect 1494 623 1495 627
rect 1499 623 1500 627
rect 927 618 931 619
rect 927 613 931 614
rect 935 618 939 619
rect 942 618 948 619
rect 1007 618 1011 619
rect 935 613 939 614
rect 1007 613 1011 614
rect 1087 618 1091 619
rect 1287 618 1291 619
rect 1087 613 1091 614
rect 1106 615 1112 616
rect 928 594 930 613
rect 1008 594 1010 613
rect 1014 607 1020 608
rect 1014 603 1015 607
rect 1019 603 1020 607
rect 1014 602 1020 603
rect 926 593 932 594
rect 846 588 852 589
rect 870 591 876 592
rect 622 586 628 587
rect 870 587 871 591
rect 875 587 876 591
rect 926 589 927 593
rect 931 589 932 593
rect 926 588 932 589
rect 1006 593 1012 594
rect 1006 589 1007 593
rect 1011 589 1012 593
rect 1006 588 1012 589
rect 870 586 876 587
rect 486 572 492 573
rect 486 568 487 572
rect 491 568 492 572
rect 486 567 492 568
rect 582 572 588 573
rect 582 568 583 572
rect 587 568 588 572
rect 582 567 588 568
rect 488 563 490 567
rect 584 563 586 567
rect 487 562 491 563
rect 487 557 491 558
rect 583 562 587 563
rect 583 557 587 558
rect 591 562 595 563
rect 591 557 595 558
rect 486 556 492 557
rect 486 552 487 556
rect 491 552 492 556
rect 486 551 492 552
rect 590 556 596 557
rect 590 552 591 556
rect 595 552 596 556
rect 590 551 596 552
rect 238 535 244 536
rect 238 531 239 535
rect 243 531 244 535
rect 238 530 244 531
rect 286 535 292 536
rect 286 531 287 535
rect 291 531 292 535
rect 286 530 292 531
rect 390 535 396 536
rect 390 531 391 535
rect 395 531 396 535
rect 390 530 396 531
rect 414 535 420 536
rect 414 531 415 535
rect 419 531 420 535
rect 414 530 420 531
rect 502 535 508 536
rect 502 531 503 535
rect 507 531 508 535
rect 502 530 508 531
rect 606 535 612 536
rect 606 531 607 535
rect 611 531 612 535
rect 606 530 612 531
rect 214 519 220 520
rect 214 515 215 519
rect 219 515 220 519
rect 214 514 220 515
rect 111 506 115 507
rect 111 501 115 502
rect 151 506 155 507
rect 151 501 155 502
rect 191 506 195 507
rect 191 501 195 502
rect 112 481 114 501
rect 152 482 154 501
rect 240 496 242 530
rect 288 507 290 530
rect 392 507 394 530
rect 494 515 500 516
rect 494 511 495 515
rect 499 511 500 515
rect 494 510 500 511
rect 247 506 251 507
rect 247 501 251 502
rect 287 506 291 507
rect 287 501 291 502
rect 367 506 371 507
rect 367 501 371 502
rect 391 506 395 507
rect 391 501 395 502
rect 487 506 491 507
rect 487 501 491 502
rect 238 495 244 496
rect 238 491 239 495
rect 243 491 244 495
rect 238 490 244 491
rect 248 482 250 501
rect 342 495 348 496
rect 342 491 343 495
rect 347 491 348 495
rect 342 490 348 491
rect 150 481 156 482
rect 110 480 116 481
rect 110 476 111 480
rect 115 476 116 480
rect 150 477 151 481
rect 155 477 156 481
rect 246 481 252 482
rect 150 476 156 477
rect 158 479 164 480
rect 110 475 116 476
rect 158 475 159 479
rect 163 475 164 479
rect 246 477 247 481
rect 251 477 252 481
rect 246 476 252 477
rect 158 474 164 475
rect 110 463 116 464
rect 110 459 111 463
rect 115 459 116 463
rect 110 458 116 459
rect 134 460 140 461
rect 112 451 114 458
rect 134 456 135 460
rect 139 456 140 460
rect 134 455 140 456
rect 136 451 138 455
rect 111 450 115 451
rect 111 445 115 446
rect 135 450 139 451
rect 135 445 139 446
rect 112 442 114 445
rect 134 444 140 445
rect 110 441 116 442
rect 110 437 111 441
rect 115 437 116 441
rect 134 440 135 444
rect 139 440 140 444
rect 134 439 140 440
rect 110 436 116 437
rect 110 424 116 425
rect 110 420 111 424
rect 115 420 116 424
rect 110 419 116 420
rect 150 423 156 424
rect 150 419 151 423
rect 155 419 156 423
rect 112 391 114 419
rect 150 418 156 419
rect 152 391 154 418
rect 160 408 162 474
rect 230 460 236 461
rect 230 456 231 460
rect 235 456 236 460
rect 230 455 236 456
rect 232 451 234 455
rect 191 450 195 451
rect 191 445 195 446
rect 231 450 235 451
rect 231 445 235 446
rect 247 450 251 451
rect 247 445 251 446
rect 303 450 307 451
rect 303 445 307 446
rect 190 444 196 445
rect 190 440 191 444
rect 195 440 196 444
rect 190 439 196 440
rect 246 444 252 445
rect 246 440 247 444
rect 251 440 252 444
rect 246 439 252 440
rect 302 444 308 445
rect 302 440 303 444
rect 307 440 308 444
rect 302 439 308 440
rect 344 424 346 490
rect 368 482 370 501
rect 488 482 490 501
rect 366 481 372 482
rect 366 477 367 481
rect 371 477 372 481
rect 366 476 372 477
rect 486 481 492 482
rect 486 477 487 481
rect 491 477 492 481
rect 496 480 498 510
rect 504 507 506 530
rect 608 507 610 530
rect 624 516 626 586
rect 670 572 676 573
rect 670 568 671 572
rect 675 568 676 572
rect 670 567 676 568
rect 750 572 756 573
rect 750 568 751 572
rect 755 568 756 572
rect 750 567 756 568
rect 830 572 836 573
rect 830 568 831 572
rect 835 568 836 572
rect 830 567 836 568
rect 910 572 916 573
rect 910 568 911 572
rect 915 568 916 572
rect 910 567 916 568
rect 990 572 996 573
rect 990 568 991 572
rect 995 568 996 572
rect 990 567 996 568
rect 672 563 674 567
rect 752 563 754 567
rect 832 563 834 567
rect 912 563 914 567
rect 992 563 994 567
rect 671 562 675 563
rect 671 557 675 558
rect 695 562 699 563
rect 695 557 699 558
rect 751 562 755 563
rect 751 557 755 558
rect 791 562 795 563
rect 791 557 795 558
rect 831 562 835 563
rect 831 557 835 558
rect 879 562 883 563
rect 879 557 883 558
rect 911 562 915 563
rect 911 557 915 558
rect 967 562 971 563
rect 967 557 971 558
rect 991 562 995 563
rect 991 557 995 558
rect 694 556 700 557
rect 694 552 695 556
rect 699 552 700 556
rect 694 551 700 552
rect 790 556 796 557
rect 790 552 791 556
rect 795 552 796 556
rect 790 551 796 552
rect 878 556 884 557
rect 878 552 879 556
rect 883 552 884 556
rect 878 551 884 552
rect 966 556 972 557
rect 966 552 967 556
rect 971 552 972 556
rect 966 551 972 552
rect 1016 536 1018 602
rect 1088 594 1090 613
rect 1106 611 1107 615
rect 1111 611 1112 615
rect 1287 613 1291 614
rect 1106 610 1112 611
rect 1086 593 1092 594
rect 1086 589 1087 593
rect 1091 589 1092 593
rect 1108 592 1110 610
rect 1288 593 1290 613
rect 1328 599 1330 623
rect 1494 622 1500 623
rect 1574 627 1580 628
rect 1574 623 1575 627
rect 1579 623 1580 627
rect 1574 622 1580 623
rect 1496 599 1498 622
rect 1576 599 1578 622
rect 1656 608 1658 682
rect 1734 668 1740 669
rect 1734 664 1735 668
rect 1739 664 1740 668
rect 1734 663 1740 664
rect 1736 655 1738 663
rect 1735 654 1739 655
rect 1735 649 1739 650
rect 1734 648 1740 649
rect 1734 644 1735 648
rect 1739 644 1740 648
rect 1734 643 1740 644
rect 1760 628 1762 698
rect 1864 690 1866 709
rect 1862 689 1868 690
rect 1862 685 1863 689
rect 1867 685 1868 689
rect 1884 688 1886 722
rect 1944 715 1946 738
rect 1975 724 1979 725
rect 1975 719 1979 720
rect 1943 714 1947 715
rect 1943 709 1947 710
rect 1967 714 1971 715
rect 1967 709 1971 710
rect 1968 690 1970 709
rect 1976 704 1978 719
rect 2056 715 2058 738
rect 2160 715 2162 738
rect 2264 715 2266 738
rect 2272 725 2274 738
rect 2271 724 2275 725
rect 2296 724 2298 794
rect 2366 780 2372 781
rect 2366 776 2367 780
rect 2371 776 2372 780
rect 2366 775 2372 776
rect 2368 771 2370 775
rect 2351 770 2355 771
rect 2351 765 2355 766
rect 2367 770 2371 771
rect 2367 765 2371 766
rect 2350 764 2356 765
rect 2350 760 2351 764
rect 2355 760 2356 764
rect 2350 759 2356 760
rect 2392 744 2394 810
rect 2408 800 2410 930
rect 2422 900 2428 901
rect 2422 896 2423 900
rect 2427 896 2428 900
rect 2422 895 2428 896
rect 2424 887 2426 895
rect 2423 886 2427 887
rect 2423 881 2427 882
rect 2432 844 2434 982
rect 2446 971 2452 972
rect 2446 967 2447 971
rect 2451 967 2452 971
rect 2446 966 2452 967
rect 2439 946 2443 947
rect 2439 941 2443 942
rect 2440 922 2442 941
rect 2438 921 2444 922
rect 2438 917 2439 921
rect 2443 917 2444 921
rect 2448 920 2450 966
rect 2456 947 2458 982
rect 2464 972 2466 1042
rect 2480 988 2482 1174
rect 2504 1165 2506 1185
rect 2502 1164 2508 1165
rect 2502 1160 2503 1164
rect 2507 1160 2508 1164
rect 2502 1159 2508 1160
rect 2502 1147 2508 1148
rect 2502 1143 2503 1147
rect 2507 1143 2508 1147
rect 2502 1142 2508 1143
rect 2504 1135 2506 1142
rect 2503 1134 2507 1135
rect 2503 1129 2507 1130
rect 2504 1126 2506 1129
rect 2502 1125 2508 1126
rect 2502 1121 2503 1125
rect 2507 1121 2508 1125
rect 2502 1120 2508 1121
rect 2502 1108 2508 1109
rect 2502 1104 2503 1108
rect 2507 1104 2508 1108
rect 2502 1103 2508 1104
rect 2504 1075 2506 1103
rect 2503 1074 2507 1075
rect 2503 1069 2507 1070
rect 2504 1049 2506 1069
rect 2502 1048 2508 1049
rect 2502 1044 2503 1048
rect 2507 1044 2508 1048
rect 2502 1043 2508 1044
rect 2502 1031 2508 1032
rect 2502 1027 2503 1031
rect 2507 1027 2508 1031
rect 2502 1026 2508 1027
rect 2504 1015 2506 1026
rect 2503 1014 2507 1015
rect 2503 1009 2507 1010
rect 2504 1006 2506 1009
rect 2502 1005 2508 1006
rect 2502 1001 2503 1005
rect 2507 1001 2508 1005
rect 2502 1000 2508 1001
rect 2502 988 2508 989
rect 2478 987 2484 988
rect 2478 983 2479 987
rect 2483 983 2484 987
rect 2502 984 2503 988
rect 2507 984 2508 988
rect 2502 983 2508 984
rect 2478 982 2484 983
rect 2462 971 2468 972
rect 2462 967 2463 971
rect 2467 967 2468 971
rect 2462 966 2468 967
rect 2504 947 2506 983
rect 2455 946 2459 947
rect 2455 941 2459 942
rect 2503 946 2507 947
rect 2503 941 2507 942
rect 2504 921 2506 941
rect 2502 920 2508 921
rect 2438 916 2444 917
rect 2446 919 2452 920
rect 2446 915 2447 919
rect 2451 915 2452 919
rect 2502 916 2503 920
rect 2507 916 2508 920
rect 2502 915 2508 916
rect 2446 914 2452 915
rect 2502 903 2508 904
rect 2502 899 2503 903
rect 2507 899 2508 903
rect 2502 898 2508 899
rect 2504 887 2506 898
rect 2439 886 2443 887
rect 2439 881 2443 882
rect 2503 886 2507 887
rect 2503 881 2507 882
rect 2438 880 2444 881
rect 2438 876 2439 880
rect 2443 876 2444 880
rect 2504 878 2506 881
rect 2438 875 2444 876
rect 2502 877 2508 878
rect 2502 873 2503 877
rect 2507 873 2508 877
rect 2502 872 2508 873
rect 2502 860 2508 861
rect 2454 859 2460 860
rect 2454 855 2455 859
rect 2459 855 2460 859
rect 2454 854 2460 855
rect 2462 859 2468 860
rect 2462 855 2463 859
rect 2467 855 2468 859
rect 2502 856 2503 860
rect 2507 856 2508 860
rect 2502 855 2508 856
rect 2462 854 2468 855
rect 2430 843 2436 844
rect 2430 839 2431 843
rect 2435 839 2436 843
rect 2430 838 2436 839
rect 2456 827 2458 854
rect 2455 826 2459 827
rect 2455 821 2459 822
rect 2456 802 2458 821
rect 2464 816 2466 854
rect 2504 827 2506 855
rect 2503 826 2507 827
rect 2503 821 2507 822
rect 2462 815 2468 816
rect 2462 811 2463 815
rect 2467 811 2468 815
rect 2462 810 2468 811
rect 2454 801 2460 802
rect 2504 801 2506 821
rect 2406 799 2412 800
rect 2406 795 2407 799
rect 2411 795 2412 799
rect 2454 797 2455 801
rect 2459 797 2460 801
rect 2502 800 2508 801
rect 2454 796 2460 797
rect 2470 799 2476 800
rect 2406 794 2412 795
rect 2470 795 2471 799
rect 2475 795 2476 799
rect 2502 796 2503 800
rect 2507 796 2508 800
rect 2502 795 2508 796
rect 2470 794 2476 795
rect 2438 780 2444 781
rect 2438 776 2439 780
rect 2443 776 2444 780
rect 2438 775 2444 776
rect 2440 771 2442 775
rect 2439 770 2443 771
rect 2439 765 2443 766
rect 2438 764 2444 765
rect 2438 760 2439 764
rect 2443 760 2444 764
rect 2438 759 2444 760
rect 2366 743 2372 744
rect 2366 739 2367 743
rect 2371 739 2372 743
rect 2366 738 2372 739
rect 2390 743 2396 744
rect 2390 739 2391 743
rect 2395 739 2396 743
rect 2390 738 2396 739
rect 2454 743 2460 744
rect 2454 739 2455 743
rect 2459 739 2460 743
rect 2454 738 2460 739
rect 2462 743 2468 744
rect 2462 739 2463 743
rect 2467 739 2468 743
rect 2462 738 2468 739
rect 2271 719 2275 720
rect 2294 723 2300 724
rect 2294 719 2295 723
rect 2299 719 2300 723
rect 2294 718 2300 719
rect 2368 715 2370 738
rect 2410 727 2416 728
rect 2410 723 2411 727
rect 2415 723 2416 727
rect 2410 722 2416 723
rect 2055 714 2059 715
rect 2055 709 2059 710
rect 2063 714 2067 715
rect 2063 709 2067 710
rect 2151 714 2155 715
rect 2151 709 2155 710
rect 2159 714 2163 715
rect 2159 709 2163 710
rect 2231 714 2235 715
rect 2231 709 2235 710
rect 2263 714 2267 715
rect 2263 709 2267 710
rect 2311 714 2315 715
rect 2311 709 2315 710
rect 2367 714 2371 715
rect 2367 709 2371 710
rect 2391 714 2395 715
rect 2391 709 2395 710
rect 1974 703 1980 704
rect 1974 699 1975 703
rect 1979 699 1980 703
rect 1974 698 1980 699
rect 2064 690 2066 709
rect 2152 690 2154 709
rect 2232 690 2234 709
rect 2274 703 2280 704
rect 2274 699 2275 703
rect 2279 699 2280 703
rect 2274 698 2280 699
rect 1966 689 1972 690
rect 1862 684 1868 685
rect 1882 687 1888 688
rect 1882 683 1883 687
rect 1887 683 1888 687
rect 1966 685 1967 689
rect 1971 685 1972 689
rect 1966 684 1972 685
rect 2062 689 2068 690
rect 2062 685 2063 689
rect 2067 685 2068 689
rect 2062 684 2068 685
rect 2150 689 2156 690
rect 2150 685 2151 689
rect 2155 685 2156 689
rect 2150 684 2156 685
rect 2230 689 2236 690
rect 2230 685 2231 689
rect 2235 685 2236 689
rect 2230 684 2236 685
rect 2246 687 2252 688
rect 1882 682 1888 683
rect 2246 683 2247 687
rect 2251 683 2252 687
rect 2246 682 2252 683
rect 1846 668 1852 669
rect 1846 664 1847 668
rect 1851 664 1852 668
rect 1846 663 1852 664
rect 1950 668 1956 669
rect 1950 664 1951 668
rect 1955 664 1956 668
rect 1950 663 1956 664
rect 2046 668 2052 669
rect 2046 664 2047 668
rect 2051 664 2052 668
rect 2046 663 2052 664
rect 2134 668 2140 669
rect 2134 664 2135 668
rect 2139 664 2140 668
rect 2134 663 2140 664
rect 2214 668 2220 669
rect 2214 664 2215 668
rect 2219 664 2220 668
rect 2214 663 2220 664
rect 1848 655 1850 663
rect 1952 655 1954 663
rect 2048 655 2050 663
rect 2136 655 2138 663
rect 2216 655 2218 663
rect 1831 654 1835 655
rect 1831 649 1835 650
rect 1847 654 1851 655
rect 1847 649 1851 650
rect 1919 654 1923 655
rect 1919 649 1923 650
rect 1951 654 1955 655
rect 1951 649 1955 650
rect 2007 654 2011 655
rect 2007 649 2011 650
rect 2047 654 2051 655
rect 2047 649 2051 650
rect 2087 654 2091 655
rect 2087 649 2091 650
rect 2135 654 2139 655
rect 2135 649 2139 650
rect 2167 654 2171 655
rect 2167 649 2171 650
rect 2215 654 2219 655
rect 2215 649 2219 650
rect 2239 654 2243 655
rect 2239 649 2243 650
rect 1830 648 1836 649
rect 1830 644 1831 648
rect 1835 644 1836 648
rect 1830 643 1836 644
rect 1918 648 1924 649
rect 1918 644 1919 648
rect 1923 644 1924 648
rect 1918 643 1924 644
rect 2006 648 2012 649
rect 2006 644 2007 648
rect 2011 644 2012 648
rect 2006 643 2012 644
rect 2086 648 2092 649
rect 2086 644 2087 648
rect 2091 644 2092 648
rect 2086 643 2092 644
rect 2166 648 2172 649
rect 2166 644 2167 648
rect 2171 644 2172 648
rect 2166 643 2172 644
rect 2238 648 2244 649
rect 2238 644 2239 648
rect 2243 644 2244 648
rect 2238 643 2244 644
rect 1662 627 1668 628
rect 1662 623 1663 627
rect 1667 623 1668 627
rect 1662 622 1668 623
rect 1678 627 1684 628
rect 1678 623 1679 627
rect 1683 623 1684 627
rect 1678 622 1684 623
rect 1750 627 1756 628
rect 1750 623 1751 627
rect 1755 623 1756 627
rect 1750 622 1756 623
rect 1758 627 1764 628
rect 1758 623 1759 627
rect 1763 623 1764 627
rect 1758 622 1764 623
rect 1846 627 1852 628
rect 1846 623 1847 627
rect 1851 623 1852 627
rect 1846 622 1852 623
rect 1862 627 1868 628
rect 1862 623 1863 627
rect 1867 623 1868 627
rect 1862 622 1868 623
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 1934 622 1940 623
rect 2022 627 2028 628
rect 2022 623 2023 627
rect 2027 623 2028 627
rect 2022 622 2028 623
rect 2102 627 2108 628
rect 2102 623 2103 627
rect 2107 623 2108 627
rect 2102 622 2108 623
rect 2174 627 2180 628
rect 2174 623 2175 627
rect 2179 623 2180 627
rect 2174 622 2180 623
rect 2182 627 2188 628
rect 2182 623 2183 627
rect 2187 623 2188 627
rect 2182 622 2188 623
rect 1654 607 1660 608
rect 1654 603 1655 607
rect 1659 603 1660 607
rect 1654 602 1660 603
rect 1664 599 1666 622
rect 1327 598 1331 599
rect 1327 593 1331 594
rect 1455 598 1459 599
rect 1455 593 1459 594
rect 1495 598 1499 599
rect 1495 593 1499 594
rect 1559 598 1563 599
rect 1559 593 1563 594
rect 1575 598 1579 599
rect 1575 593 1579 594
rect 1663 598 1667 599
rect 1663 593 1667 594
rect 1671 598 1675 599
rect 1671 593 1675 594
rect 1286 592 1292 593
rect 1086 588 1092 589
rect 1106 591 1112 592
rect 1106 587 1107 591
rect 1111 587 1112 591
rect 1286 588 1287 592
rect 1291 588 1292 592
rect 1286 587 1292 588
rect 1106 586 1112 587
rect 1286 575 1292 576
rect 1070 572 1076 573
rect 1070 568 1071 572
rect 1075 568 1076 572
rect 1286 571 1287 575
rect 1291 571 1292 575
rect 1328 573 1330 593
rect 1456 574 1458 593
rect 1560 574 1562 593
rect 1672 574 1674 593
rect 1680 588 1682 622
rect 1752 599 1754 622
rect 1848 599 1850 622
rect 1864 608 1866 622
rect 1902 611 1908 612
rect 1862 607 1868 608
rect 1862 603 1863 607
rect 1867 603 1868 607
rect 1902 607 1903 611
rect 1907 607 1908 611
rect 1902 606 1908 607
rect 1862 602 1868 603
rect 1751 598 1755 599
rect 1751 593 1755 594
rect 1775 598 1779 599
rect 1775 593 1779 594
rect 1847 598 1851 599
rect 1847 593 1851 594
rect 1879 598 1883 599
rect 1879 593 1883 594
rect 1678 587 1684 588
rect 1678 583 1679 587
rect 1683 583 1684 587
rect 1678 582 1684 583
rect 1776 574 1778 593
rect 1834 587 1840 588
rect 1834 583 1835 587
rect 1839 583 1840 587
rect 1834 582 1840 583
rect 1454 573 1460 574
rect 1286 570 1292 571
rect 1326 572 1332 573
rect 1070 567 1076 568
rect 1072 563 1074 567
rect 1288 563 1290 570
rect 1326 568 1327 572
rect 1331 568 1332 572
rect 1454 569 1455 573
rect 1459 569 1460 573
rect 1558 573 1564 574
rect 1454 568 1460 569
rect 1470 571 1476 572
rect 1326 567 1332 568
rect 1470 567 1471 571
rect 1475 567 1476 571
rect 1558 569 1559 573
rect 1563 569 1564 573
rect 1558 568 1564 569
rect 1670 573 1676 574
rect 1670 569 1671 573
rect 1675 569 1676 573
rect 1670 568 1676 569
rect 1774 573 1780 574
rect 1774 569 1775 573
rect 1779 569 1780 573
rect 1774 568 1780 569
rect 1470 566 1476 567
rect 1055 562 1059 563
rect 1055 557 1059 558
rect 1071 562 1075 563
rect 1071 557 1075 558
rect 1151 562 1155 563
rect 1151 557 1155 558
rect 1287 562 1291 563
rect 1287 557 1291 558
rect 1054 556 1060 557
rect 1054 552 1055 556
rect 1059 552 1060 556
rect 1054 551 1060 552
rect 1150 556 1156 557
rect 1150 552 1151 556
rect 1155 552 1156 556
rect 1288 554 1290 557
rect 1326 555 1332 556
rect 1150 551 1156 552
rect 1286 553 1292 554
rect 1286 549 1287 553
rect 1291 549 1292 553
rect 1326 551 1327 555
rect 1331 551 1332 555
rect 1326 550 1332 551
rect 1438 552 1444 553
rect 1286 548 1292 549
rect 1328 543 1330 550
rect 1438 548 1439 552
rect 1443 548 1444 552
rect 1438 547 1444 548
rect 1440 543 1442 547
rect 1327 542 1331 543
rect 1327 537 1331 538
rect 1367 542 1371 543
rect 1367 537 1371 538
rect 1439 542 1443 543
rect 1439 537 1443 538
rect 1447 542 1451 543
rect 1447 537 1451 538
rect 1286 536 1292 537
rect 710 535 716 536
rect 710 531 711 535
rect 715 531 716 535
rect 710 530 716 531
rect 742 535 748 536
rect 742 531 743 535
rect 747 531 748 535
rect 742 530 748 531
rect 806 535 812 536
rect 806 531 807 535
rect 811 531 812 535
rect 806 530 812 531
rect 894 535 900 536
rect 894 531 895 535
rect 899 531 900 535
rect 894 530 900 531
rect 982 535 988 536
rect 982 531 983 535
rect 987 531 988 535
rect 982 530 988 531
rect 1014 535 1020 536
rect 1014 531 1015 535
rect 1019 531 1020 535
rect 1014 530 1020 531
rect 1070 535 1076 536
rect 1070 531 1071 535
rect 1075 531 1076 535
rect 1070 530 1076 531
rect 1166 535 1172 536
rect 1166 531 1167 535
rect 1171 531 1172 535
rect 1166 530 1172 531
rect 1174 535 1180 536
rect 1174 531 1175 535
rect 1179 531 1180 535
rect 1286 532 1287 536
rect 1291 532 1292 536
rect 1328 534 1330 537
rect 1366 536 1372 537
rect 1286 531 1292 532
rect 1326 533 1332 534
rect 1174 530 1180 531
rect 622 515 628 516
rect 622 511 623 515
rect 627 511 628 515
rect 622 510 628 511
rect 712 507 714 530
rect 503 506 507 507
rect 503 501 507 502
rect 607 506 611 507
rect 607 501 611 502
rect 615 506 619 507
rect 615 501 619 502
rect 711 506 715 507
rect 711 501 715 502
rect 735 506 739 507
rect 735 501 739 502
rect 616 482 618 501
rect 736 482 738 501
rect 744 496 746 530
rect 808 507 810 530
rect 896 507 898 530
rect 984 507 986 530
rect 1072 507 1074 530
rect 1078 519 1084 520
rect 1078 515 1079 519
rect 1083 515 1084 519
rect 1078 514 1084 515
rect 807 506 811 507
rect 807 501 811 502
rect 847 506 851 507
rect 847 501 851 502
rect 895 506 899 507
rect 895 501 899 502
rect 951 506 955 507
rect 951 501 955 502
rect 983 506 987 507
rect 983 501 987 502
rect 1055 506 1059 507
rect 1055 501 1059 502
rect 1071 506 1075 507
rect 1071 501 1075 502
rect 742 495 748 496
rect 742 491 743 495
rect 747 491 748 495
rect 742 490 748 491
rect 848 482 850 501
rect 952 482 954 501
rect 1056 482 1058 501
rect 614 481 620 482
rect 486 476 492 477
rect 494 479 500 480
rect 494 475 495 479
rect 499 475 500 479
rect 614 477 615 481
rect 619 477 620 481
rect 734 481 740 482
rect 614 476 620 477
rect 622 479 628 480
rect 494 474 500 475
rect 622 475 623 479
rect 627 475 628 479
rect 734 477 735 481
rect 739 477 740 481
rect 734 476 740 477
rect 846 481 852 482
rect 846 477 847 481
rect 851 477 852 481
rect 846 476 852 477
rect 950 481 956 482
rect 950 477 951 481
rect 955 477 956 481
rect 950 476 956 477
rect 1054 481 1060 482
rect 1054 477 1055 481
rect 1059 477 1060 481
rect 1080 480 1082 514
rect 1168 507 1170 530
rect 1176 512 1178 530
rect 1174 511 1180 512
rect 1174 507 1175 511
rect 1179 507 1180 511
rect 1288 507 1290 531
rect 1326 529 1327 533
rect 1331 529 1332 533
rect 1366 532 1367 536
rect 1371 532 1372 536
rect 1366 531 1372 532
rect 1446 536 1452 537
rect 1446 532 1447 536
rect 1451 532 1452 536
rect 1446 531 1452 532
rect 1326 528 1332 529
rect 1326 516 1332 517
rect 1326 512 1327 516
rect 1331 512 1332 516
rect 1326 511 1332 512
rect 1382 515 1388 516
rect 1382 511 1383 515
rect 1387 511 1388 515
rect 1159 506 1163 507
rect 1159 501 1163 502
rect 1167 506 1171 507
rect 1174 506 1180 507
rect 1239 506 1243 507
rect 1167 501 1171 502
rect 1178 503 1184 504
rect 1160 482 1162 501
rect 1178 499 1179 503
rect 1183 499 1184 503
rect 1239 501 1243 502
rect 1287 506 1291 507
rect 1287 501 1291 502
rect 1178 498 1184 499
rect 1158 481 1164 482
rect 1054 476 1060 477
rect 1078 479 1084 480
rect 622 474 628 475
rect 1078 475 1079 479
rect 1083 475 1084 479
rect 1158 477 1159 481
rect 1163 477 1164 481
rect 1180 480 1182 498
rect 1240 482 1242 501
rect 1258 495 1264 496
rect 1258 491 1259 495
rect 1263 491 1264 495
rect 1258 490 1264 491
rect 1238 481 1244 482
rect 1158 476 1164 477
rect 1178 479 1184 480
rect 1078 474 1084 475
rect 1178 475 1179 479
rect 1183 475 1184 479
rect 1238 477 1239 481
rect 1243 477 1244 481
rect 1238 476 1244 477
rect 1178 474 1184 475
rect 350 460 356 461
rect 350 456 351 460
rect 355 456 356 460
rect 350 455 356 456
rect 470 460 476 461
rect 470 456 471 460
rect 475 456 476 460
rect 470 455 476 456
rect 598 460 604 461
rect 598 456 599 460
rect 603 456 604 460
rect 598 455 604 456
rect 352 451 354 455
rect 472 451 474 455
rect 600 451 602 455
rect 351 450 355 451
rect 351 445 355 446
rect 383 450 387 451
rect 383 445 387 446
rect 471 450 475 451
rect 471 445 475 446
rect 567 450 571 451
rect 567 445 571 446
rect 599 450 603 451
rect 599 445 603 446
rect 382 444 388 445
rect 382 440 383 444
rect 387 440 388 444
rect 382 439 388 440
rect 470 444 476 445
rect 470 440 471 444
rect 475 440 476 444
rect 470 439 476 440
rect 566 444 572 445
rect 566 440 567 444
rect 571 440 572 444
rect 566 439 572 440
rect 206 423 212 424
rect 206 419 207 423
rect 211 419 212 423
rect 206 418 212 419
rect 214 423 220 424
rect 214 419 215 423
rect 219 419 220 423
rect 214 418 220 419
rect 262 423 268 424
rect 262 419 263 423
rect 267 419 268 423
rect 262 418 268 419
rect 318 423 324 424
rect 318 419 319 423
rect 323 419 324 423
rect 318 418 324 419
rect 342 423 348 424
rect 342 419 343 423
rect 347 419 348 423
rect 342 418 348 419
rect 398 423 404 424
rect 398 419 399 423
rect 403 419 404 423
rect 398 418 404 419
rect 414 423 420 424
rect 414 419 415 423
rect 419 419 420 423
rect 414 418 420 419
rect 486 423 492 424
rect 486 419 487 423
rect 491 419 492 423
rect 486 418 492 419
rect 582 423 588 424
rect 582 419 583 423
rect 587 419 588 423
rect 582 418 588 419
rect 158 407 164 408
rect 158 403 159 407
rect 163 403 164 407
rect 158 402 164 403
rect 208 391 210 418
rect 111 390 115 391
rect 111 385 115 386
rect 151 390 155 391
rect 151 385 155 386
rect 207 390 211 391
rect 207 385 211 386
rect 112 365 114 385
rect 152 366 154 385
rect 208 366 210 385
rect 216 380 218 418
rect 264 391 266 418
rect 320 391 322 418
rect 400 391 402 418
rect 416 404 418 418
rect 414 403 420 404
rect 414 399 415 403
rect 419 399 420 403
rect 414 398 420 399
rect 488 391 490 418
rect 530 407 536 408
rect 530 403 531 407
rect 535 403 536 407
rect 530 402 536 403
rect 263 390 267 391
rect 263 385 267 386
rect 279 390 283 391
rect 319 390 323 391
rect 279 385 283 386
rect 298 387 304 388
rect 214 379 220 380
rect 214 375 215 379
rect 219 375 220 379
rect 214 374 220 375
rect 280 366 282 385
rect 298 383 299 387
rect 303 383 304 387
rect 319 385 323 386
rect 359 390 363 391
rect 359 385 363 386
rect 399 390 403 391
rect 399 385 403 386
rect 431 390 435 391
rect 487 390 491 391
rect 431 385 435 386
rect 478 387 484 388
rect 298 382 304 383
rect 150 365 156 366
rect 110 364 116 365
rect 110 360 111 364
rect 115 360 116 364
rect 150 361 151 365
rect 155 361 156 365
rect 206 365 212 366
rect 150 360 156 361
rect 158 363 164 364
rect 110 359 116 360
rect 158 359 159 363
rect 163 359 164 363
rect 206 361 207 365
rect 211 361 212 365
rect 206 360 212 361
rect 278 365 284 366
rect 278 361 279 365
rect 283 361 284 365
rect 300 364 302 382
rect 360 366 362 385
rect 432 366 434 385
rect 478 383 479 387
rect 483 383 484 387
rect 487 385 491 386
rect 511 390 515 391
rect 511 385 515 386
rect 478 382 484 383
rect 358 365 364 366
rect 278 360 284 361
rect 298 363 304 364
rect 158 358 164 359
rect 298 359 299 363
rect 303 359 304 363
rect 358 361 359 365
rect 363 361 364 365
rect 358 360 364 361
rect 430 365 436 366
rect 430 361 431 365
rect 435 361 436 365
rect 430 360 436 361
rect 298 358 304 359
rect 110 347 116 348
rect 110 343 111 347
rect 115 343 116 347
rect 110 342 116 343
rect 134 344 140 345
rect 112 331 114 342
rect 134 340 135 344
rect 139 340 140 344
rect 134 339 140 340
rect 136 331 138 339
rect 111 330 115 331
rect 111 325 115 326
rect 135 330 139 331
rect 135 325 139 326
rect 112 322 114 325
rect 134 324 140 325
rect 110 321 116 322
rect 110 317 111 321
rect 115 317 116 321
rect 134 320 135 324
rect 139 320 140 324
rect 134 319 140 320
rect 110 316 116 317
rect 110 304 116 305
rect 110 300 111 304
rect 115 300 116 304
rect 110 299 116 300
rect 150 303 156 304
rect 150 299 151 303
rect 155 299 156 303
rect 112 271 114 299
rect 150 298 156 299
rect 152 271 154 298
rect 160 288 162 358
rect 190 344 196 345
rect 190 340 191 344
rect 195 340 196 344
rect 190 339 196 340
rect 262 344 268 345
rect 262 340 263 344
rect 267 340 268 344
rect 262 339 268 340
rect 342 344 348 345
rect 342 340 343 344
rect 347 340 348 344
rect 342 339 348 340
rect 414 344 420 345
rect 414 340 415 344
rect 419 340 420 344
rect 414 339 420 340
rect 192 331 194 339
rect 264 331 266 339
rect 344 331 346 339
rect 416 331 418 339
rect 191 330 195 331
rect 191 325 195 326
rect 199 330 203 331
rect 199 325 203 326
rect 263 330 267 331
rect 263 325 267 326
rect 287 330 291 331
rect 287 325 291 326
rect 343 330 347 331
rect 343 325 347 326
rect 375 330 379 331
rect 375 325 379 326
rect 415 330 419 331
rect 415 325 419 326
rect 455 330 459 331
rect 455 325 459 326
rect 198 324 204 325
rect 198 320 199 324
rect 203 320 204 324
rect 198 319 204 320
rect 286 324 292 325
rect 286 320 287 324
rect 291 320 292 324
rect 286 319 292 320
rect 374 324 380 325
rect 374 320 375 324
rect 379 320 380 324
rect 374 319 380 320
rect 454 324 460 325
rect 454 320 455 324
rect 459 320 460 324
rect 454 319 460 320
rect 480 304 482 382
rect 512 366 514 385
rect 510 365 516 366
rect 510 361 511 365
rect 515 361 516 365
rect 532 364 534 402
rect 584 391 586 418
rect 624 408 626 474
rect 718 460 724 461
rect 718 456 719 460
rect 723 456 724 460
rect 718 455 724 456
rect 830 460 836 461
rect 830 456 831 460
rect 835 456 836 460
rect 830 455 836 456
rect 934 460 940 461
rect 934 456 935 460
rect 939 456 940 460
rect 934 455 940 456
rect 1038 460 1044 461
rect 1038 456 1039 460
rect 1043 456 1044 460
rect 1038 455 1044 456
rect 1142 460 1148 461
rect 1142 456 1143 460
rect 1147 456 1148 460
rect 1142 455 1148 456
rect 1222 460 1228 461
rect 1222 456 1223 460
rect 1227 456 1228 460
rect 1222 455 1228 456
rect 720 451 722 455
rect 832 451 834 455
rect 936 451 938 455
rect 1040 451 1042 455
rect 1144 451 1146 455
rect 1224 451 1226 455
rect 671 450 675 451
rect 671 445 675 446
rect 719 450 723 451
rect 719 445 723 446
rect 783 450 787 451
rect 783 445 787 446
rect 831 450 835 451
rect 831 445 835 446
rect 895 450 899 451
rect 895 445 899 446
rect 935 450 939 451
rect 935 445 939 446
rect 1007 450 1011 451
rect 1007 445 1011 446
rect 1039 450 1043 451
rect 1039 445 1043 446
rect 1127 450 1131 451
rect 1127 445 1131 446
rect 1143 450 1147 451
rect 1143 445 1147 446
rect 1223 450 1227 451
rect 1223 445 1227 446
rect 670 444 676 445
rect 670 440 671 444
rect 675 440 676 444
rect 670 439 676 440
rect 782 444 788 445
rect 782 440 783 444
rect 787 440 788 444
rect 782 439 788 440
rect 894 444 900 445
rect 894 440 895 444
rect 899 440 900 444
rect 894 439 900 440
rect 1006 444 1012 445
rect 1006 440 1007 444
rect 1011 440 1012 444
rect 1006 439 1012 440
rect 1126 444 1132 445
rect 1126 440 1127 444
rect 1131 440 1132 444
rect 1126 439 1132 440
rect 1222 444 1228 445
rect 1222 440 1223 444
rect 1227 440 1228 444
rect 1222 439 1228 440
rect 1260 424 1262 490
rect 1288 481 1290 501
rect 1328 487 1330 511
rect 1382 510 1388 511
rect 1390 515 1396 516
rect 1390 511 1391 515
rect 1395 511 1396 515
rect 1390 510 1396 511
rect 1462 515 1468 516
rect 1462 511 1463 515
rect 1467 511 1468 515
rect 1462 510 1468 511
rect 1384 487 1386 510
rect 1327 486 1331 487
rect 1327 481 1331 482
rect 1367 486 1371 487
rect 1367 481 1371 482
rect 1383 486 1387 487
rect 1392 484 1394 510
rect 1464 487 1466 510
rect 1472 500 1474 566
rect 1542 552 1548 553
rect 1542 548 1543 552
rect 1547 548 1548 552
rect 1542 547 1548 548
rect 1654 552 1660 553
rect 1654 548 1655 552
rect 1659 548 1660 552
rect 1654 547 1660 548
rect 1758 552 1764 553
rect 1758 548 1759 552
rect 1763 548 1764 552
rect 1758 547 1764 548
rect 1544 543 1546 547
rect 1656 543 1658 547
rect 1760 543 1762 547
rect 1527 542 1531 543
rect 1527 537 1531 538
rect 1543 542 1547 543
rect 1543 537 1547 538
rect 1615 542 1619 543
rect 1615 537 1619 538
rect 1655 542 1659 543
rect 1655 537 1659 538
rect 1711 542 1715 543
rect 1711 537 1715 538
rect 1759 542 1763 543
rect 1759 537 1763 538
rect 1799 542 1803 543
rect 1799 537 1803 538
rect 1526 536 1532 537
rect 1526 532 1527 536
rect 1531 532 1532 536
rect 1526 531 1532 532
rect 1614 536 1620 537
rect 1614 532 1615 536
rect 1619 532 1620 536
rect 1614 531 1620 532
rect 1710 536 1716 537
rect 1710 532 1711 536
rect 1715 532 1716 536
rect 1710 531 1716 532
rect 1798 536 1804 537
rect 1798 532 1799 536
rect 1803 532 1804 536
rect 1798 531 1804 532
rect 1836 516 1838 582
rect 1880 574 1882 593
rect 1878 573 1884 574
rect 1878 569 1879 573
rect 1883 569 1884 573
rect 1904 572 1906 606
rect 1936 599 1938 622
rect 2024 599 2026 622
rect 2104 599 2106 622
rect 1935 598 1939 599
rect 1935 593 1939 594
rect 1983 598 1987 599
rect 1983 593 1987 594
rect 2023 598 2027 599
rect 2023 593 2027 594
rect 2087 598 2091 599
rect 2087 593 2091 594
rect 2103 598 2107 599
rect 2103 593 2107 594
rect 1984 574 1986 593
rect 2088 574 2090 593
rect 2176 588 2178 622
rect 2184 599 2186 622
rect 2248 612 2250 682
rect 2276 628 2278 698
rect 2312 690 2314 709
rect 2392 690 2394 709
rect 2310 689 2316 690
rect 2310 685 2311 689
rect 2315 685 2316 689
rect 2310 684 2316 685
rect 2390 689 2396 690
rect 2390 685 2391 689
rect 2395 685 2396 689
rect 2412 688 2414 722
rect 2456 715 2458 738
rect 2455 714 2459 715
rect 2455 709 2459 710
rect 2456 690 2458 709
rect 2464 704 2466 738
rect 2472 728 2474 794
rect 2502 783 2508 784
rect 2502 779 2503 783
rect 2507 779 2508 783
rect 2502 778 2508 779
rect 2504 771 2506 778
rect 2503 770 2507 771
rect 2503 765 2507 766
rect 2504 762 2506 765
rect 2502 761 2508 762
rect 2502 757 2503 761
rect 2507 757 2508 761
rect 2502 756 2508 757
rect 2502 744 2508 745
rect 2502 740 2503 744
rect 2507 740 2508 744
rect 2502 739 2508 740
rect 2470 727 2476 728
rect 2470 723 2471 727
rect 2475 723 2476 727
rect 2470 722 2476 723
rect 2504 715 2506 739
rect 2503 714 2507 715
rect 2503 709 2507 710
rect 2462 703 2468 704
rect 2462 699 2463 703
rect 2467 699 2468 703
rect 2462 698 2468 699
rect 2454 689 2460 690
rect 2504 689 2506 709
rect 2390 684 2396 685
rect 2410 687 2416 688
rect 2410 683 2411 687
rect 2415 683 2416 687
rect 2454 685 2455 689
rect 2459 685 2460 689
rect 2502 688 2508 689
rect 2454 684 2460 685
rect 2470 687 2476 688
rect 2410 682 2416 683
rect 2470 683 2471 687
rect 2475 683 2476 687
rect 2502 684 2503 688
rect 2507 684 2508 688
rect 2502 683 2508 684
rect 2470 682 2476 683
rect 2294 668 2300 669
rect 2294 664 2295 668
rect 2299 664 2300 668
rect 2294 663 2300 664
rect 2374 668 2380 669
rect 2374 664 2375 668
rect 2379 664 2380 668
rect 2374 663 2380 664
rect 2438 668 2444 669
rect 2438 664 2439 668
rect 2443 664 2444 668
rect 2438 663 2444 664
rect 2296 655 2298 663
rect 2376 655 2378 663
rect 2440 655 2442 663
rect 2295 654 2299 655
rect 2295 649 2299 650
rect 2311 654 2315 655
rect 2311 649 2315 650
rect 2375 654 2379 655
rect 2375 649 2379 650
rect 2383 654 2387 655
rect 2383 649 2387 650
rect 2439 654 2443 655
rect 2439 649 2443 650
rect 2310 648 2316 649
rect 2310 644 2311 648
rect 2315 644 2316 648
rect 2310 643 2316 644
rect 2382 648 2388 649
rect 2382 644 2383 648
rect 2387 644 2388 648
rect 2382 643 2388 644
rect 2438 648 2444 649
rect 2438 644 2439 648
rect 2443 644 2444 648
rect 2438 643 2444 644
rect 2254 627 2260 628
rect 2254 623 2255 627
rect 2259 623 2260 627
rect 2254 622 2260 623
rect 2274 627 2280 628
rect 2274 623 2275 627
rect 2279 623 2280 627
rect 2274 622 2280 623
rect 2326 627 2332 628
rect 2326 623 2327 627
rect 2331 623 2332 627
rect 2326 622 2332 623
rect 2342 627 2348 628
rect 2342 623 2343 627
rect 2347 623 2348 627
rect 2342 622 2348 623
rect 2398 627 2404 628
rect 2398 623 2399 627
rect 2403 623 2404 627
rect 2398 622 2404 623
rect 2454 627 2460 628
rect 2454 623 2455 627
rect 2459 623 2460 627
rect 2454 622 2460 623
rect 2462 627 2468 628
rect 2462 623 2463 627
rect 2467 623 2468 627
rect 2462 622 2468 623
rect 2246 611 2252 612
rect 2246 607 2247 611
rect 2251 607 2252 611
rect 2246 606 2252 607
rect 2256 599 2258 622
rect 2328 599 2330 622
rect 2344 608 2346 622
rect 2342 607 2348 608
rect 2342 603 2343 607
rect 2347 603 2348 607
rect 2342 602 2348 603
rect 2400 599 2402 622
rect 2406 611 2412 612
rect 2406 607 2407 611
rect 2411 607 2412 611
rect 2406 606 2412 607
rect 2183 598 2187 599
rect 2183 593 2187 594
rect 2255 598 2259 599
rect 2255 593 2259 594
rect 2279 598 2283 599
rect 2327 598 2331 599
rect 2279 593 2283 594
rect 2298 595 2304 596
rect 2174 587 2180 588
rect 2174 583 2175 587
rect 2179 583 2180 587
rect 2174 582 2180 583
rect 2184 574 2186 593
rect 2280 574 2282 593
rect 2298 591 2299 595
rect 2303 591 2304 595
rect 2327 593 2331 594
rect 2375 598 2379 599
rect 2375 593 2379 594
rect 2399 598 2403 599
rect 2399 593 2403 594
rect 2298 590 2304 591
rect 1982 573 1988 574
rect 1878 568 1884 569
rect 1902 571 1908 572
rect 1902 567 1903 571
rect 1907 567 1908 571
rect 1982 569 1983 573
rect 1987 569 1988 573
rect 1982 568 1988 569
rect 2086 573 2092 574
rect 2086 569 2087 573
rect 2091 569 2092 573
rect 2182 573 2188 574
rect 2086 568 2092 569
rect 2158 571 2164 572
rect 1902 566 1908 567
rect 2158 567 2159 571
rect 2163 567 2164 571
rect 2182 569 2183 573
rect 2187 569 2188 573
rect 2182 568 2188 569
rect 2278 573 2284 574
rect 2278 569 2279 573
rect 2283 569 2284 573
rect 2300 572 2302 590
rect 2376 574 2378 593
rect 2382 587 2388 588
rect 2382 583 2383 587
rect 2387 583 2388 587
rect 2382 582 2388 583
rect 2374 573 2380 574
rect 2278 568 2284 569
rect 2298 571 2304 572
rect 2158 566 2164 567
rect 2298 567 2299 571
rect 2303 567 2304 571
rect 2374 569 2375 573
rect 2379 569 2380 573
rect 2374 568 2380 569
rect 2298 566 2304 567
rect 1862 552 1868 553
rect 1862 548 1863 552
rect 1867 548 1868 552
rect 1862 547 1868 548
rect 1966 552 1972 553
rect 1966 548 1967 552
rect 1971 548 1972 552
rect 1966 547 1972 548
rect 2070 552 2076 553
rect 2070 548 2071 552
rect 2075 548 2076 552
rect 2070 547 2076 548
rect 1864 543 1866 547
rect 1968 543 1970 547
rect 2072 543 2074 547
rect 1863 542 1867 543
rect 1863 537 1867 538
rect 1887 542 1891 543
rect 1887 537 1891 538
rect 1967 542 1971 543
rect 1967 537 1971 538
rect 1975 542 1979 543
rect 1975 537 1979 538
rect 2063 542 2067 543
rect 2063 537 2067 538
rect 2071 542 2075 543
rect 2071 537 2075 538
rect 2151 542 2155 543
rect 2151 537 2155 538
rect 1886 536 1892 537
rect 1886 532 1887 536
rect 1891 532 1892 536
rect 1886 531 1892 532
rect 1974 536 1980 537
rect 1974 532 1975 536
rect 1979 532 1980 536
rect 1974 531 1980 532
rect 2062 536 2068 537
rect 2062 532 2063 536
rect 2067 532 2068 536
rect 2062 531 2068 532
rect 2150 536 2156 537
rect 2150 532 2151 536
rect 2155 532 2156 536
rect 2150 531 2156 532
rect 1542 515 1548 516
rect 1542 511 1543 515
rect 1547 511 1548 515
rect 1542 510 1548 511
rect 1550 515 1556 516
rect 1550 511 1551 515
rect 1555 511 1556 515
rect 1550 510 1556 511
rect 1630 515 1636 516
rect 1630 511 1631 515
rect 1635 511 1636 515
rect 1630 510 1636 511
rect 1726 515 1732 516
rect 1726 511 1727 515
rect 1731 511 1732 515
rect 1726 510 1732 511
rect 1814 515 1820 516
rect 1814 511 1815 515
rect 1819 511 1820 515
rect 1814 510 1820 511
rect 1834 515 1840 516
rect 1834 511 1835 515
rect 1839 511 1840 515
rect 1834 510 1840 511
rect 1902 515 1908 516
rect 1902 511 1903 515
rect 1907 511 1908 515
rect 1902 510 1908 511
rect 1990 515 1996 516
rect 1990 511 1991 515
rect 1995 511 1996 515
rect 1990 510 1996 511
rect 2078 515 2084 516
rect 2078 511 2079 515
rect 2083 511 2084 515
rect 2078 510 2084 511
rect 2150 515 2156 516
rect 2150 511 2151 515
rect 2155 511 2156 515
rect 2150 510 2156 511
rect 1470 499 1476 500
rect 1470 495 1471 499
rect 1475 495 1476 499
rect 1470 494 1476 495
rect 1544 487 1546 510
rect 1552 492 1554 510
rect 1550 491 1556 492
rect 1550 487 1551 491
rect 1555 487 1556 491
rect 1632 487 1634 510
rect 1718 495 1724 496
rect 1718 491 1719 495
rect 1723 491 1724 495
rect 1718 490 1724 491
rect 1431 486 1435 487
rect 1383 481 1387 482
rect 1390 483 1396 484
rect 1286 480 1292 481
rect 1286 476 1287 480
rect 1291 476 1292 480
rect 1286 475 1292 476
rect 1286 463 1292 464
rect 1286 459 1287 463
rect 1291 459 1292 463
rect 1328 461 1330 481
rect 1368 462 1370 481
rect 1390 479 1391 483
rect 1395 479 1396 483
rect 1431 481 1435 482
rect 1463 486 1467 487
rect 1463 481 1467 482
rect 1519 486 1523 487
rect 1519 481 1523 482
rect 1543 486 1547 487
rect 1550 486 1556 487
rect 1615 486 1619 487
rect 1543 481 1547 482
rect 1615 481 1619 482
rect 1631 486 1635 487
rect 1631 481 1635 482
rect 1711 486 1715 487
rect 1711 481 1715 482
rect 1390 478 1396 479
rect 1432 462 1434 481
rect 1520 462 1522 481
rect 1550 475 1556 476
rect 1550 471 1551 475
rect 1555 471 1556 475
rect 1550 470 1556 471
rect 1366 461 1372 462
rect 1286 458 1292 459
rect 1326 460 1332 461
rect 1288 451 1290 458
rect 1326 456 1327 460
rect 1331 456 1332 460
rect 1366 457 1367 461
rect 1371 457 1372 461
rect 1366 456 1372 457
rect 1430 461 1436 462
rect 1430 457 1431 461
rect 1435 457 1436 461
rect 1430 456 1436 457
rect 1518 461 1524 462
rect 1518 457 1519 461
rect 1523 457 1524 461
rect 1518 456 1524 457
rect 1526 459 1532 460
rect 1326 455 1332 456
rect 1526 455 1527 459
rect 1531 455 1532 459
rect 1526 454 1532 455
rect 1287 450 1291 451
rect 1287 445 1291 446
rect 1288 442 1290 445
rect 1326 443 1332 444
rect 1286 441 1292 442
rect 1286 437 1287 441
rect 1291 437 1292 441
rect 1326 439 1327 443
rect 1331 439 1332 443
rect 1326 438 1332 439
rect 1350 440 1356 441
rect 1286 436 1292 437
rect 1328 431 1330 438
rect 1350 436 1351 440
rect 1355 436 1356 440
rect 1350 435 1356 436
rect 1414 440 1420 441
rect 1414 436 1415 440
rect 1419 436 1420 440
rect 1414 435 1420 436
rect 1502 440 1508 441
rect 1502 436 1503 440
rect 1507 436 1508 440
rect 1502 435 1508 436
rect 1352 431 1354 435
rect 1416 431 1418 435
rect 1504 431 1506 435
rect 1327 430 1331 431
rect 1327 425 1331 426
rect 1351 430 1355 431
rect 1351 425 1355 426
rect 1415 430 1419 431
rect 1415 425 1419 426
rect 1423 430 1427 431
rect 1423 425 1427 426
rect 1503 430 1507 431
rect 1503 425 1507 426
rect 1511 430 1515 431
rect 1511 425 1515 426
rect 1286 424 1292 425
rect 686 423 692 424
rect 686 419 687 423
rect 691 419 692 423
rect 686 418 692 419
rect 798 423 804 424
rect 798 419 799 423
rect 803 419 804 423
rect 798 418 804 419
rect 910 423 916 424
rect 910 419 911 423
rect 915 419 916 423
rect 910 418 916 419
rect 918 423 924 424
rect 918 419 919 423
rect 923 419 924 423
rect 918 418 924 419
rect 1022 423 1028 424
rect 1022 419 1023 423
rect 1027 419 1028 423
rect 1022 418 1028 419
rect 1142 423 1148 424
rect 1142 419 1143 423
rect 1147 419 1148 423
rect 1142 418 1148 419
rect 1238 423 1244 424
rect 1238 419 1239 423
rect 1243 419 1244 423
rect 1238 418 1244 419
rect 1258 423 1264 424
rect 1258 419 1259 423
rect 1263 419 1264 423
rect 1286 420 1287 424
rect 1291 420 1292 424
rect 1328 422 1330 425
rect 1350 424 1356 425
rect 1286 419 1292 420
rect 1326 421 1332 422
rect 1258 418 1264 419
rect 622 407 628 408
rect 622 403 623 407
rect 627 403 628 407
rect 622 402 628 403
rect 688 391 690 418
rect 800 391 802 418
rect 912 391 914 418
rect 583 390 587 391
rect 583 385 587 386
rect 591 390 595 391
rect 591 385 595 386
rect 671 390 675 391
rect 671 385 675 386
rect 687 390 691 391
rect 687 385 691 386
rect 751 390 755 391
rect 751 385 755 386
rect 799 390 803 391
rect 799 385 803 386
rect 823 390 827 391
rect 895 390 899 391
rect 823 385 827 386
rect 842 387 848 388
rect 592 366 594 385
rect 672 366 674 385
rect 752 366 754 385
rect 824 366 826 385
rect 842 383 843 387
rect 847 383 848 387
rect 895 385 899 386
rect 911 390 915 391
rect 911 385 915 386
rect 842 382 848 383
rect 590 365 596 366
rect 510 360 516 361
rect 530 363 536 364
rect 530 359 531 363
rect 535 359 536 363
rect 590 361 591 365
rect 595 361 596 365
rect 670 365 676 366
rect 590 360 596 361
rect 638 363 644 364
rect 530 358 536 359
rect 638 359 639 363
rect 643 359 644 363
rect 670 361 671 365
rect 675 361 676 365
rect 670 360 676 361
rect 750 365 756 366
rect 750 361 751 365
rect 755 361 756 365
rect 750 360 756 361
rect 822 365 828 366
rect 822 361 823 365
rect 827 361 828 365
rect 844 364 846 382
rect 896 366 898 385
rect 920 380 922 418
rect 990 407 996 408
rect 990 403 991 407
rect 995 403 996 407
rect 990 402 996 403
rect 967 390 971 391
rect 967 385 971 386
rect 918 379 924 380
rect 918 375 919 379
rect 923 375 924 379
rect 918 374 924 375
rect 968 366 970 385
rect 894 365 900 366
rect 822 360 828 361
rect 842 363 848 364
rect 638 358 644 359
rect 842 359 843 363
rect 847 359 848 363
rect 894 361 895 365
rect 899 361 900 365
rect 894 360 900 361
rect 966 365 972 366
rect 966 361 967 365
rect 971 361 972 365
rect 992 364 994 402
rect 1024 391 1026 418
rect 1144 391 1146 418
rect 1240 391 1242 418
rect 1288 391 1290 419
rect 1326 417 1327 421
rect 1331 417 1332 421
rect 1350 420 1351 424
rect 1355 420 1356 424
rect 1350 419 1356 420
rect 1422 424 1428 425
rect 1422 420 1423 424
rect 1427 420 1428 424
rect 1422 419 1428 420
rect 1510 424 1516 425
rect 1510 420 1511 424
rect 1515 420 1516 424
rect 1510 419 1516 420
rect 1326 416 1332 417
rect 1528 411 1530 454
rect 1520 409 1530 411
rect 1326 404 1332 405
rect 1326 400 1327 404
rect 1331 400 1332 404
rect 1326 399 1332 400
rect 1366 403 1372 404
rect 1366 399 1367 403
rect 1371 399 1372 403
rect 1023 390 1027 391
rect 1023 385 1027 386
rect 1039 390 1043 391
rect 1039 385 1043 386
rect 1111 390 1115 391
rect 1111 385 1115 386
rect 1143 390 1147 391
rect 1143 385 1147 386
rect 1183 390 1187 391
rect 1183 385 1187 386
rect 1239 390 1243 391
rect 1239 385 1243 386
rect 1287 390 1291 391
rect 1287 385 1291 386
rect 1040 366 1042 385
rect 1070 379 1076 380
rect 1070 375 1071 379
rect 1075 375 1076 379
rect 1070 374 1076 375
rect 1038 365 1044 366
rect 966 360 972 361
rect 990 363 996 364
rect 842 358 848 359
rect 990 359 991 363
rect 995 359 996 363
rect 1038 361 1039 365
rect 1043 361 1044 365
rect 1038 360 1044 361
rect 990 358 996 359
rect 494 344 500 345
rect 494 340 495 344
rect 499 340 500 344
rect 494 339 500 340
rect 574 344 580 345
rect 574 340 575 344
rect 579 340 580 344
rect 574 339 580 340
rect 496 331 498 339
rect 576 331 578 339
rect 495 330 499 331
rect 495 325 499 326
rect 543 330 547 331
rect 543 325 547 326
rect 575 330 579 331
rect 575 325 579 326
rect 631 330 635 331
rect 631 325 635 326
rect 542 324 548 325
rect 542 320 543 324
rect 547 320 548 324
rect 542 319 548 320
rect 630 324 636 325
rect 630 320 631 324
rect 635 320 636 324
rect 630 319 636 320
rect 214 303 220 304
rect 214 299 215 303
rect 219 299 220 303
rect 214 298 220 299
rect 302 303 308 304
rect 302 299 303 303
rect 307 299 308 303
rect 302 298 308 299
rect 334 303 340 304
rect 334 299 335 303
rect 339 299 340 303
rect 334 298 340 299
rect 390 303 396 304
rect 390 299 391 303
rect 395 299 396 303
rect 390 298 396 299
rect 470 303 476 304
rect 470 299 471 303
rect 475 299 476 303
rect 470 298 476 299
rect 478 303 484 304
rect 478 299 479 303
rect 483 299 484 303
rect 478 298 484 299
rect 558 303 564 304
rect 558 299 559 303
rect 563 299 564 303
rect 558 298 564 299
rect 158 287 164 288
rect 158 283 159 287
rect 163 283 164 287
rect 158 282 164 283
rect 216 271 218 298
rect 304 271 306 298
rect 111 270 115 271
rect 111 265 115 266
rect 151 270 155 271
rect 151 265 155 266
rect 215 270 219 271
rect 215 265 219 266
rect 231 270 235 271
rect 231 265 235 266
rect 303 270 307 271
rect 303 265 307 266
rect 327 270 331 271
rect 327 265 331 266
rect 112 245 114 265
rect 152 246 154 265
rect 232 246 234 265
rect 328 246 330 265
rect 336 260 338 298
rect 392 271 394 298
rect 472 271 474 298
rect 542 287 548 288
rect 542 283 543 287
rect 547 283 548 287
rect 542 282 548 283
rect 391 270 395 271
rect 346 267 352 268
rect 346 263 347 267
rect 351 263 352 267
rect 391 265 395 266
rect 423 270 427 271
rect 423 265 427 266
rect 471 270 475 271
rect 471 265 475 266
rect 519 270 523 271
rect 519 265 523 266
rect 346 262 352 263
rect 334 259 340 260
rect 334 255 335 259
rect 339 255 340 259
rect 334 254 340 255
rect 150 245 156 246
rect 110 244 116 245
rect 110 240 111 244
rect 115 240 116 244
rect 150 241 151 245
rect 155 241 156 245
rect 150 240 156 241
rect 230 245 236 246
rect 230 241 231 245
rect 235 241 236 245
rect 326 245 332 246
rect 230 240 236 241
rect 262 243 268 244
rect 110 239 116 240
rect 262 239 263 243
rect 267 239 268 243
rect 326 241 327 245
rect 331 241 332 245
rect 348 244 350 262
rect 424 246 426 265
rect 520 246 522 265
rect 422 245 428 246
rect 326 240 332 241
rect 346 243 352 244
rect 262 238 268 239
rect 346 239 347 243
rect 351 239 352 243
rect 422 241 423 245
rect 427 241 428 245
rect 422 240 428 241
rect 518 245 524 246
rect 518 241 519 245
rect 523 241 524 245
rect 544 244 546 282
rect 560 271 562 298
rect 640 288 642 358
rect 654 344 660 345
rect 654 340 655 344
rect 659 340 660 344
rect 654 339 660 340
rect 734 344 740 345
rect 734 340 735 344
rect 739 340 740 344
rect 734 339 740 340
rect 806 344 812 345
rect 806 340 807 344
rect 811 340 812 344
rect 806 339 812 340
rect 878 344 884 345
rect 878 340 879 344
rect 883 340 884 344
rect 878 339 884 340
rect 950 344 956 345
rect 950 340 951 344
rect 955 340 956 344
rect 950 339 956 340
rect 1022 344 1028 345
rect 1022 340 1023 344
rect 1027 340 1028 344
rect 1022 339 1028 340
rect 656 331 658 339
rect 736 331 738 339
rect 808 331 810 339
rect 880 331 882 339
rect 952 331 954 339
rect 1024 331 1026 339
rect 655 330 659 331
rect 655 325 659 326
rect 727 330 731 331
rect 727 325 731 326
rect 735 330 739 331
rect 735 325 739 326
rect 807 330 811 331
rect 807 325 811 326
rect 823 330 827 331
rect 823 325 827 326
rect 879 330 883 331
rect 879 325 883 326
rect 927 330 931 331
rect 927 325 931 326
rect 951 330 955 331
rect 951 325 955 326
rect 1023 330 1027 331
rect 1023 325 1027 326
rect 1031 330 1035 331
rect 1031 325 1035 326
rect 726 324 732 325
rect 726 320 727 324
rect 731 320 732 324
rect 726 319 732 320
rect 822 324 828 325
rect 822 320 823 324
rect 827 320 828 324
rect 822 319 828 320
rect 926 324 932 325
rect 926 320 927 324
rect 931 320 932 324
rect 926 319 932 320
rect 1030 324 1036 325
rect 1030 320 1031 324
rect 1035 320 1036 324
rect 1030 319 1036 320
rect 1072 304 1074 374
rect 1112 366 1114 385
rect 1184 366 1186 385
rect 1240 366 1242 385
rect 1110 365 1116 366
rect 1110 361 1111 365
rect 1115 361 1116 365
rect 1110 360 1116 361
rect 1182 365 1188 366
rect 1182 361 1183 365
rect 1187 361 1188 365
rect 1238 365 1244 366
rect 1288 365 1290 385
rect 1328 375 1330 399
rect 1366 398 1372 399
rect 1374 403 1380 404
rect 1374 399 1375 403
rect 1379 399 1380 403
rect 1374 398 1380 399
rect 1438 403 1444 404
rect 1438 399 1439 403
rect 1443 399 1444 403
rect 1438 398 1444 399
rect 1368 375 1370 398
rect 1376 380 1378 398
rect 1374 379 1380 380
rect 1374 375 1375 379
rect 1379 375 1380 379
rect 1440 375 1442 398
rect 1520 388 1522 409
rect 1552 404 1554 470
rect 1616 462 1618 481
rect 1712 462 1714 481
rect 1614 461 1620 462
rect 1614 457 1615 461
rect 1619 457 1620 461
rect 1614 456 1620 457
rect 1710 461 1716 462
rect 1710 457 1711 461
rect 1715 457 1716 461
rect 1720 460 1722 490
rect 1728 487 1730 510
rect 1816 487 1818 510
rect 1904 487 1906 510
rect 1992 487 1994 510
rect 2055 500 2059 501
rect 2054 495 2060 496
rect 2054 491 2055 495
rect 2059 491 2060 495
rect 2054 490 2060 491
rect 2080 487 2082 510
rect 1727 486 1731 487
rect 1727 481 1731 482
rect 1815 486 1819 487
rect 1815 481 1819 482
rect 1903 486 1907 487
rect 1903 481 1907 482
rect 1927 486 1931 487
rect 1927 481 1931 482
rect 1991 486 1995 487
rect 1991 481 1995 482
rect 2055 486 2059 487
rect 2079 486 2083 487
rect 2055 481 2059 482
rect 2070 483 2076 484
rect 1816 462 1818 481
rect 1928 462 1930 481
rect 2056 462 2058 481
rect 2070 479 2071 483
rect 2075 479 2076 483
rect 2079 481 2083 482
rect 2070 478 2076 479
rect 1814 461 1820 462
rect 1710 456 1716 457
rect 1718 459 1724 460
rect 1718 455 1719 459
rect 1723 455 1724 459
rect 1814 457 1815 461
rect 1819 457 1820 461
rect 1814 456 1820 457
rect 1926 461 1932 462
rect 1926 457 1927 461
rect 1931 457 1932 461
rect 2054 461 2060 462
rect 1926 456 1932 457
rect 2022 459 2028 460
rect 1718 454 1724 455
rect 2022 455 2023 459
rect 2027 455 2028 459
rect 2054 457 2055 461
rect 2059 457 2060 461
rect 2072 460 2074 478
rect 2152 476 2154 510
rect 2160 500 2162 566
rect 2166 552 2172 553
rect 2166 548 2167 552
rect 2171 548 2172 552
rect 2166 547 2172 548
rect 2262 552 2268 553
rect 2262 548 2263 552
rect 2267 548 2268 552
rect 2262 547 2268 548
rect 2358 552 2364 553
rect 2358 548 2359 552
rect 2363 548 2364 552
rect 2358 547 2364 548
rect 2168 543 2170 547
rect 2264 543 2266 547
rect 2360 543 2362 547
rect 2167 542 2171 543
rect 2167 537 2171 538
rect 2247 542 2251 543
rect 2247 537 2251 538
rect 2263 542 2267 543
rect 2263 537 2267 538
rect 2343 542 2347 543
rect 2343 537 2347 538
rect 2359 542 2363 543
rect 2359 537 2363 538
rect 2246 536 2252 537
rect 2246 532 2247 536
rect 2251 532 2252 536
rect 2246 531 2252 532
rect 2342 536 2348 537
rect 2342 532 2343 536
rect 2347 532 2348 536
rect 2342 531 2348 532
rect 2384 516 2386 582
rect 2408 572 2410 606
rect 2456 599 2458 622
rect 2455 598 2459 599
rect 2455 593 2459 594
rect 2456 574 2458 593
rect 2464 588 2466 622
rect 2472 612 2474 682
rect 2502 671 2508 672
rect 2502 667 2503 671
rect 2507 667 2508 671
rect 2502 666 2508 667
rect 2504 655 2506 666
rect 2503 654 2507 655
rect 2503 649 2507 650
rect 2504 646 2506 649
rect 2502 645 2508 646
rect 2502 641 2503 645
rect 2507 641 2508 645
rect 2502 640 2508 641
rect 2502 628 2508 629
rect 2502 624 2503 628
rect 2507 624 2508 628
rect 2502 623 2508 624
rect 2470 611 2476 612
rect 2470 607 2471 611
rect 2475 607 2476 611
rect 2470 606 2476 607
rect 2504 599 2506 623
rect 2503 598 2507 599
rect 2503 593 2507 594
rect 2462 587 2468 588
rect 2462 583 2463 587
rect 2467 583 2468 587
rect 2462 582 2468 583
rect 2454 573 2460 574
rect 2504 573 2506 593
rect 2406 571 2412 572
rect 2406 567 2407 571
rect 2411 567 2412 571
rect 2454 569 2455 573
rect 2459 569 2460 573
rect 2502 572 2508 573
rect 2454 568 2460 569
rect 2462 571 2468 572
rect 2406 566 2412 567
rect 2462 567 2463 571
rect 2467 567 2468 571
rect 2502 568 2503 572
rect 2507 568 2508 572
rect 2502 567 2508 568
rect 2462 566 2468 567
rect 2438 552 2444 553
rect 2438 548 2439 552
rect 2443 548 2444 552
rect 2438 547 2444 548
rect 2440 543 2442 547
rect 2439 542 2443 543
rect 2439 537 2443 538
rect 2438 536 2444 537
rect 2438 532 2439 536
rect 2443 532 2444 536
rect 2438 531 2444 532
rect 2166 515 2172 516
rect 2166 511 2167 515
rect 2171 511 2172 515
rect 2166 510 2172 511
rect 2262 515 2268 516
rect 2262 511 2263 515
rect 2267 511 2268 515
rect 2262 510 2268 511
rect 2270 515 2276 516
rect 2270 511 2271 515
rect 2275 511 2276 515
rect 2270 510 2276 511
rect 2358 515 2364 516
rect 2358 511 2359 515
rect 2363 511 2364 515
rect 2358 510 2364 511
rect 2382 515 2388 516
rect 2382 511 2383 515
rect 2387 511 2388 515
rect 2382 510 2388 511
rect 2454 515 2460 516
rect 2454 511 2455 515
rect 2459 511 2460 515
rect 2454 510 2460 511
rect 2158 499 2164 500
rect 2158 495 2159 499
rect 2163 495 2164 499
rect 2158 494 2164 495
rect 2168 487 2170 510
rect 2264 487 2266 510
rect 2272 501 2274 510
rect 2271 500 2275 501
rect 2271 495 2275 496
rect 2360 487 2362 510
rect 2456 487 2458 510
rect 2167 486 2171 487
rect 2167 481 2171 482
rect 2191 486 2195 487
rect 2191 481 2195 482
rect 2263 486 2267 487
rect 2263 481 2267 482
rect 2335 486 2339 487
rect 2359 486 2363 487
rect 2335 481 2339 482
rect 2350 483 2356 484
rect 2150 475 2156 476
rect 2150 471 2151 475
rect 2155 471 2156 475
rect 2150 470 2156 471
rect 2192 462 2194 481
rect 2336 462 2338 481
rect 2350 479 2351 483
rect 2355 479 2356 483
rect 2359 481 2363 482
rect 2455 486 2459 487
rect 2455 481 2459 482
rect 2350 478 2356 479
rect 2190 461 2196 462
rect 2054 456 2060 457
rect 2070 459 2076 460
rect 2022 454 2028 455
rect 2070 455 2071 459
rect 2075 455 2076 459
rect 2190 457 2191 461
rect 2195 457 2196 461
rect 2190 456 2196 457
rect 2334 461 2340 462
rect 2334 457 2335 461
rect 2339 457 2340 461
rect 2352 460 2354 478
rect 2456 462 2458 481
rect 2464 476 2466 566
rect 2502 555 2508 556
rect 2502 551 2503 555
rect 2507 551 2508 555
rect 2502 550 2508 551
rect 2504 543 2506 550
rect 2503 542 2507 543
rect 2503 537 2507 538
rect 2504 534 2506 537
rect 2502 533 2508 534
rect 2502 529 2503 533
rect 2507 529 2508 533
rect 2502 528 2508 529
rect 2502 516 2508 517
rect 2502 512 2503 516
rect 2507 512 2508 516
rect 2502 511 2508 512
rect 2478 499 2484 500
rect 2478 495 2479 499
rect 2483 495 2484 499
rect 2478 494 2484 495
rect 2462 475 2468 476
rect 2462 471 2463 475
rect 2467 471 2468 475
rect 2462 470 2468 471
rect 2454 461 2460 462
rect 2334 456 2340 457
rect 2350 459 2356 460
rect 2070 454 2076 455
rect 2350 455 2351 459
rect 2355 455 2356 459
rect 2454 457 2455 461
rect 2459 457 2460 461
rect 2454 456 2460 457
rect 2470 459 2476 460
rect 2350 454 2356 455
rect 2470 455 2471 459
rect 2475 455 2476 459
rect 2470 454 2476 455
rect 1598 440 1604 441
rect 1598 436 1599 440
rect 1603 436 1604 440
rect 1598 435 1604 436
rect 1694 440 1700 441
rect 1694 436 1695 440
rect 1699 436 1700 440
rect 1694 435 1700 436
rect 1798 440 1804 441
rect 1798 436 1799 440
rect 1803 436 1804 440
rect 1798 435 1804 436
rect 1910 440 1916 441
rect 1910 436 1911 440
rect 1915 436 1916 440
rect 1910 435 1916 436
rect 1600 431 1602 435
rect 1696 431 1698 435
rect 1800 431 1802 435
rect 1912 431 1914 435
rect 1599 430 1603 431
rect 1599 425 1603 426
rect 1679 430 1683 431
rect 1679 425 1683 426
rect 1695 430 1699 431
rect 1695 425 1699 426
rect 1775 430 1779 431
rect 1775 425 1779 426
rect 1799 430 1803 431
rect 1799 425 1803 426
rect 1887 430 1891 431
rect 1887 425 1891 426
rect 1911 430 1915 431
rect 1911 425 1915 426
rect 2015 430 2019 431
rect 2015 425 2019 426
rect 1598 424 1604 425
rect 1598 420 1599 424
rect 1603 420 1604 424
rect 1598 419 1604 420
rect 1678 424 1684 425
rect 1678 420 1679 424
rect 1683 420 1684 424
rect 1678 419 1684 420
rect 1774 424 1780 425
rect 1774 420 1775 424
rect 1779 420 1780 424
rect 1774 419 1780 420
rect 1886 424 1892 425
rect 1886 420 1887 424
rect 1891 420 1892 424
rect 1886 419 1892 420
rect 2014 424 2020 425
rect 2014 420 2015 424
rect 2019 420 2020 424
rect 2014 419 2020 420
rect 1526 403 1532 404
rect 1526 399 1527 403
rect 1531 399 1532 403
rect 1526 398 1532 399
rect 1550 403 1556 404
rect 1550 399 1551 403
rect 1555 399 1556 403
rect 1550 398 1556 399
rect 1614 403 1620 404
rect 1614 399 1615 403
rect 1619 399 1620 403
rect 1614 398 1620 399
rect 1694 403 1700 404
rect 1694 399 1695 403
rect 1699 399 1700 403
rect 1694 398 1700 399
rect 1790 403 1796 404
rect 1790 399 1791 403
rect 1795 399 1796 403
rect 1790 398 1796 399
rect 1814 403 1820 404
rect 1814 399 1815 403
rect 1819 399 1820 403
rect 1814 398 1820 399
rect 1902 403 1908 404
rect 1902 399 1903 403
rect 1907 399 1908 403
rect 1902 398 1908 399
rect 1518 387 1524 388
rect 1518 383 1519 387
rect 1523 383 1524 387
rect 1518 382 1524 383
rect 1528 375 1530 398
rect 1616 375 1618 398
rect 1696 375 1698 398
rect 1754 379 1760 380
rect 1754 375 1755 379
rect 1759 375 1760 379
rect 1792 375 1794 398
rect 1327 374 1331 375
rect 1327 369 1331 370
rect 1367 374 1371 375
rect 1374 374 1380 375
rect 1439 374 1443 375
rect 1367 369 1371 370
rect 1439 369 1443 370
rect 1527 374 1531 375
rect 1527 369 1531 370
rect 1615 374 1619 375
rect 1615 369 1619 370
rect 1679 374 1683 375
rect 1679 369 1683 370
rect 1695 374 1699 375
rect 1695 369 1699 370
rect 1735 374 1739 375
rect 1754 374 1760 375
rect 1791 374 1795 375
rect 1735 369 1739 370
rect 1182 360 1188 361
rect 1230 363 1236 364
rect 1230 359 1231 363
rect 1235 359 1236 363
rect 1238 361 1239 365
rect 1243 361 1244 365
rect 1238 360 1244 361
rect 1286 364 1292 365
rect 1286 360 1287 364
rect 1291 360 1292 364
rect 1286 359 1292 360
rect 1230 358 1236 359
rect 1094 344 1100 345
rect 1094 340 1095 344
rect 1099 340 1100 344
rect 1094 339 1100 340
rect 1166 344 1172 345
rect 1166 340 1167 344
rect 1171 340 1172 344
rect 1166 339 1172 340
rect 1222 344 1228 345
rect 1222 340 1223 344
rect 1227 340 1228 344
rect 1222 339 1228 340
rect 1096 331 1098 339
rect 1168 331 1170 339
rect 1224 331 1226 339
rect 1095 330 1099 331
rect 1095 325 1099 326
rect 1135 330 1139 331
rect 1135 325 1139 326
rect 1167 330 1171 331
rect 1167 325 1171 326
rect 1223 330 1227 331
rect 1223 325 1227 326
rect 1134 324 1140 325
rect 1134 320 1135 324
rect 1139 320 1140 324
rect 1134 319 1140 320
rect 1222 324 1228 325
rect 1222 320 1223 324
rect 1227 320 1228 324
rect 1222 319 1228 320
rect 646 303 652 304
rect 646 299 647 303
rect 651 299 652 303
rect 646 298 652 299
rect 742 303 748 304
rect 742 299 743 303
rect 747 299 748 303
rect 742 298 748 299
rect 838 303 844 304
rect 838 299 839 303
rect 843 299 844 303
rect 838 298 844 299
rect 942 303 948 304
rect 942 299 943 303
rect 947 299 948 303
rect 942 298 948 299
rect 950 303 956 304
rect 950 299 951 303
rect 955 299 956 303
rect 950 298 956 299
rect 1046 303 1052 304
rect 1046 299 1047 303
rect 1051 299 1052 303
rect 1046 298 1052 299
rect 1070 303 1076 304
rect 1070 299 1071 303
rect 1075 299 1076 303
rect 1070 298 1076 299
rect 1150 303 1156 304
rect 1150 299 1151 303
rect 1155 299 1156 303
rect 1150 298 1156 299
rect 638 287 644 288
rect 638 283 639 287
rect 643 283 644 287
rect 638 282 644 283
rect 648 271 650 298
rect 744 271 746 298
rect 840 271 842 298
rect 944 271 946 298
rect 559 270 563 271
rect 559 265 563 266
rect 615 270 619 271
rect 647 270 651 271
rect 615 265 619 266
rect 634 267 640 268
rect 616 246 618 265
rect 634 263 635 267
rect 639 263 640 267
rect 647 265 651 266
rect 711 270 715 271
rect 711 265 715 266
rect 743 270 747 271
rect 743 265 747 266
rect 807 270 811 271
rect 807 265 811 266
rect 839 270 843 271
rect 839 265 843 266
rect 903 270 907 271
rect 943 270 947 271
rect 903 265 907 266
rect 922 267 928 268
rect 634 262 640 263
rect 614 245 620 246
rect 518 240 524 241
rect 542 243 548 244
rect 346 238 352 239
rect 542 239 543 243
rect 547 239 548 243
rect 614 241 615 245
rect 619 241 620 245
rect 636 244 638 262
rect 642 259 648 260
rect 642 255 643 259
rect 647 255 648 259
rect 642 254 648 255
rect 614 240 620 241
rect 634 243 640 244
rect 542 238 548 239
rect 634 239 635 243
rect 639 239 640 243
rect 634 238 640 239
rect 110 227 116 228
rect 110 223 111 227
rect 115 223 116 227
rect 110 222 116 223
rect 134 224 140 225
rect 112 211 114 222
rect 134 220 135 224
rect 139 220 140 224
rect 134 219 140 220
rect 214 224 220 225
rect 214 220 215 224
rect 219 220 220 224
rect 214 219 220 220
rect 136 211 138 219
rect 216 211 218 219
rect 111 210 115 211
rect 111 205 115 206
rect 135 210 139 211
rect 135 205 139 206
rect 159 210 163 211
rect 159 205 163 206
rect 215 210 219 211
rect 215 205 219 206
rect 239 210 243 211
rect 239 205 243 206
rect 112 202 114 205
rect 158 204 164 205
rect 110 201 116 202
rect 110 197 111 201
rect 115 197 116 201
rect 158 200 159 204
rect 163 200 164 204
rect 158 199 164 200
rect 238 204 244 205
rect 238 200 239 204
rect 243 200 244 204
rect 238 199 244 200
rect 110 196 116 197
rect 110 184 116 185
rect 110 180 111 184
rect 115 180 116 184
rect 110 179 116 180
rect 174 183 180 184
rect 174 179 175 183
rect 179 179 180 183
rect 112 139 114 179
rect 174 178 180 179
rect 182 183 188 184
rect 182 179 183 183
rect 187 179 188 183
rect 182 178 188 179
rect 254 183 260 184
rect 254 179 255 183
rect 259 179 260 183
rect 254 178 260 179
rect 176 139 178 178
rect 111 138 115 139
rect 111 133 115 134
rect 151 138 155 139
rect 151 133 155 134
rect 175 138 179 139
rect 184 136 186 178
rect 256 139 258 178
rect 264 168 266 238
rect 310 224 316 225
rect 310 220 311 224
rect 315 220 316 224
rect 310 219 316 220
rect 406 224 412 225
rect 406 220 407 224
rect 411 220 412 224
rect 406 219 412 220
rect 502 224 508 225
rect 502 220 503 224
rect 507 220 508 224
rect 502 219 508 220
rect 598 224 604 225
rect 598 220 599 224
rect 603 220 604 224
rect 598 219 604 220
rect 312 211 314 219
rect 408 211 410 219
rect 504 211 506 219
rect 600 211 602 219
rect 311 210 315 211
rect 311 205 315 206
rect 327 210 331 211
rect 327 205 331 206
rect 407 210 411 211
rect 407 205 411 206
rect 415 210 419 211
rect 415 205 419 206
rect 503 210 507 211
rect 503 205 507 206
rect 511 210 515 211
rect 511 205 515 206
rect 599 210 603 211
rect 599 205 603 206
rect 607 210 611 211
rect 607 205 611 206
rect 326 204 332 205
rect 326 200 327 204
rect 331 200 332 204
rect 326 199 332 200
rect 414 204 420 205
rect 414 200 415 204
rect 419 200 420 204
rect 414 199 420 200
rect 510 204 516 205
rect 510 200 511 204
rect 515 200 516 204
rect 510 199 516 200
rect 606 204 612 205
rect 606 200 607 204
rect 611 200 612 204
rect 606 199 612 200
rect 644 184 646 254
rect 712 246 714 265
rect 808 246 810 265
rect 904 246 906 265
rect 922 263 923 267
rect 927 263 928 267
rect 943 265 947 266
rect 922 262 928 263
rect 710 245 716 246
rect 710 241 711 245
rect 715 241 716 245
rect 710 240 716 241
rect 806 245 812 246
rect 806 241 807 245
rect 811 241 812 245
rect 902 245 908 246
rect 806 240 812 241
rect 878 243 884 244
rect 878 239 879 243
rect 883 239 884 243
rect 902 241 903 245
rect 907 241 908 245
rect 924 244 926 262
rect 952 260 954 298
rect 1048 271 1050 298
rect 1152 271 1154 298
rect 1232 288 1234 358
rect 1328 349 1330 369
rect 1670 363 1676 364
rect 1670 359 1671 363
rect 1675 359 1676 363
rect 1670 358 1676 359
rect 1326 348 1332 349
rect 1286 347 1292 348
rect 1286 343 1287 347
rect 1291 343 1292 347
rect 1326 344 1327 348
rect 1331 344 1332 348
rect 1326 343 1332 344
rect 1286 342 1292 343
rect 1288 331 1290 342
rect 1326 331 1332 332
rect 1287 330 1291 331
rect 1326 327 1327 331
rect 1331 327 1332 331
rect 1326 326 1332 327
rect 1662 328 1668 329
rect 1287 325 1291 326
rect 1288 322 1290 325
rect 1328 323 1330 326
rect 1662 324 1663 328
rect 1667 324 1668 328
rect 1662 323 1668 324
rect 1327 322 1331 323
rect 1286 321 1292 322
rect 1286 317 1287 321
rect 1291 317 1292 321
rect 1327 317 1331 318
rect 1351 322 1355 323
rect 1351 317 1355 318
rect 1431 322 1435 323
rect 1431 317 1435 318
rect 1527 322 1531 323
rect 1527 317 1531 318
rect 1623 322 1627 323
rect 1623 317 1627 318
rect 1663 322 1667 323
rect 1663 317 1667 318
rect 1286 316 1292 317
rect 1328 314 1330 317
rect 1350 316 1356 317
rect 1326 313 1332 314
rect 1326 309 1327 313
rect 1331 309 1332 313
rect 1350 312 1351 316
rect 1355 312 1356 316
rect 1350 311 1356 312
rect 1430 316 1436 317
rect 1430 312 1431 316
rect 1435 312 1436 316
rect 1430 311 1436 312
rect 1526 316 1532 317
rect 1526 312 1527 316
rect 1531 312 1532 316
rect 1526 311 1532 312
rect 1622 316 1628 317
rect 1622 312 1623 316
rect 1627 312 1628 316
rect 1622 311 1628 312
rect 1326 308 1332 309
rect 1286 304 1292 305
rect 1238 303 1244 304
rect 1238 299 1239 303
rect 1243 299 1244 303
rect 1238 298 1244 299
rect 1278 303 1284 304
rect 1278 299 1279 303
rect 1283 299 1284 303
rect 1286 300 1287 304
rect 1291 300 1292 304
rect 1286 299 1292 300
rect 1278 298 1284 299
rect 1222 287 1228 288
rect 1222 283 1223 287
rect 1227 283 1228 287
rect 1222 282 1228 283
rect 1230 287 1236 288
rect 1230 283 1231 287
rect 1235 283 1236 287
rect 1230 282 1236 283
rect 1007 270 1011 271
rect 1007 265 1011 266
rect 1047 270 1051 271
rect 1047 265 1051 266
rect 1111 270 1115 271
rect 1111 265 1115 266
rect 1151 270 1155 271
rect 1151 265 1155 266
rect 1215 270 1219 271
rect 1215 265 1219 266
rect 950 259 956 260
rect 950 255 951 259
rect 955 255 956 259
rect 950 254 956 255
rect 998 259 1004 260
rect 998 255 999 259
rect 1003 255 1004 259
rect 998 254 1004 255
rect 902 240 908 241
rect 922 243 928 244
rect 878 238 884 239
rect 922 239 923 243
rect 927 239 928 243
rect 922 238 928 239
rect 694 224 700 225
rect 694 220 695 224
rect 699 220 700 224
rect 694 219 700 220
rect 790 224 796 225
rect 790 220 791 224
rect 795 220 796 224
rect 790 219 796 220
rect 696 211 698 219
rect 792 211 794 219
rect 695 210 699 211
rect 695 205 699 206
rect 783 210 787 211
rect 783 205 787 206
rect 791 210 795 211
rect 791 205 795 206
rect 871 210 875 211
rect 871 205 875 206
rect 694 204 700 205
rect 694 200 695 204
rect 699 200 700 204
rect 694 199 700 200
rect 782 204 788 205
rect 782 200 783 204
rect 787 200 788 204
rect 782 199 788 200
rect 870 204 876 205
rect 870 200 871 204
rect 875 200 876 204
rect 870 199 876 200
rect 342 183 348 184
rect 342 179 343 183
rect 347 179 348 183
rect 342 178 348 179
rect 350 183 356 184
rect 350 179 351 183
rect 355 179 356 183
rect 350 178 356 179
rect 430 183 436 184
rect 430 179 431 183
rect 435 179 436 183
rect 430 178 436 179
rect 526 183 532 184
rect 526 179 527 183
rect 531 179 532 183
rect 526 178 532 179
rect 622 183 628 184
rect 622 179 623 183
rect 627 179 628 183
rect 622 178 628 179
rect 642 183 648 184
rect 642 179 643 183
rect 647 179 648 183
rect 642 178 648 179
rect 710 183 716 184
rect 710 179 711 183
rect 715 179 716 183
rect 710 178 716 179
rect 718 183 724 184
rect 718 179 719 183
rect 723 179 724 183
rect 718 178 724 179
rect 798 183 804 184
rect 798 179 799 183
rect 803 179 804 183
rect 798 178 804 179
rect 814 183 820 184
rect 814 179 815 183
rect 819 179 820 183
rect 814 178 820 179
rect 262 167 268 168
rect 262 163 263 167
rect 267 163 268 167
rect 262 162 268 163
rect 344 139 346 178
rect 352 160 354 178
rect 350 159 356 160
rect 350 155 351 159
rect 355 155 356 159
rect 350 154 356 155
rect 432 139 434 178
rect 528 139 530 178
rect 624 139 626 178
rect 642 163 648 164
rect 642 159 643 163
rect 647 159 648 163
rect 642 158 648 159
rect 207 138 211 139
rect 175 133 179 134
rect 182 135 188 136
rect 112 113 114 133
rect 152 114 154 133
rect 182 131 183 135
rect 187 131 188 135
rect 207 133 211 134
rect 255 138 259 139
rect 255 133 259 134
rect 263 138 267 139
rect 263 133 267 134
rect 319 138 323 139
rect 319 133 323 134
rect 343 138 347 139
rect 343 133 347 134
rect 375 138 379 139
rect 375 133 379 134
rect 431 138 435 139
rect 431 133 435 134
rect 487 138 491 139
rect 487 133 491 134
rect 527 138 531 139
rect 527 133 531 134
rect 551 138 555 139
rect 551 133 555 134
rect 623 138 627 139
rect 623 133 627 134
rect 182 130 188 131
rect 208 114 210 133
rect 264 114 266 133
rect 320 114 322 133
rect 376 114 378 133
rect 432 114 434 133
rect 488 114 490 133
rect 552 114 554 133
rect 624 114 626 133
rect 150 113 156 114
rect 110 112 116 113
rect 110 108 111 112
rect 115 108 116 112
rect 150 109 151 113
rect 155 109 156 113
rect 150 108 156 109
rect 206 113 212 114
rect 206 109 207 113
rect 211 109 212 113
rect 206 108 212 109
rect 262 113 268 114
rect 262 109 263 113
rect 267 109 268 113
rect 262 108 268 109
rect 318 113 324 114
rect 318 109 319 113
rect 323 109 324 113
rect 318 108 324 109
rect 374 113 380 114
rect 374 109 375 113
rect 379 109 380 113
rect 374 108 380 109
rect 430 113 436 114
rect 430 109 431 113
rect 435 109 436 113
rect 430 108 436 109
rect 486 113 492 114
rect 486 109 487 113
rect 491 109 492 113
rect 486 108 492 109
rect 550 113 556 114
rect 550 109 551 113
rect 555 109 556 113
rect 550 108 556 109
rect 622 113 628 114
rect 622 109 623 113
rect 627 109 628 113
rect 644 112 646 158
rect 712 139 714 178
rect 687 138 691 139
rect 687 133 691 134
rect 711 138 715 139
rect 720 136 722 178
rect 800 139 802 178
rect 816 164 818 178
rect 880 168 882 238
rect 886 224 892 225
rect 886 220 887 224
rect 891 220 892 224
rect 886 219 892 220
rect 990 224 996 225
rect 990 220 991 224
rect 995 220 996 224
rect 990 219 996 220
rect 888 211 890 219
rect 992 211 994 219
rect 887 210 891 211
rect 887 205 891 206
rect 959 210 963 211
rect 959 205 963 206
rect 991 210 995 211
rect 991 205 995 206
rect 958 204 964 205
rect 958 200 959 204
rect 963 200 964 204
rect 958 199 964 200
rect 1000 184 1002 254
rect 1008 246 1010 265
rect 1112 246 1114 265
rect 1216 246 1218 265
rect 1006 245 1012 246
rect 1006 241 1007 245
rect 1011 241 1012 245
rect 1006 240 1012 241
rect 1110 245 1116 246
rect 1110 241 1111 245
rect 1115 241 1116 245
rect 1110 240 1116 241
rect 1214 245 1220 246
rect 1214 241 1215 245
rect 1219 241 1220 245
rect 1224 244 1226 282
rect 1240 271 1242 298
rect 1280 280 1282 298
rect 1278 279 1284 280
rect 1278 275 1279 279
rect 1283 275 1284 279
rect 1278 274 1284 275
rect 1288 271 1290 299
rect 1326 296 1332 297
rect 1672 296 1674 358
rect 1680 350 1682 369
rect 1736 350 1738 369
rect 1678 349 1684 350
rect 1678 345 1679 349
rect 1683 345 1684 349
rect 1678 344 1684 345
rect 1734 349 1740 350
rect 1734 345 1735 349
rect 1739 345 1740 349
rect 1756 348 1758 374
rect 1791 369 1795 370
rect 1807 374 1811 375
rect 1807 369 1811 370
rect 1808 350 1810 369
rect 1816 364 1818 398
rect 1904 375 1906 398
rect 2024 388 2026 454
rect 2038 440 2044 441
rect 2038 436 2039 440
rect 2043 436 2044 440
rect 2038 435 2044 436
rect 2174 440 2180 441
rect 2174 436 2175 440
rect 2179 436 2180 440
rect 2174 435 2180 436
rect 2318 440 2324 441
rect 2318 436 2319 440
rect 2323 436 2324 440
rect 2318 435 2324 436
rect 2438 440 2444 441
rect 2438 436 2439 440
rect 2443 436 2444 440
rect 2438 435 2444 436
rect 2040 431 2042 435
rect 2176 431 2178 435
rect 2320 431 2322 435
rect 2440 431 2442 435
rect 2039 430 2043 431
rect 2039 425 2043 426
rect 2159 430 2163 431
rect 2159 425 2163 426
rect 2175 430 2179 431
rect 2175 425 2179 426
rect 2311 430 2315 431
rect 2311 425 2315 426
rect 2319 430 2323 431
rect 2319 425 2323 426
rect 2439 430 2443 431
rect 2439 425 2443 426
rect 2158 424 2164 425
rect 2158 420 2159 424
rect 2163 420 2164 424
rect 2158 419 2164 420
rect 2310 424 2316 425
rect 2310 420 2311 424
rect 2315 420 2316 424
rect 2310 419 2316 420
rect 2438 424 2444 425
rect 2438 420 2439 424
rect 2443 420 2444 424
rect 2438 419 2444 420
rect 2030 403 2036 404
rect 2030 399 2031 403
rect 2035 399 2036 403
rect 2030 398 2036 399
rect 2174 403 2180 404
rect 2174 399 2175 403
rect 2179 399 2180 403
rect 2174 398 2180 399
rect 2326 403 2332 404
rect 2326 399 2327 403
rect 2331 399 2332 403
rect 2326 398 2332 399
rect 2334 403 2340 404
rect 2334 399 2335 403
rect 2339 399 2340 403
rect 2334 398 2340 399
rect 2454 403 2460 404
rect 2454 399 2455 403
rect 2459 399 2460 403
rect 2454 398 2460 399
rect 2462 403 2468 404
rect 2462 399 2463 403
rect 2467 399 2468 403
rect 2462 398 2468 399
rect 2022 387 2028 388
rect 2022 383 2023 387
rect 2027 383 2028 387
rect 2022 382 2028 383
rect 2032 375 2034 398
rect 2176 375 2178 398
rect 2328 375 2330 398
rect 2336 380 2338 398
rect 2334 379 2340 380
rect 2334 375 2335 379
rect 2339 375 2340 379
rect 2456 375 2458 398
rect 1903 374 1907 375
rect 1903 369 1907 370
rect 2023 374 2027 375
rect 2023 369 2027 370
rect 2031 374 2035 375
rect 2031 369 2035 370
rect 2159 374 2163 375
rect 2159 369 2163 370
rect 2175 374 2179 375
rect 2175 369 2179 370
rect 2303 374 2307 375
rect 2303 369 2307 370
rect 2327 374 2331 375
rect 2334 374 2340 375
rect 2455 374 2459 375
rect 2327 369 2331 370
rect 2455 369 2459 370
rect 1814 363 1820 364
rect 1814 359 1815 363
rect 1819 359 1820 363
rect 1814 358 1820 359
rect 1904 350 1906 369
rect 2024 350 2026 369
rect 2160 350 2162 369
rect 2304 350 2306 369
rect 2456 350 2458 369
rect 2464 364 2466 398
rect 2472 388 2474 454
rect 2470 387 2476 388
rect 2470 383 2471 387
rect 2475 383 2476 387
rect 2470 382 2476 383
rect 2462 363 2468 364
rect 2462 359 2463 363
rect 2467 359 2468 363
rect 2462 358 2468 359
rect 1806 349 1812 350
rect 1734 344 1740 345
rect 1754 347 1760 348
rect 1754 343 1755 347
rect 1759 343 1760 347
rect 1806 345 1807 349
rect 1811 345 1812 349
rect 1806 344 1812 345
rect 1902 349 1908 350
rect 1902 345 1903 349
rect 1907 345 1908 349
rect 1902 344 1908 345
rect 2022 349 2028 350
rect 2022 345 2023 349
rect 2027 345 2028 349
rect 2022 344 2028 345
rect 2158 349 2164 350
rect 2158 345 2159 349
rect 2163 345 2164 349
rect 2158 344 2164 345
rect 2302 349 2308 350
rect 2302 345 2303 349
rect 2307 345 2308 349
rect 2454 349 2460 350
rect 2302 344 2308 345
rect 2318 347 2324 348
rect 1754 342 1760 343
rect 2318 343 2319 347
rect 2323 343 2324 347
rect 2454 345 2455 349
rect 2459 345 2460 349
rect 2480 348 2482 494
rect 2504 487 2506 511
rect 2503 486 2507 487
rect 2503 481 2507 482
rect 2504 461 2506 481
rect 2502 460 2508 461
rect 2502 456 2503 460
rect 2507 456 2508 460
rect 2502 455 2508 456
rect 2502 443 2508 444
rect 2502 439 2503 443
rect 2507 439 2508 443
rect 2502 438 2508 439
rect 2504 431 2506 438
rect 2503 430 2507 431
rect 2503 425 2507 426
rect 2504 422 2506 425
rect 2502 421 2508 422
rect 2502 417 2503 421
rect 2507 417 2508 421
rect 2502 416 2508 417
rect 2502 404 2508 405
rect 2502 400 2503 404
rect 2507 400 2508 404
rect 2502 399 2508 400
rect 2504 375 2506 399
rect 2503 374 2507 375
rect 2503 369 2507 370
rect 2504 349 2506 369
rect 2502 348 2508 349
rect 2454 344 2460 345
rect 2478 347 2484 348
rect 2318 342 2324 343
rect 2478 343 2479 347
rect 2483 343 2484 347
rect 2502 344 2503 348
rect 2507 344 2508 348
rect 2502 343 2508 344
rect 2478 342 2484 343
rect 1718 328 1724 329
rect 1718 324 1719 328
rect 1723 324 1724 328
rect 1718 323 1724 324
rect 1790 328 1796 329
rect 1790 324 1791 328
rect 1795 324 1796 328
rect 1790 323 1796 324
rect 1886 328 1892 329
rect 1886 324 1887 328
rect 1891 324 1892 328
rect 1886 323 1892 324
rect 2006 328 2012 329
rect 2006 324 2007 328
rect 2011 324 2012 328
rect 2006 323 2012 324
rect 2142 328 2148 329
rect 2142 324 2143 328
rect 2147 324 2148 328
rect 2142 323 2148 324
rect 2286 328 2292 329
rect 2286 324 2287 328
rect 2291 324 2292 328
rect 2286 323 2292 324
rect 1711 322 1715 323
rect 1711 317 1715 318
rect 1719 322 1723 323
rect 1719 317 1723 318
rect 1791 322 1795 323
rect 1791 317 1795 318
rect 1807 322 1811 323
rect 1807 317 1811 318
rect 1887 322 1891 323
rect 1887 317 1891 318
rect 1911 322 1915 323
rect 1911 317 1915 318
rect 2007 322 2011 323
rect 2007 317 2011 318
rect 2023 322 2027 323
rect 2023 317 2027 318
rect 2143 322 2147 323
rect 2143 317 2147 318
rect 2151 322 2155 323
rect 2151 317 2155 318
rect 2287 322 2291 323
rect 2287 317 2291 318
rect 1710 316 1716 317
rect 1710 312 1711 316
rect 1715 312 1716 316
rect 1710 311 1716 312
rect 1806 316 1812 317
rect 1806 312 1807 316
rect 1811 312 1812 316
rect 1806 311 1812 312
rect 1910 316 1916 317
rect 1910 312 1911 316
rect 1915 312 1916 316
rect 1910 311 1916 312
rect 2022 316 2028 317
rect 2022 312 2023 316
rect 2027 312 2028 316
rect 2022 311 2028 312
rect 2150 316 2156 317
rect 2150 312 2151 316
rect 2155 312 2156 316
rect 2150 311 2156 312
rect 2286 316 2292 317
rect 2286 312 2287 316
rect 2291 312 2292 316
rect 2286 311 2292 312
rect 1326 292 1327 296
rect 1331 292 1332 296
rect 1326 291 1332 292
rect 1366 295 1372 296
rect 1366 291 1367 295
rect 1371 291 1372 295
rect 1239 270 1243 271
rect 1239 265 1243 266
rect 1287 270 1291 271
rect 1328 267 1330 291
rect 1366 290 1372 291
rect 1446 295 1452 296
rect 1446 291 1447 295
rect 1451 291 1452 295
rect 1446 290 1452 291
rect 1542 295 1548 296
rect 1542 291 1543 295
rect 1547 291 1548 295
rect 1542 290 1548 291
rect 1550 295 1556 296
rect 1550 291 1551 295
rect 1555 291 1556 295
rect 1550 290 1556 291
rect 1638 295 1644 296
rect 1638 291 1639 295
rect 1643 291 1644 295
rect 1638 290 1644 291
rect 1670 295 1676 296
rect 1670 291 1671 295
rect 1675 291 1676 295
rect 1670 290 1676 291
rect 1726 295 1732 296
rect 1726 291 1727 295
rect 1731 291 1732 295
rect 1726 290 1732 291
rect 1822 295 1828 296
rect 1822 291 1823 295
rect 1827 291 1828 295
rect 1822 290 1828 291
rect 1926 295 1932 296
rect 1926 291 1927 295
rect 1931 291 1932 295
rect 1926 290 1932 291
rect 2038 295 2044 296
rect 2038 291 2039 295
rect 2043 291 2044 295
rect 2038 290 2044 291
rect 2166 295 2172 296
rect 2166 291 2167 295
rect 2171 291 2172 295
rect 2166 290 2172 291
rect 2302 295 2308 296
rect 2302 291 2303 295
rect 2307 291 2308 295
rect 2302 290 2308 291
rect 2310 295 2316 296
rect 2310 291 2311 295
rect 2315 291 2316 295
rect 2310 290 2316 291
rect 1368 267 1370 290
rect 1448 267 1450 290
rect 1544 267 1546 290
rect 1287 265 1291 266
rect 1327 266 1331 267
rect 1288 245 1290 265
rect 1327 261 1331 262
rect 1367 266 1371 267
rect 1367 261 1371 262
rect 1439 266 1443 267
rect 1439 261 1443 262
rect 1447 266 1451 267
rect 1447 261 1451 262
rect 1535 266 1539 267
rect 1535 261 1539 262
rect 1543 266 1547 267
rect 1552 264 1554 290
rect 1640 267 1642 290
rect 1728 267 1730 290
rect 1806 279 1812 280
rect 1806 275 1807 279
rect 1811 275 1812 279
rect 1806 274 1812 275
rect 1631 266 1635 267
rect 1543 261 1547 262
rect 1550 263 1556 264
rect 1286 244 1292 245
rect 1214 240 1220 241
rect 1222 243 1228 244
rect 1222 239 1223 243
rect 1227 239 1228 243
rect 1286 240 1287 244
rect 1291 240 1292 244
rect 1328 241 1330 261
rect 1368 242 1370 261
rect 1440 242 1442 261
rect 1536 242 1538 261
rect 1550 259 1551 263
rect 1555 259 1556 263
rect 1631 261 1635 262
rect 1639 266 1643 267
rect 1639 261 1643 262
rect 1727 266 1731 267
rect 1727 261 1731 262
rect 1738 263 1744 264
rect 1550 258 1556 259
rect 1632 242 1634 261
rect 1728 242 1730 261
rect 1738 259 1739 263
rect 1743 259 1744 263
rect 1738 258 1744 259
rect 1366 241 1372 242
rect 1286 239 1292 240
rect 1326 240 1332 241
rect 1222 238 1228 239
rect 1326 236 1327 240
rect 1331 236 1332 240
rect 1366 237 1367 241
rect 1371 237 1372 241
rect 1366 236 1372 237
rect 1438 241 1444 242
rect 1438 237 1439 241
rect 1443 237 1444 241
rect 1438 236 1444 237
rect 1534 241 1540 242
rect 1534 237 1535 241
rect 1539 237 1540 241
rect 1630 241 1636 242
rect 1534 236 1540 237
rect 1606 239 1612 240
rect 1326 235 1332 236
rect 1606 235 1607 239
rect 1611 235 1612 239
rect 1630 237 1631 241
rect 1635 237 1636 241
rect 1630 236 1636 237
rect 1726 241 1732 242
rect 1726 237 1727 241
rect 1731 237 1732 241
rect 1726 236 1732 237
rect 1606 234 1612 235
rect 1286 227 1292 228
rect 1094 224 1100 225
rect 1094 220 1095 224
rect 1099 220 1100 224
rect 1094 219 1100 220
rect 1198 224 1204 225
rect 1198 220 1199 224
rect 1203 220 1204 224
rect 1286 223 1287 227
rect 1291 223 1292 227
rect 1286 222 1292 223
rect 1326 223 1332 224
rect 1198 219 1204 220
rect 1096 211 1098 219
rect 1200 211 1202 219
rect 1288 211 1290 222
rect 1326 219 1327 223
rect 1331 219 1332 223
rect 1326 218 1332 219
rect 1350 220 1356 221
rect 1328 211 1330 218
rect 1350 216 1351 220
rect 1355 216 1356 220
rect 1350 215 1356 216
rect 1422 220 1428 221
rect 1422 216 1423 220
rect 1427 216 1428 220
rect 1422 215 1428 216
rect 1518 220 1524 221
rect 1518 216 1519 220
rect 1523 216 1524 220
rect 1518 215 1524 216
rect 1352 211 1354 215
rect 1424 211 1426 215
rect 1520 211 1522 215
rect 1047 210 1051 211
rect 1047 205 1051 206
rect 1095 210 1099 211
rect 1095 205 1099 206
rect 1135 210 1139 211
rect 1135 205 1139 206
rect 1199 210 1203 211
rect 1199 205 1203 206
rect 1287 210 1291 211
rect 1287 205 1291 206
rect 1327 210 1331 211
rect 1327 205 1331 206
rect 1351 210 1355 211
rect 1351 205 1355 206
rect 1391 210 1395 211
rect 1391 205 1395 206
rect 1423 210 1427 211
rect 1423 205 1427 206
rect 1495 210 1499 211
rect 1495 205 1499 206
rect 1519 210 1523 211
rect 1519 205 1523 206
rect 1599 210 1603 211
rect 1599 205 1603 206
rect 1046 204 1052 205
rect 1046 200 1047 204
rect 1051 200 1052 204
rect 1046 199 1052 200
rect 1134 204 1140 205
rect 1134 200 1135 204
rect 1139 200 1140 204
rect 1288 202 1290 205
rect 1328 202 1330 205
rect 1390 204 1396 205
rect 1134 199 1140 200
rect 1286 201 1292 202
rect 1286 197 1287 201
rect 1291 197 1292 201
rect 1286 196 1292 197
rect 1326 201 1332 202
rect 1326 197 1327 201
rect 1331 197 1332 201
rect 1390 200 1391 204
rect 1395 200 1396 204
rect 1390 199 1396 200
rect 1494 204 1500 205
rect 1494 200 1495 204
rect 1499 200 1500 204
rect 1494 199 1500 200
rect 1598 204 1604 205
rect 1598 200 1599 204
rect 1603 200 1604 204
rect 1598 199 1604 200
rect 1326 196 1332 197
rect 1286 184 1292 185
rect 886 183 892 184
rect 886 179 887 183
rect 891 179 892 183
rect 886 178 892 179
rect 974 183 980 184
rect 974 179 975 183
rect 979 179 980 183
rect 974 178 980 179
rect 998 183 1004 184
rect 998 179 999 183
rect 1003 179 1004 183
rect 998 178 1004 179
rect 1062 183 1068 184
rect 1062 179 1063 183
rect 1067 179 1068 183
rect 1062 178 1068 179
rect 1150 183 1156 184
rect 1150 179 1151 183
rect 1155 179 1156 183
rect 1286 180 1287 184
rect 1291 180 1292 184
rect 1286 179 1292 180
rect 1326 184 1332 185
rect 1326 180 1327 184
rect 1331 180 1332 184
rect 1326 179 1332 180
rect 1406 183 1412 184
rect 1406 179 1407 183
rect 1411 179 1412 183
rect 1150 178 1156 179
rect 878 167 884 168
rect 814 163 820 164
rect 814 159 815 163
rect 819 159 820 163
rect 878 163 879 167
rect 883 163 884 167
rect 878 162 884 163
rect 814 158 820 159
rect 888 139 890 178
rect 976 139 978 178
rect 1064 139 1066 178
rect 1152 139 1154 178
rect 1218 167 1224 168
rect 1218 163 1219 167
rect 1223 163 1224 167
rect 1218 162 1224 163
rect 751 138 755 139
rect 711 133 715 134
rect 718 135 724 136
rect 688 114 690 133
rect 718 131 719 135
rect 723 131 724 135
rect 751 133 755 134
rect 799 138 803 139
rect 799 133 803 134
rect 815 138 819 139
rect 815 133 819 134
rect 879 138 883 139
rect 879 133 883 134
rect 887 138 891 139
rect 887 133 891 134
rect 943 138 947 139
rect 943 133 947 134
rect 975 138 979 139
rect 975 133 979 134
rect 1007 138 1011 139
rect 1007 133 1011 134
rect 1063 138 1067 139
rect 1063 133 1067 134
rect 1071 138 1075 139
rect 1071 133 1075 134
rect 1135 138 1139 139
rect 1135 133 1139 134
rect 1151 138 1155 139
rect 1151 133 1155 134
rect 1199 138 1203 139
rect 1199 133 1203 134
rect 718 130 724 131
rect 752 114 754 133
rect 816 114 818 133
rect 880 114 882 133
rect 944 114 946 133
rect 1008 114 1010 133
rect 1072 114 1074 133
rect 1136 114 1138 133
rect 1200 114 1202 133
rect 686 113 692 114
rect 622 108 628 109
rect 642 111 648 112
rect 110 107 116 108
rect 642 107 643 111
rect 647 107 648 111
rect 686 109 687 113
rect 691 109 692 113
rect 686 108 692 109
rect 750 113 756 114
rect 750 109 751 113
rect 755 109 756 113
rect 750 108 756 109
rect 814 113 820 114
rect 814 109 815 113
rect 819 109 820 113
rect 814 108 820 109
rect 878 113 884 114
rect 878 109 879 113
rect 883 109 884 113
rect 878 108 884 109
rect 942 113 948 114
rect 942 109 943 113
rect 947 109 948 113
rect 942 108 948 109
rect 1006 113 1012 114
rect 1006 109 1007 113
rect 1011 109 1012 113
rect 1006 108 1012 109
rect 1070 113 1076 114
rect 1070 109 1071 113
rect 1075 109 1076 113
rect 1070 108 1076 109
rect 1134 113 1140 114
rect 1134 109 1135 113
rect 1139 109 1140 113
rect 1134 108 1140 109
rect 1198 113 1204 114
rect 1198 109 1199 113
rect 1203 109 1204 113
rect 1220 112 1222 162
rect 1288 139 1290 179
rect 1328 139 1330 179
rect 1406 178 1412 179
rect 1414 183 1420 184
rect 1414 179 1415 183
rect 1419 179 1420 183
rect 1414 178 1420 179
rect 1510 183 1516 184
rect 1510 179 1511 183
rect 1515 179 1516 183
rect 1510 178 1516 179
rect 1526 183 1532 184
rect 1526 179 1527 183
rect 1531 179 1532 183
rect 1526 178 1532 179
rect 1408 139 1410 178
rect 1287 138 1291 139
rect 1287 133 1291 134
rect 1327 138 1331 139
rect 1327 133 1331 134
rect 1367 138 1371 139
rect 1367 133 1371 134
rect 1407 138 1411 139
rect 1416 136 1418 178
rect 1512 139 1514 178
rect 1528 164 1530 178
rect 1608 168 1610 234
rect 1614 220 1620 221
rect 1614 216 1615 220
rect 1619 216 1620 220
rect 1614 215 1620 216
rect 1710 220 1716 221
rect 1710 216 1711 220
rect 1715 216 1716 220
rect 1710 215 1716 216
rect 1616 211 1618 215
rect 1712 211 1714 215
rect 1615 210 1619 211
rect 1615 205 1619 206
rect 1711 210 1715 211
rect 1711 205 1715 206
rect 1710 204 1716 205
rect 1710 200 1711 204
rect 1715 200 1716 204
rect 1710 199 1716 200
rect 1740 184 1742 258
rect 1808 248 1810 274
rect 1824 267 1826 290
rect 1928 267 1930 290
rect 2040 267 2042 290
rect 2168 267 2170 290
rect 2304 267 2306 290
rect 1815 266 1819 267
rect 1815 261 1819 262
rect 1823 266 1827 267
rect 1823 261 1827 262
rect 1903 266 1907 267
rect 1903 261 1907 262
rect 1927 266 1931 267
rect 1927 261 1931 262
rect 1999 266 2003 267
rect 1999 261 2003 262
rect 2039 266 2043 267
rect 2039 261 2043 262
rect 2103 266 2107 267
rect 2103 261 2107 262
rect 2167 266 2171 267
rect 2167 261 2171 262
rect 2215 266 2219 267
rect 2215 261 2219 262
rect 2303 266 2307 267
rect 2312 264 2314 290
rect 2320 276 2322 342
rect 2502 331 2508 332
rect 2438 328 2444 329
rect 2438 324 2439 328
rect 2443 324 2444 328
rect 2502 327 2503 331
rect 2507 327 2508 331
rect 2502 326 2508 327
rect 2438 323 2444 324
rect 2504 323 2506 326
rect 2423 322 2427 323
rect 2423 317 2427 318
rect 2439 322 2443 323
rect 2439 317 2443 318
rect 2503 322 2507 323
rect 2503 317 2507 318
rect 2422 316 2428 317
rect 2422 312 2423 316
rect 2427 312 2428 316
rect 2504 314 2506 317
rect 2422 311 2428 312
rect 2502 313 2508 314
rect 2502 309 2503 313
rect 2507 309 2508 313
rect 2502 308 2508 309
rect 2502 296 2508 297
rect 2438 295 2444 296
rect 2438 291 2439 295
rect 2443 291 2444 295
rect 2438 290 2444 291
rect 2462 295 2468 296
rect 2462 291 2463 295
rect 2467 291 2468 295
rect 2502 292 2503 296
rect 2507 292 2508 296
rect 2502 291 2508 292
rect 2462 290 2468 291
rect 2414 279 2420 280
rect 2318 275 2324 276
rect 2318 271 2319 275
rect 2323 271 2324 275
rect 2414 275 2415 279
rect 2419 275 2420 279
rect 2414 274 2420 275
rect 2318 270 2324 271
rect 2335 266 2339 267
rect 2303 261 2307 262
rect 2310 263 2316 264
rect 1806 247 1812 248
rect 1806 243 1807 247
rect 1811 243 1812 247
rect 1806 242 1812 243
rect 1816 242 1818 261
rect 1904 242 1906 261
rect 2000 242 2002 261
rect 2104 242 2106 261
rect 2216 242 2218 261
rect 2310 259 2311 263
rect 2315 259 2316 263
rect 2335 261 2339 262
rect 2310 258 2316 259
rect 2336 242 2338 261
rect 1814 241 1820 242
rect 1814 237 1815 241
rect 1819 237 1820 241
rect 1814 236 1820 237
rect 1902 241 1908 242
rect 1902 237 1903 241
rect 1907 237 1908 241
rect 1902 236 1908 237
rect 1998 241 2004 242
rect 1998 237 1999 241
rect 2003 237 2004 241
rect 1998 236 2004 237
rect 2102 241 2108 242
rect 2102 237 2103 241
rect 2107 237 2108 241
rect 2102 236 2108 237
rect 2214 241 2220 242
rect 2214 237 2215 241
rect 2219 237 2220 241
rect 2214 236 2220 237
rect 2334 241 2340 242
rect 2334 237 2335 241
rect 2339 237 2340 241
rect 2334 236 2340 237
rect 2342 239 2348 240
rect 2342 235 2343 239
rect 2347 235 2348 239
rect 2342 234 2348 235
rect 1798 220 1804 221
rect 1798 216 1799 220
rect 1803 216 1804 220
rect 1798 215 1804 216
rect 1886 220 1892 221
rect 1886 216 1887 220
rect 1891 216 1892 220
rect 1886 215 1892 216
rect 1982 220 1988 221
rect 1982 216 1983 220
rect 1987 216 1988 220
rect 1982 215 1988 216
rect 2086 220 2092 221
rect 2086 216 2087 220
rect 2091 216 2092 220
rect 2086 215 2092 216
rect 2198 220 2204 221
rect 2198 216 2199 220
rect 2203 216 2204 220
rect 2198 215 2204 216
rect 2318 220 2324 221
rect 2318 216 2319 220
rect 2323 216 2324 220
rect 2318 215 2324 216
rect 1800 211 1802 215
rect 1888 211 1890 215
rect 1984 211 1986 215
rect 2088 211 2090 215
rect 2200 211 2202 215
rect 2320 211 2322 215
rect 1799 210 1803 211
rect 1799 205 1803 206
rect 1815 210 1819 211
rect 1815 205 1819 206
rect 1887 210 1891 211
rect 1887 205 1891 206
rect 1919 210 1923 211
rect 1919 205 1923 206
rect 1983 210 1987 211
rect 1983 205 1987 206
rect 2015 210 2019 211
rect 2015 205 2019 206
rect 2087 210 2091 211
rect 2087 205 2091 206
rect 2111 210 2115 211
rect 2111 205 2115 206
rect 2199 210 2203 211
rect 2199 205 2203 206
rect 2287 210 2291 211
rect 2287 205 2291 206
rect 2319 210 2323 211
rect 2319 205 2323 206
rect 1814 204 1820 205
rect 1814 200 1815 204
rect 1819 200 1820 204
rect 1814 199 1820 200
rect 1918 204 1924 205
rect 1918 200 1919 204
rect 1923 200 1924 204
rect 1918 199 1924 200
rect 2014 204 2020 205
rect 2014 200 2015 204
rect 2019 200 2020 204
rect 2014 199 2020 200
rect 2110 204 2116 205
rect 2110 200 2111 204
rect 2115 200 2116 204
rect 2110 199 2116 200
rect 2198 204 2204 205
rect 2198 200 2199 204
rect 2203 200 2204 204
rect 2198 199 2204 200
rect 2286 204 2292 205
rect 2286 200 2287 204
rect 2291 200 2292 204
rect 2286 199 2292 200
rect 1614 183 1620 184
rect 1614 179 1615 183
rect 1619 179 1620 183
rect 1614 178 1620 179
rect 1726 183 1732 184
rect 1726 179 1727 183
rect 1731 179 1732 183
rect 1726 178 1732 179
rect 1738 183 1744 184
rect 1738 179 1739 183
rect 1743 179 1744 183
rect 1738 178 1744 179
rect 1830 183 1836 184
rect 1830 179 1831 183
rect 1835 179 1836 183
rect 1830 178 1836 179
rect 1934 183 1940 184
rect 1934 179 1935 183
rect 1939 179 1940 183
rect 1934 178 1940 179
rect 2030 183 2036 184
rect 2030 179 2031 183
rect 2035 179 2036 183
rect 2030 178 2036 179
rect 2126 183 2132 184
rect 2126 179 2127 183
rect 2131 179 2132 183
rect 2126 178 2132 179
rect 2214 183 2220 184
rect 2214 179 2215 183
rect 2219 179 2220 183
rect 2214 178 2220 179
rect 2230 183 2236 184
rect 2230 179 2231 183
rect 2235 179 2236 183
rect 2230 178 2236 179
rect 2302 183 2308 184
rect 2302 179 2303 183
rect 2307 179 2308 183
rect 2302 178 2308 179
rect 1606 167 1612 168
rect 1526 163 1532 164
rect 1526 159 1527 163
rect 1531 159 1532 163
rect 1606 163 1607 167
rect 1611 163 1612 167
rect 1606 162 1612 163
rect 1526 158 1532 159
rect 1616 139 1618 178
rect 1728 139 1730 178
rect 1832 139 1834 178
rect 1838 167 1844 168
rect 1838 163 1839 167
rect 1843 163 1844 167
rect 1838 162 1844 163
rect 1423 138 1427 139
rect 1407 133 1411 134
rect 1414 135 1420 136
rect 1288 113 1290 133
rect 1328 113 1330 133
rect 1368 114 1370 133
rect 1414 131 1415 135
rect 1419 131 1420 135
rect 1423 133 1427 134
rect 1479 138 1483 139
rect 1479 133 1483 134
rect 1511 138 1515 139
rect 1511 133 1515 134
rect 1535 138 1539 139
rect 1535 133 1539 134
rect 1591 138 1595 139
rect 1591 133 1595 134
rect 1615 138 1619 139
rect 1615 133 1619 134
rect 1647 138 1651 139
rect 1647 133 1651 134
rect 1703 138 1707 139
rect 1703 133 1707 134
rect 1727 138 1731 139
rect 1727 133 1731 134
rect 1759 138 1763 139
rect 1759 133 1763 134
rect 1815 138 1819 139
rect 1815 133 1819 134
rect 1831 138 1835 139
rect 1831 133 1835 134
rect 1414 130 1420 131
rect 1424 114 1426 133
rect 1480 114 1482 133
rect 1536 114 1538 133
rect 1592 114 1594 133
rect 1648 114 1650 133
rect 1704 114 1706 133
rect 1760 114 1762 133
rect 1816 114 1818 133
rect 1366 113 1372 114
rect 1286 112 1292 113
rect 1198 108 1204 109
rect 1218 111 1224 112
rect 642 106 648 107
rect 1218 107 1219 111
rect 1223 107 1224 111
rect 1286 108 1287 112
rect 1291 108 1292 112
rect 1286 107 1292 108
rect 1326 112 1332 113
rect 1326 108 1327 112
rect 1331 108 1332 112
rect 1366 109 1367 113
rect 1371 109 1372 113
rect 1366 108 1372 109
rect 1422 113 1428 114
rect 1422 109 1423 113
rect 1427 109 1428 113
rect 1422 108 1428 109
rect 1478 113 1484 114
rect 1478 109 1479 113
rect 1483 109 1484 113
rect 1478 108 1484 109
rect 1534 113 1540 114
rect 1534 109 1535 113
rect 1539 109 1540 113
rect 1534 108 1540 109
rect 1590 113 1596 114
rect 1590 109 1591 113
rect 1595 109 1596 113
rect 1590 108 1596 109
rect 1646 113 1652 114
rect 1646 109 1647 113
rect 1651 109 1652 113
rect 1646 108 1652 109
rect 1702 113 1708 114
rect 1702 109 1703 113
rect 1707 109 1708 113
rect 1702 108 1708 109
rect 1758 113 1764 114
rect 1758 109 1759 113
rect 1763 109 1764 113
rect 1758 108 1764 109
rect 1814 113 1820 114
rect 1814 109 1815 113
rect 1819 109 1820 113
rect 1840 112 1842 162
rect 1936 139 1938 178
rect 2032 139 2034 178
rect 2128 139 2130 178
rect 2216 139 2218 178
rect 1871 138 1875 139
rect 1871 133 1875 134
rect 1927 138 1931 139
rect 1927 133 1931 134
rect 1935 138 1939 139
rect 1935 133 1939 134
rect 1983 138 1987 139
rect 1983 133 1987 134
rect 2031 138 2035 139
rect 2031 133 2035 134
rect 2039 138 2043 139
rect 2039 133 2043 134
rect 2095 138 2099 139
rect 2095 133 2099 134
rect 2127 138 2131 139
rect 2127 133 2131 134
rect 2159 138 2163 139
rect 2159 133 2163 134
rect 2215 138 2219 139
rect 2215 133 2219 134
rect 2223 138 2227 139
rect 2232 136 2234 178
rect 2304 139 2306 178
rect 2344 160 2346 234
rect 2375 210 2379 211
rect 2375 205 2379 206
rect 2374 204 2380 205
rect 2374 200 2375 204
rect 2379 200 2380 204
rect 2374 199 2380 200
rect 2416 184 2418 274
rect 2440 267 2442 290
rect 2439 266 2443 267
rect 2439 261 2443 262
rect 2455 266 2459 267
rect 2455 261 2459 262
rect 2456 242 2458 261
rect 2464 256 2466 290
rect 2504 267 2506 291
rect 2503 266 2507 267
rect 2503 261 2507 262
rect 2462 255 2468 256
rect 2462 251 2463 255
rect 2467 251 2468 255
rect 2462 250 2468 251
rect 2454 241 2460 242
rect 2504 241 2506 261
rect 2454 237 2455 241
rect 2459 237 2460 241
rect 2502 240 2508 241
rect 2454 236 2460 237
rect 2470 239 2476 240
rect 2470 235 2471 239
rect 2475 235 2476 239
rect 2502 236 2503 240
rect 2507 236 2508 240
rect 2502 235 2508 236
rect 2470 234 2476 235
rect 2438 220 2444 221
rect 2438 216 2439 220
rect 2443 216 2444 220
rect 2438 215 2444 216
rect 2440 211 2442 215
rect 2439 210 2443 211
rect 2439 205 2443 206
rect 2438 204 2444 205
rect 2438 200 2439 204
rect 2443 200 2444 204
rect 2438 199 2444 200
rect 2390 183 2396 184
rect 2390 179 2391 183
rect 2395 179 2396 183
rect 2390 178 2396 179
rect 2414 183 2420 184
rect 2414 179 2415 183
rect 2419 179 2420 183
rect 2414 178 2420 179
rect 2454 183 2460 184
rect 2454 179 2455 183
rect 2459 179 2460 183
rect 2454 178 2460 179
rect 2462 183 2468 184
rect 2462 179 2463 183
rect 2467 179 2468 183
rect 2462 178 2468 179
rect 2354 167 2360 168
rect 2354 163 2355 167
rect 2359 163 2360 167
rect 2354 162 2360 163
rect 2342 159 2348 160
rect 2342 155 2343 159
rect 2347 155 2348 159
rect 2342 154 2348 155
rect 2287 138 2291 139
rect 2223 133 2227 134
rect 2230 135 2236 136
rect 1872 114 1874 133
rect 1928 114 1930 133
rect 1984 114 1986 133
rect 2040 114 2042 133
rect 2096 114 2098 133
rect 2160 114 2162 133
rect 2224 114 2226 133
rect 2230 131 2231 135
rect 2235 131 2236 135
rect 2287 133 2291 134
rect 2303 138 2307 139
rect 2303 133 2307 134
rect 2343 138 2347 139
rect 2343 133 2347 134
rect 2230 130 2236 131
rect 2288 114 2290 133
rect 2344 114 2346 133
rect 1870 113 1876 114
rect 1814 108 1820 109
rect 1838 111 1844 112
rect 1326 107 1332 108
rect 1838 107 1839 111
rect 1843 107 1844 111
rect 1870 109 1871 113
rect 1875 109 1876 113
rect 1870 108 1876 109
rect 1926 113 1932 114
rect 1926 109 1927 113
rect 1931 109 1932 113
rect 1926 108 1932 109
rect 1982 113 1988 114
rect 1982 109 1983 113
rect 1987 109 1988 113
rect 1982 108 1988 109
rect 2038 113 2044 114
rect 2038 109 2039 113
rect 2043 109 2044 113
rect 2038 108 2044 109
rect 2094 113 2100 114
rect 2094 109 2095 113
rect 2099 109 2100 113
rect 2094 108 2100 109
rect 2158 113 2164 114
rect 2158 109 2159 113
rect 2163 109 2164 113
rect 2158 108 2164 109
rect 2222 113 2228 114
rect 2222 109 2223 113
rect 2227 109 2228 113
rect 2222 108 2228 109
rect 2286 113 2292 114
rect 2286 109 2287 113
rect 2291 109 2292 113
rect 2286 108 2292 109
rect 2342 113 2348 114
rect 2342 109 2343 113
rect 2347 109 2348 113
rect 2356 112 2358 162
rect 2392 139 2394 178
rect 2456 139 2458 178
rect 2391 138 2395 139
rect 2391 133 2395 134
rect 2399 138 2403 139
rect 2399 133 2403 134
rect 2455 138 2459 139
rect 2455 133 2459 134
rect 2400 114 2402 133
rect 2456 114 2458 133
rect 2464 128 2466 178
rect 2472 168 2474 234
rect 2502 223 2508 224
rect 2502 219 2503 223
rect 2507 219 2508 223
rect 2502 218 2508 219
rect 2504 211 2506 218
rect 2503 210 2507 211
rect 2503 205 2507 206
rect 2504 202 2506 205
rect 2502 201 2508 202
rect 2502 197 2503 201
rect 2507 197 2508 201
rect 2502 196 2508 197
rect 2502 184 2508 185
rect 2502 180 2503 184
rect 2507 180 2508 184
rect 2502 179 2508 180
rect 2470 167 2476 168
rect 2470 163 2471 167
rect 2475 163 2476 167
rect 2470 162 2476 163
rect 2504 139 2506 179
rect 2503 138 2507 139
rect 2503 133 2507 134
rect 2462 127 2468 128
rect 2462 123 2463 127
rect 2467 123 2468 127
rect 2462 122 2468 123
rect 2398 113 2404 114
rect 2342 108 2348 109
rect 2354 111 2360 112
rect 1218 106 1224 107
rect 1838 106 1844 107
rect 2354 107 2355 111
rect 2359 107 2360 111
rect 2398 109 2399 113
rect 2403 109 2404 113
rect 2398 108 2404 109
rect 2454 113 2460 114
rect 2504 113 2506 133
rect 2454 109 2455 113
rect 2459 109 2460 113
rect 2454 108 2460 109
rect 2502 112 2508 113
rect 2502 108 2503 112
rect 2507 108 2508 112
rect 2502 107 2508 108
rect 2354 106 2360 107
rect 110 95 116 96
rect 110 91 111 95
rect 115 91 116 95
rect 1286 95 1292 96
rect 110 90 116 91
rect 134 92 140 93
rect 112 87 114 90
rect 134 88 135 92
rect 139 88 140 92
rect 134 87 140 88
rect 190 92 196 93
rect 190 88 191 92
rect 195 88 196 92
rect 190 87 196 88
rect 246 92 252 93
rect 246 88 247 92
rect 251 88 252 92
rect 246 87 252 88
rect 302 92 308 93
rect 302 88 303 92
rect 307 88 308 92
rect 302 87 308 88
rect 358 92 364 93
rect 358 88 359 92
rect 363 88 364 92
rect 358 87 364 88
rect 414 92 420 93
rect 414 88 415 92
rect 419 88 420 92
rect 414 87 420 88
rect 470 92 476 93
rect 470 88 471 92
rect 475 88 476 92
rect 470 87 476 88
rect 534 92 540 93
rect 534 88 535 92
rect 539 88 540 92
rect 534 87 540 88
rect 606 92 612 93
rect 606 88 607 92
rect 611 88 612 92
rect 606 87 612 88
rect 670 92 676 93
rect 670 88 671 92
rect 675 88 676 92
rect 670 87 676 88
rect 734 92 740 93
rect 734 88 735 92
rect 739 88 740 92
rect 734 87 740 88
rect 798 92 804 93
rect 798 88 799 92
rect 803 88 804 92
rect 798 87 804 88
rect 862 92 868 93
rect 862 88 863 92
rect 867 88 868 92
rect 862 87 868 88
rect 926 92 932 93
rect 926 88 927 92
rect 931 88 932 92
rect 926 87 932 88
rect 990 92 996 93
rect 990 88 991 92
rect 995 88 996 92
rect 990 87 996 88
rect 1054 92 1060 93
rect 1054 88 1055 92
rect 1059 88 1060 92
rect 1054 87 1060 88
rect 1118 92 1124 93
rect 1118 88 1119 92
rect 1123 88 1124 92
rect 1118 87 1124 88
rect 1182 92 1188 93
rect 1182 88 1183 92
rect 1187 88 1188 92
rect 1286 91 1287 95
rect 1291 91 1292 95
rect 1286 90 1292 91
rect 1326 95 1332 96
rect 1326 91 1327 95
rect 1331 91 1332 95
rect 2502 95 2508 96
rect 1326 90 1332 91
rect 1350 92 1356 93
rect 1182 87 1188 88
rect 1288 87 1290 90
rect 1328 87 1330 90
rect 1350 88 1351 92
rect 1355 88 1356 92
rect 1350 87 1356 88
rect 1406 92 1412 93
rect 1406 88 1407 92
rect 1411 88 1412 92
rect 1406 87 1412 88
rect 1462 92 1468 93
rect 1462 88 1463 92
rect 1467 88 1468 92
rect 1462 87 1468 88
rect 1518 92 1524 93
rect 1518 88 1519 92
rect 1523 88 1524 92
rect 1518 87 1524 88
rect 1574 92 1580 93
rect 1574 88 1575 92
rect 1579 88 1580 92
rect 1574 87 1580 88
rect 1630 92 1636 93
rect 1630 88 1631 92
rect 1635 88 1636 92
rect 1630 87 1636 88
rect 1686 92 1692 93
rect 1686 88 1687 92
rect 1691 88 1692 92
rect 1686 87 1692 88
rect 1742 92 1748 93
rect 1742 88 1743 92
rect 1747 88 1748 92
rect 1742 87 1748 88
rect 1798 92 1804 93
rect 1798 88 1799 92
rect 1803 88 1804 92
rect 1798 87 1804 88
rect 1854 92 1860 93
rect 1854 88 1855 92
rect 1859 88 1860 92
rect 1854 87 1860 88
rect 1910 92 1916 93
rect 1910 88 1911 92
rect 1915 88 1916 92
rect 1910 87 1916 88
rect 1966 92 1972 93
rect 1966 88 1967 92
rect 1971 88 1972 92
rect 1966 87 1972 88
rect 2022 92 2028 93
rect 2022 88 2023 92
rect 2027 88 2028 92
rect 2022 87 2028 88
rect 2078 92 2084 93
rect 2078 88 2079 92
rect 2083 88 2084 92
rect 2078 87 2084 88
rect 2142 92 2148 93
rect 2142 88 2143 92
rect 2147 88 2148 92
rect 2142 87 2148 88
rect 2206 92 2212 93
rect 2206 88 2207 92
rect 2211 88 2212 92
rect 2206 87 2212 88
rect 2270 92 2276 93
rect 2270 88 2271 92
rect 2275 88 2276 92
rect 2270 87 2276 88
rect 2326 92 2332 93
rect 2326 88 2327 92
rect 2331 88 2332 92
rect 2326 87 2332 88
rect 2382 92 2388 93
rect 2382 88 2383 92
rect 2387 88 2388 92
rect 2382 87 2388 88
rect 2438 92 2444 93
rect 2438 88 2439 92
rect 2443 88 2444 92
rect 2502 91 2503 95
rect 2507 91 2508 95
rect 2502 90 2508 91
rect 2438 87 2444 88
rect 2504 87 2506 90
rect 111 86 115 87
rect 111 81 115 82
rect 135 86 139 87
rect 135 81 139 82
rect 191 86 195 87
rect 191 81 195 82
rect 247 86 251 87
rect 247 81 251 82
rect 303 86 307 87
rect 303 81 307 82
rect 359 86 363 87
rect 359 81 363 82
rect 415 86 419 87
rect 415 81 419 82
rect 471 86 475 87
rect 471 81 475 82
rect 535 86 539 87
rect 535 81 539 82
rect 607 86 611 87
rect 607 81 611 82
rect 671 86 675 87
rect 671 81 675 82
rect 735 86 739 87
rect 735 81 739 82
rect 799 86 803 87
rect 799 81 803 82
rect 863 86 867 87
rect 863 81 867 82
rect 927 86 931 87
rect 927 81 931 82
rect 991 86 995 87
rect 991 81 995 82
rect 1055 86 1059 87
rect 1055 81 1059 82
rect 1119 86 1123 87
rect 1119 81 1123 82
rect 1183 86 1187 87
rect 1183 81 1187 82
rect 1287 86 1291 87
rect 1287 81 1291 82
rect 1327 86 1331 87
rect 1327 81 1331 82
rect 1351 86 1355 87
rect 1351 81 1355 82
rect 1407 86 1411 87
rect 1407 81 1411 82
rect 1463 86 1467 87
rect 1463 81 1467 82
rect 1519 86 1523 87
rect 1519 81 1523 82
rect 1575 86 1579 87
rect 1575 81 1579 82
rect 1631 86 1635 87
rect 1631 81 1635 82
rect 1687 86 1691 87
rect 1687 81 1691 82
rect 1743 86 1747 87
rect 1743 81 1747 82
rect 1799 86 1803 87
rect 1799 81 1803 82
rect 1855 86 1859 87
rect 1855 81 1859 82
rect 1911 86 1915 87
rect 1911 81 1915 82
rect 1967 86 1971 87
rect 1967 81 1971 82
rect 2023 86 2027 87
rect 2023 81 2027 82
rect 2079 86 2083 87
rect 2079 81 2083 82
rect 2143 86 2147 87
rect 2143 81 2147 82
rect 2207 86 2211 87
rect 2207 81 2211 82
rect 2271 86 2275 87
rect 2271 81 2275 82
rect 2327 86 2331 87
rect 2327 81 2331 82
rect 2383 86 2387 87
rect 2383 81 2387 82
rect 2439 86 2443 87
rect 2439 81 2443 82
rect 2503 86 2507 87
rect 2503 81 2507 82
<< m4c >>
rect 111 2578 115 2582
rect 719 2578 723 2582
rect 775 2578 779 2582
rect 831 2578 835 2582
rect 887 2578 891 2582
rect 943 2578 947 2582
rect 1287 2578 1291 2582
rect 1327 2554 1331 2558
rect 1399 2554 1403 2558
rect 1455 2554 1459 2558
rect 1511 2554 1515 2558
rect 1567 2554 1571 2558
rect 1623 2554 1627 2558
rect 1679 2554 1683 2558
rect 111 2526 115 2530
rect 167 2526 171 2530
rect 223 2526 227 2530
rect 279 2526 283 2530
rect 343 2526 347 2530
rect 407 2526 411 2530
rect 479 2526 483 2530
rect 559 2526 563 2530
rect 639 2526 643 2530
rect 703 2526 707 2530
rect 719 2526 723 2530
rect 759 2526 763 2530
rect 799 2526 803 2530
rect 815 2526 819 2530
rect 871 2526 875 2530
rect 879 2526 883 2530
rect 927 2526 931 2530
rect 111 2474 115 2478
rect 183 2474 187 2478
rect 239 2474 243 2478
rect 247 2474 251 2478
rect 295 2474 299 2478
rect 327 2474 331 2478
rect 359 2474 363 2478
rect 415 2474 419 2478
rect 423 2474 427 2478
rect 495 2474 499 2478
rect 503 2474 507 2478
rect 575 2474 579 2478
rect 599 2474 603 2478
rect 1735 2554 1739 2558
rect 1791 2554 1795 2558
rect 1847 2554 1851 2558
rect 1903 2554 1907 2558
rect 1959 2554 1963 2558
rect 2015 2554 2019 2558
rect 2071 2554 2075 2558
rect 2127 2554 2131 2558
rect 2183 2554 2187 2558
rect 2503 2554 2507 2558
rect 959 2526 963 2530
rect 1039 2526 1043 2530
rect 1287 2526 1291 2530
rect 655 2474 659 2478
rect 695 2474 699 2478
rect 735 2474 739 2478
rect 791 2474 795 2478
rect 815 2474 819 2478
rect 879 2474 883 2478
rect 895 2474 899 2478
rect 967 2474 971 2478
rect 975 2474 979 2478
rect 1055 2474 1059 2478
rect 1063 2474 1067 2478
rect 1327 2494 1331 2498
rect 1351 2494 1355 2498
rect 1383 2494 1387 2498
rect 1423 2494 1427 2498
rect 1439 2494 1443 2498
rect 1495 2494 1499 2498
rect 1511 2494 1515 2498
rect 1551 2494 1555 2498
rect 1599 2494 1603 2498
rect 1607 2494 1611 2498
rect 1663 2494 1667 2498
rect 1687 2494 1691 2498
rect 111 2418 115 2422
rect 151 2418 155 2422
rect 167 2418 171 2422
rect 231 2418 235 2422
rect 311 2418 315 2422
rect 319 2418 323 2422
rect 399 2418 403 2422
rect 415 2418 419 2422
rect 487 2418 491 2422
rect 519 2418 523 2422
rect 583 2418 587 2422
rect 623 2418 627 2422
rect 679 2418 683 2422
rect 727 2418 731 2422
rect 1159 2474 1163 2478
rect 1287 2474 1291 2478
rect 1719 2494 1723 2498
rect 1775 2494 1779 2498
rect 1831 2494 1835 2498
rect 775 2418 779 2422
rect 831 2418 835 2422
rect 863 2418 867 2422
rect 935 2418 939 2422
rect 951 2418 955 2422
rect 1039 2418 1043 2422
rect 1047 2418 1051 2422
rect 1143 2418 1147 2422
rect 1151 2418 1155 2422
rect 111 2366 115 2370
rect 167 2366 171 2370
rect 175 2366 179 2370
rect 247 2366 251 2370
rect 279 2366 283 2370
rect 335 2366 339 2370
rect 391 2366 395 2370
rect 431 2366 435 2370
rect 503 2366 507 2370
rect 535 2366 539 2370
rect 623 2366 627 2370
rect 639 2366 643 2370
rect 743 2366 747 2370
rect 847 2366 851 2370
rect 871 2366 875 2370
rect 951 2366 955 2370
rect 999 2366 1003 2370
rect 1055 2366 1059 2370
rect 1127 2366 1131 2370
rect 111 2310 115 2314
rect 159 2310 163 2314
rect 207 2310 211 2314
rect 263 2310 267 2314
rect 287 2310 291 2314
rect 375 2310 379 2314
rect 471 2310 475 2314
rect 487 2310 491 2314
rect 111 2254 115 2258
rect 223 2254 227 2258
rect 263 2254 267 2258
rect 303 2254 307 2258
rect 319 2254 323 2258
rect 383 2254 387 2258
rect 391 2254 395 2258
rect 447 2254 451 2258
rect 487 2254 491 2258
rect 559 2310 563 2314
rect 607 2310 611 2314
rect 647 2310 651 2314
rect 727 2310 731 2314
rect 735 2310 739 2314
rect 1167 2366 1171 2370
rect 1327 2434 1331 2438
rect 1367 2434 1371 2438
rect 1439 2434 1443 2438
rect 1527 2434 1531 2438
rect 1543 2434 1547 2438
rect 1615 2434 1619 2438
rect 1639 2434 1643 2438
rect 1287 2418 1291 2422
rect 1327 2374 1331 2378
rect 1351 2374 1355 2378
rect 1287 2366 1291 2370
rect 1863 2494 1867 2498
rect 1887 2494 1891 2498
rect 1943 2494 1947 2498
rect 1951 2494 1955 2498
rect 1999 2494 2003 2498
rect 2039 2494 2043 2498
rect 2055 2494 2059 2498
rect 2111 2494 2115 2498
rect 2127 2494 2131 2498
rect 2167 2494 2171 2498
rect 2503 2494 2507 2498
rect 1703 2434 1707 2438
rect 1735 2434 1739 2438
rect 1791 2434 1795 2438
rect 1823 2434 1827 2438
rect 1879 2434 1883 2438
rect 1911 2434 1915 2438
rect 1967 2434 1971 2438
rect 2007 2434 2011 2438
rect 2055 2434 2059 2438
rect 2103 2434 2107 2438
rect 2143 2434 2147 2438
rect 2503 2434 2507 2438
rect 1407 2374 1411 2378
rect 1423 2374 1427 2378
rect 1495 2374 1499 2378
rect 1527 2374 1531 2378
rect 1583 2374 1587 2378
rect 1623 2374 1627 2378
rect 1671 2374 1675 2378
rect 1719 2374 1723 2378
rect 1751 2374 1755 2378
rect 815 2310 819 2314
rect 855 2310 859 2314
rect 903 2310 907 2314
rect 983 2310 987 2314
rect 991 2310 995 2314
rect 503 2254 507 2258
rect 559 2254 563 2258
rect 575 2254 579 2258
rect 615 2254 619 2258
rect 663 2254 667 2258
rect 671 2254 675 2258
rect 727 2254 731 2258
rect 751 2254 755 2258
rect 791 2254 795 2258
rect 831 2254 835 2258
rect 855 2254 859 2258
rect 919 2254 923 2258
rect 1327 2318 1331 2322
rect 1367 2318 1371 2322
rect 1423 2318 1427 2322
rect 1455 2318 1459 2322
rect 1511 2318 1515 2322
rect 1543 2318 1547 2322
rect 1079 2310 1083 2314
rect 1111 2310 1115 2314
rect 1287 2310 1291 2314
rect 1807 2374 1811 2378
rect 1831 2374 1835 2378
rect 1895 2374 1899 2378
rect 1919 2374 1923 2378
rect 1991 2374 1995 2378
rect 2007 2374 2011 2378
rect 2087 2374 2091 2378
rect 2095 2374 2099 2378
rect 2503 2374 2507 2378
rect 1599 2318 1603 2322
rect 1639 2318 1643 2322
rect 1687 2318 1691 2322
rect 1735 2318 1739 2322
rect 1767 2318 1771 2322
rect 1831 2318 1835 2322
rect 1847 2318 1851 2322
rect 1927 2318 1931 2322
rect 1935 2318 1939 2322
rect 2015 2318 2019 2322
rect 2023 2318 2027 2322
rect 2111 2318 2115 2322
rect 2207 2318 2211 2322
rect 2503 2318 2507 2322
rect 1327 2266 1331 2270
rect 1351 2266 1355 2270
rect 1439 2266 1443 2270
rect 1455 2266 1459 2270
rect 1527 2266 1531 2270
rect 1543 2266 1547 2270
rect 1623 2266 1627 2270
rect 1639 2266 1643 2270
rect 1719 2266 1723 2270
rect 1735 2266 1739 2270
rect 1815 2266 1819 2270
rect 1839 2266 1843 2270
rect 1911 2266 1915 2270
rect 983 2254 987 2258
rect 1007 2254 1011 2258
rect 1047 2254 1051 2258
rect 1095 2254 1099 2258
rect 1111 2254 1115 2258
rect 1287 2254 1291 2258
rect 1935 2266 1939 2270
rect 1999 2266 2003 2270
rect 2031 2266 2035 2270
rect 2095 2266 2099 2270
rect 2119 2266 2123 2270
rect 2191 2266 2195 2270
rect 2215 2266 2219 2270
rect 1327 2210 1331 2214
rect 1471 2210 1475 2214
rect 1559 2210 1563 2214
rect 1567 2210 1571 2214
rect 111 2198 115 2202
rect 247 2198 251 2202
rect 303 2198 307 2202
rect 335 2198 339 2202
rect 367 2198 371 2202
rect 391 2198 395 2202
rect 431 2198 435 2202
rect 447 2198 451 2202
rect 487 2198 491 2202
rect 503 2198 507 2202
rect 543 2198 547 2202
rect 559 2198 563 2202
rect 599 2198 603 2202
rect 655 2198 659 2202
rect 711 2198 715 2202
rect 775 2198 779 2202
rect 839 2198 843 2202
rect 903 2198 907 2202
rect 967 2198 971 2202
rect 1031 2198 1035 2202
rect 1095 2198 1099 2202
rect 1287 2198 1291 2202
rect 2311 2266 2315 2270
rect 2503 2266 2507 2270
rect 1623 2210 1627 2214
rect 1655 2210 1659 2214
rect 1679 2210 1683 2214
rect 1743 2210 1747 2214
rect 1751 2210 1755 2214
rect 1807 2210 1811 2214
rect 1855 2210 1859 2214
rect 1871 2210 1875 2214
rect 111 2146 115 2150
rect 351 2146 355 2150
rect 407 2146 411 2150
rect 415 2146 419 2150
rect 463 2146 467 2150
rect 511 2146 515 2150
rect 519 2146 523 2150
rect 575 2146 579 2150
rect 607 2146 611 2150
rect 711 2146 715 2150
rect 815 2146 819 2150
rect 927 2146 931 2150
rect 1039 2146 1043 2150
rect 1151 2146 1155 2150
rect 1239 2146 1243 2150
rect 1287 2146 1291 2150
rect 1327 2146 1331 2150
rect 1551 2146 1555 2150
rect 1607 2146 1611 2150
rect 1663 2146 1667 2150
rect 1719 2146 1723 2150
rect 1727 2146 1731 2150
rect 1791 2146 1795 2150
rect 111 2094 115 2098
rect 375 2094 379 2098
rect 399 2094 403 2098
rect 447 2094 451 2098
rect 495 2094 499 2098
rect 519 2094 523 2098
rect 591 2094 595 2098
rect 599 2094 603 2098
rect 679 2094 683 2098
rect 695 2094 699 2098
rect 759 2094 763 2098
rect 799 2094 803 2098
rect 111 2038 115 2042
rect 295 2038 299 2042
rect 375 2038 379 2042
rect 391 2038 395 2042
rect 831 2094 835 2098
rect 903 2094 907 2098
rect 911 2094 915 2098
rect 967 2094 971 2098
rect 1023 2094 1027 2098
rect 1031 2094 1035 2098
rect 1103 2094 1107 2098
rect 1927 2210 1931 2214
rect 1951 2210 1955 2214
rect 1983 2210 1987 2214
rect 2039 2210 2043 2214
rect 2047 2210 2051 2214
rect 2095 2210 2099 2214
rect 2135 2210 2139 2214
rect 2159 2210 2163 2214
rect 2223 2210 2227 2214
rect 2231 2210 2235 2214
rect 2287 2210 2291 2214
rect 2327 2210 2331 2214
rect 2343 2210 2347 2214
rect 2399 2210 2403 2214
rect 2455 2210 2459 2214
rect 2503 2210 2507 2214
rect 1855 2146 1859 2150
rect 1871 2146 1875 2150
rect 1911 2146 1915 2150
rect 1967 2146 1971 2150
rect 2023 2146 2027 2150
rect 2079 2146 2083 2150
rect 2143 2146 2147 2150
rect 2199 2146 2203 2150
rect 2207 2146 2211 2150
rect 2271 2146 2275 2150
rect 2327 2146 2331 2150
rect 2383 2146 2387 2150
rect 2439 2146 2443 2150
rect 1135 2094 1139 2098
rect 1167 2094 1171 2098
rect 1223 2094 1227 2098
rect 463 2038 467 2042
rect 535 2038 539 2042
rect 551 2038 555 2042
rect 615 2038 619 2042
rect 639 2038 643 2042
rect 695 2038 699 2042
rect 719 2038 723 2042
rect 775 2038 779 2042
rect 799 2038 803 2042
rect 847 2038 851 2042
rect 887 2038 891 2042
rect 919 2038 923 2042
rect 975 2038 979 2042
rect 983 2038 987 2042
rect 1047 2038 1051 2042
rect 1063 2038 1067 2042
rect 111 1982 115 1986
rect 135 1982 139 1986
rect 207 1982 211 1986
rect 279 1982 283 1986
rect 287 1982 291 1986
rect 359 1982 363 1986
rect 383 1982 387 1986
rect 111 1922 115 1926
rect 151 1922 155 1926
rect 223 1922 227 1926
rect 239 1922 243 1926
rect 303 1922 307 1926
rect 447 1982 451 1986
rect 487 1982 491 1986
rect 535 1982 539 1986
rect 591 1982 595 1986
rect 623 1982 627 1986
rect 695 1982 699 1986
rect 703 1982 707 1986
rect 1287 2094 1291 2098
rect 1327 2082 1331 2086
rect 1367 2082 1371 2086
rect 1423 2082 1427 2086
rect 1503 2082 1507 2086
rect 1591 2082 1595 2086
rect 1679 2082 1683 2086
rect 1735 2082 1739 2086
rect 1783 2082 1787 2086
rect 1807 2082 1811 2086
rect 1887 2082 1891 2086
rect 1895 2082 1899 2086
rect 1983 2082 1987 2086
rect 2023 2082 2027 2086
rect 2095 2082 2099 2086
rect 2167 2082 2171 2086
rect 2215 2082 2219 2086
rect 2319 2082 2323 2086
rect 1119 2038 1123 2042
rect 1183 2038 1187 2042
rect 1239 2038 1243 2042
rect 1287 2038 1291 2042
rect 1327 2030 1331 2034
rect 1351 2030 1355 2034
rect 1407 2030 1411 2034
rect 1423 2030 1427 2034
rect 1487 2030 1491 2034
rect 1519 2030 1523 2034
rect 1575 2030 1579 2034
rect 1615 2030 1619 2034
rect 1663 2030 1667 2034
rect 783 1982 787 1986
rect 799 1982 803 1986
rect 871 1982 875 1986
rect 903 1982 907 1986
rect 959 1982 963 1986
rect 1015 1982 1019 1986
rect 1047 1982 1051 1986
rect 1287 1982 1291 1986
rect 1719 2030 1723 2034
rect 1767 2030 1771 2034
rect 1823 2030 1827 2034
rect 2343 2082 2347 2086
rect 2455 2082 2459 2086
rect 2503 2146 2507 2150
rect 2503 2082 2507 2086
rect 1879 2030 1883 2034
rect 1935 2030 1939 2034
rect 2007 2030 2011 2034
rect 2055 2030 2059 2034
rect 2151 2030 2155 2034
rect 2183 2030 2187 2034
rect 2303 2030 2307 2034
rect 2319 2030 2323 2034
rect 2439 2030 2443 2034
rect 1327 1974 1331 1978
rect 1367 1974 1371 1978
rect 1439 1974 1443 1978
rect 1455 1974 1459 1978
rect 1535 1974 1539 1978
rect 1543 1974 1547 1978
rect 1631 1974 1635 1978
rect 1639 1974 1643 1978
rect 1735 1974 1739 1978
rect 375 1922 379 1926
rect 399 1922 403 1926
rect 503 1922 507 1926
rect 527 1922 531 1926
rect 607 1922 611 1926
rect 687 1922 691 1926
rect 711 1922 715 1926
rect 815 1922 819 1926
rect 863 1922 867 1926
rect 1839 1974 1843 1978
rect 1943 1974 1947 1978
rect 1951 1974 1955 1978
rect 2047 1974 2051 1978
rect 2071 1974 2075 1978
rect 2151 1974 2155 1978
rect 2199 1974 2203 1978
rect 2255 1974 2259 1978
rect 919 1922 923 1926
rect 1031 1922 1035 1926
rect 1039 1922 1043 1926
rect 1287 1922 1291 1926
rect 111 1870 115 1874
rect 135 1870 139 1874
rect 191 1870 195 1874
rect 111 1810 115 1814
rect 151 1810 155 1814
rect 223 1870 227 1874
rect 263 1870 267 1874
rect 335 1870 339 1874
rect 359 1870 363 1874
rect 407 1870 411 1874
rect 479 1870 483 1874
rect 511 1870 515 1874
rect 551 1870 555 1874
rect 615 1870 619 1874
rect 671 1870 675 1874
rect 679 1870 683 1874
rect 743 1870 747 1874
rect 815 1870 819 1874
rect 847 1870 851 1874
rect 887 1870 891 1874
rect 959 1870 963 1874
rect 1023 1870 1027 1874
rect 1039 1870 1043 1874
rect 1327 1918 1331 1922
rect 1439 1918 1443 1922
rect 1527 1918 1531 1922
rect 1615 1918 1619 1922
rect 1623 1918 1627 1922
rect 1711 1918 1715 1922
rect 1719 1918 1723 1922
rect 1815 1918 1819 1922
rect 1823 1918 1827 1922
rect 1287 1870 1291 1874
rect 1919 1918 1923 1922
rect 1927 1918 1931 1922
rect 2015 1918 2019 1922
rect 2031 1918 2035 1922
rect 2111 1918 2115 1922
rect 2135 1918 2139 1922
rect 2199 1918 2203 1922
rect 2239 1918 2243 1922
rect 2335 1974 2339 1978
rect 2367 1974 2371 1978
rect 2455 1974 2459 1978
rect 2503 2030 2507 2034
rect 2503 1974 2507 1978
rect 2287 1918 2291 1922
rect 2351 1918 2355 1922
rect 2375 1918 2379 1922
rect 2439 1918 2443 1922
rect 1327 1866 1331 1870
rect 1535 1866 1539 1870
rect 1543 1866 1547 1870
rect 1607 1866 1611 1870
rect 1631 1866 1635 1870
rect 1687 1866 1691 1870
rect 1727 1866 1731 1870
rect 1783 1866 1787 1870
rect 1831 1866 1835 1870
rect 1879 1866 1883 1870
rect 1935 1866 1939 1870
rect 207 1810 211 1814
rect 231 1810 235 1814
rect 279 1810 283 1814
rect 335 1810 339 1814
rect 351 1810 355 1814
rect 423 1810 427 1814
rect 439 1810 443 1814
rect 495 1810 499 1814
rect 535 1810 539 1814
rect 567 1810 571 1814
rect 631 1810 635 1814
rect 111 1754 115 1758
rect 135 1754 139 1758
rect 215 1754 219 1758
rect 239 1754 243 1758
rect 319 1754 323 1758
rect 351 1754 355 1758
rect 111 1698 115 1702
rect 151 1698 155 1702
rect 423 1754 427 1758
rect 463 1754 467 1758
rect 695 1810 699 1814
rect 719 1810 723 1814
rect 759 1810 763 1814
rect 799 1810 803 1814
rect 831 1810 835 1814
rect 879 1810 883 1814
rect 903 1810 907 1814
rect 959 1810 963 1814
rect 975 1810 979 1814
rect 1039 1810 1043 1814
rect 1055 1810 1059 1814
rect 2503 1918 2507 1922
rect 1983 1866 1987 1870
rect 2031 1866 2035 1870
rect 2079 1866 2083 1870
rect 2127 1866 2131 1870
rect 2175 1866 2179 1870
rect 2215 1866 2219 1870
rect 2271 1866 2275 1870
rect 2303 1866 2307 1870
rect 2367 1866 2371 1870
rect 2391 1866 2395 1870
rect 2455 1866 2459 1870
rect 1119 1810 1123 1814
rect 1287 1810 1291 1814
rect 1327 1810 1331 1814
rect 1463 1810 1467 1814
rect 1519 1810 1523 1814
rect 1559 1810 1563 1814
rect 1591 1810 1595 1814
rect 1663 1810 1667 1814
rect 1671 1810 1675 1814
rect 519 1754 523 1758
rect 575 1754 579 1758
rect 615 1754 619 1758
rect 679 1754 683 1758
rect 703 1754 707 1758
rect 783 1754 787 1758
rect 863 1754 867 1758
rect 887 1754 891 1758
rect 943 1754 947 1758
rect 991 1754 995 1758
rect 191 1698 195 1702
rect 255 1698 259 1702
rect 271 1698 275 1702
rect 351 1698 355 1702
rect 367 1698 371 1702
rect 439 1698 443 1702
rect 479 1698 483 1702
rect 535 1698 539 1702
rect 591 1698 595 1702
rect 639 1698 643 1702
rect 111 1646 115 1650
rect 175 1646 179 1650
rect 215 1646 219 1650
rect 255 1646 259 1650
rect 271 1646 275 1650
rect 335 1646 339 1650
rect 111 1594 115 1598
rect 231 1594 235 1598
rect 287 1594 291 1598
rect 407 1646 411 1650
rect 423 1646 427 1650
rect 695 1698 699 1702
rect 1023 1754 1027 1758
rect 1103 1754 1107 1758
rect 1287 1754 1291 1758
rect 1327 1754 1331 1758
rect 1375 1754 1379 1758
rect 1471 1754 1475 1758
rect 1479 1754 1483 1758
rect 1767 1810 1771 1814
rect 1863 1810 1867 1814
rect 1879 1810 1883 1814
rect 1967 1810 1971 1814
rect 1983 1810 1987 1814
rect 2063 1810 2067 1814
rect 2087 1810 2091 1814
rect 2159 1810 2163 1814
rect 2183 1810 2187 1814
rect 2255 1810 2259 1814
rect 2271 1810 2275 1814
rect 2351 1810 2355 1814
rect 2367 1810 2371 1814
rect 2439 1810 2443 1814
rect 2167 1792 2171 1796
rect 2403 1792 2407 1796
rect 1567 1754 1571 1758
rect 1575 1754 1579 1758
rect 1671 1754 1675 1758
rect 1679 1754 1683 1758
rect 1775 1754 1779 1758
rect 1783 1754 1787 1758
rect 1887 1754 1891 1758
rect 1895 1754 1899 1758
rect 1999 1754 2003 1758
rect 2103 1754 2107 1758
rect 2111 1754 2115 1758
rect 2199 1754 2203 1758
rect 2231 1754 2235 1758
rect 2287 1754 2291 1758
rect 2351 1754 2355 1758
rect 743 1698 747 1702
rect 799 1698 803 1702
rect 847 1698 851 1702
rect 903 1698 907 1702
rect 951 1698 955 1702
rect 1007 1698 1011 1702
rect 1063 1698 1067 1702
rect 1119 1698 1123 1702
rect 1175 1698 1179 1702
rect 479 1646 483 1650
rect 519 1646 523 1650
rect 559 1646 563 1650
rect 623 1646 627 1650
rect 647 1646 651 1650
rect 727 1646 731 1650
rect 743 1646 747 1650
rect 831 1646 835 1650
rect 839 1646 843 1650
rect 935 1646 939 1650
rect 943 1646 947 1650
rect 351 1594 355 1598
rect 423 1594 427 1598
rect 495 1594 499 1598
rect 503 1594 507 1598
rect 575 1594 579 1598
rect 599 1594 603 1598
rect 663 1594 667 1598
rect 703 1594 707 1598
rect 759 1594 763 1598
rect 1047 1646 1051 1650
rect 1055 1646 1059 1650
rect 1287 1698 1291 1702
rect 1327 1702 1331 1706
rect 1351 1702 1355 1706
rect 1359 1702 1363 1706
rect 1431 1702 1435 1706
rect 1159 1646 1163 1650
rect 1175 1646 1179 1650
rect 1287 1646 1291 1650
rect 1327 1642 1331 1646
rect 1367 1642 1371 1646
rect 1383 1664 1387 1668
rect 1455 1702 1459 1706
rect 1535 1702 1539 1706
rect 1551 1702 1555 1706
rect 1647 1702 1651 1706
rect 1655 1702 1659 1706
rect 1759 1702 1763 1706
rect 1871 1702 1875 1706
rect 1879 1702 1883 1706
rect 1983 1702 1987 1706
rect 2015 1702 2019 1706
rect 2095 1702 2099 1706
rect 2159 1702 2163 1706
rect 2215 1702 2219 1706
rect 2311 1702 2315 1706
rect 2335 1702 2339 1706
rect 2383 1754 2387 1758
rect 2455 1754 2459 1758
rect 2503 1866 2507 1870
rect 2503 1810 2507 1814
rect 2503 1754 2507 1758
rect 2439 1702 2443 1706
rect 1671 1664 1675 1668
rect 1431 1642 1435 1646
rect 1447 1642 1451 1646
rect 1519 1642 1523 1646
rect 1551 1642 1555 1646
rect 1599 1642 1603 1646
rect 1663 1642 1667 1646
rect 1679 1642 1683 1646
rect 1751 1642 1755 1646
rect 1775 1642 1779 1646
rect 1839 1642 1843 1646
rect 1895 1642 1899 1646
rect 1935 1642 1939 1646
rect 2031 1642 2035 1646
rect 2055 1642 2059 1646
rect 2175 1642 2179 1646
rect 2183 1642 2187 1646
rect 2327 1642 2331 1646
rect 815 1594 819 1598
rect 855 1594 859 1598
rect 935 1594 939 1598
rect 959 1594 963 1598
rect 1063 1594 1067 1598
rect 1071 1594 1075 1598
rect 1191 1594 1195 1598
rect 619 1568 623 1572
rect 955 1571 959 1572
rect 955 1568 959 1571
rect 111 1534 115 1538
rect 271 1534 275 1538
rect 335 1534 339 1538
rect 407 1534 411 1538
rect 471 1534 475 1538
rect 487 1534 491 1538
rect 551 1534 555 1538
rect 583 1534 587 1538
rect 639 1534 643 1538
rect 687 1534 691 1538
rect 735 1534 739 1538
rect 111 1482 115 1486
rect 375 1482 379 1486
rect 463 1482 467 1486
rect 487 1482 491 1486
rect 559 1482 563 1486
rect 567 1482 571 1486
rect 655 1482 659 1486
rect 799 1534 803 1538
rect 839 1534 843 1538
rect 919 1534 923 1538
rect 951 1534 955 1538
rect 1287 1594 1291 1598
rect 1327 1586 1331 1590
rect 1351 1586 1355 1590
rect 1415 1586 1419 1590
rect 1423 1586 1427 1590
rect 1503 1586 1507 1590
rect 1527 1586 1531 1590
rect 1047 1534 1051 1538
rect 1063 1534 1067 1538
rect 1175 1534 1179 1538
rect 1287 1534 1291 1538
rect 1327 1534 1331 1538
rect 1367 1534 1371 1538
rect 1583 1586 1587 1590
rect 1647 1586 1651 1590
rect 1663 1586 1667 1590
rect 1735 1586 1739 1590
rect 1783 1586 1787 1590
rect 1823 1586 1827 1590
rect 1919 1586 1923 1590
rect 1935 1586 1939 1590
rect 2039 1586 2043 1590
rect 2103 1586 2107 1590
rect 2455 1642 2459 1646
rect 2503 1702 2507 1706
rect 2503 1642 2507 1646
rect 2167 1586 2171 1590
rect 2279 1586 2283 1590
rect 2311 1586 2315 1590
rect 2439 1586 2443 1590
rect 1439 1534 1443 1538
rect 1543 1534 1547 1538
rect 1647 1534 1651 1538
rect 1663 1534 1667 1538
rect 1751 1534 1755 1538
rect 1799 1534 1803 1538
rect 1855 1534 1859 1538
rect 751 1482 755 1486
rect 855 1482 859 1486
rect 959 1482 963 1486
rect 967 1482 971 1486
rect 1063 1482 1067 1486
rect 1079 1482 1083 1486
rect 1167 1482 1171 1486
rect 1191 1482 1195 1486
rect 111 1430 115 1434
rect 231 1430 235 1434
rect 319 1430 323 1434
rect 359 1430 363 1434
rect 415 1430 419 1434
rect 447 1430 451 1434
rect 511 1430 515 1434
rect 543 1430 547 1434
rect 615 1430 619 1434
rect 111 1378 115 1382
rect 151 1378 155 1382
rect 215 1378 219 1382
rect 247 1378 251 1382
rect 311 1378 315 1382
rect 335 1378 339 1382
rect 407 1378 411 1382
rect 431 1378 435 1382
rect 639 1430 643 1434
rect 711 1430 715 1434
rect 735 1430 739 1434
rect 807 1430 811 1434
rect 839 1430 843 1434
rect 895 1430 899 1434
rect 943 1430 947 1434
rect 991 1430 995 1434
rect 1047 1430 1051 1434
rect 1087 1430 1091 1434
rect 1287 1482 1291 1486
rect 1327 1478 1331 1482
rect 1351 1478 1355 1482
rect 1423 1478 1427 1482
rect 1151 1430 1155 1434
rect 1287 1430 1291 1434
rect 1327 1422 1331 1426
rect 1367 1422 1371 1426
rect 1519 1478 1523 1482
rect 1527 1478 1531 1482
rect 1615 1478 1619 1482
rect 1631 1478 1635 1482
rect 1951 1534 1955 1538
rect 1959 1534 1963 1538
rect 2055 1534 2059 1538
rect 2119 1534 2123 1538
rect 2151 1534 2155 1538
rect 2247 1534 2251 1538
rect 2503 1586 2507 1590
rect 2295 1534 2299 1538
rect 2343 1534 2347 1538
rect 2439 1534 2443 1538
rect 2455 1534 2459 1538
rect 1711 1478 1715 1482
rect 1735 1478 1739 1482
rect 1815 1478 1819 1482
rect 1839 1478 1843 1482
rect 1927 1478 1931 1482
rect 1943 1478 1947 1482
rect 2039 1478 2043 1482
rect 2047 1478 2051 1482
rect 2135 1478 2139 1482
rect 1423 1422 1427 1426
rect 1439 1422 1443 1426
rect 1503 1422 1507 1426
rect 1535 1422 1539 1426
rect 1591 1422 1595 1426
rect 1631 1422 1635 1426
rect 1679 1422 1683 1426
rect 511 1378 515 1382
rect 527 1378 531 1382
rect 607 1378 611 1382
rect 631 1378 635 1382
rect 703 1378 707 1382
rect 727 1378 731 1382
rect 799 1378 803 1382
rect 823 1378 827 1382
rect 895 1378 899 1382
rect 911 1378 915 1382
rect 999 1378 1003 1382
rect 1007 1378 1011 1382
rect 111 1326 115 1330
rect 135 1326 139 1330
rect 199 1326 203 1330
rect 215 1326 219 1330
rect 295 1326 299 1330
rect 319 1326 323 1330
rect 391 1326 395 1330
rect 415 1326 419 1330
rect 495 1326 499 1330
rect 511 1326 515 1330
rect 591 1326 595 1330
rect 599 1326 603 1330
rect 687 1326 691 1330
rect 783 1326 787 1330
rect 879 1326 883 1330
rect 1103 1378 1107 1382
rect 1287 1378 1291 1382
rect 1327 1366 1331 1370
rect 1351 1366 1355 1370
rect 983 1326 987 1330
rect 1287 1326 1291 1330
rect 1407 1366 1411 1370
rect 1479 1366 1483 1370
rect 1487 1366 1491 1370
rect 1567 1366 1571 1370
rect 1575 1366 1579 1370
rect 1727 1422 1731 1426
rect 1775 1422 1779 1426
rect 1831 1422 1835 1426
rect 2175 1478 2179 1482
rect 2231 1478 2235 1482
rect 2303 1478 2307 1482
rect 2327 1478 2331 1482
rect 2503 1534 2507 1538
rect 2423 1478 2427 1482
rect 2439 1478 2443 1482
rect 1879 1422 1883 1426
rect 1943 1422 1947 1426
rect 1991 1422 1995 1426
rect 2063 1422 2067 1426
rect 2111 1422 2115 1426
rect 2191 1422 2195 1426
rect 2231 1422 2235 1426
rect 2503 1478 2507 1482
rect 2319 1422 2323 1426
rect 2351 1422 2355 1426
rect 2455 1422 2459 1426
rect 1655 1366 1659 1370
rect 1663 1366 1667 1370
rect 1751 1366 1755 1370
rect 1759 1366 1763 1370
rect 1855 1366 1859 1370
rect 1863 1366 1867 1370
rect 1967 1366 1971 1370
rect 1975 1366 1979 1370
rect 2079 1366 2083 1370
rect 2095 1366 2099 1370
rect 1327 1306 1331 1310
rect 1367 1306 1371 1310
rect 1423 1306 1427 1310
rect 1495 1306 1499 1310
rect 1519 1306 1523 1310
rect 111 1274 115 1278
rect 151 1274 155 1278
rect 191 1274 195 1278
rect 231 1274 235 1278
rect 247 1274 251 1278
rect 303 1274 307 1278
rect 335 1274 339 1278
rect 367 1274 371 1278
rect 431 1274 435 1278
rect 439 1274 443 1278
rect 527 1274 531 1278
rect 615 1274 619 1278
rect 639 1274 643 1278
rect 703 1274 707 1278
rect 775 1274 779 1278
rect 799 1274 803 1278
rect 895 1274 899 1278
rect 927 1274 931 1278
rect 1095 1274 1099 1278
rect 111 1222 115 1226
rect 175 1222 179 1226
rect 231 1222 235 1226
rect 287 1222 291 1226
rect 351 1222 355 1226
rect 407 1222 411 1226
rect 423 1222 427 1226
rect 463 1222 467 1226
rect 511 1222 515 1226
rect 519 1222 523 1226
rect 575 1222 579 1226
rect 623 1222 627 1226
rect 631 1222 635 1226
rect 1239 1274 1243 1278
rect 1583 1306 1587 1310
rect 1615 1306 1619 1310
rect 1671 1306 1675 1310
rect 1719 1306 1723 1310
rect 2199 1366 2203 1370
rect 2215 1366 2219 1370
rect 2327 1366 2331 1370
rect 2335 1366 2339 1370
rect 2503 1422 2507 1426
rect 2439 1366 2443 1370
rect 1767 1306 1771 1310
rect 1823 1306 1827 1310
rect 1871 1306 1875 1310
rect 1919 1306 1923 1310
rect 1983 1306 1987 1310
rect 2015 1306 2019 1310
rect 2095 1306 2099 1310
rect 2103 1306 2107 1310
rect 2183 1306 2187 1310
rect 2215 1306 2219 1310
rect 1287 1274 1291 1278
rect 687 1222 691 1226
rect 743 1222 747 1226
rect 759 1222 763 1226
rect 799 1222 803 1226
rect 855 1222 859 1226
rect 911 1222 915 1226
rect 1079 1222 1083 1226
rect 1223 1222 1227 1226
rect 1327 1238 1331 1242
rect 1351 1238 1355 1242
rect 1407 1238 1411 1242
rect 1447 1238 1451 1242
rect 1503 1238 1507 1242
rect 1575 1238 1579 1242
rect 1599 1238 1603 1242
rect 1695 1238 1699 1242
rect 1703 1238 1707 1242
rect 1807 1238 1811 1242
rect 1815 1238 1819 1242
rect 1287 1222 1291 1226
rect 2255 1306 2259 1310
rect 2327 1306 2331 1310
rect 2343 1306 2347 1310
rect 2503 1366 2507 1370
rect 2399 1306 2403 1310
rect 2455 1306 2459 1310
rect 2503 1306 2507 1310
rect 1903 1238 1907 1242
rect 1927 1238 1931 1242
rect 1999 1238 2003 1242
rect 2031 1238 2035 1242
rect 2087 1238 2091 1242
rect 2127 1238 2131 1242
rect 2167 1238 2171 1242
rect 2215 1238 2219 1242
rect 2239 1238 2243 1242
rect 111 1166 115 1170
rect 367 1166 371 1170
rect 423 1166 427 1170
rect 479 1166 483 1170
rect 535 1166 539 1170
rect 591 1166 595 1170
rect 647 1166 651 1170
rect 703 1166 707 1170
rect 759 1166 763 1170
rect 815 1166 819 1170
rect 871 1166 875 1170
rect 111 1110 115 1114
rect 223 1110 227 1114
rect 311 1110 315 1114
rect 399 1110 403 1114
rect 407 1110 411 1114
rect 463 1110 467 1114
rect 495 1110 499 1114
rect 519 1110 523 1114
rect 575 1110 579 1114
rect 111 1054 115 1058
rect 151 1054 155 1058
rect 207 1054 211 1058
rect 239 1054 243 1058
rect 303 1054 307 1058
rect 327 1054 331 1058
rect 415 1054 419 1058
rect 591 1110 595 1114
rect 631 1110 635 1114
rect 679 1110 683 1114
rect 687 1110 691 1114
rect 743 1110 747 1114
rect 767 1110 771 1114
rect 799 1110 803 1114
rect 847 1110 851 1114
rect 855 1110 859 1114
rect 1327 1186 1331 1190
rect 1367 1186 1371 1190
rect 1463 1186 1467 1190
rect 1471 1186 1475 1190
rect 1951 1200 1955 1204
rect 2295 1238 2299 1242
rect 2311 1238 2315 1242
rect 2375 1238 2379 1242
rect 2383 1238 2387 1242
rect 2439 1238 2443 1242
rect 2263 1200 2267 1204
rect 927 1166 931 1170
rect 983 1166 987 1170
rect 1287 1166 1291 1170
rect 1591 1186 1595 1190
rect 1599 1186 1603 1190
rect 1711 1186 1715 1190
rect 1735 1186 1739 1190
rect 1831 1186 1835 1190
rect 1863 1186 1867 1190
rect 1943 1186 1947 1190
rect 1983 1186 1987 1190
rect 2047 1186 2051 1190
rect 2087 1186 2091 1190
rect 2143 1186 2147 1190
rect 2191 1186 2195 1190
rect 1327 1130 1331 1134
rect 1351 1130 1355 1134
rect 1367 1130 1371 1134
rect 1447 1130 1451 1134
rect 1455 1130 1459 1134
rect 1535 1130 1539 1134
rect 1583 1130 1587 1134
rect 911 1110 915 1114
rect 927 1110 931 1114
rect 967 1110 971 1114
rect 1015 1110 1019 1114
rect 1103 1110 1107 1114
rect 1287 1110 1291 1114
rect 511 1054 515 1058
rect 535 1054 539 1058
rect 607 1054 611 1058
rect 655 1054 659 1058
rect 695 1054 699 1058
rect 767 1054 771 1058
rect 783 1054 787 1058
rect 863 1054 867 1058
rect 879 1054 883 1058
rect 943 1054 947 1058
rect 983 1054 987 1058
rect 775 1032 779 1036
rect 111 998 115 1002
rect 135 998 139 1002
rect 191 998 195 1002
rect 215 998 219 1002
rect 287 998 291 1002
rect 327 998 331 1002
rect 111 946 115 950
rect 151 946 155 950
rect 399 998 403 1002
rect 439 998 443 1002
rect 519 998 523 1002
rect 551 998 555 1002
rect 639 998 643 1002
rect 663 998 667 1002
rect 751 998 755 1002
rect 759 998 763 1002
rect 1327 1070 1331 1074
rect 1383 1070 1387 1074
rect 1031 1054 1035 1058
rect 1095 1054 1099 1058
rect 1119 1054 1123 1058
rect 1207 1054 1211 1058
rect 1287 1054 1291 1058
rect 1227 1032 1231 1036
rect 1631 1130 1635 1134
rect 1719 1130 1723 1134
rect 1807 1130 1811 1134
rect 1847 1130 1851 1134
rect 2231 1186 2235 1190
rect 2287 1186 2291 1190
rect 2311 1186 2315 1190
rect 2383 1186 2387 1190
rect 2391 1186 2395 1190
rect 2503 1238 2507 1242
rect 2455 1186 2459 1190
rect 1895 1130 1899 1134
rect 1967 1130 1971 1134
rect 1983 1130 1987 1134
rect 2071 1130 2075 1134
rect 2159 1130 2163 1134
rect 1431 1070 1435 1074
rect 1463 1070 1467 1074
rect 1495 1070 1499 1074
rect 1551 1070 1555 1074
rect 1567 1070 1571 1074
rect 1639 1070 1643 1074
rect 1647 1070 1651 1074
rect 1703 1070 1707 1074
rect 1735 1070 1739 1074
rect 1767 1070 1771 1074
rect 1327 1010 1331 1014
rect 1415 1010 1419 1014
rect 1479 1010 1483 1014
rect 1511 1010 1515 1014
rect 1551 1010 1555 1014
rect 1567 1010 1571 1014
rect 1623 1010 1627 1014
rect 847 998 851 1002
rect 863 998 867 1002
rect 935 998 939 1002
rect 967 998 971 1002
rect 1015 998 1019 1002
rect 1079 998 1083 1002
rect 1087 998 1091 1002
rect 1167 998 1171 1002
rect 1191 998 1195 1002
rect 1223 998 1227 1002
rect 1287 998 1291 1002
rect 207 946 211 950
rect 231 946 235 950
rect 295 946 299 950
rect 343 946 347 950
rect 399 946 403 950
rect 455 946 459 950
rect 511 946 515 950
rect 567 946 571 950
rect 623 946 627 950
rect 679 946 683 950
rect 735 946 739 950
rect 111 890 115 894
rect 135 890 139 894
rect 191 890 195 894
rect 247 890 251 894
rect 279 890 283 894
rect 343 890 347 894
rect 383 890 387 894
rect 775 946 779 950
rect 831 946 835 950
rect 439 890 443 894
rect 495 890 499 894
rect 543 890 547 894
rect 607 890 611 894
rect 647 890 651 894
rect 719 890 723 894
rect 743 890 747 894
rect 863 946 867 950
rect 927 946 931 950
rect 951 946 955 950
rect 1015 946 1019 950
rect 1031 946 1035 950
rect 1095 946 1099 950
rect 1103 946 1107 950
rect 1175 946 1179 950
rect 1183 946 1187 950
rect 1239 946 1243 950
rect 1287 946 1291 950
rect 815 890 819 894
rect 839 890 843 894
rect 911 890 915 894
rect 927 890 931 894
rect 999 890 1003 894
rect 1007 890 1011 894
rect 1079 890 1083 894
rect 1087 890 1091 894
rect 111 834 115 838
rect 239 834 243 838
rect 263 834 267 838
rect 303 834 307 838
rect 359 834 363 838
rect 383 834 387 838
rect 455 834 459 838
rect 463 834 467 838
rect 551 834 555 838
rect 559 834 563 838
rect 639 834 643 838
rect 663 834 667 838
rect 1159 890 1163 894
rect 1167 890 1171 894
rect 1223 890 1227 894
rect 1327 942 1331 946
rect 1367 942 1371 946
rect 1439 942 1443 946
rect 1527 942 1531 946
rect 1679 1010 1683 1014
rect 1687 1010 1691 1014
rect 1959 1091 1963 1092
rect 1959 1088 1963 1091
rect 1823 1070 1827 1074
rect 1839 1070 1843 1074
rect 1911 1070 1915 1074
rect 1919 1070 1923 1074
rect 1999 1070 2003 1074
rect 2007 1070 2011 1074
rect 2087 1070 2091 1074
rect 2111 1070 2115 1074
rect 2175 1130 2179 1134
rect 2255 1130 2259 1134
rect 2271 1130 2275 1134
rect 2359 1130 2363 1134
rect 2367 1130 2371 1134
rect 2439 1130 2443 1134
rect 2383 1088 2387 1092
rect 2175 1070 2179 1074
rect 2231 1070 2235 1074
rect 2271 1070 2275 1074
rect 2351 1070 2355 1074
rect 2375 1070 2379 1074
rect 2455 1070 2459 1074
rect 2503 1186 2507 1190
rect 1735 1010 1739 1014
rect 1751 1010 1755 1014
rect 1807 1010 1811 1014
rect 1823 1010 1827 1014
rect 1887 1010 1891 1014
rect 1903 1010 1907 1014
rect 1983 1010 1987 1014
rect 1991 1010 1995 1014
rect 2095 1010 2099 1014
rect 2215 1010 2219 1014
rect 2335 1010 2339 1014
rect 2439 1010 2443 1014
rect 1583 942 1587 946
rect 1615 942 1619 946
rect 1639 942 1643 946
rect 1695 942 1699 946
rect 1751 942 1755 946
rect 1791 942 1795 946
rect 1823 942 1827 946
rect 1895 942 1899 946
rect 1903 942 1907 946
rect 1999 942 2003 946
rect 2015 942 2019 946
rect 2111 942 2115 946
rect 2151 942 2155 946
rect 2231 942 2235 946
rect 2295 942 2299 946
rect 2351 942 2355 946
rect 1287 890 1291 894
rect 1327 882 1331 886
rect 1351 882 1355 886
rect 1423 882 1427 886
rect 1487 882 1491 886
rect 1511 882 1515 886
rect 1559 882 1563 886
rect 727 834 731 838
rect 759 834 763 838
rect 807 834 811 838
rect 855 834 859 838
rect 895 834 899 838
rect 943 834 947 838
rect 983 834 987 838
rect 1023 834 1027 838
rect 1071 834 1075 838
rect 1103 834 1107 838
rect 111 778 115 782
rect 151 778 155 782
rect 223 778 227 782
rect 247 778 251 782
rect 287 778 291 782
rect 343 778 347 782
rect 111 722 115 726
rect 167 722 171 726
rect 175 722 179 726
rect 1183 834 1187 838
rect 1239 834 1243 838
rect 1287 834 1291 838
rect 1327 822 1331 826
rect 1439 822 1443 826
rect 1503 822 1507 826
rect 1511 822 1515 826
rect 1599 882 1603 886
rect 1623 882 1627 886
rect 1679 882 1683 886
rect 1687 882 1691 886
rect 1751 882 1755 886
rect 1775 882 1779 886
rect 1815 882 1819 886
rect 1879 882 1883 886
rect 1887 882 1891 886
rect 1975 882 1979 886
rect 1999 882 2003 886
rect 2079 882 2083 886
rect 2135 882 2139 886
rect 2199 882 2203 886
rect 2279 882 2283 886
rect 1575 822 1579 826
rect 1591 822 1595 826
rect 1639 822 1643 826
rect 1671 822 1675 826
rect 1703 822 1707 826
rect 1759 822 1763 826
rect 1767 822 1771 826
rect 367 778 371 782
rect 439 778 443 782
rect 447 778 451 782
rect 527 778 531 782
rect 535 778 539 782
rect 607 778 611 782
rect 623 778 627 782
rect 679 778 683 782
rect 711 778 715 782
rect 751 778 755 782
rect 791 778 795 782
rect 823 778 827 782
rect 879 778 883 782
rect 895 778 899 782
rect 967 778 971 782
rect 975 778 979 782
rect 1055 778 1059 782
rect 1287 778 1291 782
rect 1327 766 1331 770
rect 1351 766 1355 770
rect 1423 766 1427 770
rect 1447 766 1451 770
rect 1495 766 1499 770
rect 1567 766 1571 770
rect 1575 766 1579 770
rect 263 722 267 726
rect 343 722 347 726
rect 359 722 363 726
rect 111 670 115 674
rect 159 670 163 674
rect 215 670 219 674
rect 247 670 251 674
rect 295 670 299 674
rect 423 722 427 726
rect 455 722 459 726
rect 503 722 507 726
rect 543 722 547 726
rect 575 722 579 726
rect 623 722 627 726
rect 639 722 643 726
rect 695 722 699 726
rect 703 722 707 726
rect 767 722 771 726
rect 839 722 843 726
rect 911 722 915 726
rect 327 670 331 674
rect 375 670 379 674
rect 407 670 411 674
rect 455 670 459 674
rect 487 670 491 674
rect 527 670 531 674
rect 111 614 115 618
rect 207 614 211 618
rect 231 614 235 618
rect 303 614 307 618
rect 311 614 315 618
rect 391 614 395 618
rect 407 614 411 618
rect 111 558 115 562
rect 175 558 179 562
rect 191 558 195 562
rect 271 558 275 562
rect 287 558 291 562
rect 375 558 379 562
rect 391 558 395 562
rect 471 614 475 618
rect 559 670 563 674
rect 591 670 595 674
rect 623 670 627 674
rect 991 722 995 726
rect 1287 722 1291 726
rect 1327 710 1331 714
rect 1367 710 1371 714
rect 1655 766 1659 770
rect 1687 766 1691 770
rect 1839 848 1843 852
rect 2319 882 2323 886
rect 2303 848 2307 852
rect 1831 822 1835 826
rect 1847 822 1851 826
rect 1903 822 1907 826
rect 1935 822 1939 826
rect 1991 822 1995 826
rect 2023 822 2027 826
rect 2095 822 2099 826
rect 2111 822 2115 826
rect 2199 822 2203 826
rect 2215 822 2219 826
rect 2287 822 2291 826
rect 2335 822 2339 826
rect 2383 822 2387 826
rect 1743 766 1747 770
rect 1807 766 1811 770
rect 1831 766 1835 770
rect 1919 766 1923 770
rect 1927 766 1931 770
rect 2007 766 2011 770
rect 2039 766 2043 770
rect 2095 766 2099 770
rect 2143 766 2147 770
rect 2183 766 2187 770
rect 2247 766 2251 770
rect 2271 766 2275 770
rect 1431 710 1435 714
rect 1463 710 1467 714
rect 1535 710 1539 714
rect 1583 710 1587 714
rect 1639 710 1643 714
rect 1703 710 1707 714
rect 1751 710 1755 714
rect 1823 710 1827 714
rect 1863 710 1867 714
rect 655 670 659 674
rect 687 670 691 674
rect 719 670 723 674
rect 751 670 755 674
rect 783 670 787 674
rect 823 670 827 674
rect 847 670 851 674
rect 895 670 899 674
rect 919 670 923 674
rect 1287 670 1291 674
rect 1327 650 1331 654
rect 1351 650 1355 654
rect 1415 650 1419 654
rect 1479 650 1483 654
rect 1519 650 1523 654
rect 1559 650 1563 654
rect 1623 650 1627 654
rect 1647 650 1651 654
rect 503 614 507 618
rect 543 614 547 618
rect 599 614 603 618
rect 607 614 611 618
rect 671 614 675 618
rect 687 614 691 618
rect 735 614 739 618
rect 767 614 771 618
rect 799 614 803 618
rect 847 614 851 618
rect 863 614 867 618
rect 927 614 931 618
rect 935 614 939 618
rect 1007 614 1011 618
rect 1087 614 1091 618
rect 487 558 491 562
rect 583 558 587 562
rect 591 558 595 562
rect 111 502 115 506
rect 151 502 155 506
rect 191 502 195 506
rect 247 502 251 506
rect 287 502 291 506
rect 367 502 371 506
rect 391 502 395 506
rect 487 502 491 506
rect 111 446 115 450
rect 135 446 139 450
rect 191 446 195 450
rect 231 446 235 450
rect 247 446 251 450
rect 303 446 307 450
rect 671 558 675 562
rect 695 558 699 562
rect 751 558 755 562
rect 791 558 795 562
rect 831 558 835 562
rect 879 558 883 562
rect 911 558 915 562
rect 967 558 971 562
rect 991 558 995 562
rect 1287 614 1291 618
rect 1735 650 1739 654
rect 1975 720 1979 724
rect 1943 710 1947 714
rect 1967 710 1971 714
rect 2351 766 2355 770
rect 2367 766 2371 770
rect 2423 882 2427 886
rect 2439 942 2443 946
rect 2503 1130 2507 1134
rect 2503 1070 2507 1074
rect 2503 1010 2507 1014
rect 2455 942 2459 946
rect 2503 942 2507 946
rect 2439 882 2443 886
rect 2503 882 2507 886
rect 2455 822 2459 826
rect 2503 822 2507 826
rect 2439 766 2443 770
rect 2271 720 2275 724
rect 2055 710 2059 714
rect 2063 710 2067 714
rect 2151 710 2155 714
rect 2159 710 2163 714
rect 2231 710 2235 714
rect 2263 710 2267 714
rect 2311 710 2315 714
rect 2367 710 2371 714
rect 2391 710 2395 714
rect 1831 650 1835 654
rect 1847 650 1851 654
rect 1919 650 1923 654
rect 1951 650 1955 654
rect 2007 650 2011 654
rect 2047 650 2051 654
rect 2087 650 2091 654
rect 2135 650 2139 654
rect 2167 650 2171 654
rect 2215 650 2219 654
rect 2239 650 2243 654
rect 1327 594 1331 598
rect 1455 594 1459 598
rect 1495 594 1499 598
rect 1559 594 1563 598
rect 1575 594 1579 598
rect 1663 594 1667 598
rect 1671 594 1675 598
rect 1751 594 1755 598
rect 1775 594 1779 598
rect 1847 594 1851 598
rect 1879 594 1883 598
rect 1055 558 1059 562
rect 1071 558 1075 562
rect 1151 558 1155 562
rect 1287 558 1291 562
rect 1327 538 1331 542
rect 1367 538 1371 542
rect 1439 538 1443 542
rect 1447 538 1451 542
rect 503 502 507 506
rect 607 502 611 506
rect 615 502 619 506
rect 711 502 715 506
rect 735 502 739 506
rect 807 502 811 506
rect 847 502 851 506
rect 895 502 899 506
rect 951 502 955 506
rect 983 502 987 506
rect 1055 502 1059 506
rect 1071 502 1075 506
rect 1159 502 1163 506
rect 1167 502 1171 506
rect 1239 502 1243 506
rect 1287 502 1291 506
rect 351 446 355 450
rect 383 446 387 450
rect 471 446 475 450
rect 567 446 571 450
rect 599 446 603 450
rect 111 386 115 390
rect 151 386 155 390
rect 207 386 211 390
rect 263 386 267 390
rect 279 386 283 390
rect 319 386 323 390
rect 359 386 363 390
rect 399 386 403 390
rect 431 386 435 390
rect 487 386 491 390
rect 511 386 515 390
rect 111 326 115 330
rect 135 326 139 330
rect 191 326 195 330
rect 199 326 203 330
rect 263 326 267 330
rect 287 326 291 330
rect 343 326 347 330
rect 375 326 379 330
rect 415 326 419 330
rect 455 326 459 330
rect 671 446 675 450
rect 719 446 723 450
rect 783 446 787 450
rect 831 446 835 450
rect 895 446 899 450
rect 935 446 939 450
rect 1007 446 1011 450
rect 1039 446 1043 450
rect 1127 446 1131 450
rect 1143 446 1147 450
rect 1223 446 1227 450
rect 1327 482 1331 486
rect 1367 482 1371 486
rect 1383 482 1387 486
rect 1527 538 1531 542
rect 1543 538 1547 542
rect 1615 538 1619 542
rect 1655 538 1659 542
rect 1711 538 1715 542
rect 1759 538 1763 542
rect 1799 538 1803 542
rect 1935 594 1939 598
rect 1983 594 1987 598
rect 2023 594 2027 598
rect 2087 594 2091 598
rect 2103 594 2107 598
rect 2455 710 2459 714
rect 2503 766 2507 770
rect 2503 710 2507 714
rect 2295 650 2299 654
rect 2311 650 2315 654
rect 2375 650 2379 654
rect 2383 650 2387 654
rect 2439 650 2443 654
rect 2183 594 2187 598
rect 2255 594 2259 598
rect 2279 594 2283 598
rect 2327 594 2331 598
rect 2375 594 2379 598
rect 2399 594 2403 598
rect 1863 538 1867 542
rect 1887 538 1891 542
rect 1967 538 1971 542
rect 1975 538 1979 542
rect 2063 538 2067 542
rect 2071 538 2075 542
rect 2151 538 2155 542
rect 1431 482 1435 486
rect 1463 482 1467 486
rect 1519 482 1523 486
rect 1543 482 1547 486
rect 1615 482 1619 486
rect 1631 482 1635 486
rect 1711 482 1715 486
rect 1287 446 1291 450
rect 1327 426 1331 430
rect 1351 426 1355 430
rect 1415 426 1419 430
rect 1423 426 1427 430
rect 1503 426 1507 430
rect 1511 426 1515 430
rect 583 386 587 390
rect 591 386 595 390
rect 671 386 675 390
rect 687 386 691 390
rect 751 386 755 390
rect 799 386 803 390
rect 823 386 827 390
rect 895 386 899 390
rect 911 386 915 390
rect 967 386 971 390
rect 1023 386 1027 390
rect 1039 386 1043 390
rect 1111 386 1115 390
rect 1143 386 1147 390
rect 1183 386 1187 390
rect 1239 386 1243 390
rect 1287 386 1291 390
rect 495 326 499 330
rect 543 326 547 330
rect 575 326 579 330
rect 631 326 635 330
rect 111 266 115 270
rect 151 266 155 270
rect 215 266 219 270
rect 231 266 235 270
rect 303 266 307 270
rect 327 266 331 270
rect 391 266 395 270
rect 423 266 427 270
rect 471 266 475 270
rect 519 266 523 270
rect 655 326 659 330
rect 727 326 731 330
rect 735 326 739 330
rect 807 326 811 330
rect 823 326 827 330
rect 879 326 883 330
rect 927 326 931 330
rect 951 326 955 330
rect 1023 326 1027 330
rect 1031 326 1035 330
rect 2055 496 2059 500
rect 1727 482 1731 486
rect 1815 482 1819 486
rect 1903 482 1907 486
rect 1927 482 1931 486
rect 1991 482 1995 486
rect 2055 482 2059 486
rect 2079 482 2083 486
rect 2167 538 2171 542
rect 2247 538 2251 542
rect 2263 538 2267 542
rect 2343 538 2347 542
rect 2359 538 2363 542
rect 2455 594 2459 598
rect 2503 650 2507 654
rect 2503 594 2507 598
rect 2439 538 2443 542
rect 2271 496 2275 500
rect 2167 482 2171 486
rect 2191 482 2195 486
rect 2263 482 2267 486
rect 2335 482 2339 486
rect 2359 482 2363 486
rect 2455 482 2459 486
rect 2503 538 2507 542
rect 1599 426 1603 430
rect 1679 426 1683 430
rect 1695 426 1699 430
rect 1775 426 1779 430
rect 1799 426 1803 430
rect 1887 426 1891 430
rect 1911 426 1915 430
rect 2015 426 2019 430
rect 1327 370 1331 374
rect 1367 370 1371 374
rect 1439 370 1443 374
rect 1527 370 1531 374
rect 1615 370 1619 374
rect 1679 370 1683 374
rect 1695 370 1699 374
rect 1735 370 1739 374
rect 1095 326 1099 330
rect 1135 326 1139 330
rect 1167 326 1171 330
rect 1223 326 1227 330
rect 559 266 563 270
rect 615 266 619 270
rect 647 266 651 270
rect 711 266 715 270
rect 743 266 747 270
rect 807 266 811 270
rect 839 266 843 270
rect 903 266 907 270
rect 111 206 115 210
rect 135 206 139 210
rect 159 206 163 210
rect 215 206 219 210
rect 239 206 243 210
rect 111 134 115 138
rect 151 134 155 138
rect 175 134 179 138
rect 311 206 315 210
rect 327 206 331 210
rect 407 206 411 210
rect 415 206 419 210
rect 503 206 507 210
rect 511 206 515 210
rect 599 206 603 210
rect 607 206 611 210
rect 943 266 947 270
rect 1287 326 1291 330
rect 1327 318 1331 322
rect 1351 318 1355 322
rect 1431 318 1435 322
rect 1527 318 1531 322
rect 1623 318 1627 322
rect 1663 318 1667 322
rect 1007 266 1011 270
rect 1047 266 1051 270
rect 1111 266 1115 270
rect 1151 266 1155 270
rect 1215 266 1219 270
rect 695 206 699 210
rect 783 206 787 210
rect 791 206 795 210
rect 871 206 875 210
rect 207 134 211 138
rect 255 134 259 138
rect 263 134 267 138
rect 319 134 323 138
rect 343 134 347 138
rect 375 134 379 138
rect 431 134 435 138
rect 487 134 491 138
rect 527 134 531 138
rect 551 134 555 138
rect 623 134 627 138
rect 687 134 691 138
rect 711 134 715 138
rect 887 206 891 210
rect 959 206 963 210
rect 991 206 995 210
rect 1791 370 1795 374
rect 1807 370 1811 374
rect 2039 426 2043 430
rect 2159 426 2163 430
rect 2175 426 2179 430
rect 2311 426 2315 430
rect 2319 426 2323 430
rect 2439 426 2443 430
rect 1903 370 1907 374
rect 2023 370 2027 374
rect 2031 370 2035 374
rect 2159 370 2163 374
rect 2175 370 2179 374
rect 2303 370 2307 374
rect 2327 370 2331 374
rect 2455 370 2459 374
rect 2503 482 2507 486
rect 2503 426 2507 430
rect 2503 370 2507 374
rect 1711 318 1715 322
rect 1719 318 1723 322
rect 1791 318 1795 322
rect 1807 318 1811 322
rect 1887 318 1891 322
rect 1911 318 1915 322
rect 2007 318 2011 322
rect 2023 318 2027 322
rect 2143 318 2147 322
rect 2151 318 2155 322
rect 2287 318 2291 322
rect 1239 266 1243 270
rect 1287 266 1291 270
rect 1327 262 1331 266
rect 1367 262 1371 266
rect 1439 262 1443 266
rect 1447 262 1451 266
rect 1535 262 1539 266
rect 1543 262 1547 266
rect 1631 262 1635 266
rect 1639 262 1643 266
rect 1727 262 1731 266
rect 1047 206 1051 210
rect 1095 206 1099 210
rect 1135 206 1139 210
rect 1199 206 1203 210
rect 1287 206 1291 210
rect 1327 206 1331 210
rect 1351 206 1355 210
rect 1391 206 1395 210
rect 1423 206 1427 210
rect 1495 206 1499 210
rect 1519 206 1523 210
rect 1599 206 1603 210
rect 751 134 755 138
rect 799 134 803 138
rect 815 134 819 138
rect 879 134 883 138
rect 887 134 891 138
rect 943 134 947 138
rect 975 134 979 138
rect 1007 134 1011 138
rect 1063 134 1067 138
rect 1071 134 1075 138
rect 1135 134 1139 138
rect 1151 134 1155 138
rect 1199 134 1203 138
rect 1287 134 1291 138
rect 1327 134 1331 138
rect 1367 134 1371 138
rect 1407 134 1411 138
rect 1615 206 1619 210
rect 1711 206 1715 210
rect 1815 262 1819 266
rect 1823 262 1827 266
rect 1903 262 1907 266
rect 1927 262 1931 266
rect 1999 262 2003 266
rect 2039 262 2043 266
rect 2103 262 2107 266
rect 2167 262 2171 266
rect 2215 262 2219 266
rect 2303 262 2307 266
rect 2423 318 2427 322
rect 2439 318 2443 322
rect 2503 318 2507 322
rect 2335 262 2339 266
rect 1799 206 1803 210
rect 1815 206 1819 210
rect 1887 206 1891 210
rect 1919 206 1923 210
rect 1983 206 1987 210
rect 2015 206 2019 210
rect 2087 206 2091 210
rect 2111 206 2115 210
rect 2199 206 2203 210
rect 2287 206 2291 210
rect 2319 206 2323 210
rect 1423 134 1427 138
rect 1479 134 1483 138
rect 1511 134 1515 138
rect 1535 134 1539 138
rect 1591 134 1595 138
rect 1615 134 1619 138
rect 1647 134 1651 138
rect 1703 134 1707 138
rect 1727 134 1731 138
rect 1759 134 1763 138
rect 1815 134 1819 138
rect 1831 134 1835 138
rect 1871 134 1875 138
rect 1927 134 1931 138
rect 1935 134 1939 138
rect 1983 134 1987 138
rect 2031 134 2035 138
rect 2039 134 2043 138
rect 2095 134 2099 138
rect 2127 134 2131 138
rect 2159 134 2163 138
rect 2215 134 2219 138
rect 2223 134 2227 138
rect 2375 206 2379 210
rect 2439 262 2443 266
rect 2455 262 2459 266
rect 2503 262 2507 266
rect 2439 206 2443 210
rect 2287 134 2291 138
rect 2303 134 2307 138
rect 2343 134 2347 138
rect 2391 134 2395 138
rect 2399 134 2403 138
rect 2455 134 2459 138
rect 2503 206 2507 210
rect 2503 134 2507 138
rect 111 82 115 86
rect 135 82 139 86
rect 191 82 195 86
rect 247 82 251 86
rect 303 82 307 86
rect 359 82 363 86
rect 415 82 419 86
rect 471 82 475 86
rect 535 82 539 86
rect 607 82 611 86
rect 671 82 675 86
rect 735 82 739 86
rect 799 82 803 86
rect 863 82 867 86
rect 927 82 931 86
rect 991 82 995 86
rect 1055 82 1059 86
rect 1119 82 1123 86
rect 1183 82 1187 86
rect 1287 82 1291 86
rect 1327 82 1331 86
rect 1351 82 1355 86
rect 1407 82 1411 86
rect 1463 82 1467 86
rect 1519 82 1523 86
rect 1575 82 1579 86
rect 1631 82 1635 86
rect 1687 82 1691 86
rect 1743 82 1747 86
rect 1799 82 1803 86
rect 1855 82 1859 86
rect 1911 82 1915 86
rect 1967 82 1971 86
rect 2023 82 2027 86
rect 2079 82 2083 86
rect 2143 82 2147 86
rect 2207 82 2211 86
rect 2271 82 2275 86
rect 2327 82 2331 86
rect 2383 82 2387 86
rect 2439 82 2443 86
rect 2503 82 2507 86
<< m4 >>
rect 96 2577 97 2583
rect 103 2582 1311 2583
rect 103 2578 111 2582
rect 115 2578 719 2582
rect 723 2578 775 2582
rect 779 2578 831 2582
rect 835 2578 887 2582
rect 891 2578 943 2582
rect 947 2578 1287 2582
rect 1291 2578 1311 2582
rect 103 2577 1311 2578
rect 1317 2577 1318 2583
rect 1310 2553 1311 2559
rect 1317 2558 2539 2559
rect 1317 2554 1327 2558
rect 1331 2554 1399 2558
rect 1403 2554 1455 2558
rect 1459 2554 1511 2558
rect 1515 2554 1567 2558
rect 1571 2554 1623 2558
rect 1627 2554 1679 2558
rect 1683 2554 1735 2558
rect 1739 2554 1791 2558
rect 1795 2554 1847 2558
rect 1851 2554 1903 2558
rect 1907 2554 1959 2558
rect 1963 2554 2015 2558
rect 2019 2554 2071 2558
rect 2075 2554 2127 2558
rect 2131 2554 2183 2558
rect 2187 2554 2503 2558
rect 2507 2554 2539 2558
rect 1317 2553 2539 2554
rect 2545 2553 2546 2559
rect 84 2525 85 2531
rect 91 2530 1299 2531
rect 91 2526 111 2530
rect 115 2526 167 2530
rect 171 2526 223 2530
rect 227 2526 279 2530
rect 283 2526 343 2530
rect 347 2526 407 2530
rect 411 2526 479 2530
rect 483 2526 559 2530
rect 563 2526 639 2530
rect 643 2526 703 2530
rect 707 2526 719 2530
rect 723 2526 759 2530
rect 763 2526 799 2530
rect 803 2526 815 2530
rect 819 2526 871 2530
rect 875 2526 879 2530
rect 883 2526 927 2530
rect 931 2526 959 2530
rect 963 2526 1039 2530
rect 1043 2526 1287 2530
rect 1291 2526 1299 2530
rect 91 2525 1299 2526
rect 1305 2525 1306 2531
rect 1298 2493 1299 2499
rect 1305 2498 2527 2499
rect 1305 2494 1327 2498
rect 1331 2494 1351 2498
rect 1355 2494 1383 2498
rect 1387 2494 1423 2498
rect 1427 2494 1439 2498
rect 1443 2494 1495 2498
rect 1499 2494 1511 2498
rect 1515 2494 1551 2498
rect 1555 2494 1599 2498
rect 1603 2494 1607 2498
rect 1611 2494 1663 2498
rect 1667 2494 1687 2498
rect 1691 2494 1719 2498
rect 1723 2494 1775 2498
rect 1779 2494 1831 2498
rect 1835 2494 1863 2498
rect 1867 2494 1887 2498
rect 1891 2494 1943 2498
rect 1947 2494 1951 2498
rect 1955 2494 1999 2498
rect 2003 2494 2039 2498
rect 2043 2494 2055 2498
rect 2059 2494 2111 2498
rect 2115 2494 2127 2498
rect 2131 2494 2167 2498
rect 2171 2494 2503 2498
rect 2507 2494 2527 2498
rect 1305 2493 2527 2494
rect 2533 2493 2534 2499
rect 96 2473 97 2479
rect 103 2478 1311 2479
rect 103 2474 111 2478
rect 115 2474 183 2478
rect 187 2474 239 2478
rect 243 2474 247 2478
rect 251 2474 295 2478
rect 299 2474 327 2478
rect 331 2474 359 2478
rect 363 2474 415 2478
rect 419 2474 423 2478
rect 427 2474 495 2478
rect 499 2474 503 2478
rect 507 2474 575 2478
rect 579 2474 599 2478
rect 603 2474 655 2478
rect 659 2474 695 2478
rect 699 2474 735 2478
rect 739 2474 791 2478
rect 795 2474 815 2478
rect 819 2474 879 2478
rect 883 2474 895 2478
rect 899 2474 967 2478
rect 971 2474 975 2478
rect 979 2474 1055 2478
rect 1059 2474 1063 2478
rect 1067 2474 1159 2478
rect 1163 2474 1287 2478
rect 1291 2474 1311 2478
rect 103 2473 1311 2474
rect 1317 2473 1318 2479
rect 1310 2433 1311 2439
rect 1317 2438 2539 2439
rect 1317 2434 1327 2438
rect 1331 2434 1367 2438
rect 1371 2434 1439 2438
rect 1443 2434 1527 2438
rect 1531 2434 1543 2438
rect 1547 2434 1615 2438
rect 1619 2434 1639 2438
rect 1643 2434 1703 2438
rect 1707 2434 1735 2438
rect 1739 2434 1791 2438
rect 1795 2434 1823 2438
rect 1827 2434 1879 2438
rect 1883 2434 1911 2438
rect 1915 2434 1967 2438
rect 1971 2434 2007 2438
rect 2011 2434 2055 2438
rect 2059 2434 2103 2438
rect 2107 2434 2143 2438
rect 2147 2434 2503 2438
rect 2507 2434 2539 2438
rect 1317 2433 2539 2434
rect 2545 2433 2546 2439
rect 84 2417 85 2423
rect 91 2422 1299 2423
rect 91 2418 111 2422
rect 115 2418 151 2422
rect 155 2418 167 2422
rect 171 2418 231 2422
rect 235 2418 311 2422
rect 315 2418 319 2422
rect 323 2418 399 2422
rect 403 2418 415 2422
rect 419 2418 487 2422
rect 491 2418 519 2422
rect 523 2418 583 2422
rect 587 2418 623 2422
rect 627 2418 679 2422
rect 683 2418 727 2422
rect 731 2418 775 2422
rect 779 2418 831 2422
rect 835 2418 863 2422
rect 867 2418 935 2422
rect 939 2418 951 2422
rect 955 2418 1039 2422
rect 1043 2418 1047 2422
rect 1051 2418 1143 2422
rect 1147 2418 1151 2422
rect 1155 2418 1287 2422
rect 1291 2418 1299 2422
rect 91 2417 1299 2418
rect 1305 2417 1306 2423
rect 1298 2375 1299 2381
rect 1305 2379 1330 2381
rect 1305 2378 2527 2379
rect 1305 2375 1327 2378
rect 1324 2374 1327 2375
rect 1331 2374 1351 2378
rect 1355 2374 1407 2378
rect 1411 2374 1423 2378
rect 1427 2374 1495 2378
rect 1499 2374 1527 2378
rect 1531 2374 1583 2378
rect 1587 2374 1623 2378
rect 1627 2374 1671 2378
rect 1675 2374 1719 2378
rect 1723 2374 1751 2378
rect 1755 2374 1807 2378
rect 1811 2374 1831 2378
rect 1835 2374 1895 2378
rect 1899 2374 1919 2378
rect 1923 2374 1991 2378
rect 1995 2374 2007 2378
rect 2011 2374 2087 2378
rect 2091 2374 2095 2378
rect 2099 2374 2503 2378
rect 2507 2374 2527 2378
rect 1324 2373 2527 2374
rect 2533 2373 2534 2379
rect 96 2365 97 2371
rect 103 2370 1311 2371
rect 103 2366 111 2370
rect 115 2366 167 2370
rect 171 2366 175 2370
rect 179 2366 247 2370
rect 251 2366 279 2370
rect 283 2366 335 2370
rect 339 2366 391 2370
rect 395 2366 431 2370
rect 435 2366 503 2370
rect 507 2366 535 2370
rect 539 2366 623 2370
rect 627 2366 639 2370
rect 643 2366 743 2370
rect 747 2366 847 2370
rect 851 2366 871 2370
rect 875 2366 951 2370
rect 955 2366 999 2370
rect 1003 2366 1055 2370
rect 1059 2366 1127 2370
rect 1131 2366 1167 2370
rect 1171 2366 1287 2370
rect 1291 2366 1311 2370
rect 103 2365 1311 2366
rect 1317 2365 1318 2371
rect 1310 2317 1311 2323
rect 1317 2322 2539 2323
rect 1317 2318 1327 2322
rect 1331 2318 1367 2322
rect 1371 2318 1423 2322
rect 1427 2318 1455 2322
rect 1459 2318 1511 2322
rect 1515 2318 1543 2322
rect 1547 2318 1599 2322
rect 1603 2318 1639 2322
rect 1643 2318 1687 2322
rect 1691 2318 1735 2322
rect 1739 2318 1767 2322
rect 1771 2318 1831 2322
rect 1835 2318 1847 2322
rect 1851 2318 1927 2322
rect 1931 2318 1935 2322
rect 1939 2318 2015 2322
rect 2019 2318 2023 2322
rect 2027 2318 2111 2322
rect 2115 2318 2207 2322
rect 2211 2318 2503 2322
rect 2507 2318 2539 2322
rect 1317 2317 2539 2318
rect 2545 2317 2546 2323
rect 84 2309 85 2315
rect 91 2314 1299 2315
rect 91 2310 111 2314
rect 115 2310 159 2314
rect 163 2310 207 2314
rect 211 2310 263 2314
rect 267 2310 287 2314
rect 291 2310 375 2314
rect 379 2310 471 2314
rect 475 2310 487 2314
rect 491 2310 559 2314
rect 563 2310 607 2314
rect 611 2310 647 2314
rect 651 2310 727 2314
rect 731 2310 735 2314
rect 739 2310 815 2314
rect 819 2310 855 2314
rect 859 2310 903 2314
rect 907 2310 983 2314
rect 987 2310 991 2314
rect 995 2310 1079 2314
rect 1083 2310 1111 2314
rect 1115 2310 1287 2314
rect 1291 2310 1299 2314
rect 91 2309 1299 2310
rect 1305 2309 1306 2315
rect 1298 2265 1299 2271
rect 1305 2270 2527 2271
rect 1305 2266 1327 2270
rect 1331 2266 1351 2270
rect 1355 2266 1439 2270
rect 1443 2266 1455 2270
rect 1459 2266 1527 2270
rect 1531 2266 1543 2270
rect 1547 2266 1623 2270
rect 1627 2266 1639 2270
rect 1643 2266 1719 2270
rect 1723 2266 1735 2270
rect 1739 2266 1815 2270
rect 1819 2266 1839 2270
rect 1843 2266 1911 2270
rect 1915 2266 1935 2270
rect 1939 2266 1999 2270
rect 2003 2266 2031 2270
rect 2035 2266 2095 2270
rect 2099 2266 2119 2270
rect 2123 2266 2191 2270
rect 2195 2266 2215 2270
rect 2219 2266 2311 2270
rect 2315 2266 2503 2270
rect 2507 2266 2527 2270
rect 1305 2265 2527 2266
rect 2533 2265 2534 2271
rect 96 2253 97 2259
rect 103 2258 1311 2259
rect 103 2254 111 2258
rect 115 2254 223 2258
rect 227 2254 263 2258
rect 267 2254 303 2258
rect 307 2254 319 2258
rect 323 2254 383 2258
rect 387 2254 391 2258
rect 395 2254 447 2258
rect 451 2254 487 2258
rect 491 2254 503 2258
rect 507 2254 559 2258
rect 563 2254 575 2258
rect 579 2254 615 2258
rect 619 2254 663 2258
rect 667 2254 671 2258
rect 675 2254 727 2258
rect 731 2254 751 2258
rect 755 2254 791 2258
rect 795 2254 831 2258
rect 835 2254 855 2258
rect 859 2254 919 2258
rect 923 2254 983 2258
rect 987 2254 1007 2258
rect 1011 2254 1047 2258
rect 1051 2254 1095 2258
rect 1099 2254 1111 2258
rect 1115 2254 1287 2258
rect 1291 2254 1311 2258
rect 103 2253 1311 2254
rect 1317 2253 1318 2259
rect 1310 2209 1311 2215
rect 1317 2214 2539 2215
rect 1317 2210 1327 2214
rect 1331 2210 1471 2214
rect 1475 2210 1559 2214
rect 1563 2210 1567 2214
rect 1571 2210 1623 2214
rect 1627 2210 1655 2214
rect 1659 2210 1679 2214
rect 1683 2210 1743 2214
rect 1747 2210 1751 2214
rect 1755 2210 1807 2214
rect 1811 2210 1855 2214
rect 1859 2210 1871 2214
rect 1875 2210 1927 2214
rect 1931 2210 1951 2214
rect 1955 2210 1983 2214
rect 1987 2210 2039 2214
rect 2043 2210 2047 2214
rect 2051 2210 2095 2214
rect 2099 2210 2135 2214
rect 2139 2210 2159 2214
rect 2163 2210 2223 2214
rect 2227 2210 2231 2214
rect 2235 2210 2287 2214
rect 2291 2210 2327 2214
rect 2331 2210 2343 2214
rect 2347 2210 2399 2214
rect 2403 2210 2455 2214
rect 2459 2210 2503 2214
rect 2507 2210 2539 2214
rect 1317 2209 2539 2210
rect 2545 2209 2546 2215
rect 84 2197 85 2203
rect 91 2202 1299 2203
rect 91 2198 111 2202
rect 115 2198 247 2202
rect 251 2198 303 2202
rect 307 2198 335 2202
rect 339 2198 367 2202
rect 371 2198 391 2202
rect 395 2198 431 2202
rect 435 2198 447 2202
rect 451 2198 487 2202
rect 491 2198 503 2202
rect 507 2198 543 2202
rect 547 2198 559 2202
rect 563 2198 599 2202
rect 603 2198 655 2202
rect 659 2198 711 2202
rect 715 2198 775 2202
rect 779 2198 839 2202
rect 843 2198 903 2202
rect 907 2198 967 2202
rect 971 2198 1031 2202
rect 1035 2198 1095 2202
rect 1099 2198 1287 2202
rect 1291 2198 1299 2202
rect 91 2197 1299 2198
rect 1305 2197 1306 2203
rect 1298 2155 1299 2161
rect 1305 2155 1330 2161
rect 1324 2151 1330 2155
rect 96 2145 97 2151
rect 103 2150 1311 2151
rect 103 2146 111 2150
rect 115 2146 351 2150
rect 355 2146 407 2150
rect 411 2146 415 2150
rect 419 2146 463 2150
rect 467 2146 511 2150
rect 515 2146 519 2150
rect 523 2146 575 2150
rect 579 2146 607 2150
rect 611 2146 711 2150
rect 715 2146 815 2150
rect 819 2146 927 2150
rect 931 2146 1039 2150
rect 1043 2146 1151 2150
rect 1155 2146 1239 2150
rect 1243 2146 1287 2150
rect 1291 2146 1311 2150
rect 103 2145 1311 2146
rect 1317 2145 1318 2151
rect 1324 2150 2527 2151
rect 1324 2146 1327 2150
rect 1331 2146 1551 2150
rect 1555 2146 1607 2150
rect 1611 2146 1663 2150
rect 1667 2146 1719 2150
rect 1723 2146 1727 2150
rect 1731 2146 1791 2150
rect 1795 2146 1855 2150
rect 1859 2146 1871 2150
rect 1875 2146 1911 2150
rect 1915 2146 1967 2150
rect 1971 2146 2023 2150
rect 2027 2146 2079 2150
rect 2083 2146 2143 2150
rect 2147 2146 2199 2150
rect 2203 2146 2207 2150
rect 2211 2146 2271 2150
rect 2275 2146 2327 2150
rect 2331 2146 2383 2150
rect 2387 2146 2439 2150
rect 2443 2146 2503 2150
rect 2507 2146 2527 2150
rect 1324 2145 2527 2146
rect 2533 2145 2534 2151
rect 84 2093 85 2099
rect 91 2098 1299 2099
rect 91 2094 111 2098
rect 115 2094 375 2098
rect 379 2094 399 2098
rect 403 2094 447 2098
rect 451 2094 495 2098
rect 499 2094 519 2098
rect 523 2094 591 2098
rect 595 2094 599 2098
rect 603 2094 679 2098
rect 683 2094 695 2098
rect 699 2094 759 2098
rect 763 2094 799 2098
rect 803 2094 831 2098
rect 835 2094 903 2098
rect 907 2094 911 2098
rect 915 2094 967 2098
rect 971 2094 1023 2098
rect 1027 2094 1031 2098
rect 1035 2094 1103 2098
rect 1107 2094 1135 2098
rect 1139 2094 1167 2098
rect 1171 2094 1223 2098
rect 1227 2094 1287 2098
rect 1291 2094 1299 2098
rect 91 2093 1299 2094
rect 1305 2093 1306 2099
rect 1310 2081 1311 2087
rect 1317 2086 2539 2087
rect 1317 2082 1327 2086
rect 1331 2082 1367 2086
rect 1371 2082 1423 2086
rect 1427 2082 1503 2086
rect 1507 2082 1591 2086
rect 1595 2082 1679 2086
rect 1683 2082 1735 2086
rect 1739 2082 1783 2086
rect 1787 2082 1807 2086
rect 1811 2082 1887 2086
rect 1891 2082 1895 2086
rect 1899 2082 1983 2086
rect 1987 2082 2023 2086
rect 2027 2082 2095 2086
rect 2099 2082 2167 2086
rect 2171 2082 2215 2086
rect 2219 2082 2319 2086
rect 2323 2082 2343 2086
rect 2347 2082 2455 2086
rect 2459 2082 2503 2086
rect 2507 2082 2539 2086
rect 1317 2081 2539 2082
rect 2545 2081 2546 2087
rect 1298 2047 1299 2053
rect 1305 2047 1330 2053
rect 96 2037 97 2043
rect 103 2042 1311 2043
rect 103 2038 111 2042
rect 115 2038 295 2042
rect 299 2038 375 2042
rect 379 2038 391 2042
rect 395 2038 463 2042
rect 467 2038 535 2042
rect 539 2038 551 2042
rect 555 2038 615 2042
rect 619 2038 639 2042
rect 643 2038 695 2042
rect 699 2038 719 2042
rect 723 2038 775 2042
rect 779 2038 799 2042
rect 803 2038 847 2042
rect 851 2038 887 2042
rect 891 2038 919 2042
rect 923 2038 975 2042
rect 979 2038 983 2042
rect 987 2038 1047 2042
rect 1051 2038 1063 2042
rect 1067 2038 1119 2042
rect 1123 2038 1183 2042
rect 1187 2038 1239 2042
rect 1243 2038 1287 2042
rect 1291 2038 1311 2042
rect 103 2037 1311 2038
rect 1317 2037 1318 2043
rect 1324 2035 1330 2047
rect 1324 2034 2527 2035
rect 1324 2030 1327 2034
rect 1331 2030 1351 2034
rect 1355 2030 1407 2034
rect 1411 2030 1423 2034
rect 1427 2030 1487 2034
rect 1491 2030 1519 2034
rect 1523 2030 1575 2034
rect 1579 2030 1615 2034
rect 1619 2030 1663 2034
rect 1667 2030 1719 2034
rect 1723 2030 1767 2034
rect 1771 2030 1823 2034
rect 1827 2030 1879 2034
rect 1883 2030 1935 2034
rect 1939 2030 2007 2034
rect 2011 2030 2055 2034
rect 2059 2030 2151 2034
rect 2155 2030 2183 2034
rect 2187 2030 2303 2034
rect 2307 2030 2319 2034
rect 2323 2030 2439 2034
rect 2443 2030 2503 2034
rect 2507 2030 2527 2034
rect 1324 2029 2527 2030
rect 2533 2029 2534 2035
rect 84 1981 85 1987
rect 91 1986 1299 1987
rect 91 1982 111 1986
rect 115 1982 135 1986
rect 139 1982 207 1986
rect 211 1982 279 1986
rect 283 1982 287 1986
rect 291 1982 359 1986
rect 363 1982 383 1986
rect 387 1982 447 1986
rect 451 1982 487 1986
rect 491 1982 535 1986
rect 539 1982 591 1986
rect 595 1982 623 1986
rect 627 1982 695 1986
rect 699 1982 703 1986
rect 707 1982 783 1986
rect 787 1982 799 1986
rect 803 1982 871 1986
rect 875 1982 903 1986
rect 907 1982 959 1986
rect 963 1982 1015 1986
rect 1019 1982 1047 1986
rect 1051 1982 1287 1986
rect 1291 1982 1299 1986
rect 91 1981 1299 1982
rect 1305 1981 1306 1987
rect 1310 1973 1311 1979
rect 1317 1978 2539 1979
rect 1317 1974 1327 1978
rect 1331 1974 1367 1978
rect 1371 1974 1439 1978
rect 1443 1974 1455 1978
rect 1459 1974 1535 1978
rect 1539 1974 1543 1978
rect 1547 1974 1631 1978
rect 1635 1974 1639 1978
rect 1643 1974 1735 1978
rect 1739 1974 1839 1978
rect 1843 1974 1943 1978
rect 1947 1974 1951 1978
rect 1955 1974 2047 1978
rect 2051 1974 2071 1978
rect 2075 1974 2151 1978
rect 2155 1974 2199 1978
rect 2203 1974 2255 1978
rect 2259 1974 2335 1978
rect 2339 1974 2367 1978
rect 2371 1974 2455 1978
rect 2459 1974 2503 1978
rect 2507 1974 2539 1978
rect 1317 1973 2539 1974
rect 2545 1973 2546 1979
rect 1298 1931 1299 1937
rect 1305 1931 1330 1937
rect 96 1921 97 1927
rect 103 1926 1311 1927
rect 103 1922 111 1926
rect 115 1922 151 1926
rect 155 1922 223 1926
rect 227 1922 239 1926
rect 243 1922 303 1926
rect 307 1922 375 1926
rect 379 1922 399 1926
rect 403 1922 503 1926
rect 507 1922 527 1926
rect 531 1922 607 1926
rect 611 1922 687 1926
rect 691 1922 711 1926
rect 715 1922 815 1926
rect 819 1922 863 1926
rect 867 1922 919 1926
rect 923 1922 1031 1926
rect 1035 1922 1039 1926
rect 1043 1922 1287 1926
rect 1291 1922 1311 1926
rect 103 1921 1311 1922
rect 1317 1921 1318 1927
rect 1324 1923 1330 1931
rect 1324 1922 2527 1923
rect 1324 1918 1327 1922
rect 1331 1918 1439 1922
rect 1443 1918 1527 1922
rect 1531 1918 1615 1922
rect 1619 1918 1623 1922
rect 1627 1918 1711 1922
rect 1715 1918 1719 1922
rect 1723 1918 1815 1922
rect 1819 1918 1823 1922
rect 1827 1918 1919 1922
rect 1923 1918 1927 1922
rect 1931 1918 2015 1922
rect 2019 1918 2031 1922
rect 2035 1918 2111 1922
rect 2115 1918 2135 1922
rect 2139 1918 2199 1922
rect 2203 1918 2239 1922
rect 2243 1918 2287 1922
rect 2291 1918 2351 1922
rect 2355 1918 2375 1922
rect 2379 1918 2439 1922
rect 2443 1918 2503 1922
rect 2507 1918 2527 1922
rect 1324 1917 2527 1918
rect 2533 1917 2534 1923
rect 84 1869 85 1875
rect 91 1874 1299 1875
rect 91 1870 111 1874
rect 115 1870 135 1874
rect 139 1870 191 1874
rect 195 1870 223 1874
rect 227 1870 263 1874
rect 267 1870 335 1874
rect 339 1870 359 1874
rect 363 1870 407 1874
rect 411 1870 479 1874
rect 483 1870 511 1874
rect 515 1870 551 1874
rect 555 1870 615 1874
rect 619 1870 671 1874
rect 675 1870 679 1874
rect 683 1870 743 1874
rect 747 1870 815 1874
rect 819 1870 847 1874
rect 851 1870 887 1874
rect 891 1870 959 1874
rect 963 1870 1023 1874
rect 1027 1870 1039 1874
rect 1043 1870 1287 1874
rect 1291 1870 1299 1874
rect 91 1869 1299 1870
rect 1305 1869 1306 1875
rect 1310 1865 1311 1871
rect 1317 1870 2539 1871
rect 1317 1866 1327 1870
rect 1331 1866 1535 1870
rect 1539 1866 1543 1870
rect 1547 1866 1607 1870
rect 1611 1866 1631 1870
rect 1635 1866 1687 1870
rect 1691 1866 1727 1870
rect 1731 1866 1783 1870
rect 1787 1866 1831 1870
rect 1835 1866 1879 1870
rect 1883 1866 1935 1870
rect 1939 1866 1983 1870
rect 1987 1866 2031 1870
rect 2035 1866 2079 1870
rect 2083 1866 2127 1870
rect 2131 1866 2175 1870
rect 2179 1866 2215 1870
rect 2219 1866 2271 1870
rect 2275 1866 2303 1870
rect 2307 1866 2367 1870
rect 2371 1866 2391 1870
rect 2395 1866 2455 1870
rect 2459 1866 2503 1870
rect 2507 1866 2539 1870
rect 1317 1865 2539 1866
rect 2545 1865 2546 1871
rect 1298 1819 1299 1825
rect 1305 1819 1330 1825
rect 1324 1815 1330 1819
rect 96 1809 97 1815
rect 103 1814 1311 1815
rect 103 1810 111 1814
rect 115 1810 151 1814
rect 155 1810 207 1814
rect 211 1810 231 1814
rect 235 1810 279 1814
rect 283 1810 335 1814
rect 339 1810 351 1814
rect 355 1810 423 1814
rect 427 1810 439 1814
rect 443 1810 495 1814
rect 499 1810 535 1814
rect 539 1810 567 1814
rect 571 1810 631 1814
rect 635 1810 695 1814
rect 699 1810 719 1814
rect 723 1810 759 1814
rect 763 1810 799 1814
rect 803 1810 831 1814
rect 835 1810 879 1814
rect 883 1810 903 1814
rect 907 1810 959 1814
rect 963 1810 975 1814
rect 979 1810 1039 1814
rect 1043 1810 1055 1814
rect 1059 1810 1119 1814
rect 1123 1810 1287 1814
rect 1291 1810 1311 1814
rect 103 1809 1311 1810
rect 1317 1809 1318 1815
rect 1324 1814 2527 1815
rect 1324 1810 1327 1814
rect 1331 1810 1463 1814
rect 1467 1810 1519 1814
rect 1523 1810 1559 1814
rect 1563 1810 1591 1814
rect 1595 1810 1663 1814
rect 1667 1810 1671 1814
rect 1675 1810 1767 1814
rect 1771 1810 1863 1814
rect 1867 1810 1879 1814
rect 1883 1810 1967 1814
rect 1971 1810 1983 1814
rect 1987 1810 2063 1814
rect 2067 1810 2087 1814
rect 2091 1810 2159 1814
rect 2163 1810 2183 1814
rect 2187 1810 2255 1814
rect 2259 1810 2271 1814
rect 2275 1810 2351 1814
rect 2355 1810 2367 1814
rect 2371 1810 2439 1814
rect 2443 1810 2503 1814
rect 2507 1810 2527 1814
rect 1324 1809 2527 1810
rect 2533 1809 2534 1815
rect 2166 1796 2172 1797
rect 2402 1796 2408 1797
rect 2166 1792 2167 1796
rect 2171 1792 2403 1796
rect 2407 1792 2408 1796
rect 2166 1791 2172 1792
rect 2402 1791 2408 1792
rect 84 1753 85 1759
rect 91 1758 1299 1759
rect 91 1754 111 1758
rect 115 1754 135 1758
rect 139 1754 215 1758
rect 219 1754 239 1758
rect 243 1754 319 1758
rect 323 1754 351 1758
rect 355 1754 423 1758
rect 427 1754 463 1758
rect 467 1754 519 1758
rect 523 1754 575 1758
rect 579 1754 615 1758
rect 619 1754 679 1758
rect 683 1754 703 1758
rect 707 1754 783 1758
rect 787 1754 863 1758
rect 867 1754 887 1758
rect 891 1754 943 1758
rect 947 1754 991 1758
rect 995 1754 1023 1758
rect 1027 1754 1103 1758
rect 1107 1754 1287 1758
rect 1291 1754 1299 1758
rect 91 1753 1299 1754
rect 1305 1753 1306 1759
rect 1310 1753 1311 1759
rect 1317 1758 2539 1759
rect 1317 1754 1327 1758
rect 1331 1754 1375 1758
rect 1379 1754 1471 1758
rect 1475 1754 1479 1758
rect 1483 1754 1567 1758
rect 1571 1754 1575 1758
rect 1579 1754 1671 1758
rect 1675 1754 1679 1758
rect 1683 1754 1775 1758
rect 1779 1754 1783 1758
rect 1787 1754 1887 1758
rect 1891 1754 1895 1758
rect 1899 1754 1999 1758
rect 2003 1754 2103 1758
rect 2107 1754 2111 1758
rect 2115 1754 2199 1758
rect 2203 1754 2231 1758
rect 2235 1754 2287 1758
rect 2291 1754 2351 1758
rect 2355 1754 2383 1758
rect 2387 1754 2455 1758
rect 2459 1754 2503 1758
rect 2507 1754 2539 1758
rect 1317 1753 2539 1754
rect 2545 1753 2546 1759
rect 1298 1707 1299 1713
rect 1305 1707 1330 1713
rect 1324 1706 2527 1707
rect 96 1697 97 1703
rect 103 1702 1311 1703
rect 103 1698 111 1702
rect 115 1698 151 1702
rect 155 1698 191 1702
rect 195 1698 255 1702
rect 259 1698 271 1702
rect 275 1698 351 1702
rect 355 1698 367 1702
rect 371 1698 439 1702
rect 443 1698 479 1702
rect 483 1698 535 1702
rect 539 1698 591 1702
rect 595 1698 639 1702
rect 643 1698 695 1702
rect 699 1698 743 1702
rect 747 1698 799 1702
rect 803 1698 847 1702
rect 851 1698 903 1702
rect 907 1698 951 1702
rect 955 1698 1007 1702
rect 1011 1698 1063 1702
rect 1067 1698 1119 1702
rect 1123 1698 1175 1702
rect 1179 1698 1287 1702
rect 1291 1698 1311 1702
rect 103 1697 1311 1698
rect 1317 1697 1318 1703
rect 1324 1702 1327 1706
rect 1331 1702 1351 1706
rect 1355 1702 1359 1706
rect 1363 1702 1431 1706
rect 1435 1702 1455 1706
rect 1459 1702 1535 1706
rect 1539 1702 1551 1706
rect 1555 1702 1647 1706
rect 1651 1702 1655 1706
rect 1659 1702 1759 1706
rect 1763 1702 1871 1706
rect 1875 1702 1879 1706
rect 1883 1702 1983 1706
rect 1987 1702 2015 1706
rect 2019 1702 2095 1706
rect 2099 1702 2159 1706
rect 2163 1702 2215 1706
rect 2219 1702 2311 1706
rect 2315 1702 2335 1706
rect 2339 1702 2439 1706
rect 2443 1702 2503 1706
rect 2507 1702 2527 1706
rect 1324 1701 2527 1702
rect 2533 1701 2534 1707
rect 1382 1668 1388 1669
rect 1670 1668 1676 1669
rect 1382 1664 1383 1668
rect 1387 1664 1671 1668
rect 1675 1664 1676 1668
rect 1382 1663 1388 1664
rect 1670 1663 1676 1664
rect 84 1645 85 1651
rect 91 1650 1299 1651
rect 91 1646 111 1650
rect 115 1646 175 1650
rect 179 1646 215 1650
rect 219 1646 255 1650
rect 259 1646 271 1650
rect 275 1646 335 1650
rect 339 1646 407 1650
rect 411 1646 423 1650
rect 427 1646 479 1650
rect 483 1646 519 1650
rect 523 1646 559 1650
rect 563 1646 623 1650
rect 627 1646 647 1650
rect 651 1646 727 1650
rect 731 1646 743 1650
rect 747 1646 831 1650
rect 835 1646 839 1650
rect 843 1646 935 1650
rect 939 1646 943 1650
rect 947 1646 1047 1650
rect 1051 1646 1055 1650
rect 1059 1646 1159 1650
rect 1163 1646 1175 1650
rect 1179 1646 1287 1650
rect 1291 1646 1299 1650
rect 91 1645 1299 1646
rect 1305 1645 1306 1651
rect 1310 1641 1311 1647
rect 1317 1646 2539 1647
rect 1317 1642 1327 1646
rect 1331 1642 1367 1646
rect 1371 1642 1431 1646
rect 1435 1642 1447 1646
rect 1451 1642 1519 1646
rect 1523 1642 1551 1646
rect 1555 1642 1599 1646
rect 1603 1642 1663 1646
rect 1667 1642 1679 1646
rect 1683 1642 1751 1646
rect 1755 1642 1775 1646
rect 1779 1642 1839 1646
rect 1843 1642 1895 1646
rect 1899 1642 1935 1646
rect 1939 1642 2031 1646
rect 2035 1642 2055 1646
rect 2059 1642 2175 1646
rect 2179 1642 2183 1646
rect 2187 1642 2327 1646
rect 2331 1642 2455 1646
rect 2459 1642 2503 1646
rect 2507 1642 2539 1646
rect 1317 1641 2539 1642
rect 2545 1641 2546 1647
rect 1298 1603 1299 1609
rect 1305 1603 1330 1609
rect 96 1593 97 1599
rect 103 1598 1311 1599
rect 103 1594 111 1598
rect 115 1594 231 1598
rect 235 1594 287 1598
rect 291 1594 351 1598
rect 355 1594 423 1598
rect 427 1594 495 1598
rect 499 1594 503 1598
rect 507 1594 575 1598
rect 579 1594 599 1598
rect 603 1594 663 1598
rect 667 1594 703 1598
rect 707 1594 759 1598
rect 763 1594 815 1598
rect 819 1594 855 1598
rect 859 1594 935 1598
rect 939 1594 959 1598
rect 963 1594 1063 1598
rect 1067 1594 1071 1598
rect 1075 1594 1191 1598
rect 1195 1594 1287 1598
rect 1291 1594 1311 1598
rect 103 1593 1311 1594
rect 1317 1593 1318 1599
rect 1324 1591 1330 1603
rect 1324 1590 2527 1591
rect 1324 1586 1327 1590
rect 1331 1586 1351 1590
rect 1355 1586 1415 1590
rect 1419 1586 1423 1590
rect 1427 1586 1503 1590
rect 1507 1586 1527 1590
rect 1531 1586 1583 1590
rect 1587 1586 1647 1590
rect 1651 1586 1663 1590
rect 1667 1586 1735 1590
rect 1739 1586 1783 1590
rect 1787 1586 1823 1590
rect 1827 1586 1919 1590
rect 1923 1586 1935 1590
rect 1939 1586 2039 1590
rect 2043 1586 2103 1590
rect 2107 1586 2167 1590
rect 2171 1586 2279 1590
rect 2283 1586 2311 1590
rect 2315 1586 2439 1590
rect 2443 1586 2503 1590
rect 2507 1586 2527 1590
rect 1324 1585 2527 1586
rect 2533 1585 2534 1591
rect 618 1572 624 1573
rect 954 1572 960 1573
rect 618 1568 619 1572
rect 623 1568 955 1572
rect 959 1568 960 1572
rect 618 1567 624 1568
rect 954 1567 960 1568
rect 84 1533 85 1539
rect 91 1538 1299 1539
rect 91 1534 111 1538
rect 115 1534 271 1538
rect 275 1534 335 1538
rect 339 1534 407 1538
rect 411 1534 471 1538
rect 475 1534 487 1538
rect 491 1534 551 1538
rect 555 1534 583 1538
rect 587 1534 639 1538
rect 643 1534 687 1538
rect 691 1534 735 1538
rect 739 1534 799 1538
rect 803 1534 839 1538
rect 843 1534 919 1538
rect 923 1534 951 1538
rect 955 1534 1047 1538
rect 1051 1534 1063 1538
rect 1067 1534 1175 1538
rect 1179 1534 1287 1538
rect 1291 1534 1299 1538
rect 91 1533 1299 1534
rect 1305 1533 1306 1539
rect 1310 1533 1311 1539
rect 1317 1538 2539 1539
rect 1317 1534 1327 1538
rect 1331 1534 1367 1538
rect 1371 1534 1439 1538
rect 1443 1534 1543 1538
rect 1547 1534 1647 1538
rect 1651 1534 1663 1538
rect 1667 1534 1751 1538
rect 1755 1534 1799 1538
rect 1803 1534 1855 1538
rect 1859 1534 1951 1538
rect 1955 1534 1959 1538
rect 1963 1534 2055 1538
rect 2059 1534 2119 1538
rect 2123 1534 2151 1538
rect 2155 1534 2247 1538
rect 2251 1534 2295 1538
rect 2299 1534 2343 1538
rect 2347 1534 2439 1538
rect 2443 1534 2455 1538
rect 2459 1534 2503 1538
rect 2507 1534 2539 1538
rect 1317 1533 2539 1534
rect 2545 1533 2546 1539
rect 1298 1491 1299 1497
rect 1305 1491 1330 1497
rect 96 1481 97 1487
rect 103 1486 1311 1487
rect 103 1482 111 1486
rect 115 1482 375 1486
rect 379 1482 463 1486
rect 467 1482 487 1486
rect 491 1482 559 1486
rect 563 1482 567 1486
rect 571 1482 655 1486
rect 659 1482 751 1486
rect 755 1482 855 1486
rect 859 1482 959 1486
rect 963 1482 967 1486
rect 971 1482 1063 1486
rect 1067 1482 1079 1486
rect 1083 1482 1167 1486
rect 1171 1482 1191 1486
rect 1195 1482 1287 1486
rect 1291 1482 1311 1486
rect 103 1481 1311 1482
rect 1317 1481 1318 1487
rect 1324 1483 1330 1491
rect 1324 1482 2527 1483
rect 1324 1478 1327 1482
rect 1331 1478 1351 1482
rect 1355 1478 1423 1482
rect 1427 1478 1519 1482
rect 1523 1478 1527 1482
rect 1531 1478 1615 1482
rect 1619 1478 1631 1482
rect 1635 1478 1711 1482
rect 1715 1478 1735 1482
rect 1739 1478 1815 1482
rect 1819 1478 1839 1482
rect 1843 1478 1927 1482
rect 1931 1478 1943 1482
rect 1947 1478 2039 1482
rect 2043 1478 2047 1482
rect 2051 1478 2135 1482
rect 2139 1478 2175 1482
rect 2179 1478 2231 1482
rect 2235 1478 2303 1482
rect 2307 1478 2327 1482
rect 2331 1478 2423 1482
rect 2427 1478 2439 1482
rect 2443 1478 2503 1482
rect 2507 1478 2527 1482
rect 1324 1477 2527 1478
rect 2533 1477 2534 1483
rect 84 1429 85 1435
rect 91 1434 1299 1435
rect 91 1430 111 1434
rect 115 1430 231 1434
rect 235 1430 319 1434
rect 323 1430 359 1434
rect 363 1430 415 1434
rect 419 1430 447 1434
rect 451 1430 511 1434
rect 515 1430 543 1434
rect 547 1430 615 1434
rect 619 1430 639 1434
rect 643 1430 711 1434
rect 715 1430 735 1434
rect 739 1430 807 1434
rect 811 1430 839 1434
rect 843 1430 895 1434
rect 899 1430 943 1434
rect 947 1430 991 1434
rect 995 1430 1047 1434
rect 1051 1430 1087 1434
rect 1091 1430 1151 1434
rect 1155 1430 1287 1434
rect 1291 1430 1299 1434
rect 91 1429 1299 1430
rect 1305 1429 1306 1435
rect 1310 1421 1311 1427
rect 1317 1426 2539 1427
rect 1317 1422 1327 1426
rect 1331 1422 1367 1426
rect 1371 1422 1423 1426
rect 1427 1422 1439 1426
rect 1443 1422 1503 1426
rect 1507 1422 1535 1426
rect 1539 1422 1591 1426
rect 1595 1422 1631 1426
rect 1635 1422 1679 1426
rect 1683 1422 1727 1426
rect 1731 1422 1775 1426
rect 1779 1422 1831 1426
rect 1835 1422 1879 1426
rect 1883 1422 1943 1426
rect 1947 1422 1991 1426
rect 1995 1422 2063 1426
rect 2067 1422 2111 1426
rect 2115 1422 2191 1426
rect 2195 1422 2231 1426
rect 2235 1422 2319 1426
rect 2323 1422 2351 1426
rect 2355 1422 2455 1426
rect 2459 1422 2503 1426
rect 2507 1422 2539 1426
rect 1317 1421 2539 1422
rect 2545 1421 2546 1427
rect 96 1377 97 1383
rect 103 1382 1311 1383
rect 103 1378 111 1382
rect 115 1378 151 1382
rect 155 1378 215 1382
rect 219 1378 247 1382
rect 251 1378 311 1382
rect 315 1378 335 1382
rect 339 1378 407 1382
rect 411 1378 431 1382
rect 435 1378 511 1382
rect 515 1378 527 1382
rect 531 1378 607 1382
rect 611 1378 631 1382
rect 635 1378 703 1382
rect 707 1378 727 1382
rect 731 1378 799 1382
rect 803 1378 823 1382
rect 827 1378 895 1382
rect 899 1378 911 1382
rect 915 1378 999 1382
rect 1003 1378 1007 1382
rect 1011 1378 1103 1382
rect 1107 1378 1287 1382
rect 1291 1378 1311 1382
rect 103 1377 1311 1378
rect 1317 1377 1318 1383
rect 1298 1365 1299 1371
rect 1305 1370 2527 1371
rect 1305 1366 1327 1370
rect 1331 1366 1351 1370
rect 1355 1366 1407 1370
rect 1411 1366 1479 1370
rect 1483 1366 1487 1370
rect 1491 1366 1567 1370
rect 1571 1366 1575 1370
rect 1579 1366 1655 1370
rect 1659 1366 1663 1370
rect 1667 1366 1751 1370
rect 1755 1366 1759 1370
rect 1763 1366 1855 1370
rect 1859 1366 1863 1370
rect 1867 1366 1967 1370
rect 1971 1366 1975 1370
rect 1979 1366 2079 1370
rect 2083 1366 2095 1370
rect 2099 1366 2199 1370
rect 2203 1366 2215 1370
rect 2219 1366 2327 1370
rect 2331 1366 2335 1370
rect 2339 1366 2439 1370
rect 2443 1366 2503 1370
rect 2507 1366 2527 1370
rect 1305 1365 2527 1366
rect 2533 1365 2534 1371
rect 84 1325 85 1331
rect 91 1330 1299 1331
rect 91 1326 111 1330
rect 115 1326 135 1330
rect 139 1326 199 1330
rect 203 1326 215 1330
rect 219 1326 295 1330
rect 299 1326 319 1330
rect 323 1326 391 1330
rect 395 1326 415 1330
rect 419 1326 495 1330
rect 499 1326 511 1330
rect 515 1326 591 1330
rect 595 1326 599 1330
rect 603 1326 687 1330
rect 691 1326 783 1330
rect 787 1326 879 1330
rect 883 1326 983 1330
rect 987 1326 1287 1330
rect 1291 1326 1299 1330
rect 91 1325 1299 1326
rect 1305 1325 1306 1331
rect 1310 1305 1311 1311
rect 1317 1310 2539 1311
rect 1317 1306 1327 1310
rect 1331 1306 1367 1310
rect 1371 1306 1423 1310
rect 1427 1306 1495 1310
rect 1499 1306 1519 1310
rect 1523 1306 1583 1310
rect 1587 1306 1615 1310
rect 1619 1306 1671 1310
rect 1675 1306 1719 1310
rect 1723 1306 1767 1310
rect 1771 1306 1823 1310
rect 1827 1306 1871 1310
rect 1875 1306 1919 1310
rect 1923 1306 1983 1310
rect 1987 1306 2015 1310
rect 2019 1306 2095 1310
rect 2099 1306 2103 1310
rect 2107 1306 2183 1310
rect 2187 1306 2215 1310
rect 2219 1306 2255 1310
rect 2259 1306 2327 1310
rect 2331 1306 2343 1310
rect 2347 1306 2399 1310
rect 2403 1306 2455 1310
rect 2459 1306 2503 1310
rect 2507 1306 2539 1310
rect 1317 1305 2539 1306
rect 2545 1305 2546 1311
rect 96 1273 97 1279
rect 103 1278 1311 1279
rect 103 1274 111 1278
rect 115 1274 151 1278
rect 155 1274 191 1278
rect 195 1274 231 1278
rect 235 1274 247 1278
rect 251 1274 303 1278
rect 307 1274 335 1278
rect 339 1274 367 1278
rect 371 1274 431 1278
rect 435 1274 439 1278
rect 443 1274 527 1278
rect 531 1274 615 1278
rect 619 1274 639 1278
rect 643 1274 703 1278
rect 707 1274 775 1278
rect 779 1274 799 1278
rect 803 1274 895 1278
rect 899 1274 927 1278
rect 931 1274 1095 1278
rect 1099 1274 1239 1278
rect 1243 1274 1287 1278
rect 1291 1274 1311 1278
rect 103 1273 1311 1274
rect 1317 1273 1318 1279
rect 1298 1237 1299 1243
rect 1305 1242 2527 1243
rect 1305 1238 1327 1242
rect 1331 1238 1351 1242
rect 1355 1238 1407 1242
rect 1411 1238 1447 1242
rect 1451 1238 1503 1242
rect 1507 1238 1575 1242
rect 1579 1238 1599 1242
rect 1603 1238 1695 1242
rect 1699 1238 1703 1242
rect 1707 1238 1807 1242
rect 1811 1238 1815 1242
rect 1819 1238 1903 1242
rect 1907 1238 1927 1242
rect 1931 1238 1999 1242
rect 2003 1238 2031 1242
rect 2035 1238 2087 1242
rect 2091 1238 2127 1242
rect 2131 1238 2167 1242
rect 2171 1238 2215 1242
rect 2219 1238 2239 1242
rect 2243 1238 2295 1242
rect 2299 1238 2311 1242
rect 2315 1238 2375 1242
rect 2379 1238 2383 1242
rect 2387 1238 2439 1242
rect 2443 1238 2503 1242
rect 2507 1238 2527 1242
rect 1305 1237 2527 1238
rect 2533 1237 2534 1243
rect 84 1221 85 1227
rect 91 1226 1299 1227
rect 91 1222 111 1226
rect 115 1222 175 1226
rect 179 1222 231 1226
rect 235 1222 287 1226
rect 291 1222 351 1226
rect 355 1222 407 1226
rect 411 1222 423 1226
rect 427 1222 463 1226
rect 467 1222 511 1226
rect 515 1222 519 1226
rect 523 1222 575 1226
rect 579 1222 623 1226
rect 627 1222 631 1226
rect 635 1222 687 1226
rect 691 1222 743 1226
rect 747 1222 759 1226
rect 763 1222 799 1226
rect 803 1222 855 1226
rect 859 1222 911 1226
rect 915 1222 1079 1226
rect 1083 1222 1223 1226
rect 1227 1222 1287 1226
rect 1291 1222 1299 1226
rect 91 1221 1299 1222
rect 1305 1221 1306 1227
rect 1950 1204 1956 1205
rect 2262 1204 2268 1205
rect 1950 1200 1951 1204
rect 1955 1200 2263 1204
rect 2267 1200 2268 1204
rect 1950 1199 1956 1200
rect 2262 1199 2268 1200
rect 1310 1185 1311 1191
rect 1317 1190 2539 1191
rect 1317 1186 1327 1190
rect 1331 1186 1367 1190
rect 1371 1186 1463 1190
rect 1467 1186 1471 1190
rect 1475 1186 1591 1190
rect 1595 1186 1599 1190
rect 1603 1186 1711 1190
rect 1715 1186 1735 1190
rect 1739 1186 1831 1190
rect 1835 1186 1863 1190
rect 1867 1186 1943 1190
rect 1947 1186 1983 1190
rect 1987 1186 2047 1190
rect 2051 1186 2087 1190
rect 2091 1186 2143 1190
rect 2147 1186 2191 1190
rect 2195 1186 2231 1190
rect 2235 1186 2287 1190
rect 2291 1186 2311 1190
rect 2315 1186 2383 1190
rect 2387 1186 2391 1190
rect 2395 1186 2455 1190
rect 2459 1186 2503 1190
rect 2507 1186 2539 1190
rect 1317 1185 2539 1186
rect 2545 1185 2546 1191
rect 96 1165 97 1171
rect 103 1170 1311 1171
rect 103 1166 111 1170
rect 115 1166 367 1170
rect 371 1166 423 1170
rect 427 1166 479 1170
rect 483 1166 535 1170
rect 539 1166 591 1170
rect 595 1166 647 1170
rect 651 1166 703 1170
rect 707 1166 759 1170
rect 763 1166 815 1170
rect 819 1166 871 1170
rect 875 1166 927 1170
rect 931 1166 983 1170
rect 987 1166 1287 1170
rect 1291 1166 1311 1170
rect 103 1165 1311 1166
rect 1317 1165 1318 1171
rect 1298 1129 1299 1135
rect 1305 1134 2527 1135
rect 1305 1130 1327 1134
rect 1331 1130 1351 1134
rect 1355 1130 1367 1134
rect 1371 1130 1447 1134
rect 1451 1130 1455 1134
rect 1459 1130 1535 1134
rect 1539 1130 1583 1134
rect 1587 1130 1631 1134
rect 1635 1130 1719 1134
rect 1723 1130 1807 1134
rect 1811 1130 1847 1134
rect 1851 1130 1895 1134
rect 1899 1130 1967 1134
rect 1971 1130 1983 1134
rect 1987 1130 2071 1134
rect 2075 1130 2159 1134
rect 2163 1130 2175 1134
rect 2179 1130 2255 1134
rect 2259 1130 2271 1134
rect 2275 1130 2359 1134
rect 2363 1130 2367 1134
rect 2371 1130 2439 1134
rect 2443 1130 2503 1134
rect 2507 1130 2527 1134
rect 1305 1129 2527 1130
rect 2533 1129 2534 1135
rect 84 1109 85 1115
rect 91 1114 1299 1115
rect 91 1110 111 1114
rect 115 1110 223 1114
rect 227 1110 311 1114
rect 315 1110 399 1114
rect 403 1110 407 1114
rect 411 1110 463 1114
rect 467 1110 495 1114
rect 499 1110 519 1114
rect 523 1110 575 1114
rect 579 1110 591 1114
rect 595 1110 631 1114
rect 635 1110 679 1114
rect 683 1110 687 1114
rect 691 1110 743 1114
rect 747 1110 767 1114
rect 771 1110 799 1114
rect 803 1110 847 1114
rect 851 1110 855 1114
rect 859 1110 911 1114
rect 915 1110 927 1114
rect 931 1110 967 1114
rect 971 1110 1015 1114
rect 1019 1110 1103 1114
rect 1107 1110 1287 1114
rect 1291 1110 1299 1114
rect 91 1109 1299 1110
rect 1305 1109 1306 1115
rect 1958 1092 1964 1093
rect 2382 1092 2388 1093
rect 1958 1088 1959 1092
rect 1963 1088 2383 1092
rect 2387 1088 2388 1092
rect 1958 1087 1964 1088
rect 2382 1087 2388 1088
rect 1310 1069 1311 1075
rect 1317 1074 2539 1075
rect 1317 1070 1327 1074
rect 1331 1070 1383 1074
rect 1387 1070 1431 1074
rect 1435 1070 1463 1074
rect 1467 1070 1495 1074
rect 1499 1070 1551 1074
rect 1555 1070 1567 1074
rect 1571 1070 1639 1074
rect 1643 1070 1647 1074
rect 1651 1070 1703 1074
rect 1707 1070 1735 1074
rect 1739 1070 1767 1074
rect 1771 1070 1823 1074
rect 1827 1070 1839 1074
rect 1843 1070 1911 1074
rect 1915 1070 1919 1074
rect 1923 1070 1999 1074
rect 2003 1070 2007 1074
rect 2011 1070 2087 1074
rect 2091 1070 2111 1074
rect 2115 1070 2175 1074
rect 2179 1070 2231 1074
rect 2235 1070 2271 1074
rect 2275 1070 2351 1074
rect 2355 1070 2375 1074
rect 2379 1070 2455 1074
rect 2459 1070 2503 1074
rect 2507 1070 2539 1074
rect 1317 1069 2539 1070
rect 2545 1069 2546 1075
rect 96 1053 97 1059
rect 103 1058 1311 1059
rect 103 1054 111 1058
rect 115 1054 151 1058
rect 155 1054 207 1058
rect 211 1054 239 1058
rect 243 1054 303 1058
rect 307 1054 327 1058
rect 331 1054 415 1058
rect 419 1054 511 1058
rect 515 1054 535 1058
rect 539 1054 607 1058
rect 611 1054 655 1058
rect 659 1054 695 1058
rect 699 1054 767 1058
rect 771 1054 783 1058
rect 787 1054 863 1058
rect 867 1054 879 1058
rect 883 1054 943 1058
rect 947 1054 983 1058
rect 987 1054 1031 1058
rect 1035 1054 1095 1058
rect 1099 1054 1119 1058
rect 1123 1054 1207 1058
rect 1211 1054 1287 1058
rect 1291 1054 1311 1058
rect 103 1053 1311 1054
rect 1317 1053 1318 1059
rect 774 1036 780 1037
rect 1226 1036 1232 1037
rect 774 1032 775 1036
rect 779 1032 1227 1036
rect 1231 1032 1232 1036
rect 774 1031 780 1032
rect 1226 1031 1232 1032
rect 1298 1009 1299 1015
rect 1305 1014 2527 1015
rect 1305 1010 1327 1014
rect 1331 1010 1415 1014
rect 1419 1010 1479 1014
rect 1483 1010 1511 1014
rect 1515 1010 1551 1014
rect 1555 1010 1567 1014
rect 1571 1010 1623 1014
rect 1627 1010 1679 1014
rect 1683 1010 1687 1014
rect 1691 1010 1735 1014
rect 1739 1010 1751 1014
rect 1755 1010 1807 1014
rect 1811 1010 1823 1014
rect 1827 1010 1887 1014
rect 1891 1010 1903 1014
rect 1907 1010 1983 1014
rect 1987 1010 1991 1014
rect 1995 1010 2095 1014
rect 2099 1010 2215 1014
rect 2219 1010 2335 1014
rect 2339 1010 2439 1014
rect 2443 1010 2503 1014
rect 2507 1010 2527 1014
rect 1305 1009 2527 1010
rect 2533 1009 2534 1015
rect 84 997 85 1003
rect 91 1002 1299 1003
rect 91 998 111 1002
rect 115 998 135 1002
rect 139 998 191 1002
rect 195 998 215 1002
rect 219 998 287 1002
rect 291 998 327 1002
rect 331 998 399 1002
rect 403 998 439 1002
rect 443 998 519 1002
rect 523 998 551 1002
rect 555 998 639 1002
rect 643 998 663 1002
rect 667 998 751 1002
rect 755 998 759 1002
rect 763 998 847 1002
rect 851 998 863 1002
rect 867 998 935 1002
rect 939 998 967 1002
rect 971 998 1015 1002
rect 1019 998 1079 1002
rect 1083 998 1087 1002
rect 1091 998 1167 1002
rect 1171 998 1191 1002
rect 1195 998 1223 1002
rect 1227 998 1287 1002
rect 1291 998 1299 1002
rect 91 997 1299 998
rect 1305 997 1306 1003
rect 96 945 97 951
rect 103 950 1311 951
rect 103 946 111 950
rect 115 946 151 950
rect 155 946 207 950
rect 211 946 231 950
rect 235 946 295 950
rect 299 946 343 950
rect 347 946 399 950
rect 403 946 455 950
rect 459 946 511 950
rect 515 946 567 950
rect 571 946 623 950
rect 627 946 679 950
rect 683 946 735 950
rect 739 946 775 950
rect 779 946 831 950
rect 835 946 863 950
rect 867 946 927 950
rect 931 946 951 950
rect 955 946 1015 950
rect 1019 946 1031 950
rect 1035 946 1095 950
rect 1099 946 1103 950
rect 1107 946 1175 950
rect 1179 946 1183 950
rect 1187 946 1239 950
rect 1243 946 1287 950
rect 1291 946 1311 950
rect 103 945 1311 946
rect 1317 947 1318 951
rect 1317 946 2546 947
rect 1317 945 1327 946
rect 1310 942 1327 945
rect 1331 942 1367 946
rect 1371 942 1439 946
rect 1443 942 1527 946
rect 1531 942 1583 946
rect 1587 942 1615 946
rect 1619 942 1639 946
rect 1643 942 1695 946
rect 1699 942 1751 946
rect 1755 942 1791 946
rect 1795 942 1823 946
rect 1827 942 1895 946
rect 1899 942 1903 946
rect 1907 942 1999 946
rect 2003 942 2015 946
rect 2019 942 2111 946
rect 2115 942 2151 946
rect 2155 942 2231 946
rect 2235 942 2295 946
rect 2299 942 2351 946
rect 2355 942 2439 946
rect 2443 942 2455 946
rect 2459 942 2503 946
rect 2507 942 2546 946
rect 1310 941 2546 942
rect 84 889 85 895
rect 91 894 1299 895
rect 91 890 111 894
rect 115 890 135 894
rect 139 890 191 894
rect 195 890 247 894
rect 251 890 279 894
rect 283 890 343 894
rect 347 890 383 894
rect 387 890 439 894
rect 443 890 495 894
rect 499 890 543 894
rect 547 890 607 894
rect 611 890 647 894
rect 651 890 719 894
rect 723 890 743 894
rect 747 890 815 894
rect 819 890 839 894
rect 843 890 911 894
rect 915 890 927 894
rect 931 890 999 894
rect 1003 890 1007 894
rect 1011 890 1079 894
rect 1083 890 1087 894
rect 1091 890 1159 894
rect 1163 890 1167 894
rect 1171 890 1223 894
rect 1227 890 1287 894
rect 1291 890 1299 894
rect 91 889 1299 890
rect 1305 889 1306 895
rect 1298 887 1306 889
rect 1298 881 1299 887
rect 1305 886 2527 887
rect 1305 882 1327 886
rect 1331 882 1351 886
rect 1355 882 1423 886
rect 1427 882 1487 886
rect 1491 882 1511 886
rect 1515 882 1559 886
rect 1563 882 1599 886
rect 1603 882 1623 886
rect 1627 882 1679 886
rect 1683 882 1687 886
rect 1691 882 1751 886
rect 1755 882 1775 886
rect 1779 882 1815 886
rect 1819 882 1879 886
rect 1883 882 1887 886
rect 1891 882 1975 886
rect 1979 882 1999 886
rect 2003 882 2079 886
rect 2083 882 2135 886
rect 2139 882 2199 886
rect 2203 882 2279 886
rect 2283 882 2319 886
rect 2323 882 2423 886
rect 2427 882 2439 886
rect 2443 882 2503 886
rect 2507 882 2527 886
rect 1305 881 2527 882
rect 2533 881 2534 887
rect 1838 852 1844 853
rect 2302 852 2308 853
rect 1838 848 1839 852
rect 1843 848 2303 852
rect 2307 848 2308 852
rect 1838 847 1844 848
rect 2302 847 2308 848
rect 96 833 97 839
rect 103 838 1311 839
rect 103 834 111 838
rect 115 834 239 838
rect 243 834 263 838
rect 267 834 303 838
rect 307 834 359 838
rect 363 834 383 838
rect 387 834 455 838
rect 459 834 463 838
rect 467 834 551 838
rect 555 834 559 838
rect 563 834 639 838
rect 643 834 663 838
rect 667 834 727 838
rect 731 834 759 838
rect 763 834 807 838
rect 811 834 855 838
rect 859 834 895 838
rect 899 834 943 838
rect 947 834 983 838
rect 987 834 1023 838
rect 1027 834 1071 838
rect 1075 834 1103 838
rect 1107 834 1183 838
rect 1187 834 1239 838
rect 1243 834 1287 838
rect 1291 834 1311 838
rect 103 833 1311 834
rect 1317 833 1318 839
rect 1310 821 1311 827
rect 1317 826 2539 827
rect 1317 822 1327 826
rect 1331 822 1439 826
rect 1443 822 1503 826
rect 1507 822 1511 826
rect 1515 822 1575 826
rect 1579 822 1591 826
rect 1595 822 1639 826
rect 1643 822 1671 826
rect 1675 822 1703 826
rect 1707 822 1759 826
rect 1763 822 1767 826
rect 1771 822 1831 826
rect 1835 822 1847 826
rect 1851 822 1903 826
rect 1907 822 1935 826
rect 1939 822 1991 826
rect 1995 822 2023 826
rect 2027 822 2095 826
rect 2099 822 2111 826
rect 2115 822 2199 826
rect 2203 822 2215 826
rect 2219 822 2287 826
rect 2291 822 2335 826
rect 2339 822 2383 826
rect 2387 822 2455 826
rect 2459 822 2503 826
rect 2507 822 2539 826
rect 1317 821 2539 822
rect 2545 821 2546 827
rect 84 777 85 783
rect 91 782 1299 783
rect 91 778 111 782
rect 115 778 151 782
rect 155 778 223 782
rect 227 778 247 782
rect 251 778 287 782
rect 291 778 343 782
rect 347 778 367 782
rect 371 778 439 782
rect 443 778 447 782
rect 451 778 527 782
rect 531 778 535 782
rect 539 778 607 782
rect 611 778 623 782
rect 627 778 679 782
rect 683 778 711 782
rect 715 778 751 782
rect 755 778 791 782
rect 795 778 823 782
rect 827 778 879 782
rect 883 778 895 782
rect 899 778 967 782
rect 971 778 975 782
rect 979 778 1055 782
rect 1059 778 1287 782
rect 1291 778 1299 782
rect 91 777 1299 778
rect 1305 777 1306 783
rect 1298 765 1299 771
rect 1305 770 2527 771
rect 1305 766 1327 770
rect 1331 766 1351 770
rect 1355 766 1423 770
rect 1427 766 1447 770
rect 1451 766 1495 770
rect 1499 766 1567 770
rect 1571 766 1575 770
rect 1579 766 1655 770
rect 1659 766 1687 770
rect 1691 766 1743 770
rect 1747 766 1807 770
rect 1811 766 1831 770
rect 1835 766 1919 770
rect 1923 766 1927 770
rect 1931 766 2007 770
rect 2011 766 2039 770
rect 2043 766 2095 770
rect 2099 766 2143 770
rect 2147 766 2183 770
rect 2187 766 2247 770
rect 2251 766 2271 770
rect 2275 766 2351 770
rect 2355 766 2367 770
rect 2371 766 2439 770
rect 2443 766 2503 770
rect 2507 766 2527 770
rect 1305 765 2527 766
rect 2533 765 2534 771
rect 96 721 97 727
rect 103 726 1311 727
rect 103 722 111 726
rect 115 722 167 726
rect 171 722 175 726
rect 179 722 263 726
rect 267 722 343 726
rect 347 722 359 726
rect 363 722 423 726
rect 427 722 455 726
rect 459 722 503 726
rect 507 722 543 726
rect 547 722 575 726
rect 579 722 623 726
rect 627 722 639 726
rect 643 722 695 726
rect 699 722 703 726
rect 707 722 767 726
rect 771 722 839 726
rect 843 722 911 726
rect 915 722 991 726
rect 995 722 1287 726
rect 1291 722 1311 726
rect 103 721 1311 722
rect 1317 721 1318 727
rect 1974 724 1980 725
rect 2270 724 2276 725
rect 1974 720 1975 724
rect 1979 720 2271 724
rect 2275 720 2276 724
rect 1974 719 1980 720
rect 2270 719 2276 720
rect 1310 709 1311 715
rect 1317 714 2539 715
rect 1317 710 1327 714
rect 1331 710 1367 714
rect 1371 710 1431 714
rect 1435 710 1463 714
rect 1467 710 1535 714
rect 1539 710 1583 714
rect 1587 710 1639 714
rect 1643 710 1703 714
rect 1707 710 1751 714
rect 1755 710 1823 714
rect 1827 710 1863 714
rect 1867 710 1943 714
rect 1947 710 1967 714
rect 1971 710 2055 714
rect 2059 710 2063 714
rect 2067 710 2151 714
rect 2155 710 2159 714
rect 2163 710 2231 714
rect 2235 710 2263 714
rect 2267 710 2311 714
rect 2315 710 2367 714
rect 2371 710 2391 714
rect 2395 710 2455 714
rect 2459 710 2503 714
rect 2507 710 2539 714
rect 1317 709 2539 710
rect 2545 709 2546 715
rect 84 669 85 675
rect 91 674 1299 675
rect 91 670 111 674
rect 115 670 159 674
rect 163 670 215 674
rect 219 670 247 674
rect 251 670 295 674
rect 299 670 327 674
rect 331 670 375 674
rect 379 670 407 674
rect 411 670 455 674
rect 459 670 487 674
rect 491 670 527 674
rect 531 670 559 674
rect 563 670 591 674
rect 595 670 623 674
rect 627 670 655 674
rect 659 670 687 674
rect 691 670 719 674
rect 723 670 751 674
rect 755 670 783 674
rect 787 670 823 674
rect 827 670 847 674
rect 851 670 895 674
rect 899 670 919 674
rect 923 670 1287 674
rect 1291 670 1299 674
rect 91 669 1299 670
rect 1305 669 1306 675
rect 1298 649 1299 655
rect 1305 654 2527 655
rect 1305 650 1327 654
rect 1331 650 1351 654
rect 1355 650 1415 654
rect 1419 650 1479 654
rect 1483 650 1519 654
rect 1523 650 1559 654
rect 1563 650 1623 654
rect 1627 650 1647 654
rect 1651 650 1735 654
rect 1739 650 1831 654
rect 1835 650 1847 654
rect 1851 650 1919 654
rect 1923 650 1951 654
rect 1955 650 2007 654
rect 2011 650 2047 654
rect 2051 650 2087 654
rect 2091 650 2135 654
rect 2139 650 2167 654
rect 2171 650 2215 654
rect 2219 650 2239 654
rect 2243 650 2295 654
rect 2299 650 2311 654
rect 2315 650 2375 654
rect 2379 650 2383 654
rect 2387 650 2439 654
rect 2443 650 2503 654
rect 2507 650 2527 654
rect 1305 649 2527 650
rect 2533 649 2534 655
rect 96 613 97 619
rect 103 618 1311 619
rect 103 614 111 618
rect 115 614 207 618
rect 211 614 231 618
rect 235 614 303 618
rect 307 614 311 618
rect 315 614 391 618
rect 395 614 407 618
rect 411 614 471 618
rect 475 614 503 618
rect 507 614 543 618
rect 547 614 599 618
rect 603 614 607 618
rect 611 614 671 618
rect 675 614 687 618
rect 691 614 735 618
rect 739 614 767 618
rect 771 614 799 618
rect 803 614 847 618
rect 851 614 863 618
rect 867 614 927 618
rect 931 614 935 618
rect 939 614 1007 618
rect 1011 614 1087 618
rect 1091 614 1287 618
rect 1291 614 1311 618
rect 103 613 1311 614
rect 1317 613 1318 619
rect 1310 593 1311 599
rect 1317 598 2539 599
rect 1317 594 1327 598
rect 1331 594 1455 598
rect 1459 594 1495 598
rect 1499 594 1559 598
rect 1563 594 1575 598
rect 1579 594 1663 598
rect 1667 594 1671 598
rect 1675 594 1751 598
rect 1755 594 1775 598
rect 1779 594 1847 598
rect 1851 594 1879 598
rect 1883 594 1935 598
rect 1939 594 1983 598
rect 1987 594 2023 598
rect 2027 594 2087 598
rect 2091 594 2103 598
rect 2107 594 2183 598
rect 2187 594 2255 598
rect 2259 594 2279 598
rect 2283 594 2327 598
rect 2331 594 2375 598
rect 2379 594 2399 598
rect 2403 594 2455 598
rect 2459 594 2503 598
rect 2507 594 2539 598
rect 1317 593 2539 594
rect 2545 593 2546 599
rect 84 557 85 563
rect 91 562 1299 563
rect 91 558 111 562
rect 115 558 175 562
rect 179 558 191 562
rect 195 558 271 562
rect 275 558 287 562
rect 291 558 375 562
rect 379 558 391 562
rect 395 558 487 562
rect 491 558 583 562
rect 587 558 591 562
rect 595 558 671 562
rect 675 558 695 562
rect 699 558 751 562
rect 755 558 791 562
rect 795 558 831 562
rect 835 558 879 562
rect 883 558 911 562
rect 915 558 967 562
rect 971 558 991 562
rect 995 558 1055 562
rect 1059 558 1071 562
rect 1075 558 1151 562
rect 1155 558 1287 562
rect 1291 558 1299 562
rect 91 557 1299 558
rect 1305 557 1306 563
rect 1298 537 1299 543
rect 1305 542 2527 543
rect 1305 538 1327 542
rect 1331 538 1367 542
rect 1371 538 1439 542
rect 1443 538 1447 542
rect 1451 538 1527 542
rect 1531 538 1543 542
rect 1547 538 1615 542
rect 1619 538 1655 542
rect 1659 538 1711 542
rect 1715 538 1759 542
rect 1763 538 1799 542
rect 1803 538 1863 542
rect 1867 538 1887 542
rect 1891 538 1967 542
rect 1971 538 1975 542
rect 1979 538 2063 542
rect 2067 538 2071 542
rect 2075 538 2151 542
rect 2155 538 2167 542
rect 2171 538 2247 542
rect 2251 538 2263 542
rect 2267 538 2343 542
rect 2347 538 2359 542
rect 2363 538 2439 542
rect 2443 538 2503 542
rect 2507 538 2527 542
rect 1305 537 2527 538
rect 2533 537 2534 543
rect 96 501 97 507
rect 103 506 1311 507
rect 103 502 111 506
rect 115 502 151 506
rect 155 502 191 506
rect 195 502 247 506
rect 251 502 287 506
rect 291 502 367 506
rect 371 502 391 506
rect 395 502 487 506
rect 491 502 503 506
rect 507 502 607 506
rect 611 502 615 506
rect 619 502 711 506
rect 715 502 735 506
rect 739 502 807 506
rect 811 502 847 506
rect 851 502 895 506
rect 899 502 951 506
rect 955 502 983 506
rect 987 502 1055 506
rect 1059 502 1071 506
rect 1075 502 1159 506
rect 1163 502 1167 506
rect 1171 502 1239 506
rect 1243 502 1287 506
rect 1291 502 1311 506
rect 103 501 1311 502
rect 1317 501 1318 507
rect 2054 500 2060 501
rect 2270 500 2276 501
rect 2054 496 2055 500
rect 2059 496 2271 500
rect 2275 496 2276 500
rect 2054 495 2060 496
rect 2270 495 2276 496
rect 1310 481 1311 487
rect 1317 486 2539 487
rect 1317 482 1327 486
rect 1331 482 1367 486
rect 1371 482 1383 486
rect 1387 482 1431 486
rect 1435 482 1463 486
rect 1467 482 1519 486
rect 1523 482 1543 486
rect 1547 482 1615 486
rect 1619 482 1631 486
rect 1635 482 1711 486
rect 1715 482 1727 486
rect 1731 482 1815 486
rect 1819 482 1903 486
rect 1907 482 1927 486
rect 1931 482 1991 486
rect 1995 482 2055 486
rect 2059 482 2079 486
rect 2083 482 2167 486
rect 2171 482 2191 486
rect 2195 482 2263 486
rect 2267 482 2335 486
rect 2339 482 2359 486
rect 2363 482 2455 486
rect 2459 482 2503 486
rect 2507 482 2539 486
rect 1317 481 2539 482
rect 2545 481 2546 487
rect 84 445 85 451
rect 91 450 1299 451
rect 91 446 111 450
rect 115 446 135 450
rect 139 446 191 450
rect 195 446 231 450
rect 235 446 247 450
rect 251 446 303 450
rect 307 446 351 450
rect 355 446 383 450
rect 387 446 471 450
rect 475 446 567 450
rect 571 446 599 450
rect 603 446 671 450
rect 675 446 719 450
rect 723 446 783 450
rect 787 446 831 450
rect 835 446 895 450
rect 899 446 935 450
rect 939 446 1007 450
rect 1011 446 1039 450
rect 1043 446 1127 450
rect 1131 446 1143 450
rect 1147 446 1223 450
rect 1227 446 1287 450
rect 1291 446 1299 450
rect 91 445 1299 446
rect 1305 445 1306 451
rect 1298 425 1299 431
rect 1305 430 2527 431
rect 1305 426 1327 430
rect 1331 426 1351 430
rect 1355 426 1415 430
rect 1419 426 1423 430
rect 1427 426 1503 430
rect 1507 426 1511 430
rect 1515 426 1599 430
rect 1603 426 1679 430
rect 1683 426 1695 430
rect 1699 426 1775 430
rect 1779 426 1799 430
rect 1803 426 1887 430
rect 1891 426 1911 430
rect 1915 426 2015 430
rect 2019 426 2039 430
rect 2043 426 2159 430
rect 2163 426 2175 430
rect 2179 426 2311 430
rect 2315 426 2319 430
rect 2323 426 2439 430
rect 2443 426 2503 430
rect 2507 426 2527 430
rect 1305 425 2527 426
rect 2533 425 2534 431
rect 96 385 97 391
rect 103 390 1311 391
rect 103 386 111 390
rect 115 386 151 390
rect 155 386 207 390
rect 211 386 263 390
rect 267 386 279 390
rect 283 386 319 390
rect 323 386 359 390
rect 363 386 399 390
rect 403 386 431 390
rect 435 386 487 390
rect 491 386 511 390
rect 515 386 583 390
rect 587 386 591 390
rect 595 386 671 390
rect 675 386 687 390
rect 691 386 751 390
rect 755 386 799 390
rect 803 386 823 390
rect 827 386 895 390
rect 899 386 911 390
rect 915 386 967 390
rect 971 386 1023 390
rect 1027 386 1039 390
rect 1043 386 1111 390
rect 1115 386 1143 390
rect 1147 386 1183 390
rect 1187 386 1239 390
rect 1243 386 1287 390
rect 1291 386 1311 390
rect 103 385 1311 386
rect 1317 385 1318 391
rect 1310 369 1311 375
rect 1317 374 2539 375
rect 1317 370 1327 374
rect 1331 370 1367 374
rect 1371 370 1439 374
rect 1443 370 1527 374
rect 1531 370 1615 374
rect 1619 370 1679 374
rect 1683 370 1695 374
rect 1699 370 1735 374
rect 1739 370 1791 374
rect 1795 370 1807 374
rect 1811 370 1903 374
rect 1907 370 2023 374
rect 2027 370 2031 374
rect 2035 370 2159 374
rect 2163 370 2175 374
rect 2179 370 2303 374
rect 2307 370 2327 374
rect 2331 370 2455 374
rect 2459 370 2503 374
rect 2507 370 2539 374
rect 1317 369 2539 370
rect 2545 369 2546 375
rect 84 325 85 331
rect 91 330 1299 331
rect 91 326 111 330
rect 115 326 135 330
rect 139 326 191 330
rect 195 326 199 330
rect 203 326 263 330
rect 267 326 287 330
rect 291 326 343 330
rect 347 326 375 330
rect 379 326 415 330
rect 419 326 455 330
rect 459 326 495 330
rect 499 326 543 330
rect 547 326 575 330
rect 579 326 631 330
rect 635 326 655 330
rect 659 326 727 330
rect 731 326 735 330
rect 739 326 807 330
rect 811 326 823 330
rect 827 326 879 330
rect 883 326 927 330
rect 931 326 951 330
rect 955 326 1023 330
rect 1027 326 1031 330
rect 1035 326 1095 330
rect 1099 326 1135 330
rect 1139 326 1167 330
rect 1171 326 1223 330
rect 1227 326 1287 330
rect 1291 326 1299 330
rect 91 325 1299 326
rect 1305 325 1306 331
rect 1298 323 1306 325
rect 1298 317 1299 323
rect 1305 322 2527 323
rect 1305 318 1327 322
rect 1331 318 1351 322
rect 1355 318 1431 322
rect 1435 318 1527 322
rect 1531 318 1623 322
rect 1627 318 1663 322
rect 1667 318 1711 322
rect 1715 318 1719 322
rect 1723 318 1791 322
rect 1795 318 1807 322
rect 1811 318 1887 322
rect 1891 318 1911 322
rect 1915 318 2007 322
rect 2011 318 2023 322
rect 2027 318 2143 322
rect 2147 318 2151 322
rect 2155 318 2287 322
rect 2291 318 2423 322
rect 2427 318 2439 322
rect 2443 318 2503 322
rect 2507 318 2527 322
rect 1305 317 2527 318
rect 2533 317 2534 323
rect 96 265 97 271
rect 103 270 1311 271
rect 103 266 111 270
rect 115 266 151 270
rect 155 266 215 270
rect 219 266 231 270
rect 235 266 303 270
rect 307 266 327 270
rect 331 266 391 270
rect 395 266 423 270
rect 427 266 471 270
rect 475 266 519 270
rect 523 266 559 270
rect 563 266 615 270
rect 619 266 647 270
rect 651 266 711 270
rect 715 266 743 270
rect 747 266 807 270
rect 811 266 839 270
rect 843 266 903 270
rect 907 266 943 270
rect 947 266 1007 270
rect 1011 266 1047 270
rect 1051 266 1111 270
rect 1115 266 1151 270
rect 1155 266 1215 270
rect 1219 266 1239 270
rect 1243 266 1287 270
rect 1291 266 1311 270
rect 103 265 1311 266
rect 1317 267 1318 271
rect 1317 266 2546 267
rect 1317 265 1327 266
rect 1310 262 1327 265
rect 1331 262 1367 266
rect 1371 262 1439 266
rect 1443 262 1447 266
rect 1451 262 1535 266
rect 1539 262 1543 266
rect 1547 262 1631 266
rect 1635 262 1639 266
rect 1643 262 1727 266
rect 1731 262 1815 266
rect 1819 262 1823 266
rect 1827 262 1903 266
rect 1907 262 1927 266
rect 1931 262 1999 266
rect 2003 262 2039 266
rect 2043 262 2103 266
rect 2107 262 2167 266
rect 2171 262 2215 266
rect 2219 262 2303 266
rect 2307 262 2335 266
rect 2339 262 2439 266
rect 2443 262 2455 266
rect 2459 262 2503 266
rect 2507 262 2546 266
rect 1310 261 2546 262
rect 84 205 85 211
rect 91 210 1299 211
rect 91 206 111 210
rect 115 206 135 210
rect 139 206 159 210
rect 163 206 215 210
rect 219 206 239 210
rect 243 206 311 210
rect 315 206 327 210
rect 331 206 407 210
rect 411 206 415 210
rect 419 206 503 210
rect 507 206 511 210
rect 515 206 599 210
rect 603 206 607 210
rect 611 206 695 210
rect 699 206 783 210
rect 787 206 791 210
rect 795 206 871 210
rect 875 206 887 210
rect 891 206 959 210
rect 963 206 991 210
rect 995 206 1047 210
rect 1051 206 1095 210
rect 1099 206 1135 210
rect 1139 206 1199 210
rect 1203 206 1287 210
rect 1291 206 1299 210
rect 91 205 1299 206
rect 1305 210 2534 211
rect 1305 206 1327 210
rect 1331 206 1351 210
rect 1355 206 1391 210
rect 1395 206 1423 210
rect 1427 206 1495 210
rect 1499 206 1519 210
rect 1523 206 1599 210
rect 1603 206 1615 210
rect 1619 206 1711 210
rect 1715 206 1799 210
rect 1803 206 1815 210
rect 1819 206 1887 210
rect 1891 206 1919 210
rect 1923 206 1983 210
rect 1987 206 2015 210
rect 2019 206 2087 210
rect 2091 206 2111 210
rect 2115 206 2199 210
rect 2203 206 2287 210
rect 2291 206 2319 210
rect 2323 206 2375 210
rect 2379 206 2439 210
rect 2443 206 2503 210
rect 2507 206 2534 210
rect 1305 205 2534 206
rect 96 133 97 139
rect 103 138 1311 139
rect 103 134 111 138
rect 115 134 151 138
rect 155 134 175 138
rect 179 134 207 138
rect 211 134 255 138
rect 259 134 263 138
rect 267 134 319 138
rect 323 134 343 138
rect 347 134 375 138
rect 379 134 431 138
rect 435 134 487 138
rect 491 134 527 138
rect 531 134 551 138
rect 555 134 623 138
rect 627 134 687 138
rect 691 134 711 138
rect 715 134 751 138
rect 755 134 799 138
rect 803 134 815 138
rect 819 134 879 138
rect 883 134 887 138
rect 891 134 943 138
rect 947 134 975 138
rect 979 134 1007 138
rect 1011 134 1063 138
rect 1067 134 1071 138
rect 1075 134 1135 138
rect 1139 134 1151 138
rect 1155 134 1199 138
rect 1203 134 1287 138
rect 1291 134 1311 138
rect 103 133 1311 134
rect 1317 138 2546 139
rect 1317 134 1327 138
rect 1331 134 1367 138
rect 1371 134 1407 138
rect 1411 134 1423 138
rect 1427 134 1479 138
rect 1483 134 1511 138
rect 1515 134 1535 138
rect 1539 134 1591 138
rect 1595 134 1615 138
rect 1619 134 1647 138
rect 1651 134 1703 138
rect 1707 134 1727 138
rect 1731 134 1759 138
rect 1763 134 1815 138
rect 1819 134 1831 138
rect 1835 134 1871 138
rect 1875 134 1927 138
rect 1931 134 1935 138
rect 1939 134 1983 138
rect 1987 134 2031 138
rect 2035 134 2039 138
rect 2043 134 2095 138
rect 2099 134 2127 138
rect 2131 134 2159 138
rect 2163 134 2215 138
rect 2219 134 2223 138
rect 2227 134 2287 138
rect 2291 134 2303 138
rect 2307 134 2343 138
rect 2347 134 2391 138
rect 2395 134 2399 138
rect 2403 134 2455 138
rect 2459 134 2503 138
rect 2507 134 2546 138
rect 1317 133 2546 134
rect 84 81 85 87
rect 91 86 1299 87
rect 91 82 111 86
rect 115 82 135 86
rect 139 82 191 86
rect 195 82 247 86
rect 251 82 303 86
rect 307 82 359 86
rect 363 82 415 86
rect 419 82 471 86
rect 475 82 535 86
rect 539 82 607 86
rect 611 82 671 86
rect 675 82 735 86
rect 739 82 799 86
rect 803 82 863 86
rect 867 82 927 86
rect 931 82 991 86
rect 995 82 1055 86
rect 1059 82 1119 86
rect 1123 82 1183 86
rect 1187 82 1287 86
rect 1291 82 1299 86
rect 91 81 1299 82
rect 1305 86 2534 87
rect 1305 82 1327 86
rect 1331 82 1351 86
rect 1355 82 1407 86
rect 1411 82 1463 86
rect 1467 82 1519 86
rect 1523 82 1575 86
rect 1579 82 1631 86
rect 1635 82 1687 86
rect 1691 82 1743 86
rect 1747 82 1799 86
rect 1803 82 1855 86
rect 1859 82 1911 86
rect 1915 82 1967 86
rect 1971 82 2023 86
rect 2027 82 2079 86
rect 2083 82 2143 86
rect 2147 82 2207 86
rect 2211 82 2271 86
rect 2275 82 2327 86
rect 2331 82 2383 86
rect 2387 82 2439 86
rect 2443 82 2503 86
rect 2507 82 2534 86
rect 1305 81 2534 82
<< m5c >>
rect 97 2577 103 2583
rect 1311 2577 1317 2583
rect 1311 2553 1317 2559
rect 2539 2553 2545 2559
rect 85 2525 91 2531
rect 1299 2525 1305 2531
rect 1299 2493 1305 2499
rect 2527 2493 2533 2499
rect 97 2473 103 2479
rect 1311 2473 1317 2479
rect 1311 2433 1317 2439
rect 2539 2433 2545 2439
rect 85 2417 91 2423
rect 1299 2417 1305 2423
rect 1299 2375 1305 2381
rect 2527 2373 2533 2379
rect 97 2365 103 2371
rect 1311 2365 1317 2371
rect 1311 2317 1317 2323
rect 2539 2317 2545 2323
rect 85 2309 91 2315
rect 1299 2309 1305 2315
rect 1299 2265 1305 2271
rect 2527 2265 2533 2271
rect 97 2253 103 2259
rect 1311 2253 1317 2259
rect 1311 2209 1317 2215
rect 2539 2209 2545 2215
rect 85 2197 91 2203
rect 1299 2197 1305 2203
rect 1299 2155 1305 2161
rect 97 2145 103 2151
rect 1311 2145 1317 2151
rect 2527 2145 2533 2151
rect 85 2093 91 2099
rect 1299 2093 1305 2099
rect 1311 2081 1317 2087
rect 2539 2081 2545 2087
rect 1299 2047 1305 2053
rect 97 2037 103 2043
rect 1311 2037 1317 2043
rect 2527 2029 2533 2035
rect 85 1981 91 1987
rect 1299 1981 1305 1987
rect 1311 1973 1317 1979
rect 2539 1973 2545 1979
rect 1299 1931 1305 1937
rect 97 1921 103 1927
rect 1311 1921 1317 1927
rect 2527 1917 2533 1923
rect 85 1869 91 1875
rect 1299 1869 1305 1875
rect 1311 1865 1317 1871
rect 2539 1865 2545 1871
rect 1299 1819 1305 1825
rect 97 1809 103 1815
rect 1311 1809 1317 1815
rect 2527 1809 2533 1815
rect 85 1753 91 1759
rect 1299 1753 1305 1759
rect 1311 1753 1317 1759
rect 2539 1753 2545 1759
rect 1299 1707 1305 1713
rect 97 1697 103 1703
rect 1311 1697 1317 1703
rect 2527 1701 2533 1707
rect 85 1645 91 1651
rect 1299 1645 1305 1651
rect 1311 1641 1317 1647
rect 2539 1641 2545 1647
rect 1299 1603 1305 1609
rect 97 1593 103 1599
rect 1311 1593 1317 1599
rect 2527 1585 2533 1591
rect 85 1533 91 1539
rect 1299 1533 1305 1539
rect 1311 1533 1317 1539
rect 2539 1533 2545 1539
rect 1299 1491 1305 1497
rect 97 1481 103 1487
rect 1311 1481 1317 1487
rect 2527 1477 2533 1483
rect 85 1429 91 1435
rect 1299 1429 1305 1435
rect 1311 1421 1317 1427
rect 2539 1421 2545 1427
rect 97 1377 103 1383
rect 1311 1377 1317 1383
rect 1299 1365 1305 1371
rect 2527 1365 2533 1371
rect 85 1325 91 1331
rect 1299 1325 1305 1331
rect 1311 1305 1317 1311
rect 2539 1305 2545 1311
rect 97 1273 103 1279
rect 1311 1273 1317 1279
rect 1299 1237 1305 1243
rect 2527 1237 2533 1243
rect 85 1221 91 1227
rect 1299 1221 1305 1227
rect 1311 1185 1317 1191
rect 2539 1185 2545 1191
rect 97 1165 103 1171
rect 1311 1165 1317 1171
rect 1299 1129 1305 1135
rect 2527 1129 2533 1135
rect 85 1109 91 1115
rect 1299 1109 1305 1115
rect 1311 1069 1317 1075
rect 2539 1069 2545 1075
rect 97 1053 103 1059
rect 1311 1053 1317 1059
rect 1299 1009 1305 1015
rect 2527 1009 2533 1015
rect 85 997 91 1003
rect 1299 997 1305 1003
rect 97 945 103 951
rect 1311 945 1317 951
rect 85 889 91 895
rect 1299 889 1305 895
rect 1299 881 1305 887
rect 2527 881 2533 887
rect 97 833 103 839
rect 1311 833 1317 839
rect 1311 821 1317 827
rect 2539 821 2545 827
rect 85 777 91 783
rect 1299 777 1305 783
rect 1299 765 1305 771
rect 2527 765 2533 771
rect 97 721 103 727
rect 1311 721 1317 727
rect 1311 709 1317 715
rect 2539 709 2545 715
rect 85 669 91 675
rect 1299 669 1305 675
rect 1299 649 1305 655
rect 2527 649 2533 655
rect 97 613 103 619
rect 1311 613 1317 619
rect 1311 593 1317 599
rect 2539 593 2545 599
rect 85 557 91 563
rect 1299 557 1305 563
rect 1299 537 1305 543
rect 2527 537 2533 543
rect 97 501 103 507
rect 1311 501 1317 507
rect 1311 481 1317 487
rect 2539 481 2545 487
rect 85 445 91 451
rect 1299 445 1305 451
rect 1299 425 1305 431
rect 2527 425 2533 431
rect 97 385 103 391
rect 1311 385 1317 391
rect 1311 369 1317 375
rect 2539 369 2545 375
rect 85 325 91 331
rect 1299 325 1305 331
rect 1299 317 1305 323
rect 2527 317 2533 323
rect 97 265 103 271
rect 1311 265 1317 271
rect 85 205 91 211
rect 1299 205 1305 211
rect 97 133 103 139
rect 1311 133 1317 139
rect 85 81 91 87
rect 1299 81 1305 87
<< m5 >>
rect 84 2531 92 2592
rect 84 2525 85 2531
rect 91 2525 92 2531
rect 84 2423 92 2525
rect 84 2417 85 2423
rect 91 2417 92 2423
rect 84 2315 92 2417
rect 84 2309 85 2315
rect 91 2309 92 2315
rect 84 2203 92 2309
rect 84 2197 85 2203
rect 91 2197 92 2203
rect 84 2099 92 2197
rect 84 2093 85 2099
rect 91 2093 92 2099
rect 84 1987 92 2093
rect 84 1981 85 1987
rect 91 1981 92 1987
rect 84 1875 92 1981
rect 84 1869 85 1875
rect 91 1869 92 1875
rect 84 1759 92 1869
rect 84 1753 85 1759
rect 91 1753 92 1759
rect 84 1651 92 1753
rect 84 1645 85 1651
rect 91 1645 92 1651
rect 84 1539 92 1645
rect 84 1533 85 1539
rect 91 1533 92 1539
rect 84 1435 92 1533
rect 84 1429 85 1435
rect 91 1429 92 1435
rect 84 1331 92 1429
rect 84 1325 85 1331
rect 91 1325 92 1331
rect 84 1227 92 1325
rect 84 1221 85 1227
rect 91 1221 92 1227
rect 84 1115 92 1221
rect 84 1109 85 1115
rect 91 1109 92 1115
rect 84 1003 92 1109
rect 84 997 85 1003
rect 91 997 92 1003
rect 84 895 92 997
rect 84 889 85 895
rect 91 889 92 895
rect 84 783 92 889
rect 84 777 85 783
rect 91 777 92 783
rect 84 675 92 777
rect 84 669 85 675
rect 91 669 92 675
rect 84 563 92 669
rect 84 557 85 563
rect 91 557 92 563
rect 84 451 92 557
rect 84 445 85 451
rect 91 445 92 451
rect 84 331 92 445
rect 84 325 85 331
rect 91 325 92 331
rect 84 211 92 325
rect 84 205 85 211
rect 91 205 92 211
rect 84 87 92 205
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 2583 104 2592
rect 96 2577 97 2583
rect 103 2577 104 2583
rect 96 2479 104 2577
rect 96 2473 97 2479
rect 103 2473 104 2479
rect 96 2371 104 2473
rect 96 2365 97 2371
rect 103 2365 104 2371
rect 96 2259 104 2365
rect 96 2253 97 2259
rect 103 2253 104 2259
rect 96 2151 104 2253
rect 96 2145 97 2151
rect 103 2145 104 2151
rect 96 2043 104 2145
rect 96 2037 97 2043
rect 103 2037 104 2043
rect 96 1927 104 2037
rect 96 1921 97 1927
rect 103 1921 104 1927
rect 96 1815 104 1921
rect 96 1809 97 1815
rect 103 1809 104 1815
rect 96 1703 104 1809
rect 96 1697 97 1703
rect 103 1697 104 1703
rect 96 1599 104 1697
rect 96 1593 97 1599
rect 103 1593 104 1599
rect 96 1487 104 1593
rect 96 1481 97 1487
rect 103 1481 104 1487
rect 96 1383 104 1481
rect 96 1377 97 1383
rect 103 1377 104 1383
rect 96 1279 104 1377
rect 96 1273 97 1279
rect 103 1273 104 1279
rect 96 1171 104 1273
rect 96 1165 97 1171
rect 103 1165 104 1171
rect 96 1059 104 1165
rect 96 1053 97 1059
rect 103 1053 104 1059
rect 96 951 104 1053
rect 96 945 97 951
rect 103 945 104 951
rect 96 839 104 945
rect 96 833 97 839
rect 103 833 104 839
rect 96 727 104 833
rect 96 721 97 727
rect 103 721 104 727
rect 96 619 104 721
rect 96 613 97 619
rect 103 613 104 619
rect 96 507 104 613
rect 96 501 97 507
rect 103 501 104 507
rect 96 391 104 501
rect 96 385 97 391
rect 103 385 104 391
rect 96 271 104 385
rect 96 265 97 271
rect 103 265 104 271
rect 96 139 104 265
rect 96 133 97 139
rect 103 133 104 139
rect 96 72 104 133
rect 1298 2531 1306 2592
rect 1298 2525 1299 2531
rect 1305 2525 1306 2531
rect 1298 2499 1306 2525
rect 1298 2493 1299 2499
rect 1305 2493 1306 2499
rect 1298 2423 1306 2493
rect 1298 2417 1299 2423
rect 1305 2417 1306 2423
rect 1298 2381 1306 2417
rect 1298 2375 1299 2381
rect 1305 2375 1306 2381
rect 1298 2315 1306 2375
rect 1298 2309 1299 2315
rect 1305 2309 1306 2315
rect 1298 2271 1306 2309
rect 1298 2265 1299 2271
rect 1305 2265 1306 2271
rect 1298 2203 1306 2265
rect 1298 2197 1299 2203
rect 1305 2197 1306 2203
rect 1298 2161 1306 2197
rect 1298 2155 1299 2161
rect 1305 2155 1306 2161
rect 1298 2099 1306 2155
rect 1298 2093 1299 2099
rect 1305 2093 1306 2099
rect 1298 2053 1306 2093
rect 1298 2047 1299 2053
rect 1305 2047 1306 2053
rect 1298 1987 1306 2047
rect 1298 1981 1299 1987
rect 1305 1981 1306 1987
rect 1298 1937 1306 1981
rect 1298 1931 1299 1937
rect 1305 1931 1306 1937
rect 1298 1875 1306 1931
rect 1298 1869 1299 1875
rect 1305 1869 1306 1875
rect 1298 1825 1306 1869
rect 1298 1819 1299 1825
rect 1305 1819 1306 1825
rect 1298 1759 1306 1819
rect 1298 1753 1299 1759
rect 1305 1753 1306 1759
rect 1298 1713 1306 1753
rect 1298 1707 1299 1713
rect 1305 1707 1306 1713
rect 1298 1651 1306 1707
rect 1298 1645 1299 1651
rect 1305 1645 1306 1651
rect 1298 1609 1306 1645
rect 1298 1603 1299 1609
rect 1305 1603 1306 1609
rect 1298 1539 1306 1603
rect 1298 1533 1299 1539
rect 1305 1533 1306 1539
rect 1298 1497 1306 1533
rect 1298 1491 1299 1497
rect 1305 1491 1306 1497
rect 1298 1435 1306 1491
rect 1298 1429 1299 1435
rect 1305 1429 1306 1435
rect 1298 1371 1306 1429
rect 1298 1365 1299 1371
rect 1305 1365 1306 1371
rect 1298 1331 1306 1365
rect 1298 1325 1299 1331
rect 1305 1325 1306 1331
rect 1298 1243 1306 1325
rect 1298 1237 1299 1243
rect 1305 1237 1306 1243
rect 1298 1227 1306 1237
rect 1298 1221 1299 1227
rect 1305 1221 1306 1227
rect 1298 1135 1306 1221
rect 1298 1129 1299 1135
rect 1305 1129 1306 1135
rect 1298 1115 1306 1129
rect 1298 1109 1299 1115
rect 1305 1109 1306 1115
rect 1298 1015 1306 1109
rect 1298 1009 1299 1015
rect 1305 1009 1306 1015
rect 1298 1003 1306 1009
rect 1298 997 1299 1003
rect 1305 997 1306 1003
rect 1298 895 1306 997
rect 1298 889 1299 895
rect 1305 889 1306 895
rect 1298 887 1306 889
rect 1298 881 1299 887
rect 1305 881 1306 887
rect 1298 783 1306 881
rect 1298 777 1299 783
rect 1305 777 1306 783
rect 1298 771 1306 777
rect 1298 765 1299 771
rect 1305 765 1306 771
rect 1298 675 1306 765
rect 1298 669 1299 675
rect 1305 669 1306 675
rect 1298 655 1306 669
rect 1298 649 1299 655
rect 1305 649 1306 655
rect 1298 563 1306 649
rect 1298 557 1299 563
rect 1305 557 1306 563
rect 1298 543 1306 557
rect 1298 537 1299 543
rect 1305 537 1306 543
rect 1298 451 1306 537
rect 1298 445 1299 451
rect 1305 445 1306 451
rect 1298 431 1306 445
rect 1298 425 1299 431
rect 1305 425 1306 431
rect 1298 331 1306 425
rect 1298 325 1299 331
rect 1305 325 1306 331
rect 1298 323 1306 325
rect 1298 317 1299 323
rect 1305 317 1306 323
rect 1298 211 1306 317
rect 1298 205 1299 211
rect 1305 205 1306 211
rect 1298 87 1306 205
rect 1298 81 1299 87
rect 1305 81 1306 87
rect 1298 72 1306 81
rect 1310 2583 1318 2592
rect 1310 2577 1311 2583
rect 1317 2577 1318 2583
rect 1310 2559 1318 2577
rect 1310 2553 1311 2559
rect 1317 2553 1318 2559
rect 1310 2479 1318 2553
rect 1310 2473 1311 2479
rect 1317 2473 1318 2479
rect 1310 2439 1318 2473
rect 1310 2433 1311 2439
rect 1317 2433 1318 2439
rect 1310 2371 1318 2433
rect 1310 2365 1311 2371
rect 1317 2365 1318 2371
rect 1310 2323 1318 2365
rect 1310 2317 1311 2323
rect 1317 2317 1318 2323
rect 1310 2259 1318 2317
rect 1310 2253 1311 2259
rect 1317 2253 1318 2259
rect 1310 2215 1318 2253
rect 1310 2209 1311 2215
rect 1317 2209 1318 2215
rect 1310 2151 1318 2209
rect 1310 2145 1311 2151
rect 1317 2145 1318 2151
rect 1310 2087 1318 2145
rect 1310 2081 1311 2087
rect 1317 2081 1318 2087
rect 1310 2043 1318 2081
rect 1310 2037 1311 2043
rect 1317 2037 1318 2043
rect 1310 1979 1318 2037
rect 1310 1973 1311 1979
rect 1317 1973 1318 1979
rect 1310 1927 1318 1973
rect 1310 1921 1311 1927
rect 1317 1921 1318 1927
rect 1310 1871 1318 1921
rect 1310 1865 1311 1871
rect 1317 1865 1318 1871
rect 1310 1815 1318 1865
rect 1310 1809 1311 1815
rect 1317 1809 1318 1815
rect 1310 1759 1318 1809
rect 1310 1753 1311 1759
rect 1317 1753 1318 1759
rect 1310 1703 1318 1753
rect 1310 1697 1311 1703
rect 1317 1697 1318 1703
rect 1310 1647 1318 1697
rect 1310 1641 1311 1647
rect 1317 1641 1318 1647
rect 1310 1599 1318 1641
rect 1310 1593 1311 1599
rect 1317 1593 1318 1599
rect 1310 1539 1318 1593
rect 1310 1533 1311 1539
rect 1317 1533 1318 1539
rect 1310 1487 1318 1533
rect 1310 1481 1311 1487
rect 1317 1481 1318 1487
rect 1310 1427 1318 1481
rect 1310 1421 1311 1427
rect 1317 1421 1318 1427
rect 1310 1383 1318 1421
rect 1310 1377 1311 1383
rect 1317 1377 1318 1383
rect 1310 1311 1318 1377
rect 1310 1305 1311 1311
rect 1317 1305 1318 1311
rect 1310 1279 1318 1305
rect 1310 1273 1311 1279
rect 1317 1273 1318 1279
rect 1310 1191 1318 1273
rect 1310 1185 1311 1191
rect 1317 1185 1318 1191
rect 1310 1171 1318 1185
rect 1310 1165 1311 1171
rect 1317 1165 1318 1171
rect 1310 1075 1318 1165
rect 1310 1069 1311 1075
rect 1317 1069 1318 1075
rect 1310 1059 1318 1069
rect 1310 1053 1311 1059
rect 1317 1053 1318 1059
rect 1310 951 1318 1053
rect 1310 945 1311 951
rect 1317 945 1318 951
rect 1310 839 1318 945
rect 1310 833 1311 839
rect 1317 833 1318 839
rect 1310 827 1318 833
rect 1310 821 1311 827
rect 1317 821 1318 827
rect 1310 727 1318 821
rect 1310 721 1311 727
rect 1317 721 1318 727
rect 1310 715 1318 721
rect 1310 709 1311 715
rect 1317 709 1318 715
rect 1310 619 1318 709
rect 1310 613 1311 619
rect 1317 613 1318 619
rect 1310 599 1318 613
rect 1310 593 1311 599
rect 1317 593 1318 599
rect 1310 507 1318 593
rect 1310 501 1311 507
rect 1317 501 1318 507
rect 1310 487 1318 501
rect 1310 481 1311 487
rect 1317 481 1318 487
rect 1310 391 1318 481
rect 1310 385 1311 391
rect 1317 385 1318 391
rect 1310 375 1318 385
rect 1310 369 1311 375
rect 1317 369 1318 375
rect 1310 271 1318 369
rect 1310 265 1311 271
rect 1317 265 1318 271
rect 1310 139 1318 265
rect 1310 133 1311 139
rect 1317 133 1318 139
rect 1310 72 1318 133
rect 2526 2499 2534 2592
rect 2526 2493 2527 2499
rect 2533 2493 2534 2499
rect 2526 2379 2534 2493
rect 2526 2373 2527 2379
rect 2533 2373 2534 2379
rect 2526 2271 2534 2373
rect 2526 2265 2527 2271
rect 2533 2265 2534 2271
rect 2526 2151 2534 2265
rect 2526 2145 2527 2151
rect 2533 2145 2534 2151
rect 2526 2035 2534 2145
rect 2526 2029 2527 2035
rect 2533 2029 2534 2035
rect 2526 1923 2534 2029
rect 2526 1917 2527 1923
rect 2533 1917 2534 1923
rect 2526 1815 2534 1917
rect 2526 1809 2527 1815
rect 2533 1809 2534 1815
rect 2526 1707 2534 1809
rect 2526 1701 2527 1707
rect 2533 1701 2534 1707
rect 2526 1591 2534 1701
rect 2526 1585 2527 1591
rect 2533 1585 2534 1591
rect 2526 1483 2534 1585
rect 2526 1477 2527 1483
rect 2533 1477 2534 1483
rect 2526 1371 2534 1477
rect 2526 1365 2527 1371
rect 2533 1365 2534 1371
rect 2526 1243 2534 1365
rect 2526 1237 2527 1243
rect 2533 1237 2534 1243
rect 2526 1135 2534 1237
rect 2526 1129 2527 1135
rect 2533 1129 2534 1135
rect 2526 1015 2534 1129
rect 2526 1009 2527 1015
rect 2533 1009 2534 1015
rect 2526 887 2534 1009
rect 2526 881 2527 887
rect 2533 881 2534 887
rect 2526 771 2534 881
rect 2526 765 2527 771
rect 2533 765 2534 771
rect 2526 655 2534 765
rect 2526 649 2527 655
rect 2533 649 2534 655
rect 2526 543 2534 649
rect 2526 537 2527 543
rect 2533 537 2534 543
rect 2526 431 2534 537
rect 2526 425 2527 431
rect 2533 425 2534 431
rect 2526 323 2534 425
rect 2526 317 2527 323
rect 2533 317 2534 323
rect 2526 72 2534 317
rect 2538 2559 2546 2592
rect 2538 2553 2539 2559
rect 2545 2553 2546 2559
rect 2538 2439 2546 2553
rect 2538 2433 2539 2439
rect 2545 2433 2546 2439
rect 2538 2323 2546 2433
rect 2538 2317 2539 2323
rect 2545 2317 2546 2323
rect 2538 2215 2546 2317
rect 2538 2209 2539 2215
rect 2545 2209 2546 2215
rect 2538 2087 2546 2209
rect 2538 2081 2539 2087
rect 2545 2081 2546 2087
rect 2538 1979 2546 2081
rect 2538 1973 2539 1979
rect 2545 1973 2546 1979
rect 2538 1871 2546 1973
rect 2538 1865 2539 1871
rect 2545 1865 2546 1871
rect 2538 1759 2546 1865
rect 2538 1753 2539 1759
rect 2545 1753 2546 1759
rect 2538 1647 2546 1753
rect 2538 1641 2539 1647
rect 2545 1641 2546 1647
rect 2538 1539 2546 1641
rect 2538 1533 2539 1539
rect 2545 1533 2546 1539
rect 2538 1427 2546 1533
rect 2538 1421 2539 1427
rect 2545 1421 2546 1427
rect 2538 1311 2546 1421
rect 2538 1305 2539 1311
rect 2545 1305 2546 1311
rect 2538 1191 2546 1305
rect 2538 1185 2539 1191
rect 2545 1185 2546 1191
rect 2538 1075 2546 1185
rect 2538 1069 2539 1075
rect 2545 1069 2546 1075
rect 2538 827 2546 1069
rect 2538 821 2539 827
rect 2545 821 2546 827
rect 2538 715 2546 821
rect 2538 709 2539 715
rect 2545 709 2546 715
rect 2538 599 2546 709
rect 2538 593 2539 599
rect 2545 593 2546 599
rect 2538 487 2546 593
rect 2538 481 2539 487
rect 2545 481 2546 487
rect 2538 375 2546 481
rect 2538 369 2539 375
rect 2545 369 2546 375
rect 2538 72 2546 369
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__175
timestamp 1731220663
transform 1 0 2496 0 1 2508
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220663
transform 1 0 1320 0 1 2508
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220663
transform 1 0 2496 0 -1 2492
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220663
transform 1 0 1320 0 -1 2492
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220663
transform 1 0 2496 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220663
transform 1 0 1320 0 1 2388
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220663
transform 1 0 2496 0 -1 2372
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220663
transform 1 0 1320 0 -1 2372
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220663
transform 1 0 2496 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220663
transform 1 0 1320 0 1 2272
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220663
transform 1 0 2496 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220663
transform 1 0 1320 0 -1 2264
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220663
transform 1 0 2496 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220663
transform 1 0 1320 0 1 2164
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220663
transform 1 0 2496 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220663
transform 1 0 1320 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220663
transform 1 0 2496 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220663
transform 1 0 1320 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220663
transform 1 0 2496 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220663
transform 1 0 1320 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220663
transform 1 0 2496 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220663
transform 1 0 1320 0 1 1928
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220663
transform 1 0 2496 0 -1 1916
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220663
transform 1 0 1320 0 -1 1916
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220663
transform 1 0 2496 0 1 1820
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220663
transform 1 0 1320 0 1 1820
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220663
transform 1 0 2496 0 -1 1808
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220663
transform 1 0 1320 0 -1 1808
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220663
transform 1 0 2496 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220663
transform 1 0 1320 0 1 1708
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220663
transform 1 0 2496 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220663
transform 1 0 1320 0 -1 1700
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220663
transform 1 0 2496 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220663
transform 1 0 1320 0 1 1596
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220663
transform 1 0 2496 0 -1 1584
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220663
transform 1 0 1320 0 -1 1584
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220663
transform 1 0 2496 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220663
transform 1 0 1320 0 1 1488
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220663
transform 1 0 2496 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220663
transform 1 0 1320 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220663
transform 1 0 2496 0 1 1376
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220663
transform 1 0 1320 0 1 1376
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220663
transform 1 0 2496 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220663
transform 1 0 1320 0 -1 1364
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220663
transform 1 0 2496 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220663
transform 1 0 1320 0 1 1260
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220663
transform 1 0 2496 0 -1 1236
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220663
transform 1 0 1320 0 -1 1236
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220663
transform 1 0 2496 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220663
transform 1 0 1320 0 1 1140
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220663
transform 1 0 2496 0 -1 1128
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220663
transform 1 0 1320 0 -1 1128
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220663
transform 1 0 2496 0 1 1024
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220663
transform 1 0 1320 0 1 1024
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220663
transform 1 0 2496 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220663
transform 1 0 1320 0 -1 1008
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220663
transform 1 0 2496 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220663
transform 1 0 1320 0 1 896
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220663
transform 1 0 2496 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220663
transform 1 0 1320 0 -1 880
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220663
transform 1 0 2496 0 1 776
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220663
transform 1 0 1320 0 1 776
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220663
transform 1 0 2496 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220663
transform 1 0 1320 0 -1 764
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220663
transform 1 0 2496 0 1 664
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220663
transform 1 0 1320 0 1 664
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220663
transform 1 0 2496 0 -1 648
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220663
transform 1 0 1320 0 -1 648
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220663
transform 1 0 2496 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220663
transform 1 0 1320 0 1 548
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220663
transform 1 0 2496 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220663
transform 1 0 1320 0 -1 536
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220663
transform 1 0 2496 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220663
transform 1 0 1320 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220663
transform 1 0 2496 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220663
transform 1 0 1320 0 -1 424
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220663
transform 1 0 2496 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220663
transform 1 0 1320 0 1 324
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220663
transform 1 0 2496 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220663
transform 1 0 1320 0 -1 316
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220663
transform 1 0 2496 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220663
transform 1 0 1320 0 1 216
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220663
transform 1 0 2496 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220663
transform 1 0 1320 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220663
transform 1 0 2496 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220663
transform 1 0 1320 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220663
transform 1 0 1280 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220663
transform 1 0 104 0 1 2532
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220663
transform 1 0 1280 0 -1 2524
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220663
transform 1 0 104 0 -1 2524
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220663
transform 1 0 1280 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220663
transform 1 0 104 0 1 2428
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220663
transform 1 0 1280 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220663
transform 1 0 104 0 -1 2416
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220663
transform 1 0 1280 0 1 2320
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220663
transform 1 0 104 0 1 2320
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220663
transform 1 0 1280 0 -1 2308
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220663
transform 1 0 104 0 -1 2308
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220663
transform 1 0 1280 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220663
transform 1 0 104 0 1 2208
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220663
transform 1 0 1280 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220663
transform 1 0 104 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220663
transform 1 0 1280 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220663
transform 1 0 104 0 1 2100
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220663
transform 1 0 1280 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220663
transform 1 0 104 0 -1 2092
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220663
transform 1 0 1280 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220663
transform 1 0 104 0 1 1992
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220663
transform 1 0 1280 0 -1 1980
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220663
transform 1 0 104 0 -1 1980
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220663
transform 1 0 1280 0 1 1876
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220663
transform 1 0 104 0 1 1876
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220663
transform 1 0 1280 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220663
transform 1 0 104 0 -1 1868
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220663
transform 1 0 1280 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220663
transform 1 0 104 0 1 1764
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220663
transform 1 0 1280 0 -1 1752
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220663
transform 1 0 104 0 -1 1752
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220663
transform 1 0 1280 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220663
transform 1 0 104 0 1 1652
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220663
transform 1 0 1280 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220663
transform 1 0 104 0 -1 1644
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220663
transform 1 0 1280 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220663
transform 1 0 104 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220663
transform 1 0 1280 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220663
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220663
transform 1 0 1280 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220663
transform 1 0 104 0 1 1436
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220663
transform 1 0 1280 0 -1 1428
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220663
transform 1 0 104 0 -1 1428
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220663
transform 1 0 1280 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220663
transform 1 0 104 0 1 1332
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220663
transform 1 0 1280 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220663
transform 1 0 104 0 -1 1324
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220663
transform 1 0 1280 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220663
transform 1 0 104 0 1 1228
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220663
transform 1 0 1280 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220663
transform 1 0 104 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220663
transform 1 0 1280 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220663
transform 1 0 104 0 1 1120
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220663
transform 1 0 1280 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220663
transform 1 0 104 0 -1 1108
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220663
transform 1 0 1280 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220663
transform 1 0 104 0 1 1008
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220663
transform 1 0 1280 0 -1 996
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220663
transform 1 0 104 0 -1 996
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220663
transform 1 0 1280 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220663
transform 1 0 104 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220663
transform 1 0 1280 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220663
transform 1 0 104 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220663
transform 1 0 1280 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220663
transform 1 0 104 0 1 788
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220663
transform 1 0 1280 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220663
transform 1 0 104 0 -1 776
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220663
transform 1 0 1280 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220663
transform 1 0 104 0 1 676
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220663
transform 1 0 1280 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220663
transform 1 0 104 0 -1 668
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220663
transform 1 0 1280 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220663
transform 1 0 104 0 1 568
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220663
transform 1 0 1280 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220663
transform 1 0 104 0 -1 556
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220663
transform 1 0 1280 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220663
transform 1 0 104 0 1 456
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220663
transform 1 0 1280 0 -1 444
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220663
transform 1 0 104 0 -1 444
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220663
transform 1 0 1280 0 1 340
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220663
transform 1 0 104 0 1 340
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220663
transform 1 0 1280 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220663
transform 1 0 104 0 -1 324
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220663
transform 1 0 1280 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220663
transform 1 0 104 0 1 220
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220663
transform 1 0 1280 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220663
transform 1 0 104 0 -1 204
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220663
transform 1 0 1280 0 1 88
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220663
transform 1 0 104 0 1 88
box 7 3 12 24
use _0_0std_0_0cells_0_0OR2X1  tst_5999_6
timestamp 1731220663
transform 1 0 2376 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5998_6
timestamp 1731220663
transform 1 0 2432 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5997_6
timestamp 1731220663
transform 1 0 2432 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5996_6
timestamp 1731220663
transform 1 0 2432 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5995_6
timestamp 1731220663
transform 1 0 2416 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5994_6
timestamp 1731220663
transform 1 0 2368 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5993_6
timestamp 1731220663
transform 1 0 2280 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5992_6
timestamp 1731220663
transform 1 0 2320 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5991_6
timestamp 1731220663
transform 1 0 2264 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5990_6
timestamp 1731220663
transform 1 0 2200 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5989_6
timestamp 1731220663
transform 1 0 2136 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5988_6
timestamp 1731220663
transform 1 0 2072 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5987_6
timestamp 1731220663
transform 1 0 2016 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5986_6
timestamp 1731220663
transform 1 0 1960 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5985_6
timestamp 1731220663
transform 1 0 1904 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5984_6
timestamp 1731220663
transform 1 0 1848 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5983_6
timestamp 1731220663
transform 1 0 2192 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5982_6
timestamp 1731220663
transform 1 0 2104 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5981_6
timestamp 1731220663
transform 1 0 2008 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5980_6
timestamp 1731220663
transform 1 0 1912 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5979_6
timestamp 1731220663
transform 1 0 2312 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5978_6
timestamp 1731220663
transform 1 0 2192 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5977_6
timestamp 1731220663
transform 1 0 2080 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5976_6
timestamp 1731220663
transform 1 0 1976 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5975_6
timestamp 1731220663
transform 1 0 1880 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5974_6
timestamp 1731220663
transform 1 0 2280 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5973_6
timestamp 1731220663
transform 1 0 2144 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5972_6
timestamp 1731220663
transform 1 0 2016 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5971_6
timestamp 1731220663
transform 1 0 1904 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5970_6
timestamp 1731220663
transform 1 0 1800 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5969_6
timestamp 1731220663
transform 1 0 2280 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5968_6
timestamp 1731220663
transform 1 0 2136 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5967_6
timestamp 1731220663
transform 1 0 2000 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5966_6
timestamp 1731220663
transform 1 0 1880 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5965_6
timestamp 1731220663
transform 1 0 1784 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5964_6
timestamp 1731220663
transform 1 0 1768 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5963_6
timestamp 1731220663
transform 1 0 1672 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5962_6
timestamp 1731220663
transform 1 0 1880 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5961_6
timestamp 1731220663
transform 1 0 2304 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5960_6
timestamp 1731220663
transform 1 0 2152 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5959_6
timestamp 1731220663
transform 1 0 2008 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5958_6
timestamp 1731220663
transform 1 0 1904 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5957_6
timestamp 1731220663
transform 1 0 1792 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5956_6
timestamp 1731220663
transform 1 0 2032 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5955_6
timestamp 1731220663
transform 1 0 2312 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5954_6
timestamp 1731220663
transform 1 0 2168 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5953_6
timestamp 1731220663
transform 1 0 2056 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5952_6
timestamp 1731220663
transform 1 0 1968 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5951_6
timestamp 1731220663
transform 1 0 1880 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5950_6
timestamp 1731220663
transform 1 0 2240 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5949_6
timestamp 1731220663
transform 1 0 2144 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5948_6
timestamp 1731220663
transform 1 0 2064 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5947_6
timestamp 1731220663
transform 1 0 1960 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5946_6
timestamp 1731220663
transform 1 0 2256 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5945_6
timestamp 1731220663
transform 1 0 2160 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5944_6
timestamp 1731220663
transform 1 0 2080 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5943_6
timestamp 1731220663
transform 1 0 2000 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5942_6
timestamp 1731220663
transform 1 0 2160 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5941_6
timestamp 1731220663
transform 1 0 2208 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5940_6
timestamp 1731220663
transform 1 0 2232 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5939_6
timestamp 1731220663
transform 1 0 2304 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5938_6
timestamp 1731220663
transform 1 0 2376 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5937_6
timestamp 1731220663
transform 1 0 2352 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5936_6
timestamp 1731220663
transform 1 0 2336 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5935_6
timestamp 1731220663
transform 1 0 2432 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5934_6
timestamp 1731220663
transform 1 0 2432 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5933_6
timestamp 1731220663
transform 1 0 2432 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5932_6
timestamp 1731220663
transform 1 0 2432 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5931_6
timestamp 1731220663
transform 1 0 2432 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5930_6
timestamp 1731220663
transform 1 0 2432 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5929_6
timestamp 1731220663
transform 1 0 2432 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5928_6
timestamp 1731220663
transform 1 0 2432 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5927_6
timestamp 1731220663
transform 1 0 2432 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5926_6
timestamp 1731220663
transform 1 0 2432 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5925_6
timestamp 1731220663
transform 1 0 2328 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5924_6
timestamp 1731220663
transform 1 0 2416 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5923_6
timestamp 1731220663
transform 1 0 2360 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5922_6
timestamp 1731220663
transform 1 0 2344 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5921_6
timestamp 1731220663
transform 1 0 2368 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5920_6
timestamp 1731220663
transform 1 0 2288 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5919_6
timestamp 1731220663
transform 1 0 2128 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5918_6
timestamp 1731220663
transform 1 0 2040 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5917_6
timestamp 1731220663
transform 1 0 1944 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5916_6
timestamp 1731220663
transform 1 0 2240 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5915_6
timestamp 1731220663
transform 1 0 2136 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5914_6
timestamp 1731220663
transform 1 0 2032 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5913_6
timestamp 1731220663
transform 1 0 1920 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5912_6
timestamp 1731220663
transform 1 0 2264 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5911_6
timestamp 1731220663
transform 1 0 2176 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5910_6
timestamp 1731220663
transform 1 0 2088 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5909_6
timestamp 1731220663
transform 1 0 2000 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5908_6
timestamp 1731220663
transform 1 0 1912 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5907_6
timestamp 1731220663
transform 1 0 2312 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5906_6
timestamp 1731220663
transform 1 0 2192 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5905_6
timestamp 1731220663
transform 1 0 2072 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5904_6
timestamp 1731220663
transform 1 0 1968 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5903_6
timestamp 1731220663
transform 1 0 1880 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5902_6
timestamp 1731220663
transform 1 0 1808 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5901_6
timestamp 1731220663
transform 1 0 2272 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5900_6
timestamp 1731220663
transform 1 0 2128 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5899_6
timestamp 1731220663
transform 1 0 1992 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5898_6
timestamp 1731220663
transform 1 0 1872 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5897_6
timestamp 1731220663
transform 1 0 1768 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5896_6
timestamp 1731220663
transform 1 0 1728 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5895_6
timestamp 1731220663
transform 1 0 1800 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5894_6
timestamp 1731220663
transform 1 0 1880 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5893_6
timestamp 1731220663
transform 1 0 2208 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5892_6
timestamp 1731220663
transform 1 0 2088 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5891_6
timestamp 1731220663
transform 1 0 1976 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5890_6
timestamp 1731220663
transform 1 0 1984 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5889_6
timestamp 1731220663
transform 1 0 1896 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5888_6
timestamp 1731220663
transform 1 0 1816 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5887_6
timestamp 1731220663
transform 1 0 2328 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5886_6
timestamp 1731220663
transform 1 0 2208 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5885_6
timestamp 1731220663
transform 1 0 2088 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5884_6
timestamp 1731220663
transform 1 0 2064 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5883_6
timestamp 1731220663
transform 1 0 1976 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5882_6
timestamp 1731220663
transform 1 0 1888 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5881_6
timestamp 1731220663
transform 1 0 2352 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5880_6
timestamp 1731220663
transform 1 0 2248 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5879_6
timestamp 1731220663
transform 1 0 2152 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5878_6
timestamp 1731220663
transform 1 0 2064 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5877_6
timestamp 1731220663
transform 1 0 1960 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5876_6
timestamp 1731220663
transform 1 0 2168 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5875_6
timestamp 1731220663
transform 1 0 2264 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5874_6
timestamp 1731220663
transform 1 0 2360 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5873_6
timestamp 1731220663
transform 1 0 2288 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5872_6
timestamp 1731220663
transform 1 0 2208 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5871_6
timestamp 1731220663
transform 1 0 2120 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5870_6
timestamp 1731220663
transform 1 0 2024 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5869_6
timestamp 1731220663
transform 1 0 1920 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5868_6
timestamp 1731220663
transform 1 0 2232 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5867_6
timestamp 1731220663
transform 1 0 2160 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5866_6
timestamp 1731220663
transform 1 0 2080 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5865_6
timestamp 1731220663
transform 1 0 1992 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5864_6
timestamp 1731220663
transform 1 0 1896 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5863_6
timestamp 1731220663
transform 1 0 2192 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5862_6
timestamp 1731220663
transform 1 0 2072 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5861_6
timestamp 1731220663
transform 1 0 1960 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5860_6
timestamp 1731220663
transform 1 0 1848 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5859_6
timestamp 1731220663
transform 1 0 2088 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5858_6
timestamp 1731220663
transform 1 0 1968 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5857_6
timestamp 1731220663
transform 1 0 1856 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5856_6
timestamp 1731220663
transform 1 0 1752 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5855_6
timestamp 1731220663
transform 1 0 1808 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5854_6
timestamp 1731220663
transform 1 0 1920 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5853_6
timestamp 1731220663
transform 1 0 2040 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5852_6
timestamp 1731220663
transform 1 0 2168 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5851_6
timestamp 1731220663
transform 1 0 2032 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5850_6
timestamp 1731220663
transform 1 0 1936 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5849_6
timestamp 1731220663
transform 1 0 2272 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5848_6
timestamp 1731220663
transform 1 0 2224 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5847_6
timestamp 1731220663
transform 1 0 2128 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5846_6
timestamp 1731220663
transform 1 0 2320 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5845_6
timestamp 1731220663
transform 1 0 2296 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5844_6
timestamp 1731220663
transform 1 0 2208 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5843_6
timestamp 1731220663
transform 1 0 2328 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5842_6
timestamp 1731220663
transform 1 0 2320 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5841_6
timestamp 1731220663
transform 1 0 2304 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5840_6
timestamp 1731220663
transform 1 0 2368 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5839_6
timestamp 1731220663
transform 1 0 2432 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5838_6
timestamp 1731220663
transform 1 0 2432 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5837_6
timestamp 1731220663
transform 1 0 2432 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5836_6
timestamp 1731220663
transform 1 0 2432 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5835_6
timestamp 1731220663
transform 1 0 2432 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5834_6
timestamp 1731220663
transform 1 0 2432 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5833_6
timestamp 1731220663
transform 1 0 2376 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5832_6
timestamp 1731220663
transform 1 0 2432 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5831_6
timestamp 1731220663
transform 1 0 2432 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5830_6
timestamp 1731220663
transform 1 0 2432 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5829_6
timestamp 1731220663
transform 1 0 2416 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5828_6
timestamp 1731220663
transform 1 0 2432 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5827_6
timestamp 1731220663
transform 1 0 2432 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5826_6
timestamp 1731220663
transform 1 0 2432 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5825_6
timestamp 1731220663
transform 1 0 2432 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5824_6
timestamp 1731220663
transform 1 0 2432 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5823_6
timestamp 1731220663
transform 1 0 2432 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5822_6
timestamp 1731220663
transform 1 0 2432 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5821_6
timestamp 1731220663
transform 1 0 2432 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5820_6
timestamp 1731220663
transform 1 0 2432 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5819_6
timestamp 1731220663
transform 1 0 2432 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5818_6
timestamp 1731220663
transform 1 0 2320 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5817_6
timestamp 1731220663
transform 1 0 2432 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5816_6
timestamp 1731220663
transform 1 0 2376 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5815_6
timestamp 1731220663
transform 1 0 2320 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5814_6
timestamp 1731220663
transform 1 0 2264 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5813_6
timestamp 1731220663
transform 1 0 2200 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5812_6
timestamp 1731220663
transform 1 0 2136 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5811_6
timestamp 1731220663
transform 1 0 2072 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5810_6
timestamp 1731220663
transform 1 0 2016 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5809_6
timestamp 1731220663
transform 1 0 1960 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5808_6
timestamp 1731220663
transform 1 0 1904 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5807_6
timestamp 1731220663
transform 1 0 2304 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5806_6
timestamp 1731220663
transform 1 0 2208 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5805_6
timestamp 1731220663
transform 1 0 2112 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5804_6
timestamp 1731220663
transform 1 0 2024 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5803_6
timestamp 1731220663
transform 1 0 1928 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5802_6
timestamp 1731220663
transform 1 0 2184 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5801_6
timestamp 1731220663
transform 1 0 2088 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5800_6
timestamp 1731220663
transform 1 0 1992 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5799_6
timestamp 1731220663
transform 1 0 1904 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5798_6
timestamp 1731220663
transform 1 0 1808 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5797_6
timestamp 1731220663
transform 1 0 2088 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5796_6
timestamp 1731220663
transform 1 0 2000 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5795_6
timestamp 1731220663
transform 1 0 1912 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5794_6
timestamp 1731220663
transform 1 0 1824 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5793_6
timestamp 1731220663
transform 1 0 1744 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5792_6
timestamp 1731220663
transform 1 0 1712 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5791_6
timestamp 1731220663
transform 1 0 1800 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5790_6
timestamp 1731220663
transform 1 0 1888 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5789_6
timestamp 1731220663
transform 1 0 1984 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5788_6
timestamp 1731220663
transform 1 0 2080 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5787_6
timestamp 1731220663
transform 1 0 2120 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5786_6
timestamp 1731220663
transform 1 0 2032 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5785_6
timestamp 1731220663
transform 1 0 1944 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5784_6
timestamp 1731220663
transform 1 0 1856 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5783_6
timestamp 1731220663
transform 1 0 1768 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5782_6
timestamp 1731220663
transform 1 0 2160 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5781_6
timestamp 1731220663
transform 1 0 2104 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5780_6
timestamp 1731220663
transform 1 0 2048 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5779_6
timestamp 1731220663
transform 1 0 1992 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5778_6
timestamp 1731220663
transform 1 0 1936 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5777_6
timestamp 1731220663
transform 1 0 1880 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5776_6
timestamp 1731220663
transform 1 0 1824 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5775_6
timestamp 1731220663
transform 1 0 1768 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5774_6
timestamp 1731220663
transform 1 0 1712 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5773_6
timestamp 1731220663
transform 1 0 1656 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5772_6
timestamp 1731220663
transform 1 0 1600 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5771_6
timestamp 1731220663
transform 1 0 1544 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5770_6
timestamp 1731220663
transform 1 0 1488 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5769_6
timestamp 1731220663
transform 1 0 1432 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5768_6
timestamp 1731220663
transform 1 0 1376 0 1 2504
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5767_6
timestamp 1731220663
transform 1 0 1680 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5766_6
timestamp 1731220663
transform 1 0 1592 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5765_6
timestamp 1731220663
transform 1 0 1504 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5764_6
timestamp 1731220663
transform 1 0 1416 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5763_6
timestamp 1731220663
transform 1 0 1344 0 -1 2496
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5762_6
timestamp 1731220663
transform 1 0 1616 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5761_6
timestamp 1731220663
transform 1 0 1520 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5760_6
timestamp 1731220663
transform 1 0 1416 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5759_6
timestamp 1731220663
transform 1 0 1344 0 1 2384
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5758_6
timestamp 1731220663
transform 1 0 1344 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5757_6
timestamp 1731220663
transform 1 0 1400 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5756_6
timestamp 1731220663
transform 1 0 1488 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5755_6
timestamp 1731220663
transform 1 0 1664 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5754_6
timestamp 1731220663
transform 1 0 1576 0 -1 2376
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5753_6
timestamp 1731220663
transform 1 0 1520 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5752_6
timestamp 1731220663
transform 1 0 1432 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5751_6
timestamp 1731220663
transform 1 0 1344 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5750_6
timestamp 1731220663
transform 1 0 1616 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5749_6
timestamp 1731220663
transform 1 0 1712 0 1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5748_6
timestamp 1731220663
transform 1 0 1832 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5747_6
timestamp 1731220663
transform 1 0 1728 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5746_6
timestamp 1731220663
transform 1 0 1632 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5745_6
timestamp 1731220663
transform 1 0 1536 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5744_6
timestamp 1731220663
transform 1 0 1448 0 -1 2268
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5743_6
timestamp 1731220663
transform 1 0 1544 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5742_6
timestamp 1731220663
transform 1 0 1600 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5741_6
timestamp 1731220663
transform 1 0 1656 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5740_6
timestamp 1731220663
transform 1 0 1720 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5739_6
timestamp 1731220663
transform 1 0 1848 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5738_6
timestamp 1731220663
transform 1 0 1784 0 1 2160
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5737_6
timestamp 1731220663
transform 1 0 1784 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5736_6
timestamp 1731220663
transform 1 0 1712 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5735_6
timestamp 1731220663
transform 1 0 1656 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5734_6
timestamp 1731220663
transform 1 0 1864 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5733_6
timestamp 1731220663
transform 1 0 1960 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5732_6
timestamp 1731220663
transform 1 0 2072 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5731_6
timestamp 1731220663
transform 1 0 2192 0 -1 2148
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5730_6
timestamp 1731220663
transform 1 0 2296 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5729_6
timestamp 1731220663
transform 1 0 2144 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5728_6
timestamp 1731220663
transform 1 0 2000 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5727_6
timestamp 1731220663
transform 1 0 1872 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5726_6
timestamp 1731220663
transform 1 0 1760 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5725_6
timestamp 1731220663
transform 1 0 1816 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5724_6
timestamp 1731220663
transform 1 0 1928 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5723_6
timestamp 1731220663
transform 1 0 2048 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5722_6
timestamp 1731220663
transform 1 0 2312 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5721_6
timestamp 1731220663
transform 1 0 2176 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5720_6
timestamp 1731220663
transform 1 0 2128 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5719_6
timestamp 1731220663
transform 1 0 2024 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5718_6
timestamp 1731220663
transform 1 0 1920 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5717_6
timestamp 1731220663
transform 1 0 2344 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5716_6
timestamp 1731220663
transform 1 0 2232 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5715_6
timestamp 1731220663
transform 1 0 2192 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5714_6
timestamp 1731220663
transform 1 0 2104 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5713_6
timestamp 1731220663
transform 1 0 2008 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5712_6
timestamp 1731220663
transform 1 0 2280 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5711_6
timestamp 1731220663
transform 1 0 2368 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5710_6
timestamp 1731220663
transform 1 0 2432 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5709_6
timestamp 1731220663
transform 1 0 2344 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5708_6
timestamp 1731220663
transform 1 0 2248 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5707_6
timestamp 1731220663
transform 1 0 2152 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5706_6
timestamp 1731220663
transform 1 0 2056 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5705_6
timestamp 1731220663
transform 1 0 2360 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5704_6
timestamp 1731220663
transform 1 0 2264 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5703_6
timestamp 1731220663
transform 1 0 2176 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5702_6
timestamp 1731220663
transform 1 0 2080 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5701_6
timestamp 1731220663
transform 1 0 1976 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5700_6
timestamp 1731220663
transform 1 0 2328 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5699_6
timestamp 1731220663
transform 1 0 2208 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5698_6
timestamp 1731220663
transform 1 0 2088 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5697_6
timestamp 1731220663
transform 1 0 1976 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5696_6
timestamp 1731220663
transform 1 0 1864 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5695_6
timestamp 1731220663
transform 1 0 2304 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5694_6
timestamp 1731220663
transform 1 0 2152 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5693_6
timestamp 1731220663
transform 1 0 2008 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5692_6
timestamp 1731220663
transform 1 0 1872 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5691_6
timestamp 1731220663
transform 1 0 1752 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5690_6
timestamp 1731220663
transform 1 0 2304 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5689_6
timestamp 1731220663
transform 1 0 2160 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5688_6
timestamp 1731220663
transform 1 0 2032 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5687_6
timestamp 1731220663
transform 1 0 1912 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5686_6
timestamp 1731220663
transform 1 0 1816 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5685_6
timestamp 1731220663
transform 1 0 1728 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5684_6
timestamp 1731220663
transform 1 0 1656 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5683_6
timestamp 1731220663
transform 1 0 1576 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5682_6
timestamp 1731220663
transform 1 0 2096 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5681_6
timestamp 1731220663
transform 1 0 1928 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5680_6
timestamp 1731220663
transform 1 0 1776 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5679_6
timestamp 1731220663
transform 1 0 1640 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5678_6
timestamp 1731220663
transform 1 0 1520 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5677_6
timestamp 1731220663
transform 1 0 1832 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5676_6
timestamp 1731220663
transform 1 0 1728 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5675_6
timestamp 1731220663
transform 1 0 1624 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5674_6
timestamp 1731220663
transform 1 0 1608 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5673_6
timestamp 1731220663
transform 1 0 1512 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5672_6
timestamp 1731220663
transform 1 0 1704 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5671_6
timestamp 1731220663
transform 1 0 1656 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5670_6
timestamp 1731220663
transform 1 0 1568 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5669_6
timestamp 1731220663
transform 1 0 1480 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5668_6
timestamp 1731220663
transform 1 0 1560 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5667_6
timestamp 1731220663
transform 1 0 1648 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5666_6
timestamp 1731220663
transform 1 0 1744 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5665_6
timestamp 1731220663
transform 1 0 1696 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5664_6
timestamp 1731220663
transform 1 0 1592 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5663_6
timestamp 1731220663
transform 1 0 1800 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5662_6
timestamp 1731220663
transform 1 0 1808 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5661_6
timestamp 1731220663
transform 1 0 1688 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5660_6
timestamp 1731220663
transform 1 0 1568 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5659_6
timestamp 1731220663
transform 1 0 1712 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5658_6
timestamp 1731220663
transform 1 0 1840 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5657_6
timestamp 1731220663
transform 1 0 1800 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5656_6
timestamp 1731220663
transform 1 0 1712 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5655_6
timestamp 1731220663
transform 1 0 1624 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5654_6
timestamp 1731220663
transform 1 0 1744 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5653_6
timestamp 1731220663
transform 1 0 1680 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5652_6
timestamp 1731220663
transform 1 0 1672 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5651_6
timestamp 1731220663
transform 1 0 1592 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5650_6
timestamp 1731220663
transform 1 0 1672 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5649_6
timestamp 1731220663
transform 1 0 1680 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5648_6
timestamp 1731220663
transform 1 0 1744 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5647_6
timestamp 1731220663
transform 1 0 1824 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5646_6
timestamp 1731220663
transform 1 0 1736 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5645_6
timestamp 1731220663
transform 1 0 1648 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5644_6
timestamp 1731220663
transform 1 0 1680 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5643_6
timestamp 1731220663
transform 1 0 1800 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5642_6
timestamp 1731220663
transform 1 0 1840 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5641_6
timestamp 1731220663
transform 1 0 1728 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5640_6
timestamp 1731220663
transform 1 0 1728 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5639_6
timestamp 1731220663
transform 1 0 1824 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5638_6
timestamp 1731220663
transform 1 0 1912 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5637_6
timestamp 1731220663
transform 1 0 1856 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5636_6
timestamp 1731220663
transform 1 0 1752 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5635_6
timestamp 1731220663
transform 1 0 1792 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5634_6
timestamp 1731220663
transform 1 0 1704 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5633_6
timestamp 1731220663
transform 1 0 1608 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5632_6
timestamp 1731220663
transform 1 0 1688 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5631_6
timestamp 1731220663
transform 1 0 1592 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5630_6
timestamp 1731220663
transform 1 0 1504 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5629_6
timestamp 1731220663
transform 1 0 1592 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5628_6
timestamp 1731220663
transform 1 0 1712 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5627_6
timestamp 1731220663
transform 1 0 1656 0 1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5626_6
timestamp 1731220663
transform 1 0 1616 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5625_6
timestamp 1731220663
transform 1 0 1704 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5624_6
timestamp 1731220663
transform 1 0 1792 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5623_6
timestamp 1731220663
transform 1 0 1704 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5622_6
timestamp 1731220663
transform 1 0 1608 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5621_6
timestamp 1731220663
transform 1 0 1704 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5620_6
timestamp 1731220663
transform 1 0 1808 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5619_6
timestamp 1731220663
transform 1 0 1792 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5618_6
timestamp 1731220663
transform 1 0 1736 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5617_6
timestamp 1731220663
transform 1 0 1680 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5616_6
timestamp 1731220663
transform 1 0 1624 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5615_6
timestamp 1731220663
transform 1 0 1568 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5614_6
timestamp 1731220663
transform 1 0 1512 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5613_6
timestamp 1731220663
transform 1 0 1456 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5612_6
timestamp 1731220663
transform 1 0 1400 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5611_6
timestamp 1731220663
transform 1 0 1344 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5610_6
timestamp 1731220663
transform 1 0 1384 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5609_6
timestamp 1731220663
transform 1 0 1488 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5608_6
timestamp 1731220663
transform 1 0 1592 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5607_6
timestamp 1731220663
transform 1 0 1512 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5606_6
timestamp 1731220663
transform 1 0 1416 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5605_6
timestamp 1731220663
transform 1 0 1344 0 1 212
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5604_6
timestamp 1731220663
transform 1 0 1520 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5603_6
timestamp 1731220663
transform 1 0 1424 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5602_6
timestamp 1731220663
transform 1 0 1344 0 -1 320
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5601_6
timestamp 1731220663
transform 1 0 1216 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5600_6
timestamp 1731220663
transform 1 0 1160 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5599_6
timestamp 1731220663
transform 1 0 1216 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5598_6
timestamp 1731220663
transform 1 0 1344 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5597_6
timestamp 1731220663
transform 1 0 1416 0 -1 428
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5596_6
timestamp 1731220663
transform 1 0 1496 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5595_6
timestamp 1731220663
transform 1 0 1408 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5594_6
timestamp 1731220663
transform 1 0 1344 0 1 432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5593_6
timestamp 1731220663
transform 1 0 1360 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5592_6
timestamp 1731220663
transform 1 0 1520 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5591_6
timestamp 1731220663
transform 1 0 1440 0 -1 540
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5590_6
timestamp 1731220663
transform 1 0 1432 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5589_6
timestamp 1731220663
transform 1 0 1536 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5588_6
timestamp 1731220663
transform 1 0 1648 0 1 544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5587_6
timestamp 1731220663
transform 1 0 1640 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5586_6
timestamp 1731220663
transform 1 0 1552 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5585_6
timestamp 1731220663
transform 1 0 1472 0 -1 652
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5584_6
timestamp 1731220663
transform 1 0 1616 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5583_6
timestamp 1731220663
transform 1 0 1512 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5582_6
timestamp 1731220663
transform 1 0 1408 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5581_6
timestamp 1731220663
transform 1 0 1344 0 1 660
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5580_6
timestamp 1731220663
transform 1 0 1344 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5579_6
timestamp 1731220663
transform 1 0 1440 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5578_6
timestamp 1731220663
transform 1 0 1560 0 -1 768
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5577_6
timestamp 1731220663
transform 1 0 1568 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5576_6
timestamp 1731220663
transform 1 0 1488 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5575_6
timestamp 1731220663
transform 1 0 1416 0 1 772
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5574_6
timestamp 1731220663
transform 1 0 1480 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5573_6
timestamp 1731220663
transform 1 0 1616 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5572_6
timestamp 1731220663
transform 1 0 1552 0 -1 884
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5571_6
timestamp 1731220663
transform 1 0 1504 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5570_6
timestamp 1731220663
transform 1 0 1416 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5569_6
timestamp 1731220663
transform 1 0 1504 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5568_6
timestamp 1731220663
transform 1 0 1560 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5567_6
timestamp 1731220663
transform 1 0 1616 0 -1 1012
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5566_6
timestamp 1731220663
transform 1 0 1616 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5565_6
timestamp 1731220663
transform 1 0 1544 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5564_6
timestamp 1731220663
transform 1 0 1472 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5563_6
timestamp 1731220663
transform 1 0 1408 0 1 1020
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5562_6
timestamp 1731220663
transform 1 0 1360 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5561_6
timestamp 1731220663
transform 1 0 1440 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5560_6
timestamp 1731220663
transform 1 0 1528 0 -1 1132
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5559_6
timestamp 1731220663
transform 1 0 1576 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5558_6
timestamp 1731220663
transform 1 0 1448 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5557_6
timestamp 1731220663
transform 1 0 1344 0 1 1136
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5556_6
timestamp 1731220663
transform 1 0 1440 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5555_6
timestamp 1731220663
transform 1 0 1344 0 -1 1240
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5554_6
timestamp 1731220663
transform 1 0 1216 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5553_6
timestamp 1731220663
transform 1 0 1344 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5552_6
timestamp 1731220663
transform 1 0 1400 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5551_6
timestamp 1731220663
transform 1 0 1496 0 1 1256
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5550_6
timestamp 1731220663
transform 1 0 1472 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5549_6
timestamp 1731220663
transform 1 0 1400 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5548_6
timestamp 1731220663
transform 1 0 1344 0 -1 1368
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5547_6
timestamp 1731220663
transform 1 0 1344 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5546_6
timestamp 1731220663
transform 1 0 1400 0 1 1372
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5545_6
timestamp 1731220663
transform 1 0 1344 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5544_6
timestamp 1731220663
transform 1 0 1416 0 -1 1480
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5543_6
timestamp 1731220663
transform 1 0 1520 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5542_6
timestamp 1731220663
transform 1 0 1416 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5541_6
timestamp 1731220663
transform 1 0 1344 0 1 1484
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5540_6
timestamp 1731220663
transform 1 0 1344 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5539_6
timestamp 1731220663
transform 1 0 1416 0 -1 1588
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5538_6
timestamp 1731220663
transform 1 0 1496 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5537_6
timestamp 1731220663
transform 1 0 1408 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5536_6
timestamp 1731220663
transform 1 0 1344 0 1 1592
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5535_6
timestamp 1731220663
transform 1 0 1344 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5534_6
timestamp 1731220663
transform 1 0 1640 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5533_6
timestamp 1731220663
transform 1 0 1528 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5532_6
timestamp 1731220663
transform 1 0 1424 0 -1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5531_6
timestamp 1731220663
transform 1 0 1352 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5530_6
timestamp 1731220663
transform 1 0 1448 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5529_6
timestamp 1731220663
transform 1 0 1752 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5528_6
timestamp 1731220663
transform 1 0 1648 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5527_6
timestamp 1731220663
transform 1 0 1544 0 1 1704
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5526_6
timestamp 1731220663
transform 1 0 1456 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5525_6
timestamp 1731220663
transform 1 0 1552 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5524_6
timestamp 1731220663
transform 1 0 1872 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5523_6
timestamp 1731220663
transform 1 0 1760 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5522_6
timestamp 1731220663
transform 1 0 1656 0 -1 1812
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5521_6
timestamp 1731220663
transform 1 0 1664 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5520_6
timestamp 1731220663
transform 1 0 1584 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5519_6
timestamp 1731220663
transform 1 0 1512 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5518_6
timestamp 1731220663
transform 1 0 1760 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5517_6
timestamp 1731220663
transform 1 0 1856 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5516_6
timestamp 1731220663
transform 1 0 1960 0 1 1816
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5515_6
timestamp 1731220663
transform 1 0 1912 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5514_6
timestamp 1731220663
transform 1 0 1808 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5513_6
timestamp 1731220663
transform 1 0 1704 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5512_6
timestamp 1731220663
transform 1 0 1608 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5511_6
timestamp 1731220663
transform 1 0 1520 0 -1 1920
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5510_6
timestamp 1731220663
transform 1 0 1816 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5509_6
timestamp 1731220663
transform 1 0 1712 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5508_6
timestamp 1731220663
transform 1 0 1616 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5507_6
timestamp 1731220663
transform 1 0 1520 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5506_6
timestamp 1731220663
transform 1 0 1432 0 1 1924
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5505_6
timestamp 1731220663
transform 1 0 1712 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5504_6
timestamp 1731220663
transform 1 0 1608 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5503_6
timestamp 1731220663
transform 1 0 1512 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5502_6
timestamp 1731220663
transform 1 0 1416 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5501_6
timestamp 1731220663
transform 1 0 1344 0 -1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5500_6
timestamp 1731220663
transform 1 0 1656 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5499_6
timestamp 1731220663
transform 1 0 1568 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5498_6
timestamp 1731220663
transform 1 0 1480 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5497_6
timestamp 1731220663
transform 1 0 1400 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5496_6
timestamp 1731220663
transform 1 0 1344 0 1 2032
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5495_6
timestamp 1731220663
transform 1 0 1216 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5494_6
timestamp 1731220663
transform 1 0 1160 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5493_6
timestamp 1731220663
transform 1 0 1216 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5492_6
timestamp 1731220663
transform 1 0 1128 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5491_6
timestamp 1731220663
transform 1 0 1016 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5490_6
timestamp 1731220663
transform 1 0 904 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5489_6
timestamp 1731220663
transform 1 0 1096 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5488_6
timestamp 1731220663
transform 1 0 1024 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5487_6
timestamp 1731220663
transform 1 0 960 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5486_6
timestamp 1731220663
transform 1 0 896 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5485_6
timestamp 1731220663
transform 1 0 824 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5484_6
timestamp 1731220663
transform 1 0 752 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5483_6
timestamp 1731220663
transform 1 0 1040 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5482_6
timestamp 1731220663
transform 1 0 952 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5481_6
timestamp 1731220663
transform 1 0 864 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5480_6
timestamp 1731220663
transform 1 0 776 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5479_6
timestamp 1731220663
transform 1 0 696 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5478_6
timestamp 1731220663
transform 1 0 688 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5477_6
timestamp 1731220663
transform 1 0 792 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5476_6
timestamp 1731220663
transform 1 0 1008 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5475_6
timestamp 1731220663
transform 1 0 896 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5474_6
timestamp 1731220663
transform 1 0 840 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5473_6
timestamp 1731220663
transform 1 0 1016 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5472_6
timestamp 1731220663
transform 1 0 1032 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5471_6
timestamp 1731220663
transform 1 0 1016 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5470_6
timestamp 1731220663
transform 1 0 1096 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5469_6
timestamp 1731220663
transform 1 0 1096 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5468_6
timestamp 1731220663
transform 1 0 1152 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5467_6
timestamp 1731220663
transform 1 0 1040 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5466_6
timestamp 1731220663
transform 1 0 1048 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5465_6
timestamp 1731220663
transform 1 0 1168 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5464_6
timestamp 1731220663
transform 1 0 1168 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5463_6
timestamp 1731220663
transform 1 0 1040 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5462_6
timestamp 1731220663
transform 1 0 944 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5461_6
timestamp 1731220663
transform 1 0 1056 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5460_6
timestamp 1731220663
transform 1 0 1168 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5459_6
timestamp 1731220663
transform 1 0 1144 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5458_6
timestamp 1731220663
transform 1 0 1040 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5457_6
timestamp 1731220663
transform 1 0 936 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5456_6
timestamp 1731220663
transform 1 0 832 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5455_6
timestamp 1731220663
transform 1 0 1080 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5454_6
timestamp 1731220663
transform 1 0 984 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5453_6
timestamp 1731220663
transform 1 0 888 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5452_6
timestamp 1731220663
transform 1 0 800 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5451_6
timestamp 1731220663
transform 1 0 704 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5450_6
timestamp 1731220663
transform 1 0 976 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5449_6
timestamp 1731220663
transform 1 0 872 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5448_6
timestamp 1731220663
transform 1 0 776 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5447_6
timestamp 1731220663
transform 1 0 680 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5446_6
timestamp 1731220663
transform 1 0 584 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5445_6
timestamp 1731220663
transform 1 0 872 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5444_6
timestamp 1731220663
transform 1 0 776 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5443_6
timestamp 1731220663
transform 1 0 680 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5442_6
timestamp 1731220663
transform 1 0 592 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5441_6
timestamp 1731220663
transform 1 0 504 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5440_6
timestamp 1731220663
transform 1 0 1072 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5439_6
timestamp 1731220663
transform 1 0 904 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5438_6
timestamp 1731220663
transform 1 0 752 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5437_6
timestamp 1731220663
transform 1 0 616 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5436_6
timestamp 1731220663
transform 1 0 624 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5435_6
timestamp 1731220663
transform 1 0 680 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5434_6
timestamp 1731220663
transform 1 0 736 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5433_6
timestamp 1731220663
transform 1 0 792 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5432_6
timestamp 1731220663
transform 1 0 848 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5431_6
timestamp 1731220663
transform 1 0 904 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5430_6
timestamp 1731220663
transform 1 0 848 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5429_6
timestamp 1731220663
transform 1 0 792 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5428_6
timestamp 1731220663
transform 1 0 736 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5427_6
timestamp 1731220663
transform 1 0 960 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5426_6
timestamp 1731220663
transform 1 0 904 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5425_6
timestamp 1731220663
transform 1 0 840 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5424_6
timestamp 1731220663
transform 1 0 760 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5423_6
timestamp 1731220663
transform 1 0 672 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5422_6
timestamp 1731220663
transform 1 0 920 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5421_6
timestamp 1731220663
transform 1 0 1096 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5420_6
timestamp 1731220663
transform 1 0 1008 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5419_6
timestamp 1731220663
transform 1 0 960 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5418_6
timestamp 1731220663
transform 1 0 856 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5417_6
timestamp 1731220663
transform 1 0 744 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5416_6
timestamp 1731220663
transform 1 0 1184 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5415_6
timestamp 1731220663
transform 1 0 1072 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5414_6
timestamp 1731220663
transform 1 0 752 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5413_6
timestamp 1731220663
transform 1 0 656 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5412_6
timestamp 1731220663
transform 1 0 928 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5411_6
timestamp 1731220663
transform 1 0 1008 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5410_6
timestamp 1731220663
transform 1 0 1080 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5409_6
timestamp 1731220663
transform 1 0 1216 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5408_6
timestamp 1731220663
transform 1 0 1160 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5407_6
timestamp 1731220663
transform 1 0 1152 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5406_6
timestamp 1731220663
transform 1 0 1344 0 1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5405_6
timestamp 1731220663
transform 1 0 1216 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5404_6
timestamp 1731220663
transform 1 0 1216 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5403_6
timestamp 1731220663
transform 1 0 1160 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5402_6
timestamp 1731220663
transform 1 0 1080 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5401_6
timestamp 1731220663
transform 1 0 1000 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5400_6
timestamp 1731220663
transform 1 0 920 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5399_6
timestamp 1731220663
transform 1 0 832 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5398_6
timestamp 1731220663
transform 1 0 1072 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5397_6
timestamp 1731220663
transform 1 0 992 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5396_6
timestamp 1731220663
transform 1 0 904 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5395_6
timestamp 1731220663
transform 1 0 840 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5394_6
timestamp 1731220663
transform 1 0 808 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5393_6
timestamp 1731220663
transform 1 0 712 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5392_6
timestamp 1731220663
transform 1 0 736 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5391_6
timestamp 1731220663
transform 1 0 1048 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5390_6
timestamp 1731220663
transform 1 0 960 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5389_6
timestamp 1731220663
transform 1 0 872 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5388_6
timestamp 1731220663
transform 1 0 784 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5387_6
timestamp 1731220663
transform 1 0 704 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5386_6
timestamp 1731220663
transform 1 0 968 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5385_6
timestamp 1731220663
transform 1 0 888 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5384_6
timestamp 1731220663
transform 1 0 816 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5383_6
timestamp 1731220663
transform 1 0 744 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5382_6
timestamp 1731220663
transform 1 0 672 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5381_6
timestamp 1731220663
transform 1 0 600 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5380_6
timestamp 1731220663
transform 1 0 888 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5379_6
timestamp 1731220663
transform 1 0 816 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5378_6
timestamp 1731220663
transform 1 0 744 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5377_6
timestamp 1731220663
transform 1 0 680 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5376_6
timestamp 1731220663
transform 1 0 616 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5375_6
timestamp 1731220663
transform 1 0 584 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5374_6
timestamp 1731220663
transform 1 0 648 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5373_6
timestamp 1731220663
transform 1 0 712 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5372_6
timestamp 1731220663
transform 1 0 776 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5371_6
timestamp 1731220663
transform 1 0 912 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5370_6
timestamp 1731220663
transform 1 0 840 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5369_6
timestamp 1731220663
transform 1 0 824 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5368_6
timestamp 1731220663
transform 1 0 744 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5367_6
timestamp 1731220663
transform 1 0 664 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5366_6
timestamp 1731220663
transform 1 0 904 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5365_6
timestamp 1731220663
transform 1 0 1064 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5364_6
timestamp 1731220663
transform 1 0 984 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5363_6
timestamp 1731220663
transform 1 0 960 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5362_6
timestamp 1731220663
transform 1 0 872 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5361_6
timestamp 1731220663
transform 1 0 784 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5360_6
timestamp 1731220663
transform 1 0 1144 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5359_6
timestamp 1731220663
transform 1 0 1048 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5358_6
timestamp 1731220663
transform 1 0 1032 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5357_6
timestamp 1731220663
transform 1 0 928 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5356_6
timestamp 1731220663
transform 1 0 824 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5355_6
timestamp 1731220663
transform 1 0 1136 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5354_6
timestamp 1731220663
transform 1 0 1216 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5353_6
timestamp 1731220663
transform 1 0 1216 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5352_6
timestamp 1731220663
transform 1 0 1120 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5351_6
timestamp 1731220663
transform 1 0 1000 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5350_6
timestamp 1731220663
transform 1 0 944 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5349_6
timestamp 1731220663
transform 1 0 1016 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5348_6
timestamp 1731220663
transform 1 0 1088 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5347_6
timestamp 1731220663
transform 1 0 1024 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5346_6
timestamp 1731220663
transform 1 0 1128 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5345_6
timestamp 1731220663
transform 1 0 1192 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5344_6
timestamp 1731220663
transform 1 0 1088 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5343_6
timestamp 1731220663
transform 1 0 984 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5342_6
timestamp 1731220663
transform 1 0 952 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5341_6
timestamp 1731220663
transform 1 0 1040 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5340_6
timestamp 1731220663
transform 1 0 1128 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5339_6
timestamp 1731220663
transform 1 0 1176 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5338_6
timestamp 1731220663
transform 1 0 1112 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5337_6
timestamp 1731220663
transform 1 0 1048 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5336_6
timestamp 1731220663
transform 1 0 984 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5335_6
timestamp 1731220663
transform 1 0 920 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5334_6
timestamp 1731220663
transform 1 0 856 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5333_6
timestamp 1731220663
transform 1 0 792 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5332_6
timestamp 1731220663
transform 1 0 728 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5331_6
timestamp 1731220663
transform 1 0 664 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5330_6
timestamp 1731220663
transform 1 0 688 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5329_6
timestamp 1731220663
transform 1 0 776 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5328_6
timestamp 1731220663
transform 1 0 864 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5327_6
timestamp 1731220663
transform 1 0 784 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5326_6
timestamp 1731220663
transform 1 0 688 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5325_6
timestamp 1731220663
transform 1 0 880 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5324_6
timestamp 1731220663
transform 1 0 920 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5323_6
timestamp 1731220663
transform 1 0 816 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5322_6
timestamp 1731220663
transform 1 0 720 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5321_6
timestamp 1731220663
transform 1 0 624 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5320_6
timestamp 1731220663
transform 1 0 568 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5319_6
timestamp 1731220663
transform 1 0 648 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5318_6
timestamp 1731220663
transform 1 0 728 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5317_6
timestamp 1731220663
transform 1 0 800 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5316_6
timestamp 1731220663
transform 1 0 872 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5315_6
timestamp 1731220663
transform 1 0 888 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5314_6
timestamp 1731220663
transform 1 0 776 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5313_6
timestamp 1731220663
transform 1 0 664 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5312_6
timestamp 1731220663
transform 1 0 560 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5311_6
timestamp 1731220663
transform 1 0 592 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5310_6
timestamp 1731220663
transform 1 0 712 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5309_6
timestamp 1731220663
transform 1 0 688 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5308_6
timestamp 1731220663
transform 1 0 584 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5307_6
timestamp 1731220663
transform 1 0 480 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5306_6
timestamp 1731220663
transform 1 0 576 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5305_6
timestamp 1731220663
transform 1 0 480 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5304_6
timestamp 1731220663
transform 1 0 448 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5303_6
timestamp 1731220663
transform 1 0 520 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5302_6
timestamp 1731220663
transform 1 0 480 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5301_6
timestamp 1731220663
transform 1 0 400 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5300_6
timestamp 1731220663
transform 1 0 552 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5299_6
timestamp 1731220663
transform 1 0 520 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5298_6
timestamp 1731220663
transform 1 0 432 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5297_6
timestamp 1731220663
transform 1 0 320 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5296_6
timestamp 1731220663
transform 1 0 240 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5295_6
timestamp 1731220663
transform 1 0 288 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5294_6
timestamp 1731220663
transform 1 0 368 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5293_6
timestamp 1731220663
transform 1 0 384 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5292_6
timestamp 1731220663
transform 1 0 368 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5291_6
timestamp 1731220663
transform 1 0 264 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5290_6
timestamp 1731220663
transform 1 0 464 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5289_6
timestamp 1731220663
transform 1 0 344 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5288_6
timestamp 1731220663
transform 1 0 296 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5287_6
timestamp 1731220663
transform 1 0 240 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5286_6
timestamp 1731220663
transform 1 0 376 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5285_6
timestamp 1731220663
transform 1 0 464 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5284_6
timestamp 1731220663
transform 1 0 488 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5283_6
timestamp 1731220663
transform 1 0 408 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5282_6
timestamp 1731220663
transform 1 0 336 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5281_6
timestamp 1731220663
transform 1 0 448 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5280_6
timestamp 1731220663
transform 1 0 368 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5279_6
timestamp 1731220663
transform 1 0 536 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5278_6
timestamp 1731220663
transform 1 0 496 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5277_6
timestamp 1731220663
transform 1 0 400 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5276_6
timestamp 1731220663
transform 1 0 592 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5275_6
timestamp 1731220663
transform 1 0 600 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5274_6
timestamp 1731220663
transform 1 0 504 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5273_6
timestamp 1731220663
transform 1 0 408 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5272_6
timestamp 1731220663
transform 1 0 600 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5271_6
timestamp 1731220663
transform 1 0 528 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5270_6
timestamp 1731220663
transform 1 0 464 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5269_6
timestamp 1731220663
transform 1 0 408 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5268_6
timestamp 1731220663
transform 1 0 352 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5267_6
timestamp 1731220663
transform 1 0 296 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5266_6
timestamp 1731220663
transform 1 0 240 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5265_6
timestamp 1731220663
transform 1 0 184 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5264_6
timestamp 1731220663
transform 1 0 128 0 1 84
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5263_6
timestamp 1731220663
transform 1 0 152 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5262_6
timestamp 1731220663
transform 1 0 320 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5261_6
timestamp 1731220663
transform 1 0 232 0 -1 208
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5260_6
timestamp 1731220663
transform 1 0 208 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5259_6
timestamp 1731220663
transform 1 0 128 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5258_6
timestamp 1731220663
transform 1 0 304 0 1 216
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5257_6
timestamp 1731220663
transform 1 0 280 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5256_6
timestamp 1731220663
transform 1 0 192 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5255_6
timestamp 1731220663
transform 1 0 128 0 -1 328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5254_6
timestamp 1731220663
transform 1 0 128 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5253_6
timestamp 1731220663
transform 1 0 256 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5252_6
timestamp 1731220663
transform 1 0 184 0 1 336
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5251_6
timestamp 1731220663
transform 1 0 184 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5250_6
timestamp 1731220663
transform 1 0 128 0 -1 448
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5249_6
timestamp 1731220663
transform 1 0 128 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5248_6
timestamp 1731220663
transform 1 0 224 0 1 452
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5247_6
timestamp 1731220663
transform 1 0 168 0 -1 560
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5246_6
timestamp 1731220663
transform 1 0 184 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5245_6
timestamp 1731220663
transform 1 0 280 0 1 564
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5244_6
timestamp 1731220663
transform 1 0 208 0 -1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5243_6
timestamp 1731220663
transform 1 0 152 0 1 672
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5242_6
timestamp 1731220663
transform 1 0 144 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5241_6
timestamp 1731220663
transform 1 0 240 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5240_6
timestamp 1731220663
transform 1 0 336 0 -1 780
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5239_6
timestamp 1731220663
transform 1 0 280 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5238_6
timestamp 1731220663
transform 1 0 216 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5237_6
timestamp 1731220663
transform 1 0 360 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5236_6
timestamp 1731220663
transform 1 0 440 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5235_6
timestamp 1731220663
transform 1 0 528 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5234_6
timestamp 1731220663
transform 1 0 616 0 1 784
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5233_6
timestamp 1731220663
transform 1 0 640 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5232_6
timestamp 1731220663
transform 1 0 536 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5231_6
timestamp 1731220663
transform 1 0 432 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5230_6
timestamp 1731220663
transform 1 0 336 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5229_6
timestamp 1731220663
transform 1 0 240 0 -1 892
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5228_6
timestamp 1731220663
transform 1 0 600 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5227_6
timestamp 1731220663
transform 1 0 488 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5226_6
timestamp 1731220663
transform 1 0 376 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5225_6
timestamp 1731220663
transform 1 0 272 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5224_6
timestamp 1731220663
transform 1 0 184 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5223_6
timestamp 1731220663
transform 1 0 128 0 1 896
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5222_6
timestamp 1731220663
transform 1 0 128 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5221_6
timestamp 1731220663
transform 1 0 208 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5220_6
timestamp 1731220663
transform 1 0 544 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5219_6
timestamp 1731220663
transform 1 0 432 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5218_6
timestamp 1731220663
transform 1 0 320 0 -1 1000
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5217_6
timestamp 1731220663
transform 1 0 280 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5216_6
timestamp 1731220663
transform 1 0 184 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5215_6
timestamp 1731220663
transform 1 0 128 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5214_6
timestamp 1731220663
transform 1 0 632 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5213_6
timestamp 1731220663
transform 1 0 512 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5212_6
timestamp 1731220663
transform 1 0 392 0 1 1004
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5211_6
timestamp 1731220663
transform 1 0 392 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5210_6
timestamp 1731220663
transform 1 0 304 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5209_6
timestamp 1731220663
transform 1 0 216 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5208_6
timestamp 1731220663
transform 1 0 488 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5207_6
timestamp 1731220663
transform 1 0 584 0 -1 1112
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5206_6
timestamp 1731220663
transform 1 0 512 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5205_6
timestamp 1731220663
transform 1 0 456 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5204_6
timestamp 1731220663
transform 1 0 400 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5203_6
timestamp 1731220663
transform 1 0 568 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5202_6
timestamp 1731220663
transform 1 0 680 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5201_6
timestamp 1731220663
transform 1 0 624 0 1 1116
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5200_6
timestamp 1731220663
transform 1 0 568 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5199_6
timestamp 1731220663
transform 1 0 512 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5198_6
timestamp 1731220663
transform 1 0 456 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5197_6
timestamp 1731220663
transform 1 0 400 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5196_6
timestamp 1731220663
transform 1 0 344 0 -1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5195_6
timestamp 1731220663
transform 1 0 504 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5194_6
timestamp 1731220663
transform 1 0 416 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5193_6
timestamp 1731220663
transform 1 0 344 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5192_6
timestamp 1731220663
transform 1 0 280 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5191_6
timestamp 1731220663
transform 1 0 224 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5190_6
timestamp 1731220663
transform 1 0 168 0 1 1224
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5189_6
timestamp 1731220663
transform 1 0 408 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5188_6
timestamp 1731220663
transform 1 0 312 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5187_6
timestamp 1731220663
transform 1 0 208 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5186_6
timestamp 1731220663
transform 1 0 128 0 -1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5185_6
timestamp 1731220663
transform 1 0 128 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5184_6
timestamp 1731220663
transform 1 0 192 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5183_6
timestamp 1731220663
transform 1 0 288 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5182_6
timestamp 1731220663
transform 1 0 384 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5181_6
timestamp 1731220663
transform 1 0 488 0 1 1328
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5180_6
timestamp 1731220663
transform 1 0 408 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5179_6
timestamp 1731220663
transform 1 0 312 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5178_6
timestamp 1731220663
transform 1 0 224 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5177_6
timestamp 1731220663
transform 1 0 504 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5176_6
timestamp 1731220663
transform 1 0 608 0 -1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5175_6
timestamp 1731220663
transform 1 0 536 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5174_6
timestamp 1731220663
transform 1 0 440 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5173_6
timestamp 1731220663
transform 1 0 352 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5172_6
timestamp 1731220663
transform 1 0 728 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5171_6
timestamp 1731220663
transform 1 0 632 0 1 1432
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5170_6
timestamp 1731220663
transform 1 0 632 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5169_6
timestamp 1731220663
transform 1 0 544 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5168_6
timestamp 1731220663
transform 1 0 464 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5167_6
timestamp 1731220663
transform 1 0 832 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5166_6
timestamp 1731220663
transform 1 0 728 0 -1 1536
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5165_6
timestamp 1731220663
transform 1 0 680 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5164_6
timestamp 1731220663
transform 1 0 576 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5163_6
timestamp 1731220663
transform 1 0 912 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5162_6
timestamp 1731220663
transform 1 0 792 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5161_6
timestamp 1731220663
transform 1 0 736 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5160_6
timestamp 1731220663
transform 1 0 640 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5159_6
timestamp 1731220663
transform 1 0 832 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5158_6
timestamp 1731220663
transform 1 0 936 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5157_6
timestamp 1731220663
transform 1 0 928 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5156_6
timestamp 1731220663
transform 1 0 824 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5155_6
timestamp 1731220663
transform 1 0 720 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5154_6
timestamp 1731220663
transform 1 0 672 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5153_6
timestamp 1731220663
transform 1 0 776 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5152_6
timestamp 1731220663
transform 1 0 880 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5151_6
timestamp 1731220663
transform 1 0 984 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5150_6
timestamp 1731220663
transform 1 0 936 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5149_6
timestamp 1731220663
transform 1 0 856 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5148_6
timestamp 1731220663
transform 1 0 776 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5147_6
timestamp 1731220663
transform 1 0 696 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5146_6
timestamp 1731220663
transform 1 0 952 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5145_6
timestamp 1731220663
transform 1 0 880 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5144_6
timestamp 1731220663
transform 1 0 808 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5143_6
timestamp 1731220663
transform 1 0 736 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5142_6
timestamp 1731220663
transform 1 0 672 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5141_6
timestamp 1731220663
transform 1 0 608 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5140_6
timestamp 1731220663
transform 1 0 544 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5139_6
timestamp 1731220663
transform 1 0 472 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5138_6
timestamp 1731220663
transform 1 0 400 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5137_6
timestamp 1731220663
transform 1 0 416 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5136_6
timestamp 1731220663
transform 1 0 608 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5135_6
timestamp 1731220663
transform 1 0 512 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5134_6
timestamp 1731220663
transform 1 0 456 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5133_6
timestamp 1731220663
transform 1 0 568 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5132_6
timestamp 1731220663
transform 1 0 616 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5131_6
timestamp 1731220663
transform 1 0 512 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5130_6
timestamp 1731220663
transform 1 0 416 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5129_6
timestamp 1731220663
transform 1 0 400 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5128_6
timestamp 1731220663
transform 1 0 472 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5127_6
timestamp 1731220663
transform 1 0 552 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5126_6
timestamp 1731220663
transform 1 0 480 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5125_6
timestamp 1731220663
transform 1 0 400 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5124_6
timestamp 1731220663
transform 1 0 328 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5123_6
timestamp 1731220663
transform 1 0 264 0 1 1544
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5122_6
timestamp 1731220663
transform 1 0 264 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5121_6
timestamp 1731220663
transform 1 0 208 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5120_6
timestamp 1731220663
transform 1 0 328 0 -1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5119_6
timestamp 1731220663
transform 1 0 328 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5118_6
timestamp 1731220663
transform 1 0 248 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5117_6
timestamp 1731220663
transform 1 0 168 0 1 1648
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5116_6
timestamp 1731220663
transform 1 0 128 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5115_6
timestamp 1731220663
transform 1 0 232 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5114_6
timestamp 1731220663
transform 1 0 344 0 -1 1756
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5113_6
timestamp 1731220663
transform 1 0 312 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5112_6
timestamp 1731220663
transform 1 0 208 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5111_6
timestamp 1731220663
transform 1 0 128 0 1 1760
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5110_6
timestamp 1731220663
transform 1 0 128 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5109_6
timestamp 1731220663
transform 1 0 328 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5108_6
timestamp 1731220663
transform 1 0 256 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5107_6
timestamp 1731220663
transform 1 0 184 0 -1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5106_6
timestamp 1731220663
transform 1 0 128 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5105_6
timestamp 1731220663
transform 1 0 216 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5104_6
timestamp 1731220663
transform 1 0 664 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5103_6
timestamp 1731220663
transform 1 0 504 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5102_6
timestamp 1731220663
transform 1 0 352 0 1 1872
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5101_6
timestamp 1731220663
transform 1 0 280 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_5100_6
timestamp 1731220663
transform 1 0 200 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_599_6
timestamp 1731220663
transform 1 0 128 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_598_6
timestamp 1731220663
transform 1 0 584 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_597_6
timestamp 1731220663
transform 1 0 480 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_596_6
timestamp 1731220663
transform 1 0 376 0 -1 1984
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_595_6
timestamp 1731220663
transform 1 0 352 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_594_6
timestamp 1731220663
transform 1 0 272 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_593_6
timestamp 1731220663
transform 1 0 616 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_592_6
timestamp 1731220663
transform 1 0 528 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_591_6
timestamp 1731220663
transform 1 0 440 0 1 1988
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_590_6
timestamp 1731220663
transform 1 0 368 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_589_6
timestamp 1731220663
transform 1 0 440 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_588_6
timestamp 1731220663
transform 1 0 512 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_587_6
timestamp 1731220663
transform 1 0 592 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_586_6
timestamp 1731220663
transform 1 0 672 0 -1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_585_6
timestamp 1731220663
transform 1 0 792 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_584_6
timestamp 1731220663
transform 1 0 688 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_583_6
timestamp 1731220663
transform 1 0 584 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_582_6
timestamp 1731220663
transform 1 0 488 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_581_6
timestamp 1731220663
transform 1 0 392 0 1 2096
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_580_6
timestamp 1731220663
transform 1 0 552 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_579_6
timestamp 1731220663
transform 1 0 496 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_578_6
timestamp 1731220663
transform 1 0 440 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_577_6
timestamp 1731220663
transform 1 0 384 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_576_6
timestamp 1731220663
transform 1 0 328 0 -1 2200
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_575_6
timestamp 1731220663
transform 1 0 480 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_574_6
timestamp 1731220663
transform 1 0 424 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_573_6
timestamp 1731220663
transform 1 0 360 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_572_6
timestamp 1731220663
transform 1 0 296 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_571_6
timestamp 1731220663
transform 1 0 240 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_570_6
timestamp 1731220663
transform 1 0 464 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_569_6
timestamp 1731220663
transform 1 0 368 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_568_6
timestamp 1731220663
transform 1 0 280 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_567_6
timestamp 1731220663
transform 1 0 200 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_566_6
timestamp 1731220663
transform 1 0 480 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_565_6
timestamp 1731220663
transform 1 0 368 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_564_6
timestamp 1731220663
transform 1 0 256 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_563_6
timestamp 1731220663
transform 1 0 152 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_562_6
timestamp 1731220663
transform 1 0 408 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_561_6
timestamp 1731220663
transform 1 0 312 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_560_6
timestamp 1731220663
transform 1 0 224 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_559_6
timestamp 1731220663
transform 1 0 144 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_558_6
timestamp 1731220663
transform 1 0 160 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_557_6
timestamp 1731220663
transform 1 0 392 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_556_6
timestamp 1731220663
transform 1 0 304 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_555_6
timestamp 1731220663
transform 1 0 224 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_554_6
timestamp 1731220663
transform 1 0 216 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_553_6
timestamp 1731220663
transform 1 0 160 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_552_6
timestamp 1731220663
transform 1 0 272 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_551_6
timestamp 1731220663
transform 1 0 336 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_550_6
timestamp 1731220663
transform 1 0 400 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_549_6
timestamp 1731220663
transform 1 0 472 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_548_6
timestamp 1731220663
transform 1 0 552 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_547_6
timestamp 1731220663
transform 1 0 632 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_546_6
timestamp 1731220663
transform 1 0 576 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_545_6
timestamp 1731220663
transform 1 0 480 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_544_6
timestamp 1731220663
transform 1 0 672 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_543_6
timestamp 1731220663
transform 1 0 720 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_542_6
timestamp 1731220663
transform 1 0 616 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_541_6
timestamp 1731220663
transform 1 0 512 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_540_6
timestamp 1731220663
transform 1 0 600 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_539_6
timestamp 1731220663
transform 1 0 720 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_538_6
timestamp 1731220663
transform 1 0 728 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_537_6
timestamp 1731220663
transform 1 0 640 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_536_6
timestamp 1731220663
transform 1 0 552 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_535_6
timestamp 1731220663
transform 1 0 536 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_534_6
timestamp 1731220663
transform 1 0 592 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_533_6
timestamp 1731220663
transform 1 0 648 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_532_6
timestamp 1731220663
transform 1 0 704 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_531_6
timestamp 1731220663
transform 1 0 768 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_530_6
timestamp 1731220663
transform 1 0 832 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_529_6
timestamp 1731220663
transform 1 0 896 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_528_6
timestamp 1731220663
transform 1 0 1088 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_527_6
timestamp 1731220663
transform 1 0 1024 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_526_6
timestamp 1731220663
transform 1 0 960 0 1 2204
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_525_6
timestamp 1731220663
transform 1 0 896 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_524_6
timestamp 1731220663
transform 1 0 808 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_523_6
timestamp 1731220663
transform 1 0 1072 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_522_6
timestamp 1731220663
transform 1 0 984 0 -1 2312
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_521_6
timestamp 1731220663
transform 1 0 976 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_520_6
timestamp 1731220663
transform 1 0 848 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_519_6
timestamp 1731220663
transform 1 0 1104 0 1 2316
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_518_6
timestamp 1731220663
transform 1 0 1144 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_517_6
timestamp 1731220663
transform 1 0 1032 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_516_6
timestamp 1731220663
transform 1 0 928 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_515_6
timestamp 1731220663
transform 1 0 824 0 -1 2420
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_514_6
timestamp 1731220663
transform 1 0 1136 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_513_6
timestamp 1731220663
transform 1 0 1040 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_512_6
timestamp 1731220663
transform 1 0 944 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_511_6
timestamp 1731220663
transform 1 0 856 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_510_6
timestamp 1731220663
transform 1 0 768 0 1 2424
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_59_6
timestamp 1731220663
transform 1 0 1032 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_58_6
timestamp 1731220663
transform 1 0 952 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_57_6
timestamp 1731220663
transform 1 0 872 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_56_6
timestamp 1731220663
transform 1 0 792 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_55_6
timestamp 1731220663
transform 1 0 712 0 -1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_54_6
timestamp 1731220663
transform 1 0 920 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_53_6
timestamp 1731220663
transform 1 0 864 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_52_6
timestamp 1731220663
transform 1 0 808 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_51_6
timestamp 1731220663
transform 1 0 752 0 1 2528
box 4 4 48 48
use _0_0std_0_0cells_0_0OR2X1  tst_50_6
timestamp 1731220663
transform 1 0 696 0 1 2528
box 4 4 48 48
<< end >>
