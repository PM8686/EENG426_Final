magic
tech sky130l
timestamp 1731220555
<< m1 >>
rect 1136 3999 1140 4015
rect 296 3967 300 3995
rect 1072 3695 1076 3711
rect 2336 3671 2340 3707
rect 384 3235 388 3287
rect 1336 3207 1340 3335
rect 3872 2899 3876 2935
rect 1336 2551 1340 2571
rect 2424 2551 2428 2571
rect 1184 2295 1188 2411
rect 1176 2275 1180 2291
rect 3760 2275 3764 2395
rect 2192 2235 2196 2251
rect 1256 2107 1260 2123
rect 232 1947 236 1963
rect 2976 1891 2980 1923
rect 3392 1907 3396 1923
rect 232 1783 236 1799
rect 560 1763 564 1799
rect 1368 1651 1372 1667
rect 2672 1275 2676 1311
rect 232 995 236 1123
rect 2504 1115 2508 1147
rect 2424 951 2428 983
rect 3568 967 3572 983
rect 1216 859 1220 907
rect 3056 815 3060 931
rect 744 487 748 531
rect 1104 515 1108 531
rect 824 487 828 511
rect 3584 499 3588 515
rect 3104 355 3108 411
rect 1768 151 1772 203
rect 2768 191 2772 207
rect 2856 151 2860 195
rect 3496 159 3500 207
<< m2c >>
rect 1136 4015 1140 4019
rect 296 3995 300 3999
rect 400 3995 404 3999
rect 504 3995 508 3999
rect 608 3995 612 3999
rect 712 3995 716 3999
rect 816 3995 820 3999
rect 920 3995 924 3999
rect 1024 3995 1028 3999
rect 1128 3995 1132 3999
rect 1136 3995 1140 3999
rect 1232 3995 1236 3999
rect 1248 3995 1252 3999
rect 1336 3995 1340 3999
rect 1352 3995 1356 3999
rect 1440 3995 1444 3999
rect 1456 3995 1460 3999
rect 1544 3995 1548 3999
rect 2336 3995 2340 3999
rect 2352 3995 2356 3999
rect 2440 3995 2444 3999
rect 2544 3995 2548 3999
rect 2648 3995 2652 3999
rect 2664 3995 2668 3999
rect 2752 3995 2756 3999
rect 248 3979 252 3983
rect 2304 3983 2308 3987
rect 2464 3983 2468 3987
rect 2624 3983 2628 3987
rect 2776 3983 2780 3987
rect 2920 3983 2924 3987
rect 2968 3983 2972 3987
rect 3056 3983 3060 3987
rect 3104 3983 3108 3987
rect 3192 3983 3196 3987
rect 3232 3983 3236 3987
rect 3320 3983 3324 3987
rect 3352 3983 3356 3987
rect 3440 3983 3444 3987
rect 3464 3983 3468 3987
rect 3552 3983 3556 3987
rect 3584 3983 3588 3987
rect 3672 3983 3676 3987
rect 3704 3983 3708 3987
rect 3792 3983 3796 3987
rect 3824 3983 3828 3987
rect 3912 3983 3916 3987
rect 368 3979 372 3983
rect 456 3979 460 3983
rect 576 3979 580 3983
rect 664 3979 668 3983
rect 776 3979 780 3983
rect 864 3979 868 3983
rect 1056 3979 1060 3983
rect 1152 3979 1156 3983
rect 1240 3979 1244 3983
rect 1416 3979 1420 3983
rect 1592 3979 1596 3983
rect 1688 3979 1692 3983
rect 1776 3979 1780 3983
rect 296 3963 300 3967
rect 2296 3851 2300 3855
rect 2528 3851 2532 3855
rect 2656 3851 2660 3855
rect 2744 3851 2748 3855
rect 2952 3851 2956 3855
rect 3056 3851 3060 3855
rect 3144 3851 3148 3855
rect 3232 3851 3236 3855
rect 3320 3851 3324 3855
rect 3400 3851 3404 3855
rect 3488 3851 3492 3855
rect 3656 3851 3660 3855
rect 3824 3851 3828 3855
rect 432 3847 436 3851
rect 536 3847 540 3851
rect 624 3847 628 3851
rect 720 3847 724 3851
rect 808 3847 812 3851
rect 904 3847 908 3851
rect 992 3847 996 3851
rect 1160 3847 1164 3851
rect 1232 3847 1236 3851
rect 1320 3847 1324 3851
rect 1384 3847 1388 3851
rect 1472 3847 1476 3851
rect 1616 3847 1620 3851
rect 1752 3847 1756 3851
rect 1888 3847 1892 3851
rect 2008 3847 2012 3851
rect 2264 3839 2268 3843
rect 2560 3839 2564 3843
rect 2832 3839 2836 3843
rect 2984 3839 2988 3843
rect 3072 3841 3076 3845
rect 3288 3839 3292 3843
rect 3480 3839 3484 3843
rect 3568 3839 3572 3843
rect 3656 3839 3660 3843
rect 3968 3839 3972 3843
rect 656 3835 660 3839
rect 720 3835 724 3839
rect 808 3835 812 3839
rect 872 3835 876 3839
rect 960 3835 964 3839
rect 1016 3835 1020 3839
rect 1104 3835 1108 3839
rect 1248 3835 1252 3839
rect 1296 3835 1300 3839
rect 1384 3835 1388 3839
rect 1432 3835 1436 3839
rect 1520 3835 1524 3839
rect 1560 3835 1564 3839
rect 1648 3835 1652 3839
rect 1688 3835 1692 3839
rect 1776 3835 1780 3839
rect 1816 3835 1820 3839
rect 1904 3835 1908 3839
rect 1920 3835 1924 3839
rect 2008 3835 2012 3839
rect 1072 3711 1076 3715
rect 2184 3707 2188 3711
rect 2320 3707 2324 3711
rect 2336 3707 2340 3711
rect 2408 3707 2412 3711
rect 2632 3707 2636 3711
rect 2848 3707 2852 3711
rect 3048 3707 3052 3711
rect 3144 3707 3148 3711
rect 3232 3707 3236 3711
rect 3312 3707 3316 3711
rect 3400 3707 3404 3711
rect 3464 3707 3468 3711
rect 3552 3707 3556 3711
rect 3696 3707 3700 3711
rect 3752 3707 3756 3711
rect 3840 3707 3844 3711
rect 3880 3707 3884 3711
rect 3968 3707 3972 3711
rect 672 3691 676 3695
rect 704 3691 708 3695
rect 792 3691 796 3695
rect 920 3691 924 3695
rect 1056 3691 1060 3695
rect 1072 3691 1076 3695
rect 1184 3691 1188 3695
rect 1312 3691 1316 3695
rect 1352 3691 1356 3695
rect 1440 3691 1444 3695
rect 1480 3691 1484 3695
rect 1568 3691 1572 3695
rect 1616 3691 1620 3695
rect 1704 3691 1708 3695
rect 1752 3691 1756 3695
rect 1840 3691 1844 3695
rect 2184 3683 2188 3687
rect 2328 3683 2332 3687
rect 544 3675 548 3679
rect 600 3675 604 3679
rect 688 3675 692 3679
rect 832 3675 836 3679
rect 888 3675 892 3679
rect 976 3675 980 3679
rect 1120 3675 1124 3679
rect 1176 3675 1180 3679
rect 1264 3675 1268 3679
rect 1320 3675 1324 3679
rect 1408 3675 1412 3679
rect 1464 3675 1468 3679
rect 1552 3675 1556 3679
rect 2512 3683 2516 3687
rect 2608 3683 2612 3687
rect 2696 3683 2700 3687
rect 2800 3683 2804 3687
rect 2888 3683 2892 3687
rect 3080 3683 3084 3687
rect 3184 3683 3188 3687
rect 3272 3683 3276 3687
rect 3376 3683 3380 3687
rect 3464 3683 3468 3687
rect 3568 3683 3572 3687
rect 3656 3683 3660 3687
rect 2336 3667 2340 3671
rect 320 3543 324 3547
rect 360 3543 364 3547
rect 448 3543 452 3547
rect 592 3543 596 3547
rect 752 3543 756 3547
rect 832 3543 836 3547
rect 920 3543 924 3547
rect 1096 3543 1100 3547
rect 1192 3543 1196 3547
rect 1280 3543 1284 3547
rect 1376 3543 1380 3547
rect 1464 3543 1468 3547
rect 1648 3543 1652 3547
rect 1840 3543 1844 3547
rect 2008 3543 2012 3547
rect 2432 3539 2436 3543
rect 2656 3539 2660 3543
rect 2872 3539 2876 3543
rect 2992 3539 2996 3543
rect 3080 3539 3084 3543
rect 3200 3539 3204 3543
rect 3288 3539 3292 3543
rect 3416 3539 3420 3543
rect 3504 3539 3508 3543
rect 2512 3523 2516 3527
rect 2560 3523 2564 3527
rect 2648 3523 2652 3527
rect 2776 3523 2780 3527
rect 2816 3523 2820 3527
rect 2904 3523 2908 3527
rect 2936 3523 2940 3527
rect 3024 3523 3028 3527
rect 3056 3523 3060 3527
rect 3144 3523 3148 3527
rect 3184 3523 3188 3527
rect 3272 3523 3276 3527
rect 3312 3523 3316 3527
rect 3400 3523 3404 3527
rect 224 3519 228 3523
rect 248 3519 252 3523
rect 336 3519 340 3523
rect 472 3519 476 3523
rect 528 3519 532 3523
rect 616 3519 620 3523
rect 672 3519 676 3523
rect 760 3519 764 3523
rect 904 3519 908 3523
rect 952 3519 956 3523
rect 1040 3519 1044 3523
rect 1168 3519 1172 3523
rect 1296 3519 1300 3523
rect 1416 3519 1420 3523
rect 1536 3519 1540 3523
rect 1656 3519 1660 3523
rect 1696 3519 1700 3523
rect 1784 3519 1788 3523
rect 2432 3391 2436 3395
rect 2536 3391 2540 3395
rect 2640 3391 2644 3395
rect 2656 3391 2660 3395
rect 2744 3391 2748 3395
rect 2760 3391 2764 3395
rect 2848 3391 2852 3395
rect 2864 3391 2868 3395
rect 2952 3391 2956 3395
rect 2968 3391 2972 3395
rect 3056 3391 3060 3395
rect 3072 3391 3076 3395
rect 3160 3391 3164 3395
rect 3176 3391 3180 3395
rect 3264 3391 3268 3395
rect 224 3387 228 3391
rect 496 3387 500 3391
rect 728 3387 732 3391
rect 816 3387 820 3391
rect 1056 3387 1060 3391
rect 1144 3387 1148 3391
rect 1472 3387 1476 3391
rect 224 3351 228 3355
rect 304 3351 308 3355
rect 392 3351 396 3355
rect 512 3351 516 3355
rect 600 3351 604 3355
rect 728 3351 732 3355
rect 816 3351 820 3355
rect 944 3351 948 3355
rect 1032 3351 1036 3355
rect 1240 3351 1244 3355
rect 1352 3351 1356 3355
rect 1440 3351 1444 3355
rect 1544 3351 1548 3355
rect 1632 3351 1636 3355
rect 1736 3351 1740 3355
rect 1824 3351 1828 3355
rect 1920 3351 1924 3355
rect 2008 3351 2012 3355
rect 2512 3351 2516 3355
rect 2616 3351 2620 3355
rect 2720 3351 2724 3355
rect 2824 3351 2828 3355
rect 2928 3351 2932 3355
rect 2944 3351 2948 3355
rect 3032 3351 3036 3355
rect 1336 3335 1340 3339
rect 384 3287 388 3291
rect 384 3231 388 3235
rect 384 3211 388 3215
rect 464 3211 468 3215
rect 552 3211 556 3215
rect 640 3211 644 3215
rect 728 3211 732 3215
rect 832 3211 836 3215
rect 920 3211 924 3215
rect 1024 3211 1028 3215
rect 1112 3211 1116 3215
rect 1304 3211 1308 3215
rect 2600 3219 2604 3223
rect 2704 3219 2708 3223
rect 2720 3219 2724 3223
rect 2808 3219 2812 3223
rect 2824 3219 2828 3223
rect 2912 3219 2916 3223
rect 3016 3219 3020 3223
rect 3120 3219 3124 3223
rect 3224 3219 3228 3223
rect 3240 3219 3244 3223
rect 3328 3219 3332 3223
rect 1416 3211 1420 3215
rect 1504 3211 1508 3215
rect 1616 3211 1620 3215
rect 1704 3211 1708 3215
rect 1904 3211 1908 3215
rect 2472 3207 2476 3211
rect 2536 3207 2540 3211
rect 2624 3207 2628 3211
rect 2680 3207 2684 3211
rect 2768 3207 2772 3211
rect 2912 3207 2916 3211
rect 2960 3207 2964 3211
rect 3048 3207 3052 3211
rect 3096 3207 3100 3211
rect 3184 3207 3188 3211
rect 3320 3207 3324 3211
rect 3376 3207 3380 3211
rect 3464 3207 3468 3211
rect 1336 3203 1340 3207
rect 696 3195 700 3199
rect 744 3195 748 3199
rect 832 3195 836 3199
rect 888 3195 892 3199
rect 976 3195 980 3199
rect 1040 3195 1044 3199
rect 1128 3195 1132 3199
rect 1280 3195 1284 3199
rect 1424 3195 1428 3199
rect 1576 3195 1580 3199
rect 1728 3195 1732 3199
rect 1792 3195 1796 3199
rect 1880 3195 1884 3199
rect 1920 3195 1924 3199
rect 2008 3195 2012 3199
rect 672 3063 676 3067
rect 776 3063 780 3067
rect 880 3063 884 3067
rect 984 3063 988 3067
rect 1112 3063 1116 3067
rect 1168 3063 1172 3067
rect 1256 3063 1260 3067
rect 1344 3063 1348 3067
rect 1432 3063 1436 3067
rect 1536 3063 1540 3067
rect 1624 3063 1628 3067
rect 1736 3063 1740 3067
rect 1824 3063 1828 3067
rect 2008 3063 2012 3067
rect 2096 3063 2100 3067
rect 2184 3063 2188 3067
rect 2416 3063 2420 3067
rect 2656 3063 2660 3067
rect 2872 3063 2876 3067
rect 2984 3063 2988 3067
rect 3072 3063 3076 3067
rect 3176 3063 3180 3067
rect 3264 3063 3268 3067
rect 3448 3063 3452 3067
rect 3640 3063 3644 3067
rect 2184 3047 2188 3051
rect 2248 3047 2252 3051
rect 2336 3047 2340 3051
rect 2440 3047 2444 3051
rect 2528 3047 2532 3051
rect 2728 3047 2732 3051
rect 2928 3047 2932 3051
rect 3128 3047 3132 3051
rect 3240 3047 3244 3051
rect 3328 3047 3332 3051
rect 3440 3047 3444 3051
rect 3528 3047 3532 3051
rect 3640 3047 3644 3051
rect 3728 3047 3732 3051
rect 384 3043 388 3047
rect 400 3043 404 3047
rect 488 3043 492 3047
rect 512 3043 516 3047
rect 600 3043 604 3047
rect 712 3043 716 3047
rect 736 3043 740 3047
rect 824 3043 828 3047
rect 936 3043 940 3047
rect 960 3043 964 3047
rect 1048 3043 1052 3047
rect 1080 3043 1084 3047
rect 1168 3043 1172 3047
rect 1288 3043 1292 3047
rect 1320 3043 1324 3047
rect 1408 3043 1412 3047
rect 3872 2935 3876 2939
rect 2592 2923 2596 2927
rect 2184 2915 2188 2919
rect 2344 2915 2348 2919
rect 2432 2915 2436 2919
rect 2680 2915 2684 2919
rect 2832 2915 2836 2919
rect 2920 2915 2924 2919
rect 3152 2915 3156 2919
rect 3376 2915 3380 2919
rect 3608 2915 3612 2919
rect 3840 2915 3844 2919
rect 224 2903 228 2907
rect 256 2903 260 2907
rect 344 2903 348 2907
rect 416 2903 420 2907
rect 504 2903 508 2907
rect 680 2903 684 2907
rect 768 2903 772 2907
rect 856 2903 860 2907
rect 1032 2903 1036 2907
rect 1208 2903 1212 2907
rect 1376 2903 1380 2907
rect 1544 2903 1548 2907
rect 1720 2903 1724 2907
rect 2184 2895 2188 2899
rect 2264 2895 2268 2899
rect 2352 2895 2356 2899
rect 2472 2895 2476 2899
rect 2560 2895 2564 2899
rect 2680 2895 2684 2899
rect 2768 2895 2772 2899
rect 2888 2895 2892 2899
rect 2976 2895 2980 2899
rect 3184 2895 3188 2899
rect 3288 2895 3292 2899
rect 3376 2895 3380 2899
rect 3480 2895 3484 2899
rect 3568 2895 3572 2899
rect 3672 2895 3676 2899
rect 3760 2895 3764 2899
rect 3864 2895 3868 2899
rect 3872 2895 3876 2899
rect 3952 2895 3956 2899
rect 224 2879 228 2883
rect 360 2879 364 2883
rect 520 2879 524 2883
rect 672 2879 676 2883
rect 744 2879 748 2883
rect 832 2879 836 2883
rect 912 2879 916 2883
rect 1000 2879 1004 2883
rect 1088 2879 1092 2883
rect 1176 2879 1180 2883
rect 1272 2879 1276 2883
rect 1360 2879 1364 2883
rect 1464 2879 1468 2883
rect 1552 2879 1556 2883
rect 1744 2879 1748 2883
rect 2216 2751 2220 2755
rect 2304 2751 2308 2755
rect 2392 2751 2396 2755
rect 2576 2751 2580 2755
rect 2768 2751 2772 2755
rect 2960 2751 2964 2755
rect 3152 2751 3156 2755
rect 3248 2751 3252 2755
rect 3336 2751 3340 2755
rect 3424 2751 3428 2755
rect 3512 2751 3516 2755
rect 3600 2751 3604 2755
rect 3688 2751 3692 2755
rect 3776 2751 3780 2755
rect 3864 2751 3868 2755
rect 224 2735 228 2739
rect 304 2735 308 2739
rect 392 2735 396 2739
rect 576 2735 580 2739
rect 760 2735 764 2739
rect 856 2735 860 2739
rect 944 2735 948 2739
rect 1128 2735 1132 2739
rect 1312 2735 1316 2739
rect 1504 2735 1508 2739
rect 1704 2735 1708 2739
rect 1904 2735 1908 2739
rect 2184 2727 2188 2731
rect 2352 2727 2356 2731
rect 2528 2727 2532 2731
rect 2624 2727 2628 2731
rect 2712 2727 2716 2731
rect 2800 2727 2804 2731
rect 2888 2727 2892 2731
rect 3056 2727 3060 2731
rect 3128 2727 3132 2731
rect 3216 2727 3220 2731
rect 3288 2727 3292 2731
rect 3376 2727 3380 2731
rect 3448 2727 3452 2731
rect 3536 2727 3540 2731
rect 3608 2727 3612 2731
rect 3696 2727 3700 2731
rect 256 2720 260 2724
rect 456 2719 460 2723
rect 656 2719 660 2723
rect 768 2719 772 2723
rect 856 2719 860 2723
rect 1056 2719 1060 2723
rect 1184 2719 1188 2723
rect 1272 2719 1276 2723
rect 1400 2719 1404 2723
rect 1488 2719 1492 2723
rect 1624 2719 1628 2723
rect 1712 2719 1716 2723
rect 1944 2719 1948 2723
rect 2184 2583 2188 2587
rect 2248 2583 2252 2587
rect 2336 2583 2340 2587
rect 2504 2583 2508 2587
rect 2584 2583 2588 2587
rect 2672 2583 2676 2587
rect 2824 2583 2828 2587
rect 2968 2583 2972 2587
rect 3024 2583 3028 2587
rect 3112 2583 3116 2587
rect 3160 2583 3164 2587
rect 3248 2583 3252 2587
rect 3296 2583 3300 2587
rect 3384 2583 3388 2587
rect 3440 2583 3444 2587
rect 3528 2583 3532 2587
rect 328 2579 332 2583
rect 408 2579 412 2583
rect 496 2579 500 2583
rect 672 2579 676 2583
rect 848 2579 852 2583
rect 944 2579 948 2583
rect 1032 2579 1036 2583
rect 1224 2579 1228 2583
rect 1328 2579 1332 2583
rect 1416 2579 1420 2583
rect 1520 2579 1524 2583
rect 1608 2579 1612 2583
rect 1800 2579 1804 2583
rect 1912 2579 1916 2583
rect 2000 2579 2004 2583
rect 1336 2571 1340 2575
rect 392 2563 396 2567
rect 520 2563 524 2567
rect 608 2563 612 2567
rect 816 2563 820 2567
rect 1024 2563 1028 2567
rect 1232 2563 1236 2567
rect 2424 2571 2428 2575
rect 1344 2563 1348 2567
rect 1432 2563 1436 2567
rect 1632 2563 1636 2567
rect 1832 2563 1836 2567
rect 2008 2563 2012 2567
rect 2096 2563 2100 2567
rect 2184 2563 2188 2567
rect 2344 2563 2348 2567
rect 1336 2547 1340 2551
rect 2432 2563 2436 2567
rect 2520 2563 2524 2567
rect 2688 2563 2692 2567
rect 2840 2563 2844 2567
rect 2896 2563 2900 2567
rect 2984 2563 2988 2567
rect 3032 2563 3036 2567
rect 3120 2563 3124 2567
rect 3168 2563 3172 2567
rect 3256 2563 3260 2567
rect 3304 2563 3308 2567
rect 3392 2563 3396 2567
rect 2424 2547 2428 2551
rect 352 2431 356 2435
rect 512 2431 516 2435
rect 680 2431 684 2435
rect 768 2431 772 2435
rect 856 2431 860 2435
rect 944 2431 948 2435
rect 1032 2431 1036 2435
rect 1200 2431 1204 2435
rect 1280 2431 1284 2435
rect 1368 2431 1372 2435
rect 1536 2431 1540 2435
rect 1696 2431 1700 2435
rect 1776 2431 1780 2435
rect 1864 2431 1868 2435
rect 1920 2431 1924 2435
rect 2008 2431 2012 2435
rect 2696 2419 2700 2423
rect 2728 2419 2732 2423
rect 2816 2419 2820 2423
rect 2944 2419 2948 2423
rect 3000 2419 3004 2423
rect 3088 2419 3092 2423
rect 3144 2419 3148 2423
rect 3232 2419 3236 2423
rect 3296 2419 3300 2423
rect 3384 2419 3388 2423
rect 3536 2419 3540 2423
rect 3600 2419 3604 2423
rect 3688 2419 3692 2423
rect 3840 2419 3844 2423
rect 3968 2419 3972 2423
rect 400 2411 404 2415
rect 456 2411 460 2415
rect 544 2411 548 2415
rect 608 2411 612 2415
rect 696 2411 700 2415
rect 856 2411 860 2415
rect 928 2411 932 2415
rect 1016 2411 1020 2415
rect 1168 2411 1172 2415
rect 1184 2411 1188 2415
rect 1320 2411 1324 2415
rect 1376 2411 1380 2415
rect 1464 2411 1468 2415
rect 1608 2411 1612 2415
rect 1656 2411 1660 2415
rect 1744 2411 1748 2415
rect 1888 2411 1892 2415
rect 2008 2411 2012 2415
rect 2560 2395 2564 2399
rect 2584 2395 2588 2399
rect 2672 2396 2676 2400
rect 2800 2395 2804 2399
rect 2952 2395 2956 2399
rect 3128 2395 3132 2399
rect 3232 2395 3236 2399
rect 3320 2395 3324 2399
rect 3440 2395 3444 2399
rect 3528 2395 3532 2399
rect 3752 2395 3756 2399
rect 3760 2395 3764 2399
rect 3968 2395 3972 2399
rect 1176 2291 1180 2295
rect 1184 2291 1188 2295
rect 432 2271 436 2275
rect 480 2271 484 2275
rect 568 2271 572 2275
rect 712 2271 716 2275
rect 856 2271 860 2275
rect 1008 2271 1012 2275
rect 1160 2271 1164 2275
rect 1176 2271 1180 2275
rect 1320 2271 1324 2275
rect 1488 2271 1492 2275
rect 1664 2271 1668 2275
rect 1848 2271 1852 2275
rect 2008 2271 2012 2275
rect 3760 2271 3764 2275
rect 2184 2251 2188 2255
rect 2192 2251 2196 2255
rect 2208 2251 2212 2255
rect 2296 2251 2300 2255
rect 2432 2251 2436 2255
rect 2584 2251 2588 2255
rect 2744 2251 2748 2255
rect 2920 2251 2924 2255
rect 3024 2251 3028 2255
rect 3112 2251 3116 2255
rect 3232 2251 3236 2255
rect 3320 2251 3324 2255
rect 3448 2251 3452 2255
rect 3536 2251 3540 2255
rect 3760 2251 3764 2255
rect 3968 2251 3972 2255
rect 312 2247 316 2251
rect 376 2247 380 2251
rect 464 2247 468 2251
rect 536 2247 540 2251
rect 624 2247 628 2251
rect 784 2247 788 2251
rect 856 2247 860 2251
rect 944 2247 948 2251
rect 1104 2247 1108 2251
rect 1176 2247 1180 2251
rect 1264 2247 1268 2251
rect 1344 2247 1348 2251
rect 1432 2247 1436 2251
rect 1600 2247 1604 2251
rect 1680 2247 1684 2251
rect 1768 2247 1772 2251
rect 2184 2231 2188 2235
rect 2192 2231 2196 2235
rect 2352 2231 2356 2235
rect 2464 2231 2468 2235
rect 2552 2231 2556 2235
rect 2664 2231 2668 2235
rect 2752 2231 2756 2235
rect 2952 2231 2956 2235
rect 3064 2231 3068 2235
rect 3152 2231 3156 2235
rect 3352 2231 3356 2235
rect 3560 2231 3564 2235
rect 3776 2231 3780 2235
rect 3968 2231 3972 2235
rect 1256 2123 1260 2127
rect 224 2103 228 2107
rect 392 2103 396 2107
rect 584 2103 588 2107
rect 776 2103 780 2107
rect 968 2103 972 2107
rect 1160 2103 1164 2107
rect 1256 2103 1260 2107
rect 1352 2103 1356 2107
rect 1536 2103 1540 2107
rect 1728 2103 1732 2107
rect 1832 2103 1836 2107
rect 1920 2103 1924 2107
rect 2216 2091 2220 2095
rect 2304 2091 2308 2095
rect 2392 2091 2396 2095
rect 2568 2091 2572 2095
rect 2664 2091 2668 2095
rect 2752 2091 2756 2095
rect 2848 2091 2852 2095
rect 2936 2091 2940 2095
rect 3112 2091 3116 2095
rect 3200 2091 3204 2095
rect 3288 2091 3292 2095
rect 3376 2091 3380 2095
rect 3464 2091 3468 2095
rect 3640 2091 3644 2095
rect 3728 2091 3732 2095
rect 3816 2091 3820 2095
rect 3968 2091 3972 2095
rect 224 2083 228 2087
rect 288 2083 292 2087
rect 376 2083 380 2087
rect 464 2083 468 2087
rect 552 2083 556 2087
rect 736 2083 740 2087
rect 832 2083 836 2087
rect 920 2083 924 2087
rect 1112 2083 1116 2087
rect 1224 2083 1228 2087
rect 1312 2083 1316 2087
rect 1432 2083 1436 2087
rect 1520 2083 1524 2087
rect 1736 2083 1740 2087
rect 1952 2083 1956 2087
rect 2280 2067 2284 2071
rect 2464 2067 2468 2071
rect 2648 2067 2652 2071
rect 2832 2067 2836 2071
rect 3008 2067 3012 2071
rect 3176 2067 3180 2071
rect 3336 2067 3340 2071
rect 3408 2067 3412 2071
rect 3496 2067 3500 2071
rect 3656 2067 3660 2071
rect 3824 2067 3828 2071
rect 3968 2067 3972 2071
rect 232 1963 236 1967
rect 224 1943 228 1947
rect 232 1943 236 1947
rect 376 1943 380 1947
rect 560 1943 564 1947
rect 760 1943 764 1947
rect 968 1943 972 1947
rect 1176 1943 1180 1947
rect 1384 1943 1388 1947
rect 1600 1943 1604 1947
rect 1728 1943 1732 1947
rect 1816 1943 1820 1947
rect 1920 1943 1924 1947
rect 2008 1943 2012 1947
rect 3752 1931 3756 1935
rect 2352 1923 2356 1927
rect 2536 1923 2540 1927
rect 2712 1923 2716 1927
rect 2800 1923 2804 1927
rect 2888 1923 2892 1927
rect 2968 1923 2972 1927
rect 2976 1923 2980 1927
rect 3056 1923 3060 1927
rect 3224 1923 3228 1927
rect 3384 1923 3388 1927
rect 3392 1923 3396 1927
rect 3448 1923 3452 1927
rect 3536 1923 3540 1927
rect 3688 1923 3692 1927
rect 3840 1923 3844 1927
rect 3968 1923 3972 1927
rect 224 1919 228 1923
rect 256 1919 260 1923
rect 344 1919 348 1923
rect 392 1919 396 1923
rect 480 1919 484 1923
rect 616 1919 620 1923
rect 752 1919 756 1923
rect 896 1919 900 1923
rect 968 1919 972 1923
rect 1056 1919 1060 1923
rect 1144 1919 1148 1923
rect 1232 1919 1236 1923
rect 1328 1919 1332 1923
rect 1416 1919 1420 1923
rect 1528 1919 1532 1923
rect 1616 1919 1620 1923
rect 1824 1919 1828 1923
rect 2008 1919 2012 1923
rect 2480 1903 2484 1907
rect 2640 1903 2644 1907
rect 2728 1903 2732 1907
rect 2960 1903 2964 1907
rect 3176 1903 3180 1907
rect 3296 1903 3300 1907
rect 3384 1903 3388 1907
rect 3392 1903 3396 1907
rect 3584 1903 3588 1907
rect 3784 1903 3788 1907
rect 3968 1903 3972 1907
rect 2976 1887 2980 1891
rect 232 1799 236 1803
rect 560 1799 564 1803
rect 224 1779 228 1783
rect 232 1779 236 1783
rect 360 1779 364 1783
rect 520 1779 524 1783
rect 672 1779 676 1783
rect 736 1779 740 1783
rect 824 1779 828 1783
rect 992 1779 996 1783
rect 1088 1779 1092 1783
rect 1176 1779 1180 1783
rect 1288 1779 1292 1783
rect 1376 1779 1380 1783
rect 1496 1779 1500 1783
rect 1584 1779 1588 1783
rect 1720 1779 1724 1783
rect 1808 1779 1812 1783
rect 2008 1779 2012 1783
rect 2184 1771 2188 1775
rect 2456 1771 2460 1775
rect 2720 1771 2724 1775
rect 2960 1771 2964 1775
rect 3080 1771 3084 1775
rect 3168 1771 3172 1775
rect 3360 1771 3364 1775
rect 3528 1771 3532 1775
rect 3688 1771 3692 1775
rect 3840 1771 3844 1775
rect 3968 1771 3972 1775
rect 280 1759 284 1763
rect 368 1759 372 1763
rect 456 1759 460 1763
rect 552 1759 556 1763
rect 560 1759 564 1763
rect 640 1759 644 1763
rect 824 1759 828 1763
rect 920 1759 924 1763
rect 1008 1759 1012 1763
rect 1184 1759 1188 1763
rect 1264 1759 1268 1763
rect 1352 1759 1356 1763
rect 1440 1759 1444 1763
rect 1528 1759 1532 1763
rect 1616 1759 1620 1763
rect 1704 1759 1708 1763
rect 2184 1759 2188 1763
rect 2360 1759 2364 1763
rect 2568 1759 2572 1763
rect 2784 1759 2788 1763
rect 2904 1759 2908 1763
rect 2992 1760 2996 1764
rect 3192 1759 3196 1763
rect 3304 1759 3308 1763
rect 3392 1759 3396 1763
rect 3584 1759 3588 1763
rect 3688 1759 3692 1763
rect 3776 1759 3780 1763
rect 3880 1759 3884 1763
rect 3968 1759 3972 1763
rect 1368 1667 1372 1671
rect 1368 1647 1372 1651
rect 376 1627 380 1631
rect 608 1627 612 1631
rect 840 1627 844 1631
rect 1056 1627 1060 1631
rect 1264 1627 1268 1631
rect 1368 1627 1372 1631
rect 1456 1627 1460 1631
rect 1552 1627 1556 1631
rect 1640 1627 1644 1631
rect 1728 1627 1732 1631
rect 1816 1627 1820 1631
rect 1912 1627 1916 1631
rect 2000 1627 2004 1631
rect 2184 1619 2188 1623
rect 2224 1619 2228 1623
rect 2312 1619 2316 1623
rect 2368 1619 2372 1623
rect 2456 1619 2460 1623
rect 2592 1619 2596 1623
rect 2640 1619 2644 1623
rect 2728 1619 2732 1623
rect 2864 1619 2868 1623
rect 3000 1619 3004 1623
rect 3136 1619 3140 1623
rect 3280 1619 3284 1623
rect 3336 1619 3340 1623
rect 3424 1619 3428 1623
rect 472 1611 476 1615
rect 560 1611 564 1615
rect 648 1611 652 1615
rect 736 1611 740 1615
rect 824 1611 828 1615
rect 1008 1611 1012 1615
rect 1096 1611 1100 1615
rect 1184 1611 1188 1615
rect 1352 1611 1356 1615
rect 1432 1611 1436 1615
rect 1520 1611 1524 1615
rect 1680 1611 1684 1615
rect 1840 1611 1844 1615
rect 2008 1611 2012 1615
rect 2240 1595 2244 1599
rect 2360 1595 2364 1599
rect 2480 1595 2484 1599
rect 2600 1595 2604 1599
rect 2720 1595 2724 1599
rect 2840 1595 2844 1599
rect 2960 1595 2964 1599
rect 2992 1595 2996 1599
rect 3080 1595 3084 1599
rect 3112 1595 3116 1599
rect 3200 1595 3204 1599
rect 3240 1595 3244 1599
rect 3328 1595 3332 1599
rect 576 1471 580 1475
rect 688 1471 692 1475
rect 808 1471 812 1475
rect 928 1471 932 1475
rect 1040 1471 1044 1475
rect 1152 1471 1156 1475
rect 1184 1471 1188 1475
rect 1272 1471 1276 1475
rect 1392 1471 1396 1475
rect 1512 1471 1516 1475
rect 1632 1471 1636 1475
rect 2424 1455 2428 1459
rect 2448 1455 2452 1459
rect 2536 1455 2540 1459
rect 2648 1455 2652 1459
rect 2680 1455 2684 1459
rect 2768 1455 2772 1459
rect 2888 1455 2892 1459
rect 3000 1455 3004 1459
rect 3120 1455 3124 1459
rect 3240 1455 3244 1459
rect 3360 1455 3364 1459
rect 3392 1455 3396 1459
rect 3480 1455 3484 1459
rect 656 1447 660 1451
rect 672 1447 676 1451
rect 760 1447 764 1451
rect 864 1447 868 1451
rect 968 1447 972 1451
rect 984 1447 988 1451
rect 1072 1447 1076 1451
rect 1088 1447 1092 1451
rect 1176 1447 1180 1451
rect 1280 1447 1284 1451
rect 1296 1447 1300 1451
rect 1384 1447 1388 1451
rect 1400 1447 1404 1451
rect 1488 1447 1492 1451
rect 1504 1447 1508 1451
rect 1592 1447 1596 1451
rect 2416 1431 2420 1435
rect 2432 1431 2436 1435
rect 2520 1431 2524 1435
rect 2552 1431 2556 1435
rect 2640 1431 2644 1435
rect 2768 1431 2772 1435
rect 2824 1431 2828 1435
rect 2912 1431 2916 1435
rect 3064 1431 3068 1435
rect 3128 1431 3132 1435
rect 3216 1431 3220 1435
rect 3376 1431 3380 1435
rect 3544 1431 3548 1435
rect 3720 1431 3724 1435
rect 3896 1431 3900 1435
rect 2672 1311 2676 1315
rect 624 1307 628 1311
rect 640 1307 644 1311
rect 728 1307 732 1311
rect 744 1307 748 1311
rect 832 1307 836 1311
rect 848 1307 852 1311
rect 936 1307 940 1311
rect 960 1307 964 1311
rect 1048 1307 1052 1311
rect 1160 1307 1164 1311
rect 1184 1307 1188 1311
rect 1272 1307 1276 1311
rect 1384 1307 1388 1311
rect 1416 1307 1420 1311
rect 1504 1307 1508 1311
rect 1536 1307 1540 1311
rect 1624 1307 1628 1311
rect 416 1291 420 1295
rect 448 1291 452 1295
rect 536 1291 540 1295
rect 584 1291 588 1295
rect 672 1291 676 1295
rect 728 1291 732 1295
rect 816 1291 820 1295
rect 888 1291 892 1295
rect 976 1291 980 1295
rect 1136 1291 1140 1295
rect 1304 1291 1308 1295
rect 1480 1291 1484 1295
rect 1656 1291 1660 1295
rect 2360 1291 2364 1295
rect 2480 1291 2484 1295
rect 2616 1291 2620 1295
rect 2768 1291 2772 1295
rect 2928 1291 2932 1295
rect 3088 1291 3092 1295
rect 3256 1291 3260 1295
rect 3336 1291 3340 1295
rect 3424 1291 3428 1295
rect 3504 1291 3508 1295
rect 3592 1291 3596 1295
rect 3672 1291 3676 1295
rect 3760 1291 3764 1295
rect 3928 1291 3932 1295
rect 2200 1271 2204 1275
rect 2280 1271 2284 1275
rect 2368 1271 2372 1275
rect 2464 1271 2468 1275
rect 2552 1271 2556 1275
rect 2664 1271 2668 1275
rect 2672 1271 2676 1275
rect 2752 1271 2756 1275
rect 2952 1271 2956 1275
rect 3144 1271 3148 1275
rect 3320 1271 3324 1275
rect 3488 1271 3492 1275
rect 3656 1271 3660 1275
rect 3824 1271 3828 1275
rect 3968 1271 3972 1275
rect 256 1159 260 1163
rect 336 1159 340 1163
rect 424 1159 428 1163
rect 520 1159 524 1163
rect 608 1159 612 1163
rect 712 1159 716 1163
rect 800 1159 804 1163
rect 904 1159 908 1163
rect 992 1159 996 1163
rect 1176 1159 1180 1163
rect 1360 1159 1364 1163
rect 1456 1159 1460 1163
rect 1544 1159 1548 1163
rect 1640 1159 1644 1163
rect 1728 1159 1732 1163
rect 1824 1159 1828 1163
rect 1912 1159 1916 1163
rect 2504 1147 2508 1151
rect 224 1139 228 1143
rect 288 1139 292 1143
rect 376 1139 380 1143
rect 480 1139 484 1143
rect 568 1139 572 1143
rect 688 1139 692 1143
rect 776 1139 780 1143
rect 896 1139 900 1143
rect 984 1139 988 1143
rect 1192 1139 1196 1143
rect 1392 1139 1396 1143
rect 1592 1139 1596 1143
rect 1792 1139 1796 1143
rect 1992 1139 1996 1143
rect 2184 1128 2188 1132
rect 2320 1127 2324 1131
rect 2480 1127 2484 1131
rect 232 1123 236 1127
rect 224 999 228 1003
rect 2632 1127 2636 1131
rect 2688 1127 2692 1131
rect 2776 1127 2780 1131
rect 2936 1127 2940 1131
rect 3024 1127 3028 1131
rect 3112 1127 3116 1131
rect 3224 1127 3228 1131
rect 3312 1127 3316 1131
rect 3440 1127 3444 1131
rect 3528 1127 3532 1131
rect 3672 1127 3676 1131
rect 3760 1127 3764 1131
rect 3968 1127 3972 1131
rect 2184 1111 2188 1115
rect 2288 1111 2292 1115
rect 2376 1111 2380 1115
rect 2496 1111 2500 1115
rect 2504 1111 2508 1115
rect 2584 1111 2588 1115
rect 2776 1111 2780 1115
rect 2968 1111 2972 1115
rect 3072 1111 3076 1115
rect 3160 1111 3164 1115
rect 3272 1111 3276 1115
rect 3360 1111 3364 1115
rect 3480 1111 3484 1115
rect 3568 1111 3572 1115
rect 3688 1111 3692 1115
rect 3776 1111 3780 1115
rect 3968 1111 3972 1115
rect 264 999 268 1003
rect 352 999 356 1003
rect 432 999 436 1003
rect 520 999 524 1003
rect 608 999 612 1003
rect 696 999 700 1003
rect 784 999 788 1003
rect 872 999 876 1003
rect 1040 999 1044 1003
rect 1200 999 1204 1003
rect 1352 999 1356 1003
rect 1408 999 1412 1003
rect 1496 999 1500 1003
rect 1544 999 1548 1003
rect 1632 999 1636 1003
rect 1680 999 1684 1003
rect 1768 999 1772 1003
rect 1808 999 1812 1003
rect 1896 999 1900 1003
rect 1920 999 1924 1003
rect 2008 999 2012 1003
rect 232 991 236 995
rect 2424 983 2428 987
rect 224 975 228 979
rect 360 975 364 979
rect 544 975 548 979
rect 744 975 748 979
rect 856 975 860 979
rect 944 975 948 979
rect 1064 975 1068 979
rect 1152 975 1156 979
rect 1272 975 1276 979
rect 1360 975 1364 979
rect 1480 975 1484 979
rect 1568 975 1572 979
rect 1776 975 1780 979
rect 1984 975 1988 979
rect 2392 963 2396 967
rect 3568 983 3572 987
rect 2472 963 2476 967
rect 2560 963 2564 967
rect 2648 963 2652 967
rect 2736 963 2740 967
rect 2920 963 2924 967
rect 3024 963 3028 967
rect 3112 963 3116 967
rect 3320 963 3324 967
rect 3536 963 3540 967
rect 3568 963 3572 967
rect 3760 963 3764 967
rect 3968 963 3972 967
rect 2224 947 2228 951
rect 2272 947 2276 951
rect 2360 947 2364 951
rect 2416 947 2420 951
rect 2424 947 2428 951
rect 2504 947 2508 951
rect 2664 947 2668 951
rect 2744 947 2748 951
rect 2832 947 2836 951
rect 3008 947 3012 951
rect 3192 947 3196 951
rect 3296 947 3300 951
rect 3384 947 3388 951
rect 3496 947 3500 951
rect 3584 947 3588 951
rect 3696 947 3700 951
rect 3784 947 3788 951
rect 3968 947 3972 951
rect 3056 931 3060 935
rect 1216 907 1220 911
rect 1216 855 1220 859
rect 224 835 228 839
rect 304 835 308 839
rect 392 835 396 839
rect 504 835 508 839
rect 592 835 596 839
rect 800 835 804 839
rect 920 835 924 839
rect 1008 835 1012 839
rect 1216 835 1220 839
rect 1320 835 1324 839
rect 1408 835 1412 839
rect 1512 835 1516 839
rect 1600 835 1604 839
rect 1704 835 1708 839
rect 1792 835 1796 839
rect 1896 835 1900 839
rect 1984 835 1988 839
rect 336 811 340 815
rect 352 811 356 815
rect 440 811 444 815
rect 464 811 468 815
rect 552 811 556 815
rect 576 811 580 815
rect 664 811 668 815
rect 696 811 700 815
rect 784 811 788 815
rect 928 811 932 815
rect 1016 811 1020 815
rect 1104 811 1108 815
rect 1224 811 1228 815
rect 1312 811 1316 815
rect 1456 811 1460 815
rect 1544 811 1548 815
rect 1696 811 1700 815
rect 1784 811 1788 815
rect 2008 811 2012 815
rect 3056 811 3060 815
rect 2184 803 2188 807
rect 2224 803 2228 807
rect 2312 803 2316 807
rect 2480 803 2484 807
rect 2648 803 2652 807
rect 2824 803 2828 807
rect 2920 803 2924 807
rect 3008 803 3012 807
rect 3104 803 3108 807
rect 3192 803 3196 807
rect 3384 803 3388 807
rect 3584 803 3588 807
rect 3784 803 3788 807
rect 3968 803 3972 807
rect 2096 791 2100 795
rect 2184 791 2188 795
rect 2464 791 2468 795
rect 2752 791 2756 795
rect 3024 791 3028 795
rect 3272 791 3276 795
rect 3424 791 3428 795
rect 3512 791 3516 795
rect 3656 791 3660 795
rect 3744 791 3748 795
rect 3968 791 3972 795
rect 496 675 500 679
rect 600 675 604 679
rect 712 675 716 679
rect 832 675 836 679
rect 952 675 956 679
rect 1080 675 1084 679
rect 1128 675 1132 679
rect 1216 675 1220 679
rect 1272 675 1276 679
rect 1360 675 1364 679
rect 1432 675 1436 679
rect 1520 675 1524 679
rect 1600 675 1604 679
rect 1688 675 1692 679
rect 1856 675 1860 679
rect 2008 675 2012 679
rect 664 651 668 655
rect 680 651 684 655
rect 768 651 772 655
rect 792 651 796 655
rect 880 653 884 657
rect 992 651 996 655
rect 1016 651 1020 655
rect 1104 651 1108 655
rect 1216 651 1220 655
rect 1248 651 1252 655
rect 1336 651 1340 655
rect 1368 651 1372 655
rect 1456 651 1460 655
rect 1488 651 1492 655
rect 1576 651 1580 655
rect 1608 651 1612 655
rect 1696 651 1700 655
rect 2184 651 2188 655
rect 2400 651 2404 655
rect 2536 651 2540 655
rect 2624 651 2628 655
rect 2760 651 2764 655
rect 2848 651 2852 655
rect 3064 651 3068 655
rect 3280 651 3284 655
rect 3488 651 3492 655
rect 3608 651 3612 655
rect 3696 651 3700 655
rect 3904 651 3908 655
rect 2200 635 2204 639
rect 2368 635 2372 639
rect 2528 635 2532 639
rect 2688 635 2692 639
rect 2768 635 2772 639
rect 2856 635 2860 639
rect 3024 635 3028 639
rect 3112 635 3116 639
rect 3200 635 3204 639
rect 3376 635 3380 639
rect 3560 635 3564 639
rect 3752 635 3756 639
rect 3952 636 3956 640
rect 744 531 748 535
rect 736 511 740 515
rect 1104 531 1108 535
rect 3584 515 3588 519
rect 824 511 828 515
rect 848 511 852 515
rect 880 511 884 515
rect 968 511 972 515
rect 1096 511 1100 515
rect 1104 511 1108 515
rect 1232 511 1236 515
rect 1376 511 1380 515
rect 1520 511 1524 515
rect 1576 511 1580 515
rect 1664 511 1668 515
rect 1720 511 1724 515
rect 1808 511 1812 515
rect 1864 511 1868 515
rect 1952 511 1956 515
rect 2376 495 2380 499
rect 2432 495 2436 499
rect 2520 495 2524 499
rect 2664 495 2668 499
rect 2808 495 2812 499
rect 2952 495 2956 499
rect 3104 495 3108 499
rect 3168 495 3172 499
rect 3256 495 3260 499
rect 3320 495 3324 499
rect 3408 495 3412 499
rect 3568 495 3572 499
rect 3584 495 3588 499
rect 3728 495 3732 499
rect 3896 495 3900 499
rect 608 483 612 487
rect 624 483 628 487
rect 712 483 716 487
rect 728 483 732 487
rect 744 483 748 487
rect 816 483 820 487
rect 824 483 828 487
rect 832 483 836 487
rect 920 483 924 487
rect 952 483 956 487
rect 1040 483 1044 487
rect 1176 483 1180 487
rect 1240 483 1244 487
rect 1328 483 1332 487
rect 1488 483 1492 487
rect 1576 483 1580 487
rect 1664 483 1668 487
rect 1848 483 1852 487
rect 2008 483 2012 487
rect 2584 475 2588 479
rect 2600 475 2604 479
rect 2688 475 2692 479
rect 2720 475 2724 479
rect 2808 475 2812 479
rect 2936 475 2940 479
rect 2992 475 2996 479
rect 3080 475 3084 479
rect 3144 475 3148 479
rect 3232 475 3236 479
rect 3304 475 3308 479
rect 3392 475 3396 479
rect 3552 475 3556 479
rect 3632 475 3636 479
rect 3720 475 3724 479
rect 3896 475 3900 479
rect 3104 411 3108 415
rect 3104 351 3108 355
rect 568 347 572 351
rect 704 347 708 351
rect 840 347 844 351
rect 984 347 988 351
rect 1120 347 1124 351
rect 1256 347 1260 351
rect 1304 347 1308 351
rect 1392 347 1396 351
rect 1520 347 1524 351
rect 1648 347 1652 351
rect 1776 347 1780 351
rect 1904 347 1908 351
rect 1920 347 1924 351
rect 2008 347 2012 351
rect 2576 331 2580 335
rect 2664 331 2668 335
rect 2680 331 2684 335
rect 2768 331 2772 335
rect 2800 331 2804 335
rect 2888 331 2892 335
rect 3032 331 3036 335
rect 3104 331 3108 335
rect 3192 331 3196 335
rect 3288 331 3292 335
rect 3376 331 3380 335
rect 3488 331 3492 335
rect 3576 331 3580 335
rect 3784 331 3788 335
rect 3968 331 3972 335
rect 408 323 412 327
rect 448 323 452 327
rect 536 323 540 327
rect 592 323 596 327
rect 680 323 684 327
rect 752 323 756 327
rect 840 323 844 327
rect 1016 323 1020 327
rect 1112 323 1116 327
rect 1200 323 1204 327
rect 1296 323 1300 327
rect 1384 323 1388 327
rect 1576 323 1580 327
rect 1688 323 1692 327
rect 1776 323 1780 327
rect 1976 323 1980 327
rect 2096 319 2100 323
rect 2184 319 2188 323
rect 2256 319 2260 323
rect 2344 319 2348 323
rect 2528 319 2532 323
rect 2704 319 2708 323
rect 2880 319 2884 323
rect 2984 319 2988 323
rect 3072 319 3076 323
rect 3200 319 3204 323
rect 3288 319 3292 323
rect 3424 319 3428 323
rect 3512 319 3516 323
rect 3664 319 3668 323
rect 3752 319 3756 323
rect 3968 319 3972 323
rect 2768 207 2772 211
rect 1768 203 1772 207
rect 224 183 228 187
rect 264 183 268 187
rect 352 183 356 187
rect 416 183 420 187
rect 504 183 508 187
rect 584 183 588 187
rect 672 183 676 187
rect 768 183 772 187
rect 856 183 860 187
rect 1048 183 1052 187
rect 1248 183 1252 187
rect 1448 183 1452 187
rect 1656 183 1660 187
rect 3496 207 3500 211
rect 2184 187 2188 191
rect 2344 187 2348 191
rect 2544 187 2548 191
rect 2760 187 2764 191
rect 2768 187 2772 191
rect 2856 195 2860 199
rect 2888 195 2892 199
rect 1784 183 1788 187
rect 1872 183 1876 187
rect 2976 187 2980 191
rect 3184 187 3188 191
rect 3392 187 3396 191
rect 3504 187 3508 191
rect 3592 187 3596 191
rect 3704 187 3708 191
rect 3792 187 3796 191
rect 3968 187 3972 191
rect 3496 155 3500 159
rect 224 147 228 151
rect 240 147 244 151
rect 328 147 332 151
rect 344 147 348 151
rect 432 147 436 151
rect 456 147 460 151
rect 544 147 548 151
rect 592 147 596 151
rect 680 147 684 151
rect 728 147 732 151
rect 816 147 820 151
rect 864 147 868 151
rect 952 147 956 151
rect 1088 147 1092 151
rect 1136 147 1140 151
rect 1224 147 1228 151
rect 1264 147 1268 151
rect 1352 147 1356 151
rect 1384 147 1388 151
rect 1472 147 1476 151
rect 1504 147 1508 151
rect 1592 147 1596 151
rect 1632 147 1636 151
rect 1720 147 1724 151
rect 1760 147 1764 151
rect 1768 147 1772 151
rect 1848 147 1852 151
rect 2184 147 2188 151
rect 2200 147 2204 151
rect 2288 147 2292 151
rect 2304 147 2308 151
rect 2392 147 2396 151
rect 2408 147 2412 151
rect 2496 147 2500 151
rect 2512 147 2516 151
rect 2600 147 2604 151
rect 2640 147 2644 151
rect 2728 147 2732 151
rect 2760 147 2764 151
rect 2848 147 2852 151
rect 2856 147 2860 151
rect 2968 147 2972 151
rect 3000 147 3004 151
rect 3088 147 3092 151
rect 3120 147 3124 151
rect 3208 147 3212 151
rect 3232 147 3236 151
rect 3320 147 3324 151
rect 3344 147 3348 151
rect 3432 147 3436 151
rect 3456 147 3460 151
rect 3544 147 3548 151
rect 3568 147 3572 151
rect 3656 147 3660 151
rect 3672 147 3676 151
rect 3760 147 3764 151
rect 3864 147 3868 151
rect 3880 147 3884 151
rect 3968 147 3972 151
<< m2 >>
rect 326 4050 332 4051
rect 326 4046 327 4050
rect 331 4046 332 4050
rect 110 4045 116 4046
rect 326 4045 332 4046
rect 430 4050 436 4051
rect 430 4046 431 4050
rect 435 4046 436 4050
rect 430 4045 436 4046
rect 534 4050 540 4051
rect 534 4046 535 4050
rect 539 4046 540 4050
rect 534 4045 540 4046
rect 638 4050 644 4051
rect 638 4046 639 4050
rect 643 4046 644 4050
rect 638 4045 644 4046
rect 742 4050 748 4051
rect 742 4046 743 4050
rect 747 4046 748 4050
rect 742 4045 748 4046
rect 846 4050 852 4051
rect 846 4046 847 4050
rect 851 4046 852 4050
rect 846 4045 852 4046
rect 950 4050 956 4051
rect 950 4046 951 4050
rect 955 4046 956 4050
rect 950 4045 956 4046
rect 1054 4050 1060 4051
rect 1054 4046 1055 4050
rect 1059 4046 1060 4050
rect 1054 4045 1060 4046
rect 1158 4050 1164 4051
rect 1158 4046 1159 4050
rect 1163 4046 1164 4050
rect 1158 4045 1164 4046
rect 1262 4050 1268 4051
rect 1262 4046 1263 4050
rect 1267 4046 1268 4050
rect 1262 4045 1268 4046
rect 1366 4050 1372 4051
rect 1366 4046 1367 4050
rect 1371 4046 1372 4050
rect 1366 4045 1372 4046
rect 1470 4050 1476 4051
rect 1470 4046 1471 4050
rect 1475 4046 1476 4050
rect 2262 4050 2268 4051
rect 2262 4046 2263 4050
rect 2267 4046 2268 4050
rect 1470 4045 1476 4046
rect 2030 4045 2036 4046
rect 110 4041 111 4045
rect 115 4041 116 4045
rect 110 4040 116 4041
rect 2030 4041 2031 4045
rect 2035 4041 2036 4045
rect 2030 4040 2036 4041
rect 2070 4045 2076 4046
rect 2262 4045 2268 4046
rect 2366 4050 2372 4051
rect 2366 4046 2367 4050
rect 2371 4046 2372 4050
rect 2366 4045 2372 4046
rect 2470 4050 2476 4051
rect 2470 4046 2471 4050
rect 2475 4046 2476 4050
rect 2470 4045 2476 4046
rect 2574 4050 2580 4051
rect 2574 4046 2575 4050
rect 2579 4046 2580 4050
rect 2574 4045 2580 4046
rect 2678 4050 2684 4051
rect 2678 4046 2679 4050
rect 2683 4046 2684 4050
rect 2678 4045 2684 4046
rect 3990 4045 3996 4046
rect 2070 4041 2071 4045
rect 2075 4041 2076 4045
rect 2070 4040 2076 4041
rect 3990 4041 3991 4045
rect 3995 4041 3996 4045
rect 3990 4040 3996 4041
rect 110 4028 116 4029
rect 110 4024 111 4028
rect 115 4024 116 4028
rect 110 4023 116 4024
rect 2030 4028 2036 4029
rect 2030 4024 2031 4028
rect 2035 4024 2036 4028
rect 2030 4023 2036 4024
rect 2070 4028 2076 4029
rect 2070 4024 2071 4028
rect 2075 4024 2076 4028
rect 2070 4023 2076 4024
rect 3990 4028 3996 4029
rect 3990 4024 3991 4028
rect 3995 4024 3996 4028
rect 3990 4023 3996 4024
rect 410 4019 416 4020
rect 410 4018 411 4019
rect 377 4016 411 4018
rect 410 4015 411 4016
rect 415 4015 416 4019
rect 518 4019 524 4020
rect 518 4018 519 4019
rect 481 4016 519 4018
rect 410 4014 416 4015
rect 518 4015 519 4016
rect 523 4015 524 4019
rect 622 4019 628 4020
rect 622 4018 623 4019
rect 585 4016 623 4018
rect 518 4014 524 4015
rect 622 4015 623 4016
rect 627 4015 628 4019
rect 726 4019 732 4020
rect 726 4018 727 4019
rect 689 4016 727 4018
rect 622 4014 628 4015
rect 726 4015 727 4016
rect 731 4015 732 4019
rect 830 4019 836 4020
rect 830 4018 831 4019
rect 793 4016 831 4018
rect 726 4014 732 4015
rect 830 4015 831 4016
rect 835 4015 836 4019
rect 934 4019 940 4020
rect 934 4018 935 4019
rect 897 4016 935 4018
rect 830 4014 836 4015
rect 934 4015 935 4016
rect 939 4015 940 4019
rect 1038 4019 1044 4020
rect 1038 4018 1039 4019
rect 1001 4016 1039 4018
rect 934 4014 940 4015
rect 1038 4015 1039 4016
rect 1043 4015 1044 4019
rect 1135 4019 1141 4020
rect 1135 4018 1136 4019
rect 1105 4016 1136 4018
rect 1038 4014 1044 4015
rect 1135 4015 1136 4016
rect 1140 4015 1141 4019
rect 1246 4019 1252 4020
rect 1246 4018 1247 4019
rect 1209 4016 1247 4018
rect 1135 4014 1141 4015
rect 1246 4015 1247 4016
rect 1251 4015 1252 4019
rect 2334 4019 2340 4020
rect 2334 4018 2335 4019
rect 2313 4016 2335 4018
rect 1246 4014 1252 4015
rect 2334 4015 2335 4016
rect 2339 4015 2340 4019
rect 2598 4019 2604 4020
rect 2521 4016 2566 4018
rect 2334 4014 2340 4015
rect 326 4009 332 4010
rect 326 4005 327 4009
rect 331 4005 332 4009
rect 326 4004 332 4005
rect 430 4009 436 4010
rect 430 4005 431 4009
rect 435 4005 436 4009
rect 430 4004 436 4005
rect 534 4009 540 4010
rect 534 4005 535 4009
rect 539 4005 540 4009
rect 534 4004 540 4005
rect 638 4009 644 4010
rect 638 4005 639 4009
rect 643 4005 644 4009
rect 638 4004 644 4005
rect 742 4009 748 4010
rect 742 4005 743 4009
rect 747 4005 748 4009
rect 742 4004 748 4005
rect 846 4009 852 4010
rect 846 4005 847 4009
rect 851 4005 852 4009
rect 846 4004 852 4005
rect 950 4009 956 4010
rect 950 4005 951 4009
rect 955 4005 956 4009
rect 950 4004 956 4005
rect 1054 4009 1060 4010
rect 1054 4005 1055 4009
rect 1059 4005 1060 4009
rect 1054 4004 1060 4005
rect 1158 4009 1164 4010
rect 1158 4005 1159 4009
rect 1163 4005 1164 4009
rect 1158 4004 1164 4005
rect 1262 4009 1268 4010
rect 1262 4005 1263 4009
rect 1267 4005 1268 4009
rect 1262 4004 1268 4005
rect 1366 4009 1372 4010
rect 1366 4005 1367 4009
rect 1371 4005 1372 4009
rect 1366 4004 1372 4005
rect 1470 4009 1476 4010
rect 1470 4005 1471 4009
rect 1475 4005 1476 4009
rect 1470 4004 1476 4005
rect 2262 4009 2268 4010
rect 2262 4005 2263 4009
rect 2267 4005 2268 4009
rect 2262 4004 2268 4005
rect 2366 4009 2372 4010
rect 2366 4005 2367 4009
rect 2371 4005 2372 4009
rect 2366 4004 2372 4005
rect 2470 4009 2476 4010
rect 2470 4005 2471 4009
rect 2475 4005 2476 4009
rect 2470 4004 2476 4005
rect 2564 4002 2566 4016
rect 2598 4015 2599 4019
rect 2603 4015 2604 4019
rect 2598 4014 2604 4015
rect 2574 4009 2580 4010
rect 2574 4005 2575 4009
rect 2579 4005 2580 4009
rect 2678 4009 2684 4010
rect 2574 4004 2580 4005
rect 2640 4004 2674 4006
rect 2678 4005 2679 4009
rect 2683 4005 2684 4009
rect 2678 4004 2684 4005
rect 2640 4002 2642 4004
rect 2564 4000 2642 4002
rect 295 3999 301 4000
rect 295 3995 296 3999
rect 300 3998 301 3999
rect 399 3999 405 4000
rect 399 3998 400 3999
rect 300 3996 400 3998
rect 300 3995 301 3996
rect 295 3994 301 3995
rect 399 3995 400 3996
rect 404 3995 405 3999
rect 399 3994 405 3995
rect 410 3999 416 4000
rect 410 3995 411 3999
rect 415 3998 416 3999
rect 503 3999 509 4000
rect 503 3998 504 3999
rect 415 3996 504 3998
rect 415 3995 416 3996
rect 410 3994 416 3995
rect 503 3995 504 3996
rect 508 3995 509 3999
rect 503 3994 509 3995
rect 518 3999 524 4000
rect 518 3995 519 3999
rect 523 3998 524 3999
rect 607 3999 613 4000
rect 607 3998 608 3999
rect 523 3996 608 3998
rect 523 3995 524 3996
rect 518 3994 524 3995
rect 607 3995 608 3996
rect 612 3995 613 3999
rect 607 3994 613 3995
rect 622 3999 628 4000
rect 622 3995 623 3999
rect 627 3998 628 3999
rect 711 3999 717 4000
rect 711 3998 712 3999
rect 627 3996 712 3998
rect 627 3995 628 3996
rect 622 3994 628 3995
rect 711 3995 712 3996
rect 716 3995 717 3999
rect 711 3994 717 3995
rect 726 3999 732 4000
rect 726 3995 727 3999
rect 731 3998 732 3999
rect 815 3999 821 4000
rect 815 3998 816 3999
rect 731 3996 816 3998
rect 731 3995 732 3996
rect 726 3994 732 3995
rect 815 3995 816 3996
rect 820 3995 821 3999
rect 815 3994 821 3995
rect 830 3999 836 4000
rect 830 3995 831 3999
rect 835 3998 836 3999
rect 919 3999 925 4000
rect 919 3998 920 3999
rect 835 3996 920 3998
rect 835 3995 836 3996
rect 830 3994 836 3995
rect 919 3995 920 3996
rect 924 3995 925 3999
rect 919 3994 925 3995
rect 934 3999 940 4000
rect 934 3995 935 3999
rect 939 3998 940 3999
rect 1023 3999 1029 4000
rect 1023 3998 1024 3999
rect 939 3996 1024 3998
rect 939 3995 940 3996
rect 934 3994 940 3995
rect 1023 3995 1024 3996
rect 1028 3995 1029 3999
rect 1023 3994 1029 3995
rect 1038 3999 1044 4000
rect 1038 3995 1039 3999
rect 1043 3998 1044 3999
rect 1127 3999 1133 4000
rect 1127 3998 1128 3999
rect 1043 3996 1128 3998
rect 1043 3995 1044 3996
rect 1038 3994 1044 3995
rect 1127 3995 1128 3996
rect 1132 3995 1133 3999
rect 1127 3994 1133 3995
rect 1135 3999 1141 4000
rect 1135 3995 1136 3999
rect 1140 3998 1141 3999
rect 1231 3999 1237 4000
rect 1231 3998 1232 3999
rect 1140 3996 1232 3998
rect 1140 3995 1141 3996
rect 1135 3994 1141 3995
rect 1231 3995 1232 3996
rect 1236 3995 1237 3999
rect 1231 3994 1237 3995
rect 1247 3999 1253 4000
rect 1247 3995 1248 3999
rect 1252 3995 1253 3999
rect 1247 3994 1253 3995
rect 1335 3999 1341 4000
rect 1335 3995 1336 3999
rect 1340 3998 1341 3999
rect 1351 3999 1357 4000
rect 1351 3998 1352 3999
rect 1340 3996 1352 3998
rect 1340 3995 1341 3996
rect 1335 3994 1341 3995
rect 1351 3995 1352 3996
rect 1356 3995 1357 3999
rect 1351 3994 1357 3995
rect 1439 3999 1445 4000
rect 1439 3995 1440 3999
rect 1444 3998 1445 3999
rect 1455 3999 1461 4000
rect 1455 3998 1456 3999
rect 1444 3996 1456 3998
rect 1444 3995 1445 3996
rect 1439 3994 1445 3995
rect 1455 3995 1456 3996
rect 1460 3995 1461 3999
rect 1543 3999 1549 4000
rect 1543 3998 1544 3999
rect 1455 3994 1461 3995
rect 1464 3996 1544 3998
rect 247 3983 253 3984
rect 247 3979 248 3983
rect 252 3982 253 3983
rect 367 3983 373 3984
rect 367 3982 368 3983
rect 252 3980 368 3982
rect 252 3979 253 3980
rect 247 3978 253 3979
rect 367 3979 368 3980
rect 372 3979 373 3983
rect 367 3978 373 3979
rect 455 3983 461 3984
rect 455 3979 456 3983
rect 460 3982 461 3983
rect 575 3983 581 3984
rect 575 3982 576 3983
rect 460 3980 576 3982
rect 460 3979 461 3980
rect 455 3978 461 3979
rect 575 3979 576 3980
rect 580 3979 581 3983
rect 575 3978 581 3979
rect 663 3983 669 3984
rect 663 3979 664 3983
rect 668 3982 669 3983
rect 775 3983 781 3984
rect 775 3982 776 3983
rect 668 3980 776 3982
rect 668 3979 669 3980
rect 663 3978 669 3979
rect 775 3979 776 3980
rect 780 3979 781 3983
rect 775 3978 781 3979
rect 862 3983 869 3984
rect 862 3979 863 3983
rect 868 3979 869 3983
rect 862 3978 869 3979
rect 1055 3983 1061 3984
rect 1055 3979 1056 3983
rect 1060 3982 1061 3983
rect 1151 3983 1157 3984
rect 1151 3982 1152 3983
rect 1060 3980 1152 3982
rect 1060 3979 1061 3980
rect 1055 3978 1061 3979
rect 1151 3979 1152 3980
rect 1156 3979 1157 3983
rect 1151 3978 1157 3979
rect 1239 3983 1245 3984
rect 1239 3979 1240 3983
rect 1244 3982 1245 3983
rect 1248 3982 1250 3994
rect 1254 3991 1260 3992
rect 1254 3987 1255 3991
rect 1259 3990 1260 3991
rect 1464 3990 1466 3996
rect 1543 3995 1544 3996
rect 1548 3995 1549 3999
rect 1543 3994 1549 3995
rect 2335 3999 2341 4000
rect 2335 3995 2336 3999
rect 2340 3998 2341 3999
rect 2351 3999 2357 4000
rect 2351 3998 2352 3999
rect 2340 3996 2352 3998
rect 2340 3995 2341 3996
rect 2335 3994 2341 3995
rect 2351 3995 2352 3996
rect 2356 3995 2357 3999
rect 2351 3994 2357 3995
rect 2414 3999 2420 4000
rect 2414 3995 2415 3999
rect 2419 3998 2420 3999
rect 2439 3999 2445 4000
rect 2439 3998 2440 3999
rect 2419 3996 2440 3998
rect 2419 3995 2420 3996
rect 2414 3994 2420 3995
rect 2439 3995 2440 3996
rect 2444 3995 2445 3999
rect 2543 3999 2549 4000
rect 2543 3998 2544 3999
rect 2439 3994 2445 3995
rect 2448 3996 2544 3998
rect 1259 3988 1466 3990
rect 2334 3991 2340 3992
rect 1259 3987 1260 3988
rect 1254 3986 1260 3987
rect 2294 3987 2300 3988
rect 1244 3980 1250 3982
rect 1286 3983 1292 3984
rect 1244 3979 1245 3980
rect 1239 3978 1245 3979
rect 1286 3979 1287 3983
rect 1291 3982 1292 3983
rect 1415 3983 1421 3984
rect 1415 3982 1416 3983
rect 1291 3980 1416 3982
rect 1291 3979 1292 3980
rect 1286 3978 1292 3979
rect 1415 3979 1416 3980
rect 1420 3979 1421 3983
rect 1415 3978 1421 3979
rect 1591 3983 1597 3984
rect 1591 3979 1592 3983
rect 1596 3982 1597 3983
rect 1687 3983 1693 3984
rect 1687 3982 1688 3983
rect 1596 3980 1688 3982
rect 1596 3979 1597 3980
rect 1591 3978 1597 3979
rect 1687 3979 1688 3980
rect 1692 3979 1693 3983
rect 1687 3978 1693 3979
rect 1774 3983 1781 3984
rect 1774 3979 1775 3983
rect 1780 3979 1781 3983
rect 2294 3983 2295 3987
rect 2299 3986 2300 3987
rect 2303 3987 2309 3988
rect 2303 3986 2304 3987
rect 2299 3984 2304 3986
rect 2299 3983 2300 3984
rect 2294 3982 2300 3983
rect 2303 3983 2304 3984
rect 2308 3983 2309 3987
rect 2334 3987 2335 3991
rect 2339 3990 2340 3991
rect 2448 3990 2450 3996
rect 2543 3995 2544 3996
rect 2548 3995 2549 3999
rect 2543 3994 2549 3995
rect 2647 3999 2653 4000
rect 2647 3995 2648 3999
rect 2652 3998 2653 3999
rect 2663 3999 2669 4000
rect 2663 3998 2664 3999
rect 2652 3996 2664 3998
rect 2652 3995 2653 3996
rect 2647 3994 2653 3995
rect 2663 3995 2664 3996
rect 2668 3995 2669 3999
rect 2672 3998 2674 4004
rect 2751 3999 2757 4000
rect 2751 3998 2752 3999
rect 2672 3996 2752 3998
rect 2663 3994 2669 3995
rect 2751 3995 2752 3996
rect 2756 3995 2757 3999
rect 2751 3994 2757 3995
rect 2339 3988 2450 3990
rect 2339 3987 2340 3988
rect 2334 3986 2340 3987
rect 2463 3987 2469 3988
rect 2463 3986 2464 3987
rect 2303 3982 2309 3983
rect 2344 3984 2464 3986
rect 1774 3978 1781 3979
rect 2230 3979 2236 3980
rect 174 3975 180 3976
rect 174 3971 175 3975
rect 179 3971 180 3975
rect 174 3970 180 3971
rect 382 3975 388 3976
rect 382 3971 383 3975
rect 387 3971 388 3975
rect 382 3970 388 3971
rect 590 3975 596 3976
rect 590 3971 591 3975
rect 595 3971 596 3975
rect 590 3970 596 3971
rect 790 3975 796 3976
rect 790 3971 791 3975
rect 795 3971 796 3975
rect 790 3970 796 3971
rect 982 3975 988 3976
rect 982 3971 983 3975
rect 987 3971 988 3975
rect 982 3970 988 3971
rect 1166 3975 1172 3976
rect 1166 3971 1167 3975
rect 1171 3971 1172 3975
rect 1166 3970 1172 3971
rect 1342 3975 1348 3976
rect 1342 3971 1343 3975
rect 1347 3971 1348 3975
rect 1342 3970 1348 3971
rect 1518 3975 1524 3976
rect 1518 3971 1519 3975
rect 1523 3971 1524 3975
rect 1518 3970 1524 3971
rect 1702 3975 1708 3976
rect 1702 3971 1703 3975
rect 1707 3971 1708 3975
rect 2230 3975 2231 3979
rect 2235 3975 2236 3979
rect 2230 3974 2236 3975
rect 1702 3970 1708 3971
rect 2344 3970 2346 3984
rect 2463 3983 2464 3984
rect 2468 3983 2469 3987
rect 2463 3982 2469 3983
rect 2598 3987 2604 3988
rect 2598 3983 2599 3987
rect 2603 3986 2604 3987
rect 2623 3987 2629 3988
rect 2623 3986 2624 3987
rect 2603 3984 2624 3986
rect 2603 3983 2604 3984
rect 2598 3982 2604 3983
rect 2623 3983 2624 3984
rect 2628 3983 2629 3987
rect 2775 3987 2781 3988
rect 2775 3986 2776 3987
rect 2623 3982 2629 3983
rect 2660 3984 2776 3986
rect 2390 3979 2396 3980
rect 2390 3975 2391 3979
rect 2395 3975 2396 3979
rect 2390 3974 2396 3975
rect 2550 3979 2556 3980
rect 2550 3975 2551 3979
rect 2555 3975 2556 3979
rect 2550 3974 2556 3975
rect 2660 3970 2662 3984
rect 2775 3983 2776 3984
rect 2780 3983 2781 3987
rect 2775 3982 2781 3983
rect 2919 3987 2925 3988
rect 2919 3983 2920 3987
rect 2924 3986 2925 3987
rect 2967 3987 2973 3988
rect 2967 3986 2968 3987
rect 2924 3984 2968 3986
rect 2924 3983 2925 3984
rect 2919 3982 2925 3983
rect 2967 3983 2968 3984
rect 2972 3983 2973 3987
rect 2967 3982 2973 3983
rect 3055 3987 3061 3988
rect 3055 3983 3056 3987
rect 3060 3986 3061 3987
rect 3103 3987 3109 3988
rect 3103 3986 3104 3987
rect 3060 3984 3104 3986
rect 3060 3983 3061 3984
rect 3055 3982 3061 3983
rect 3103 3983 3104 3984
rect 3108 3983 3109 3987
rect 3103 3982 3109 3983
rect 3191 3987 3197 3988
rect 3191 3983 3192 3987
rect 3196 3986 3197 3987
rect 3231 3987 3237 3988
rect 3231 3986 3232 3987
rect 3196 3984 3232 3986
rect 3196 3983 3197 3984
rect 3191 3982 3197 3983
rect 3231 3983 3232 3984
rect 3236 3983 3237 3987
rect 3231 3982 3237 3983
rect 3319 3987 3325 3988
rect 3319 3983 3320 3987
rect 3324 3986 3325 3987
rect 3351 3987 3357 3988
rect 3351 3986 3352 3987
rect 3324 3984 3352 3986
rect 3324 3983 3325 3984
rect 3319 3982 3325 3983
rect 3351 3983 3352 3984
rect 3356 3983 3357 3987
rect 3351 3982 3357 3983
rect 3439 3987 3445 3988
rect 3439 3983 3440 3987
rect 3444 3986 3445 3987
rect 3463 3987 3469 3988
rect 3463 3986 3464 3987
rect 3444 3984 3464 3986
rect 3444 3983 3445 3984
rect 3439 3982 3445 3983
rect 3463 3983 3464 3984
rect 3468 3983 3469 3987
rect 3463 3982 3469 3983
rect 3551 3987 3557 3988
rect 3551 3983 3552 3987
rect 3556 3986 3557 3987
rect 3583 3987 3589 3988
rect 3583 3986 3584 3987
rect 3556 3984 3584 3986
rect 3556 3983 3557 3984
rect 3551 3982 3557 3983
rect 3583 3983 3584 3984
rect 3588 3983 3589 3987
rect 3583 3982 3589 3983
rect 3671 3987 3677 3988
rect 3671 3983 3672 3987
rect 3676 3986 3677 3987
rect 3703 3987 3709 3988
rect 3703 3986 3704 3987
rect 3676 3984 3704 3986
rect 3676 3983 3677 3984
rect 3671 3982 3677 3983
rect 3703 3983 3704 3984
rect 3708 3983 3709 3987
rect 3703 3982 3709 3983
rect 3791 3987 3797 3988
rect 3791 3983 3792 3987
rect 3796 3986 3797 3987
rect 3823 3987 3829 3988
rect 3823 3986 3824 3987
rect 3796 3984 3824 3986
rect 3796 3983 3797 3984
rect 3791 3982 3797 3983
rect 3823 3983 3824 3984
rect 3828 3983 3829 3987
rect 3823 3982 3829 3983
rect 3882 3987 3888 3988
rect 3882 3983 3883 3987
rect 3887 3986 3888 3987
rect 3911 3987 3917 3988
rect 3911 3986 3912 3987
rect 3887 3984 3912 3986
rect 3887 3983 3888 3984
rect 3882 3982 3888 3983
rect 3911 3983 3912 3984
rect 3916 3983 3917 3987
rect 3911 3982 3917 3983
rect 2702 3979 2708 3980
rect 2702 3975 2703 3979
rect 2707 3975 2708 3979
rect 2702 3974 2708 3975
rect 2846 3979 2852 3980
rect 2846 3975 2847 3979
rect 2851 3975 2852 3979
rect 2846 3974 2852 3975
rect 2982 3979 2988 3980
rect 2982 3975 2983 3979
rect 2987 3975 2988 3979
rect 2982 3974 2988 3975
rect 3118 3979 3124 3980
rect 3118 3975 3119 3979
rect 3123 3975 3124 3979
rect 3118 3974 3124 3975
rect 3246 3979 3252 3980
rect 3246 3975 3247 3979
rect 3251 3975 3252 3979
rect 3246 3974 3252 3975
rect 3366 3979 3372 3980
rect 3366 3975 3367 3979
rect 3371 3975 3372 3979
rect 3366 3974 3372 3975
rect 3478 3979 3484 3980
rect 3478 3975 3479 3979
rect 3483 3975 3484 3979
rect 3478 3974 3484 3975
rect 3598 3979 3604 3980
rect 3598 3975 3599 3979
rect 3603 3975 3604 3979
rect 3598 3974 3604 3975
rect 3718 3979 3724 3980
rect 3718 3975 3719 3979
rect 3723 3975 3724 3979
rect 3718 3974 3724 3975
rect 3838 3979 3844 3980
rect 3838 3975 3839 3979
rect 3843 3975 3844 3979
rect 3838 3974 3844 3975
rect 2950 3971 2956 3972
rect 2950 3970 2951 3971
rect 2281 3968 2346 3970
rect 2601 3968 2662 3970
rect 2897 3968 2951 3970
rect 295 3967 301 3968
rect 295 3966 296 3967
rect 225 3964 296 3966
rect 295 3963 296 3964
rect 300 3963 301 3967
rect 1074 3967 1080 3968
rect 1074 3966 1075 3967
rect 1033 3964 1075 3966
rect 295 3962 301 3963
rect 1074 3963 1075 3964
rect 1079 3963 1080 3967
rect 1502 3967 1508 3968
rect 1502 3966 1503 3967
rect 1393 3964 1503 3966
rect 1074 3962 1080 3963
rect 1502 3963 1503 3964
rect 1507 3963 1508 3967
rect 2414 3967 2420 3968
rect 1502 3962 1508 3963
rect 1510 3963 1516 3964
rect 1510 3959 1511 3963
rect 1515 3959 1516 3963
rect 2414 3963 2415 3967
rect 2419 3963 2420 3967
rect 2414 3962 2420 3963
rect 2726 3967 2732 3968
rect 2726 3963 2727 3967
rect 2731 3963 2732 3967
rect 2950 3967 2951 3968
rect 2955 3967 2956 3971
rect 2950 3966 2956 3967
rect 2726 3962 2732 3963
rect 1510 3958 1516 3959
rect 2070 3960 2076 3961
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 110 3951 116 3952
rect 2030 3956 2036 3957
rect 2030 3952 2031 3956
rect 2035 3952 2036 3956
rect 2070 3956 2071 3960
rect 2075 3956 2076 3960
rect 2070 3955 2076 3956
rect 3990 3960 3996 3961
rect 3990 3956 3991 3960
rect 3995 3956 3996 3960
rect 3990 3955 3996 3956
rect 2030 3951 2036 3952
rect 2070 3943 2076 3944
rect 110 3939 116 3940
rect 110 3935 111 3939
rect 115 3935 116 3939
rect 2030 3939 2036 3940
rect 2030 3935 2031 3939
rect 2035 3935 2036 3939
rect 2070 3939 2071 3943
rect 2075 3939 2076 3943
rect 3990 3943 3996 3944
rect 3990 3939 3991 3943
rect 3995 3939 3996 3943
rect 2070 3938 2076 3939
rect 2230 3938 2236 3939
rect 110 3934 116 3935
rect 174 3934 180 3935
rect 174 3930 175 3934
rect 179 3930 180 3934
rect 174 3929 180 3930
rect 382 3934 388 3935
rect 382 3930 383 3934
rect 387 3930 388 3934
rect 382 3929 388 3930
rect 590 3934 596 3935
rect 590 3930 591 3934
rect 595 3930 596 3934
rect 590 3929 596 3930
rect 790 3934 796 3935
rect 790 3930 791 3934
rect 795 3930 796 3934
rect 790 3929 796 3930
rect 982 3934 988 3935
rect 982 3930 983 3934
rect 987 3930 988 3934
rect 982 3929 988 3930
rect 1166 3934 1172 3935
rect 1166 3930 1167 3934
rect 1171 3930 1172 3934
rect 1166 3929 1172 3930
rect 1342 3934 1348 3935
rect 1342 3930 1343 3934
rect 1347 3930 1348 3934
rect 1342 3929 1348 3930
rect 1518 3934 1524 3935
rect 1518 3930 1519 3934
rect 1523 3930 1524 3934
rect 1518 3929 1524 3930
rect 1702 3934 1708 3935
rect 2030 3934 2036 3935
rect 2230 3934 2231 3938
rect 2235 3934 2236 3938
rect 1702 3930 1703 3934
rect 1707 3930 1708 3934
rect 2230 3933 2236 3934
rect 2390 3938 2396 3939
rect 2390 3934 2391 3938
rect 2395 3934 2396 3938
rect 2390 3933 2396 3934
rect 2550 3938 2556 3939
rect 2550 3934 2551 3938
rect 2555 3934 2556 3938
rect 2550 3933 2556 3934
rect 2702 3938 2708 3939
rect 2702 3934 2703 3938
rect 2707 3934 2708 3938
rect 2702 3933 2708 3934
rect 2846 3938 2852 3939
rect 2846 3934 2847 3938
rect 2851 3934 2852 3938
rect 2846 3933 2852 3934
rect 2982 3938 2988 3939
rect 2982 3934 2983 3938
rect 2987 3934 2988 3938
rect 2982 3933 2988 3934
rect 3118 3938 3124 3939
rect 3118 3934 3119 3938
rect 3123 3934 3124 3938
rect 3118 3933 3124 3934
rect 3246 3938 3252 3939
rect 3246 3934 3247 3938
rect 3251 3934 3252 3938
rect 3246 3933 3252 3934
rect 3366 3938 3372 3939
rect 3366 3934 3367 3938
rect 3371 3934 3372 3938
rect 3366 3933 3372 3934
rect 3478 3938 3484 3939
rect 3478 3934 3479 3938
rect 3483 3934 3484 3938
rect 3478 3933 3484 3934
rect 3598 3938 3604 3939
rect 3598 3934 3599 3938
rect 3603 3934 3604 3938
rect 3598 3933 3604 3934
rect 3718 3938 3724 3939
rect 3718 3934 3719 3938
rect 3723 3934 3724 3938
rect 3718 3933 3724 3934
rect 3838 3938 3844 3939
rect 3990 3938 3996 3939
rect 3838 3934 3839 3938
rect 3843 3934 3844 3938
rect 3838 3933 3844 3934
rect 1702 3929 1708 3930
rect 2222 3906 2228 3907
rect 358 3902 364 3903
rect 358 3898 359 3902
rect 363 3898 364 3902
rect 110 3897 116 3898
rect 358 3897 364 3898
rect 550 3902 556 3903
rect 550 3898 551 3902
rect 555 3898 556 3902
rect 550 3897 556 3898
rect 734 3902 740 3903
rect 734 3898 735 3902
rect 739 3898 740 3902
rect 734 3897 740 3898
rect 918 3902 924 3903
rect 918 3898 919 3902
rect 923 3898 924 3902
rect 918 3897 924 3898
rect 1086 3902 1092 3903
rect 1086 3898 1087 3902
rect 1091 3898 1092 3902
rect 1086 3897 1092 3898
rect 1246 3902 1252 3903
rect 1246 3898 1247 3902
rect 1251 3898 1252 3902
rect 1246 3897 1252 3898
rect 1398 3902 1404 3903
rect 1398 3898 1399 3902
rect 1403 3898 1404 3902
rect 1398 3897 1404 3898
rect 1542 3902 1548 3903
rect 1542 3898 1543 3902
rect 1547 3898 1548 3902
rect 1542 3897 1548 3898
rect 1678 3902 1684 3903
rect 1678 3898 1679 3902
rect 1683 3898 1684 3902
rect 1678 3897 1684 3898
rect 1814 3902 1820 3903
rect 1814 3898 1815 3902
rect 1819 3898 1820 3902
rect 1814 3897 1820 3898
rect 1934 3902 1940 3903
rect 2222 3902 2223 3906
rect 2227 3902 2228 3906
rect 1934 3898 1935 3902
rect 1939 3898 1940 3902
rect 2070 3901 2076 3902
rect 2222 3901 2228 3902
rect 2454 3906 2460 3907
rect 2454 3902 2455 3906
rect 2459 3902 2460 3906
rect 2454 3901 2460 3902
rect 2670 3906 2676 3907
rect 2670 3902 2671 3906
rect 2675 3902 2676 3906
rect 2670 3901 2676 3902
rect 2878 3906 2884 3907
rect 2878 3902 2879 3906
rect 2883 3902 2884 3906
rect 2878 3901 2884 3902
rect 3070 3906 3076 3907
rect 3070 3902 3071 3906
rect 3075 3902 3076 3906
rect 3070 3901 3076 3902
rect 3246 3906 3252 3907
rect 3246 3902 3247 3906
rect 3251 3902 3252 3906
rect 3246 3901 3252 3902
rect 3414 3906 3420 3907
rect 3414 3902 3415 3906
rect 3419 3902 3420 3906
rect 3414 3901 3420 3902
rect 3582 3906 3588 3907
rect 3582 3902 3583 3906
rect 3587 3902 3588 3906
rect 3582 3901 3588 3902
rect 3750 3906 3756 3907
rect 3750 3902 3751 3906
rect 3755 3902 3756 3906
rect 3750 3901 3756 3902
rect 3990 3901 3996 3902
rect 1934 3897 1940 3898
rect 2030 3897 2036 3898
rect 110 3893 111 3897
rect 115 3893 116 3897
rect 110 3892 116 3893
rect 2030 3893 2031 3897
rect 2035 3893 2036 3897
rect 2070 3897 2071 3901
rect 2075 3897 2076 3901
rect 2070 3896 2076 3897
rect 3990 3897 3991 3901
rect 3995 3897 3996 3901
rect 3990 3896 3996 3897
rect 2030 3892 2036 3893
rect 2070 3884 2076 3885
rect 110 3880 116 3881
rect 110 3876 111 3880
rect 115 3876 116 3880
rect 110 3875 116 3876
rect 2030 3880 2036 3881
rect 2030 3876 2031 3880
rect 2035 3876 2036 3880
rect 2070 3880 2071 3884
rect 2075 3880 2076 3884
rect 2070 3879 2076 3880
rect 3990 3884 3996 3885
rect 3990 3880 3991 3884
rect 3995 3880 3996 3884
rect 3990 3879 3996 3880
rect 2030 3875 2036 3876
rect 2294 3875 2300 3876
rect 2294 3874 2295 3875
rect 2273 3872 2295 3874
rect 534 3871 540 3872
rect 534 3870 535 3871
rect 409 3868 535 3870
rect 534 3867 535 3868
rect 539 3867 540 3871
rect 1662 3871 1668 3872
rect 1662 3870 1663 3871
rect 1137 3868 1161 3870
rect 1593 3868 1663 3870
rect 534 3866 540 3867
rect 358 3861 364 3862
rect 358 3857 359 3861
rect 363 3857 364 3861
rect 358 3856 364 3857
rect 550 3861 556 3862
rect 550 3857 551 3861
rect 555 3857 556 3861
rect 734 3861 740 3862
rect 550 3856 556 3857
rect 718 3859 724 3860
rect 718 3855 719 3859
rect 723 3858 724 3859
rect 723 3856 730 3858
rect 734 3857 735 3861
rect 739 3857 740 3861
rect 918 3861 924 3862
rect 734 3856 740 3857
rect 796 3856 914 3858
rect 918 3857 919 3861
rect 923 3857 924 3861
rect 918 3856 924 3857
rect 1086 3861 1092 3862
rect 1086 3857 1087 3861
rect 1091 3857 1092 3861
rect 1086 3856 1092 3857
rect 1159 3858 1161 3868
rect 1662 3867 1663 3868
rect 1667 3867 1668 3871
rect 1798 3871 1804 3872
rect 1798 3870 1799 3871
rect 1729 3868 1799 3870
rect 1662 3866 1668 3867
rect 1798 3867 1799 3868
rect 1803 3867 1804 3871
rect 1902 3871 1908 3872
rect 1902 3870 1903 3871
rect 1865 3868 1903 3870
rect 1798 3866 1804 3867
rect 1902 3867 1903 3868
rect 1907 3867 1908 3871
rect 2006 3871 2012 3872
rect 2006 3870 2007 3871
rect 1985 3868 2007 3870
rect 1902 3866 1908 3867
rect 2006 3867 2007 3868
rect 2011 3867 2012 3871
rect 2294 3871 2295 3872
rect 2299 3871 2300 3875
rect 2526 3875 2532 3876
rect 2526 3874 2527 3875
rect 2505 3872 2527 3874
rect 2294 3870 2300 3871
rect 2526 3871 2527 3872
rect 2531 3871 2532 3875
rect 3054 3875 3060 3876
rect 3054 3874 3055 3875
rect 2929 3872 3055 3874
rect 2526 3870 2532 3871
rect 3054 3871 3055 3872
rect 3059 3871 3060 3875
rect 3734 3875 3740 3876
rect 3734 3874 3735 3875
rect 3633 3872 3735 3874
rect 3054 3870 3060 3871
rect 3734 3871 3735 3872
rect 3739 3871 3740 3875
rect 3882 3875 3888 3876
rect 3882 3874 3883 3875
rect 3801 3872 3883 3874
rect 3734 3870 3740 3871
rect 3882 3871 3883 3872
rect 3887 3871 3888 3875
rect 3882 3870 3888 3871
rect 2006 3866 2012 3867
rect 2222 3865 2228 3866
rect 1246 3861 1252 3862
rect 1159 3856 1242 3858
rect 1246 3857 1247 3861
rect 1251 3857 1252 3861
rect 1398 3861 1404 3862
rect 1246 3856 1252 3857
rect 1312 3856 1394 3858
rect 1398 3857 1399 3861
rect 1403 3857 1404 3861
rect 1542 3861 1548 3862
rect 1398 3856 1404 3857
rect 1464 3856 1522 3858
rect 1542 3857 1543 3861
rect 1547 3857 1548 3861
rect 1542 3856 1548 3857
rect 1678 3861 1684 3862
rect 1678 3857 1679 3861
rect 1683 3857 1684 3861
rect 1678 3856 1684 3857
rect 1814 3861 1820 3862
rect 1814 3857 1815 3861
rect 1819 3857 1820 3861
rect 1814 3856 1820 3857
rect 1934 3861 1940 3862
rect 1934 3857 1935 3861
rect 1939 3857 1940 3861
rect 2222 3861 2223 3865
rect 2227 3861 2228 3865
rect 2222 3860 2228 3861
rect 2454 3865 2460 3866
rect 2454 3861 2455 3865
rect 2459 3861 2460 3865
rect 2454 3860 2460 3861
rect 2670 3865 2676 3866
rect 2670 3861 2671 3865
rect 2675 3861 2676 3865
rect 2670 3860 2676 3861
rect 2878 3865 2884 3866
rect 2878 3861 2879 3865
rect 2883 3861 2884 3865
rect 2878 3860 2884 3861
rect 3070 3865 3076 3866
rect 3070 3861 3071 3865
rect 3075 3861 3076 3865
rect 3070 3860 3076 3861
rect 3246 3865 3252 3866
rect 3246 3861 3247 3865
rect 3251 3861 3252 3865
rect 3246 3860 3252 3861
rect 3414 3865 3420 3866
rect 3414 3861 3415 3865
rect 3419 3861 3420 3865
rect 3414 3860 3420 3861
rect 3582 3865 3588 3866
rect 3582 3861 3583 3865
rect 3587 3861 3588 3865
rect 3582 3860 3588 3861
rect 3750 3865 3756 3866
rect 3750 3861 3751 3865
rect 3755 3861 3756 3865
rect 3750 3860 3756 3861
rect 1934 3856 1940 3857
rect 723 3855 724 3856
rect 718 3854 724 3855
rect 728 3854 730 3856
rect 796 3854 798 3856
rect 728 3852 798 3854
rect 431 3851 437 3852
rect 431 3847 432 3851
rect 436 3850 437 3851
rect 535 3851 541 3852
rect 535 3850 536 3851
rect 436 3848 536 3850
rect 436 3847 437 3848
rect 431 3846 437 3847
rect 535 3847 536 3848
rect 540 3847 541 3851
rect 535 3846 541 3847
rect 623 3851 629 3852
rect 623 3847 624 3851
rect 628 3850 629 3851
rect 719 3851 725 3852
rect 719 3850 720 3851
rect 628 3848 720 3850
rect 628 3847 629 3848
rect 623 3846 629 3847
rect 719 3847 720 3848
rect 724 3847 725 3851
rect 719 3846 725 3847
rect 807 3851 813 3852
rect 807 3847 808 3851
rect 812 3850 813 3851
rect 903 3851 909 3852
rect 903 3850 904 3851
rect 812 3848 904 3850
rect 812 3847 813 3848
rect 807 3846 813 3847
rect 903 3847 904 3848
rect 908 3847 909 3851
rect 912 3850 914 3856
rect 1240 3854 1242 3856
rect 1312 3854 1314 3856
rect 1240 3852 1314 3854
rect 1392 3854 1394 3856
rect 1464 3854 1466 3856
rect 1392 3852 1466 3854
rect 991 3851 997 3852
rect 991 3850 992 3851
rect 912 3848 992 3850
rect 903 3846 909 3847
rect 991 3847 992 3848
rect 996 3847 997 3851
rect 991 3846 997 3847
rect 1159 3851 1165 3852
rect 1159 3847 1160 3851
rect 1164 3850 1165 3851
rect 1231 3851 1237 3852
rect 1231 3850 1232 3851
rect 1164 3848 1232 3850
rect 1164 3847 1165 3848
rect 1159 3846 1165 3847
rect 1231 3847 1232 3848
rect 1236 3847 1237 3851
rect 1231 3846 1237 3847
rect 1319 3851 1325 3852
rect 1319 3847 1320 3851
rect 1324 3850 1325 3851
rect 1383 3851 1389 3852
rect 1383 3850 1384 3851
rect 1324 3848 1384 3850
rect 1324 3847 1325 3848
rect 1319 3846 1325 3847
rect 1383 3847 1384 3848
rect 1388 3847 1389 3851
rect 1383 3846 1389 3847
rect 1471 3851 1477 3852
rect 1471 3847 1472 3851
rect 1476 3850 1477 3851
rect 1510 3851 1516 3852
rect 1510 3850 1511 3851
rect 1476 3848 1511 3850
rect 1476 3847 1477 3848
rect 1471 3846 1477 3847
rect 1510 3847 1511 3848
rect 1515 3847 1516 3851
rect 1520 3850 1522 3856
rect 2254 3855 2260 3856
rect 1615 3851 1621 3852
rect 1615 3850 1616 3851
rect 1520 3848 1616 3850
rect 1510 3846 1516 3847
rect 1615 3847 1616 3848
rect 1620 3847 1621 3851
rect 1615 3846 1621 3847
rect 1662 3851 1668 3852
rect 1662 3847 1663 3851
rect 1667 3850 1668 3851
rect 1751 3851 1757 3852
rect 1751 3850 1752 3851
rect 1667 3848 1752 3850
rect 1667 3847 1668 3848
rect 1662 3846 1668 3847
rect 1751 3847 1752 3848
rect 1756 3847 1757 3851
rect 1751 3846 1757 3847
rect 1798 3851 1804 3852
rect 1798 3847 1799 3851
rect 1803 3850 1804 3851
rect 1887 3851 1893 3852
rect 1887 3850 1888 3851
rect 1803 3848 1888 3850
rect 1803 3847 1804 3848
rect 1798 3846 1804 3847
rect 1887 3847 1888 3848
rect 1892 3847 1893 3851
rect 1887 3846 1893 3847
rect 1902 3851 1908 3852
rect 1902 3847 1903 3851
rect 1907 3850 1908 3851
rect 2007 3851 2013 3852
rect 2007 3850 2008 3851
rect 1907 3848 2008 3850
rect 1907 3847 1908 3848
rect 1902 3846 1908 3847
rect 2007 3847 2008 3848
rect 2012 3847 2013 3851
rect 2254 3851 2255 3855
rect 2259 3854 2260 3855
rect 2295 3855 2301 3856
rect 2295 3854 2296 3855
rect 2259 3852 2296 3854
rect 2259 3851 2260 3852
rect 2254 3850 2260 3851
rect 2295 3851 2296 3852
rect 2300 3851 2301 3855
rect 2295 3850 2301 3851
rect 2527 3855 2533 3856
rect 2527 3851 2528 3855
rect 2532 3854 2533 3855
rect 2655 3855 2661 3856
rect 2655 3854 2656 3855
rect 2532 3852 2656 3854
rect 2532 3851 2533 3852
rect 2527 3850 2533 3851
rect 2655 3851 2656 3852
rect 2660 3851 2661 3855
rect 2655 3850 2661 3851
rect 2726 3855 2732 3856
rect 2726 3851 2727 3855
rect 2731 3854 2732 3855
rect 2743 3855 2749 3856
rect 2743 3854 2744 3855
rect 2731 3852 2744 3854
rect 2731 3851 2732 3852
rect 2726 3850 2732 3851
rect 2743 3851 2744 3852
rect 2748 3851 2749 3855
rect 2743 3850 2749 3851
rect 2950 3855 2957 3856
rect 2950 3851 2951 3855
rect 2956 3851 2957 3855
rect 2950 3850 2957 3851
rect 3055 3855 3061 3856
rect 3055 3851 3056 3855
rect 3060 3854 3061 3855
rect 3143 3855 3149 3856
rect 3060 3852 3070 3854
rect 3060 3851 3061 3852
rect 3055 3850 3061 3851
rect 3068 3850 3070 3852
rect 3143 3851 3144 3855
rect 3148 3854 3149 3855
rect 3231 3855 3237 3856
rect 3231 3854 3232 3855
rect 3148 3852 3232 3854
rect 3148 3851 3149 3852
rect 3143 3850 3149 3851
rect 3231 3851 3232 3852
rect 3236 3851 3237 3855
rect 3231 3850 3237 3851
rect 3319 3855 3325 3856
rect 3319 3851 3320 3855
rect 3324 3854 3325 3855
rect 3399 3855 3405 3856
rect 3399 3854 3400 3855
rect 3324 3852 3400 3854
rect 3324 3851 3325 3852
rect 3319 3850 3325 3851
rect 3399 3851 3400 3852
rect 3404 3851 3405 3855
rect 3399 3850 3405 3851
rect 3486 3855 3493 3856
rect 3486 3851 3487 3855
rect 3492 3851 3493 3855
rect 3486 3850 3493 3851
rect 3510 3855 3516 3856
rect 3510 3851 3511 3855
rect 3515 3854 3516 3855
rect 3655 3855 3661 3856
rect 3655 3854 3656 3855
rect 3515 3852 3656 3854
rect 3515 3851 3516 3852
rect 3510 3850 3516 3851
rect 3655 3851 3656 3852
rect 3660 3851 3661 3855
rect 3655 3850 3661 3851
rect 3734 3855 3740 3856
rect 3734 3851 3735 3855
rect 3739 3854 3740 3855
rect 3823 3855 3829 3856
rect 3823 3854 3824 3855
rect 3739 3852 3824 3854
rect 3739 3851 3740 3852
rect 3734 3850 3740 3851
rect 3823 3851 3824 3852
rect 3828 3851 3829 3855
rect 3823 3850 3829 3851
rect 3068 3848 3074 3850
rect 2007 3846 2013 3847
rect 3072 3846 3074 3848
rect 3071 3845 3077 3846
rect 2262 3843 2269 3844
rect 655 3839 661 3840
rect 655 3835 656 3839
rect 660 3838 661 3839
rect 719 3839 725 3840
rect 719 3838 720 3839
rect 660 3836 720 3838
rect 660 3835 661 3836
rect 655 3834 661 3835
rect 719 3835 720 3836
rect 724 3835 725 3839
rect 719 3834 725 3835
rect 807 3839 813 3840
rect 807 3835 808 3839
rect 812 3838 813 3839
rect 871 3839 877 3840
rect 871 3838 872 3839
rect 812 3836 872 3838
rect 812 3835 813 3836
rect 807 3834 813 3835
rect 871 3835 872 3836
rect 876 3835 877 3839
rect 871 3834 877 3835
rect 959 3839 965 3840
rect 959 3835 960 3839
rect 964 3838 965 3839
rect 1015 3839 1021 3840
rect 1015 3838 1016 3839
rect 964 3836 1016 3838
rect 964 3835 965 3836
rect 959 3834 965 3835
rect 1015 3835 1016 3836
rect 1020 3835 1021 3839
rect 1015 3834 1021 3835
rect 1102 3839 1109 3840
rect 1102 3835 1103 3839
rect 1108 3835 1109 3839
rect 1102 3834 1109 3835
rect 1247 3839 1253 3840
rect 1247 3835 1248 3839
rect 1252 3838 1253 3839
rect 1295 3839 1301 3840
rect 1295 3838 1296 3839
rect 1252 3836 1296 3838
rect 1252 3835 1253 3836
rect 1247 3834 1253 3835
rect 1295 3835 1296 3836
rect 1300 3835 1301 3839
rect 1295 3834 1301 3835
rect 1383 3839 1389 3840
rect 1383 3835 1384 3839
rect 1388 3838 1389 3839
rect 1431 3839 1437 3840
rect 1431 3838 1432 3839
rect 1388 3836 1432 3838
rect 1388 3835 1389 3836
rect 1383 3834 1389 3835
rect 1431 3835 1432 3836
rect 1436 3835 1437 3839
rect 1431 3834 1437 3835
rect 1519 3839 1525 3840
rect 1519 3835 1520 3839
rect 1524 3838 1525 3839
rect 1559 3839 1565 3840
rect 1559 3838 1560 3839
rect 1524 3836 1560 3838
rect 1524 3835 1525 3836
rect 1519 3834 1525 3835
rect 1559 3835 1560 3836
rect 1564 3835 1565 3839
rect 1559 3834 1565 3835
rect 1647 3839 1653 3840
rect 1647 3835 1648 3839
rect 1652 3838 1653 3839
rect 1687 3839 1693 3840
rect 1687 3838 1688 3839
rect 1652 3836 1688 3838
rect 1652 3835 1653 3836
rect 1647 3834 1653 3835
rect 1687 3835 1688 3836
rect 1692 3835 1693 3839
rect 1687 3834 1693 3835
rect 1775 3839 1781 3840
rect 1775 3835 1776 3839
rect 1780 3838 1781 3839
rect 1815 3839 1821 3840
rect 1815 3838 1816 3839
rect 1780 3836 1816 3838
rect 1780 3835 1781 3836
rect 1775 3834 1781 3835
rect 1815 3835 1816 3836
rect 1820 3835 1821 3839
rect 1815 3834 1821 3835
rect 1903 3839 1909 3840
rect 1903 3835 1904 3839
rect 1908 3838 1909 3839
rect 1919 3839 1925 3840
rect 1919 3838 1920 3839
rect 1908 3836 1920 3838
rect 1908 3835 1909 3836
rect 1903 3834 1909 3835
rect 1919 3835 1920 3836
rect 1924 3835 1925 3839
rect 1919 3834 1925 3835
rect 2006 3839 2013 3840
rect 2006 3835 2007 3839
rect 2012 3835 2013 3839
rect 2262 3839 2263 3843
rect 2268 3839 2269 3843
rect 2262 3838 2269 3839
rect 2526 3843 2532 3844
rect 2526 3839 2527 3843
rect 2531 3842 2532 3843
rect 2559 3843 2565 3844
rect 2559 3842 2560 3843
rect 2531 3840 2560 3842
rect 2531 3839 2532 3840
rect 2526 3838 2532 3839
rect 2559 3839 2560 3840
rect 2564 3839 2565 3843
rect 2559 3838 2565 3839
rect 2831 3843 2837 3844
rect 2831 3839 2832 3843
rect 2836 3842 2837 3843
rect 2983 3843 2989 3844
rect 2983 3842 2984 3843
rect 2836 3840 2984 3842
rect 2836 3839 2837 3840
rect 2831 3838 2837 3839
rect 2983 3839 2984 3840
rect 2988 3839 2989 3843
rect 2983 3838 2989 3839
rect 2992 3840 3062 3842
rect 3071 3841 3072 3845
rect 3076 3841 3077 3845
rect 3287 3843 3293 3844
rect 3287 3842 3288 3843
rect 3071 3840 3077 3841
rect 3080 3840 3288 3842
rect 2006 3834 2013 3835
rect 2190 3835 2196 3836
rect 582 3831 588 3832
rect 582 3827 583 3831
rect 587 3827 588 3831
rect 582 3826 588 3827
rect 734 3831 740 3832
rect 734 3827 735 3831
rect 739 3827 740 3831
rect 734 3826 740 3827
rect 886 3831 892 3832
rect 886 3827 887 3831
rect 891 3827 892 3831
rect 886 3826 892 3827
rect 1030 3831 1036 3832
rect 1030 3827 1031 3831
rect 1035 3827 1036 3831
rect 1030 3826 1036 3827
rect 1174 3831 1180 3832
rect 1174 3827 1175 3831
rect 1179 3827 1180 3831
rect 1174 3826 1180 3827
rect 1310 3831 1316 3832
rect 1310 3827 1311 3831
rect 1315 3827 1316 3831
rect 1310 3826 1316 3827
rect 1446 3831 1452 3832
rect 1446 3827 1447 3831
rect 1451 3827 1452 3831
rect 1446 3826 1452 3827
rect 1574 3831 1580 3832
rect 1574 3827 1575 3831
rect 1579 3827 1580 3831
rect 1574 3826 1580 3827
rect 1702 3831 1708 3832
rect 1702 3827 1703 3831
rect 1707 3827 1708 3831
rect 1702 3826 1708 3827
rect 1830 3831 1836 3832
rect 1830 3827 1831 3831
rect 1835 3827 1836 3831
rect 1830 3826 1836 3827
rect 1934 3831 1940 3832
rect 1934 3827 1935 3831
rect 1939 3827 1940 3831
rect 2190 3831 2191 3835
rect 2195 3831 2196 3835
rect 2190 3830 2196 3831
rect 2486 3835 2492 3836
rect 2486 3831 2487 3835
rect 2491 3831 2492 3835
rect 2486 3830 2492 3831
rect 2758 3835 2764 3836
rect 2758 3831 2759 3835
rect 2763 3831 2764 3835
rect 2992 3834 2994 3840
rect 2758 3830 2764 3831
rect 2839 3832 2994 3834
rect 2998 3835 3004 3836
rect 1934 3826 1940 3827
rect 2254 3827 2260 3828
rect 2254 3826 2255 3827
rect 2241 3824 2255 3826
rect 718 3823 724 3824
rect 718 3822 719 3823
rect 633 3820 719 3822
rect 718 3819 719 3820
rect 723 3819 724 3823
rect 1294 3823 1300 3824
rect 1294 3822 1295 3823
rect 1225 3820 1295 3822
rect 718 3818 724 3819
rect 1294 3819 1295 3820
rect 1299 3819 1300 3823
rect 2254 3823 2255 3824
rect 2259 3823 2260 3827
rect 2630 3827 2636 3828
rect 2630 3826 2631 3827
rect 2537 3824 2631 3826
rect 2254 3822 2260 3823
rect 2630 3823 2631 3824
rect 2635 3823 2636 3827
rect 2839 3826 2841 3832
rect 2998 3831 2999 3835
rect 3003 3831 3004 3835
rect 3060 3834 3062 3840
rect 3080 3834 3082 3840
rect 3287 3839 3288 3840
rect 3292 3839 3293 3843
rect 3287 3838 3293 3839
rect 3479 3843 3485 3844
rect 3479 3839 3480 3843
rect 3484 3842 3485 3843
rect 3567 3843 3573 3844
rect 3567 3842 3568 3843
rect 3484 3840 3568 3842
rect 3484 3839 3485 3840
rect 3479 3838 3485 3839
rect 3567 3839 3568 3840
rect 3572 3839 3573 3843
rect 3567 3838 3573 3839
rect 3646 3843 3652 3844
rect 3646 3839 3647 3843
rect 3651 3842 3652 3843
rect 3655 3843 3661 3844
rect 3655 3842 3656 3843
rect 3651 3840 3656 3842
rect 3651 3839 3652 3840
rect 3646 3838 3652 3839
rect 3655 3839 3656 3840
rect 3660 3839 3661 3843
rect 3967 3843 3973 3844
rect 3967 3842 3968 3843
rect 3655 3838 3661 3839
rect 3852 3840 3968 3842
rect 3060 3832 3082 3834
rect 3214 3835 3220 3836
rect 2998 3830 3004 3831
rect 3214 3831 3215 3835
rect 3219 3831 3220 3835
rect 3214 3830 3220 3831
rect 3406 3835 3412 3836
rect 3406 3831 3407 3835
rect 3411 3831 3412 3835
rect 3406 3830 3412 3831
rect 3582 3835 3588 3836
rect 3582 3831 3583 3835
rect 3587 3831 3588 3835
rect 3582 3830 3588 3831
rect 3750 3835 3756 3836
rect 3750 3831 3751 3835
rect 3755 3831 3756 3835
rect 3750 3830 3756 3831
rect 3390 3827 3396 3828
rect 3390 3826 3391 3827
rect 2809 3824 2841 3826
rect 3265 3824 3391 3826
rect 2630 3822 2636 3823
rect 3390 3823 3391 3824
rect 3395 3823 3396 3827
rect 3510 3827 3516 3828
rect 3510 3826 3511 3827
rect 3457 3824 3511 3826
rect 3390 3822 3396 3823
rect 3510 3823 3511 3824
rect 3515 3823 3516 3827
rect 3852 3826 3854 3840
rect 3967 3839 3968 3840
rect 3972 3839 3973 3843
rect 3967 3838 3973 3839
rect 3894 3835 3900 3836
rect 3894 3831 3895 3835
rect 3899 3831 3900 3835
rect 3894 3830 3900 3831
rect 3966 3827 3972 3828
rect 3966 3826 3967 3827
rect 3801 3824 3854 3826
rect 3945 3824 3967 3826
rect 3510 3822 3516 3823
rect 3966 3823 3967 3824
rect 3971 3823 3972 3827
rect 3966 3822 3972 3823
rect 1294 3818 1300 3819
rect 2070 3816 2076 3817
rect 110 3812 116 3813
rect 110 3808 111 3812
rect 115 3808 116 3812
rect 110 3807 116 3808
rect 2030 3812 2036 3813
rect 2030 3808 2031 3812
rect 2035 3808 2036 3812
rect 2070 3812 2071 3816
rect 2075 3812 2076 3816
rect 2070 3811 2076 3812
rect 3990 3816 3996 3817
rect 3990 3812 3991 3816
rect 3995 3812 3996 3816
rect 3990 3811 3996 3812
rect 2030 3807 2036 3808
rect 2070 3799 2076 3800
rect 110 3795 116 3796
rect 110 3791 111 3795
rect 115 3791 116 3795
rect 2030 3795 2036 3796
rect 2030 3791 2031 3795
rect 2035 3791 2036 3795
rect 2070 3795 2071 3799
rect 2075 3795 2076 3799
rect 3990 3799 3996 3800
rect 3990 3795 3991 3799
rect 3995 3795 3996 3799
rect 2070 3794 2076 3795
rect 2190 3794 2196 3795
rect 110 3790 116 3791
rect 582 3790 588 3791
rect 582 3786 583 3790
rect 587 3786 588 3790
rect 582 3785 588 3786
rect 734 3790 740 3791
rect 734 3786 735 3790
rect 739 3786 740 3790
rect 734 3785 740 3786
rect 886 3790 892 3791
rect 886 3786 887 3790
rect 891 3786 892 3790
rect 886 3785 892 3786
rect 1030 3790 1036 3791
rect 1030 3786 1031 3790
rect 1035 3786 1036 3790
rect 1030 3785 1036 3786
rect 1174 3790 1180 3791
rect 1174 3786 1175 3790
rect 1179 3786 1180 3790
rect 1174 3785 1180 3786
rect 1310 3790 1316 3791
rect 1310 3786 1311 3790
rect 1315 3786 1316 3790
rect 1310 3785 1316 3786
rect 1446 3790 1452 3791
rect 1446 3786 1447 3790
rect 1451 3786 1452 3790
rect 1446 3785 1452 3786
rect 1574 3790 1580 3791
rect 1574 3786 1575 3790
rect 1579 3786 1580 3790
rect 1574 3785 1580 3786
rect 1702 3790 1708 3791
rect 1702 3786 1703 3790
rect 1707 3786 1708 3790
rect 1702 3785 1708 3786
rect 1830 3790 1836 3791
rect 1830 3786 1831 3790
rect 1835 3786 1836 3790
rect 1830 3785 1836 3786
rect 1934 3790 1940 3791
rect 2030 3790 2036 3791
rect 2190 3790 2191 3794
rect 2195 3790 2196 3794
rect 1934 3786 1935 3790
rect 1939 3786 1940 3790
rect 2190 3789 2196 3790
rect 2486 3794 2492 3795
rect 2486 3790 2487 3794
rect 2491 3790 2492 3794
rect 2486 3789 2492 3790
rect 2758 3794 2764 3795
rect 2758 3790 2759 3794
rect 2763 3790 2764 3794
rect 2758 3789 2764 3790
rect 2998 3794 3004 3795
rect 2998 3790 2999 3794
rect 3003 3790 3004 3794
rect 2998 3789 3004 3790
rect 3214 3794 3220 3795
rect 3214 3790 3215 3794
rect 3219 3790 3220 3794
rect 3214 3789 3220 3790
rect 3406 3794 3412 3795
rect 3406 3790 3407 3794
rect 3411 3790 3412 3794
rect 3406 3789 3412 3790
rect 3582 3794 3588 3795
rect 3582 3790 3583 3794
rect 3587 3790 3588 3794
rect 3582 3789 3588 3790
rect 3750 3794 3756 3795
rect 3750 3790 3751 3794
rect 3755 3790 3756 3794
rect 3750 3789 3756 3790
rect 3894 3794 3900 3795
rect 3990 3794 3996 3795
rect 3894 3790 3895 3794
rect 3899 3790 3900 3794
rect 3894 3789 3900 3790
rect 1934 3785 1940 3786
rect 3390 3779 3396 3780
rect 3390 3775 3391 3779
rect 3395 3778 3396 3779
rect 3550 3779 3556 3780
rect 3550 3778 3551 3779
rect 3395 3776 3551 3778
rect 3395 3775 3396 3776
rect 3390 3774 3396 3775
rect 3550 3775 3551 3776
rect 3555 3775 3556 3779
rect 3550 3774 3556 3775
rect 1294 3763 1300 3764
rect 1294 3759 1295 3763
rect 1299 3762 1300 3763
rect 1838 3763 1844 3764
rect 1838 3762 1839 3763
rect 1299 3760 1839 3762
rect 1299 3759 1300 3760
rect 1294 3758 1300 3759
rect 1838 3759 1839 3760
rect 1843 3759 1844 3763
rect 1838 3758 1844 3759
rect 2110 3762 2116 3763
rect 2110 3758 2111 3762
rect 2115 3758 2116 3762
rect 2070 3757 2076 3758
rect 2110 3757 2116 3758
rect 2334 3762 2340 3763
rect 2334 3758 2335 3762
rect 2339 3758 2340 3762
rect 2334 3757 2340 3758
rect 2558 3762 2564 3763
rect 2558 3758 2559 3762
rect 2563 3758 2564 3762
rect 2558 3757 2564 3758
rect 2774 3762 2780 3763
rect 2774 3758 2775 3762
rect 2779 3758 2780 3762
rect 2774 3757 2780 3758
rect 2974 3762 2980 3763
rect 2974 3758 2975 3762
rect 2979 3758 2980 3762
rect 2974 3757 2980 3758
rect 3158 3762 3164 3763
rect 3158 3758 3159 3762
rect 3163 3758 3164 3762
rect 3158 3757 3164 3758
rect 3326 3762 3332 3763
rect 3326 3758 3327 3762
rect 3331 3758 3332 3762
rect 3326 3757 3332 3758
rect 3478 3762 3484 3763
rect 3478 3758 3479 3762
rect 3483 3758 3484 3762
rect 3478 3757 3484 3758
rect 3622 3762 3628 3763
rect 3622 3758 3623 3762
rect 3627 3758 3628 3762
rect 3622 3757 3628 3758
rect 3766 3762 3772 3763
rect 3766 3758 3767 3762
rect 3771 3758 3772 3762
rect 3766 3757 3772 3758
rect 3894 3762 3900 3763
rect 3894 3758 3895 3762
rect 3899 3758 3900 3762
rect 3894 3757 3900 3758
rect 3990 3757 3996 3758
rect 2070 3753 2071 3757
rect 2075 3753 2076 3757
rect 2070 3752 2076 3753
rect 3990 3753 3991 3757
rect 3995 3753 3996 3757
rect 3990 3752 3996 3753
rect 598 3746 604 3747
rect 598 3742 599 3746
rect 603 3742 604 3746
rect 110 3741 116 3742
rect 598 3741 604 3742
rect 718 3746 724 3747
rect 718 3742 719 3746
rect 723 3742 724 3746
rect 718 3741 724 3742
rect 846 3746 852 3747
rect 846 3742 847 3746
rect 851 3742 852 3746
rect 846 3741 852 3742
rect 982 3746 988 3747
rect 982 3742 983 3746
rect 987 3742 988 3746
rect 982 3741 988 3742
rect 1110 3746 1116 3747
rect 1110 3742 1111 3746
rect 1115 3742 1116 3746
rect 1110 3741 1116 3742
rect 1238 3746 1244 3747
rect 1238 3742 1239 3746
rect 1243 3742 1244 3746
rect 1238 3741 1244 3742
rect 1366 3746 1372 3747
rect 1366 3742 1367 3746
rect 1371 3742 1372 3746
rect 1366 3741 1372 3742
rect 1494 3746 1500 3747
rect 1494 3742 1495 3746
rect 1499 3742 1500 3746
rect 1494 3741 1500 3742
rect 1630 3746 1636 3747
rect 1630 3742 1631 3746
rect 1635 3742 1636 3746
rect 1630 3741 1636 3742
rect 1766 3746 1772 3747
rect 1766 3742 1767 3746
rect 1771 3742 1772 3746
rect 1766 3741 1772 3742
rect 2030 3741 2036 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 110 3736 116 3737
rect 2030 3737 2031 3741
rect 2035 3737 2036 3741
rect 2030 3736 2036 3737
rect 2070 3740 2076 3741
rect 2070 3736 2071 3740
rect 2075 3736 2076 3740
rect 2070 3735 2076 3736
rect 3990 3740 3996 3741
rect 3990 3736 3991 3740
rect 3995 3736 3996 3740
rect 3990 3735 3996 3736
rect 2262 3731 2268 3732
rect 2262 3730 2263 3731
rect 2161 3728 2263 3730
rect 2262 3727 2263 3728
rect 2267 3727 2268 3731
rect 2698 3731 2704 3732
rect 2698 3730 2699 3731
rect 2609 3728 2699 3730
rect 2262 3726 2268 3727
rect 2698 3727 2699 3728
rect 2703 3727 2704 3731
rect 2886 3731 2892 3732
rect 2886 3730 2887 3731
rect 2825 3728 2887 3730
rect 2698 3726 2704 3727
rect 2886 3727 2887 3728
rect 2891 3727 2892 3731
rect 3142 3731 3148 3732
rect 3142 3730 3143 3731
rect 3025 3728 3143 3730
rect 2886 3726 2892 3727
rect 3142 3727 3143 3728
rect 3147 3727 3148 3731
rect 3142 3726 3148 3727
rect 3646 3731 3652 3732
rect 3646 3727 3647 3731
rect 3651 3727 3652 3731
rect 3646 3726 3652 3727
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 110 3719 116 3720
rect 2030 3724 2036 3725
rect 2030 3720 2031 3724
rect 2035 3720 2036 3724
rect 2030 3719 2036 3720
rect 2110 3721 2116 3722
rect 2110 3717 2111 3721
rect 2115 3717 2116 3721
rect 2110 3716 2116 3717
rect 2334 3721 2340 3722
rect 2334 3717 2335 3721
rect 2339 3717 2340 3721
rect 2334 3716 2340 3717
rect 2558 3721 2564 3722
rect 2558 3717 2559 3721
rect 2563 3717 2564 3721
rect 2558 3716 2564 3717
rect 2774 3721 2780 3722
rect 2774 3717 2775 3721
rect 2779 3717 2780 3721
rect 2774 3716 2780 3717
rect 2974 3721 2980 3722
rect 2974 3717 2975 3721
rect 2979 3717 2980 3721
rect 2974 3716 2980 3717
rect 3158 3721 3164 3722
rect 3158 3717 3159 3721
rect 3163 3717 3164 3721
rect 3158 3716 3164 3717
rect 3326 3721 3332 3722
rect 3326 3717 3327 3721
rect 3331 3717 3332 3721
rect 3326 3716 3332 3717
rect 3478 3721 3484 3722
rect 3478 3717 3479 3721
rect 3483 3717 3484 3721
rect 3478 3716 3484 3717
rect 3622 3721 3628 3722
rect 3622 3717 3623 3721
rect 3627 3717 3628 3721
rect 3622 3716 3628 3717
rect 3766 3721 3772 3722
rect 3766 3717 3767 3721
rect 3771 3717 3772 3721
rect 3766 3716 3772 3717
rect 3894 3721 3900 3722
rect 3894 3717 3895 3721
rect 3899 3717 3900 3721
rect 3894 3716 3900 3717
rect 702 3715 708 3716
rect 702 3714 703 3715
rect 649 3712 703 3714
rect 702 3711 703 3712
rect 707 3711 708 3715
rect 966 3715 972 3716
rect 966 3714 967 3715
rect 897 3712 967 3714
rect 702 3710 708 3711
rect 966 3711 967 3712
rect 971 3711 972 3715
rect 1071 3715 1077 3716
rect 1071 3714 1072 3715
rect 1033 3712 1072 3714
rect 966 3710 972 3711
rect 1071 3711 1072 3712
rect 1076 3711 1077 3715
rect 1071 3710 1077 3711
rect 1102 3715 1108 3716
rect 1102 3711 1103 3715
rect 1107 3711 1108 3715
rect 1350 3715 1356 3716
rect 1350 3714 1351 3715
rect 1289 3712 1351 3714
rect 1102 3710 1108 3711
rect 1350 3711 1351 3712
rect 1355 3711 1356 3715
rect 1350 3710 1356 3711
rect 2183 3711 2189 3712
rect 2183 3707 2184 3711
rect 2188 3710 2189 3711
rect 2319 3711 2325 3712
rect 2319 3710 2320 3711
rect 2188 3708 2320 3710
rect 2188 3707 2189 3708
rect 2183 3706 2189 3707
rect 2319 3707 2320 3708
rect 2324 3707 2325 3711
rect 2319 3706 2325 3707
rect 2335 3711 2341 3712
rect 2335 3707 2336 3711
rect 2340 3710 2341 3711
rect 2407 3711 2413 3712
rect 2407 3710 2408 3711
rect 2340 3708 2408 3710
rect 2340 3707 2341 3708
rect 2335 3706 2341 3707
rect 2407 3707 2408 3708
rect 2412 3707 2413 3711
rect 2407 3706 2413 3707
rect 2630 3711 2637 3712
rect 2630 3707 2631 3711
rect 2636 3707 2637 3711
rect 2630 3706 2637 3707
rect 2698 3711 2704 3712
rect 2698 3707 2699 3711
rect 2703 3710 2704 3711
rect 2847 3711 2853 3712
rect 2847 3710 2848 3711
rect 2703 3708 2848 3710
rect 2703 3707 2704 3708
rect 2698 3706 2704 3707
rect 2847 3707 2848 3708
rect 2852 3707 2853 3711
rect 2847 3706 2853 3707
rect 3047 3711 3053 3712
rect 3047 3707 3048 3711
rect 3052 3710 3053 3711
rect 3143 3711 3149 3712
rect 3143 3710 3144 3711
rect 3052 3708 3144 3710
rect 3052 3707 3053 3708
rect 3047 3706 3053 3707
rect 3143 3707 3144 3708
rect 3148 3707 3149 3711
rect 3143 3706 3149 3707
rect 3231 3711 3237 3712
rect 3231 3707 3232 3711
rect 3236 3710 3237 3711
rect 3311 3711 3317 3712
rect 3311 3710 3312 3711
rect 3236 3708 3312 3710
rect 3236 3707 3237 3708
rect 3231 3706 3237 3707
rect 3311 3707 3312 3708
rect 3316 3707 3317 3711
rect 3311 3706 3317 3707
rect 3399 3711 3405 3712
rect 3399 3707 3400 3711
rect 3404 3710 3405 3711
rect 3463 3711 3469 3712
rect 3463 3710 3464 3711
rect 3404 3708 3464 3710
rect 3404 3707 3405 3708
rect 3399 3706 3405 3707
rect 3463 3707 3464 3708
rect 3468 3707 3469 3711
rect 3463 3706 3469 3707
rect 3550 3711 3557 3712
rect 3550 3707 3551 3711
rect 3556 3707 3557 3711
rect 3550 3706 3557 3707
rect 3695 3711 3701 3712
rect 3695 3707 3696 3711
rect 3700 3710 3701 3711
rect 3751 3711 3757 3712
rect 3751 3710 3752 3711
rect 3700 3708 3752 3710
rect 3700 3707 3701 3708
rect 3695 3706 3701 3707
rect 3751 3707 3752 3708
rect 3756 3707 3757 3711
rect 3751 3706 3757 3707
rect 3839 3711 3845 3712
rect 3839 3707 3840 3711
rect 3844 3710 3845 3711
rect 3879 3711 3885 3712
rect 3879 3710 3880 3711
rect 3844 3708 3880 3710
rect 3844 3707 3845 3708
rect 3839 3706 3845 3707
rect 3879 3707 3880 3708
rect 3884 3707 3885 3711
rect 3879 3706 3885 3707
rect 3966 3711 3973 3712
rect 3966 3707 3967 3711
rect 3972 3707 3973 3711
rect 3966 3706 3973 3707
rect 598 3705 604 3706
rect 598 3701 599 3705
rect 603 3701 604 3705
rect 598 3700 604 3701
rect 718 3705 724 3706
rect 718 3701 719 3705
rect 723 3701 724 3705
rect 718 3700 724 3701
rect 846 3705 852 3706
rect 846 3701 847 3705
rect 851 3701 852 3705
rect 846 3700 852 3701
rect 982 3705 988 3706
rect 982 3701 983 3705
rect 987 3701 988 3705
rect 982 3700 988 3701
rect 1110 3705 1116 3706
rect 1110 3701 1111 3705
rect 1115 3701 1116 3705
rect 1110 3700 1116 3701
rect 1238 3705 1244 3706
rect 1238 3701 1239 3705
rect 1243 3701 1244 3705
rect 1238 3700 1244 3701
rect 1366 3705 1372 3706
rect 1366 3701 1367 3705
rect 1371 3701 1372 3705
rect 1366 3700 1372 3701
rect 1494 3705 1500 3706
rect 1494 3701 1495 3705
rect 1499 3701 1500 3705
rect 1494 3700 1500 3701
rect 1630 3705 1636 3706
rect 1630 3701 1631 3705
rect 1635 3701 1636 3705
rect 1630 3700 1636 3701
rect 1766 3705 1772 3706
rect 1766 3701 1767 3705
rect 1771 3701 1772 3705
rect 1766 3700 1772 3701
rect 671 3695 677 3696
rect 671 3691 672 3695
rect 676 3694 677 3695
rect 703 3695 709 3696
rect 703 3694 704 3695
rect 676 3692 704 3694
rect 676 3691 677 3692
rect 671 3690 677 3691
rect 703 3691 704 3692
rect 708 3691 709 3695
rect 703 3690 709 3691
rect 782 3695 788 3696
rect 782 3691 783 3695
rect 787 3694 788 3695
rect 791 3695 797 3696
rect 791 3694 792 3695
rect 787 3692 792 3694
rect 787 3691 788 3692
rect 782 3690 788 3691
rect 791 3691 792 3692
rect 796 3691 797 3695
rect 919 3695 925 3696
rect 919 3694 920 3695
rect 791 3690 797 3691
rect 800 3692 920 3694
rect 702 3687 708 3688
rect 702 3683 703 3687
rect 707 3686 708 3687
rect 800 3686 802 3692
rect 919 3691 920 3692
rect 924 3691 925 3695
rect 919 3690 925 3691
rect 966 3695 972 3696
rect 966 3691 967 3695
rect 971 3694 972 3695
rect 1055 3695 1061 3696
rect 1055 3694 1056 3695
rect 971 3692 1056 3694
rect 971 3691 972 3692
rect 966 3690 972 3691
rect 1055 3691 1056 3692
rect 1060 3691 1061 3695
rect 1055 3690 1061 3691
rect 1071 3695 1077 3696
rect 1071 3691 1072 3695
rect 1076 3694 1077 3695
rect 1183 3695 1189 3696
rect 1183 3694 1184 3695
rect 1076 3692 1184 3694
rect 1076 3691 1077 3692
rect 1071 3690 1077 3691
rect 1183 3691 1184 3692
rect 1188 3691 1189 3695
rect 1183 3690 1189 3691
rect 1311 3695 1317 3696
rect 1311 3691 1312 3695
rect 1316 3694 1317 3695
rect 1351 3695 1357 3696
rect 1351 3694 1352 3695
rect 1316 3692 1352 3694
rect 1316 3691 1317 3692
rect 1311 3690 1317 3691
rect 1351 3691 1352 3692
rect 1356 3691 1357 3695
rect 1351 3690 1357 3691
rect 1439 3695 1445 3696
rect 1439 3691 1440 3695
rect 1444 3694 1445 3695
rect 1479 3695 1485 3696
rect 1479 3694 1480 3695
rect 1444 3692 1480 3694
rect 1444 3691 1445 3692
rect 1439 3690 1445 3691
rect 1479 3691 1480 3692
rect 1484 3691 1485 3695
rect 1479 3690 1485 3691
rect 1567 3695 1573 3696
rect 1567 3691 1568 3695
rect 1572 3694 1573 3695
rect 1615 3695 1621 3696
rect 1615 3694 1616 3695
rect 1572 3692 1616 3694
rect 1572 3691 1573 3692
rect 1567 3690 1573 3691
rect 1615 3691 1616 3692
rect 1620 3691 1621 3695
rect 1615 3690 1621 3691
rect 1703 3695 1709 3696
rect 1703 3691 1704 3695
rect 1708 3694 1709 3695
rect 1751 3695 1757 3696
rect 1751 3694 1752 3695
rect 1708 3692 1752 3694
rect 1708 3691 1709 3692
rect 1703 3690 1709 3691
rect 1751 3691 1752 3692
rect 1756 3691 1757 3695
rect 1751 3690 1757 3691
rect 1838 3695 1845 3696
rect 1838 3691 1839 3695
rect 1844 3691 1845 3695
rect 1838 3690 1845 3691
rect 3142 3695 3148 3696
rect 3142 3691 3143 3695
rect 3147 3694 3148 3695
rect 3147 3692 3578 3694
rect 3147 3691 3148 3692
rect 3142 3690 3148 3691
rect 707 3684 802 3686
rect 1350 3687 1356 3688
rect 707 3683 708 3684
rect 702 3682 708 3683
rect 1350 3683 1351 3687
rect 1355 3686 1356 3687
rect 2050 3687 2056 3688
rect 1355 3684 1474 3686
rect 1355 3683 1356 3684
rect 1350 3682 1356 3683
rect 543 3679 549 3680
rect 543 3675 544 3679
rect 548 3678 549 3679
rect 599 3679 605 3680
rect 599 3678 600 3679
rect 548 3676 600 3678
rect 548 3675 549 3676
rect 543 3674 549 3675
rect 599 3675 600 3676
rect 604 3675 605 3679
rect 599 3674 605 3675
rect 686 3679 693 3680
rect 686 3675 687 3679
rect 692 3675 693 3679
rect 686 3674 693 3675
rect 831 3679 837 3680
rect 831 3675 832 3679
rect 836 3678 837 3679
rect 887 3679 893 3680
rect 887 3678 888 3679
rect 836 3676 888 3678
rect 836 3675 837 3676
rect 831 3674 837 3675
rect 887 3675 888 3676
rect 892 3675 893 3679
rect 887 3674 893 3675
rect 910 3679 916 3680
rect 910 3675 911 3679
rect 915 3678 916 3679
rect 975 3679 981 3680
rect 975 3678 976 3679
rect 915 3676 976 3678
rect 915 3675 916 3676
rect 910 3674 916 3675
rect 975 3675 976 3676
rect 980 3675 981 3679
rect 975 3674 981 3675
rect 1119 3679 1125 3680
rect 1119 3675 1120 3679
rect 1124 3678 1125 3679
rect 1175 3679 1181 3680
rect 1175 3678 1176 3679
rect 1124 3676 1176 3678
rect 1124 3675 1125 3676
rect 1119 3674 1125 3675
rect 1175 3675 1176 3676
rect 1180 3675 1181 3679
rect 1175 3674 1181 3675
rect 1263 3679 1269 3680
rect 1263 3675 1264 3679
rect 1268 3678 1269 3679
rect 1319 3679 1325 3680
rect 1319 3678 1320 3679
rect 1268 3676 1320 3678
rect 1268 3675 1269 3676
rect 1263 3674 1269 3675
rect 1319 3675 1320 3676
rect 1324 3675 1325 3679
rect 1319 3674 1325 3675
rect 1407 3679 1413 3680
rect 1407 3675 1408 3679
rect 1412 3678 1413 3679
rect 1463 3679 1469 3680
rect 1463 3678 1464 3679
rect 1412 3676 1464 3678
rect 1412 3675 1413 3676
rect 1407 3674 1413 3675
rect 1463 3675 1464 3676
rect 1468 3675 1469 3679
rect 1472 3678 1474 3684
rect 2050 3683 2051 3687
rect 2055 3686 2056 3687
rect 2183 3687 2189 3688
rect 2183 3686 2184 3687
rect 2055 3684 2184 3686
rect 2055 3683 2056 3684
rect 2050 3682 2056 3683
rect 2183 3683 2184 3684
rect 2188 3683 2189 3687
rect 2327 3687 2333 3688
rect 2327 3686 2328 3687
rect 2183 3682 2189 3683
rect 2216 3684 2328 3686
rect 1551 3679 1557 3680
rect 1551 3678 1552 3679
rect 1472 3676 1552 3678
rect 1463 3674 1469 3675
rect 1551 3675 1552 3676
rect 1556 3675 1557 3679
rect 1551 3674 1557 3675
rect 2110 3679 2116 3680
rect 2110 3675 2111 3679
rect 2115 3675 2116 3679
rect 2110 3674 2116 3675
rect 470 3671 476 3672
rect 470 3667 471 3671
rect 475 3667 476 3671
rect 470 3666 476 3667
rect 614 3671 620 3672
rect 614 3667 615 3671
rect 619 3667 620 3671
rect 614 3666 620 3667
rect 758 3671 764 3672
rect 758 3667 759 3671
rect 763 3667 764 3671
rect 758 3666 764 3667
rect 902 3671 908 3672
rect 902 3667 903 3671
rect 907 3667 908 3671
rect 902 3666 908 3667
rect 1046 3671 1052 3672
rect 1046 3667 1047 3671
rect 1051 3667 1052 3671
rect 1046 3666 1052 3667
rect 1190 3671 1196 3672
rect 1190 3667 1191 3671
rect 1195 3667 1196 3671
rect 1190 3666 1196 3667
rect 1334 3671 1340 3672
rect 1334 3667 1335 3671
rect 1339 3667 1340 3671
rect 1334 3666 1340 3667
rect 1478 3671 1484 3672
rect 1478 3667 1479 3671
rect 1483 3667 1484 3671
rect 2216 3670 2218 3684
rect 2327 3683 2328 3684
rect 2332 3683 2333 3687
rect 2327 3682 2333 3683
rect 2511 3687 2517 3688
rect 2511 3683 2512 3687
rect 2516 3686 2517 3687
rect 2607 3687 2613 3688
rect 2607 3686 2608 3687
rect 2516 3684 2608 3686
rect 2516 3683 2517 3684
rect 2511 3682 2517 3683
rect 2607 3683 2608 3684
rect 2612 3683 2613 3687
rect 2607 3682 2613 3683
rect 2695 3687 2701 3688
rect 2695 3683 2696 3687
rect 2700 3686 2701 3687
rect 2799 3687 2805 3688
rect 2799 3686 2800 3687
rect 2700 3684 2800 3686
rect 2700 3683 2701 3684
rect 2695 3682 2701 3683
rect 2799 3683 2800 3684
rect 2804 3683 2805 3687
rect 2799 3682 2805 3683
rect 2886 3687 2893 3688
rect 2886 3683 2887 3687
rect 2892 3683 2893 3687
rect 2886 3682 2893 3683
rect 3079 3687 3085 3688
rect 3079 3683 3080 3687
rect 3084 3686 3085 3687
rect 3183 3687 3189 3688
rect 3183 3686 3184 3687
rect 3084 3684 3184 3686
rect 3084 3683 3085 3684
rect 3079 3682 3085 3683
rect 3183 3683 3184 3684
rect 3188 3683 3189 3687
rect 3183 3682 3189 3683
rect 3271 3687 3277 3688
rect 3271 3683 3272 3687
rect 3276 3686 3277 3687
rect 3375 3687 3381 3688
rect 3375 3686 3376 3687
rect 3276 3684 3376 3686
rect 3276 3683 3277 3684
rect 3271 3682 3277 3683
rect 3375 3683 3376 3684
rect 3380 3683 3381 3687
rect 3375 3682 3381 3683
rect 3463 3687 3469 3688
rect 3463 3683 3464 3687
rect 3468 3686 3469 3687
rect 3567 3687 3573 3688
rect 3567 3686 3568 3687
rect 3468 3684 3568 3686
rect 3468 3683 3469 3684
rect 3463 3682 3469 3683
rect 3567 3683 3568 3684
rect 3572 3683 3573 3687
rect 3576 3686 3578 3692
rect 3655 3687 3661 3688
rect 3655 3686 3656 3687
rect 3576 3684 3656 3686
rect 3567 3682 3573 3683
rect 3655 3683 3656 3684
rect 3660 3683 3661 3687
rect 3655 3682 3661 3683
rect 2254 3679 2260 3680
rect 2254 3675 2255 3679
rect 2259 3675 2260 3679
rect 2254 3674 2260 3675
rect 2438 3679 2444 3680
rect 2438 3675 2439 3679
rect 2443 3675 2444 3679
rect 2438 3674 2444 3675
rect 2622 3679 2628 3680
rect 2622 3675 2623 3679
rect 2627 3675 2628 3679
rect 2622 3674 2628 3675
rect 2814 3679 2820 3680
rect 2814 3675 2815 3679
rect 2819 3675 2820 3679
rect 2814 3674 2820 3675
rect 3006 3679 3012 3680
rect 3006 3675 3007 3679
rect 3011 3675 3012 3679
rect 3006 3674 3012 3675
rect 3198 3679 3204 3680
rect 3198 3675 3199 3679
rect 3203 3675 3204 3679
rect 3198 3674 3204 3675
rect 3390 3679 3396 3680
rect 3390 3675 3391 3679
rect 3395 3675 3396 3679
rect 3390 3674 3396 3675
rect 3582 3679 3588 3680
rect 3582 3675 3583 3679
rect 3587 3675 3588 3679
rect 3582 3674 3588 3675
rect 2335 3671 2341 3672
rect 2335 3670 2336 3671
rect 2161 3668 2218 3670
rect 2305 3668 2336 3670
rect 1478 3666 1484 3667
rect 2335 3667 2336 3668
rect 2340 3667 2341 3671
rect 3182 3671 3188 3672
rect 3182 3670 3183 3671
rect 3057 3668 3183 3670
rect 2335 3666 2341 3667
rect 2430 3667 2436 3668
rect 598 3663 604 3664
rect 598 3662 599 3663
rect 521 3660 599 3662
rect 598 3659 599 3660
rect 603 3659 604 3663
rect 1174 3663 1180 3664
rect 1174 3662 1175 3663
rect 1097 3660 1175 3662
rect 598 3658 604 3659
rect 782 3659 788 3660
rect 782 3655 783 3659
rect 787 3655 788 3659
rect 1174 3659 1175 3660
rect 1179 3659 1180 3663
rect 2430 3663 2431 3667
rect 2435 3663 2436 3667
rect 3182 3667 3183 3668
rect 3187 3667 3188 3671
rect 3182 3666 3188 3667
rect 2430 3662 2436 3663
rect 1174 3658 1180 3659
rect 2070 3660 2076 3661
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 3990 3660 3996 3661
rect 3990 3656 3991 3660
rect 3995 3656 3996 3660
rect 3990 3655 3996 3656
rect 782 3654 788 3655
rect 110 3652 116 3653
rect 110 3648 111 3652
rect 115 3648 116 3652
rect 110 3647 116 3648
rect 2030 3652 2036 3653
rect 2030 3648 2031 3652
rect 2035 3648 2036 3652
rect 2030 3647 2036 3648
rect 2070 3643 2076 3644
rect 2070 3639 2071 3643
rect 2075 3639 2076 3643
rect 3990 3643 3996 3644
rect 3990 3639 3991 3643
rect 3995 3639 3996 3643
rect 2070 3638 2076 3639
rect 2110 3638 2116 3639
rect 110 3635 116 3636
rect 110 3631 111 3635
rect 115 3631 116 3635
rect 2030 3635 2036 3636
rect 2030 3631 2031 3635
rect 2035 3631 2036 3635
rect 2110 3634 2111 3638
rect 2115 3634 2116 3638
rect 2110 3633 2116 3634
rect 2254 3638 2260 3639
rect 2254 3634 2255 3638
rect 2259 3634 2260 3638
rect 2254 3633 2260 3634
rect 2438 3638 2444 3639
rect 2438 3634 2439 3638
rect 2443 3634 2444 3638
rect 2438 3633 2444 3634
rect 2622 3638 2628 3639
rect 2622 3634 2623 3638
rect 2627 3634 2628 3638
rect 2622 3633 2628 3634
rect 2814 3638 2820 3639
rect 2814 3634 2815 3638
rect 2819 3634 2820 3638
rect 2814 3633 2820 3634
rect 3006 3638 3012 3639
rect 3006 3634 3007 3638
rect 3011 3634 3012 3638
rect 3006 3633 3012 3634
rect 3198 3638 3204 3639
rect 3198 3634 3199 3638
rect 3203 3634 3204 3638
rect 3198 3633 3204 3634
rect 3390 3638 3396 3639
rect 3390 3634 3391 3638
rect 3395 3634 3396 3638
rect 3390 3633 3396 3634
rect 3582 3638 3588 3639
rect 3990 3638 3996 3639
rect 3582 3634 3583 3638
rect 3587 3634 3588 3638
rect 3582 3633 3588 3634
rect 110 3630 116 3631
rect 470 3630 476 3631
rect 470 3626 471 3630
rect 475 3626 476 3630
rect 470 3625 476 3626
rect 614 3630 620 3631
rect 614 3626 615 3630
rect 619 3626 620 3630
rect 614 3625 620 3626
rect 758 3630 764 3631
rect 758 3626 759 3630
rect 763 3626 764 3630
rect 758 3625 764 3626
rect 902 3630 908 3631
rect 902 3626 903 3630
rect 907 3626 908 3630
rect 902 3625 908 3626
rect 1046 3630 1052 3631
rect 1046 3626 1047 3630
rect 1051 3626 1052 3630
rect 1046 3625 1052 3626
rect 1190 3630 1196 3631
rect 1190 3626 1191 3630
rect 1195 3626 1196 3630
rect 1190 3625 1196 3626
rect 1334 3630 1340 3631
rect 1334 3626 1335 3630
rect 1339 3626 1340 3630
rect 1334 3625 1340 3626
rect 1478 3630 1484 3631
rect 2030 3630 2036 3631
rect 1478 3626 1479 3630
rect 1483 3626 1484 3630
rect 1478 3625 1484 3626
rect 246 3598 252 3599
rect 246 3594 247 3598
rect 251 3594 252 3598
rect 110 3593 116 3594
rect 246 3593 252 3594
rect 374 3598 380 3599
rect 374 3594 375 3598
rect 379 3594 380 3598
rect 374 3593 380 3594
rect 518 3598 524 3599
rect 518 3594 519 3598
rect 523 3594 524 3598
rect 518 3593 524 3594
rect 678 3598 684 3599
rect 678 3594 679 3598
rect 683 3594 684 3598
rect 678 3593 684 3594
rect 846 3598 852 3599
rect 846 3594 847 3598
rect 851 3594 852 3598
rect 846 3593 852 3594
rect 1022 3598 1028 3599
rect 1022 3594 1023 3598
rect 1027 3594 1028 3598
rect 1022 3593 1028 3594
rect 1206 3598 1212 3599
rect 1206 3594 1207 3598
rect 1211 3594 1212 3598
rect 1206 3593 1212 3594
rect 1390 3598 1396 3599
rect 1390 3594 1391 3598
rect 1395 3594 1396 3598
rect 1390 3593 1396 3594
rect 1574 3598 1580 3599
rect 1574 3594 1575 3598
rect 1579 3594 1580 3598
rect 1574 3593 1580 3594
rect 1766 3598 1772 3599
rect 1766 3594 1767 3598
rect 1771 3594 1772 3598
rect 1766 3593 1772 3594
rect 1934 3598 1940 3599
rect 1934 3594 1935 3598
rect 1939 3594 1940 3598
rect 2358 3594 2364 3595
rect 1934 3593 1940 3594
rect 2030 3593 2036 3594
rect 110 3589 111 3593
rect 115 3589 116 3593
rect 110 3588 116 3589
rect 2030 3589 2031 3593
rect 2035 3589 2036 3593
rect 2358 3590 2359 3594
rect 2363 3590 2364 3594
rect 2030 3588 2036 3589
rect 2070 3589 2076 3590
rect 2358 3589 2364 3590
rect 2582 3594 2588 3595
rect 2582 3590 2583 3594
rect 2587 3590 2588 3594
rect 2582 3589 2588 3590
rect 2798 3594 2804 3595
rect 2798 3590 2799 3594
rect 2803 3590 2804 3594
rect 2798 3589 2804 3590
rect 3006 3594 3012 3595
rect 3006 3590 3007 3594
rect 3011 3590 3012 3594
rect 3006 3589 3012 3590
rect 3214 3594 3220 3595
rect 3214 3590 3215 3594
rect 3219 3590 3220 3594
rect 3214 3589 3220 3590
rect 3430 3594 3436 3595
rect 3430 3590 3431 3594
rect 3435 3590 3436 3594
rect 3430 3589 3436 3590
rect 3990 3589 3996 3590
rect 2070 3585 2071 3589
rect 2075 3585 2076 3589
rect 2070 3584 2076 3585
rect 3990 3585 3991 3589
rect 3995 3585 3996 3589
rect 3990 3584 3996 3585
rect 3182 3583 3188 3584
rect 3182 3579 3183 3583
rect 3187 3582 3188 3583
rect 3502 3583 3508 3584
rect 3502 3582 3503 3583
rect 3187 3580 3503 3582
rect 3187 3579 3188 3580
rect 3182 3578 3188 3579
rect 3502 3579 3503 3580
rect 3507 3579 3508 3583
rect 3502 3578 3508 3579
rect 110 3576 116 3577
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 2030 3576 2036 3577
rect 2030 3572 2031 3576
rect 2035 3572 2036 3576
rect 2030 3571 2036 3572
rect 2070 3572 2076 3573
rect 2070 3568 2071 3572
rect 2075 3568 2076 3572
rect 358 3567 364 3568
rect 358 3566 359 3567
rect 297 3564 359 3566
rect 358 3563 359 3564
rect 363 3563 364 3567
rect 662 3567 668 3568
rect 662 3566 663 3567
rect 569 3564 663 3566
rect 358 3562 364 3563
rect 662 3563 663 3564
rect 667 3563 668 3567
rect 662 3562 668 3563
rect 686 3567 692 3568
rect 686 3563 687 3567
rect 691 3563 692 3567
rect 686 3562 692 3563
rect 1038 3567 1044 3568
rect 1038 3563 1039 3567
rect 1043 3563 1044 3567
rect 1750 3567 1756 3568
rect 1750 3566 1751 3567
rect 1625 3564 1751 3566
rect 1038 3562 1044 3563
rect 1750 3563 1751 3564
rect 1755 3563 1756 3567
rect 1878 3567 1884 3568
rect 1878 3566 1879 3567
rect 1817 3564 1879 3566
rect 1750 3562 1756 3563
rect 1878 3563 1879 3564
rect 1883 3563 1884 3567
rect 2050 3567 2056 3568
rect 2070 3567 2076 3568
rect 3990 3572 3996 3573
rect 3990 3568 3991 3572
rect 3995 3568 3996 3572
rect 3990 3567 3996 3568
rect 2050 3566 2051 3567
rect 1985 3564 2051 3566
rect 1878 3562 1884 3563
rect 2050 3563 2051 3564
rect 2055 3563 2056 3567
rect 2050 3562 2056 3563
rect 2566 3563 2572 3564
rect 2566 3562 2567 3563
rect 2409 3560 2567 3562
rect 2566 3559 2567 3560
rect 2571 3559 2572 3563
rect 2990 3563 2996 3564
rect 2990 3562 2991 3563
rect 2633 3560 2650 3562
rect 2849 3560 2991 3562
rect 2566 3558 2572 3559
rect 2646 3559 2652 3560
rect 246 3557 252 3558
rect 246 3553 247 3557
rect 251 3553 252 3557
rect 246 3552 252 3553
rect 374 3557 380 3558
rect 374 3553 375 3557
rect 379 3553 380 3557
rect 374 3552 380 3553
rect 518 3557 524 3558
rect 518 3553 519 3557
rect 523 3553 524 3557
rect 518 3552 524 3553
rect 678 3557 684 3558
rect 678 3553 679 3557
rect 683 3553 684 3557
rect 678 3552 684 3553
rect 846 3557 852 3558
rect 846 3553 847 3557
rect 851 3553 852 3557
rect 846 3552 852 3553
rect 1022 3557 1028 3558
rect 1022 3553 1023 3557
rect 1027 3553 1028 3557
rect 1022 3552 1028 3553
rect 1206 3557 1212 3558
rect 1206 3553 1207 3557
rect 1211 3553 1212 3557
rect 1206 3552 1212 3553
rect 1390 3557 1396 3558
rect 1390 3553 1391 3557
rect 1395 3553 1396 3557
rect 1390 3552 1396 3553
rect 1574 3557 1580 3558
rect 1574 3553 1575 3557
rect 1579 3553 1580 3557
rect 1574 3552 1580 3553
rect 1766 3557 1772 3558
rect 1766 3553 1767 3557
rect 1771 3553 1772 3557
rect 1766 3552 1772 3553
rect 1934 3557 1940 3558
rect 1934 3553 1935 3557
rect 1939 3553 1940 3557
rect 2646 3555 2647 3559
rect 2651 3555 2652 3559
rect 2990 3559 2991 3560
rect 2995 3559 2996 3563
rect 2990 3558 2996 3559
rect 2646 3554 2652 3555
rect 1934 3552 1940 3553
rect 2358 3553 2364 3554
rect 2358 3549 2359 3553
rect 2363 3549 2364 3553
rect 2358 3548 2364 3549
rect 2582 3553 2588 3554
rect 2582 3549 2583 3553
rect 2587 3549 2588 3553
rect 2582 3548 2588 3549
rect 2798 3553 2804 3554
rect 2798 3549 2799 3553
rect 2803 3549 2804 3553
rect 2798 3548 2804 3549
rect 3006 3553 3012 3554
rect 3006 3549 3007 3553
rect 3011 3549 3012 3553
rect 3006 3548 3012 3549
rect 3214 3553 3220 3554
rect 3214 3549 3215 3553
rect 3219 3549 3220 3553
rect 3214 3548 3220 3549
rect 3430 3553 3436 3554
rect 3430 3549 3431 3553
rect 3435 3549 3436 3553
rect 3430 3548 3436 3549
rect 319 3547 325 3548
rect 319 3543 320 3547
rect 324 3546 325 3547
rect 359 3547 365 3548
rect 359 3546 360 3547
rect 324 3544 360 3546
rect 324 3543 325 3544
rect 319 3542 325 3543
rect 359 3543 360 3544
rect 364 3543 365 3547
rect 359 3542 365 3543
rect 422 3547 428 3548
rect 422 3543 423 3547
rect 427 3546 428 3547
rect 447 3547 453 3548
rect 447 3546 448 3547
rect 427 3544 448 3546
rect 427 3543 428 3544
rect 422 3542 428 3543
rect 447 3543 448 3544
rect 452 3543 453 3547
rect 591 3547 597 3548
rect 591 3546 592 3547
rect 447 3542 453 3543
rect 456 3544 592 3546
rect 358 3539 364 3540
rect 358 3535 359 3539
rect 363 3538 364 3539
rect 456 3538 458 3544
rect 591 3543 592 3544
rect 596 3543 597 3547
rect 591 3542 597 3543
rect 751 3547 757 3548
rect 751 3543 752 3547
rect 756 3546 757 3547
rect 831 3547 837 3548
rect 831 3546 832 3547
rect 756 3544 832 3546
rect 756 3543 757 3544
rect 751 3542 757 3543
rect 831 3543 832 3544
rect 836 3543 837 3547
rect 831 3542 837 3543
rect 919 3547 925 3548
rect 919 3543 920 3547
rect 924 3543 925 3547
rect 919 3542 925 3543
rect 1095 3547 1101 3548
rect 1095 3543 1096 3547
rect 1100 3546 1101 3547
rect 1191 3547 1197 3548
rect 1191 3546 1192 3547
rect 1100 3544 1192 3546
rect 1100 3543 1101 3544
rect 1095 3542 1101 3543
rect 1191 3543 1192 3544
rect 1196 3543 1197 3547
rect 1191 3542 1197 3543
rect 1279 3547 1285 3548
rect 1279 3543 1280 3547
rect 1284 3546 1285 3547
rect 1375 3547 1381 3548
rect 1375 3546 1376 3547
rect 1284 3544 1376 3546
rect 1284 3543 1285 3544
rect 1279 3542 1285 3543
rect 1375 3543 1376 3544
rect 1380 3543 1381 3547
rect 1375 3542 1381 3543
rect 1462 3547 1469 3548
rect 1462 3543 1463 3547
rect 1468 3543 1469 3547
rect 1462 3542 1469 3543
rect 1646 3547 1653 3548
rect 1646 3543 1647 3547
rect 1652 3543 1653 3547
rect 1646 3542 1653 3543
rect 1750 3547 1756 3548
rect 1750 3543 1751 3547
rect 1755 3546 1756 3547
rect 1839 3547 1845 3548
rect 1839 3546 1840 3547
rect 1755 3544 1840 3546
rect 1755 3543 1756 3544
rect 1750 3542 1756 3543
rect 1839 3543 1840 3544
rect 1844 3543 1845 3547
rect 1839 3542 1845 3543
rect 1878 3547 1884 3548
rect 1878 3543 1879 3547
rect 1883 3546 1884 3547
rect 2007 3547 2013 3548
rect 2007 3546 2008 3547
rect 1883 3544 2008 3546
rect 1883 3543 1884 3544
rect 1878 3542 1884 3543
rect 2007 3543 2008 3544
rect 2012 3543 2013 3547
rect 2007 3542 2013 3543
rect 2430 3543 2437 3544
rect 363 3536 458 3538
rect 662 3539 668 3540
rect 363 3535 364 3536
rect 358 3534 364 3535
rect 662 3535 663 3539
rect 667 3538 668 3539
rect 921 3538 923 3542
rect 2430 3539 2431 3543
rect 2436 3539 2437 3543
rect 2430 3538 2437 3539
rect 2566 3543 2572 3544
rect 2566 3539 2567 3543
rect 2571 3542 2572 3543
rect 2655 3543 2661 3544
rect 2655 3542 2656 3543
rect 2571 3540 2656 3542
rect 2571 3539 2572 3540
rect 2566 3538 2572 3539
rect 2655 3539 2656 3540
rect 2660 3539 2661 3543
rect 2655 3538 2661 3539
rect 2871 3543 2877 3544
rect 2871 3539 2872 3543
rect 2876 3542 2877 3543
rect 2991 3543 2997 3544
rect 2991 3542 2992 3543
rect 2876 3540 2992 3542
rect 2876 3539 2877 3540
rect 2871 3538 2877 3539
rect 2991 3539 2992 3540
rect 2996 3539 2997 3543
rect 2991 3538 2997 3539
rect 3079 3543 3085 3544
rect 3079 3539 3080 3543
rect 3084 3542 3085 3543
rect 3199 3543 3205 3544
rect 3199 3542 3200 3543
rect 3084 3540 3200 3542
rect 3084 3539 3085 3540
rect 3079 3538 3085 3539
rect 3199 3539 3200 3540
rect 3204 3539 3205 3543
rect 3199 3538 3205 3539
rect 3287 3543 3293 3544
rect 3287 3539 3288 3543
rect 3292 3542 3293 3543
rect 3415 3543 3421 3544
rect 3415 3542 3416 3543
rect 3292 3540 3416 3542
rect 3292 3539 3293 3540
rect 3287 3538 3293 3539
rect 3415 3539 3416 3540
rect 3420 3539 3421 3543
rect 3415 3538 3421 3539
rect 3502 3543 3509 3544
rect 3502 3539 3503 3543
rect 3508 3539 3509 3543
rect 3502 3538 3509 3539
rect 667 3536 923 3538
rect 667 3535 668 3536
rect 662 3534 668 3535
rect 2990 3535 2996 3536
rect 230 3531 236 3532
rect 230 3527 231 3531
rect 235 3530 236 3531
rect 950 3531 956 3532
rect 235 3528 682 3530
rect 235 3527 236 3528
rect 230 3526 236 3527
rect 223 3523 229 3524
rect 223 3519 224 3523
rect 228 3522 229 3523
rect 247 3523 253 3524
rect 247 3522 248 3523
rect 228 3520 248 3522
rect 228 3519 229 3520
rect 223 3518 229 3519
rect 247 3519 248 3520
rect 252 3519 253 3523
rect 247 3518 253 3519
rect 335 3523 341 3524
rect 335 3519 336 3523
rect 340 3522 341 3523
rect 414 3523 420 3524
rect 414 3522 415 3523
rect 340 3520 415 3522
rect 340 3519 341 3520
rect 335 3518 341 3519
rect 414 3519 415 3520
rect 419 3519 420 3523
rect 414 3518 420 3519
rect 471 3523 477 3524
rect 471 3519 472 3523
rect 476 3522 477 3523
rect 527 3523 533 3524
rect 527 3522 528 3523
rect 476 3520 528 3522
rect 476 3519 477 3520
rect 471 3518 477 3519
rect 527 3519 528 3520
rect 532 3519 533 3523
rect 527 3518 533 3519
rect 615 3523 621 3524
rect 615 3519 616 3523
rect 620 3522 621 3523
rect 671 3523 677 3524
rect 671 3522 672 3523
rect 620 3520 672 3522
rect 620 3519 621 3520
rect 615 3518 621 3519
rect 671 3519 672 3520
rect 676 3519 677 3523
rect 680 3522 682 3528
rect 950 3527 951 3531
rect 955 3530 956 3531
rect 1566 3531 1572 3532
rect 955 3528 1161 3530
rect 955 3527 956 3528
rect 950 3526 956 3527
rect 759 3523 765 3524
rect 759 3522 760 3523
rect 680 3520 760 3522
rect 671 3518 677 3519
rect 759 3519 760 3520
rect 764 3519 765 3523
rect 759 3518 765 3519
rect 903 3523 909 3524
rect 903 3519 904 3523
rect 908 3522 909 3523
rect 951 3523 957 3524
rect 951 3522 952 3523
rect 908 3520 952 3522
rect 908 3519 909 3520
rect 903 3518 909 3519
rect 951 3519 952 3520
rect 956 3519 957 3523
rect 951 3518 957 3519
rect 1038 3523 1045 3524
rect 1038 3519 1039 3523
rect 1044 3519 1045 3523
rect 1159 3522 1161 3528
rect 1566 3527 1567 3531
rect 1571 3530 1572 3531
rect 2990 3531 2991 3535
rect 2995 3534 2996 3535
rect 2995 3532 3322 3534
rect 2995 3531 2996 3532
rect 2990 3530 2996 3531
rect 1571 3528 1706 3530
rect 1571 3527 1572 3528
rect 1566 3526 1572 3527
rect 1167 3523 1173 3524
rect 1167 3522 1168 3523
rect 1159 3520 1168 3522
rect 1038 3518 1045 3519
rect 1167 3519 1168 3520
rect 1172 3519 1173 3523
rect 1295 3523 1301 3524
rect 1295 3522 1296 3523
rect 1167 3518 1173 3519
rect 1177 3520 1296 3522
rect 150 3515 156 3516
rect 150 3511 151 3515
rect 155 3511 156 3515
rect 150 3510 156 3511
rect 262 3515 268 3516
rect 262 3511 263 3515
rect 267 3511 268 3515
rect 262 3510 268 3511
rect 398 3515 404 3516
rect 398 3511 399 3515
rect 403 3511 404 3515
rect 398 3510 404 3511
rect 542 3515 548 3516
rect 542 3511 543 3515
rect 547 3511 548 3515
rect 542 3510 548 3511
rect 686 3515 692 3516
rect 686 3511 687 3515
rect 691 3511 692 3515
rect 686 3510 692 3511
rect 830 3515 836 3516
rect 830 3511 831 3515
rect 835 3511 836 3515
rect 830 3510 836 3511
rect 966 3515 972 3516
rect 966 3511 967 3515
rect 971 3511 972 3515
rect 966 3510 972 3511
rect 1094 3515 1100 3516
rect 1094 3511 1095 3515
rect 1099 3511 1100 3515
rect 1094 3510 1100 3511
rect 230 3507 236 3508
rect 230 3506 231 3507
rect 201 3504 231 3506
rect 230 3503 231 3504
rect 235 3503 236 3507
rect 950 3507 956 3508
rect 950 3506 951 3507
rect 881 3504 951 3506
rect 230 3502 236 3503
rect 422 3503 428 3504
rect 422 3499 423 3503
rect 427 3499 428 3503
rect 950 3503 951 3504
rect 955 3503 956 3507
rect 1177 3506 1179 3520
rect 1295 3519 1296 3520
rect 1300 3519 1301 3523
rect 1415 3523 1421 3524
rect 1415 3522 1416 3523
rect 1295 3518 1301 3519
rect 1313 3520 1416 3522
rect 1222 3515 1228 3516
rect 1222 3511 1223 3515
rect 1227 3511 1228 3515
rect 1222 3510 1228 3511
rect 1313 3506 1315 3520
rect 1415 3519 1416 3520
rect 1420 3519 1421 3523
rect 1415 3518 1421 3519
rect 1534 3523 1541 3524
rect 1534 3519 1535 3523
rect 1540 3519 1541 3523
rect 1534 3518 1541 3519
rect 1655 3523 1661 3524
rect 1655 3519 1656 3523
rect 1660 3522 1661 3523
rect 1695 3523 1701 3524
rect 1695 3522 1696 3523
rect 1660 3520 1696 3522
rect 1660 3519 1661 3520
rect 1655 3518 1661 3519
rect 1695 3519 1696 3520
rect 1700 3519 1701 3523
rect 1704 3522 1706 3528
rect 2511 3527 2517 3528
rect 1783 3523 1789 3524
rect 1783 3522 1784 3523
rect 1704 3520 1784 3522
rect 1695 3518 1701 3519
rect 1783 3519 1784 3520
rect 1788 3519 1789 3523
rect 2511 3523 2512 3527
rect 2516 3526 2517 3527
rect 2559 3527 2565 3528
rect 2559 3526 2560 3527
rect 2516 3524 2560 3526
rect 2516 3523 2517 3524
rect 2511 3522 2517 3523
rect 2559 3523 2560 3524
rect 2564 3523 2565 3527
rect 2559 3522 2565 3523
rect 2646 3527 2653 3528
rect 2646 3523 2647 3527
rect 2652 3523 2653 3527
rect 2646 3522 2653 3523
rect 2775 3527 2781 3528
rect 2775 3523 2776 3527
rect 2780 3526 2781 3527
rect 2815 3527 2821 3528
rect 2815 3526 2816 3527
rect 2780 3524 2816 3526
rect 2780 3523 2781 3524
rect 2775 3522 2781 3523
rect 2815 3523 2816 3524
rect 2820 3523 2821 3527
rect 2815 3522 2821 3523
rect 2903 3527 2909 3528
rect 2903 3523 2904 3527
rect 2908 3526 2909 3527
rect 2935 3527 2941 3528
rect 2935 3526 2936 3527
rect 2908 3524 2936 3526
rect 2908 3523 2909 3524
rect 2903 3522 2909 3523
rect 2935 3523 2936 3524
rect 2940 3523 2941 3527
rect 2935 3522 2941 3523
rect 3023 3527 3029 3528
rect 3023 3523 3024 3527
rect 3028 3526 3029 3527
rect 3055 3527 3061 3528
rect 3055 3526 3056 3527
rect 3028 3524 3056 3526
rect 3028 3523 3029 3524
rect 3023 3522 3029 3523
rect 3055 3523 3056 3524
rect 3060 3523 3061 3527
rect 3055 3522 3061 3523
rect 3143 3527 3149 3528
rect 3143 3523 3144 3527
rect 3148 3526 3149 3527
rect 3183 3527 3189 3528
rect 3183 3526 3184 3527
rect 3148 3524 3184 3526
rect 3148 3523 3149 3524
rect 3143 3522 3149 3523
rect 3183 3523 3184 3524
rect 3188 3523 3189 3527
rect 3183 3522 3189 3523
rect 3271 3527 3277 3528
rect 3271 3523 3272 3527
rect 3276 3526 3277 3527
rect 3311 3527 3317 3528
rect 3311 3526 3312 3527
rect 3276 3524 3312 3526
rect 3276 3523 3277 3524
rect 3271 3522 3277 3523
rect 3311 3523 3312 3524
rect 3316 3523 3317 3527
rect 3320 3526 3322 3532
rect 3399 3527 3405 3528
rect 3399 3526 3400 3527
rect 3320 3524 3400 3526
rect 3311 3522 3317 3523
rect 3399 3523 3400 3524
rect 3404 3523 3405 3527
rect 3399 3522 3405 3523
rect 1783 3518 1789 3519
rect 2438 3519 2444 3520
rect 1342 3515 1348 3516
rect 1342 3511 1343 3515
rect 1347 3511 1348 3515
rect 1342 3510 1348 3511
rect 1462 3515 1468 3516
rect 1462 3511 1463 3515
rect 1467 3511 1468 3515
rect 1462 3510 1468 3511
rect 1582 3515 1588 3516
rect 1582 3511 1583 3515
rect 1587 3511 1588 3515
rect 1582 3510 1588 3511
rect 1710 3515 1716 3516
rect 1710 3511 1711 3515
rect 1715 3511 1716 3515
rect 2438 3515 2439 3519
rect 2443 3515 2444 3519
rect 2438 3514 2444 3515
rect 2574 3519 2580 3520
rect 2574 3515 2575 3519
rect 2579 3515 2580 3519
rect 2574 3514 2580 3515
rect 2702 3519 2708 3520
rect 2702 3515 2703 3519
rect 2707 3515 2708 3519
rect 2702 3514 2708 3515
rect 2830 3519 2836 3520
rect 2830 3515 2831 3519
rect 2835 3515 2836 3519
rect 2830 3514 2836 3515
rect 2950 3519 2956 3520
rect 2950 3515 2951 3519
rect 2955 3515 2956 3519
rect 2950 3514 2956 3515
rect 3070 3519 3076 3520
rect 3070 3515 3071 3519
rect 3075 3515 3076 3519
rect 3070 3514 3076 3515
rect 3198 3519 3204 3520
rect 3198 3515 3199 3519
rect 3203 3515 3204 3519
rect 3198 3514 3204 3515
rect 3326 3519 3332 3520
rect 3326 3515 3327 3519
rect 3331 3515 3332 3519
rect 3326 3514 3332 3515
rect 1710 3510 1716 3511
rect 2786 3511 2792 3512
rect 2786 3510 2787 3511
rect 2753 3508 2787 3510
rect 1446 3507 1452 3508
rect 1446 3506 1447 3507
rect 1145 3504 1179 3506
rect 1273 3504 1315 3506
rect 1393 3504 1447 3506
rect 950 3502 956 3503
rect 1446 3503 1447 3504
rect 1451 3503 1452 3507
rect 1566 3507 1572 3508
rect 1566 3506 1567 3507
rect 1513 3504 1567 3506
rect 1446 3502 1452 3503
rect 1566 3503 1567 3504
rect 1571 3503 1572 3507
rect 1646 3507 1652 3508
rect 1646 3506 1647 3507
rect 1633 3504 1647 3506
rect 1566 3502 1572 3503
rect 1646 3503 1647 3504
rect 1651 3503 1652 3507
rect 1646 3502 1652 3503
rect 2430 3507 2436 3508
rect 2430 3503 2431 3507
rect 2435 3503 2436 3507
rect 2786 3507 2787 3508
rect 2791 3507 2792 3511
rect 2786 3506 2792 3507
rect 2430 3502 2436 3503
rect 422 3498 428 3499
rect 2070 3500 2076 3501
rect 110 3496 116 3497
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 110 3491 116 3492
rect 2030 3496 2036 3497
rect 2030 3492 2031 3496
rect 2035 3492 2036 3496
rect 2070 3496 2071 3500
rect 2075 3496 2076 3500
rect 2070 3495 2076 3496
rect 3990 3500 3996 3501
rect 3990 3496 3991 3500
rect 3995 3496 3996 3500
rect 3990 3495 3996 3496
rect 2030 3491 2036 3492
rect 2070 3483 2076 3484
rect 110 3479 116 3480
rect 110 3475 111 3479
rect 115 3475 116 3479
rect 2030 3479 2036 3480
rect 2030 3475 2031 3479
rect 2035 3475 2036 3479
rect 2070 3479 2071 3483
rect 2075 3479 2076 3483
rect 3990 3483 3996 3484
rect 3990 3479 3991 3483
rect 3995 3479 3996 3483
rect 2070 3478 2076 3479
rect 2438 3478 2444 3479
rect 110 3474 116 3475
rect 150 3474 156 3475
rect 150 3470 151 3474
rect 155 3470 156 3474
rect 150 3469 156 3470
rect 262 3474 268 3475
rect 262 3470 263 3474
rect 267 3470 268 3474
rect 262 3469 268 3470
rect 398 3474 404 3475
rect 398 3470 399 3474
rect 403 3470 404 3474
rect 398 3469 404 3470
rect 542 3474 548 3475
rect 542 3470 543 3474
rect 547 3470 548 3474
rect 542 3469 548 3470
rect 686 3474 692 3475
rect 686 3470 687 3474
rect 691 3470 692 3474
rect 686 3469 692 3470
rect 830 3474 836 3475
rect 830 3470 831 3474
rect 835 3470 836 3474
rect 830 3469 836 3470
rect 966 3474 972 3475
rect 966 3470 967 3474
rect 971 3470 972 3474
rect 966 3469 972 3470
rect 1094 3474 1100 3475
rect 1094 3470 1095 3474
rect 1099 3470 1100 3474
rect 1094 3469 1100 3470
rect 1222 3474 1228 3475
rect 1222 3470 1223 3474
rect 1227 3470 1228 3474
rect 1222 3469 1228 3470
rect 1342 3474 1348 3475
rect 1342 3470 1343 3474
rect 1347 3470 1348 3474
rect 1342 3469 1348 3470
rect 1462 3474 1468 3475
rect 1462 3470 1463 3474
rect 1467 3470 1468 3474
rect 1462 3469 1468 3470
rect 1582 3474 1588 3475
rect 1582 3470 1583 3474
rect 1587 3470 1588 3474
rect 1582 3469 1588 3470
rect 1710 3474 1716 3475
rect 2030 3474 2036 3475
rect 2438 3474 2439 3478
rect 2443 3474 2444 3478
rect 1710 3470 1711 3474
rect 1715 3470 1716 3474
rect 2438 3473 2444 3474
rect 2574 3478 2580 3479
rect 2574 3474 2575 3478
rect 2579 3474 2580 3478
rect 2574 3473 2580 3474
rect 2702 3478 2708 3479
rect 2702 3474 2703 3478
rect 2707 3474 2708 3478
rect 2702 3473 2708 3474
rect 2830 3478 2836 3479
rect 2830 3474 2831 3478
rect 2835 3474 2836 3478
rect 2830 3473 2836 3474
rect 2950 3478 2956 3479
rect 2950 3474 2951 3478
rect 2955 3474 2956 3478
rect 2950 3473 2956 3474
rect 3070 3478 3076 3479
rect 3070 3474 3071 3478
rect 3075 3474 3076 3478
rect 3070 3473 3076 3474
rect 3198 3478 3204 3479
rect 3198 3474 3199 3478
rect 3203 3474 3204 3478
rect 3198 3473 3204 3474
rect 3326 3478 3332 3479
rect 3990 3478 3996 3479
rect 3326 3474 3327 3478
rect 3331 3474 3332 3478
rect 3326 3473 3332 3474
rect 1710 3469 1716 3470
rect 2358 3446 2364 3447
rect 150 3442 156 3443
rect 150 3438 151 3442
rect 155 3438 156 3442
rect 110 3437 116 3438
rect 150 3437 156 3438
rect 422 3442 428 3443
rect 422 3438 423 3442
rect 427 3438 428 3442
rect 422 3437 428 3438
rect 742 3442 748 3443
rect 742 3438 743 3442
rect 747 3438 748 3442
rect 742 3437 748 3438
rect 1070 3442 1076 3443
rect 1070 3438 1071 3442
rect 1075 3438 1076 3442
rect 1070 3437 1076 3438
rect 1398 3442 1404 3443
rect 2358 3442 2359 3446
rect 2363 3442 2364 3446
rect 1398 3438 1399 3442
rect 1403 3438 1404 3442
rect 2070 3441 2076 3442
rect 2358 3441 2364 3442
rect 2462 3446 2468 3447
rect 2462 3442 2463 3446
rect 2467 3442 2468 3446
rect 2462 3441 2468 3442
rect 2566 3446 2572 3447
rect 2566 3442 2567 3446
rect 2571 3442 2572 3446
rect 2566 3441 2572 3442
rect 2670 3446 2676 3447
rect 2670 3442 2671 3446
rect 2675 3442 2676 3446
rect 2670 3441 2676 3442
rect 2774 3446 2780 3447
rect 2774 3442 2775 3446
rect 2779 3442 2780 3446
rect 2774 3441 2780 3442
rect 2878 3446 2884 3447
rect 2878 3442 2879 3446
rect 2883 3442 2884 3446
rect 2878 3441 2884 3442
rect 2982 3446 2988 3447
rect 2982 3442 2983 3446
rect 2987 3442 2988 3446
rect 2982 3441 2988 3442
rect 3086 3446 3092 3447
rect 3086 3442 3087 3446
rect 3091 3442 3092 3446
rect 3086 3441 3092 3442
rect 3190 3446 3196 3447
rect 3190 3442 3191 3446
rect 3195 3442 3196 3446
rect 3190 3441 3196 3442
rect 3990 3441 3996 3442
rect 1398 3437 1404 3438
rect 2030 3437 2036 3438
rect 110 3433 111 3437
rect 115 3433 116 3437
rect 110 3432 116 3433
rect 2030 3433 2031 3437
rect 2035 3433 2036 3437
rect 2070 3437 2071 3441
rect 2075 3437 2076 3441
rect 2070 3436 2076 3437
rect 3990 3437 3991 3441
rect 3995 3437 3996 3441
rect 3990 3436 3996 3437
rect 2030 3432 2036 3433
rect 2070 3424 2076 3425
rect 110 3420 116 3421
rect 110 3416 111 3420
rect 115 3416 116 3420
rect 110 3415 116 3416
rect 2030 3420 2036 3421
rect 2030 3416 2031 3420
rect 2035 3416 2036 3420
rect 2070 3420 2071 3424
rect 2075 3420 2076 3424
rect 2070 3419 2076 3420
rect 3990 3424 3996 3425
rect 3990 3420 3991 3424
rect 3995 3420 3996 3424
rect 3990 3419 3996 3420
rect 2030 3415 2036 3416
rect 2446 3415 2452 3416
rect 2446 3414 2447 3415
rect 2409 3412 2447 3414
rect 406 3411 412 3412
rect 406 3410 407 3411
rect 201 3408 407 3410
rect 406 3407 407 3408
rect 411 3407 412 3411
rect 406 3406 412 3407
rect 414 3411 420 3412
rect 414 3407 415 3411
rect 419 3407 420 3411
rect 1534 3411 1540 3412
rect 1534 3410 1535 3411
rect 1449 3408 1535 3410
rect 414 3406 420 3407
rect 1534 3407 1535 3408
rect 1539 3407 1540 3411
rect 2446 3411 2447 3412
rect 2451 3411 2452 3415
rect 2446 3410 2452 3411
rect 2486 3415 2492 3416
rect 2486 3411 2487 3415
rect 2491 3411 2492 3415
rect 2638 3415 2644 3416
rect 2638 3414 2639 3415
rect 2617 3412 2639 3414
rect 2486 3410 2492 3411
rect 2638 3411 2639 3412
rect 2643 3411 2644 3415
rect 2638 3410 2644 3411
rect 1534 3406 1540 3407
rect 2358 3405 2364 3406
rect 150 3401 156 3402
rect 150 3397 151 3401
rect 155 3397 156 3401
rect 150 3396 156 3397
rect 422 3401 428 3402
rect 422 3397 423 3401
rect 427 3397 428 3401
rect 422 3396 428 3397
rect 742 3401 748 3402
rect 742 3397 743 3401
rect 747 3397 748 3401
rect 742 3396 748 3397
rect 1070 3401 1076 3402
rect 1070 3397 1071 3401
rect 1075 3397 1076 3401
rect 1070 3396 1076 3397
rect 1398 3401 1404 3402
rect 1398 3397 1399 3401
rect 1403 3397 1404 3401
rect 2358 3401 2359 3405
rect 2363 3401 2364 3405
rect 2358 3400 2364 3401
rect 2462 3405 2468 3406
rect 2462 3401 2463 3405
rect 2467 3401 2468 3405
rect 2462 3400 2468 3401
rect 2566 3405 2572 3406
rect 2566 3401 2567 3405
rect 2571 3401 2572 3405
rect 2566 3400 2572 3401
rect 2670 3405 2676 3406
rect 2670 3401 2671 3405
rect 2675 3401 2676 3405
rect 2670 3400 2676 3401
rect 2774 3405 2780 3406
rect 2774 3401 2775 3405
rect 2779 3401 2780 3405
rect 2774 3400 2780 3401
rect 2878 3405 2884 3406
rect 2878 3401 2879 3405
rect 2883 3401 2884 3405
rect 2878 3400 2884 3401
rect 2982 3405 2988 3406
rect 2982 3401 2983 3405
rect 2987 3401 2988 3405
rect 2982 3400 2988 3401
rect 3086 3405 3092 3406
rect 3086 3401 3087 3405
rect 3091 3401 3092 3405
rect 3086 3400 3092 3401
rect 3190 3405 3196 3406
rect 3190 3401 3191 3405
rect 3195 3401 3196 3405
rect 3190 3400 3196 3401
rect 1398 3396 1404 3397
rect 2430 3395 2437 3396
rect 214 3391 220 3392
rect 214 3387 215 3391
rect 219 3390 220 3391
rect 223 3391 229 3392
rect 223 3390 224 3391
rect 219 3388 224 3390
rect 219 3387 220 3388
rect 214 3386 220 3387
rect 223 3387 224 3388
rect 228 3387 229 3391
rect 223 3386 229 3387
rect 495 3391 501 3392
rect 495 3387 496 3391
rect 500 3390 501 3391
rect 727 3391 733 3392
rect 727 3390 728 3391
rect 500 3388 728 3390
rect 500 3387 501 3388
rect 495 3386 501 3387
rect 727 3387 728 3388
rect 732 3387 733 3391
rect 727 3386 733 3387
rect 815 3391 821 3392
rect 815 3387 816 3391
rect 820 3390 821 3391
rect 1055 3391 1061 3392
rect 1055 3390 1056 3391
rect 820 3388 1056 3390
rect 820 3387 821 3388
rect 815 3386 821 3387
rect 1055 3387 1056 3388
rect 1060 3387 1061 3391
rect 1143 3391 1149 3392
rect 1143 3390 1144 3391
rect 1055 3386 1061 3387
rect 1064 3388 1144 3390
rect 406 3383 412 3384
rect 406 3379 407 3383
rect 411 3382 412 3383
rect 1064 3382 1066 3388
rect 1143 3387 1144 3388
rect 1148 3387 1149 3391
rect 1143 3386 1149 3387
rect 1446 3391 1452 3392
rect 1446 3387 1447 3391
rect 1451 3390 1452 3391
rect 1471 3391 1477 3392
rect 1471 3390 1472 3391
rect 1451 3388 1472 3390
rect 1451 3387 1452 3388
rect 1446 3386 1452 3387
rect 1471 3387 1472 3388
rect 1476 3387 1477 3391
rect 2430 3391 2431 3395
rect 2436 3391 2437 3395
rect 2430 3390 2437 3391
rect 2446 3395 2452 3396
rect 2446 3391 2447 3395
rect 2451 3394 2452 3395
rect 2535 3395 2541 3396
rect 2535 3394 2536 3395
rect 2451 3392 2536 3394
rect 2451 3391 2452 3392
rect 2446 3390 2452 3391
rect 2535 3391 2536 3392
rect 2540 3391 2541 3395
rect 2535 3390 2541 3391
rect 2639 3395 2645 3396
rect 2639 3391 2640 3395
rect 2644 3394 2645 3395
rect 2655 3395 2661 3396
rect 2655 3394 2656 3395
rect 2644 3392 2656 3394
rect 2644 3391 2645 3392
rect 2639 3390 2645 3391
rect 2655 3391 2656 3392
rect 2660 3391 2661 3395
rect 2655 3390 2661 3391
rect 2743 3395 2749 3396
rect 2743 3391 2744 3395
rect 2748 3394 2749 3395
rect 2759 3395 2765 3396
rect 2759 3394 2760 3395
rect 2748 3392 2760 3394
rect 2748 3391 2749 3392
rect 2743 3390 2749 3391
rect 2759 3391 2760 3392
rect 2764 3391 2765 3395
rect 2759 3390 2765 3391
rect 2847 3395 2853 3396
rect 2847 3391 2848 3395
rect 2852 3394 2853 3395
rect 2863 3395 2869 3396
rect 2863 3394 2864 3395
rect 2852 3392 2864 3394
rect 2852 3391 2853 3392
rect 2847 3390 2853 3391
rect 2863 3391 2864 3392
rect 2868 3391 2869 3395
rect 2863 3390 2869 3391
rect 2951 3395 2957 3396
rect 2951 3391 2952 3395
rect 2956 3394 2957 3395
rect 2967 3395 2973 3396
rect 2967 3394 2968 3395
rect 2956 3392 2968 3394
rect 2956 3391 2957 3392
rect 2951 3390 2957 3391
rect 2967 3391 2968 3392
rect 2972 3391 2973 3395
rect 2967 3390 2973 3391
rect 3055 3395 3061 3396
rect 3055 3391 3056 3395
rect 3060 3394 3061 3395
rect 3071 3395 3077 3396
rect 3071 3394 3072 3395
rect 3060 3392 3072 3394
rect 3060 3391 3061 3392
rect 3055 3390 3061 3391
rect 3071 3391 3072 3392
rect 3076 3391 3077 3395
rect 3071 3390 3077 3391
rect 3159 3395 3165 3396
rect 3159 3391 3160 3395
rect 3164 3394 3165 3395
rect 3175 3395 3181 3396
rect 3175 3394 3176 3395
rect 3164 3392 3176 3394
rect 3164 3391 3165 3392
rect 3159 3390 3165 3391
rect 3175 3391 3176 3392
rect 3180 3391 3181 3395
rect 3263 3395 3269 3396
rect 3263 3394 3264 3395
rect 3175 3390 3181 3391
rect 3184 3392 3264 3394
rect 1471 3386 1477 3387
rect 2786 3387 2792 3388
rect 2786 3383 2787 3387
rect 2791 3386 2792 3387
rect 3184 3386 3186 3392
rect 3263 3391 3264 3392
rect 3268 3391 3269 3395
rect 3263 3390 3269 3391
rect 2791 3384 3186 3386
rect 2791 3383 2792 3384
rect 2786 3382 2792 3383
rect 411 3380 1066 3382
rect 411 3379 412 3380
rect 406 3378 412 3379
rect 2838 3363 2844 3364
rect 2838 3359 2839 3363
rect 2843 3362 2844 3363
rect 2843 3360 2954 3362
rect 2843 3359 2844 3360
rect 2838 3358 2844 3359
rect 223 3355 229 3356
rect 223 3351 224 3355
rect 228 3354 229 3355
rect 303 3355 309 3356
rect 303 3354 304 3355
rect 228 3352 304 3354
rect 228 3351 229 3352
rect 223 3350 229 3351
rect 303 3351 304 3352
rect 308 3351 309 3355
rect 303 3350 309 3351
rect 391 3355 397 3356
rect 391 3351 392 3355
rect 396 3354 397 3355
rect 511 3355 517 3356
rect 511 3354 512 3355
rect 396 3352 512 3354
rect 396 3351 397 3352
rect 391 3350 397 3351
rect 511 3351 512 3352
rect 516 3351 517 3355
rect 511 3350 517 3351
rect 599 3355 605 3356
rect 599 3351 600 3355
rect 604 3354 605 3355
rect 727 3355 733 3356
rect 727 3354 728 3355
rect 604 3352 728 3354
rect 604 3351 605 3352
rect 599 3350 605 3351
rect 727 3351 728 3352
rect 732 3351 733 3355
rect 727 3350 733 3351
rect 815 3355 821 3356
rect 815 3351 816 3355
rect 820 3354 821 3355
rect 943 3355 949 3356
rect 943 3354 944 3355
rect 820 3352 944 3354
rect 820 3351 821 3352
rect 815 3350 821 3351
rect 943 3351 944 3352
rect 948 3351 949 3355
rect 943 3350 949 3351
rect 994 3355 1000 3356
rect 994 3351 995 3355
rect 999 3354 1000 3355
rect 1031 3355 1037 3356
rect 1031 3354 1032 3355
rect 999 3352 1032 3354
rect 999 3351 1000 3352
rect 994 3350 1000 3351
rect 1031 3351 1032 3352
rect 1036 3351 1037 3355
rect 1031 3350 1037 3351
rect 1239 3355 1245 3356
rect 1239 3351 1240 3355
rect 1244 3354 1245 3355
rect 1351 3355 1357 3356
rect 1351 3354 1352 3355
rect 1244 3352 1352 3354
rect 1244 3351 1245 3352
rect 1239 3350 1245 3351
rect 1351 3351 1352 3352
rect 1356 3351 1357 3355
rect 1351 3350 1357 3351
rect 1439 3355 1445 3356
rect 1439 3351 1440 3355
rect 1444 3354 1445 3355
rect 1543 3355 1549 3356
rect 1543 3354 1544 3355
rect 1444 3352 1544 3354
rect 1444 3351 1445 3352
rect 1439 3350 1445 3351
rect 1543 3351 1544 3352
rect 1548 3351 1549 3355
rect 1543 3350 1549 3351
rect 1631 3355 1637 3356
rect 1631 3351 1632 3355
rect 1636 3354 1637 3355
rect 1735 3355 1741 3356
rect 1735 3354 1736 3355
rect 1636 3352 1736 3354
rect 1636 3351 1637 3352
rect 1631 3350 1637 3351
rect 1735 3351 1736 3352
rect 1740 3351 1741 3355
rect 1735 3350 1741 3351
rect 1823 3355 1829 3356
rect 1823 3351 1824 3355
rect 1828 3354 1829 3355
rect 1919 3355 1925 3356
rect 1919 3354 1920 3355
rect 1828 3352 1920 3354
rect 1828 3351 1829 3352
rect 1823 3350 1829 3351
rect 1919 3351 1920 3352
rect 1924 3351 1925 3355
rect 1919 3350 1925 3351
rect 2002 3355 2013 3356
rect 2002 3351 2003 3355
rect 2007 3351 2008 3355
rect 2012 3351 2013 3355
rect 2002 3350 2013 3351
rect 2486 3355 2492 3356
rect 2486 3351 2487 3355
rect 2491 3354 2492 3355
rect 2511 3355 2517 3356
rect 2511 3354 2512 3355
rect 2491 3352 2512 3354
rect 2491 3351 2492 3352
rect 2486 3350 2492 3351
rect 2511 3351 2512 3352
rect 2516 3351 2517 3355
rect 2615 3355 2621 3356
rect 2615 3354 2616 3355
rect 2511 3350 2517 3351
rect 2524 3352 2616 3354
rect 150 3347 156 3348
rect 150 3343 151 3347
rect 155 3343 156 3347
rect 150 3342 156 3343
rect 318 3347 324 3348
rect 318 3343 319 3347
rect 323 3343 324 3347
rect 318 3342 324 3343
rect 526 3347 532 3348
rect 526 3343 527 3347
rect 531 3343 532 3347
rect 526 3342 532 3343
rect 742 3347 748 3348
rect 742 3343 743 3347
rect 747 3343 748 3347
rect 742 3342 748 3343
rect 958 3347 964 3348
rect 958 3343 959 3347
rect 963 3343 964 3347
rect 958 3342 964 3343
rect 1166 3347 1172 3348
rect 1166 3343 1167 3347
rect 1171 3343 1172 3347
rect 1166 3342 1172 3343
rect 1366 3347 1372 3348
rect 1366 3343 1367 3347
rect 1371 3343 1372 3347
rect 1366 3342 1372 3343
rect 1558 3347 1564 3348
rect 1558 3343 1559 3347
rect 1563 3343 1564 3347
rect 1558 3342 1564 3343
rect 1750 3347 1756 3348
rect 1750 3343 1751 3347
rect 1755 3343 1756 3347
rect 1750 3342 1756 3343
rect 1934 3347 1940 3348
rect 1934 3343 1935 3347
rect 1939 3343 1940 3347
rect 1934 3342 1940 3343
rect 2438 3347 2444 3348
rect 2438 3343 2439 3347
rect 2443 3343 2444 3347
rect 2438 3342 2444 3343
rect 214 3339 220 3340
rect 214 3338 215 3339
rect 201 3336 215 3338
rect 214 3335 215 3336
rect 219 3335 220 3339
rect 1335 3339 1341 3340
rect 1335 3338 1336 3339
rect 1217 3336 1336 3338
rect 214 3334 220 3335
rect 1335 3335 1336 3336
rect 1340 3335 1341 3339
rect 2524 3338 2526 3352
rect 2615 3351 2616 3352
rect 2620 3351 2621 3355
rect 2615 3350 2621 3351
rect 2638 3355 2644 3356
rect 2638 3351 2639 3355
rect 2643 3354 2644 3355
rect 2719 3355 2725 3356
rect 2719 3354 2720 3355
rect 2643 3352 2720 3354
rect 2643 3351 2644 3352
rect 2638 3350 2644 3351
rect 2719 3351 2720 3352
rect 2724 3351 2725 3355
rect 2823 3355 2829 3356
rect 2823 3354 2824 3355
rect 2719 3350 2725 3351
rect 2732 3352 2824 3354
rect 2542 3347 2548 3348
rect 2542 3343 2543 3347
rect 2547 3343 2548 3347
rect 2542 3342 2548 3343
rect 2646 3347 2652 3348
rect 2646 3343 2647 3347
rect 2651 3343 2652 3347
rect 2646 3342 2652 3343
rect 2606 3339 2612 3340
rect 2606 3338 2607 3339
rect 2489 3336 2526 3338
rect 2593 3336 2607 3338
rect 1335 3334 1341 3335
rect 2606 3335 2607 3336
rect 2611 3335 2612 3339
rect 2732 3338 2734 3352
rect 2823 3351 2824 3352
rect 2828 3351 2829 3355
rect 2823 3350 2829 3351
rect 2927 3355 2933 3356
rect 2927 3351 2928 3355
rect 2932 3354 2933 3355
rect 2943 3355 2949 3356
rect 2943 3354 2944 3355
rect 2932 3352 2944 3354
rect 2932 3351 2933 3352
rect 2927 3350 2933 3351
rect 2943 3351 2944 3352
rect 2948 3351 2949 3355
rect 2952 3354 2954 3360
rect 3031 3355 3037 3356
rect 3031 3354 3032 3355
rect 2952 3352 3032 3354
rect 2943 3350 2949 3351
rect 3031 3351 3032 3352
rect 3036 3351 3037 3355
rect 3031 3350 3037 3351
rect 2750 3347 2756 3348
rect 2750 3343 2751 3347
rect 2755 3343 2756 3347
rect 2750 3342 2756 3343
rect 2854 3347 2860 3348
rect 2854 3343 2855 3347
rect 2859 3343 2860 3347
rect 2854 3342 2860 3343
rect 2958 3347 2964 3348
rect 2958 3343 2959 3347
rect 2963 3343 2964 3347
rect 2958 3342 2964 3343
rect 2838 3339 2844 3340
rect 2838 3338 2839 3339
rect 2697 3336 2734 3338
rect 2801 3336 2839 3338
rect 2606 3334 2612 3335
rect 2838 3335 2839 3336
rect 2843 3335 2844 3339
rect 2918 3339 2924 3340
rect 2918 3338 2919 3339
rect 2905 3336 2919 3338
rect 2838 3334 2844 3335
rect 2918 3335 2919 3336
rect 2923 3335 2924 3339
rect 2918 3334 2924 3335
rect 110 3328 116 3329
rect 110 3324 111 3328
rect 115 3324 116 3328
rect 110 3323 116 3324
rect 2030 3328 2036 3329
rect 2030 3324 2031 3328
rect 2035 3324 2036 3328
rect 2030 3323 2036 3324
rect 2070 3328 2076 3329
rect 2070 3324 2071 3328
rect 2075 3324 2076 3328
rect 2070 3323 2076 3324
rect 3990 3328 3996 3329
rect 3990 3324 3991 3328
rect 3995 3324 3996 3328
rect 3990 3323 3996 3324
rect 110 3311 116 3312
rect 110 3307 111 3311
rect 115 3307 116 3311
rect 2030 3311 2036 3312
rect 2030 3307 2031 3311
rect 2035 3307 2036 3311
rect 110 3306 116 3307
rect 150 3306 156 3307
rect 150 3302 151 3306
rect 155 3302 156 3306
rect 150 3301 156 3302
rect 318 3306 324 3307
rect 318 3302 319 3306
rect 323 3302 324 3306
rect 318 3301 324 3302
rect 526 3306 532 3307
rect 526 3302 527 3306
rect 531 3302 532 3306
rect 526 3301 532 3302
rect 742 3306 748 3307
rect 742 3302 743 3306
rect 747 3302 748 3306
rect 742 3301 748 3302
rect 958 3306 964 3307
rect 958 3302 959 3306
rect 963 3302 964 3306
rect 958 3301 964 3302
rect 1166 3306 1172 3307
rect 1166 3302 1167 3306
rect 1171 3302 1172 3306
rect 1166 3301 1172 3302
rect 1366 3306 1372 3307
rect 1366 3302 1367 3306
rect 1371 3302 1372 3306
rect 1366 3301 1372 3302
rect 1558 3306 1564 3307
rect 1558 3302 1559 3306
rect 1563 3302 1564 3306
rect 1558 3301 1564 3302
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 1934 3306 1940 3307
rect 2030 3306 2036 3307
rect 2070 3311 2076 3312
rect 2070 3307 2071 3311
rect 2075 3307 2076 3311
rect 3990 3311 3996 3312
rect 3990 3307 3991 3311
rect 3995 3307 3996 3311
rect 2070 3306 2076 3307
rect 2438 3306 2444 3307
rect 1934 3302 1935 3306
rect 1939 3302 1940 3306
rect 1934 3301 1940 3302
rect 2438 3302 2439 3306
rect 2443 3302 2444 3306
rect 2438 3301 2444 3302
rect 2542 3306 2548 3307
rect 2542 3302 2543 3306
rect 2547 3302 2548 3306
rect 2542 3301 2548 3302
rect 2646 3306 2652 3307
rect 2646 3302 2647 3306
rect 2651 3302 2652 3306
rect 2646 3301 2652 3302
rect 2750 3306 2756 3307
rect 2750 3302 2751 3306
rect 2755 3302 2756 3306
rect 2750 3301 2756 3302
rect 2854 3306 2860 3307
rect 2854 3302 2855 3306
rect 2859 3302 2860 3306
rect 2854 3301 2860 3302
rect 2958 3306 2964 3307
rect 3990 3306 3996 3307
rect 2958 3302 2959 3306
rect 2963 3302 2964 3306
rect 2958 3301 2964 3302
rect 383 3291 389 3292
rect 383 3287 384 3291
rect 388 3290 389 3291
rect 994 3291 1000 3292
rect 994 3290 995 3291
rect 388 3288 995 3290
rect 388 3287 389 3288
rect 383 3286 389 3287
rect 994 3287 995 3288
rect 999 3287 1000 3291
rect 994 3286 1000 3287
rect 2526 3274 2532 3275
rect 2526 3270 2527 3274
rect 2531 3270 2532 3274
rect 2070 3269 2076 3270
rect 2526 3269 2532 3270
rect 2630 3274 2636 3275
rect 2630 3270 2631 3274
rect 2635 3270 2636 3274
rect 2630 3269 2636 3270
rect 2734 3274 2740 3275
rect 2734 3270 2735 3274
rect 2739 3270 2740 3274
rect 2734 3269 2740 3270
rect 2838 3274 2844 3275
rect 2838 3270 2839 3274
rect 2843 3270 2844 3274
rect 2838 3269 2844 3270
rect 2942 3274 2948 3275
rect 2942 3270 2943 3274
rect 2947 3270 2948 3274
rect 2942 3269 2948 3270
rect 3046 3274 3052 3275
rect 3046 3270 3047 3274
rect 3051 3270 3052 3274
rect 3046 3269 3052 3270
rect 3150 3274 3156 3275
rect 3150 3270 3151 3274
rect 3155 3270 3156 3274
rect 3150 3269 3156 3270
rect 3254 3274 3260 3275
rect 3254 3270 3255 3274
rect 3259 3270 3260 3274
rect 3254 3269 3260 3270
rect 3990 3269 3996 3270
rect 310 3266 316 3267
rect 310 3262 311 3266
rect 315 3262 316 3266
rect 110 3261 116 3262
rect 310 3261 316 3262
rect 478 3266 484 3267
rect 478 3262 479 3266
rect 483 3262 484 3266
rect 478 3261 484 3262
rect 654 3266 660 3267
rect 654 3262 655 3266
rect 659 3262 660 3266
rect 654 3261 660 3262
rect 846 3266 852 3267
rect 846 3262 847 3266
rect 851 3262 852 3266
rect 846 3261 852 3262
rect 1038 3266 1044 3267
rect 1038 3262 1039 3266
rect 1043 3262 1044 3266
rect 1038 3261 1044 3262
rect 1230 3266 1236 3267
rect 1230 3262 1231 3266
rect 1235 3262 1236 3266
rect 1230 3261 1236 3262
rect 1430 3266 1436 3267
rect 1430 3262 1431 3266
rect 1435 3262 1436 3266
rect 1430 3261 1436 3262
rect 1630 3266 1636 3267
rect 1630 3262 1631 3266
rect 1635 3262 1636 3266
rect 1630 3261 1636 3262
rect 1830 3266 1836 3267
rect 1830 3262 1831 3266
rect 1835 3262 1836 3266
rect 2070 3265 2071 3269
rect 2075 3265 2076 3269
rect 2070 3264 2076 3265
rect 3990 3265 3991 3269
rect 3995 3265 3996 3269
rect 3990 3264 3996 3265
rect 1830 3261 1836 3262
rect 2030 3261 2036 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 110 3256 116 3257
rect 2030 3257 2031 3261
rect 2035 3257 2036 3261
rect 2030 3256 2036 3257
rect 2070 3252 2076 3253
rect 2070 3248 2071 3252
rect 2075 3248 2076 3252
rect 2070 3247 2076 3248
rect 3990 3252 3996 3253
rect 3990 3248 3991 3252
rect 3995 3248 3996 3252
rect 3990 3247 3996 3248
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 110 3239 116 3240
rect 2030 3244 2036 3245
rect 2030 3240 2031 3244
rect 2035 3240 2036 3244
rect 2614 3243 2620 3244
rect 2614 3242 2615 3243
rect 2577 3240 2615 3242
rect 2030 3239 2036 3240
rect 2614 3239 2615 3240
rect 2619 3239 2620 3243
rect 2718 3243 2724 3244
rect 2718 3242 2719 3243
rect 2681 3240 2719 3242
rect 2614 3238 2620 3239
rect 2718 3239 2719 3240
rect 2723 3239 2724 3243
rect 3030 3243 3036 3244
rect 3030 3242 3031 3243
rect 2993 3240 3031 3242
rect 2718 3238 2724 3239
rect 3030 3239 3031 3240
rect 3035 3239 3036 3243
rect 3174 3243 3180 3244
rect 3097 3240 3142 3242
rect 3030 3238 3036 3239
rect 383 3235 389 3236
rect 383 3234 384 3235
rect 361 3232 384 3234
rect 383 3231 384 3232
rect 388 3231 389 3235
rect 383 3230 389 3231
rect 1254 3235 1260 3236
rect 1254 3231 1255 3235
rect 1259 3231 1260 3235
rect 2002 3235 2008 3236
rect 2002 3234 2003 3235
rect 1881 3232 2003 3234
rect 1254 3230 1260 3231
rect 2002 3231 2003 3232
rect 2007 3231 2008 3235
rect 2002 3230 2008 3231
rect 2526 3233 2532 3234
rect 2526 3229 2527 3233
rect 2531 3229 2532 3233
rect 2526 3228 2532 3229
rect 2630 3233 2636 3234
rect 2630 3229 2631 3233
rect 2635 3229 2636 3233
rect 2630 3228 2636 3229
rect 2734 3233 2740 3234
rect 2734 3229 2735 3233
rect 2739 3229 2740 3233
rect 2734 3228 2740 3229
rect 2838 3233 2844 3234
rect 2838 3229 2839 3233
rect 2843 3229 2844 3233
rect 2838 3228 2844 3229
rect 2942 3233 2948 3234
rect 2942 3229 2943 3233
rect 2947 3229 2948 3233
rect 2942 3228 2948 3229
rect 3046 3233 3052 3234
rect 3046 3229 3047 3233
rect 3051 3229 3052 3233
rect 3046 3228 3052 3229
rect 3140 3226 3142 3240
rect 3174 3239 3175 3243
rect 3179 3239 3180 3243
rect 3174 3238 3180 3239
rect 3150 3233 3156 3234
rect 3150 3229 3151 3233
rect 3155 3229 3156 3233
rect 3254 3233 3260 3234
rect 3150 3228 3156 3229
rect 3216 3228 3250 3230
rect 3254 3229 3255 3233
rect 3259 3229 3260 3233
rect 3254 3228 3260 3229
rect 3216 3226 3218 3228
rect 310 3225 316 3226
rect 310 3221 311 3225
rect 315 3221 316 3225
rect 310 3220 316 3221
rect 478 3225 484 3226
rect 478 3221 479 3225
rect 483 3221 484 3225
rect 478 3220 484 3221
rect 654 3225 660 3226
rect 654 3221 655 3225
rect 659 3221 660 3225
rect 654 3220 660 3221
rect 846 3225 852 3226
rect 846 3221 847 3225
rect 851 3221 852 3225
rect 846 3220 852 3221
rect 1038 3225 1044 3226
rect 1038 3221 1039 3225
rect 1043 3221 1044 3225
rect 1038 3220 1044 3221
rect 1230 3225 1236 3226
rect 1230 3221 1231 3225
rect 1235 3221 1236 3225
rect 1230 3220 1236 3221
rect 1430 3225 1436 3226
rect 1430 3221 1431 3225
rect 1435 3221 1436 3225
rect 1430 3220 1436 3221
rect 1630 3225 1636 3226
rect 1630 3221 1631 3225
rect 1635 3221 1636 3225
rect 1630 3220 1636 3221
rect 1830 3225 1836 3226
rect 1830 3221 1831 3225
rect 1835 3221 1836 3225
rect 3140 3224 3218 3226
rect 1830 3220 1836 3221
rect 2599 3223 2605 3224
rect 2599 3219 2600 3223
rect 2604 3219 2605 3223
rect 2703 3223 2709 3224
rect 2599 3218 2605 3219
rect 2614 3219 2620 3220
rect 383 3215 389 3216
rect 383 3211 384 3215
rect 388 3214 389 3215
rect 463 3215 469 3216
rect 463 3214 464 3215
rect 388 3212 464 3214
rect 388 3211 389 3212
rect 383 3210 389 3211
rect 463 3211 464 3212
rect 468 3211 469 3215
rect 463 3210 469 3211
rect 551 3215 557 3216
rect 551 3211 552 3215
rect 556 3214 557 3215
rect 639 3215 645 3216
rect 639 3214 640 3215
rect 556 3212 640 3214
rect 556 3211 557 3212
rect 551 3210 557 3211
rect 639 3211 640 3212
rect 644 3211 645 3215
rect 639 3210 645 3211
rect 727 3215 733 3216
rect 727 3211 728 3215
rect 732 3214 733 3215
rect 831 3215 837 3216
rect 831 3214 832 3215
rect 732 3212 832 3214
rect 732 3211 733 3212
rect 727 3210 733 3211
rect 831 3211 832 3212
rect 836 3211 837 3215
rect 831 3210 837 3211
rect 919 3215 925 3216
rect 919 3211 920 3215
rect 924 3214 925 3215
rect 1023 3215 1029 3216
rect 1023 3214 1024 3215
rect 924 3212 1024 3214
rect 924 3211 925 3212
rect 919 3210 925 3211
rect 1023 3211 1024 3212
rect 1028 3211 1029 3215
rect 1023 3210 1029 3211
rect 1046 3215 1052 3216
rect 1046 3211 1047 3215
rect 1051 3214 1052 3215
rect 1111 3215 1117 3216
rect 1111 3214 1112 3215
rect 1051 3212 1112 3214
rect 1051 3211 1052 3212
rect 1046 3210 1052 3211
rect 1111 3211 1112 3212
rect 1116 3211 1117 3215
rect 1111 3210 1117 3211
rect 1303 3215 1309 3216
rect 1303 3211 1304 3215
rect 1308 3214 1309 3215
rect 1415 3215 1421 3216
rect 1415 3214 1416 3215
rect 1308 3212 1416 3214
rect 1308 3211 1309 3212
rect 1303 3210 1309 3211
rect 1415 3211 1416 3212
rect 1420 3211 1421 3215
rect 1415 3210 1421 3211
rect 1503 3215 1509 3216
rect 1503 3211 1504 3215
rect 1508 3214 1509 3215
rect 1615 3215 1621 3216
rect 1615 3214 1616 3215
rect 1508 3212 1616 3214
rect 1508 3211 1509 3212
rect 1503 3210 1509 3211
rect 1615 3211 1616 3212
rect 1620 3211 1621 3215
rect 1615 3210 1621 3211
rect 1703 3215 1709 3216
rect 1703 3211 1704 3215
rect 1708 3211 1709 3215
rect 1703 3210 1709 3211
rect 1774 3215 1780 3216
rect 1774 3211 1775 3215
rect 1779 3214 1780 3215
rect 1903 3215 1909 3216
rect 1903 3214 1904 3215
rect 1779 3212 1904 3214
rect 1779 3211 1780 3212
rect 1774 3210 1780 3211
rect 1903 3211 1904 3212
rect 1908 3211 1909 3215
rect 2614 3215 2615 3219
rect 2619 3218 2620 3219
rect 2703 3219 2704 3223
rect 2708 3222 2709 3223
rect 2719 3223 2725 3224
rect 2719 3222 2720 3223
rect 2708 3220 2720 3222
rect 2708 3219 2709 3220
rect 2703 3218 2709 3219
rect 2719 3219 2720 3220
rect 2724 3219 2725 3223
rect 2719 3218 2725 3219
rect 2807 3223 2813 3224
rect 2807 3219 2808 3223
rect 2812 3222 2813 3223
rect 2823 3223 2829 3224
rect 2823 3222 2824 3223
rect 2812 3220 2824 3222
rect 2812 3219 2813 3220
rect 2807 3218 2813 3219
rect 2823 3219 2824 3220
rect 2828 3219 2829 3223
rect 2823 3218 2829 3219
rect 2911 3223 2917 3224
rect 2911 3219 2912 3223
rect 2916 3219 2917 3223
rect 2911 3218 2917 3219
rect 3014 3223 3021 3224
rect 3014 3219 3015 3223
rect 3020 3219 3021 3223
rect 3014 3218 3021 3219
rect 3030 3223 3036 3224
rect 3030 3219 3031 3223
rect 3035 3222 3036 3223
rect 3119 3223 3125 3224
rect 3119 3222 3120 3223
rect 3035 3220 3120 3222
rect 3035 3219 3036 3220
rect 3030 3218 3036 3219
rect 3119 3219 3120 3220
rect 3124 3219 3125 3223
rect 3119 3218 3125 3219
rect 3223 3223 3229 3224
rect 3223 3219 3224 3223
rect 3228 3222 3229 3223
rect 3239 3223 3245 3224
rect 3239 3222 3240 3223
rect 3228 3220 3240 3222
rect 3228 3219 3229 3220
rect 3223 3218 3229 3219
rect 3239 3219 3240 3220
rect 3244 3219 3245 3223
rect 3248 3222 3250 3228
rect 3327 3223 3333 3224
rect 3327 3222 3328 3223
rect 3248 3220 3328 3222
rect 3239 3218 3245 3219
rect 3327 3219 3328 3220
rect 3332 3219 3333 3223
rect 3327 3218 3333 3219
rect 2619 3216 2690 3218
rect 2619 3215 2620 3216
rect 2614 3214 2620 3215
rect 1903 3210 1909 3211
rect 2471 3211 2477 3212
rect 1335 3207 1341 3208
rect 1335 3203 1336 3207
rect 1340 3206 1341 3207
rect 1705 3206 1707 3210
rect 2471 3207 2472 3211
rect 2476 3210 2477 3211
rect 2535 3211 2541 3212
rect 2535 3210 2536 3211
rect 2476 3208 2536 3210
rect 2476 3207 2477 3208
rect 2471 3206 2477 3207
rect 2535 3207 2536 3208
rect 2540 3207 2541 3211
rect 2535 3206 2541 3207
rect 2623 3211 2629 3212
rect 2623 3207 2624 3211
rect 2628 3210 2629 3211
rect 2679 3211 2685 3212
rect 2679 3210 2680 3211
rect 2628 3208 2680 3210
rect 2628 3207 2629 3208
rect 2623 3206 2629 3207
rect 2679 3207 2680 3208
rect 2684 3207 2685 3211
rect 2688 3210 2690 3216
rect 2767 3211 2773 3212
rect 2767 3210 2768 3211
rect 2688 3208 2768 3210
rect 2679 3206 2685 3207
rect 2767 3207 2768 3208
rect 2772 3207 2773 3211
rect 2767 3206 2773 3207
rect 2911 3211 2917 3212
rect 2911 3207 2912 3211
rect 2916 3210 2917 3211
rect 2959 3211 2965 3212
rect 2959 3210 2960 3211
rect 2916 3208 2960 3210
rect 2916 3207 2917 3208
rect 2911 3206 2917 3207
rect 2959 3207 2960 3208
rect 2964 3207 2965 3211
rect 2959 3206 2965 3207
rect 3047 3211 3053 3212
rect 3047 3207 3048 3211
rect 3052 3210 3053 3211
rect 3095 3211 3101 3212
rect 3095 3210 3096 3211
rect 3052 3208 3096 3210
rect 3052 3207 3053 3208
rect 3047 3206 3053 3207
rect 3095 3207 3096 3208
rect 3100 3207 3101 3211
rect 3095 3206 3101 3207
rect 3174 3211 3180 3212
rect 3174 3207 3175 3211
rect 3179 3210 3180 3211
rect 3183 3211 3189 3212
rect 3183 3210 3184 3211
rect 3179 3208 3184 3210
rect 3179 3207 3180 3208
rect 3174 3206 3180 3207
rect 3183 3207 3184 3208
rect 3188 3207 3189 3211
rect 3183 3206 3189 3207
rect 3319 3211 3325 3212
rect 3319 3207 3320 3211
rect 3324 3210 3325 3211
rect 3375 3211 3381 3212
rect 3375 3210 3376 3211
rect 3324 3208 3376 3210
rect 3324 3207 3325 3208
rect 3319 3206 3325 3207
rect 3375 3207 3376 3208
rect 3380 3207 3381 3211
rect 3375 3206 3381 3207
rect 3398 3211 3404 3212
rect 3398 3207 3399 3211
rect 3403 3210 3404 3211
rect 3463 3211 3469 3212
rect 3463 3210 3464 3211
rect 3403 3208 3464 3210
rect 3403 3207 3404 3208
rect 3398 3206 3404 3207
rect 3463 3207 3464 3208
rect 3468 3207 3469 3211
rect 3463 3206 3469 3207
rect 1340 3204 1707 3206
rect 1340 3203 1341 3204
rect 1335 3202 1341 3203
rect 2398 3203 2404 3204
rect 695 3199 701 3200
rect 695 3195 696 3199
rect 700 3198 701 3199
rect 743 3199 749 3200
rect 743 3198 744 3199
rect 700 3196 744 3198
rect 700 3195 701 3196
rect 695 3194 701 3195
rect 743 3195 744 3196
rect 748 3195 749 3199
rect 743 3194 749 3195
rect 831 3199 837 3200
rect 831 3195 832 3199
rect 836 3198 837 3199
rect 887 3199 893 3200
rect 887 3198 888 3199
rect 836 3196 888 3198
rect 836 3195 837 3196
rect 831 3194 837 3195
rect 887 3195 888 3196
rect 892 3195 893 3199
rect 887 3194 893 3195
rect 975 3199 981 3200
rect 975 3195 976 3199
rect 980 3198 981 3199
rect 1039 3199 1045 3200
rect 1039 3198 1040 3199
rect 980 3196 1040 3198
rect 980 3195 981 3196
rect 975 3194 981 3195
rect 1039 3195 1040 3196
rect 1044 3195 1045 3199
rect 1039 3194 1045 3195
rect 1126 3199 1133 3200
rect 1126 3195 1127 3199
rect 1132 3195 1133 3199
rect 1126 3194 1133 3195
rect 1254 3199 1260 3200
rect 1254 3195 1255 3199
rect 1259 3198 1260 3199
rect 1279 3199 1285 3200
rect 1279 3198 1280 3199
rect 1259 3196 1280 3198
rect 1259 3195 1260 3196
rect 1254 3194 1260 3195
rect 1279 3195 1280 3196
rect 1284 3195 1285 3199
rect 1423 3199 1429 3200
rect 1423 3198 1424 3199
rect 1279 3194 1285 3195
rect 1308 3196 1424 3198
rect 622 3191 628 3192
rect 622 3187 623 3191
rect 627 3187 628 3191
rect 622 3186 628 3187
rect 758 3191 764 3192
rect 758 3187 759 3191
rect 763 3187 764 3191
rect 758 3186 764 3187
rect 902 3191 908 3192
rect 902 3187 903 3191
rect 907 3187 908 3191
rect 902 3186 908 3187
rect 1054 3191 1060 3192
rect 1054 3187 1055 3191
rect 1059 3187 1060 3191
rect 1054 3186 1060 3187
rect 1206 3191 1212 3192
rect 1206 3187 1207 3191
rect 1211 3187 1212 3191
rect 1206 3186 1212 3187
rect 742 3183 748 3184
rect 742 3182 743 3183
rect 673 3180 743 3182
rect 742 3179 743 3180
rect 747 3179 748 3183
rect 1308 3182 1310 3196
rect 1423 3195 1424 3196
rect 1428 3195 1429 3199
rect 1575 3199 1581 3200
rect 1575 3198 1576 3199
rect 1423 3194 1429 3195
rect 1460 3196 1576 3198
rect 1350 3191 1356 3192
rect 1350 3187 1351 3191
rect 1355 3187 1356 3191
rect 1350 3186 1356 3187
rect 1460 3182 1462 3196
rect 1575 3195 1576 3196
rect 1580 3195 1581 3199
rect 1575 3194 1581 3195
rect 1727 3199 1733 3200
rect 1727 3195 1728 3199
rect 1732 3198 1733 3199
rect 1791 3199 1797 3200
rect 1791 3198 1792 3199
rect 1732 3196 1792 3198
rect 1732 3195 1733 3196
rect 1727 3194 1733 3195
rect 1791 3195 1792 3196
rect 1796 3195 1797 3199
rect 1791 3194 1797 3195
rect 1879 3199 1885 3200
rect 1879 3195 1880 3199
rect 1884 3198 1885 3199
rect 1919 3199 1925 3200
rect 1919 3198 1920 3199
rect 1884 3196 1920 3198
rect 1884 3195 1885 3196
rect 1879 3194 1885 3195
rect 1919 3195 1920 3196
rect 1924 3195 1925 3199
rect 1919 3194 1925 3195
rect 2006 3199 2013 3200
rect 2006 3195 2007 3199
rect 2012 3195 2013 3199
rect 2398 3199 2399 3203
rect 2403 3199 2404 3203
rect 2398 3198 2404 3199
rect 2550 3203 2556 3204
rect 2550 3199 2551 3203
rect 2555 3199 2556 3203
rect 2550 3198 2556 3199
rect 2694 3203 2700 3204
rect 2694 3199 2695 3203
rect 2699 3199 2700 3203
rect 2694 3198 2700 3199
rect 2838 3203 2844 3204
rect 2838 3199 2839 3203
rect 2843 3199 2844 3203
rect 2838 3198 2844 3199
rect 2974 3203 2980 3204
rect 2974 3199 2975 3203
rect 2979 3199 2980 3203
rect 2974 3198 2980 3199
rect 3110 3203 3116 3204
rect 3110 3199 3111 3203
rect 3115 3199 3116 3203
rect 3110 3198 3116 3199
rect 3246 3203 3252 3204
rect 3246 3199 3247 3203
rect 3251 3199 3252 3203
rect 3246 3198 3252 3199
rect 3390 3203 3396 3204
rect 3390 3199 3391 3203
rect 3395 3199 3396 3203
rect 3390 3198 3396 3199
rect 2006 3194 2013 3195
rect 2958 3195 2964 3196
rect 2958 3194 2959 3195
rect 2889 3192 2959 3194
rect 1502 3191 1508 3192
rect 1502 3187 1503 3191
rect 1507 3187 1508 3191
rect 1502 3186 1508 3187
rect 1654 3191 1660 3192
rect 1654 3187 1655 3191
rect 1659 3187 1660 3191
rect 1654 3186 1660 3187
rect 1806 3191 1812 3192
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 1806 3186 1812 3187
rect 1934 3191 1940 3192
rect 1934 3187 1935 3191
rect 1939 3187 1940 3191
rect 1934 3186 1940 3187
rect 2414 3191 2420 3192
rect 2414 3187 2415 3191
rect 2419 3187 2420 3191
rect 2958 3191 2959 3192
rect 2963 3191 2964 3195
rect 2958 3190 2964 3191
rect 3262 3191 3268 3192
rect 2414 3186 2420 3187
rect 3262 3187 3263 3191
rect 3267 3187 3268 3191
rect 3262 3186 3268 3187
rect 2070 3184 2076 3185
rect 1638 3183 1644 3184
rect 1638 3182 1639 3183
rect 1257 3180 1310 3182
rect 1401 3180 1462 3182
rect 1553 3180 1639 3182
rect 742 3178 748 3179
rect 1638 3179 1639 3180
rect 1643 3179 1644 3183
rect 1774 3183 1780 3184
rect 1774 3182 1775 3183
rect 1705 3180 1775 3182
rect 1638 3178 1644 3179
rect 1774 3179 1775 3180
rect 1779 3179 1780 3183
rect 2070 3180 2071 3184
rect 2075 3180 2076 3184
rect 2070 3179 2076 3180
rect 3990 3184 3996 3185
rect 3990 3180 3991 3184
rect 3995 3180 3996 3184
rect 3990 3179 3996 3180
rect 1774 3178 1780 3179
rect 110 3172 116 3173
rect 110 3168 111 3172
rect 115 3168 116 3172
rect 110 3167 116 3168
rect 2030 3172 2036 3173
rect 2030 3168 2031 3172
rect 2035 3168 2036 3172
rect 2030 3167 2036 3168
rect 2070 3167 2076 3168
rect 2070 3163 2071 3167
rect 2075 3163 2076 3167
rect 3990 3167 3996 3168
rect 3990 3163 3991 3167
rect 3995 3163 3996 3167
rect 2070 3162 2076 3163
rect 2398 3162 2404 3163
rect 2398 3158 2399 3162
rect 2403 3158 2404 3162
rect 2398 3157 2404 3158
rect 2550 3162 2556 3163
rect 2550 3158 2551 3162
rect 2555 3158 2556 3162
rect 2550 3157 2556 3158
rect 2694 3162 2700 3163
rect 2694 3158 2695 3162
rect 2699 3158 2700 3162
rect 2694 3157 2700 3158
rect 2838 3162 2844 3163
rect 2838 3158 2839 3162
rect 2843 3158 2844 3162
rect 2838 3157 2844 3158
rect 2974 3162 2980 3163
rect 2974 3158 2975 3162
rect 2979 3158 2980 3162
rect 2974 3157 2980 3158
rect 3110 3162 3116 3163
rect 3110 3158 3111 3162
rect 3115 3158 3116 3162
rect 3110 3157 3116 3158
rect 3246 3162 3252 3163
rect 3246 3158 3247 3162
rect 3251 3158 3252 3162
rect 3246 3157 3252 3158
rect 3390 3162 3396 3163
rect 3990 3162 3996 3163
rect 3390 3158 3391 3162
rect 3395 3158 3396 3162
rect 3390 3157 3396 3158
rect 110 3155 116 3156
rect 110 3151 111 3155
rect 115 3151 116 3155
rect 2030 3155 2036 3156
rect 2030 3151 2031 3155
rect 2035 3151 2036 3155
rect 110 3150 116 3151
rect 622 3150 628 3151
rect 622 3146 623 3150
rect 627 3146 628 3150
rect 622 3145 628 3146
rect 758 3150 764 3151
rect 758 3146 759 3150
rect 763 3146 764 3150
rect 758 3145 764 3146
rect 902 3150 908 3151
rect 902 3146 903 3150
rect 907 3146 908 3150
rect 902 3145 908 3146
rect 1054 3150 1060 3151
rect 1054 3146 1055 3150
rect 1059 3146 1060 3150
rect 1054 3145 1060 3146
rect 1206 3150 1212 3151
rect 1206 3146 1207 3150
rect 1211 3146 1212 3150
rect 1206 3145 1212 3146
rect 1350 3150 1356 3151
rect 1350 3146 1351 3150
rect 1355 3146 1356 3150
rect 1350 3145 1356 3146
rect 1502 3150 1508 3151
rect 1502 3146 1503 3150
rect 1507 3146 1508 3150
rect 1502 3145 1508 3146
rect 1654 3150 1660 3151
rect 1654 3146 1655 3150
rect 1659 3146 1660 3150
rect 1654 3145 1660 3146
rect 1806 3150 1812 3151
rect 1806 3146 1807 3150
rect 1811 3146 1812 3150
rect 1806 3145 1812 3146
rect 1934 3150 1940 3151
rect 2030 3150 2036 3151
rect 1934 3146 1935 3150
rect 1939 3146 1940 3150
rect 1934 3145 1940 3146
rect 598 3118 604 3119
rect 598 3114 599 3118
rect 603 3114 604 3118
rect 110 3113 116 3114
rect 598 3113 604 3114
rect 702 3118 708 3119
rect 702 3114 703 3118
rect 707 3114 708 3118
rect 702 3113 708 3114
rect 806 3118 812 3119
rect 806 3114 807 3118
rect 811 3114 812 3118
rect 806 3113 812 3114
rect 910 3118 916 3119
rect 910 3114 911 3118
rect 915 3114 916 3118
rect 910 3113 916 3114
rect 1038 3118 1044 3119
rect 1038 3114 1039 3118
rect 1043 3114 1044 3118
rect 1038 3113 1044 3114
rect 1182 3118 1188 3119
rect 1182 3114 1183 3118
rect 1187 3114 1188 3118
rect 1182 3113 1188 3114
rect 1358 3118 1364 3119
rect 1358 3114 1359 3118
rect 1363 3114 1364 3118
rect 1358 3113 1364 3114
rect 1550 3118 1556 3119
rect 1550 3114 1551 3118
rect 1555 3114 1556 3118
rect 1550 3113 1556 3114
rect 1750 3118 1756 3119
rect 1750 3114 1751 3118
rect 1755 3114 1756 3118
rect 1750 3113 1756 3114
rect 1934 3118 1940 3119
rect 1934 3114 1935 3118
rect 1939 3114 1940 3118
rect 2110 3118 2116 3119
rect 2110 3114 2111 3118
rect 2115 3114 2116 3118
rect 1934 3113 1940 3114
rect 2030 3113 2036 3114
rect 110 3109 111 3113
rect 115 3109 116 3113
rect 110 3108 116 3109
rect 2030 3109 2031 3113
rect 2035 3109 2036 3113
rect 2030 3108 2036 3109
rect 2070 3113 2076 3114
rect 2110 3113 2116 3114
rect 2342 3118 2348 3119
rect 2342 3114 2343 3118
rect 2347 3114 2348 3118
rect 2342 3113 2348 3114
rect 2582 3118 2588 3119
rect 2582 3114 2583 3118
rect 2587 3114 2588 3118
rect 2582 3113 2588 3114
rect 2798 3118 2804 3119
rect 2798 3114 2799 3118
rect 2803 3114 2804 3118
rect 2798 3113 2804 3114
rect 2998 3118 3004 3119
rect 2998 3114 2999 3118
rect 3003 3114 3004 3118
rect 2998 3113 3004 3114
rect 3190 3118 3196 3119
rect 3190 3114 3191 3118
rect 3195 3114 3196 3118
rect 3190 3113 3196 3114
rect 3374 3118 3380 3119
rect 3374 3114 3375 3118
rect 3379 3114 3380 3118
rect 3374 3113 3380 3114
rect 3566 3118 3572 3119
rect 3566 3114 3567 3118
rect 3571 3114 3572 3118
rect 3566 3113 3572 3114
rect 3990 3113 3996 3114
rect 2070 3109 2071 3113
rect 2075 3109 2076 3113
rect 2070 3108 2076 3109
rect 3990 3109 3991 3113
rect 3995 3109 3996 3113
rect 3990 3108 3996 3109
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 2030 3096 2036 3097
rect 2030 3092 2031 3096
rect 2035 3092 2036 3096
rect 2030 3091 2036 3092
rect 2070 3096 2076 3097
rect 2070 3092 2071 3096
rect 2075 3092 2076 3096
rect 2070 3091 2076 3092
rect 3990 3096 3996 3097
rect 3990 3092 3991 3096
rect 3995 3092 3996 3096
rect 3990 3091 3996 3092
rect 686 3087 692 3088
rect 686 3086 687 3087
rect 649 3084 687 3086
rect 686 3083 687 3084
rect 691 3083 692 3087
rect 790 3087 796 3088
rect 790 3086 791 3087
rect 753 3084 791 3086
rect 686 3082 692 3083
rect 790 3083 791 3084
rect 795 3083 796 3087
rect 894 3087 900 3088
rect 894 3086 895 3087
rect 857 3084 895 3086
rect 790 3082 796 3083
rect 894 3083 895 3084
rect 899 3083 900 3087
rect 1022 3087 1028 3088
rect 1022 3086 1023 3087
rect 961 3084 1023 3086
rect 894 3082 900 3083
rect 1022 3083 1023 3084
rect 1027 3083 1028 3087
rect 1126 3087 1132 3088
rect 1126 3086 1127 3087
rect 1089 3084 1127 3086
rect 1022 3082 1028 3083
rect 1126 3083 1127 3084
rect 1131 3083 1132 3087
rect 2006 3087 2012 3088
rect 2006 3086 2007 3087
rect 1985 3084 2007 3086
rect 1126 3082 1132 3083
rect 2006 3083 2007 3084
rect 2011 3083 2012 3087
rect 2566 3087 2572 3088
rect 2566 3086 2567 3087
rect 2393 3084 2567 3086
rect 2006 3082 2012 3083
rect 2566 3083 2567 3084
rect 2571 3083 2572 3087
rect 2662 3087 2668 3088
rect 2662 3086 2663 3087
rect 2633 3084 2663 3086
rect 2566 3082 2572 3083
rect 2662 3083 2663 3084
rect 2667 3083 2668 3087
rect 2982 3087 2988 3088
rect 2982 3086 2983 3087
rect 2849 3084 2983 3086
rect 2662 3082 2668 3083
rect 2982 3083 2983 3084
rect 2987 3083 2988 3087
rect 3550 3087 3556 3088
rect 3550 3086 3551 3087
rect 3425 3084 3551 3086
rect 2982 3082 2988 3083
rect 3550 3083 3551 3084
rect 3555 3083 3556 3087
rect 3662 3087 3668 3088
rect 3662 3086 3663 3087
rect 3617 3084 3663 3086
rect 3550 3082 3556 3083
rect 3662 3083 3663 3084
rect 3667 3083 3668 3087
rect 3662 3082 3668 3083
rect 598 3077 604 3078
rect 598 3073 599 3077
rect 603 3073 604 3077
rect 598 3072 604 3073
rect 702 3077 708 3078
rect 702 3073 703 3077
rect 707 3073 708 3077
rect 702 3072 708 3073
rect 806 3077 812 3078
rect 806 3073 807 3077
rect 811 3073 812 3077
rect 806 3072 812 3073
rect 910 3077 916 3078
rect 910 3073 911 3077
rect 915 3073 916 3077
rect 910 3072 916 3073
rect 1038 3077 1044 3078
rect 1038 3073 1039 3077
rect 1043 3073 1044 3077
rect 1038 3072 1044 3073
rect 1182 3077 1188 3078
rect 1182 3073 1183 3077
rect 1187 3073 1188 3077
rect 1182 3072 1188 3073
rect 1358 3077 1364 3078
rect 1358 3073 1359 3077
rect 1363 3073 1364 3077
rect 1358 3072 1364 3073
rect 1550 3077 1556 3078
rect 1550 3073 1551 3077
rect 1555 3073 1556 3077
rect 1750 3077 1756 3078
rect 1550 3072 1556 3073
rect 1638 3075 1644 3076
rect 1638 3071 1639 3075
rect 1643 3074 1644 3075
rect 1643 3072 1746 3074
rect 1750 3073 1751 3077
rect 1755 3073 1756 3077
rect 1750 3072 1756 3073
rect 1934 3077 1940 3078
rect 1934 3073 1935 3077
rect 1939 3073 1940 3077
rect 1934 3072 1940 3073
rect 2110 3077 2116 3078
rect 2110 3073 2111 3077
rect 2115 3073 2116 3077
rect 2110 3072 2116 3073
rect 2342 3077 2348 3078
rect 2342 3073 2343 3077
rect 2347 3073 2348 3077
rect 2342 3072 2348 3073
rect 2582 3077 2588 3078
rect 2582 3073 2583 3077
rect 2587 3073 2588 3077
rect 2582 3072 2588 3073
rect 2798 3077 2804 3078
rect 2798 3073 2799 3077
rect 2803 3073 2804 3077
rect 2798 3072 2804 3073
rect 2998 3077 3004 3078
rect 2998 3073 2999 3077
rect 3003 3073 3004 3077
rect 2998 3072 3004 3073
rect 3190 3077 3196 3078
rect 3190 3073 3191 3077
rect 3195 3073 3196 3077
rect 3190 3072 3196 3073
rect 3374 3077 3380 3078
rect 3374 3073 3375 3077
rect 3379 3073 3380 3077
rect 3374 3072 3380 3073
rect 3566 3077 3572 3078
rect 3566 3073 3567 3077
rect 3571 3073 3572 3077
rect 3566 3072 3572 3073
rect 1643 3071 1644 3072
rect 1638 3070 1644 3071
rect 662 3067 668 3068
rect 662 3063 663 3067
rect 667 3066 668 3067
rect 671 3067 677 3068
rect 671 3066 672 3067
rect 667 3064 672 3066
rect 667 3063 668 3064
rect 662 3062 668 3063
rect 671 3063 672 3064
rect 676 3063 677 3067
rect 671 3062 677 3063
rect 686 3067 692 3068
rect 686 3063 687 3067
rect 691 3066 692 3067
rect 775 3067 781 3068
rect 775 3066 776 3067
rect 691 3064 776 3066
rect 691 3063 692 3064
rect 686 3062 692 3063
rect 775 3063 776 3064
rect 780 3063 781 3067
rect 775 3062 781 3063
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3066 796 3067
rect 879 3067 885 3068
rect 879 3066 880 3067
rect 795 3064 880 3066
rect 795 3063 796 3064
rect 790 3062 796 3063
rect 879 3063 880 3064
rect 884 3063 885 3067
rect 879 3062 885 3063
rect 894 3067 900 3068
rect 894 3063 895 3067
rect 899 3066 900 3067
rect 983 3067 989 3068
rect 983 3066 984 3067
rect 899 3064 984 3066
rect 899 3063 900 3064
rect 894 3062 900 3063
rect 983 3063 984 3064
rect 988 3063 989 3067
rect 983 3062 989 3063
rect 1022 3067 1028 3068
rect 1022 3063 1023 3067
rect 1027 3066 1028 3067
rect 1111 3067 1117 3068
rect 1111 3066 1112 3067
rect 1027 3064 1112 3066
rect 1027 3063 1028 3064
rect 1022 3062 1028 3063
rect 1111 3063 1112 3064
rect 1116 3063 1117 3067
rect 1111 3062 1117 3063
rect 1166 3067 1173 3068
rect 1166 3063 1167 3067
rect 1172 3063 1173 3067
rect 1166 3062 1173 3063
rect 1255 3067 1261 3068
rect 1255 3063 1256 3067
rect 1260 3066 1261 3067
rect 1343 3067 1349 3068
rect 1343 3066 1344 3067
rect 1260 3064 1344 3066
rect 1260 3063 1261 3064
rect 1255 3062 1261 3063
rect 1343 3063 1344 3064
rect 1348 3063 1349 3067
rect 1343 3062 1349 3063
rect 1431 3067 1437 3068
rect 1431 3063 1432 3067
rect 1436 3066 1437 3067
rect 1535 3067 1541 3068
rect 1535 3066 1536 3067
rect 1436 3064 1536 3066
rect 1436 3063 1437 3064
rect 1431 3062 1437 3063
rect 1535 3063 1536 3064
rect 1540 3063 1541 3067
rect 1535 3062 1541 3063
rect 1623 3067 1629 3068
rect 1623 3063 1624 3067
rect 1628 3066 1629 3067
rect 1735 3067 1741 3068
rect 1735 3066 1736 3067
rect 1628 3064 1736 3066
rect 1628 3063 1629 3064
rect 1623 3062 1629 3063
rect 1735 3063 1736 3064
rect 1740 3063 1741 3067
rect 1744 3066 1746 3072
rect 1823 3067 1829 3068
rect 1823 3066 1824 3067
rect 1744 3064 1824 3066
rect 1735 3062 1741 3063
rect 1823 3063 1824 3064
rect 1828 3063 1829 3067
rect 1823 3062 1829 3063
rect 2007 3067 2013 3068
rect 2007 3063 2008 3067
rect 2012 3066 2013 3067
rect 2095 3067 2101 3068
rect 2095 3066 2096 3067
rect 2012 3064 2096 3066
rect 2012 3063 2013 3064
rect 2007 3062 2013 3063
rect 2095 3063 2096 3064
rect 2100 3063 2101 3067
rect 2095 3062 2101 3063
rect 2174 3067 2180 3068
rect 2174 3063 2175 3067
rect 2179 3066 2180 3067
rect 2183 3067 2189 3068
rect 2183 3066 2184 3067
rect 2179 3064 2184 3066
rect 2179 3063 2180 3064
rect 2174 3062 2180 3063
rect 2183 3063 2184 3064
rect 2188 3063 2189 3067
rect 2183 3062 2189 3063
rect 2414 3067 2421 3068
rect 2414 3063 2415 3067
rect 2420 3063 2421 3067
rect 2414 3062 2421 3063
rect 2566 3067 2572 3068
rect 2566 3063 2567 3067
rect 2571 3066 2572 3067
rect 2655 3067 2661 3068
rect 2655 3066 2656 3067
rect 2571 3064 2656 3066
rect 2571 3063 2572 3064
rect 2566 3062 2572 3063
rect 2655 3063 2656 3064
rect 2660 3063 2661 3067
rect 2655 3062 2661 3063
rect 2871 3067 2877 3068
rect 2871 3063 2872 3067
rect 2876 3066 2877 3067
rect 2983 3067 2989 3068
rect 2983 3066 2984 3067
rect 2876 3064 2984 3066
rect 2876 3063 2877 3064
rect 2871 3062 2877 3063
rect 2983 3063 2984 3064
rect 2988 3063 2989 3067
rect 2983 3062 2989 3063
rect 3071 3067 3077 3068
rect 3071 3063 3072 3067
rect 3076 3066 3077 3067
rect 3175 3067 3181 3068
rect 3175 3066 3176 3067
rect 3076 3064 3176 3066
rect 3076 3063 3077 3064
rect 3071 3062 3077 3063
rect 3175 3063 3176 3064
rect 3180 3063 3181 3067
rect 3175 3062 3181 3063
rect 3262 3067 3269 3068
rect 3262 3063 3263 3067
rect 3268 3063 3269 3067
rect 3447 3067 3453 3068
rect 3447 3066 3448 3067
rect 3262 3062 3269 3063
rect 3272 3064 3448 3066
rect 2982 3059 2988 3060
rect 398 3055 404 3056
rect 398 3051 399 3055
rect 403 3054 404 3055
rect 958 3055 964 3056
rect 403 3052 746 3054
rect 403 3051 404 3052
rect 398 3050 404 3051
rect 383 3047 389 3048
rect 383 3043 384 3047
rect 388 3046 389 3047
rect 399 3047 405 3048
rect 399 3046 400 3047
rect 388 3044 400 3046
rect 388 3043 389 3044
rect 383 3042 389 3043
rect 399 3043 400 3044
rect 404 3043 405 3047
rect 399 3042 405 3043
rect 487 3047 493 3048
rect 487 3043 488 3047
rect 492 3046 493 3047
rect 511 3047 517 3048
rect 511 3046 512 3047
rect 492 3044 512 3046
rect 492 3043 493 3044
rect 487 3042 493 3043
rect 511 3043 512 3044
rect 516 3043 517 3047
rect 599 3047 605 3048
rect 599 3044 600 3047
rect 511 3042 517 3043
rect 598 3043 600 3044
rect 604 3043 605 3047
rect 310 3039 316 3040
rect 310 3035 311 3039
rect 315 3035 316 3039
rect 310 3034 316 3035
rect 414 3039 420 3040
rect 414 3035 415 3039
rect 419 3035 420 3039
rect 414 3034 420 3035
rect 526 3039 532 3040
rect 526 3035 527 3039
rect 531 3035 532 3039
rect 598 3039 599 3043
rect 603 3042 605 3043
rect 711 3047 717 3048
rect 711 3043 712 3047
rect 716 3046 717 3047
rect 735 3047 741 3048
rect 735 3046 736 3047
rect 716 3044 736 3046
rect 716 3043 717 3044
rect 711 3042 717 3043
rect 735 3043 736 3044
rect 740 3043 741 3047
rect 744 3046 746 3052
rect 958 3051 959 3055
rect 963 3054 964 3055
rect 2982 3055 2983 3059
rect 2987 3058 2988 3059
rect 3272 3058 3274 3064
rect 3447 3063 3448 3064
rect 3452 3063 3453 3067
rect 3447 3062 3453 3063
rect 3550 3067 3556 3068
rect 3550 3063 3551 3067
rect 3555 3066 3556 3067
rect 3639 3067 3645 3068
rect 3639 3066 3640 3067
rect 3555 3064 3640 3066
rect 3555 3063 3556 3064
rect 3550 3062 3556 3063
rect 3639 3063 3640 3064
rect 3644 3063 3645 3067
rect 3639 3062 3645 3063
rect 2987 3056 3274 3058
rect 2987 3055 2988 3056
rect 2982 3054 2988 3055
rect 963 3052 1411 3054
rect 963 3051 964 3052
rect 958 3050 964 3051
rect 1409 3048 1411 3052
rect 2183 3051 2189 3052
rect 823 3047 829 3048
rect 823 3046 824 3047
rect 744 3044 824 3046
rect 735 3042 741 3043
rect 823 3043 824 3044
rect 828 3043 829 3047
rect 823 3042 829 3043
rect 935 3047 941 3048
rect 935 3043 936 3047
rect 940 3046 941 3047
rect 959 3047 965 3048
rect 959 3046 960 3047
rect 940 3044 960 3046
rect 940 3043 941 3044
rect 935 3042 941 3043
rect 959 3043 960 3044
rect 964 3043 965 3047
rect 959 3042 965 3043
rect 1047 3047 1053 3048
rect 1047 3043 1048 3047
rect 1052 3046 1053 3047
rect 1079 3047 1085 3048
rect 1079 3046 1080 3047
rect 1052 3044 1080 3046
rect 1052 3043 1053 3044
rect 1047 3042 1053 3043
rect 1079 3043 1080 3044
rect 1084 3043 1085 3047
rect 1079 3042 1085 3043
rect 1166 3047 1173 3048
rect 1166 3043 1167 3047
rect 1172 3043 1173 3047
rect 1166 3042 1173 3043
rect 1287 3047 1293 3048
rect 1287 3043 1288 3047
rect 1292 3046 1293 3047
rect 1319 3047 1325 3048
rect 1319 3046 1320 3047
rect 1292 3044 1320 3046
rect 1292 3043 1293 3044
rect 1287 3042 1293 3043
rect 1319 3043 1320 3044
rect 1324 3043 1325 3047
rect 1319 3042 1325 3043
rect 1407 3047 1413 3048
rect 1407 3043 1408 3047
rect 1412 3043 1413 3047
rect 2183 3047 2184 3051
rect 2188 3050 2189 3051
rect 2247 3051 2253 3052
rect 2247 3050 2248 3051
rect 2188 3048 2248 3050
rect 2188 3047 2189 3048
rect 2183 3046 2189 3047
rect 2247 3047 2248 3048
rect 2252 3047 2253 3051
rect 2247 3046 2253 3047
rect 2335 3051 2341 3052
rect 2335 3047 2336 3051
rect 2340 3050 2341 3051
rect 2439 3051 2445 3052
rect 2439 3050 2440 3051
rect 2340 3048 2440 3050
rect 2340 3047 2341 3048
rect 2335 3046 2341 3047
rect 2439 3047 2440 3048
rect 2444 3047 2445 3051
rect 2439 3046 2445 3047
rect 2526 3051 2533 3052
rect 2526 3047 2527 3051
rect 2532 3047 2533 3051
rect 2526 3046 2533 3047
rect 2662 3051 2668 3052
rect 2662 3047 2663 3051
rect 2667 3050 2668 3051
rect 2727 3051 2733 3052
rect 2727 3050 2728 3051
rect 2667 3048 2728 3050
rect 2667 3047 2668 3048
rect 2662 3046 2668 3047
rect 2727 3047 2728 3048
rect 2732 3047 2733 3051
rect 2927 3051 2933 3052
rect 2927 3050 2928 3051
rect 2727 3046 2733 3047
rect 2839 3048 2928 3050
rect 1407 3042 1413 3043
rect 2110 3043 2116 3044
rect 603 3039 604 3042
rect 598 3038 604 3039
rect 638 3039 644 3040
rect 526 3034 532 3035
rect 638 3035 639 3039
rect 643 3035 644 3039
rect 638 3034 644 3035
rect 750 3039 756 3040
rect 750 3035 751 3039
rect 755 3035 756 3039
rect 750 3034 756 3035
rect 862 3039 868 3040
rect 862 3035 863 3039
rect 867 3035 868 3039
rect 862 3034 868 3035
rect 974 3039 980 3040
rect 974 3035 975 3039
rect 979 3035 980 3039
rect 974 3034 980 3035
rect 1094 3039 1100 3040
rect 1094 3035 1095 3039
rect 1099 3035 1100 3039
rect 1094 3034 1100 3035
rect 1214 3039 1220 3040
rect 1214 3035 1215 3039
rect 1219 3035 1220 3039
rect 1214 3034 1220 3035
rect 1334 3039 1340 3040
rect 1334 3035 1335 3039
rect 1339 3035 1340 3039
rect 2110 3039 2111 3043
rect 2115 3039 2116 3043
rect 2110 3038 2116 3039
rect 2262 3043 2268 3044
rect 2262 3039 2263 3043
rect 2267 3039 2268 3043
rect 2262 3038 2268 3039
rect 2454 3043 2460 3044
rect 2454 3039 2455 3043
rect 2459 3039 2460 3043
rect 2454 3038 2460 3039
rect 2654 3043 2660 3044
rect 2654 3039 2655 3043
rect 2659 3039 2660 3043
rect 2654 3038 2660 3039
rect 1334 3034 1340 3035
rect 2174 3035 2180 3036
rect 2174 3034 2175 3035
rect 2161 3032 2175 3034
rect 398 3031 404 3032
rect 398 3030 399 3031
rect 361 3028 399 3030
rect 398 3027 399 3028
rect 403 3027 404 3031
rect 958 3031 964 3032
rect 958 3030 959 3031
rect 913 3028 959 3030
rect 398 3026 404 3027
rect 662 3027 668 3028
rect 662 3023 663 3027
rect 667 3023 668 3027
rect 958 3027 959 3028
rect 963 3027 964 3031
rect 2174 3031 2175 3032
rect 2179 3031 2180 3035
rect 2839 3034 2841 3048
rect 2927 3047 2928 3048
rect 2932 3047 2933 3051
rect 2927 3046 2933 3047
rect 3127 3051 3133 3052
rect 3127 3047 3128 3051
rect 3132 3050 3133 3051
rect 3239 3051 3245 3052
rect 3239 3050 3240 3051
rect 3132 3048 3240 3050
rect 3132 3047 3133 3048
rect 3127 3046 3133 3047
rect 3239 3047 3240 3048
rect 3244 3047 3245 3051
rect 3239 3046 3245 3047
rect 3327 3051 3333 3052
rect 3327 3047 3328 3051
rect 3332 3050 3333 3051
rect 3439 3051 3445 3052
rect 3439 3050 3440 3051
rect 3332 3048 3440 3050
rect 3332 3047 3333 3048
rect 3327 3046 3333 3047
rect 3439 3047 3440 3048
rect 3444 3047 3445 3051
rect 3439 3046 3445 3047
rect 3527 3051 3533 3052
rect 3527 3047 3528 3051
rect 3532 3050 3533 3051
rect 3639 3051 3645 3052
rect 3639 3050 3640 3051
rect 3532 3048 3640 3050
rect 3532 3047 3533 3048
rect 3527 3046 3533 3047
rect 3639 3047 3640 3048
rect 3644 3047 3645 3051
rect 3639 3046 3645 3047
rect 3662 3051 3668 3052
rect 3662 3047 3663 3051
rect 3667 3050 3668 3051
rect 3727 3051 3733 3052
rect 3727 3050 3728 3051
rect 3667 3048 3728 3050
rect 3667 3047 3668 3048
rect 3662 3046 3668 3047
rect 3727 3047 3728 3048
rect 3732 3047 3733 3051
rect 3727 3046 3733 3047
rect 2854 3043 2860 3044
rect 2854 3039 2855 3043
rect 2859 3039 2860 3043
rect 2854 3038 2860 3039
rect 3054 3043 3060 3044
rect 3054 3039 3055 3043
rect 3059 3039 3060 3043
rect 3054 3038 3060 3039
rect 3254 3043 3260 3044
rect 3254 3039 3255 3043
rect 3259 3039 3260 3043
rect 3254 3038 3260 3039
rect 3454 3043 3460 3044
rect 3454 3039 3455 3043
rect 3459 3039 3460 3043
rect 3454 3038 3460 3039
rect 3654 3043 3660 3044
rect 3654 3039 3655 3043
rect 3659 3039 3660 3043
rect 3654 3038 3660 3039
rect 2918 3035 2924 3036
rect 2918 3034 2919 3035
rect 2705 3032 2841 3034
rect 2905 3032 2919 3034
rect 2174 3030 2180 3031
rect 2918 3031 2919 3032
rect 2923 3031 2924 3035
rect 3150 3035 3156 3036
rect 3150 3034 3151 3035
rect 3105 3032 3151 3034
rect 2918 3030 2924 3031
rect 3150 3031 3151 3032
rect 3155 3031 3156 3035
rect 3150 3030 3156 3031
rect 958 3026 964 3027
rect 1206 3027 1212 3028
rect 662 3022 668 3023
rect 1206 3023 1207 3027
rect 1211 3023 1212 3027
rect 1206 3022 1212 3023
rect 2070 3024 2076 3025
rect 110 3020 116 3021
rect 110 3016 111 3020
rect 115 3016 116 3020
rect 110 3015 116 3016
rect 2030 3020 2036 3021
rect 2030 3016 2031 3020
rect 2035 3016 2036 3020
rect 2070 3020 2071 3024
rect 2075 3020 2076 3024
rect 2070 3019 2076 3020
rect 3990 3024 3996 3025
rect 3990 3020 3991 3024
rect 3995 3020 3996 3024
rect 3990 3019 3996 3020
rect 2030 3015 2036 3016
rect 2070 3007 2076 3008
rect 110 3003 116 3004
rect 110 2999 111 3003
rect 115 2999 116 3003
rect 2030 3003 2036 3004
rect 2030 2999 2031 3003
rect 2035 2999 2036 3003
rect 2070 3003 2071 3007
rect 2075 3003 2076 3007
rect 3990 3007 3996 3008
rect 3990 3003 3991 3007
rect 3995 3003 3996 3007
rect 2070 3002 2076 3003
rect 2110 3002 2116 3003
rect 110 2998 116 2999
rect 310 2998 316 2999
rect 310 2994 311 2998
rect 315 2994 316 2998
rect 310 2993 316 2994
rect 414 2998 420 2999
rect 414 2994 415 2998
rect 419 2994 420 2998
rect 414 2993 420 2994
rect 526 2998 532 2999
rect 526 2994 527 2998
rect 531 2994 532 2998
rect 526 2993 532 2994
rect 638 2998 644 2999
rect 638 2994 639 2998
rect 643 2994 644 2998
rect 638 2993 644 2994
rect 750 2998 756 2999
rect 750 2994 751 2998
rect 755 2994 756 2998
rect 750 2993 756 2994
rect 862 2998 868 2999
rect 862 2994 863 2998
rect 867 2994 868 2998
rect 862 2993 868 2994
rect 974 2998 980 2999
rect 974 2994 975 2998
rect 979 2994 980 2998
rect 974 2993 980 2994
rect 1094 2998 1100 2999
rect 1094 2994 1095 2998
rect 1099 2994 1100 2998
rect 1094 2993 1100 2994
rect 1214 2998 1220 2999
rect 1214 2994 1215 2998
rect 1219 2994 1220 2998
rect 1214 2993 1220 2994
rect 1334 2998 1340 2999
rect 2030 2998 2036 2999
rect 2110 2998 2111 3002
rect 2115 2998 2116 3002
rect 1334 2994 1335 2998
rect 1339 2994 1340 2998
rect 2110 2997 2116 2998
rect 2262 3002 2268 3003
rect 2262 2998 2263 3002
rect 2267 2998 2268 3002
rect 2262 2997 2268 2998
rect 2454 3002 2460 3003
rect 2454 2998 2455 3002
rect 2459 2998 2460 3002
rect 2454 2997 2460 2998
rect 2654 3002 2660 3003
rect 2654 2998 2655 3002
rect 2659 2998 2660 3002
rect 2654 2997 2660 2998
rect 2854 3002 2860 3003
rect 2854 2998 2855 3002
rect 2859 2998 2860 3002
rect 2854 2997 2860 2998
rect 3054 3002 3060 3003
rect 3054 2998 3055 3002
rect 3059 2998 3060 3002
rect 3054 2997 3060 2998
rect 3254 3002 3260 3003
rect 3254 2998 3255 3002
rect 3259 2998 3260 3002
rect 3254 2997 3260 2998
rect 3454 3002 3460 3003
rect 3454 2998 3455 3002
rect 3459 2998 3460 3002
rect 3454 2997 3460 2998
rect 3654 3002 3660 3003
rect 3990 3002 3996 3003
rect 3654 2998 3655 3002
rect 3659 2998 3660 3002
rect 3654 2997 3660 2998
rect 1334 2993 1340 2994
rect 2338 2987 2344 2988
rect 2338 2983 2339 2987
rect 2343 2986 2344 2987
rect 2526 2987 2532 2988
rect 2526 2986 2527 2987
rect 2343 2984 2527 2986
rect 2343 2983 2344 2984
rect 2338 2982 2344 2983
rect 2526 2983 2527 2984
rect 2531 2983 2532 2987
rect 2526 2982 2532 2983
rect 2110 2970 2116 2971
rect 2110 2966 2111 2970
rect 2115 2966 2116 2970
rect 2070 2965 2076 2966
rect 2110 2965 2116 2966
rect 2358 2970 2364 2971
rect 2358 2966 2359 2970
rect 2363 2966 2364 2970
rect 2358 2965 2364 2966
rect 2606 2970 2612 2971
rect 2606 2966 2607 2970
rect 2611 2966 2612 2970
rect 2606 2965 2612 2966
rect 2846 2970 2852 2971
rect 2846 2966 2847 2970
rect 2851 2966 2852 2970
rect 2846 2965 2852 2966
rect 3078 2970 3084 2971
rect 3078 2966 3079 2970
rect 3083 2966 3084 2970
rect 3078 2965 3084 2966
rect 3302 2970 3308 2971
rect 3302 2966 3303 2970
rect 3307 2966 3308 2970
rect 3302 2965 3308 2966
rect 3534 2970 3540 2971
rect 3534 2966 3535 2970
rect 3539 2966 3540 2970
rect 3534 2965 3540 2966
rect 3766 2970 3772 2971
rect 3766 2966 3767 2970
rect 3771 2966 3772 2970
rect 3766 2965 3772 2966
rect 3990 2965 3996 2966
rect 2070 2961 2071 2965
rect 2075 2961 2076 2965
rect 2070 2960 2076 2961
rect 3990 2961 3991 2965
rect 3995 2961 3996 2965
rect 3990 2960 3996 2961
rect 150 2958 156 2959
rect 150 2954 151 2958
rect 155 2954 156 2958
rect 110 2953 116 2954
rect 150 2953 156 2954
rect 270 2958 276 2959
rect 270 2954 271 2958
rect 275 2954 276 2958
rect 270 2953 276 2954
rect 430 2958 436 2959
rect 430 2954 431 2958
rect 435 2954 436 2958
rect 430 2953 436 2954
rect 606 2958 612 2959
rect 606 2954 607 2958
rect 611 2954 612 2958
rect 606 2953 612 2954
rect 782 2958 788 2959
rect 782 2954 783 2958
rect 787 2954 788 2958
rect 782 2953 788 2954
rect 958 2958 964 2959
rect 958 2954 959 2958
rect 963 2954 964 2958
rect 958 2953 964 2954
rect 1134 2958 1140 2959
rect 1134 2954 1135 2958
rect 1139 2954 1140 2958
rect 1134 2953 1140 2954
rect 1302 2958 1308 2959
rect 1302 2954 1303 2958
rect 1307 2954 1308 2958
rect 1302 2953 1308 2954
rect 1470 2958 1476 2959
rect 1470 2954 1471 2958
rect 1475 2954 1476 2958
rect 1470 2953 1476 2954
rect 1646 2958 1652 2959
rect 1646 2954 1647 2958
rect 1651 2954 1652 2958
rect 1646 2953 1652 2954
rect 2030 2953 2036 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 110 2948 116 2949
rect 2030 2949 2031 2953
rect 2035 2949 2036 2953
rect 2030 2948 2036 2949
rect 2070 2948 2076 2949
rect 2070 2944 2071 2948
rect 2075 2944 2076 2948
rect 2070 2943 2076 2944
rect 3990 2948 3996 2949
rect 3990 2944 3991 2948
rect 3995 2944 3996 2948
rect 3990 2943 3996 2944
rect 2338 2939 2344 2940
rect 2338 2938 2339 2939
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 110 2931 116 2932
rect 2030 2936 2036 2937
rect 2161 2936 2339 2938
rect 2030 2932 2031 2936
rect 2035 2932 2036 2936
rect 2338 2935 2339 2936
rect 2343 2935 2344 2939
rect 3286 2939 3292 2940
rect 3286 2938 3287 2939
rect 3129 2936 3287 2938
rect 2338 2934 2344 2935
rect 3286 2935 3287 2936
rect 3291 2935 3292 2939
rect 3518 2939 3524 2940
rect 3518 2938 3519 2939
rect 3353 2936 3519 2938
rect 3286 2934 3292 2935
rect 3518 2935 3519 2936
rect 3523 2935 3524 2939
rect 3750 2939 3756 2940
rect 3750 2938 3751 2939
rect 3585 2936 3751 2938
rect 3518 2934 3524 2935
rect 3750 2935 3751 2936
rect 3755 2935 3756 2939
rect 3871 2939 3877 2940
rect 3871 2938 3872 2939
rect 3817 2936 3872 2938
rect 3750 2934 3756 2935
rect 3871 2935 3872 2936
rect 3876 2935 3877 2939
rect 3871 2934 3877 2935
rect 2030 2931 2036 2932
rect 2110 2929 2116 2930
rect 230 2927 236 2928
rect 230 2926 231 2927
rect 201 2924 231 2926
rect 230 2923 231 2924
rect 235 2923 236 2927
rect 230 2922 236 2923
rect 598 2927 604 2928
rect 598 2923 599 2927
rect 603 2923 604 2927
rect 598 2922 604 2923
rect 982 2927 988 2928
rect 982 2923 983 2927
rect 987 2923 988 2927
rect 1266 2927 1272 2928
rect 1266 2926 1267 2927
rect 1185 2924 1267 2926
rect 982 2922 988 2923
rect 1266 2923 1267 2924
rect 1271 2923 1272 2927
rect 1454 2927 1460 2928
rect 1454 2926 1455 2927
rect 1353 2924 1455 2926
rect 1266 2922 1272 2923
rect 1454 2923 1455 2924
rect 1459 2923 1460 2927
rect 1630 2927 1636 2928
rect 1630 2926 1631 2927
rect 1521 2924 1631 2926
rect 1454 2922 1460 2923
rect 1630 2923 1631 2924
rect 1635 2923 1636 2927
rect 1718 2927 1724 2928
rect 1718 2926 1719 2927
rect 1697 2924 1719 2926
rect 1630 2922 1636 2923
rect 1718 2923 1719 2924
rect 1723 2923 1724 2927
rect 2110 2925 2111 2929
rect 2115 2925 2116 2929
rect 2110 2924 2116 2925
rect 2358 2929 2364 2930
rect 2358 2925 2359 2929
rect 2363 2925 2364 2929
rect 2606 2929 2612 2930
rect 2358 2924 2364 2925
rect 2422 2927 2428 2928
rect 1718 2922 1724 2923
rect 2422 2923 2423 2927
rect 2427 2926 2428 2927
rect 2591 2927 2597 2928
rect 2591 2926 2592 2927
rect 2427 2924 2592 2926
rect 2427 2923 2428 2924
rect 2422 2922 2428 2923
rect 2591 2923 2592 2924
rect 2596 2923 2597 2927
rect 2606 2925 2607 2929
rect 2611 2925 2612 2929
rect 2606 2924 2612 2925
rect 2846 2929 2852 2930
rect 2846 2925 2847 2929
rect 2851 2925 2852 2929
rect 2846 2924 2852 2925
rect 3078 2929 3084 2930
rect 3078 2925 3079 2929
rect 3083 2925 3084 2929
rect 3078 2924 3084 2925
rect 3302 2929 3308 2930
rect 3302 2925 3303 2929
rect 3307 2925 3308 2929
rect 3302 2924 3308 2925
rect 3534 2929 3540 2930
rect 3534 2925 3535 2929
rect 3539 2925 3540 2929
rect 3534 2924 3540 2925
rect 3766 2929 3772 2930
rect 3766 2925 3767 2929
rect 3771 2925 3772 2929
rect 3766 2924 3772 2925
rect 2591 2922 2597 2923
rect 2183 2919 2189 2920
rect 150 2917 156 2918
rect 150 2913 151 2917
rect 155 2913 156 2917
rect 150 2912 156 2913
rect 270 2917 276 2918
rect 270 2913 271 2917
rect 275 2913 276 2917
rect 270 2912 276 2913
rect 430 2917 436 2918
rect 430 2913 431 2917
rect 435 2913 436 2917
rect 430 2912 436 2913
rect 606 2917 612 2918
rect 606 2913 607 2917
rect 611 2913 612 2917
rect 606 2912 612 2913
rect 782 2917 788 2918
rect 782 2913 783 2917
rect 787 2913 788 2917
rect 782 2912 788 2913
rect 958 2917 964 2918
rect 958 2913 959 2917
rect 963 2913 964 2917
rect 958 2912 964 2913
rect 1134 2917 1140 2918
rect 1134 2913 1135 2917
rect 1139 2913 1140 2917
rect 1134 2912 1140 2913
rect 1302 2917 1308 2918
rect 1302 2913 1303 2917
rect 1307 2913 1308 2917
rect 1302 2912 1308 2913
rect 1470 2917 1476 2918
rect 1470 2913 1471 2917
rect 1475 2913 1476 2917
rect 1470 2912 1476 2913
rect 1646 2917 1652 2918
rect 1646 2913 1647 2917
rect 1651 2913 1652 2917
rect 2183 2915 2184 2919
rect 2188 2918 2189 2919
rect 2343 2919 2349 2920
rect 2343 2918 2344 2919
rect 2188 2916 2344 2918
rect 2188 2915 2189 2916
rect 2183 2914 2189 2915
rect 2343 2915 2344 2916
rect 2348 2915 2349 2919
rect 2343 2914 2349 2915
rect 2431 2919 2440 2920
rect 2431 2915 2432 2919
rect 2439 2915 2440 2919
rect 2431 2914 2440 2915
rect 2679 2919 2685 2920
rect 2679 2915 2680 2919
rect 2684 2918 2685 2919
rect 2831 2919 2837 2920
rect 2831 2918 2832 2919
rect 2684 2916 2832 2918
rect 2684 2915 2685 2916
rect 2679 2914 2685 2915
rect 2831 2915 2832 2916
rect 2836 2915 2837 2919
rect 2831 2914 2837 2915
rect 2918 2919 2925 2920
rect 2918 2915 2919 2919
rect 2924 2915 2925 2919
rect 2918 2914 2925 2915
rect 3150 2919 3157 2920
rect 3150 2915 3151 2919
rect 3156 2915 3157 2919
rect 3150 2914 3157 2915
rect 3286 2919 3292 2920
rect 3286 2915 3287 2919
rect 3291 2918 3292 2919
rect 3375 2919 3381 2920
rect 3375 2918 3376 2919
rect 3291 2916 3376 2918
rect 3291 2915 3292 2916
rect 3286 2914 3292 2915
rect 3375 2915 3376 2916
rect 3380 2915 3381 2919
rect 3375 2914 3381 2915
rect 3518 2919 3524 2920
rect 3518 2915 3519 2919
rect 3523 2918 3524 2919
rect 3607 2919 3613 2920
rect 3607 2918 3608 2919
rect 3523 2916 3608 2918
rect 3523 2915 3524 2916
rect 3518 2914 3524 2915
rect 3607 2915 3608 2916
rect 3612 2915 3613 2919
rect 3607 2914 3613 2915
rect 3750 2919 3756 2920
rect 3750 2915 3751 2919
rect 3755 2918 3756 2919
rect 3839 2919 3845 2920
rect 3839 2918 3840 2919
rect 3755 2916 3840 2918
rect 3755 2915 3756 2916
rect 3750 2914 3756 2915
rect 3839 2915 3840 2916
rect 3844 2915 3845 2919
rect 3839 2914 3845 2915
rect 1646 2912 1652 2913
rect 223 2907 229 2908
rect 223 2903 224 2907
rect 228 2906 229 2907
rect 255 2907 261 2908
rect 255 2906 256 2907
rect 228 2904 256 2906
rect 228 2903 229 2904
rect 223 2902 229 2903
rect 255 2903 256 2904
rect 260 2903 261 2907
rect 255 2902 261 2903
rect 343 2907 349 2908
rect 343 2903 344 2907
rect 348 2906 349 2907
rect 415 2907 421 2908
rect 415 2906 416 2907
rect 348 2904 416 2906
rect 348 2903 349 2904
rect 343 2902 349 2903
rect 415 2903 416 2904
rect 420 2903 421 2907
rect 415 2902 421 2903
rect 503 2907 509 2908
rect 503 2903 504 2907
rect 508 2906 509 2907
rect 514 2907 520 2908
rect 514 2906 515 2907
rect 508 2904 515 2906
rect 508 2903 509 2904
rect 503 2902 509 2903
rect 514 2903 515 2904
rect 519 2903 520 2907
rect 514 2902 520 2903
rect 679 2907 685 2908
rect 679 2903 680 2907
rect 684 2906 685 2907
rect 767 2907 773 2908
rect 767 2906 768 2907
rect 684 2904 768 2906
rect 684 2903 685 2904
rect 679 2902 685 2903
rect 767 2903 768 2904
rect 772 2903 773 2907
rect 855 2907 861 2908
rect 855 2906 856 2907
rect 767 2902 773 2903
rect 776 2904 856 2906
rect 230 2899 236 2900
rect 230 2895 231 2899
rect 235 2898 236 2899
rect 776 2898 778 2904
rect 855 2903 856 2904
rect 860 2903 861 2907
rect 855 2902 861 2903
rect 1031 2907 1040 2908
rect 1031 2903 1032 2907
rect 1039 2903 1040 2907
rect 1031 2902 1040 2903
rect 1206 2907 1213 2908
rect 1206 2903 1207 2907
rect 1212 2903 1213 2907
rect 1206 2902 1213 2903
rect 1266 2907 1272 2908
rect 1266 2903 1267 2907
rect 1271 2906 1272 2907
rect 1375 2907 1381 2908
rect 1375 2906 1376 2907
rect 1271 2904 1376 2906
rect 1271 2903 1272 2904
rect 1266 2902 1272 2903
rect 1375 2903 1376 2904
rect 1380 2903 1381 2907
rect 1375 2902 1381 2903
rect 1454 2907 1460 2908
rect 1454 2903 1455 2907
rect 1459 2906 1460 2907
rect 1543 2907 1549 2908
rect 1543 2906 1544 2907
rect 1459 2904 1544 2906
rect 1459 2903 1460 2904
rect 1454 2902 1460 2903
rect 1543 2903 1544 2904
rect 1548 2903 1549 2907
rect 1543 2902 1549 2903
rect 1630 2907 1636 2908
rect 1630 2903 1631 2907
rect 1635 2906 1636 2907
rect 1719 2907 1725 2908
rect 1719 2906 1720 2907
rect 1635 2904 1720 2906
rect 1635 2903 1636 2904
rect 1630 2902 1636 2903
rect 1719 2903 1720 2904
rect 1724 2903 1725 2907
rect 1719 2902 1725 2903
rect 235 2896 778 2898
rect 2183 2899 2189 2900
rect 235 2895 236 2896
rect 230 2894 236 2895
rect 2183 2895 2184 2899
rect 2188 2898 2189 2899
rect 2263 2899 2269 2900
rect 2263 2898 2264 2899
rect 2188 2896 2264 2898
rect 2188 2895 2189 2896
rect 2183 2894 2189 2895
rect 2263 2895 2264 2896
rect 2268 2895 2269 2899
rect 2263 2894 2269 2895
rect 2351 2899 2357 2900
rect 2351 2895 2352 2899
rect 2356 2898 2357 2899
rect 2422 2899 2428 2900
rect 2422 2898 2423 2899
rect 2356 2896 2423 2898
rect 2356 2895 2357 2896
rect 2351 2894 2357 2895
rect 2422 2895 2423 2896
rect 2427 2895 2428 2899
rect 2422 2894 2428 2895
rect 2434 2899 2440 2900
rect 2434 2895 2435 2899
rect 2439 2898 2440 2899
rect 2471 2899 2477 2900
rect 2471 2898 2472 2899
rect 2439 2896 2472 2898
rect 2439 2895 2440 2896
rect 2434 2894 2440 2895
rect 2471 2895 2472 2896
rect 2476 2895 2477 2899
rect 2471 2894 2477 2895
rect 2559 2899 2565 2900
rect 2559 2895 2560 2899
rect 2564 2898 2565 2899
rect 2679 2899 2685 2900
rect 2679 2898 2680 2899
rect 2564 2896 2680 2898
rect 2564 2895 2565 2896
rect 2559 2894 2565 2895
rect 2679 2895 2680 2896
rect 2684 2895 2685 2899
rect 2679 2894 2685 2895
rect 2767 2899 2773 2900
rect 2767 2895 2768 2899
rect 2772 2898 2773 2899
rect 2887 2899 2893 2900
rect 2887 2898 2888 2899
rect 2772 2896 2888 2898
rect 2772 2895 2773 2896
rect 2767 2894 2773 2895
rect 2887 2895 2888 2896
rect 2892 2895 2893 2899
rect 2887 2894 2893 2895
rect 2974 2899 2981 2900
rect 2974 2895 2975 2899
rect 2980 2895 2981 2899
rect 2974 2894 2981 2895
rect 3183 2899 3189 2900
rect 3183 2895 3184 2899
rect 3188 2898 3189 2899
rect 3287 2899 3293 2900
rect 3287 2898 3288 2899
rect 3188 2896 3288 2898
rect 3188 2895 3189 2896
rect 3183 2894 3189 2895
rect 3287 2895 3288 2896
rect 3292 2895 3293 2899
rect 3287 2894 3293 2895
rect 3375 2899 3381 2900
rect 3375 2895 3376 2899
rect 3380 2898 3381 2899
rect 3479 2899 3485 2900
rect 3479 2898 3480 2899
rect 3380 2896 3480 2898
rect 3380 2895 3381 2896
rect 3375 2894 3381 2895
rect 3479 2895 3480 2896
rect 3484 2895 3485 2899
rect 3479 2894 3485 2895
rect 3567 2899 3573 2900
rect 3567 2895 3568 2899
rect 3572 2898 3573 2899
rect 3671 2899 3677 2900
rect 3671 2898 3672 2899
rect 3572 2896 3672 2898
rect 3572 2895 3573 2896
rect 3567 2894 3573 2895
rect 3671 2895 3672 2896
rect 3676 2895 3677 2899
rect 3671 2894 3677 2895
rect 3759 2899 3765 2900
rect 3759 2895 3760 2899
rect 3764 2898 3765 2899
rect 3863 2899 3869 2900
rect 3863 2898 3864 2899
rect 3764 2896 3864 2898
rect 3764 2895 3765 2896
rect 3759 2894 3765 2895
rect 3863 2895 3864 2896
rect 3868 2895 3869 2899
rect 3863 2894 3869 2895
rect 3871 2899 3877 2900
rect 3871 2895 3872 2899
rect 3876 2898 3877 2899
rect 3951 2899 3957 2900
rect 3951 2898 3952 2899
rect 3876 2896 3952 2898
rect 3876 2895 3877 2896
rect 3871 2894 3877 2895
rect 3951 2895 3952 2896
rect 3956 2895 3957 2899
rect 3951 2894 3957 2895
rect 2110 2891 2116 2892
rect 2110 2887 2111 2891
rect 2115 2887 2116 2891
rect 2110 2886 2116 2887
rect 2278 2891 2284 2892
rect 2278 2887 2279 2891
rect 2283 2887 2284 2891
rect 2278 2886 2284 2887
rect 2486 2891 2492 2892
rect 2486 2887 2487 2891
rect 2491 2887 2492 2891
rect 2486 2886 2492 2887
rect 2694 2891 2700 2892
rect 2694 2887 2695 2891
rect 2699 2887 2700 2891
rect 2694 2886 2700 2887
rect 2902 2891 2908 2892
rect 2902 2887 2903 2891
rect 2907 2887 2908 2891
rect 2902 2886 2908 2887
rect 3110 2891 3116 2892
rect 3110 2887 3111 2891
rect 3115 2887 3116 2891
rect 3110 2886 3116 2887
rect 3302 2891 3308 2892
rect 3302 2887 3303 2891
rect 3307 2887 3308 2891
rect 3302 2886 3308 2887
rect 3494 2891 3500 2892
rect 3494 2887 3495 2891
rect 3499 2887 3500 2891
rect 3494 2886 3500 2887
rect 3686 2891 3692 2892
rect 3686 2887 3687 2891
rect 3691 2887 3692 2891
rect 3686 2886 3692 2887
rect 3878 2891 3884 2892
rect 3878 2887 3879 2891
rect 3883 2887 3884 2891
rect 3878 2886 3884 2887
rect 222 2883 229 2884
rect 222 2879 223 2883
rect 228 2879 229 2883
rect 359 2883 365 2884
rect 359 2882 360 2883
rect 222 2878 229 2879
rect 232 2880 360 2882
rect 150 2875 156 2876
rect 150 2871 151 2875
rect 155 2871 156 2875
rect 150 2870 156 2871
rect 232 2866 234 2880
rect 359 2879 360 2880
rect 364 2879 365 2883
rect 519 2883 525 2884
rect 519 2882 520 2883
rect 359 2878 365 2879
rect 428 2880 520 2882
rect 286 2875 292 2876
rect 286 2871 287 2875
rect 291 2871 292 2875
rect 286 2870 292 2871
rect 428 2866 430 2880
rect 519 2879 520 2880
rect 524 2879 525 2883
rect 519 2878 525 2879
rect 671 2883 677 2884
rect 671 2879 672 2883
rect 676 2882 677 2883
rect 743 2883 749 2884
rect 743 2882 744 2883
rect 676 2880 744 2882
rect 676 2879 677 2880
rect 671 2878 677 2879
rect 743 2879 744 2880
rect 748 2879 749 2883
rect 743 2878 749 2879
rect 831 2883 837 2884
rect 831 2879 832 2883
rect 836 2882 837 2883
rect 911 2883 917 2884
rect 911 2882 912 2883
rect 836 2880 912 2882
rect 836 2879 837 2880
rect 831 2878 837 2879
rect 911 2879 912 2880
rect 916 2879 917 2883
rect 911 2878 917 2879
rect 982 2883 988 2884
rect 982 2879 983 2883
rect 987 2882 988 2883
rect 999 2883 1005 2884
rect 999 2882 1000 2883
rect 987 2880 1000 2882
rect 987 2879 988 2880
rect 982 2878 988 2879
rect 999 2879 1000 2880
rect 1004 2879 1005 2883
rect 999 2878 1005 2879
rect 1034 2883 1040 2884
rect 1034 2879 1035 2883
rect 1039 2882 1040 2883
rect 1087 2883 1093 2884
rect 1087 2882 1088 2883
rect 1039 2880 1088 2882
rect 1039 2879 1040 2880
rect 1034 2878 1040 2879
rect 1087 2879 1088 2880
rect 1092 2879 1093 2883
rect 1087 2878 1093 2879
rect 1175 2883 1181 2884
rect 1175 2879 1176 2883
rect 1180 2882 1181 2883
rect 1271 2883 1277 2884
rect 1271 2882 1272 2883
rect 1180 2880 1272 2882
rect 1180 2879 1181 2880
rect 1175 2878 1181 2879
rect 1271 2879 1272 2880
rect 1276 2879 1277 2883
rect 1271 2878 1277 2879
rect 1359 2883 1365 2884
rect 1359 2879 1360 2883
rect 1364 2882 1365 2883
rect 1463 2883 1469 2884
rect 1463 2882 1464 2883
rect 1364 2880 1464 2882
rect 1364 2879 1365 2880
rect 1359 2878 1365 2879
rect 1463 2879 1464 2880
rect 1468 2879 1469 2883
rect 1463 2878 1469 2879
rect 1534 2883 1540 2884
rect 1534 2879 1535 2883
rect 1539 2882 1540 2883
rect 1551 2883 1557 2884
rect 1551 2882 1552 2883
rect 1539 2880 1552 2882
rect 1539 2879 1540 2880
rect 1534 2878 1540 2879
rect 1551 2879 1552 2880
rect 1556 2879 1557 2883
rect 1551 2878 1557 2879
rect 1718 2883 1724 2884
rect 1718 2879 1719 2883
rect 1723 2882 1724 2883
rect 1743 2883 1749 2884
rect 1743 2882 1744 2883
rect 1723 2880 1744 2882
rect 1723 2879 1724 2880
rect 1718 2878 1724 2879
rect 1743 2879 1744 2880
rect 1748 2879 1749 2883
rect 2230 2883 2236 2884
rect 2230 2882 2231 2883
rect 2161 2880 2231 2882
rect 1743 2878 1749 2879
rect 2230 2879 2231 2880
rect 2235 2879 2236 2883
rect 3286 2883 3292 2884
rect 3286 2882 3287 2883
rect 3161 2880 3287 2882
rect 2230 2878 2236 2879
rect 3286 2879 3287 2880
rect 3291 2879 3292 2883
rect 3286 2878 3292 2879
rect 446 2875 452 2876
rect 446 2871 447 2875
rect 451 2871 452 2875
rect 446 2870 452 2871
rect 598 2875 604 2876
rect 598 2871 599 2875
rect 603 2871 604 2875
rect 598 2870 604 2871
rect 758 2875 764 2876
rect 758 2871 759 2875
rect 763 2871 764 2875
rect 758 2870 764 2871
rect 926 2875 932 2876
rect 926 2871 927 2875
rect 931 2871 932 2875
rect 926 2870 932 2871
rect 1102 2875 1108 2876
rect 1102 2871 1103 2875
rect 1107 2871 1108 2875
rect 1102 2870 1108 2871
rect 1286 2875 1292 2876
rect 1286 2871 1287 2875
rect 1291 2871 1292 2875
rect 1286 2870 1292 2871
rect 1478 2875 1484 2876
rect 1478 2871 1479 2875
rect 1483 2871 1484 2875
rect 1478 2870 1484 2871
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 2070 2872 2076 2873
rect 2070 2868 2071 2872
rect 2075 2868 2076 2872
rect 514 2867 520 2868
rect 2070 2867 2076 2868
rect 3990 2872 3996 2873
rect 3990 2868 3991 2872
rect 3995 2868 3996 2872
rect 3990 2867 3996 2868
rect 514 2866 515 2867
rect 201 2864 234 2866
rect 337 2864 430 2866
rect 497 2864 515 2866
rect 514 2863 515 2864
rect 519 2863 520 2867
rect 514 2862 520 2863
rect 590 2863 596 2864
rect 590 2859 591 2863
rect 595 2859 596 2863
rect 590 2858 596 2859
rect 1694 2863 1700 2864
rect 1694 2859 1695 2863
rect 1699 2859 1700 2863
rect 1694 2858 1700 2859
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 110 2851 116 2852
rect 2030 2856 2036 2857
rect 2030 2852 2031 2856
rect 2035 2852 2036 2856
rect 2030 2851 2036 2852
rect 2070 2855 2076 2856
rect 2070 2851 2071 2855
rect 2075 2851 2076 2855
rect 3990 2855 3996 2856
rect 3990 2851 3991 2855
rect 3995 2851 3996 2855
rect 2070 2850 2076 2851
rect 2110 2850 2116 2851
rect 2110 2846 2111 2850
rect 2115 2846 2116 2850
rect 2110 2845 2116 2846
rect 2278 2850 2284 2851
rect 2278 2846 2279 2850
rect 2283 2846 2284 2850
rect 2278 2845 2284 2846
rect 2486 2850 2492 2851
rect 2486 2846 2487 2850
rect 2491 2846 2492 2850
rect 2486 2845 2492 2846
rect 2694 2850 2700 2851
rect 2694 2846 2695 2850
rect 2699 2846 2700 2850
rect 2694 2845 2700 2846
rect 2902 2850 2908 2851
rect 2902 2846 2903 2850
rect 2907 2846 2908 2850
rect 2902 2845 2908 2846
rect 3110 2850 3116 2851
rect 3110 2846 3111 2850
rect 3115 2846 3116 2850
rect 3110 2845 3116 2846
rect 3302 2850 3308 2851
rect 3302 2846 3303 2850
rect 3307 2846 3308 2850
rect 3302 2845 3308 2846
rect 3494 2850 3500 2851
rect 3494 2846 3495 2850
rect 3499 2846 3500 2850
rect 3494 2845 3500 2846
rect 3686 2850 3692 2851
rect 3686 2846 3687 2850
rect 3691 2846 3692 2850
rect 3686 2845 3692 2846
rect 3878 2850 3884 2851
rect 3990 2850 3996 2851
rect 3878 2846 3879 2850
rect 3883 2846 3884 2850
rect 3878 2845 3884 2846
rect 110 2839 116 2840
rect 110 2835 111 2839
rect 115 2835 116 2839
rect 2030 2839 2036 2840
rect 2030 2835 2031 2839
rect 2035 2835 2036 2839
rect 110 2834 116 2835
rect 150 2834 156 2835
rect 150 2830 151 2834
rect 155 2830 156 2834
rect 150 2829 156 2830
rect 286 2834 292 2835
rect 286 2830 287 2834
rect 291 2830 292 2834
rect 286 2829 292 2830
rect 446 2834 452 2835
rect 446 2830 447 2834
rect 451 2830 452 2834
rect 446 2829 452 2830
rect 598 2834 604 2835
rect 598 2830 599 2834
rect 603 2830 604 2834
rect 598 2829 604 2830
rect 758 2834 764 2835
rect 758 2830 759 2834
rect 763 2830 764 2834
rect 758 2829 764 2830
rect 926 2834 932 2835
rect 926 2830 927 2834
rect 931 2830 932 2834
rect 926 2829 932 2830
rect 1102 2834 1108 2835
rect 1102 2830 1103 2834
rect 1107 2830 1108 2834
rect 1102 2829 1108 2830
rect 1286 2834 1292 2835
rect 1286 2830 1287 2834
rect 1291 2830 1292 2834
rect 1286 2829 1292 2830
rect 1478 2834 1484 2835
rect 1478 2830 1479 2834
rect 1483 2830 1484 2834
rect 1478 2829 1484 2830
rect 1670 2834 1676 2835
rect 2030 2834 2036 2835
rect 1670 2830 1671 2834
rect 1675 2830 1676 2834
rect 1670 2829 1676 2830
rect 3286 2823 3292 2824
rect 3286 2819 3287 2823
rect 3291 2822 3292 2823
rect 3838 2823 3844 2824
rect 3838 2822 3839 2823
rect 3291 2820 3839 2822
rect 3291 2819 3292 2820
rect 3286 2818 3292 2819
rect 3838 2819 3839 2820
rect 3843 2819 3844 2823
rect 3838 2818 3844 2819
rect 2142 2806 2148 2807
rect 2142 2802 2143 2806
rect 2147 2802 2148 2806
rect 2070 2801 2076 2802
rect 2142 2801 2148 2802
rect 2318 2806 2324 2807
rect 2318 2802 2319 2806
rect 2323 2802 2324 2806
rect 2318 2801 2324 2802
rect 2502 2806 2508 2807
rect 2502 2802 2503 2806
rect 2507 2802 2508 2806
rect 2502 2801 2508 2802
rect 2694 2806 2700 2807
rect 2694 2802 2695 2806
rect 2699 2802 2700 2806
rect 2694 2801 2700 2802
rect 2886 2806 2892 2807
rect 2886 2802 2887 2806
rect 2891 2802 2892 2806
rect 2886 2801 2892 2802
rect 3078 2806 3084 2807
rect 3078 2802 3079 2806
rect 3083 2802 3084 2806
rect 3078 2801 3084 2802
rect 3262 2806 3268 2807
rect 3262 2802 3263 2806
rect 3267 2802 3268 2806
rect 3262 2801 3268 2802
rect 3438 2806 3444 2807
rect 3438 2802 3439 2806
rect 3443 2802 3444 2806
rect 3438 2801 3444 2802
rect 3614 2806 3620 2807
rect 3614 2802 3615 2806
rect 3619 2802 3620 2806
rect 3614 2801 3620 2802
rect 3790 2806 3796 2807
rect 3790 2802 3791 2806
rect 3795 2802 3796 2806
rect 3790 2801 3796 2802
rect 3990 2801 3996 2802
rect 2070 2797 2071 2801
rect 2075 2797 2076 2801
rect 2070 2796 2076 2797
rect 3990 2797 3991 2801
rect 3995 2797 3996 2801
rect 3990 2796 3996 2797
rect 150 2790 156 2791
rect 150 2786 151 2790
rect 155 2786 156 2790
rect 110 2785 116 2786
rect 150 2785 156 2786
rect 318 2790 324 2791
rect 318 2786 319 2790
rect 323 2786 324 2790
rect 318 2785 324 2786
rect 502 2790 508 2791
rect 502 2786 503 2790
rect 507 2786 508 2790
rect 502 2785 508 2786
rect 686 2790 692 2791
rect 686 2786 687 2790
rect 691 2786 692 2790
rect 686 2785 692 2786
rect 870 2790 876 2791
rect 870 2786 871 2790
rect 875 2786 876 2790
rect 870 2785 876 2786
rect 1054 2790 1060 2791
rect 1054 2786 1055 2790
rect 1059 2786 1060 2790
rect 1054 2785 1060 2786
rect 1238 2790 1244 2791
rect 1238 2786 1239 2790
rect 1243 2786 1244 2790
rect 1238 2785 1244 2786
rect 1430 2790 1436 2791
rect 1430 2786 1431 2790
rect 1435 2786 1436 2790
rect 1430 2785 1436 2786
rect 1630 2790 1636 2791
rect 1630 2786 1631 2790
rect 1635 2786 1636 2790
rect 1630 2785 1636 2786
rect 1830 2790 1836 2791
rect 1830 2786 1831 2790
rect 1835 2786 1836 2790
rect 1830 2785 1836 2786
rect 2030 2785 2036 2786
rect 110 2781 111 2785
rect 115 2781 116 2785
rect 110 2780 116 2781
rect 2030 2781 2031 2785
rect 2035 2781 2036 2785
rect 2030 2780 2036 2781
rect 2070 2784 2076 2785
rect 2070 2780 2071 2784
rect 2075 2780 2076 2784
rect 2070 2779 2076 2780
rect 3990 2784 3996 2785
rect 3990 2780 3991 2784
rect 3995 2780 3996 2784
rect 3990 2779 3996 2780
rect 2166 2775 2172 2776
rect 2166 2771 2167 2775
rect 2171 2771 2172 2775
rect 2678 2775 2684 2776
rect 2678 2774 2679 2775
rect 2553 2772 2679 2774
rect 2166 2770 2172 2771
rect 2678 2771 2679 2772
rect 2683 2771 2684 2775
rect 2870 2775 2876 2776
rect 2870 2774 2871 2775
rect 2745 2772 2871 2774
rect 2678 2770 2684 2771
rect 2870 2771 2871 2772
rect 2875 2771 2876 2775
rect 2974 2775 2980 2776
rect 2974 2774 2975 2775
rect 2937 2772 2975 2774
rect 2870 2770 2876 2771
rect 2974 2771 2975 2772
rect 2979 2771 2980 2775
rect 3246 2775 3252 2776
rect 3246 2774 3247 2775
rect 3129 2772 3247 2774
rect 2974 2770 2980 2771
rect 3246 2771 3247 2772
rect 3251 2771 3252 2775
rect 3246 2770 3252 2771
rect 110 2768 116 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 2030 2768 2036 2769
rect 2030 2764 2031 2768
rect 2035 2764 2036 2768
rect 2030 2763 2036 2764
rect 2142 2765 2148 2766
rect 2142 2761 2143 2765
rect 2147 2761 2148 2765
rect 2318 2765 2324 2766
rect 2142 2760 2148 2761
rect 2230 2763 2236 2764
rect 222 2759 228 2760
rect 222 2758 223 2759
rect 201 2756 223 2758
rect 222 2755 223 2756
rect 227 2755 228 2759
rect 670 2759 676 2760
rect 670 2758 671 2759
rect 553 2756 671 2758
rect 222 2754 228 2755
rect 670 2755 671 2756
rect 675 2755 676 2759
rect 1222 2759 1228 2760
rect 1222 2758 1223 2759
rect 737 2756 814 2758
rect 1105 2756 1223 2758
rect 670 2754 676 2755
rect 150 2749 156 2750
rect 150 2745 151 2749
rect 155 2745 156 2749
rect 150 2744 156 2745
rect 318 2749 324 2750
rect 318 2745 319 2749
rect 323 2745 324 2749
rect 318 2744 324 2745
rect 502 2749 508 2750
rect 502 2745 503 2749
rect 507 2745 508 2749
rect 502 2744 508 2745
rect 686 2749 692 2750
rect 686 2745 687 2749
rect 691 2745 692 2749
rect 686 2744 692 2745
rect 812 2746 814 2756
rect 1222 2755 1223 2756
rect 1227 2755 1228 2759
rect 1414 2759 1420 2760
rect 1414 2758 1415 2759
rect 1289 2756 1415 2758
rect 1222 2754 1228 2755
rect 1414 2755 1415 2756
rect 1419 2755 1420 2759
rect 1534 2759 1540 2760
rect 1534 2758 1535 2759
rect 1481 2756 1535 2758
rect 1414 2754 1420 2755
rect 1534 2755 1535 2756
rect 1539 2755 1540 2759
rect 1814 2759 1820 2760
rect 1814 2758 1815 2759
rect 1681 2756 1815 2758
rect 1534 2754 1540 2755
rect 1814 2755 1815 2756
rect 1819 2755 1820 2759
rect 1902 2759 1908 2760
rect 1902 2758 1903 2759
rect 1881 2756 1903 2758
rect 1814 2754 1820 2755
rect 1902 2755 1903 2756
rect 1907 2755 1908 2759
rect 2230 2759 2231 2763
rect 2235 2762 2236 2763
rect 2235 2760 2314 2762
rect 2318 2761 2319 2765
rect 2323 2761 2324 2765
rect 2318 2760 2324 2761
rect 2502 2765 2508 2766
rect 2502 2761 2503 2765
rect 2507 2761 2508 2765
rect 2502 2760 2508 2761
rect 2694 2765 2700 2766
rect 2694 2761 2695 2765
rect 2699 2761 2700 2765
rect 2694 2760 2700 2761
rect 2886 2765 2892 2766
rect 2886 2761 2887 2765
rect 2891 2761 2892 2765
rect 2886 2760 2892 2761
rect 3078 2765 3084 2766
rect 3078 2761 3079 2765
rect 3083 2761 3084 2765
rect 3078 2760 3084 2761
rect 3262 2765 3268 2766
rect 3262 2761 3263 2765
rect 3267 2761 3268 2765
rect 3262 2760 3268 2761
rect 3438 2765 3444 2766
rect 3438 2761 3439 2765
rect 3443 2761 3444 2765
rect 3438 2760 3444 2761
rect 3614 2765 3620 2766
rect 3614 2761 3615 2765
rect 3619 2761 3620 2765
rect 3614 2760 3620 2761
rect 3790 2765 3796 2766
rect 3790 2761 3791 2765
rect 3795 2761 3796 2765
rect 3790 2760 3796 2761
rect 2235 2759 2236 2760
rect 2230 2758 2236 2759
rect 1902 2754 1908 2755
rect 2215 2755 2221 2756
rect 2215 2751 2216 2755
rect 2220 2754 2221 2755
rect 2303 2755 2309 2756
rect 2303 2754 2304 2755
rect 2220 2752 2304 2754
rect 2220 2751 2221 2752
rect 2215 2750 2221 2751
rect 2303 2751 2304 2752
rect 2308 2751 2309 2755
rect 2312 2754 2314 2760
rect 2391 2755 2397 2756
rect 2391 2754 2392 2755
rect 2312 2752 2392 2754
rect 2303 2750 2309 2751
rect 2391 2751 2392 2752
rect 2396 2751 2397 2755
rect 2391 2750 2397 2751
rect 2518 2755 2524 2756
rect 2518 2751 2519 2755
rect 2523 2754 2524 2755
rect 2575 2755 2581 2756
rect 2575 2754 2576 2755
rect 2523 2752 2576 2754
rect 2523 2751 2524 2752
rect 2518 2750 2524 2751
rect 2575 2751 2576 2752
rect 2580 2751 2581 2755
rect 2575 2750 2581 2751
rect 2678 2755 2684 2756
rect 2678 2751 2679 2755
rect 2683 2754 2684 2755
rect 2767 2755 2773 2756
rect 2767 2754 2768 2755
rect 2683 2752 2768 2754
rect 2683 2751 2684 2752
rect 2678 2750 2684 2751
rect 2767 2751 2768 2752
rect 2772 2751 2773 2755
rect 2767 2750 2773 2751
rect 2870 2755 2876 2756
rect 2870 2751 2871 2755
rect 2875 2754 2876 2755
rect 2959 2755 2965 2756
rect 2959 2754 2960 2755
rect 2875 2752 2960 2754
rect 2875 2751 2876 2752
rect 2870 2750 2876 2751
rect 2959 2751 2960 2752
rect 2964 2751 2965 2755
rect 2959 2750 2965 2751
rect 3151 2755 3157 2756
rect 3151 2751 3152 2755
rect 3156 2754 3157 2755
rect 3247 2755 3253 2756
rect 3247 2754 3248 2755
rect 3156 2752 3248 2754
rect 3156 2751 3157 2752
rect 3151 2750 3157 2751
rect 3247 2751 3248 2752
rect 3252 2751 3253 2755
rect 3247 2750 3253 2751
rect 3335 2755 3341 2756
rect 3335 2751 3336 2755
rect 3340 2754 3341 2755
rect 3423 2755 3429 2756
rect 3423 2754 3424 2755
rect 3340 2752 3424 2754
rect 3340 2751 3341 2752
rect 3335 2750 3341 2751
rect 3423 2751 3424 2752
rect 3428 2751 3429 2755
rect 3423 2750 3429 2751
rect 3511 2755 3517 2756
rect 3511 2751 3512 2755
rect 3516 2754 3517 2755
rect 3599 2755 3605 2756
rect 3599 2754 3600 2755
rect 3516 2752 3600 2754
rect 3516 2751 3517 2752
rect 3511 2750 3517 2751
rect 3599 2751 3600 2752
rect 3604 2751 3605 2755
rect 3599 2750 3605 2751
rect 3687 2755 3693 2756
rect 3687 2751 3688 2755
rect 3692 2754 3693 2755
rect 3775 2755 3781 2756
rect 3775 2754 3776 2755
rect 3692 2752 3776 2754
rect 3692 2751 3693 2752
rect 3687 2750 3693 2751
rect 3775 2751 3776 2752
rect 3780 2751 3781 2755
rect 3775 2750 3781 2751
rect 3838 2755 3844 2756
rect 3838 2751 3839 2755
rect 3843 2754 3844 2755
rect 3863 2755 3869 2756
rect 3863 2754 3864 2755
rect 3843 2752 3864 2754
rect 3843 2751 3844 2752
rect 3838 2750 3844 2751
rect 3863 2751 3864 2752
rect 3868 2751 3869 2755
rect 3863 2750 3869 2751
rect 870 2749 876 2750
rect 812 2744 866 2746
rect 870 2745 871 2749
rect 875 2745 876 2749
rect 870 2744 876 2745
rect 1054 2749 1060 2750
rect 1054 2745 1055 2749
rect 1059 2745 1060 2749
rect 1054 2744 1060 2745
rect 1238 2749 1244 2750
rect 1238 2745 1239 2749
rect 1243 2745 1244 2749
rect 1238 2744 1244 2745
rect 1430 2749 1436 2750
rect 1430 2745 1431 2749
rect 1435 2745 1436 2749
rect 1430 2744 1436 2745
rect 1630 2749 1636 2750
rect 1630 2745 1631 2749
rect 1635 2745 1636 2749
rect 1630 2744 1636 2745
rect 1830 2749 1836 2750
rect 1830 2745 1831 2749
rect 1835 2745 1836 2749
rect 1830 2744 1836 2745
rect 223 2739 229 2740
rect 223 2735 224 2739
rect 228 2738 229 2739
rect 303 2739 309 2740
rect 303 2738 304 2739
rect 228 2736 304 2738
rect 228 2735 229 2736
rect 223 2734 229 2735
rect 303 2735 304 2736
rect 308 2735 309 2739
rect 303 2734 309 2735
rect 390 2739 397 2740
rect 390 2735 391 2739
rect 396 2735 397 2739
rect 390 2734 397 2735
rect 575 2739 581 2740
rect 575 2735 576 2739
rect 580 2738 581 2739
rect 590 2739 596 2740
rect 590 2738 591 2739
rect 580 2736 591 2738
rect 580 2735 581 2736
rect 575 2734 581 2735
rect 590 2735 591 2736
rect 595 2735 596 2739
rect 590 2734 596 2735
rect 670 2739 676 2740
rect 670 2735 671 2739
rect 675 2738 676 2739
rect 759 2739 765 2740
rect 759 2738 760 2739
rect 675 2736 760 2738
rect 675 2735 676 2736
rect 670 2734 676 2735
rect 759 2735 760 2736
rect 764 2735 765 2739
rect 759 2734 765 2735
rect 855 2739 861 2740
rect 855 2735 856 2739
rect 860 2735 861 2739
rect 864 2738 866 2744
rect 943 2739 949 2740
rect 943 2738 944 2739
rect 864 2736 944 2738
rect 855 2734 861 2735
rect 943 2735 944 2736
rect 948 2735 949 2739
rect 943 2734 949 2735
rect 1046 2739 1052 2740
rect 1046 2735 1047 2739
rect 1051 2738 1052 2739
rect 1127 2739 1133 2740
rect 1127 2738 1128 2739
rect 1051 2736 1128 2738
rect 1051 2735 1052 2736
rect 1046 2734 1052 2735
rect 1127 2735 1128 2736
rect 1132 2735 1133 2739
rect 1127 2734 1133 2735
rect 1222 2739 1228 2740
rect 1222 2735 1223 2739
rect 1227 2738 1228 2739
rect 1311 2739 1317 2740
rect 1311 2738 1312 2739
rect 1227 2736 1312 2738
rect 1227 2735 1228 2736
rect 1222 2734 1228 2735
rect 1311 2735 1312 2736
rect 1316 2735 1317 2739
rect 1311 2734 1317 2735
rect 1414 2739 1420 2740
rect 1414 2735 1415 2739
rect 1419 2738 1420 2739
rect 1503 2739 1509 2740
rect 1503 2738 1504 2739
rect 1419 2736 1504 2738
rect 1419 2735 1420 2736
rect 1414 2734 1420 2735
rect 1503 2735 1504 2736
rect 1508 2735 1509 2739
rect 1503 2734 1509 2735
rect 1694 2739 1700 2740
rect 1694 2735 1695 2739
rect 1699 2738 1700 2739
rect 1703 2739 1709 2740
rect 1703 2738 1704 2739
rect 1699 2736 1704 2738
rect 1699 2735 1700 2736
rect 1694 2734 1700 2735
rect 1703 2735 1704 2736
rect 1708 2735 1709 2739
rect 1703 2734 1709 2735
rect 1814 2739 1820 2740
rect 1814 2735 1815 2739
rect 1819 2738 1820 2739
rect 1903 2739 1909 2740
rect 1903 2738 1904 2739
rect 1819 2736 1904 2738
rect 1819 2735 1820 2736
rect 1814 2734 1820 2735
rect 1903 2735 1904 2736
rect 1908 2735 1909 2739
rect 1903 2734 1909 2735
rect 3246 2739 3252 2740
rect 3246 2735 3247 2739
rect 3251 2738 3252 2739
rect 3251 2736 3681 2738
rect 3251 2735 3252 2736
rect 3246 2734 3252 2735
rect 255 2724 261 2725
rect 856 2724 858 2734
rect 2166 2731 2172 2732
rect 2166 2727 2167 2731
rect 2171 2730 2172 2731
rect 2183 2731 2189 2732
rect 2183 2730 2184 2731
rect 2171 2728 2184 2730
rect 2171 2727 2172 2728
rect 2166 2726 2172 2727
rect 2183 2727 2184 2728
rect 2188 2727 2189 2731
rect 2351 2731 2357 2732
rect 2351 2730 2352 2731
rect 2183 2726 2189 2727
rect 2228 2728 2352 2730
rect 246 2723 252 2724
rect 246 2719 247 2723
rect 251 2722 252 2723
rect 255 2722 256 2724
rect 251 2720 256 2722
rect 260 2720 261 2724
rect 455 2723 461 2724
rect 455 2722 456 2723
rect 251 2719 252 2720
rect 255 2719 261 2720
rect 319 2720 456 2722
rect 246 2718 252 2719
rect 182 2715 188 2716
rect 182 2711 183 2715
rect 187 2711 188 2715
rect 182 2710 188 2711
rect 319 2706 321 2720
rect 455 2719 456 2720
rect 460 2719 461 2723
rect 455 2718 461 2719
rect 655 2723 661 2724
rect 655 2719 656 2723
rect 660 2722 661 2723
rect 767 2723 773 2724
rect 767 2722 768 2723
rect 660 2720 768 2722
rect 660 2719 661 2720
rect 655 2718 661 2719
rect 767 2719 768 2720
rect 772 2719 773 2723
rect 767 2718 773 2719
rect 855 2723 861 2724
rect 855 2719 856 2723
rect 860 2719 861 2723
rect 855 2718 861 2719
rect 1055 2723 1061 2724
rect 1055 2719 1056 2723
rect 1060 2722 1061 2723
rect 1183 2723 1189 2724
rect 1183 2722 1184 2723
rect 1060 2720 1184 2722
rect 1060 2719 1061 2720
rect 1055 2718 1061 2719
rect 1183 2719 1184 2720
rect 1188 2719 1189 2723
rect 1183 2718 1189 2719
rect 1271 2723 1277 2724
rect 1271 2719 1272 2723
rect 1276 2722 1277 2723
rect 1399 2723 1405 2724
rect 1399 2722 1400 2723
rect 1276 2720 1400 2722
rect 1276 2719 1277 2720
rect 1271 2718 1277 2719
rect 1399 2719 1400 2720
rect 1404 2719 1405 2723
rect 1399 2718 1405 2719
rect 1487 2723 1493 2724
rect 1487 2719 1488 2723
rect 1492 2722 1493 2723
rect 1623 2723 1629 2724
rect 1623 2722 1624 2723
rect 1492 2720 1624 2722
rect 1492 2719 1493 2720
rect 1487 2718 1493 2719
rect 1623 2719 1624 2720
rect 1628 2719 1629 2723
rect 1623 2718 1629 2719
rect 1646 2723 1652 2724
rect 1646 2719 1647 2723
rect 1651 2722 1652 2723
rect 1711 2723 1717 2724
rect 1711 2722 1712 2723
rect 1651 2720 1712 2722
rect 1651 2719 1652 2720
rect 1646 2718 1652 2719
rect 1711 2719 1712 2720
rect 1716 2719 1717 2723
rect 1711 2718 1717 2719
rect 1902 2723 1908 2724
rect 1902 2719 1903 2723
rect 1907 2722 1908 2723
rect 1943 2723 1949 2724
rect 1943 2722 1944 2723
rect 1907 2720 1944 2722
rect 1907 2719 1908 2720
rect 1902 2718 1908 2719
rect 1943 2719 1944 2720
rect 1948 2719 1949 2723
rect 1943 2718 1949 2719
rect 2110 2723 2116 2724
rect 2110 2719 2111 2723
rect 2115 2719 2116 2723
rect 2110 2718 2116 2719
rect 382 2715 388 2716
rect 382 2711 383 2715
rect 387 2711 388 2715
rect 382 2710 388 2711
rect 582 2715 588 2716
rect 582 2711 583 2715
rect 587 2711 588 2715
rect 582 2710 588 2711
rect 782 2715 788 2716
rect 782 2711 783 2715
rect 787 2711 788 2715
rect 782 2710 788 2711
rect 982 2715 988 2716
rect 982 2711 983 2715
rect 987 2711 988 2715
rect 982 2710 988 2711
rect 1198 2715 1204 2716
rect 1198 2711 1199 2715
rect 1203 2711 1204 2715
rect 1198 2710 1204 2711
rect 1414 2715 1420 2716
rect 1414 2711 1415 2715
rect 1419 2711 1420 2715
rect 1414 2710 1420 2711
rect 1638 2715 1644 2716
rect 1638 2711 1639 2715
rect 1643 2711 1644 2715
rect 1638 2710 1644 2711
rect 1870 2715 1876 2716
rect 1870 2711 1871 2715
rect 1875 2711 1876 2715
rect 2228 2714 2230 2728
rect 2351 2727 2352 2728
rect 2356 2727 2357 2731
rect 2351 2726 2357 2727
rect 2527 2731 2533 2732
rect 2527 2727 2528 2731
rect 2532 2730 2533 2731
rect 2623 2731 2629 2732
rect 2623 2730 2624 2731
rect 2532 2728 2624 2730
rect 2532 2727 2533 2728
rect 2527 2726 2533 2727
rect 2623 2727 2624 2728
rect 2628 2727 2629 2731
rect 2623 2726 2629 2727
rect 2711 2731 2717 2732
rect 2711 2727 2712 2731
rect 2716 2730 2717 2731
rect 2799 2731 2805 2732
rect 2799 2730 2800 2731
rect 2716 2728 2800 2730
rect 2716 2727 2717 2728
rect 2711 2726 2717 2727
rect 2799 2727 2800 2728
rect 2804 2727 2805 2731
rect 2799 2726 2805 2727
rect 2862 2731 2868 2732
rect 2862 2727 2863 2731
rect 2867 2730 2868 2731
rect 2887 2731 2893 2732
rect 2887 2730 2888 2731
rect 2867 2728 2888 2730
rect 2867 2727 2868 2728
rect 2862 2726 2868 2727
rect 2887 2727 2888 2728
rect 2892 2727 2893 2731
rect 2887 2726 2893 2727
rect 3055 2731 3061 2732
rect 3055 2727 3056 2731
rect 3060 2730 3061 2731
rect 3127 2731 3133 2732
rect 3127 2730 3128 2731
rect 3060 2728 3128 2730
rect 3060 2727 3061 2728
rect 3055 2726 3061 2727
rect 3127 2727 3128 2728
rect 3132 2727 3133 2731
rect 3127 2726 3133 2727
rect 3215 2731 3221 2732
rect 3215 2727 3216 2731
rect 3220 2730 3221 2731
rect 3287 2731 3293 2732
rect 3287 2730 3288 2731
rect 3220 2728 3288 2730
rect 3220 2727 3221 2728
rect 3215 2726 3221 2727
rect 3287 2727 3288 2728
rect 3292 2727 3293 2731
rect 3287 2726 3293 2727
rect 3375 2731 3381 2732
rect 3375 2727 3376 2731
rect 3380 2730 3381 2731
rect 3447 2731 3453 2732
rect 3447 2730 3448 2731
rect 3380 2728 3448 2730
rect 3380 2727 3381 2728
rect 3375 2726 3381 2727
rect 3447 2727 3448 2728
rect 3452 2727 3453 2731
rect 3447 2726 3453 2727
rect 3535 2731 3541 2732
rect 3535 2727 3536 2731
rect 3540 2730 3541 2731
rect 3607 2731 3613 2732
rect 3607 2730 3608 2731
rect 3540 2728 3608 2730
rect 3540 2727 3541 2728
rect 3535 2726 3541 2727
rect 3607 2727 3608 2728
rect 3612 2727 3613 2731
rect 3679 2730 3681 2736
rect 3695 2731 3701 2732
rect 3695 2730 3696 2731
rect 3679 2728 3696 2730
rect 3607 2726 3613 2727
rect 3695 2727 3696 2728
rect 3700 2727 3701 2731
rect 3695 2726 3701 2727
rect 2278 2723 2284 2724
rect 2278 2719 2279 2723
rect 2283 2719 2284 2723
rect 2278 2718 2284 2719
rect 2454 2723 2460 2724
rect 2454 2719 2455 2723
rect 2459 2719 2460 2723
rect 2454 2718 2460 2719
rect 2638 2723 2644 2724
rect 2638 2719 2639 2723
rect 2643 2719 2644 2723
rect 2638 2718 2644 2719
rect 2814 2723 2820 2724
rect 2814 2719 2815 2723
rect 2819 2719 2820 2723
rect 2814 2718 2820 2719
rect 2982 2723 2988 2724
rect 2982 2719 2983 2723
rect 2987 2719 2988 2723
rect 2982 2718 2988 2719
rect 3142 2723 3148 2724
rect 3142 2719 3143 2723
rect 3147 2719 3148 2723
rect 3142 2718 3148 2719
rect 3302 2723 3308 2724
rect 3302 2719 3303 2723
rect 3307 2719 3308 2723
rect 3302 2718 3308 2719
rect 3462 2723 3468 2724
rect 3462 2719 3463 2723
rect 3467 2719 3468 2723
rect 3462 2718 3468 2719
rect 3622 2723 3628 2724
rect 3622 2719 3623 2723
rect 3627 2719 3628 2723
rect 3622 2718 3628 2719
rect 2342 2715 2348 2716
rect 2342 2714 2343 2715
rect 2161 2712 2230 2714
rect 2329 2712 2343 2714
rect 1870 2710 1876 2711
rect 2342 2711 2343 2712
rect 2347 2711 2348 2715
rect 2518 2715 2524 2716
rect 2518 2714 2519 2715
rect 2505 2712 2519 2714
rect 2342 2710 2348 2711
rect 2518 2711 2519 2712
rect 2523 2711 2524 2715
rect 3126 2715 3132 2716
rect 3126 2714 3127 2715
rect 3033 2712 3127 2714
rect 2518 2710 2524 2711
rect 3126 2711 3127 2712
rect 3131 2711 3132 2715
rect 3126 2710 3132 2711
rect 670 2707 676 2708
rect 670 2706 671 2707
rect 233 2704 321 2706
rect 633 2704 671 2706
rect 390 2703 396 2704
rect 390 2699 391 2703
rect 395 2699 396 2703
rect 670 2703 671 2704
rect 675 2703 676 2707
rect 1046 2707 1052 2708
rect 1046 2706 1047 2707
rect 1033 2704 1047 2706
rect 670 2702 676 2703
rect 1046 2703 1047 2704
rect 1051 2703 1052 2707
rect 1998 2707 2004 2708
rect 1998 2706 1999 2707
rect 1921 2704 1999 2706
rect 1046 2702 1052 2703
rect 1998 2703 1999 2704
rect 2003 2703 2004 2707
rect 1998 2702 2004 2703
rect 2070 2704 2076 2705
rect 2070 2700 2071 2704
rect 2075 2700 2076 2704
rect 2070 2699 2076 2700
rect 3990 2704 3996 2705
rect 3990 2700 3991 2704
rect 3995 2700 3996 2704
rect 3990 2699 3996 2700
rect 390 2698 396 2699
rect 110 2696 116 2697
rect 110 2692 111 2696
rect 115 2692 116 2696
rect 110 2691 116 2692
rect 2030 2696 2036 2697
rect 2030 2692 2031 2696
rect 2035 2692 2036 2696
rect 2030 2691 2036 2692
rect 2070 2687 2076 2688
rect 2070 2683 2071 2687
rect 2075 2683 2076 2687
rect 3990 2687 3996 2688
rect 3990 2683 3991 2687
rect 3995 2683 3996 2687
rect 2070 2682 2076 2683
rect 2110 2682 2116 2683
rect 110 2679 116 2680
rect 110 2675 111 2679
rect 115 2675 116 2679
rect 2030 2679 2036 2680
rect 2030 2675 2031 2679
rect 2035 2675 2036 2679
rect 2110 2678 2111 2682
rect 2115 2678 2116 2682
rect 2110 2677 2116 2678
rect 2278 2682 2284 2683
rect 2278 2678 2279 2682
rect 2283 2678 2284 2682
rect 2278 2677 2284 2678
rect 2454 2682 2460 2683
rect 2454 2678 2455 2682
rect 2459 2678 2460 2682
rect 2454 2677 2460 2678
rect 2638 2682 2644 2683
rect 2638 2678 2639 2682
rect 2643 2678 2644 2682
rect 2638 2677 2644 2678
rect 2814 2682 2820 2683
rect 2814 2678 2815 2682
rect 2819 2678 2820 2682
rect 2814 2677 2820 2678
rect 2982 2682 2988 2683
rect 2982 2678 2983 2682
rect 2987 2678 2988 2682
rect 2982 2677 2988 2678
rect 3142 2682 3148 2683
rect 3142 2678 3143 2682
rect 3147 2678 3148 2682
rect 3142 2677 3148 2678
rect 3302 2682 3308 2683
rect 3302 2678 3303 2682
rect 3307 2678 3308 2682
rect 3302 2677 3308 2678
rect 3462 2682 3468 2683
rect 3462 2678 3463 2682
rect 3467 2678 3468 2682
rect 3462 2677 3468 2678
rect 3622 2682 3628 2683
rect 3990 2682 3996 2683
rect 3622 2678 3623 2682
rect 3627 2678 3628 2682
rect 3622 2677 3628 2678
rect 110 2674 116 2675
rect 182 2674 188 2675
rect 182 2670 183 2674
rect 187 2670 188 2674
rect 182 2669 188 2670
rect 382 2674 388 2675
rect 382 2670 383 2674
rect 387 2670 388 2674
rect 382 2669 388 2670
rect 582 2674 588 2675
rect 582 2670 583 2674
rect 587 2670 588 2674
rect 582 2669 588 2670
rect 782 2674 788 2675
rect 782 2670 783 2674
rect 787 2670 788 2674
rect 782 2669 788 2670
rect 982 2674 988 2675
rect 982 2670 983 2674
rect 987 2670 988 2674
rect 982 2669 988 2670
rect 1198 2674 1204 2675
rect 1198 2670 1199 2674
rect 1203 2670 1204 2674
rect 1198 2669 1204 2670
rect 1414 2674 1420 2675
rect 1414 2670 1415 2674
rect 1419 2670 1420 2674
rect 1414 2669 1420 2670
rect 1638 2674 1644 2675
rect 1638 2670 1639 2674
rect 1643 2670 1644 2674
rect 1638 2669 1644 2670
rect 1870 2674 1876 2675
rect 2030 2674 2036 2675
rect 1870 2670 1871 2674
rect 1875 2670 1876 2674
rect 1870 2669 1876 2670
rect 2110 2638 2116 2639
rect 254 2634 260 2635
rect 254 2630 255 2634
rect 259 2630 260 2634
rect 110 2629 116 2630
rect 254 2629 260 2630
rect 422 2634 428 2635
rect 422 2630 423 2634
rect 427 2630 428 2634
rect 422 2629 428 2630
rect 598 2634 604 2635
rect 598 2630 599 2634
rect 603 2630 604 2634
rect 598 2629 604 2630
rect 774 2634 780 2635
rect 774 2630 775 2634
rect 779 2630 780 2634
rect 774 2629 780 2630
rect 958 2634 964 2635
rect 958 2630 959 2634
rect 963 2630 964 2634
rect 958 2629 964 2630
rect 1150 2634 1156 2635
rect 1150 2630 1151 2634
rect 1155 2630 1156 2634
rect 1150 2629 1156 2630
rect 1342 2634 1348 2635
rect 1342 2630 1343 2634
rect 1347 2630 1348 2634
rect 1342 2629 1348 2630
rect 1534 2634 1540 2635
rect 1534 2630 1535 2634
rect 1539 2630 1540 2634
rect 1534 2629 1540 2630
rect 1726 2634 1732 2635
rect 1726 2630 1727 2634
rect 1731 2630 1732 2634
rect 1726 2629 1732 2630
rect 1926 2634 1932 2635
rect 2110 2634 2111 2638
rect 2115 2634 2116 2638
rect 1926 2630 1927 2634
rect 1931 2630 1932 2634
rect 2070 2633 2076 2634
rect 2110 2633 2116 2634
rect 2262 2638 2268 2639
rect 2262 2634 2263 2638
rect 2267 2634 2268 2638
rect 2262 2633 2268 2634
rect 2430 2638 2436 2639
rect 2430 2634 2431 2638
rect 2435 2634 2436 2638
rect 2430 2633 2436 2634
rect 2598 2638 2604 2639
rect 2598 2634 2599 2638
rect 2603 2634 2604 2638
rect 2598 2633 2604 2634
rect 2750 2638 2756 2639
rect 2750 2634 2751 2638
rect 2755 2634 2756 2638
rect 2750 2633 2756 2634
rect 2894 2638 2900 2639
rect 2894 2634 2895 2638
rect 2899 2634 2900 2638
rect 2894 2633 2900 2634
rect 3038 2638 3044 2639
rect 3038 2634 3039 2638
rect 3043 2634 3044 2638
rect 3038 2633 3044 2634
rect 3174 2638 3180 2639
rect 3174 2634 3175 2638
rect 3179 2634 3180 2638
rect 3174 2633 3180 2634
rect 3310 2638 3316 2639
rect 3310 2634 3311 2638
rect 3315 2634 3316 2638
rect 3310 2633 3316 2634
rect 3454 2638 3460 2639
rect 3454 2634 3455 2638
rect 3459 2634 3460 2638
rect 3454 2633 3460 2634
rect 3990 2633 3996 2634
rect 1926 2629 1932 2630
rect 2030 2629 2036 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 110 2624 116 2625
rect 2030 2625 2031 2629
rect 2035 2625 2036 2629
rect 2070 2629 2071 2633
rect 2075 2629 2076 2633
rect 2070 2628 2076 2629
rect 3990 2629 3991 2633
rect 3995 2629 3996 2633
rect 3990 2628 3996 2629
rect 2030 2624 2036 2625
rect 1222 2623 1228 2624
rect 1222 2619 1223 2623
rect 1227 2622 1228 2623
rect 1646 2623 1652 2624
rect 1646 2622 1647 2623
rect 1227 2620 1647 2622
rect 1227 2619 1228 2620
rect 1222 2618 1228 2619
rect 1646 2619 1647 2620
rect 1651 2619 1652 2623
rect 1646 2618 1652 2619
rect 2070 2616 2076 2617
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 110 2607 116 2608
rect 2030 2612 2036 2613
rect 2030 2608 2031 2612
rect 2035 2608 2036 2612
rect 2070 2612 2071 2616
rect 2075 2612 2076 2616
rect 2070 2611 2076 2612
rect 3990 2616 3996 2617
rect 3990 2612 3991 2616
rect 3995 2612 3996 2616
rect 3990 2611 3996 2612
rect 2030 2607 2036 2608
rect 2182 2607 2188 2608
rect 2182 2606 2183 2607
rect 2161 2604 2183 2606
rect 246 2603 252 2604
rect 246 2599 247 2603
rect 251 2599 252 2603
rect 798 2603 804 2604
rect 649 2600 766 2602
rect 246 2598 252 2599
rect 254 2593 260 2594
rect 254 2589 255 2593
rect 259 2589 260 2593
rect 254 2588 260 2589
rect 422 2593 428 2594
rect 422 2589 423 2593
rect 427 2589 428 2593
rect 422 2588 428 2589
rect 598 2593 604 2594
rect 598 2589 599 2593
rect 603 2589 604 2593
rect 598 2588 604 2589
rect 764 2586 766 2600
rect 798 2599 799 2603
rect 803 2599 804 2603
rect 1222 2603 1228 2604
rect 1222 2602 1223 2603
rect 1201 2600 1223 2602
rect 798 2598 804 2599
rect 1222 2599 1223 2600
rect 1227 2599 1228 2603
rect 1798 2603 1804 2604
rect 1798 2602 1799 2603
rect 1777 2600 1799 2602
rect 1222 2598 1228 2599
rect 1798 2599 1799 2600
rect 1803 2599 1804 2603
rect 2182 2603 2183 2604
rect 2187 2603 2188 2607
rect 2582 2607 2588 2608
rect 2582 2606 2583 2607
rect 2481 2604 2583 2606
rect 2182 2602 2188 2603
rect 2582 2603 2583 2604
rect 2587 2603 2588 2607
rect 2862 2607 2868 2608
rect 2862 2606 2863 2607
rect 2801 2604 2863 2606
rect 2582 2602 2588 2603
rect 2862 2603 2863 2604
rect 2867 2603 2868 2607
rect 3022 2607 3028 2608
rect 3022 2606 3023 2607
rect 2945 2604 3023 2606
rect 2862 2602 2868 2603
rect 3022 2603 3023 2604
rect 3027 2603 3028 2607
rect 3022 2602 3028 2603
rect 1798 2598 1804 2599
rect 2110 2597 2116 2598
rect 774 2593 780 2594
rect 774 2589 775 2593
rect 779 2589 780 2593
rect 958 2593 964 2594
rect 774 2588 780 2589
rect 840 2588 954 2590
rect 958 2589 959 2593
rect 963 2589 964 2593
rect 958 2588 964 2589
rect 1150 2593 1156 2594
rect 1150 2589 1151 2593
rect 1155 2589 1156 2593
rect 1150 2588 1156 2589
rect 1342 2593 1348 2594
rect 1342 2589 1343 2593
rect 1347 2589 1348 2593
rect 1342 2588 1348 2589
rect 1534 2593 1540 2594
rect 1534 2589 1535 2593
rect 1539 2589 1540 2593
rect 1534 2588 1540 2589
rect 1726 2593 1732 2594
rect 1726 2589 1727 2593
rect 1731 2589 1732 2593
rect 1726 2588 1732 2589
rect 1926 2593 1932 2594
rect 1926 2589 1927 2593
rect 1931 2589 1932 2593
rect 2110 2593 2111 2597
rect 2115 2593 2116 2597
rect 2110 2592 2116 2593
rect 2262 2597 2268 2598
rect 2262 2593 2263 2597
rect 2267 2593 2268 2597
rect 2262 2592 2268 2593
rect 2430 2597 2436 2598
rect 2430 2593 2431 2597
rect 2435 2593 2436 2597
rect 2430 2592 2436 2593
rect 2598 2597 2604 2598
rect 2598 2593 2599 2597
rect 2603 2593 2604 2597
rect 2598 2592 2604 2593
rect 2750 2597 2756 2598
rect 2750 2593 2751 2597
rect 2755 2593 2756 2597
rect 2750 2592 2756 2593
rect 2894 2597 2900 2598
rect 2894 2593 2895 2597
rect 2899 2593 2900 2597
rect 2894 2592 2900 2593
rect 3038 2597 3044 2598
rect 3038 2593 3039 2597
rect 3043 2593 3044 2597
rect 3038 2592 3044 2593
rect 3174 2597 3180 2598
rect 3174 2593 3175 2597
rect 3179 2593 3180 2597
rect 3174 2592 3180 2593
rect 3310 2597 3316 2598
rect 3310 2593 3311 2597
rect 3315 2593 3316 2597
rect 3310 2592 3316 2593
rect 3454 2597 3460 2598
rect 3454 2593 3455 2597
rect 3459 2593 3460 2597
rect 3454 2592 3460 2593
rect 1926 2588 1932 2589
rect 840 2586 842 2588
rect 764 2584 842 2586
rect 327 2583 333 2584
rect 327 2579 328 2583
rect 332 2582 333 2583
rect 407 2583 413 2584
rect 407 2582 408 2583
rect 332 2580 408 2582
rect 332 2579 333 2580
rect 327 2578 333 2579
rect 407 2579 408 2580
rect 412 2579 413 2583
rect 407 2578 413 2579
rect 495 2583 501 2584
rect 495 2579 496 2583
rect 500 2582 501 2583
rect 670 2583 677 2584
rect 500 2580 514 2582
rect 500 2579 501 2580
rect 495 2578 501 2579
rect 391 2567 397 2568
rect 391 2563 392 2567
rect 396 2566 397 2567
rect 430 2567 436 2568
rect 430 2566 431 2567
rect 396 2564 431 2566
rect 396 2563 397 2564
rect 391 2562 397 2563
rect 430 2563 431 2564
rect 435 2563 436 2567
rect 512 2566 514 2580
rect 670 2579 671 2583
rect 676 2579 677 2583
rect 670 2578 677 2579
rect 847 2583 853 2584
rect 847 2579 848 2583
rect 852 2582 853 2583
rect 943 2583 949 2584
rect 943 2582 944 2583
rect 852 2580 944 2582
rect 852 2579 853 2580
rect 847 2578 853 2579
rect 943 2579 944 2580
rect 948 2579 949 2583
rect 952 2582 954 2588
rect 2183 2587 2189 2588
rect 1031 2583 1037 2584
rect 1031 2582 1032 2583
rect 952 2580 1032 2582
rect 943 2578 949 2579
rect 1031 2579 1032 2580
rect 1036 2579 1037 2583
rect 1031 2578 1037 2579
rect 1223 2583 1229 2584
rect 1223 2579 1224 2583
rect 1228 2582 1229 2583
rect 1327 2583 1333 2584
rect 1327 2582 1328 2583
rect 1228 2580 1328 2582
rect 1228 2579 1229 2580
rect 1223 2578 1229 2579
rect 1327 2579 1328 2580
rect 1332 2579 1333 2583
rect 1327 2578 1333 2579
rect 1415 2583 1421 2584
rect 1415 2579 1416 2583
rect 1420 2582 1421 2583
rect 1519 2583 1525 2584
rect 1519 2582 1520 2583
rect 1420 2580 1520 2582
rect 1420 2579 1421 2580
rect 1415 2578 1421 2579
rect 1519 2579 1520 2580
rect 1524 2579 1525 2583
rect 1519 2578 1525 2579
rect 1582 2583 1588 2584
rect 1582 2579 1583 2583
rect 1587 2582 1588 2583
rect 1607 2583 1613 2584
rect 1607 2582 1608 2583
rect 1587 2580 1608 2582
rect 1587 2579 1588 2580
rect 1582 2578 1588 2579
rect 1607 2579 1608 2580
rect 1612 2579 1613 2583
rect 1607 2578 1613 2579
rect 1799 2583 1805 2584
rect 1799 2579 1800 2583
rect 1804 2582 1805 2583
rect 1911 2583 1917 2584
rect 1911 2582 1912 2583
rect 1804 2580 1912 2582
rect 1804 2579 1805 2580
rect 1799 2578 1805 2579
rect 1911 2579 1912 2580
rect 1916 2579 1917 2583
rect 1911 2578 1917 2579
rect 1998 2583 2005 2584
rect 1998 2579 1999 2583
rect 2004 2579 2005 2583
rect 2183 2583 2184 2587
rect 2188 2586 2189 2587
rect 2247 2587 2253 2588
rect 2247 2586 2248 2587
rect 2188 2584 2248 2586
rect 2188 2583 2189 2584
rect 2183 2582 2189 2583
rect 2247 2583 2248 2584
rect 2252 2583 2253 2587
rect 2247 2582 2253 2583
rect 2335 2587 2341 2588
rect 2335 2583 2336 2587
rect 2340 2583 2341 2587
rect 2335 2582 2341 2583
rect 2503 2587 2509 2588
rect 2503 2583 2504 2587
rect 2508 2586 2509 2587
rect 2583 2587 2589 2588
rect 2583 2586 2584 2587
rect 2508 2584 2584 2586
rect 2508 2583 2509 2584
rect 2503 2582 2509 2583
rect 2583 2583 2584 2584
rect 2588 2583 2589 2587
rect 2583 2582 2589 2583
rect 2671 2587 2677 2588
rect 2671 2583 2672 2587
rect 2676 2586 2677 2587
rect 2682 2587 2688 2588
rect 2682 2586 2683 2587
rect 2676 2584 2683 2586
rect 2676 2583 2677 2584
rect 2671 2582 2677 2583
rect 2682 2583 2683 2584
rect 2687 2583 2688 2587
rect 2823 2587 2829 2588
rect 2823 2586 2824 2587
rect 2682 2582 2688 2583
rect 2692 2584 2824 2586
rect 1998 2578 2005 2579
rect 2582 2579 2588 2580
rect 1335 2575 1341 2576
rect 1335 2571 1336 2575
rect 1340 2574 1341 2575
rect 2423 2575 2429 2576
rect 1340 2572 1466 2574
rect 1340 2571 1341 2572
rect 1335 2570 1341 2571
rect 519 2567 525 2568
rect 519 2566 520 2567
rect 512 2564 520 2566
rect 430 2562 436 2563
rect 519 2563 520 2564
rect 524 2563 525 2567
rect 607 2567 613 2568
rect 607 2566 608 2567
rect 519 2562 525 2563
rect 528 2564 608 2566
rect 318 2559 324 2560
rect 318 2555 319 2559
rect 323 2555 324 2559
rect 318 2554 324 2555
rect 528 2554 530 2564
rect 607 2563 608 2564
rect 612 2563 613 2567
rect 607 2562 613 2563
rect 798 2567 804 2568
rect 798 2563 799 2567
rect 803 2566 804 2567
rect 815 2567 821 2568
rect 815 2566 816 2567
rect 803 2564 816 2566
rect 803 2563 804 2564
rect 798 2562 804 2563
rect 815 2563 816 2564
rect 820 2563 821 2567
rect 1023 2567 1029 2568
rect 1023 2566 1024 2567
rect 815 2562 821 2563
rect 876 2564 1024 2566
rect 534 2559 540 2560
rect 534 2555 535 2559
rect 539 2555 540 2559
rect 534 2554 540 2555
rect 742 2559 748 2560
rect 742 2555 743 2559
rect 747 2555 748 2559
rect 742 2554 748 2555
rect 464 2552 530 2554
rect 464 2550 466 2552
rect 876 2550 878 2564
rect 1023 2563 1024 2564
rect 1028 2563 1029 2567
rect 1023 2562 1029 2563
rect 1231 2567 1237 2568
rect 1231 2563 1232 2567
rect 1236 2566 1237 2567
rect 1343 2567 1349 2568
rect 1343 2566 1344 2567
rect 1236 2564 1344 2566
rect 1236 2563 1237 2564
rect 1231 2562 1237 2563
rect 1343 2563 1344 2564
rect 1348 2563 1349 2567
rect 1343 2562 1349 2563
rect 1431 2567 1437 2568
rect 1431 2563 1432 2567
rect 1436 2566 1437 2567
rect 1454 2567 1460 2568
rect 1454 2566 1455 2567
rect 1436 2564 1455 2566
rect 1436 2563 1437 2564
rect 1431 2562 1437 2563
rect 1454 2563 1455 2564
rect 1459 2563 1460 2567
rect 1464 2566 1466 2572
rect 2423 2571 2424 2575
rect 2428 2574 2429 2575
rect 2582 2575 2583 2579
rect 2587 2578 2588 2579
rect 2692 2578 2694 2584
rect 2823 2583 2824 2584
rect 2828 2583 2829 2587
rect 2823 2582 2829 2583
rect 2967 2587 2973 2588
rect 2967 2583 2968 2587
rect 2972 2586 2973 2587
rect 3023 2587 3029 2588
rect 3023 2586 3024 2587
rect 2972 2584 3024 2586
rect 2972 2583 2973 2584
rect 2967 2582 2973 2583
rect 3023 2583 3024 2584
rect 3028 2583 3029 2587
rect 3023 2582 3029 2583
rect 3111 2587 3117 2588
rect 3111 2583 3112 2587
rect 3116 2586 3117 2587
rect 3159 2587 3165 2588
rect 3159 2586 3160 2587
rect 3116 2584 3160 2586
rect 3116 2583 3117 2584
rect 3111 2582 3117 2583
rect 3159 2583 3160 2584
rect 3164 2583 3165 2587
rect 3159 2582 3165 2583
rect 3247 2587 3253 2588
rect 3247 2583 3248 2587
rect 3252 2586 3253 2587
rect 3295 2587 3301 2588
rect 3295 2586 3296 2587
rect 3252 2584 3296 2586
rect 3252 2583 3253 2584
rect 3247 2582 3253 2583
rect 3295 2583 3296 2584
rect 3300 2583 3301 2587
rect 3295 2582 3301 2583
rect 3383 2587 3389 2588
rect 3383 2583 3384 2587
rect 3388 2586 3389 2587
rect 3439 2587 3445 2588
rect 3439 2586 3440 2587
rect 3388 2584 3440 2586
rect 3388 2583 3389 2584
rect 3383 2582 3389 2583
rect 3439 2583 3440 2584
rect 3444 2583 3445 2587
rect 3439 2582 3445 2583
rect 3526 2587 3533 2588
rect 3526 2583 3527 2587
rect 3532 2583 3533 2587
rect 3526 2582 3533 2583
rect 2587 2576 2694 2578
rect 2587 2575 2588 2576
rect 2582 2574 2588 2575
rect 3022 2575 3028 2576
rect 2428 2572 2550 2574
rect 2428 2571 2429 2572
rect 2423 2570 2429 2571
rect 1631 2567 1637 2568
rect 1631 2566 1632 2567
rect 1464 2564 1632 2566
rect 1454 2562 1460 2563
rect 1631 2563 1632 2564
rect 1636 2563 1637 2567
rect 1631 2562 1637 2563
rect 1798 2567 1804 2568
rect 1798 2563 1799 2567
rect 1803 2566 1804 2567
rect 1831 2567 1837 2568
rect 1831 2566 1832 2567
rect 1803 2564 1832 2566
rect 1803 2563 1804 2564
rect 1798 2562 1804 2563
rect 1831 2563 1832 2564
rect 1836 2563 1837 2567
rect 1831 2562 1837 2563
rect 2007 2567 2013 2568
rect 2007 2563 2008 2567
rect 2012 2566 2013 2567
rect 2095 2567 2101 2568
rect 2095 2566 2096 2567
rect 2012 2564 2096 2566
rect 2012 2563 2013 2564
rect 2007 2562 2013 2563
rect 2095 2563 2096 2564
rect 2100 2563 2101 2567
rect 2095 2562 2101 2563
rect 2182 2567 2189 2568
rect 2182 2563 2183 2567
rect 2188 2563 2189 2567
rect 2182 2562 2189 2563
rect 2343 2567 2349 2568
rect 2343 2563 2344 2567
rect 2348 2566 2349 2567
rect 2431 2567 2437 2568
rect 2431 2566 2432 2567
rect 2348 2564 2432 2566
rect 2348 2563 2349 2564
rect 2343 2562 2349 2563
rect 2431 2563 2432 2564
rect 2436 2563 2437 2567
rect 2431 2562 2437 2563
rect 2519 2567 2525 2568
rect 2519 2563 2520 2567
rect 2524 2566 2525 2567
rect 2538 2567 2544 2568
rect 2538 2566 2539 2567
rect 2524 2564 2539 2566
rect 2524 2563 2525 2564
rect 2519 2562 2525 2563
rect 2538 2563 2539 2564
rect 2543 2563 2544 2567
rect 2548 2566 2550 2572
rect 3022 2571 3023 2575
rect 3027 2574 3028 2575
rect 3027 2572 3314 2574
rect 3027 2571 3028 2572
rect 3022 2570 3028 2571
rect 2687 2567 2693 2568
rect 2687 2566 2688 2567
rect 2548 2564 2688 2566
rect 2538 2562 2544 2563
rect 2687 2563 2688 2564
rect 2692 2563 2693 2567
rect 2687 2562 2693 2563
rect 2839 2567 2845 2568
rect 2839 2563 2840 2567
rect 2844 2566 2845 2567
rect 2895 2567 2901 2568
rect 2895 2566 2896 2567
rect 2844 2564 2896 2566
rect 2844 2563 2845 2564
rect 2839 2562 2845 2563
rect 2895 2563 2896 2564
rect 2900 2563 2901 2567
rect 2895 2562 2901 2563
rect 2983 2567 2989 2568
rect 2983 2563 2984 2567
rect 2988 2566 2989 2567
rect 3031 2567 3037 2568
rect 3031 2566 3032 2567
rect 2988 2564 3032 2566
rect 2988 2563 2989 2564
rect 2983 2562 2989 2563
rect 3031 2563 3032 2564
rect 3036 2563 3037 2567
rect 3031 2562 3037 2563
rect 3119 2567 3125 2568
rect 3119 2563 3120 2567
rect 3124 2566 3125 2567
rect 3167 2567 3173 2568
rect 3167 2566 3168 2567
rect 3124 2564 3168 2566
rect 3124 2563 3125 2564
rect 3119 2562 3125 2563
rect 3167 2563 3168 2564
rect 3172 2563 3173 2567
rect 3167 2562 3173 2563
rect 3255 2567 3261 2568
rect 3255 2563 3256 2567
rect 3260 2566 3261 2567
rect 3303 2567 3309 2568
rect 3303 2566 3304 2567
rect 3260 2564 3304 2566
rect 3260 2563 3261 2564
rect 3255 2562 3261 2563
rect 3303 2563 3304 2564
rect 3308 2563 3309 2567
rect 3312 2566 3314 2572
rect 3391 2567 3397 2568
rect 3391 2566 3392 2567
rect 3312 2564 3392 2566
rect 3303 2562 3309 2563
rect 3391 2563 3392 2564
rect 3396 2563 3397 2567
rect 3391 2562 3397 2563
rect 950 2559 956 2560
rect 950 2555 951 2559
rect 955 2555 956 2559
rect 950 2554 956 2555
rect 1158 2559 1164 2560
rect 1158 2555 1159 2559
rect 1163 2555 1164 2559
rect 1158 2554 1164 2555
rect 1358 2559 1364 2560
rect 1358 2555 1359 2559
rect 1363 2555 1364 2559
rect 1358 2554 1364 2555
rect 1558 2559 1564 2560
rect 1558 2555 1559 2559
rect 1563 2555 1564 2559
rect 1558 2554 1564 2555
rect 1758 2559 1764 2560
rect 1758 2555 1759 2559
rect 1763 2555 1764 2559
rect 1758 2554 1764 2555
rect 1934 2559 1940 2560
rect 1934 2555 1935 2559
rect 1939 2555 1940 2559
rect 1934 2554 1940 2555
rect 2110 2559 2116 2560
rect 2110 2555 2111 2559
rect 2115 2555 2116 2559
rect 2110 2554 2116 2555
rect 2270 2559 2276 2560
rect 2270 2555 2271 2559
rect 2275 2555 2276 2559
rect 2270 2554 2276 2555
rect 2446 2559 2452 2560
rect 2446 2555 2447 2559
rect 2451 2555 2452 2559
rect 2446 2554 2452 2555
rect 2614 2559 2620 2560
rect 2614 2555 2615 2559
rect 2619 2555 2620 2559
rect 2614 2554 2620 2555
rect 2766 2559 2772 2560
rect 2766 2555 2767 2559
rect 2771 2555 2772 2559
rect 2766 2554 2772 2555
rect 2910 2559 2916 2560
rect 2910 2555 2911 2559
rect 2915 2555 2916 2559
rect 2910 2554 2916 2555
rect 3046 2559 3052 2560
rect 3046 2555 3047 2559
rect 3051 2555 3052 2559
rect 3046 2554 3052 2555
rect 3182 2559 3188 2560
rect 3182 2555 3183 2559
rect 3187 2555 3188 2559
rect 3182 2554 3188 2555
rect 3318 2559 3324 2560
rect 3318 2555 3319 2559
rect 3323 2555 3324 2559
rect 3318 2554 3324 2555
rect 1030 2551 1036 2552
rect 1030 2550 1031 2551
rect 369 2548 466 2550
rect 793 2548 878 2550
rect 1001 2548 1031 2550
rect 1030 2547 1031 2548
rect 1035 2547 1036 2551
rect 1335 2551 1341 2552
rect 1335 2550 1336 2551
rect 1209 2548 1336 2550
rect 1030 2546 1036 2547
rect 1335 2547 1336 2548
rect 1340 2547 1341 2551
rect 1858 2551 1864 2552
rect 1858 2550 1859 2551
rect 1809 2548 1859 2550
rect 1335 2546 1341 2547
rect 1582 2547 1588 2548
rect 1582 2543 1583 2547
rect 1587 2543 1588 2547
rect 1858 2547 1859 2548
rect 1863 2547 1864 2551
rect 2006 2551 2012 2552
rect 2006 2550 2007 2551
rect 1985 2548 2007 2550
rect 1858 2546 1864 2547
rect 2006 2547 2007 2548
rect 2011 2547 2012 2551
rect 2423 2551 2429 2552
rect 2423 2550 2424 2551
rect 2321 2548 2424 2550
rect 2006 2546 2012 2547
rect 2423 2547 2424 2548
rect 2428 2547 2429 2551
rect 2682 2551 2688 2552
rect 2682 2550 2683 2551
rect 2665 2548 2683 2550
rect 2423 2546 2429 2547
rect 2682 2547 2683 2548
rect 2687 2547 2688 2551
rect 2894 2551 2900 2552
rect 2894 2550 2895 2551
rect 2817 2548 2895 2550
rect 2682 2546 2688 2547
rect 2894 2547 2895 2548
rect 2899 2547 2900 2551
rect 2894 2546 2900 2547
rect 1582 2542 1588 2543
rect 110 2540 116 2541
rect 110 2536 111 2540
rect 115 2536 116 2540
rect 110 2535 116 2536
rect 2030 2540 2036 2541
rect 2030 2536 2031 2540
rect 2035 2536 2036 2540
rect 2030 2535 2036 2536
rect 2070 2540 2076 2541
rect 2070 2536 2071 2540
rect 2075 2536 2076 2540
rect 2070 2535 2076 2536
rect 3990 2540 3996 2541
rect 3990 2536 3991 2540
rect 3995 2536 3996 2540
rect 3990 2535 3996 2536
rect 110 2523 116 2524
rect 110 2519 111 2523
rect 115 2519 116 2523
rect 2030 2523 2036 2524
rect 2030 2519 2031 2523
rect 2035 2519 2036 2523
rect 110 2518 116 2519
rect 318 2518 324 2519
rect 318 2514 319 2518
rect 323 2514 324 2518
rect 318 2513 324 2514
rect 534 2518 540 2519
rect 534 2514 535 2518
rect 539 2514 540 2518
rect 534 2513 540 2514
rect 742 2518 748 2519
rect 742 2514 743 2518
rect 747 2514 748 2518
rect 742 2513 748 2514
rect 950 2518 956 2519
rect 950 2514 951 2518
rect 955 2514 956 2518
rect 950 2513 956 2514
rect 1158 2518 1164 2519
rect 1158 2514 1159 2518
rect 1163 2514 1164 2518
rect 1158 2513 1164 2514
rect 1358 2518 1364 2519
rect 1358 2514 1359 2518
rect 1363 2514 1364 2518
rect 1358 2513 1364 2514
rect 1558 2518 1564 2519
rect 1558 2514 1559 2518
rect 1563 2514 1564 2518
rect 1558 2513 1564 2514
rect 1758 2518 1764 2519
rect 1758 2514 1759 2518
rect 1763 2514 1764 2518
rect 1758 2513 1764 2514
rect 1934 2518 1940 2519
rect 2030 2518 2036 2519
rect 2070 2523 2076 2524
rect 2070 2519 2071 2523
rect 2075 2519 2076 2523
rect 3990 2523 3996 2524
rect 3990 2519 3991 2523
rect 3995 2519 3996 2523
rect 2070 2518 2076 2519
rect 2110 2518 2116 2519
rect 1934 2514 1935 2518
rect 1939 2514 1940 2518
rect 1934 2513 1940 2514
rect 2110 2514 2111 2518
rect 2115 2514 2116 2518
rect 2110 2513 2116 2514
rect 2270 2518 2276 2519
rect 2270 2514 2271 2518
rect 2275 2514 2276 2518
rect 2270 2513 2276 2514
rect 2446 2518 2452 2519
rect 2446 2514 2447 2518
rect 2451 2514 2452 2518
rect 2446 2513 2452 2514
rect 2614 2518 2620 2519
rect 2614 2514 2615 2518
rect 2619 2514 2620 2518
rect 2614 2513 2620 2514
rect 2766 2518 2772 2519
rect 2766 2514 2767 2518
rect 2771 2514 2772 2518
rect 2766 2513 2772 2514
rect 2910 2518 2916 2519
rect 2910 2514 2911 2518
rect 2915 2514 2916 2518
rect 2910 2513 2916 2514
rect 3046 2518 3052 2519
rect 3046 2514 3047 2518
rect 3051 2514 3052 2518
rect 3046 2513 3052 2514
rect 3182 2518 3188 2519
rect 3182 2514 3183 2518
rect 3187 2514 3188 2518
rect 3182 2513 3188 2514
rect 3318 2518 3324 2519
rect 3990 2518 3996 2519
rect 3318 2514 3319 2518
rect 3323 2514 3324 2518
rect 3318 2513 3324 2514
rect 278 2486 284 2487
rect 278 2482 279 2486
rect 283 2482 284 2486
rect 110 2481 116 2482
rect 278 2481 284 2482
rect 438 2486 444 2487
rect 438 2482 439 2486
rect 443 2482 444 2486
rect 438 2481 444 2482
rect 606 2486 612 2487
rect 606 2482 607 2486
rect 611 2482 612 2486
rect 606 2481 612 2482
rect 782 2486 788 2487
rect 782 2482 783 2486
rect 787 2482 788 2486
rect 782 2481 788 2482
rect 958 2486 964 2487
rect 958 2482 959 2486
rect 963 2482 964 2486
rect 958 2481 964 2482
rect 1126 2486 1132 2487
rect 1126 2482 1127 2486
rect 1131 2482 1132 2486
rect 1126 2481 1132 2482
rect 1294 2486 1300 2487
rect 1294 2482 1295 2486
rect 1299 2482 1300 2486
rect 1294 2481 1300 2482
rect 1462 2486 1468 2487
rect 1462 2482 1463 2486
rect 1467 2482 1468 2486
rect 1462 2481 1468 2482
rect 1622 2486 1628 2487
rect 1622 2482 1623 2486
rect 1627 2482 1628 2486
rect 1622 2481 1628 2482
rect 1790 2486 1796 2487
rect 1790 2482 1791 2486
rect 1795 2482 1796 2486
rect 1790 2481 1796 2482
rect 1934 2486 1940 2487
rect 1934 2482 1935 2486
rect 1939 2482 1940 2486
rect 1934 2481 1940 2482
rect 2030 2481 2036 2482
rect 110 2477 111 2481
rect 115 2477 116 2481
rect 110 2476 116 2477
rect 2030 2477 2031 2481
rect 2035 2477 2036 2481
rect 2030 2476 2036 2477
rect 2622 2474 2628 2475
rect 2622 2470 2623 2474
rect 2627 2470 2628 2474
rect 2070 2469 2076 2470
rect 2622 2469 2628 2470
rect 2742 2474 2748 2475
rect 2742 2470 2743 2474
rect 2747 2470 2748 2474
rect 2742 2469 2748 2470
rect 2870 2474 2876 2475
rect 2870 2470 2871 2474
rect 2875 2470 2876 2474
rect 2870 2469 2876 2470
rect 3014 2474 3020 2475
rect 3014 2470 3015 2474
rect 3019 2470 3020 2474
rect 3014 2469 3020 2470
rect 3158 2474 3164 2475
rect 3158 2470 3159 2474
rect 3163 2470 3164 2474
rect 3158 2469 3164 2470
rect 3310 2474 3316 2475
rect 3310 2470 3311 2474
rect 3315 2470 3316 2474
rect 3310 2469 3316 2470
rect 3462 2474 3468 2475
rect 3462 2470 3463 2474
rect 3467 2470 3468 2474
rect 3462 2469 3468 2470
rect 3614 2474 3620 2475
rect 3614 2470 3615 2474
rect 3619 2470 3620 2474
rect 3614 2469 3620 2470
rect 3766 2474 3772 2475
rect 3766 2470 3767 2474
rect 3771 2470 3772 2474
rect 3766 2469 3772 2470
rect 3894 2474 3900 2475
rect 3894 2470 3895 2474
rect 3899 2470 3900 2474
rect 3894 2469 3900 2470
rect 3990 2469 3996 2470
rect 2070 2465 2071 2469
rect 2075 2465 2076 2469
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 110 2459 116 2460
rect 2030 2464 2036 2465
rect 2070 2464 2076 2465
rect 3990 2465 3991 2469
rect 3995 2465 3996 2469
rect 3990 2464 3996 2465
rect 2030 2460 2031 2464
rect 2035 2460 2036 2464
rect 2030 2459 2036 2460
rect 418 2455 424 2456
rect 418 2454 419 2455
rect 329 2452 419 2454
rect 418 2451 419 2452
rect 423 2451 424 2455
rect 418 2450 424 2451
rect 430 2455 436 2456
rect 430 2451 431 2455
rect 435 2451 436 2455
rect 678 2455 684 2456
rect 678 2454 679 2455
rect 657 2452 679 2454
rect 430 2450 436 2451
rect 678 2451 679 2452
rect 683 2451 684 2455
rect 1278 2455 1284 2456
rect 1278 2454 1279 2455
rect 1177 2452 1279 2454
rect 678 2450 684 2451
rect 1278 2451 1279 2452
rect 1283 2451 1284 2455
rect 1278 2450 1284 2451
rect 1454 2455 1460 2456
rect 1454 2451 1455 2455
rect 1459 2451 1460 2455
rect 1694 2455 1700 2456
rect 1694 2454 1695 2455
rect 1673 2452 1695 2454
rect 1454 2450 1460 2451
rect 1694 2451 1695 2452
rect 1699 2451 1700 2455
rect 1694 2450 1700 2451
rect 2070 2452 2076 2453
rect 2070 2448 2071 2452
rect 2075 2448 2076 2452
rect 2070 2447 2076 2448
rect 3990 2452 3996 2453
rect 3990 2448 3991 2452
rect 3995 2448 3996 2452
rect 3990 2447 3996 2448
rect 278 2445 284 2446
rect 278 2441 279 2445
rect 283 2441 284 2445
rect 278 2440 284 2441
rect 438 2445 444 2446
rect 438 2441 439 2445
rect 443 2441 444 2445
rect 438 2440 444 2441
rect 606 2445 612 2446
rect 606 2441 607 2445
rect 611 2441 612 2445
rect 606 2440 612 2441
rect 782 2445 788 2446
rect 782 2441 783 2445
rect 787 2441 788 2445
rect 782 2440 788 2441
rect 958 2445 964 2446
rect 958 2441 959 2445
rect 963 2441 964 2445
rect 958 2440 964 2441
rect 1126 2445 1132 2446
rect 1126 2441 1127 2445
rect 1131 2441 1132 2445
rect 1126 2440 1132 2441
rect 1294 2445 1300 2446
rect 1294 2441 1295 2445
rect 1299 2441 1300 2445
rect 1294 2440 1300 2441
rect 1462 2445 1468 2446
rect 1462 2441 1463 2445
rect 1467 2441 1468 2445
rect 1462 2440 1468 2441
rect 1622 2445 1628 2446
rect 1622 2441 1623 2445
rect 1627 2441 1628 2445
rect 1622 2440 1628 2441
rect 1790 2445 1796 2446
rect 1790 2441 1791 2445
rect 1795 2441 1796 2445
rect 1790 2440 1796 2441
rect 1934 2445 1940 2446
rect 1934 2441 1935 2445
rect 1939 2441 1940 2445
rect 1934 2440 1940 2441
rect 2538 2443 2544 2444
rect 2538 2439 2539 2443
rect 2543 2442 2544 2443
rect 2942 2443 2948 2444
rect 2942 2442 2943 2443
rect 2543 2440 2617 2442
rect 2921 2440 2943 2442
rect 2543 2439 2544 2440
rect 2538 2438 2544 2439
rect 2942 2439 2943 2440
rect 2947 2439 2948 2443
rect 3566 2443 3572 2444
rect 3566 2442 3567 2443
rect 3513 2440 3567 2442
rect 2942 2438 2948 2439
rect 3566 2439 3567 2440
rect 3571 2439 3572 2443
rect 3878 2443 3884 2444
rect 3878 2442 3879 2443
rect 3817 2440 3879 2442
rect 3566 2438 3572 2439
rect 3878 2439 3879 2440
rect 3883 2439 3884 2443
rect 3966 2443 3972 2444
rect 3966 2442 3967 2443
rect 3945 2440 3967 2442
rect 3878 2438 3884 2439
rect 3966 2439 3967 2440
rect 3971 2439 3972 2443
rect 3966 2438 3972 2439
rect 350 2435 357 2436
rect 350 2431 351 2435
rect 356 2431 357 2435
rect 350 2430 357 2431
rect 418 2435 424 2436
rect 418 2431 419 2435
rect 423 2434 424 2435
rect 511 2435 517 2436
rect 511 2434 512 2435
rect 423 2432 512 2434
rect 423 2431 424 2432
rect 418 2430 424 2431
rect 511 2431 512 2432
rect 516 2431 517 2435
rect 511 2430 517 2431
rect 679 2435 685 2436
rect 679 2431 680 2435
rect 684 2434 685 2435
rect 767 2435 773 2436
rect 767 2434 768 2435
rect 684 2432 768 2434
rect 684 2431 685 2432
rect 679 2430 685 2431
rect 767 2431 768 2432
rect 772 2431 773 2435
rect 767 2430 773 2431
rect 855 2435 861 2436
rect 855 2431 856 2435
rect 860 2434 861 2435
rect 943 2435 949 2436
rect 943 2434 944 2435
rect 860 2432 944 2434
rect 860 2431 861 2432
rect 855 2430 861 2431
rect 943 2431 944 2432
rect 948 2431 949 2435
rect 943 2430 949 2431
rect 1030 2435 1037 2436
rect 1030 2431 1031 2435
rect 1036 2431 1037 2435
rect 1030 2430 1037 2431
rect 1199 2435 1205 2436
rect 1199 2431 1200 2435
rect 1204 2434 1205 2435
rect 1279 2435 1285 2436
rect 1279 2434 1280 2435
rect 1204 2432 1280 2434
rect 1204 2431 1205 2432
rect 1199 2430 1205 2431
rect 1279 2431 1280 2432
rect 1284 2431 1285 2435
rect 1279 2430 1285 2431
rect 1367 2435 1376 2436
rect 1367 2431 1368 2435
rect 1375 2431 1376 2435
rect 1535 2435 1541 2436
rect 1535 2434 1536 2435
rect 1367 2430 1376 2431
rect 1380 2432 1536 2434
rect 1278 2427 1284 2428
rect 1278 2423 1279 2427
rect 1283 2426 1284 2427
rect 1380 2426 1382 2432
rect 1535 2431 1536 2432
rect 1540 2431 1541 2435
rect 1535 2430 1541 2431
rect 1695 2435 1701 2436
rect 1695 2431 1696 2435
rect 1700 2434 1701 2435
rect 1775 2435 1781 2436
rect 1775 2434 1776 2435
rect 1700 2432 1776 2434
rect 1700 2431 1701 2432
rect 1695 2430 1701 2431
rect 1775 2431 1776 2432
rect 1780 2431 1781 2435
rect 1775 2430 1781 2431
rect 1858 2435 1869 2436
rect 1858 2431 1859 2435
rect 1863 2431 1864 2435
rect 1868 2431 1869 2435
rect 1858 2430 1869 2431
rect 1890 2435 1896 2436
rect 1890 2431 1891 2435
rect 1895 2434 1896 2435
rect 1919 2435 1925 2436
rect 1919 2434 1920 2435
rect 1895 2432 1920 2434
rect 1895 2431 1896 2432
rect 1890 2430 1896 2431
rect 1919 2431 1920 2432
rect 1924 2431 1925 2435
rect 1919 2430 1925 2431
rect 2006 2435 2013 2436
rect 2006 2431 2007 2435
rect 2012 2431 2013 2435
rect 2006 2430 2013 2431
rect 2622 2433 2628 2434
rect 2622 2429 2623 2433
rect 2627 2429 2628 2433
rect 2622 2428 2628 2429
rect 2742 2433 2748 2434
rect 2742 2429 2743 2433
rect 2747 2429 2748 2433
rect 2742 2428 2748 2429
rect 2870 2433 2876 2434
rect 2870 2429 2871 2433
rect 2875 2429 2876 2433
rect 2870 2428 2876 2429
rect 3014 2433 3020 2434
rect 3014 2429 3015 2433
rect 3019 2429 3020 2433
rect 3014 2428 3020 2429
rect 3158 2433 3164 2434
rect 3158 2429 3159 2433
rect 3163 2429 3164 2433
rect 3158 2428 3164 2429
rect 3310 2433 3316 2434
rect 3310 2429 3311 2433
rect 3315 2429 3316 2433
rect 3310 2428 3316 2429
rect 3462 2433 3468 2434
rect 3462 2429 3463 2433
rect 3467 2429 3468 2433
rect 3462 2428 3468 2429
rect 3614 2433 3620 2434
rect 3614 2429 3615 2433
rect 3619 2429 3620 2433
rect 3614 2428 3620 2429
rect 3766 2433 3772 2434
rect 3766 2429 3767 2433
rect 3771 2429 3772 2433
rect 3766 2428 3772 2429
rect 3894 2433 3900 2434
rect 3894 2429 3895 2433
rect 3899 2429 3900 2433
rect 3894 2428 3900 2429
rect 1283 2424 1382 2426
rect 1283 2423 1284 2424
rect 1278 2422 1284 2423
rect 2695 2423 2701 2424
rect 2695 2419 2696 2423
rect 2700 2422 2701 2423
rect 2727 2423 2733 2424
rect 2727 2422 2728 2423
rect 2700 2420 2728 2422
rect 2700 2419 2701 2420
rect 2695 2418 2701 2419
rect 2727 2419 2728 2420
rect 2732 2419 2733 2423
rect 2727 2418 2733 2419
rect 2790 2423 2796 2424
rect 2790 2419 2791 2423
rect 2795 2422 2796 2423
rect 2815 2423 2821 2424
rect 2815 2422 2816 2423
rect 2795 2420 2816 2422
rect 2795 2419 2796 2420
rect 2790 2418 2796 2419
rect 2815 2419 2816 2420
rect 2820 2419 2821 2423
rect 2815 2418 2821 2419
rect 2943 2423 2949 2424
rect 2943 2419 2944 2423
rect 2948 2422 2949 2423
rect 2999 2423 3005 2424
rect 2999 2422 3000 2423
rect 2948 2420 3000 2422
rect 2948 2419 2949 2420
rect 2943 2418 2949 2419
rect 2999 2419 3000 2420
rect 3004 2419 3005 2423
rect 2999 2418 3005 2419
rect 3087 2423 3093 2424
rect 3087 2419 3088 2423
rect 3092 2422 3093 2423
rect 3143 2423 3149 2424
rect 3143 2422 3144 2423
rect 3092 2420 3144 2422
rect 3092 2419 3093 2420
rect 3087 2418 3093 2419
rect 3143 2419 3144 2420
rect 3148 2419 3149 2423
rect 3143 2418 3149 2419
rect 3231 2423 3237 2424
rect 3231 2419 3232 2423
rect 3236 2422 3237 2423
rect 3295 2423 3301 2424
rect 3295 2422 3296 2423
rect 3236 2420 3296 2422
rect 3236 2419 3237 2420
rect 3231 2418 3237 2419
rect 3295 2419 3296 2420
rect 3300 2419 3301 2423
rect 3383 2423 3389 2424
rect 3383 2422 3384 2423
rect 3295 2418 3301 2419
rect 3304 2420 3384 2422
rect 399 2415 405 2416
rect 399 2411 400 2415
rect 404 2414 405 2415
rect 455 2415 461 2416
rect 455 2414 456 2415
rect 404 2412 456 2414
rect 404 2411 405 2412
rect 399 2410 405 2411
rect 455 2411 456 2412
rect 460 2411 461 2415
rect 455 2410 461 2411
rect 543 2415 549 2416
rect 543 2411 544 2415
rect 548 2414 549 2415
rect 607 2415 613 2416
rect 607 2414 608 2415
rect 548 2412 608 2414
rect 548 2411 549 2412
rect 543 2410 549 2411
rect 607 2411 608 2412
rect 612 2411 613 2415
rect 607 2410 613 2411
rect 678 2415 684 2416
rect 678 2411 679 2415
rect 683 2414 684 2415
rect 695 2415 701 2416
rect 695 2414 696 2415
rect 683 2412 696 2414
rect 683 2411 684 2412
rect 678 2410 684 2411
rect 695 2411 696 2412
rect 700 2411 701 2415
rect 695 2410 701 2411
rect 855 2415 861 2416
rect 855 2411 856 2415
rect 860 2414 861 2415
rect 927 2415 933 2416
rect 927 2414 928 2415
rect 860 2412 928 2414
rect 860 2411 861 2412
rect 855 2410 861 2411
rect 927 2411 928 2412
rect 932 2411 933 2415
rect 927 2410 933 2411
rect 1006 2415 1012 2416
rect 1006 2411 1007 2415
rect 1011 2414 1012 2415
rect 1015 2415 1021 2416
rect 1015 2414 1016 2415
rect 1011 2412 1016 2414
rect 1011 2411 1012 2412
rect 1006 2410 1012 2411
rect 1015 2411 1016 2412
rect 1020 2411 1021 2415
rect 1015 2410 1021 2411
rect 1167 2415 1173 2416
rect 1167 2411 1168 2415
rect 1172 2414 1173 2415
rect 1183 2415 1189 2416
rect 1183 2414 1184 2415
rect 1172 2412 1184 2414
rect 1172 2411 1173 2412
rect 1167 2410 1173 2411
rect 1183 2411 1184 2412
rect 1188 2411 1189 2415
rect 1319 2415 1325 2416
rect 1319 2414 1320 2415
rect 1183 2410 1189 2411
rect 1232 2412 1320 2414
rect 326 2407 332 2408
rect 326 2403 327 2407
rect 331 2403 332 2407
rect 326 2402 332 2403
rect 470 2407 476 2408
rect 470 2403 471 2407
rect 475 2403 476 2407
rect 470 2402 476 2403
rect 622 2407 628 2408
rect 622 2403 623 2407
rect 627 2403 628 2407
rect 622 2402 628 2403
rect 782 2407 788 2408
rect 782 2403 783 2407
rect 787 2403 788 2407
rect 782 2402 788 2403
rect 942 2407 948 2408
rect 942 2403 943 2407
rect 947 2403 948 2407
rect 942 2402 948 2403
rect 1094 2407 1100 2408
rect 1094 2403 1095 2407
rect 1099 2403 1100 2407
rect 1232 2406 1234 2412
rect 1319 2411 1320 2412
rect 1324 2411 1325 2415
rect 1319 2410 1325 2411
rect 1370 2415 1381 2416
rect 1370 2411 1371 2415
rect 1375 2411 1376 2415
rect 1380 2411 1381 2415
rect 1463 2415 1469 2416
rect 1463 2414 1464 2415
rect 1370 2410 1381 2411
rect 1384 2412 1464 2414
rect 1094 2402 1100 2403
rect 1159 2404 1234 2406
rect 1246 2407 1252 2408
rect 686 2399 692 2400
rect 350 2395 356 2396
rect 350 2391 351 2395
rect 355 2391 356 2395
rect 686 2395 687 2399
rect 691 2398 692 2399
rect 1159 2398 1161 2404
rect 1246 2403 1247 2407
rect 1251 2403 1252 2407
rect 1384 2406 1386 2412
rect 1463 2411 1464 2412
rect 1468 2411 1469 2415
rect 1463 2410 1469 2411
rect 1607 2415 1613 2416
rect 1607 2411 1608 2415
rect 1612 2414 1613 2415
rect 1655 2415 1661 2416
rect 1655 2414 1656 2415
rect 1612 2412 1656 2414
rect 1612 2411 1613 2412
rect 1607 2410 1613 2411
rect 1655 2411 1656 2412
rect 1660 2411 1661 2415
rect 1655 2410 1661 2411
rect 1694 2415 1700 2416
rect 1694 2411 1695 2415
rect 1699 2414 1700 2415
rect 1743 2415 1749 2416
rect 1743 2414 1744 2415
rect 1699 2412 1744 2414
rect 1699 2411 1700 2412
rect 1694 2410 1700 2411
rect 1743 2411 1744 2412
rect 1748 2411 1749 2415
rect 1743 2410 1749 2411
rect 1887 2415 1896 2416
rect 1887 2411 1888 2415
rect 1895 2411 1896 2415
rect 2007 2415 2013 2416
rect 2007 2414 2008 2415
rect 1887 2410 1896 2411
rect 1904 2412 2008 2414
rect 1246 2402 1252 2403
rect 1352 2404 1386 2406
rect 1390 2407 1396 2408
rect 1352 2398 1354 2404
rect 1390 2403 1391 2407
rect 1395 2403 1396 2407
rect 1390 2402 1396 2403
rect 1534 2407 1540 2408
rect 1534 2403 1535 2407
rect 1539 2403 1540 2407
rect 1534 2402 1540 2403
rect 1670 2407 1676 2408
rect 1670 2403 1671 2407
rect 1675 2403 1676 2407
rect 1670 2402 1676 2403
rect 1814 2407 1820 2408
rect 1814 2403 1815 2407
rect 1819 2403 1820 2407
rect 1814 2402 1820 2403
rect 1904 2398 1906 2412
rect 2007 2411 2008 2412
rect 2012 2411 2013 2415
rect 2007 2410 2013 2411
rect 2894 2415 2900 2416
rect 2894 2411 2895 2415
rect 2899 2414 2900 2415
rect 3304 2414 3306 2420
rect 3383 2419 3384 2420
rect 3388 2419 3389 2423
rect 3383 2418 3389 2419
rect 3535 2423 3541 2424
rect 3535 2419 3536 2423
rect 3540 2422 3541 2423
rect 3599 2423 3605 2424
rect 3599 2422 3600 2423
rect 3540 2420 3600 2422
rect 3540 2419 3541 2420
rect 3535 2418 3541 2419
rect 3599 2419 3600 2420
rect 3604 2419 3605 2423
rect 3599 2418 3605 2419
rect 3686 2423 3693 2424
rect 3686 2419 3687 2423
rect 3692 2419 3693 2423
rect 3839 2423 3845 2424
rect 3839 2422 3840 2423
rect 3686 2418 3693 2419
rect 3760 2420 3840 2422
rect 2899 2412 3306 2414
rect 3566 2415 3572 2416
rect 2899 2411 2900 2412
rect 2894 2410 2900 2411
rect 3566 2411 3567 2415
rect 3571 2414 3572 2415
rect 3760 2414 3762 2420
rect 3839 2419 3840 2420
rect 3844 2419 3845 2423
rect 3839 2418 3845 2419
rect 3878 2423 3884 2424
rect 3878 2419 3879 2423
rect 3883 2422 3884 2423
rect 3967 2423 3973 2424
rect 3967 2422 3968 2423
rect 3883 2420 3968 2422
rect 3883 2419 3884 2420
rect 3878 2418 3884 2419
rect 3967 2419 3968 2420
rect 3972 2419 3973 2423
rect 3967 2418 3973 2419
rect 3571 2412 3762 2414
rect 3571 2411 3572 2412
rect 3566 2410 3572 2411
rect 1934 2407 1940 2408
rect 1934 2403 1935 2407
rect 1939 2403 1940 2407
rect 1934 2402 1940 2403
rect 2582 2407 2588 2408
rect 2582 2403 2583 2407
rect 2587 2406 2588 2407
rect 3038 2407 3044 2408
rect 2587 2404 2690 2406
rect 2587 2403 2588 2404
rect 2582 2402 2588 2403
rect 2671 2400 2677 2401
rect 2006 2399 2012 2400
rect 2006 2398 2007 2399
rect 691 2396 777 2398
rect 1145 2396 1161 2398
rect 1297 2396 1354 2398
rect 1865 2396 1906 2398
rect 1985 2396 2007 2398
rect 691 2395 692 2396
rect 686 2394 692 2395
rect 1526 2395 1532 2396
rect 350 2390 356 2391
rect 1526 2391 1527 2395
rect 1531 2391 1532 2395
rect 2006 2395 2007 2396
rect 2011 2395 2012 2399
rect 2006 2394 2012 2395
rect 2559 2399 2565 2400
rect 2559 2395 2560 2399
rect 2564 2398 2565 2399
rect 2583 2399 2589 2400
rect 2583 2398 2584 2399
rect 2564 2396 2584 2398
rect 2564 2395 2565 2396
rect 2559 2394 2565 2395
rect 2583 2395 2584 2396
rect 2588 2395 2589 2399
rect 2583 2394 2589 2395
rect 2662 2399 2668 2400
rect 2662 2395 2663 2399
rect 2667 2398 2668 2399
rect 2671 2398 2672 2400
rect 2667 2396 2672 2398
rect 2676 2396 2677 2400
rect 2688 2398 2690 2404
rect 3038 2403 3039 2407
rect 3043 2406 3044 2407
rect 3043 2404 3450 2406
rect 3043 2403 3044 2404
rect 3038 2402 3044 2403
rect 2799 2399 2805 2400
rect 2799 2398 2800 2399
rect 2688 2396 2800 2398
rect 2667 2395 2668 2396
rect 2671 2395 2677 2396
rect 2799 2395 2800 2396
rect 2804 2395 2805 2399
rect 2662 2394 2668 2395
rect 2799 2394 2805 2395
rect 2942 2399 2948 2400
rect 2942 2395 2943 2399
rect 2947 2398 2948 2399
rect 2951 2399 2957 2400
rect 2951 2398 2952 2399
rect 2947 2396 2952 2398
rect 2947 2395 2948 2396
rect 2942 2394 2948 2395
rect 2951 2395 2952 2396
rect 2956 2395 2957 2399
rect 2951 2394 2957 2395
rect 3127 2399 3133 2400
rect 3127 2395 3128 2399
rect 3132 2398 3133 2399
rect 3231 2399 3237 2400
rect 3231 2398 3232 2399
rect 3132 2396 3232 2398
rect 3132 2395 3133 2396
rect 3127 2394 3133 2395
rect 3231 2395 3232 2396
rect 3236 2395 3237 2399
rect 3231 2394 3237 2395
rect 3319 2399 3325 2400
rect 3319 2395 3320 2399
rect 3324 2398 3325 2399
rect 3439 2399 3445 2400
rect 3439 2398 3440 2399
rect 3324 2396 3440 2398
rect 3324 2395 3325 2396
rect 3319 2394 3325 2395
rect 3439 2395 3440 2396
rect 3444 2395 3445 2399
rect 3448 2398 3450 2404
rect 3527 2399 3533 2400
rect 3527 2398 3528 2399
rect 3448 2396 3528 2398
rect 3439 2394 3445 2395
rect 3527 2395 3528 2396
rect 3532 2395 3533 2399
rect 3527 2394 3533 2395
rect 3751 2399 3757 2400
rect 3751 2395 3752 2399
rect 3756 2398 3757 2399
rect 3759 2399 3765 2400
rect 3759 2398 3760 2399
rect 3756 2396 3760 2398
rect 3756 2395 3757 2396
rect 3751 2394 3757 2395
rect 3759 2395 3760 2396
rect 3764 2395 3765 2399
rect 3759 2394 3765 2395
rect 3966 2399 3973 2400
rect 3966 2395 3967 2399
rect 3972 2395 3973 2399
rect 3966 2394 3973 2395
rect 1526 2390 1532 2391
rect 2486 2391 2492 2392
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 2030 2388 2036 2389
rect 2030 2384 2031 2388
rect 2035 2384 2036 2388
rect 2486 2387 2487 2391
rect 2491 2387 2492 2391
rect 2486 2386 2492 2387
rect 2598 2391 2604 2392
rect 2598 2387 2599 2391
rect 2603 2387 2604 2391
rect 2598 2386 2604 2387
rect 2726 2391 2732 2392
rect 2726 2387 2727 2391
rect 2731 2387 2732 2391
rect 2726 2386 2732 2387
rect 2878 2391 2884 2392
rect 2878 2387 2879 2391
rect 2883 2387 2884 2391
rect 2878 2386 2884 2387
rect 3054 2391 3060 2392
rect 3054 2387 3055 2391
rect 3059 2387 3060 2391
rect 3054 2386 3060 2387
rect 3246 2391 3252 2392
rect 3246 2387 3247 2391
rect 3251 2387 3252 2391
rect 3246 2386 3252 2387
rect 3454 2391 3460 2392
rect 3454 2387 3455 2391
rect 3459 2387 3460 2391
rect 3454 2386 3460 2387
rect 3678 2391 3684 2392
rect 3678 2387 3679 2391
rect 3683 2387 3684 2391
rect 3678 2386 3684 2387
rect 3894 2391 3900 2392
rect 3894 2387 3895 2391
rect 3899 2387 3900 2391
rect 3894 2386 3900 2387
rect 2030 2383 2036 2384
rect 2582 2383 2588 2384
rect 2582 2382 2583 2383
rect 2537 2380 2583 2382
rect 2582 2379 2583 2380
rect 2587 2379 2588 2383
rect 2790 2383 2796 2384
rect 2790 2382 2791 2383
rect 2777 2380 2791 2382
rect 2582 2378 2588 2379
rect 2790 2379 2791 2380
rect 2795 2379 2796 2383
rect 3038 2383 3044 2384
rect 3038 2382 3039 2383
rect 2929 2380 3039 2382
rect 2790 2378 2796 2379
rect 3038 2379 3039 2380
rect 3043 2379 3044 2383
rect 3118 2383 3124 2384
rect 3118 2382 3119 2383
rect 3105 2380 3119 2382
rect 3038 2378 3044 2379
rect 3118 2379 3119 2380
rect 3123 2379 3124 2383
rect 3958 2383 3964 2384
rect 3958 2382 3959 2383
rect 3945 2380 3959 2382
rect 3118 2378 3124 2379
rect 3686 2379 3692 2380
rect 3686 2375 3687 2379
rect 3691 2375 3692 2379
rect 3958 2379 3959 2380
rect 3963 2379 3964 2383
rect 3958 2378 3964 2379
rect 3686 2374 3692 2375
rect 2070 2372 2076 2373
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 2030 2371 2036 2372
rect 2030 2367 2031 2371
rect 2035 2367 2036 2371
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 3990 2372 3996 2373
rect 3990 2368 3991 2372
rect 3995 2368 3996 2372
rect 3990 2367 3996 2368
rect 110 2366 116 2367
rect 326 2366 332 2367
rect 326 2362 327 2366
rect 331 2362 332 2366
rect 326 2361 332 2362
rect 470 2366 476 2367
rect 470 2362 471 2366
rect 475 2362 476 2366
rect 470 2361 476 2362
rect 622 2366 628 2367
rect 622 2362 623 2366
rect 627 2362 628 2366
rect 622 2361 628 2362
rect 782 2366 788 2367
rect 782 2362 783 2366
rect 787 2362 788 2366
rect 782 2361 788 2362
rect 942 2366 948 2367
rect 942 2362 943 2366
rect 947 2362 948 2366
rect 942 2361 948 2362
rect 1094 2366 1100 2367
rect 1094 2362 1095 2366
rect 1099 2362 1100 2366
rect 1094 2361 1100 2362
rect 1246 2366 1252 2367
rect 1246 2362 1247 2366
rect 1251 2362 1252 2366
rect 1246 2361 1252 2362
rect 1390 2366 1396 2367
rect 1390 2362 1391 2366
rect 1395 2362 1396 2366
rect 1390 2361 1396 2362
rect 1534 2366 1540 2367
rect 1534 2362 1535 2366
rect 1539 2362 1540 2366
rect 1534 2361 1540 2362
rect 1670 2366 1676 2367
rect 1670 2362 1671 2366
rect 1675 2362 1676 2366
rect 1670 2361 1676 2362
rect 1814 2366 1820 2367
rect 1814 2362 1815 2366
rect 1819 2362 1820 2366
rect 1814 2361 1820 2362
rect 1934 2366 1940 2367
rect 2030 2366 2036 2367
rect 1934 2362 1935 2366
rect 1939 2362 1940 2366
rect 1934 2361 1940 2362
rect 2070 2355 2076 2356
rect 2070 2351 2071 2355
rect 2075 2351 2076 2355
rect 3990 2355 3996 2356
rect 3990 2351 3991 2355
rect 3995 2351 3996 2355
rect 2070 2350 2076 2351
rect 2486 2350 2492 2351
rect 2486 2346 2487 2350
rect 2491 2346 2492 2350
rect 2486 2345 2492 2346
rect 2598 2350 2604 2351
rect 2598 2346 2599 2350
rect 2603 2346 2604 2350
rect 2598 2345 2604 2346
rect 2726 2350 2732 2351
rect 2726 2346 2727 2350
rect 2731 2346 2732 2350
rect 2726 2345 2732 2346
rect 2878 2350 2884 2351
rect 2878 2346 2879 2350
rect 2883 2346 2884 2350
rect 2878 2345 2884 2346
rect 3054 2350 3060 2351
rect 3054 2346 3055 2350
rect 3059 2346 3060 2350
rect 3054 2345 3060 2346
rect 3246 2350 3252 2351
rect 3246 2346 3247 2350
rect 3251 2346 3252 2350
rect 3246 2345 3252 2346
rect 3454 2350 3460 2351
rect 3454 2346 3455 2350
rect 3459 2346 3460 2350
rect 3454 2345 3460 2346
rect 3678 2350 3684 2351
rect 3678 2346 3679 2350
rect 3683 2346 3684 2350
rect 3678 2345 3684 2346
rect 3894 2350 3900 2351
rect 3990 2350 3996 2351
rect 3894 2346 3895 2350
rect 3899 2346 3900 2350
rect 3894 2345 3900 2346
rect 358 2326 364 2327
rect 358 2322 359 2326
rect 363 2322 364 2326
rect 110 2321 116 2322
rect 358 2321 364 2322
rect 494 2326 500 2327
rect 494 2322 495 2326
rect 499 2322 500 2326
rect 494 2321 500 2322
rect 638 2326 644 2327
rect 638 2322 639 2326
rect 643 2322 644 2326
rect 638 2321 644 2322
rect 782 2326 788 2327
rect 782 2322 783 2326
rect 787 2322 788 2326
rect 782 2321 788 2322
rect 934 2326 940 2327
rect 934 2322 935 2326
rect 939 2322 940 2326
rect 934 2321 940 2322
rect 1086 2326 1092 2327
rect 1086 2322 1087 2326
rect 1091 2322 1092 2326
rect 1086 2321 1092 2322
rect 1246 2326 1252 2327
rect 1246 2322 1247 2326
rect 1251 2322 1252 2326
rect 1246 2321 1252 2322
rect 1414 2326 1420 2327
rect 1414 2322 1415 2326
rect 1419 2322 1420 2326
rect 1414 2321 1420 2322
rect 1590 2326 1596 2327
rect 1590 2322 1591 2326
rect 1595 2322 1596 2326
rect 1590 2321 1596 2322
rect 1774 2326 1780 2327
rect 1774 2322 1775 2326
rect 1779 2322 1780 2326
rect 1774 2321 1780 2322
rect 1934 2326 1940 2327
rect 1934 2322 1935 2326
rect 1939 2322 1940 2326
rect 1934 2321 1940 2322
rect 2030 2321 2036 2322
rect 110 2317 111 2321
rect 115 2317 116 2321
rect 110 2316 116 2317
rect 2030 2317 2031 2321
rect 2035 2317 2036 2321
rect 2030 2316 2036 2317
rect 2110 2306 2116 2307
rect 110 2304 116 2305
rect 110 2300 111 2304
rect 115 2300 116 2304
rect 110 2299 116 2300
rect 2030 2304 2036 2305
rect 2030 2300 2031 2304
rect 2035 2300 2036 2304
rect 2110 2302 2111 2306
rect 2115 2302 2116 2306
rect 2030 2299 2036 2300
rect 2070 2301 2076 2302
rect 2110 2301 2116 2302
rect 2222 2306 2228 2307
rect 2222 2302 2223 2306
rect 2227 2302 2228 2306
rect 2222 2301 2228 2302
rect 2358 2306 2364 2307
rect 2358 2302 2359 2306
rect 2363 2302 2364 2306
rect 2358 2301 2364 2302
rect 2510 2306 2516 2307
rect 2510 2302 2511 2306
rect 2515 2302 2516 2306
rect 2510 2301 2516 2302
rect 2670 2306 2676 2307
rect 2670 2302 2671 2306
rect 2675 2302 2676 2306
rect 2670 2301 2676 2302
rect 2846 2306 2852 2307
rect 2846 2302 2847 2306
rect 2851 2302 2852 2306
rect 2846 2301 2852 2302
rect 3038 2306 3044 2307
rect 3038 2302 3039 2306
rect 3043 2302 3044 2306
rect 3038 2301 3044 2302
rect 3246 2306 3252 2307
rect 3246 2302 3247 2306
rect 3251 2302 3252 2306
rect 3246 2301 3252 2302
rect 3462 2306 3468 2307
rect 3462 2302 3463 2306
rect 3467 2302 3468 2306
rect 3462 2301 3468 2302
rect 3686 2306 3692 2307
rect 3686 2302 3687 2306
rect 3691 2302 3692 2306
rect 3686 2301 3692 2302
rect 3894 2306 3900 2307
rect 3894 2302 3895 2306
rect 3899 2302 3900 2306
rect 3894 2301 3900 2302
rect 3990 2301 3996 2302
rect 2070 2297 2071 2301
rect 2075 2297 2076 2301
rect 2070 2296 2076 2297
rect 3990 2297 3991 2301
rect 3995 2297 3996 2301
rect 3990 2296 3996 2297
rect 478 2295 484 2296
rect 478 2294 479 2295
rect 409 2292 479 2294
rect 478 2291 479 2292
rect 483 2291 484 2295
rect 766 2295 772 2296
rect 766 2294 767 2295
rect 689 2292 767 2294
rect 478 2290 484 2291
rect 766 2291 767 2292
rect 771 2291 772 2295
rect 918 2295 924 2296
rect 918 2294 919 2295
rect 833 2292 919 2294
rect 766 2290 772 2291
rect 918 2291 919 2292
rect 923 2291 924 2295
rect 1006 2295 1012 2296
rect 1006 2294 1007 2295
rect 985 2292 1007 2294
rect 918 2290 924 2291
rect 1006 2291 1007 2292
rect 1011 2291 1012 2295
rect 1175 2295 1181 2296
rect 1175 2294 1176 2295
rect 1137 2292 1176 2294
rect 1006 2290 1012 2291
rect 1175 2291 1176 2292
rect 1180 2291 1181 2295
rect 1175 2290 1181 2291
rect 1183 2295 1189 2296
rect 1183 2291 1184 2295
rect 1188 2294 1189 2295
rect 1574 2295 1580 2296
rect 1574 2294 1575 2295
rect 1188 2292 1241 2294
rect 1465 2292 1575 2294
rect 1188 2291 1189 2292
rect 1183 2290 1189 2291
rect 1574 2291 1575 2292
rect 1579 2291 1580 2295
rect 1758 2295 1764 2296
rect 1758 2294 1759 2295
rect 1641 2292 1759 2294
rect 1574 2290 1580 2291
rect 1758 2291 1759 2292
rect 1763 2291 1764 2295
rect 1758 2290 1764 2291
rect 1766 2295 1772 2296
rect 1766 2291 1767 2295
rect 1771 2291 1772 2295
rect 2182 2295 2188 2296
rect 2182 2294 2183 2295
rect 1985 2292 2183 2294
rect 1766 2290 1772 2291
rect 2182 2291 2183 2292
rect 2187 2291 2188 2295
rect 2182 2290 2188 2291
rect 358 2285 364 2286
rect 358 2281 359 2285
rect 363 2281 364 2285
rect 358 2280 364 2281
rect 494 2285 500 2286
rect 494 2281 495 2285
rect 499 2281 500 2285
rect 494 2280 500 2281
rect 638 2285 644 2286
rect 638 2281 639 2285
rect 643 2281 644 2285
rect 638 2280 644 2281
rect 782 2285 788 2286
rect 782 2281 783 2285
rect 787 2281 788 2285
rect 782 2280 788 2281
rect 934 2285 940 2286
rect 934 2281 935 2285
rect 939 2281 940 2285
rect 934 2280 940 2281
rect 1086 2285 1092 2286
rect 1086 2281 1087 2285
rect 1091 2281 1092 2285
rect 1086 2280 1092 2281
rect 1246 2285 1252 2286
rect 1246 2281 1247 2285
rect 1251 2281 1252 2285
rect 1246 2280 1252 2281
rect 1414 2285 1420 2286
rect 1414 2281 1415 2285
rect 1419 2281 1420 2285
rect 1414 2280 1420 2281
rect 1590 2285 1596 2286
rect 1590 2281 1591 2285
rect 1595 2281 1596 2285
rect 1590 2280 1596 2281
rect 1774 2285 1780 2286
rect 1774 2281 1775 2285
rect 1779 2281 1780 2285
rect 1774 2280 1780 2281
rect 1934 2285 1940 2286
rect 1934 2281 1935 2285
rect 1939 2281 1940 2285
rect 1934 2280 1940 2281
rect 2070 2284 2076 2285
rect 2070 2280 2071 2284
rect 2075 2280 2076 2284
rect 2070 2279 2076 2280
rect 3990 2284 3996 2285
rect 3990 2280 3991 2284
rect 3995 2280 3996 2284
rect 3990 2279 3996 2280
rect 431 2275 437 2276
rect 431 2271 432 2275
rect 436 2274 437 2275
rect 479 2275 485 2276
rect 479 2274 480 2275
rect 436 2272 480 2274
rect 436 2271 437 2272
rect 431 2270 437 2271
rect 479 2271 480 2272
rect 484 2271 485 2275
rect 479 2270 485 2271
rect 567 2275 573 2276
rect 567 2271 568 2275
rect 572 2274 573 2275
rect 686 2275 692 2276
rect 686 2274 687 2275
rect 572 2272 687 2274
rect 572 2271 573 2272
rect 567 2270 573 2271
rect 686 2271 687 2272
rect 691 2271 692 2275
rect 686 2270 692 2271
rect 702 2275 708 2276
rect 702 2271 703 2275
rect 707 2274 708 2275
rect 711 2275 717 2276
rect 711 2274 712 2275
rect 707 2272 712 2274
rect 707 2271 708 2272
rect 702 2270 708 2271
rect 711 2271 712 2272
rect 716 2271 717 2275
rect 711 2270 717 2271
rect 766 2275 772 2276
rect 766 2271 767 2275
rect 771 2274 772 2275
rect 855 2275 861 2276
rect 855 2274 856 2275
rect 771 2272 856 2274
rect 771 2271 772 2272
rect 766 2270 772 2271
rect 855 2271 856 2272
rect 860 2271 861 2275
rect 855 2270 861 2271
rect 918 2275 924 2276
rect 918 2271 919 2275
rect 923 2274 924 2275
rect 1007 2275 1013 2276
rect 1007 2274 1008 2275
rect 923 2272 1008 2274
rect 923 2271 924 2272
rect 918 2270 924 2271
rect 1007 2271 1008 2272
rect 1012 2271 1013 2275
rect 1007 2270 1013 2271
rect 1094 2275 1100 2276
rect 1094 2271 1095 2275
rect 1099 2274 1100 2275
rect 1159 2275 1165 2276
rect 1159 2274 1160 2275
rect 1099 2272 1160 2274
rect 1099 2271 1100 2272
rect 1094 2270 1100 2271
rect 1159 2271 1160 2272
rect 1164 2271 1165 2275
rect 1159 2270 1165 2271
rect 1175 2275 1181 2276
rect 1175 2271 1176 2275
rect 1180 2274 1181 2275
rect 1319 2275 1325 2276
rect 1319 2274 1320 2275
rect 1180 2272 1320 2274
rect 1180 2271 1181 2272
rect 1175 2270 1181 2271
rect 1319 2271 1320 2272
rect 1324 2271 1325 2275
rect 1319 2270 1325 2271
rect 1487 2275 1493 2276
rect 1487 2271 1488 2275
rect 1492 2274 1493 2275
rect 1526 2275 1532 2276
rect 1526 2274 1527 2275
rect 1492 2272 1527 2274
rect 1492 2271 1493 2272
rect 1487 2270 1493 2271
rect 1526 2271 1527 2272
rect 1531 2271 1532 2275
rect 1526 2270 1532 2271
rect 1574 2275 1580 2276
rect 1574 2271 1575 2275
rect 1579 2274 1580 2275
rect 1663 2275 1669 2276
rect 1663 2274 1664 2275
rect 1579 2272 1664 2274
rect 1579 2271 1580 2272
rect 1574 2270 1580 2271
rect 1663 2271 1664 2272
rect 1668 2271 1669 2275
rect 1663 2270 1669 2271
rect 1758 2275 1764 2276
rect 1758 2271 1759 2275
rect 1763 2274 1764 2275
rect 1847 2275 1853 2276
rect 1847 2274 1848 2275
rect 1763 2272 1848 2274
rect 1763 2271 1764 2272
rect 1758 2270 1764 2271
rect 1847 2271 1848 2272
rect 1852 2271 1853 2275
rect 1847 2270 1853 2271
rect 2006 2275 2013 2276
rect 2006 2271 2007 2275
rect 2012 2271 2013 2275
rect 2494 2275 2500 2276
rect 2494 2274 2495 2275
rect 2161 2272 2202 2274
rect 2409 2272 2495 2274
rect 2006 2270 2013 2271
rect 2110 2265 2116 2266
rect 2110 2261 2111 2265
rect 2115 2261 2116 2265
rect 2110 2260 2116 2261
rect 2200 2262 2202 2272
rect 2494 2271 2495 2272
rect 2499 2271 2500 2275
rect 2654 2275 2660 2276
rect 2654 2274 2655 2275
rect 2561 2272 2655 2274
rect 2494 2270 2500 2271
rect 2654 2271 2655 2272
rect 2659 2271 2660 2275
rect 2654 2270 2660 2271
rect 2662 2275 2668 2276
rect 2662 2271 2663 2275
rect 2667 2271 2668 2275
rect 3022 2275 3028 2276
rect 3022 2274 3023 2275
rect 2897 2272 3023 2274
rect 2662 2270 2668 2271
rect 3022 2271 3023 2272
rect 3027 2271 3028 2275
rect 3759 2275 3765 2276
rect 3759 2274 3760 2275
rect 3737 2272 3760 2274
rect 3022 2270 3028 2271
rect 3759 2271 3760 2272
rect 3764 2271 3765 2275
rect 3966 2275 3972 2276
rect 3966 2274 3967 2275
rect 3945 2272 3967 2274
rect 3759 2270 3765 2271
rect 3966 2271 3967 2272
rect 3971 2271 3972 2275
rect 3966 2270 3972 2271
rect 2222 2265 2228 2266
rect 2200 2260 2218 2262
rect 2222 2261 2223 2265
rect 2227 2261 2228 2265
rect 2222 2260 2228 2261
rect 2358 2265 2364 2266
rect 2358 2261 2359 2265
rect 2363 2261 2364 2265
rect 2358 2260 2364 2261
rect 2510 2265 2516 2266
rect 2510 2261 2511 2265
rect 2515 2261 2516 2265
rect 2510 2260 2516 2261
rect 2670 2265 2676 2266
rect 2670 2261 2671 2265
rect 2675 2261 2676 2265
rect 2670 2260 2676 2261
rect 2846 2265 2852 2266
rect 2846 2261 2847 2265
rect 2851 2261 2852 2265
rect 2846 2260 2852 2261
rect 3038 2265 3044 2266
rect 3038 2261 3039 2265
rect 3043 2261 3044 2265
rect 3038 2260 3044 2261
rect 3246 2265 3252 2266
rect 3246 2261 3247 2265
rect 3251 2261 3252 2265
rect 3246 2260 3252 2261
rect 3462 2265 3468 2266
rect 3462 2261 3463 2265
rect 3467 2261 3468 2265
rect 3462 2260 3468 2261
rect 3686 2265 3692 2266
rect 3686 2261 3687 2265
rect 3691 2261 3692 2265
rect 3686 2260 3692 2261
rect 3894 2265 3900 2266
rect 3894 2261 3895 2265
rect 3899 2261 3900 2265
rect 3894 2260 3900 2261
rect 478 2259 484 2260
rect 478 2255 479 2259
rect 483 2258 484 2259
rect 483 2256 546 2258
rect 483 2255 484 2256
rect 478 2254 484 2255
rect 311 2251 317 2252
rect 311 2247 312 2251
rect 316 2250 317 2251
rect 375 2251 381 2252
rect 375 2250 376 2251
rect 316 2248 376 2250
rect 316 2247 317 2248
rect 311 2246 317 2247
rect 375 2247 376 2248
rect 380 2247 381 2251
rect 375 2246 381 2247
rect 463 2251 469 2252
rect 463 2247 464 2251
rect 468 2250 469 2251
rect 535 2251 541 2252
rect 535 2250 536 2251
rect 468 2248 536 2250
rect 468 2247 469 2248
rect 463 2246 469 2247
rect 535 2247 536 2248
rect 540 2247 541 2251
rect 544 2250 546 2256
rect 2182 2255 2189 2256
rect 623 2251 629 2252
rect 623 2250 624 2251
rect 544 2248 624 2250
rect 535 2246 541 2247
rect 623 2247 624 2248
rect 628 2247 629 2251
rect 623 2246 629 2247
rect 783 2251 789 2252
rect 783 2247 784 2251
rect 788 2250 789 2251
rect 855 2251 861 2252
rect 855 2250 856 2251
rect 788 2248 856 2250
rect 788 2247 789 2248
rect 783 2246 789 2247
rect 855 2247 856 2248
rect 860 2247 861 2251
rect 855 2246 861 2247
rect 918 2251 924 2252
rect 918 2247 919 2251
rect 923 2250 924 2251
rect 943 2251 949 2252
rect 943 2250 944 2251
rect 923 2248 944 2250
rect 923 2247 924 2248
rect 918 2246 924 2247
rect 943 2247 944 2248
rect 948 2247 949 2251
rect 943 2246 949 2247
rect 1103 2251 1109 2252
rect 1103 2247 1104 2251
rect 1108 2250 1109 2251
rect 1175 2251 1181 2252
rect 1175 2250 1176 2251
rect 1108 2248 1176 2250
rect 1108 2247 1109 2248
rect 1103 2246 1109 2247
rect 1175 2247 1176 2248
rect 1180 2247 1181 2251
rect 1175 2246 1181 2247
rect 1263 2251 1269 2252
rect 1263 2247 1264 2251
rect 1268 2250 1269 2251
rect 1343 2251 1349 2252
rect 1343 2250 1344 2251
rect 1268 2248 1344 2250
rect 1268 2247 1269 2248
rect 1263 2246 1269 2247
rect 1343 2247 1344 2248
rect 1348 2247 1349 2251
rect 1343 2246 1349 2247
rect 1406 2251 1412 2252
rect 1406 2247 1407 2251
rect 1411 2250 1412 2251
rect 1431 2251 1437 2252
rect 1431 2250 1432 2251
rect 1411 2248 1432 2250
rect 1411 2247 1412 2248
rect 1406 2246 1412 2247
rect 1431 2247 1432 2248
rect 1436 2247 1437 2251
rect 1431 2246 1437 2247
rect 1599 2251 1605 2252
rect 1599 2247 1600 2251
rect 1604 2250 1605 2251
rect 1679 2251 1685 2252
rect 1679 2250 1680 2251
rect 1604 2248 1680 2250
rect 1604 2247 1605 2248
rect 1599 2246 1605 2247
rect 1679 2247 1680 2248
rect 1684 2247 1685 2251
rect 1679 2246 1685 2247
rect 1766 2251 1773 2252
rect 1766 2247 1767 2251
rect 1772 2247 1773 2251
rect 2182 2251 2183 2255
rect 2188 2251 2189 2255
rect 2182 2250 2189 2251
rect 2191 2255 2197 2256
rect 2191 2251 2192 2255
rect 2196 2254 2197 2255
rect 2207 2255 2213 2256
rect 2207 2254 2208 2255
rect 2196 2252 2208 2254
rect 2196 2251 2197 2252
rect 2191 2250 2197 2251
rect 2207 2251 2208 2252
rect 2212 2251 2213 2255
rect 2216 2254 2218 2260
rect 2295 2255 2301 2256
rect 2295 2254 2296 2255
rect 2216 2252 2296 2254
rect 2207 2250 2213 2251
rect 2295 2251 2296 2252
rect 2300 2251 2301 2255
rect 2295 2250 2301 2251
rect 2431 2255 2440 2256
rect 2431 2251 2432 2255
rect 2439 2251 2440 2255
rect 2431 2250 2440 2251
rect 2494 2255 2500 2256
rect 2494 2251 2495 2255
rect 2499 2254 2500 2255
rect 2583 2255 2589 2256
rect 2583 2254 2584 2255
rect 2499 2252 2584 2254
rect 2499 2251 2500 2252
rect 2494 2250 2500 2251
rect 2583 2251 2584 2252
rect 2588 2251 2589 2255
rect 2583 2250 2589 2251
rect 2654 2255 2660 2256
rect 2654 2251 2655 2255
rect 2659 2254 2660 2255
rect 2743 2255 2749 2256
rect 2743 2254 2744 2255
rect 2659 2252 2744 2254
rect 2659 2251 2660 2252
rect 2654 2250 2660 2251
rect 2743 2251 2744 2252
rect 2748 2251 2749 2255
rect 2743 2250 2749 2251
rect 2919 2255 2925 2256
rect 2919 2251 2920 2255
rect 2924 2254 2925 2255
rect 3023 2255 3029 2256
rect 3023 2254 3024 2255
rect 2924 2252 3024 2254
rect 2924 2251 2925 2252
rect 2919 2250 2925 2251
rect 3023 2251 3024 2252
rect 3028 2251 3029 2255
rect 3023 2250 3029 2251
rect 3111 2255 3117 2256
rect 3111 2251 3112 2255
rect 3116 2251 3117 2255
rect 3111 2250 3117 2251
rect 3154 2255 3160 2256
rect 3154 2251 3155 2255
rect 3159 2254 3160 2255
rect 3231 2255 3237 2256
rect 3231 2254 3232 2255
rect 3159 2252 3232 2254
rect 3159 2251 3160 2252
rect 3154 2250 3160 2251
rect 3231 2251 3232 2252
rect 3236 2251 3237 2255
rect 3231 2250 3237 2251
rect 3319 2255 3325 2256
rect 3319 2251 3320 2255
rect 3324 2254 3325 2255
rect 3447 2255 3453 2256
rect 3447 2254 3448 2255
rect 3324 2252 3448 2254
rect 3324 2251 3325 2252
rect 3319 2250 3325 2251
rect 3447 2251 3448 2252
rect 3452 2251 3453 2255
rect 3535 2255 3541 2256
rect 3535 2254 3536 2255
rect 3447 2250 3453 2251
rect 3456 2252 3536 2254
rect 1766 2246 1773 2247
rect 3022 2247 3028 2248
rect 238 2243 244 2244
rect 238 2239 239 2243
rect 243 2239 244 2243
rect 238 2238 244 2239
rect 390 2243 396 2244
rect 390 2239 391 2243
rect 395 2239 396 2243
rect 390 2238 396 2239
rect 550 2243 556 2244
rect 550 2239 551 2243
rect 555 2239 556 2243
rect 550 2238 556 2239
rect 710 2243 716 2244
rect 710 2239 711 2243
rect 715 2239 716 2243
rect 710 2238 716 2239
rect 870 2243 876 2244
rect 870 2239 871 2243
rect 875 2239 876 2243
rect 870 2238 876 2239
rect 1030 2243 1036 2244
rect 1030 2239 1031 2243
rect 1035 2239 1036 2243
rect 1030 2238 1036 2239
rect 1190 2243 1196 2244
rect 1190 2239 1191 2243
rect 1195 2239 1196 2243
rect 1190 2238 1196 2239
rect 1358 2243 1364 2244
rect 1358 2239 1359 2243
rect 1363 2239 1364 2243
rect 1358 2238 1364 2239
rect 1526 2243 1532 2244
rect 1526 2239 1527 2243
rect 1531 2239 1532 2243
rect 1526 2238 1532 2239
rect 1694 2243 1700 2244
rect 1694 2239 1695 2243
rect 1699 2239 1700 2243
rect 3022 2243 3023 2247
rect 3027 2246 3028 2247
rect 3456 2246 3458 2252
rect 3535 2251 3536 2252
rect 3540 2251 3541 2255
rect 3535 2250 3541 2251
rect 3759 2255 3765 2256
rect 3759 2251 3760 2255
rect 3764 2254 3765 2255
rect 3770 2255 3776 2256
rect 3770 2254 3771 2255
rect 3764 2252 3771 2254
rect 3764 2251 3765 2252
rect 3759 2250 3765 2251
rect 3770 2251 3771 2252
rect 3775 2251 3776 2255
rect 3770 2250 3776 2251
rect 3958 2255 3964 2256
rect 3958 2251 3959 2255
rect 3963 2254 3964 2255
rect 3967 2255 3973 2256
rect 3967 2254 3968 2255
rect 3963 2252 3968 2254
rect 3963 2251 3964 2252
rect 3958 2250 3964 2251
rect 3967 2251 3968 2252
rect 3972 2251 3973 2255
rect 3967 2250 3973 2251
rect 3027 2244 3458 2246
rect 3027 2243 3028 2244
rect 3022 2242 3028 2243
rect 1694 2238 1700 2239
rect 222 2235 228 2236
rect 222 2231 223 2235
rect 227 2234 228 2235
rect 702 2235 708 2236
rect 227 2232 233 2234
rect 227 2231 228 2232
rect 222 2230 228 2231
rect 702 2231 703 2235
rect 707 2231 708 2235
rect 1094 2235 1100 2236
rect 1094 2234 1095 2235
rect 1081 2232 1095 2234
rect 702 2230 708 2231
rect 1094 2231 1095 2232
rect 1099 2231 1100 2235
rect 2183 2235 2189 2236
rect 1094 2230 1100 2231
rect 1534 2231 1540 2232
rect 1534 2227 1535 2231
rect 1539 2227 1540 2231
rect 2183 2231 2184 2235
rect 2188 2234 2189 2235
rect 2191 2235 2197 2236
rect 2191 2234 2192 2235
rect 2188 2232 2192 2234
rect 2188 2231 2189 2232
rect 2183 2230 2189 2231
rect 2191 2231 2192 2232
rect 2196 2231 2197 2235
rect 2351 2235 2357 2236
rect 2351 2234 2352 2235
rect 2191 2230 2197 2231
rect 2228 2232 2352 2234
rect 1534 2226 1540 2227
rect 2110 2227 2116 2228
rect 110 2224 116 2225
rect 110 2220 111 2224
rect 115 2220 116 2224
rect 110 2219 116 2220
rect 2030 2224 2036 2225
rect 2030 2220 2031 2224
rect 2035 2220 2036 2224
rect 2110 2223 2111 2227
rect 2115 2223 2116 2227
rect 2110 2222 2116 2223
rect 2030 2219 2036 2220
rect 2228 2218 2230 2232
rect 2351 2231 2352 2232
rect 2356 2231 2357 2235
rect 2351 2230 2357 2231
rect 2434 2235 2440 2236
rect 2434 2231 2435 2235
rect 2439 2234 2440 2235
rect 2463 2235 2469 2236
rect 2463 2234 2464 2235
rect 2439 2232 2464 2234
rect 2439 2231 2440 2232
rect 2434 2230 2440 2231
rect 2463 2231 2464 2232
rect 2468 2231 2469 2235
rect 2463 2230 2469 2231
rect 2551 2235 2557 2236
rect 2551 2231 2552 2235
rect 2556 2234 2557 2235
rect 2663 2235 2669 2236
rect 2663 2234 2664 2235
rect 2556 2232 2664 2234
rect 2556 2231 2557 2232
rect 2551 2230 2557 2231
rect 2663 2231 2664 2232
rect 2668 2231 2669 2235
rect 2663 2230 2669 2231
rect 2686 2235 2692 2236
rect 2686 2231 2687 2235
rect 2691 2234 2692 2235
rect 2751 2235 2757 2236
rect 2751 2234 2752 2235
rect 2691 2232 2752 2234
rect 2691 2231 2692 2232
rect 2686 2230 2692 2231
rect 2751 2231 2752 2232
rect 2756 2231 2757 2235
rect 2751 2230 2757 2231
rect 2951 2235 2957 2236
rect 2951 2231 2952 2235
rect 2956 2234 2957 2235
rect 3063 2235 3069 2236
rect 3063 2234 3064 2235
rect 2956 2232 3064 2234
rect 2956 2231 2957 2232
rect 2951 2230 2957 2231
rect 3063 2231 3064 2232
rect 3068 2231 3069 2235
rect 3063 2230 3069 2231
rect 3151 2235 3160 2236
rect 3151 2231 3152 2235
rect 3159 2231 3160 2235
rect 3351 2235 3357 2236
rect 3351 2234 3352 2235
rect 3260 2232 3352 2234
rect 3151 2230 3160 2231
rect 3258 2231 3264 2232
rect 2278 2227 2284 2228
rect 2278 2223 2279 2227
rect 2283 2223 2284 2227
rect 2278 2222 2284 2223
rect 2478 2227 2484 2228
rect 2478 2223 2479 2227
rect 2483 2223 2484 2227
rect 2478 2222 2484 2223
rect 2678 2227 2684 2228
rect 2678 2223 2679 2227
rect 2683 2223 2684 2227
rect 2678 2222 2684 2223
rect 2878 2227 2884 2228
rect 2878 2223 2879 2227
rect 2883 2223 2884 2227
rect 2878 2222 2884 2223
rect 3078 2227 3084 2228
rect 3078 2223 3079 2227
rect 3083 2223 3084 2227
rect 3258 2227 3259 2231
rect 3263 2227 3264 2231
rect 3351 2231 3352 2232
rect 3356 2231 3357 2235
rect 3559 2235 3565 2236
rect 3559 2234 3560 2235
rect 3351 2230 3357 2231
rect 3412 2232 3560 2234
rect 3258 2226 3264 2227
rect 3278 2227 3284 2228
rect 3078 2222 3084 2223
rect 3278 2223 3279 2227
rect 3283 2223 3284 2227
rect 3278 2222 3284 2223
rect 2390 2219 2396 2220
rect 2390 2218 2391 2219
rect 2161 2216 2230 2218
rect 2329 2216 2391 2218
rect 2390 2215 2391 2216
rect 2395 2215 2396 2219
rect 3062 2219 3068 2220
rect 3062 2218 3063 2219
rect 2929 2216 3063 2218
rect 2390 2214 2396 2215
rect 3062 2215 3063 2216
rect 3067 2215 3068 2219
rect 3412 2218 3414 2232
rect 3559 2231 3560 2232
rect 3564 2231 3565 2235
rect 3559 2230 3565 2231
rect 3718 2235 3724 2236
rect 3718 2231 3719 2235
rect 3723 2234 3724 2235
rect 3775 2235 3781 2236
rect 3775 2234 3776 2235
rect 3723 2232 3776 2234
rect 3723 2231 3724 2232
rect 3718 2230 3724 2231
rect 3775 2231 3776 2232
rect 3780 2231 3781 2235
rect 3775 2230 3781 2231
rect 3966 2235 3973 2236
rect 3966 2231 3967 2235
rect 3972 2231 3973 2235
rect 3966 2230 3973 2231
rect 3486 2227 3492 2228
rect 3486 2223 3487 2227
rect 3491 2223 3492 2227
rect 3486 2222 3492 2223
rect 3702 2227 3708 2228
rect 3702 2223 3703 2227
rect 3707 2223 3708 2227
rect 3702 2222 3708 2223
rect 3894 2227 3900 2228
rect 3894 2223 3895 2227
rect 3899 2223 3900 2227
rect 3894 2222 3900 2223
rect 3770 2219 3776 2220
rect 3770 2218 3771 2219
rect 3329 2216 3414 2218
rect 3753 2216 3771 2218
rect 3062 2214 3068 2215
rect 3478 2215 3484 2216
rect 3478 2211 3479 2215
rect 3483 2211 3484 2215
rect 3770 2215 3771 2216
rect 3775 2215 3776 2219
rect 3958 2219 3964 2220
rect 3958 2218 3959 2219
rect 3945 2216 3959 2218
rect 3770 2214 3776 2215
rect 3958 2215 3959 2216
rect 3963 2215 3964 2219
rect 3958 2214 3964 2215
rect 3478 2210 3484 2211
rect 2070 2208 2076 2209
rect 110 2207 116 2208
rect 110 2203 111 2207
rect 115 2203 116 2207
rect 2030 2207 2036 2208
rect 2030 2203 2031 2207
rect 2035 2203 2036 2207
rect 2070 2204 2071 2208
rect 2075 2204 2076 2208
rect 2070 2203 2076 2204
rect 3990 2208 3996 2209
rect 3990 2204 3991 2208
rect 3995 2204 3996 2208
rect 3990 2203 3996 2204
rect 110 2202 116 2203
rect 238 2202 244 2203
rect 238 2198 239 2202
rect 243 2198 244 2202
rect 238 2197 244 2198
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 550 2202 556 2203
rect 550 2198 551 2202
rect 555 2198 556 2202
rect 550 2197 556 2198
rect 710 2202 716 2203
rect 710 2198 711 2202
rect 715 2198 716 2202
rect 710 2197 716 2198
rect 870 2202 876 2203
rect 870 2198 871 2202
rect 875 2198 876 2202
rect 870 2197 876 2198
rect 1030 2202 1036 2203
rect 1030 2198 1031 2202
rect 1035 2198 1036 2202
rect 1030 2197 1036 2198
rect 1190 2202 1196 2203
rect 1190 2198 1191 2202
rect 1195 2198 1196 2202
rect 1190 2197 1196 2198
rect 1358 2202 1364 2203
rect 1358 2198 1359 2202
rect 1363 2198 1364 2202
rect 1358 2197 1364 2198
rect 1526 2202 1532 2203
rect 1526 2198 1527 2202
rect 1531 2198 1532 2202
rect 1526 2197 1532 2198
rect 1694 2202 1700 2203
rect 2030 2202 2036 2203
rect 1694 2198 1695 2202
rect 1699 2198 1700 2202
rect 1694 2197 1700 2198
rect 2070 2191 2076 2192
rect 2070 2187 2071 2191
rect 2075 2187 2076 2191
rect 3990 2191 3996 2192
rect 3990 2187 3991 2191
rect 3995 2187 3996 2191
rect 2070 2186 2076 2187
rect 2110 2186 2116 2187
rect 2110 2182 2111 2186
rect 2115 2182 2116 2186
rect 2110 2181 2116 2182
rect 2278 2186 2284 2187
rect 2278 2182 2279 2186
rect 2283 2182 2284 2186
rect 2278 2181 2284 2182
rect 2478 2186 2484 2187
rect 2478 2182 2479 2186
rect 2483 2182 2484 2186
rect 2478 2181 2484 2182
rect 2678 2186 2684 2187
rect 2678 2182 2679 2186
rect 2683 2182 2684 2186
rect 2678 2181 2684 2182
rect 2878 2186 2884 2187
rect 2878 2182 2879 2186
rect 2883 2182 2884 2186
rect 2878 2181 2884 2182
rect 3078 2186 3084 2187
rect 3078 2182 3079 2186
rect 3083 2182 3084 2186
rect 3078 2181 3084 2182
rect 3278 2186 3284 2187
rect 3278 2182 3279 2186
rect 3283 2182 3284 2186
rect 3278 2181 3284 2182
rect 3486 2186 3492 2187
rect 3486 2182 3487 2186
rect 3491 2182 3492 2186
rect 3486 2181 3492 2182
rect 3702 2186 3708 2187
rect 3702 2182 3703 2186
rect 3707 2182 3708 2186
rect 3702 2181 3708 2182
rect 3894 2186 3900 2187
rect 3990 2186 3996 2187
rect 3894 2182 3895 2186
rect 3899 2182 3900 2186
rect 3894 2181 3900 2182
rect 150 2158 156 2159
rect 150 2154 151 2158
rect 155 2154 156 2158
rect 110 2153 116 2154
rect 150 2153 156 2154
rect 318 2158 324 2159
rect 318 2154 319 2158
rect 323 2154 324 2158
rect 318 2153 324 2154
rect 510 2158 516 2159
rect 510 2154 511 2158
rect 515 2154 516 2158
rect 510 2153 516 2154
rect 702 2158 708 2159
rect 702 2154 703 2158
rect 707 2154 708 2158
rect 702 2153 708 2154
rect 894 2158 900 2159
rect 894 2154 895 2158
rect 899 2154 900 2158
rect 894 2153 900 2154
rect 1086 2158 1092 2159
rect 1086 2154 1087 2158
rect 1091 2154 1092 2158
rect 1086 2153 1092 2154
rect 1278 2158 1284 2159
rect 1278 2154 1279 2158
rect 1283 2154 1284 2158
rect 1278 2153 1284 2154
rect 1462 2158 1468 2159
rect 1462 2154 1463 2158
rect 1467 2154 1468 2158
rect 1462 2153 1468 2154
rect 1654 2158 1660 2159
rect 1654 2154 1655 2158
rect 1659 2154 1660 2158
rect 1654 2153 1660 2154
rect 1846 2158 1852 2159
rect 1846 2154 1847 2158
rect 1851 2154 1852 2158
rect 1846 2153 1852 2154
rect 2030 2153 2036 2154
rect 110 2149 111 2153
rect 115 2149 116 2153
rect 110 2148 116 2149
rect 2030 2149 2031 2153
rect 2035 2149 2036 2153
rect 2030 2148 2036 2149
rect 2142 2146 2148 2147
rect 2142 2142 2143 2146
rect 2147 2142 2148 2146
rect 2070 2141 2076 2142
rect 2142 2141 2148 2142
rect 2318 2146 2324 2147
rect 2318 2142 2319 2146
rect 2323 2142 2324 2146
rect 2318 2141 2324 2142
rect 2494 2146 2500 2147
rect 2494 2142 2495 2146
rect 2499 2142 2500 2146
rect 2494 2141 2500 2142
rect 2678 2146 2684 2147
rect 2678 2142 2679 2146
rect 2683 2142 2684 2146
rect 2678 2141 2684 2142
rect 2862 2146 2868 2147
rect 2862 2142 2863 2146
rect 2867 2142 2868 2146
rect 2862 2141 2868 2142
rect 3038 2146 3044 2147
rect 3038 2142 3039 2146
rect 3043 2142 3044 2146
rect 3038 2141 3044 2142
rect 3214 2146 3220 2147
rect 3214 2142 3215 2146
rect 3219 2142 3220 2146
rect 3214 2141 3220 2142
rect 3390 2146 3396 2147
rect 3390 2142 3391 2146
rect 3395 2142 3396 2146
rect 3390 2141 3396 2142
rect 3566 2146 3572 2147
rect 3566 2142 3567 2146
rect 3571 2142 3572 2146
rect 3566 2141 3572 2142
rect 3742 2146 3748 2147
rect 3742 2142 3743 2146
rect 3747 2142 3748 2146
rect 3742 2141 3748 2142
rect 3894 2146 3900 2147
rect 3894 2142 3895 2146
rect 3899 2142 3900 2146
rect 3894 2141 3900 2142
rect 3990 2141 3996 2142
rect 2070 2137 2071 2141
rect 2075 2137 2076 2141
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 2030 2136 2036 2137
rect 2070 2136 2076 2137
rect 3990 2137 3991 2141
rect 3995 2137 3996 2141
rect 3990 2136 3996 2137
rect 2030 2132 2031 2136
rect 2035 2132 2036 2136
rect 2030 2131 2036 2132
rect 238 2127 244 2128
rect 238 2126 239 2127
rect 201 2124 239 2126
rect 238 2123 239 2124
rect 243 2123 244 2127
rect 450 2127 456 2128
rect 450 2126 451 2127
rect 369 2124 451 2126
rect 238 2122 244 2123
rect 450 2123 451 2124
rect 455 2123 456 2127
rect 450 2122 456 2123
rect 534 2127 540 2128
rect 534 2123 535 2127
rect 539 2123 540 2127
rect 878 2127 884 2128
rect 878 2126 879 2127
rect 753 2124 879 2126
rect 534 2122 540 2123
rect 878 2123 879 2124
rect 883 2123 884 2127
rect 878 2122 884 2123
rect 918 2127 924 2128
rect 918 2123 919 2127
rect 923 2123 924 2127
rect 1255 2127 1261 2128
rect 1255 2126 1256 2127
rect 1137 2124 1256 2126
rect 918 2122 924 2123
rect 1255 2123 1256 2124
rect 1260 2123 1261 2127
rect 1406 2127 1412 2128
rect 1406 2126 1407 2127
rect 1329 2124 1407 2126
rect 1255 2122 1261 2123
rect 1406 2123 1407 2124
rect 1411 2123 1412 2127
rect 1638 2127 1644 2128
rect 1638 2126 1639 2127
rect 1513 2124 1639 2126
rect 1406 2122 1412 2123
rect 1638 2123 1639 2124
rect 1643 2123 1644 2127
rect 1705 2124 1786 2126
rect 1638 2122 1644 2123
rect 150 2117 156 2118
rect 150 2113 151 2117
rect 155 2113 156 2117
rect 150 2112 156 2113
rect 318 2117 324 2118
rect 318 2113 319 2117
rect 323 2113 324 2117
rect 318 2112 324 2113
rect 510 2117 516 2118
rect 510 2113 511 2117
rect 515 2113 516 2117
rect 510 2112 516 2113
rect 702 2117 708 2118
rect 702 2113 703 2117
rect 707 2113 708 2117
rect 702 2112 708 2113
rect 894 2117 900 2118
rect 894 2113 895 2117
rect 899 2113 900 2117
rect 894 2112 900 2113
rect 1086 2117 1092 2118
rect 1086 2113 1087 2117
rect 1091 2113 1092 2117
rect 1086 2112 1092 2113
rect 1278 2117 1284 2118
rect 1278 2113 1279 2117
rect 1283 2113 1284 2117
rect 1278 2112 1284 2113
rect 1462 2117 1468 2118
rect 1462 2113 1463 2117
rect 1467 2113 1468 2117
rect 1462 2112 1468 2113
rect 1654 2117 1660 2118
rect 1654 2113 1655 2117
rect 1659 2113 1660 2117
rect 1654 2112 1660 2113
rect 1784 2114 1786 2124
rect 2070 2124 2076 2125
rect 3990 2124 3996 2125
rect 2070 2120 2071 2124
rect 2075 2120 2076 2124
rect 2686 2123 2692 2124
rect 2686 2122 2687 2123
rect 2070 2119 2076 2120
rect 2620 2120 2687 2122
rect 1846 2117 1852 2118
rect 1784 2112 1842 2114
rect 1846 2113 1847 2117
rect 1851 2113 1852 2117
rect 2214 2115 2220 2116
rect 2214 2114 2215 2115
rect 1846 2112 1852 2113
rect 2193 2112 2215 2114
rect 222 2107 229 2108
rect 222 2103 223 2107
rect 228 2103 229 2107
rect 222 2102 229 2103
rect 238 2107 244 2108
rect 238 2103 239 2107
rect 243 2106 244 2107
rect 391 2107 397 2108
rect 391 2106 392 2107
rect 243 2104 392 2106
rect 243 2103 244 2104
rect 238 2102 244 2103
rect 391 2103 392 2104
rect 396 2103 397 2107
rect 391 2102 397 2103
rect 450 2107 456 2108
rect 450 2103 451 2107
rect 455 2106 456 2107
rect 583 2107 589 2108
rect 583 2106 584 2107
rect 455 2104 584 2106
rect 455 2103 456 2104
rect 450 2102 456 2103
rect 583 2103 584 2104
rect 588 2103 589 2107
rect 583 2102 589 2103
rect 726 2107 732 2108
rect 726 2103 727 2107
rect 731 2106 732 2107
rect 775 2107 781 2108
rect 775 2106 776 2107
rect 731 2104 776 2106
rect 731 2103 732 2104
rect 726 2102 732 2103
rect 775 2103 776 2104
rect 780 2103 781 2107
rect 775 2102 781 2103
rect 878 2107 884 2108
rect 878 2103 879 2107
rect 883 2106 884 2107
rect 967 2107 973 2108
rect 967 2106 968 2107
rect 883 2104 968 2106
rect 883 2103 884 2104
rect 878 2102 884 2103
rect 967 2103 968 2104
rect 972 2103 973 2107
rect 967 2102 973 2103
rect 1114 2107 1120 2108
rect 1114 2103 1115 2107
rect 1119 2106 1120 2107
rect 1159 2107 1165 2108
rect 1159 2106 1160 2107
rect 1119 2104 1160 2106
rect 1119 2103 1120 2104
rect 1114 2102 1120 2103
rect 1159 2103 1160 2104
rect 1164 2103 1165 2107
rect 1159 2102 1165 2103
rect 1255 2107 1261 2108
rect 1255 2103 1256 2107
rect 1260 2106 1261 2107
rect 1351 2107 1357 2108
rect 1351 2106 1352 2107
rect 1260 2104 1352 2106
rect 1260 2103 1261 2104
rect 1255 2102 1261 2103
rect 1351 2103 1352 2104
rect 1356 2103 1357 2107
rect 1351 2102 1357 2103
rect 1534 2107 1541 2108
rect 1534 2103 1535 2107
rect 1540 2103 1541 2107
rect 1534 2102 1541 2103
rect 1638 2107 1644 2108
rect 1638 2103 1639 2107
rect 1643 2106 1644 2107
rect 1727 2107 1733 2108
rect 1727 2106 1728 2107
rect 1643 2104 1728 2106
rect 1643 2103 1644 2104
rect 1638 2102 1644 2103
rect 1727 2103 1728 2104
rect 1732 2103 1733 2107
rect 1727 2102 1733 2103
rect 1738 2107 1744 2108
rect 1738 2103 1739 2107
rect 1743 2106 1744 2107
rect 1831 2107 1837 2108
rect 1831 2106 1832 2107
rect 1743 2104 1832 2106
rect 1743 2103 1744 2104
rect 1738 2102 1744 2103
rect 1831 2103 1832 2104
rect 1836 2103 1837 2107
rect 1840 2106 1842 2112
rect 2214 2111 2215 2112
rect 2219 2111 2220 2115
rect 2620 2114 2622 2120
rect 2686 2119 2687 2120
rect 2691 2119 2692 2123
rect 3990 2120 3991 2124
rect 3995 2120 3996 2124
rect 3990 2119 3996 2120
rect 2686 2118 2692 2119
rect 3110 2115 3116 2116
rect 3110 2114 3111 2115
rect 2545 2112 2622 2114
rect 3089 2112 3111 2114
rect 2214 2110 2220 2111
rect 3110 2111 3111 2112
rect 3115 2111 3116 2115
rect 3718 2115 3724 2116
rect 3718 2114 3719 2115
rect 3617 2112 3719 2114
rect 3110 2110 3116 2111
rect 3718 2111 3719 2112
rect 3723 2111 3724 2115
rect 3966 2115 3972 2116
rect 3966 2114 3967 2115
rect 3945 2112 3967 2114
rect 3718 2110 3724 2111
rect 3966 2111 3967 2112
rect 3971 2111 3972 2115
rect 3966 2110 3972 2111
rect 1919 2107 1925 2108
rect 1919 2106 1920 2107
rect 1840 2104 1920 2106
rect 1831 2102 1837 2103
rect 1919 2103 1920 2104
rect 1924 2103 1925 2107
rect 1919 2102 1925 2103
rect 2142 2105 2148 2106
rect 2142 2101 2143 2105
rect 2147 2101 2148 2105
rect 2142 2100 2148 2101
rect 2318 2105 2324 2106
rect 2318 2101 2319 2105
rect 2323 2101 2324 2105
rect 2318 2100 2324 2101
rect 2494 2105 2500 2106
rect 2494 2101 2495 2105
rect 2499 2101 2500 2105
rect 2494 2100 2500 2101
rect 2678 2105 2684 2106
rect 2678 2101 2679 2105
rect 2683 2101 2684 2105
rect 2678 2100 2684 2101
rect 2862 2105 2868 2106
rect 2862 2101 2863 2105
rect 2867 2101 2868 2105
rect 2862 2100 2868 2101
rect 3038 2105 3044 2106
rect 3038 2101 3039 2105
rect 3043 2101 3044 2105
rect 3038 2100 3044 2101
rect 3214 2105 3220 2106
rect 3214 2101 3215 2105
rect 3219 2101 3220 2105
rect 3214 2100 3220 2101
rect 3390 2105 3396 2106
rect 3390 2101 3391 2105
rect 3395 2101 3396 2105
rect 3390 2100 3396 2101
rect 3566 2105 3572 2106
rect 3566 2101 3567 2105
rect 3571 2101 3572 2105
rect 3566 2100 3572 2101
rect 3742 2105 3748 2106
rect 3742 2101 3743 2105
rect 3747 2101 3748 2105
rect 3742 2100 3748 2101
rect 3894 2105 3900 2106
rect 3894 2101 3895 2105
rect 3899 2101 3900 2105
rect 3894 2100 3900 2101
rect 2215 2095 2221 2096
rect 2215 2091 2216 2095
rect 2220 2094 2221 2095
rect 2303 2095 2309 2096
rect 2303 2094 2304 2095
rect 2220 2092 2304 2094
rect 2220 2091 2221 2092
rect 2215 2090 2221 2091
rect 2303 2091 2304 2092
rect 2308 2091 2309 2095
rect 2303 2090 2309 2091
rect 2390 2095 2397 2096
rect 2390 2091 2391 2095
rect 2396 2091 2397 2095
rect 2390 2090 2397 2091
rect 2567 2095 2573 2096
rect 2567 2091 2568 2095
rect 2572 2094 2573 2095
rect 2663 2095 2669 2096
rect 2663 2094 2664 2095
rect 2572 2092 2664 2094
rect 2572 2091 2573 2092
rect 2567 2090 2573 2091
rect 2663 2091 2664 2092
rect 2668 2091 2669 2095
rect 2663 2090 2669 2091
rect 2751 2095 2757 2096
rect 2751 2091 2752 2095
rect 2756 2094 2757 2095
rect 2847 2095 2853 2096
rect 2847 2094 2848 2095
rect 2756 2092 2848 2094
rect 2756 2091 2757 2092
rect 2751 2090 2757 2091
rect 2847 2091 2848 2092
rect 2852 2091 2853 2095
rect 2847 2090 2853 2091
rect 2926 2095 2932 2096
rect 2926 2091 2927 2095
rect 2931 2094 2932 2095
rect 2935 2095 2941 2096
rect 2935 2094 2936 2095
rect 2931 2092 2936 2094
rect 2931 2091 2932 2092
rect 2926 2090 2932 2091
rect 2935 2091 2936 2092
rect 2940 2091 2941 2095
rect 2935 2090 2941 2091
rect 3111 2095 3117 2096
rect 3111 2091 3112 2095
rect 3116 2094 3117 2095
rect 3199 2095 3205 2096
rect 3199 2094 3200 2095
rect 3116 2092 3200 2094
rect 3116 2091 3117 2092
rect 3111 2090 3117 2091
rect 3199 2091 3200 2092
rect 3204 2091 3205 2095
rect 3199 2090 3205 2091
rect 3287 2095 3293 2096
rect 3287 2091 3288 2095
rect 3292 2094 3293 2095
rect 3375 2095 3381 2096
rect 3375 2094 3376 2095
rect 3292 2092 3376 2094
rect 3292 2091 3293 2092
rect 3287 2090 3293 2091
rect 3375 2091 3376 2092
rect 3380 2091 3381 2095
rect 3375 2090 3381 2091
rect 3463 2095 3469 2096
rect 3463 2091 3464 2095
rect 3468 2094 3469 2095
rect 3478 2095 3484 2096
rect 3478 2094 3479 2095
rect 3468 2092 3479 2094
rect 3468 2091 3469 2092
rect 3463 2090 3469 2091
rect 3478 2091 3479 2092
rect 3483 2091 3484 2095
rect 3478 2090 3484 2091
rect 3639 2095 3645 2096
rect 3639 2091 3640 2095
rect 3644 2094 3645 2095
rect 3727 2095 3733 2096
rect 3727 2094 3728 2095
rect 3644 2092 3728 2094
rect 3644 2091 3645 2092
rect 3639 2090 3645 2091
rect 3727 2091 3728 2092
rect 3732 2091 3733 2095
rect 3727 2090 3733 2091
rect 3814 2095 3821 2096
rect 3814 2091 3815 2095
rect 3820 2091 3821 2095
rect 3814 2090 3821 2091
rect 3958 2095 3964 2096
rect 3958 2091 3959 2095
rect 3963 2094 3964 2095
rect 3967 2095 3973 2096
rect 3967 2094 3968 2095
rect 3963 2092 3968 2094
rect 3963 2091 3964 2092
rect 3958 2090 3964 2091
rect 3967 2091 3968 2092
rect 3972 2091 3973 2095
rect 3967 2090 3973 2091
rect 223 2087 229 2088
rect 223 2083 224 2087
rect 228 2086 229 2087
rect 287 2087 293 2088
rect 287 2086 288 2087
rect 228 2084 288 2086
rect 228 2083 229 2084
rect 223 2082 229 2083
rect 287 2083 288 2084
rect 292 2083 293 2087
rect 287 2082 293 2083
rect 375 2087 381 2088
rect 375 2083 376 2087
rect 380 2086 381 2087
rect 463 2087 469 2088
rect 463 2086 464 2087
rect 380 2084 464 2086
rect 380 2083 381 2084
rect 375 2082 381 2083
rect 463 2083 464 2084
rect 468 2083 469 2087
rect 463 2082 469 2083
rect 534 2087 540 2088
rect 534 2083 535 2087
rect 539 2086 540 2087
rect 551 2087 557 2088
rect 551 2086 552 2087
rect 539 2084 552 2086
rect 539 2083 540 2084
rect 534 2082 540 2083
rect 551 2083 552 2084
rect 556 2083 557 2087
rect 551 2082 557 2083
rect 735 2087 741 2088
rect 735 2083 736 2087
rect 740 2086 741 2087
rect 831 2087 837 2088
rect 831 2086 832 2087
rect 740 2084 832 2086
rect 740 2083 741 2084
rect 735 2082 741 2083
rect 831 2083 832 2084
rect 836 2083 837 2087
rect 831 2082 837 2083
rect 918 2087 925 2088
rect 918 2083 919 2087
rect 924 2083 925 2087
rect 918 2082 925 2083
rect 1111 2087 1117 2088
rect 1111 2083 1112 2087
rect 1116 2086 1117 2087
rect 1223 2087 1229 2088
rect 1223 2086 1224 2087
rect 1116 2084 1224 2086
rect 1116 2083 1117 2084
rect 1111 2082 1117 2083
rect 1223 2083 1224 2084
rect 1228 2083 1229 2087
rect 1223 2082 1229 2083
rect 1311 2087 1317 2088
rect 1311 2083 1312 2087
rect 1316 2086 1317 2087
rect 1431 2087 1437 2088
rect 1431 2086 1432 2087
rect 1316 2084 1432 2086
rect 1316 2083 1317 2084
rect 1311 2082 1317 2083
rect 1431 2083 1432 2084
rect 1436 2083 1437 2087
rect 1431 2082 1437 2083
rect 1454 2087 1460 2088
rect 1454 2083 1455 2087
rect 1459 2086 1460 2087
rect 1519 2087 1525 2088
rect 1519 2086 1520 2087
rect 1459 2084 1520 2086
rect 1459 2083 1460 2084
rect 1454 2082 1460 2083
rect 1519 2083 1520 2084
rect 1524 2083 1525 2087
rect 1519 2082 1525 2083
rect 1735 2087 1744 2088
rect 1735 2083 1736 2087
rect 1743 2083 1744 2087
rect 1951 2087 1957 2088
rect 1951 2086 1952 2087
rect 1735 2082 1744 2083
rect 1804 2084 1952 2086
rect 150 2079 156 2080
rect 150 2075 151 2079
rect 155 2075 156 2079
rect 150 2074 156 2075
rect 302 2079 308 2080
rect 302 2075 303 2079
rect 307 2075 308 2079
rect 302 2074 308 2075
rect 478 2079 484 2080
rect 478 2075 479 2079
rect 483 2075 484 2079
rect 478 2074 484 2075
rect 662 2079 668 2080
rect 662 2075 663 2079
rect 667 2075 668 2079
rect 662 2074 668 2075
rect 846 2079 852 2080
rect 846 2075 847 2079
rect 851 2075 852 2079
rect 846 2074 852 2075
rect 1038 2079 1044 2080
rect 1038 2075 1039 2079
rect 1043 2075 1044 2079
rect 1038 2074 1044 2075
rect 1238 2079 1244 2080
rect 1238 2075 1239 2079
rect 1243 2075 1244 2079
rect 1238 2074 1244 2075
rect 1446 2079 1452 2080
rect 1446 2075 1447 2079
rect 1451 2075 1452 2079
rect 1446 2074 1452 2075
rect 1662 2079 1668 2080
rect 1662 2075 1663 2079
rect 1667 2075 1668 2079
rect 1662 2074 1668 2075
rect 222 2071 228 2072
rect 222 2070 223 2071
rect 201 2068 223 2070
rect 222 2067 223 2068
rect 227 2067 228 2071
rect 726 2071 732 2072
rect 726 2070 727 2071
rect 713 2068 727 2070
rect 222 2066 228 2067
rect 726 2067 727 2068
rect 731 2067 732 2071
rect 1114 2071 1120 2072
rect 1114 2070 1115 2071
rect 1089 2068 1115 2070
rect 726 2066 732 2067
rect 1114 2067 1115 2068
rect 1119 2067 1120 2071
rect 1804 2070 1806 2084
rect 1951 2083 1952 2084
rect 1956 2083 1957 2087
rect 1951 2082 1957 2083
rect 1878 2079 1884 2080
rect 1878 2075 1879 2079
rect 1883 2075 1884 2079
rect 1878 2074 1884 2075
rect 3246 2079 3252 2080
rect 3246 2075 3247 2079
rect 3251 2078 3252 2079
rect 3251 2076 3418 2078
rect 3251 2075 3252 2076
rect 3246 2074 3252 2075
rect 2006 2071 2012 2072
rect 2006 2070 2007 2071
rect 1713 2068 1806 2070
rect 1929 2068 2007 2070
rect 1114 2066 1120 2067
rect 2006 2067 2007 2068
rect 2011 2067 2012 2071
rect 2006 2066 2012 2067
rect 2214 2071 2220 2072
rect 2214 2067 2215 2071
rect 2219 2070 2220 2071
rect 2279 2071 2285 2072
rect 2279 2070 2280 2071
rect 2219 2068 2280 2070
rect 2219 2067 2220 2068
rect 2214 2066 2220 2067
rect 2279 2067 2280 2068
rect 2284 2067 2285 2071
rect 2463 2071 2469 2072
rect 2463 2070 2464 2071
rect 2279 2066 2285 2067
rect 2332 2068 2464 2070
rect 2206 2063 2212 2064
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 2030 2060 2036 2061
rect 2030 2056 2031 2060
rect 2035 2056 2036 2060
rect 2206 2059 2207 2063
rect 2211 2059 2212 2063
rect 2206 2058 2212 2059
rect 2030 2055 2036 2056
rect 2332 2054 2334 2068
rect 2463 2067 2464 2068
rect 2468 2067 2469 2071
rect 2463 2066 2469 2067
rect 2646 2071 2653 2072
rect 2646 2067 2647 2071
rect 2652 2067 2653 2071
rect 2831 2071 2837 2072
rect 2831 2070 2832 2071
rect 2646 2066 2653 2067
rect 2700 2068 2832 2070
rect 2390 2063 2396 2064
rect 2390 2059 2391 2063
rect 2395 2059 2396 2063
rect 2390 2058 2396 2059
rect 2574 2063 2580 2064
rect 2574 2059 2575 2063
rect 2579 2059 2580 2063
rect 2574 2058 2580 2059
rect 2700 2054 2702 2068
rect 2831 2067 2832 2068
rect 2836 2067 2837 2071
rect 3007 2071 3013 2072
rect 3007 2070 3008 2071
rect 2831 2066 2837 2067
rect 2839 2068 3008 2070
rect 2758 2063 2764 2064
rect 2758 2059 2759 2063
rect 2763 2059 2764 2063
rect 2758 2058 2764 2059
rect 2839 2054 2841 2068
rect 3007 2067 3008 2068
rect 3012 2067 3013 2071
rect 3007 2066 3013 2067
rect 3110 2071 3116 2072
rect 3110 2067 3111 2071
rect 3115 2070 3116 2071
rect 3175 2071 3181 2072
rect 3175 2070 3176 2071
rect 3115 2068 3176 2070
rect 3115 2067 3116 2068
rect 3110 2066 3116 2067
rect 3175 2067 3176 2068
rect 3180 2067 3181 2071
rect 3175 2066 3181 2067
rect 3335 2071 3341 2072
rect 3335 2067 3336 2071
rect 3340 2070 3341 2071
rect 3407 2071 3413 2072
rect 3407 2070 3408 2071
rect 3340 2068 3408 2070
rect 3340 2067 3341 2068
rect 3335 2066 3341 2067
rect 3407 2067 3408 2068
rect 3412 2067 3413 2071
rect 3416 2070 3418 2076
rect 3495 2071 3501 2072
rect 3495 2070 3496 2071
rect 3416 2068 3496 2070
rect 3407 2066 3413 2067
rect 3495 2067 3496 2068
rect 3500 2067 3501 2071
rect 3495 2066 3501 2067
rect 3638 2071 3644 2072
rect 3638 2067 3639 2071
rect 3643 2070 3644 2071
rect 3655 2071 3661 2072
rect 3655 2070 3656 2071
rect 3643 2068 3656 2070
rect 3643 2067 3644 2068
rect 3638 2066 3644 2067
rect 3655 2067 3656 2068
rect 3660 2067 3661 2071
rect 3823 2071 3829 2072
rect 3823 2070 3824 2071
rect 3655 2066 3661 2067
rect 3679 2068 3824 2070
rect 2934 2063 2940 2064
rect 2934 2059 2935 2063
rect 2939 2059 2940 2063
rect 2934 2058 2940 2059
rect 3102 2063 3108 2064
rect 3102 2059 3103 2063
rect 3107 2059 3108 2063
rect 3102 2058 3108 2059
rect 3262 2063 3268 2064
rect 3262 2059 3263 2063
rect 3267 2059 3268 2063
rect 3262 2058 3268 2059
rect 3422 2063 3428 2064
rect 3422 2059 3423 2063
rect 3427 2059 3428 2063
rect 3422 2058 3428 2059
rect 3582 2063 3588 2064
rect 3582 2059 3583 2063
rect 3587 2059 3588 2063
rect 3582 2058 3588 2059
rect 2257 2052 2334 2054
rect 2625 2052 2702 2054
rect 2809 2052 2841 2054
rect 2926 2055 2932 2056
rect 2382 2051 2388 2052
rect 2382 2047 2383 2051
rect 2387 2047 2388 2051
rect 2926 2051 2927 2055
rect 2931 2051 2932 2055
rect 3246 2055 3252 2056
rect 3246 2054 3247 2055
rect 3153 2052 3247 2054
rect 2926 2050 2932 2051
rect 3246 2051 3247 2052
rect 3251 2051 3252 2055
rect 3679 2054 3681 2068
rect 3823 2067 3824 2068
rect 3828 2067 3829 2071
rect 3823 2066 3829 2067
rect 3966 2071 3973 2072
rect 3966 2067 3967 2071
rect 3972 2067 3973 2071
rect 3966 2066 3973 2067
rect 3750 2063 3756 2064
rect 3750 2059 3751 2063
rect 3755 2059 3756 2063
rect 3750 2058 3756 2059
rect 3894 2063 3900 2064
rect 3894 2059 3895 2063
rect 3899 2059 3900 2063
rect 3894 2058 3900 2059
rect 3814 2055 3820 2056
rect 3814 2054 3815 2055
rect 3633 2052 3681 2054
rect 3801 2052 3815 2054
rect 3246 2050 3252 2051
rect 3254 2051 3260 2052
rect 2382 2046 2388 2047
rect 3254 2047 3255 2051
rect 3259 2047 3260 2051
rect 3814 2051 3815 2052
rect 3819 2051 3820 2055
rect 3958 2055 3964 2056
rect 3958 2054 3959 2055
rect 3945 2052 3959 2054
rect 3814 2050 3820 2051
rect 3958 2051 3959 2052
rect 3963 2051 3964 2055
rect 3958 2050 3964 2051
rect 3254 2046 3260 2047
rect 2070 2044 2076 2045
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 2030 2043 2036 2044
rect 2030 2039 2031 2043
rect 2035 2039 2036 2043
rect 2070 2040 2071 2044
rect 2075 2040 2076 2044
rect 2070 2039 2076 2040
rect 3990 2044 3996 2045
rect 3990 2040 3991 2044
rect 3995 2040 3996 2044
rect 3990 2039 3996 2040
rect 110 2038 116 2039
rect 150 2038 156 2039
rect 150 2034 151 2038
rect 155 2034 156 2038
rect 150 2033 156 2034
rect 302 2038 308 2039
rect 302 2034 303 2038
rect 307 2034 308 2038
rect 302 2033 308 2034
rect 478 2038 484 2039
rect 478 2034 479 2038
rect 483 2034 484 2038
rect 478 2033 484 2034
rect 662 2038 668 2039
rect 662 2034 663 2038
rect 667 2034 668 2038
rect 662 2033 668 2034
rect 846 2038 852 2039
rect 846 2034 847 2038
rect 851 2034 852 2038
rect 846 2033 852 2034
rect 1038 2038 1044 2039
rect 1038 2034 1039 2038
rect 1043 2034 1044 2038
rect 1038 2033 1044 2034
rect 1238 2038 1244 2039
rect 1238 2034 1239 2038
rect 1243 2034 1244 2038
rect 1238 2033 1244 2034
rect 1446 2038 1452 2039
rect 1446 2034 1447 2038
rect 1451 2034 1452 2038
rect 1446 2033 1452 2034
rect 1662 2038 1668 2039
rect 1662 2034 1663 2038
rect 1667 2034 1668 2038
rect 1662 2033 1668 2034
rect 1878 2038 1884 2039
rect 2030 2038 2036 2039
rect 1878 2034 1879 2038
rect 1883 2034 1884 2038
rect 1878 2033 1884 2034
rect 2070 2027 2076 2028
rect 2070 2023 2071 2027
rect 2075 2023 2076 2027
rect 3990 2027 3996 2028
rect 3990 2023 3991 2027
rect 3995 2023 3996 2027
rect 2070 2022 2076 2023
rect 2206 2022 2212 2023
rect 2206 2018 2207 2022
rect 2211 2018 2212 2022
rect 2206 2017 2212 2018
rect 2390 2022 2396 2023
rect 2390 2018 2391 2022
rect 2395 2018 2396 2022
rect 2390 2017 2396 2018
rect 2574 2022 2580 2023
rect 2574 2018 2575 2022
rect 2579 2018 2580 2022
rect 2574 2017 2580 2018
rect 2758 2022 2764 2023
rect 2758 2018 2759 2022
rect 2763 2018 2764 2022
rect 2758 2017 2764 2018
rect 2934 2022 2940 2023
rect 2934 2018 2935 2022
rect 2939 2018 2940 2022
rect 2934 2017 2940 2018
rect 3102 2022 3108 2023
rect 3102 2018 3103 2022
rect 3107 2018 3108 2022
rect 3102 2017 3108 2018
rect 3262 2022 3268 2023
rect 3262 2018 3263 2022
rect 3267 2018 3268 2022
rect 3262 2017 3268 2018
rect 3422 2022 3428 2023
rect 3422 2018 3423 2022
rect 3427 2018 3428 2022
rect 3422 2017 3428 2018
rect 3582 2022 3588 2023
rect 3582 2018 3583 2022
rect 3587 2018 3588 2022
rect 3582 2017 3588 2018
rect 3750 2022 3756 2023
rect 3750 2018 3751 2022
rect 3755 2018 3756 2022
rect 3750 2017 3756 2018
rect 3894 2022 3900 2023
rect 3990 2022 3996 2023
rect 3894 2018 3895 2022
rect 3899 2018 3900 2022
rect 3894 2017 3900 2018
rect 150 1998 156 1999
rect 150 1994 151 1998
rect 155 1994 156 1998
rect 110 1993 116 1994
rect 150 1993 156 1994
rect 302 1998 308 1999
rect 302 1994 303 1998
rect 307 1994 308 1998
rect 302 1993 308 1994
rect 486 1998 492 1999
rect 486 1994 487 1998
rect 491 1994 492 1998
rect 486 1993 492 1994
rect 686 1998 692 1999
rect 686 1994 687 1998
rect 691 1994 692 1998
rect 686 1993 692 1994
rect 894 1998 900 1999
rect 894 1994 895 1998
rect 899 1994 900 1998
rect 894 1993 900 1994
rect 1102 1998 1108 1999
rect 1102 1994 1103 1998
rect 1107 1994 1108 1998
rect 1102 1993 1108 1994
rect 1310 1998 1316 1999
rect 1310 1994 1311 1998
rect 1315 1994 1316 1998
rect 1310 1993 1316 1994
rect 1526 1998 1532 1999
rect 1526 1994 1527 1998
rect 1531 1994 1532 1998
rect 1526 1993 1532 1994
rect 1742 1998 1748 1999
rect 1742 1994 1743 1998
rect 1747 1994 1748 1998
rect 1742 1993 1748 1994
rect 1934 1998 1940 1999
rect 1934 1994 1935 1998
rect 1939 1994 1940 1998
rect 1934 1993 1940 1994
rect 2030 1993 2036 1994
rect 110 1989 111 1993
rect 115 1989 116 1993
rect 110 1988 116 1989
rect 2030 1989 2031 1993
rect 2035 1989 2036 1993
rect 2030 1988 2036 1989
rect 2278 1978 2284 1979
rect 110 1976 116 1977
rect 110 1972 111 1976
rect 115 1972 116 1976
rect 110 1971 116 1972
rect 2030 1976 2036 1977
rect 2030 1972 2031 1976
rect 2035 1972 2036 1976
rect 2278 1974 2279 1978
rect 2283 1974 2284 1978
rect 2030 1971 2036 1972
rect 2070 1973 2076 1974
rect 2278 1973 2284 1974
rect 2462 1978 2468 1979
rect 2462 1974 2463 1978
rect 2467 1974 2468 1978
rect 2462 1973 2468 1974
rect 2638 1978 2644 1979
rect 2638 1974 2639 1978
rect 2643 1974 2644 1978
rect 2638 1973 2644 1974
rect 2814 1978 2820 1979
rect 2814 1974 2815 1978
rect 2819 1974 2820 1978
rect 2814 1973 2820 1974
rect 2982 1978 2988 1979
rect 2982 1974 2983 1978
rect 2987 1974 2988 1978
rect 2982 1973 2988 1974
rect 3150 1978 3156 1979
rect 3150 1974 3151 1978
rect 3155 1974 3156 1978
rect 3150 1973 3156 1974
rect 3310 1978 3316 1979
rect 3310 1974 3311 1978
rect 3315 1974 3316 1978
rect 3310 1973 3316 1974
rect 3462 1978 3468 1979
rect 3462 1974 3463 1978
rect 3467 1974 3468 1978
rect 3462 1973 3468 1974
rect 3614 1978 3620 1979
rect 3614 1974 3615 1978
rect 3619 1974 3620 1978
rect 3614 1973 3620 1974
rect 3766 1978 3772 1979
rect 3766 1974 3767 1978
rect 3771 1974 3772 1978
rect 3766 1973 3772 1974
rect 3894 1978 3900 1979
rect 3894 1974 3895 1978
rect 3899 1974 3900 1978
rect 3894 1973 3900 1974
rect 3990 1973 3996 1974
rect 2070 1969 2071 1973
rect 2075 1969 2076 1973
rect 2070 1968 2076 1969
rect 3990 1969 3991 1973
rect 3995 1969 3996 1973
rect 3990 1968 3996 1969
rect 231 1967 237 1968
rect 231 1966 232 1967
rect 201 1964 232 1966
rect 231 1963 232 1964
rect 236 1963 237 1967
rect 438 1967 444 1968
rect 438 1966 439 1967
rect 353 1964 439 1966
rect 231 1962 237 1963
rect 438 1963 439 1964
rect 443 1963 444 1967
rect 438 1962 444 1963
rect 478 1967 484 1968
rect 478 1963 479 1967
rect 483 1963 484 1967
rect 878 1967 884 1968
rect 878 1966 879 1967
rect 737 1964 879 1966
rect 478 1962 484 1963
rect 878 1963 879 1964
rect 883 1963 884 1967
rect 878 1962 884 1963
rect 918 1967 924 1968
rect 918 1963 919 1967
rect 923 1963 924 1967
rect 1294 1967 1300 1968
rect 1294 1966 1295 1967
rect 1153 1964 1295 1966
rect 918 1962 924 1963
rect 1294 1963 1295 1964
rect 1299 1963 1300 1967
rect 1454 1967 1460 1968
rect 1454 1966 1455 1967
rect 1361 1964 1455 1966
rect 1294 1962 1300 1963
rect 1454 1963 1455 1964
rect 1459 1963 1460 1967
rect 1670 1967 1676 1968
rect 1670 1966 1671 1967
rect 1577 1964 1671 1966
rect 1454 1962 1460 1963
rect 1670 1963 1671 1964
rect 1675 1963 1676 1967
rect 1670 1962 1676 1963
rect 150 1957 156 1958
rect 150 1953 151 1957
rect 155 1953 156 1957
rect 150 1952 156 1953
rect 302 1957 308 1958
rect 302 1953 303 1957
rect 307 1953 308 1957
rect 302 1952 308 1953
rect 486 1957 492 1958
rect 486 1953 487 1957
rect 491 1953 492 1957
rect 486 1952 492 1953
rect 686 1957 692 1958
rect 686 1953 687 1957
rect 691 1953 692 1957
rect 686 1952 692 1953
rect 894 1957 900 1958
rect 894 1953 895 1957
rect 899 1953 900 1957
rect 894 1952 900 1953
rect 1102 1957 1108 1958
rect 1102 1953 1103 1957
rect 1107 1953 1108 1957
rect 1102 1952 1108 1953
rect 1310 1957 1316 1958
rect 1310 1953 1311 1957
rect 1315 1953 1316 1957
rect 1310 1952 1316 1953
rect 1526 1957 1532 1958
rect 1526 1953 1527 1957
rect 1531 1953 1532 1957
rect 1526 1952 1532 1953
rect 1742 1957 1748 1958
rect 1742 1953 1743 1957
rect 1747 1953 1748 1957
rect 1742 1952 1748 1953
rect 1934 1957 1940 1958
rect 1934 1953 1935 1957
rect 1939 1953 1940 1957
rect 1934 1952 1940 1953
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2070 1951 2076 1952
rect 3990 1956 3996 1957
rect 3990 1952 3991 1956
rect 3995 1952 3996 1956
rect 3990 1951 3996 1952
rect 222 1947 229 1948
rect 222 1943 223 1947
rect 228 1943 229 1947
rect 222 1942 229 1943
rect 231 1947 237 1948
rect 231 1943 232 1947
rect 236 1946 237 1947
rect 375 1947 381 1948
rect 375 1946 376 1947
rect 236 1944 376 1946
rect 236 1943 237 1944
rect 231 1942 237 1943
rect 375 1943 376 1944
rect 380 1943 381 1947
rect 375 1942 381 1943
rect 438 1947 444 1948
rect 438 1943 439 1947
rect 443 1946 444 1947
rect 559 1947 565 1948
rect 559 1946 560 1947
rect 443 1944 560 1946
rect 443 1943 444 1944
rect 438 1942 444 1943
rect 559 1943 560 1944
rect 564 1943 565 1947
rect 559 1942 565 1943
rect 742 1947 748 1948
rect 742 1943 743 1947
rect 747 1946 748 1947
rect 759 1947 765 1948
rect 759 1946 760 1947
rect 747 1944 760 1946
rect 747 1943 748 1944
rect 742 1942 748 1943
rect 759 1943 760 1944
rect 764 1943 765 1947
rect 759 1942 765 1943
rect 878 1947 884 1948
rect 878 1943 879 1947
rect 883 1946 884 1947
rect 967 1947 973 1948
rect 967 1946 968 1947
rect 883 1944 968 1946
rect 883 1943 884 1944
rect 878 1942 884 1943
rect 967 1943 968 1944
rect 972 1943 973 1947
rect 1175 1947 1181 1948
rect 1175 1946 1176 1947
rect 967 1942 973 1943
rect 1159 1944 1176 1946
rect 966 1939 972 1940
rect 966 1935 967 1939
rect 971 1938 972 1939
rect 1159 1938 1161 1944
rect 1175 1943 1176 1944
rect 1180 1943 1181 1947
rect 1175 1942 1181 1943
rect 1294 1947 1300 1948
rect 1294 1943 1295 1947
rect 1299 1946 1300 1947
rect 1383 1947 1389 1948
rect 1383 1946 1384 1947
rect 1299 1944 1384 1946
rect 1299 1943 1300 1944
rect 1294 1942 1300 1943
rect 1383 1943 1384 1944
rect 1388 1943 1389 1947
rect 1383 1942 1389 1943
rect 1599 1947 1605 1948
rect 1599 1943 1600 1947
rect 1604 1946 1605 1947
rect 1727 1947 1733 1948
rect 1727 1946 1728 1947
rect 1604 1944 1728 1946
rect 1604 1943 1605 1944
rect 1599 1942 1605 1943
rect 1727 1943 1728 1944
rect 1732 1943 1733 1947
rect 1727 1942 1733 1943
rect 1815 1947 1821 1948
rect 1815 1943 1816 1947
rect 1820 1946 1821 1947
rect 1919 1947 1925 1948
rect 1919 1946 1920 1947
rect 1820 1944 1920 1946
rect 1820 1943 1821 1944
rect 1815 1942 1821 1943
rect 1919 1943 1920 1944
rect 1924 1943 1925 1947
rect 1919 1942 1925 1943
rect 2006 1947 2013 1948
rect 2006 1943 2007 1947
rect 2012 1943 2013 1947
rect 2446 1947 2452 1948
rect 2446 1946 2447 1947
rect 2329 1944 2447 1946
rect 2006 1942 2013 1943
rect 2446 1943 2447 1944
rect 2451 1943 2452 1947
rect 2590 1947 2596 1948
rect 2590 1946 2591 1947
rect 2513 1944 2591 1946
rect 2446 1942 2452 1943
rect 2590 1943 2591 1944
rect 2595 1943 2596 1947
rect 2590 1942 2596 1943
rect 2646 1947 2652 1948
rect 2646 1943 2647 1947
rect 2651 1943 2652 1947
rect 3294 1947 3300 1948
rect 3294 1946 3295 1947
rect 3201 1944 3295 1946
rect 2646 1942 2652 1943
rect 3294 1943 3295 1944
rect 3299 1943 3300 1947
rect 3446 1947 3452 1948
rect 3446 1946 3447 1947
rect 3361 1944 3447 1946
rect 3294 1942 3300 1943
rect 3446 1943 3447 1944
rect 3451 1943 3452 1947
rect 3446 1942 3452 1943
rect 3638 1947 3644 1948
rect 3638 1943 3639 1947
rect 3643 1943 3644 1947
rect 3966 1947 3972 1948
rect 3966 1946 3967 1947
rect 3945 1944 3967 1946
rect 3638 1942 3644 1943
rect 3966 1943 3967 1944
rect 3971 1943 3972 1947
rect 3966 1942 3972 1943
rect 971 1936 1161 1938
rect 2278 1937 2284 1938
rect 971 1935 972 1936
rect 966 1934 972 1935
rect 2278 1933 2279 1937
rect 2283 1933 2284 1937
rect 2278 1932 2284 1933
rect 2462 1937 2468 1938
rect 2462 1933 2463 1937
rect 2467 1933 2468 1937
rect 2462 1932 2468 1933
rect 2638 1937 2644 1938
rect 2638 1933 2639 1937
rect 2643 1933 2644 1937
rect 2638 1932 2644 1933
rect 2814 1937 2820 1938
rect 2814 1933 2815 1937
rect 2819 1933 2820 1937
rect 2814 1932 2820 1933
rect 2982 1937 2988 1938
rect 2982 1933 2983 1937
rect 2987 1933 2988 1937
rect 2982 1932 2988 1933
rect 3150 1937 3156 1938
rect 3150 1933 3151 1937
rect 3155 1933 3156 1937
rect 3150 1932 3156 1933
rect 3310 1937 3316 1938
rect 3310 1933 3311 1937
rect 3315 1933 3316 1937
rect 3310 1932 3316 1933
rect 3462 1937 3468 1938
rect 3462 1933 3463 1937
rect 3467 1933 3468 1937
rect 3462 1932 3468 1933
rect 3614 1937 3620 1938
rect 3614 1933 3615 1937
rect 3619 1933 3620 1937
rect 3766 1937 3772 1938
rect 3751 1935 3757 1936
rect 3751 1934 3752 1935
rect 3614 1932 3620 1933
rect 3679 1932 3752 1934
rect 3679 1930 3681 1932
rect 3751 1931 3752 1932
rect 3756 1931 3757 1935
rect 3766 1933 3767 1937
rect 3771 1933 3772 1937
rect 3766 1932 3772 1933
rect 3894 1937 3900 1938
rect 3894 1933 3895 1937
rect 3899 1933 3900 1937
rect 3894 1932 3900 1933
rect 3751 1930 3757 1931
rect 3608 1928 3681 1930
rect 2351 1927 2357 1928
rect 223 1923 229 1924
rect 223 1919 224 1923
rect 228 1922 229 1923
rect 255 1923 261 1924
rect 255 1922 256 1923
rect 228 1920 256 1922
rect 228 1919 229 1920
rect 223 1918 229 1919
rect 255 1919 256 1920
rect 260 1919 261 1923
rect 255 1918 261 1919
rect 343 1923 349 1924
rect 343 1919 344 1923
rect 348 1922 349 1923
rect 391 1923 397 1924
rect 391 1922 392 1923
rect 348 1920 392 1922
rect 348 1919 349 1920
rect 343 1918 349 1919
rect 391 1919 392 1920
rect 396 1919 397 1923
rect 391 1918 397 1919
rect 478 1923 485 1924
rect 478 1919 479 1923
rect 484 1919 485 1923
rect 478 1918 485 1919
rect 614 1923 621 1924
rect 614 1919 615 1923
rect 620 1919 621 1923
rect 751 1923 757 1924
rect 751 1922 752 1923
rect 614 1918 621 1919
rect 644 1920 752 1922
rect 150 1915 156 1916
rect 150 1911 151 1915
rect 155 1911 156 1915
rect 150 1910 156 1911
rect 270 1915 276 1916
rect 270 1911 271 1915
rect 275 1911 276 1915
rect 270 1910 276 1911
rect 406 1915 412 1916
rect 406 1911 407 1915
rect 411 1911 412 1915
rect 406 1910 412 1911
rect 542 1915 548 1916
rect 542 1911 543 1915
rect 547 1911 548 1915
rect 542 1910 548 1911
rect 222 1907 228 1908
rect 222 1906 223 1907
rect 201 1904 223 1906
rect 222 1903 223 1904
rect 227 1903 228 1907
rect 644 1906 646 1920
rect 751 1919 752 1920
rect 756 1919 757 1923
rect 751 1918 757 1919
rect 895 1923 901 1924
rect 895 1919 896 1923
rect 900 1922 901 1923
rect 967 1923 973 1924
rect 967 1922 968 1923
rect 900 1920 968 1922
rect 900 1919 901 1920
rect 895 1918 901 1919
rect 967 1919 968 1920
rect 972 1919 973 1923
rect 967 1918 973 1919
rect 1055 1923 1061 1924
rect 1055 1919 1056 1923
rect 1060 1922 1061 1923
rect 1143 1923 1149 1924
rect 1143 1922 1144 1923
rect 1060 1920 1144 1922
rect 1060 1919 1061 1920
rect 1055 1918 1061 1919
rect 1143 1919 1144 1920
rect 1148 1919 1149 1923
rect 1143 1918 1149 1919
rect 1231 1923 1237 1924
rect 1231 1919 1232 1923
rect 1236 1922 1237 1923
rect 1327 1923 1333 1924
rect 1327 1922 1328 1923
rect 1236 1920 1328 1922
rect 1236 1919 1237 1920
rect 1231 1918 1237 1919
rect 1327 1919 1328 1920
rect 1332 1919 1333 1923
rect 1327 1918 1333 1919
rect 1415 1923 1421 1924
rect 1415 1919 1416 1923
rect 1420 1922 1421 1923
rect 1527 1923 1533 1924
rect 1527 1922 1528 1923
rect 1420 1920 1528 1922
rect 1420 1919 1421 1920
rect 1415 1918 1421 1919
rect 1527 1919 1528 1920
rect 1532 1919 1533 1923
rect 1527 1918 1533 1919
rect 1550 1923 1556 1924
rect 1550 1919 1551 1923
rect 1555 1922 1556 1923
rect 1615 1923 1621 1924
rect 1615 1922 1616 1923
rect 1555 1920 1616 1922
rect 1555 1919 1556 1920
rect 1550 1918 1556 1919
rect 1615 1919 1616 1920
rect 1620 1919 1621 1923
rect 1615 1918 1621 1919
rect 1670 1923 1676 1924
rect 1670 1919 1671 1923
rect 1675 1922 1676 1923
rect 1823 1923 1829 1924
rect 1823 1922 1824 1923
rect 1675 1920 1824 1922
rect 1675 1919 1676 1920
rect 1670 1918 1676 1919
rect 1823 1919 1824 1920
rect 1828 1919 1829 1923
rect 2007 1923 2013 1924
rect 2007 1922 2008 1923
rect 1823 1918 1829 1919
rect 1872 1920 2008 1922
rect 678 1915 684 1916
rect 678 1911 679 1915
rect 683 1911 684 1915
rect 678 1910 684 1911
rect 822 1915 828 1916
rect 822 1911 823 1915
rect 827 1911 828 1915
rect 822 1910 828 1911
rect 982 1915 988 1916
rect 982 1911 983 1915
rect 987 1911 988 1915
rect 982 1910 988 1911
rect 1158 1915 1164 1916
rect 1158 1911 1159 1915
rect 1163 1911 1164 1915
rect 1158 1910 1164 1911
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1342 1910 1348 1911
rect 1542 1915 1548 1916
rect 1542 1911 1543 1915
rect 1547 1911 1548 1915
rect 1542 1910 1548 1911
rect 1750 1915 1756 1916
rect 1750 1911 1751 1915
rect 1755 1911 1756 1915
rect 1750 1910 1756 1911
rect 742 1907 748 1908
rect 742 1906 743 1907
rect 593 1904 646 1906
rect 729 1904 743 1906
rect 222 1902 228 1903
rect 742 1903 743 1904
rect 747 1903 748 1907
rect 966 1907 972 1908
rect 966 1906 967 1907
rect 873 1904 967 1906
rect 742 1902 748 1903
rect 966 1903 967 1904
rect 971 1903 972 1907
rect 1872 1906 1874 1920
rect 2007 1919 2008 1920
rect 2012 1919 2013 1923
rect 2351 1923 2352 1927
rect 2356 1926 2357 1927
rect 2382 1927 2388 1928
rect 2382 1926 2383 1927
rect 2356 1924 2383 1926
rect 2356 1923 2357 1924
rect 2351 1922 2357 1923
rect 2382 1923 2383 1924
rect 2387 1923 2388 1927
rect 2382 1922 2388 1923
rect 2446 1927 2452 1928
rect 2446 1923 2447 1927
rect 2451 1926 2452 1927
rect 2535 1927 2541 1928
rect 2535 1926 2536 1927
rect 2451 1924 2536 1926
rect 2451 1923 2452 1924
rect 2446 1922 2452 1923
rect 2535 1923 2536 1924
rect 2540 1923 2541 1927
rect 2535 1922 2541 1923
rect 2711 1927 2717 1928
rect 2711 1923 2712 1927
rect 2716 1926 2717 1927
rect 2799 1927 2805 1928
rect 2799 1926 2800 1927
rect 2716 1924 2800 1926
rect 2716 1923 2717 1924
rect 2711 1922 2717 1923
rect 2799 1923 2800 1924
rect 2804 1923 2805 1927
rect 2799 1922 2805 1923
rect 2887 1927 2893 1928
rect 2887 1923 2888 1927
rect 2892 1926 2893 1927
rect 2967 1927 2973 1928
rect 2967 1926 2968 1927
rect 2892 1924 2968 1926
rect 2892 1923 2893 1924
rect 2887 1922 2893 1923
rect 2967 1923 2968 1924
rect 2972 1923 2973 1927
rect 2967 1922 2973 1923
rect 2975 1927 2981 1928
rect 2975 1923 2976 1927
rect 2980 1926 2981 1927
rect 3055 1927 3061 1928
rect 3055 1926 3056 1927
rect 2980 1924 3056 1926
rect 2980 1923 2981 1924
rect 2975 1922 2981 1923
rect 3055 1923 3056 1924
rect 3060 1923 3061 1927
rect 3055 1922 3061 1923
rect 3223 1927 3229 1928
rect 3223 1923 3224 1927
rect 3228 1926 3229 1927
rect 3254 1927 3260 1928
rect 3254 1926 3255 1927
rect 3228 1924 3255 1926
rect 3228 1923 3229 1924
rect 3223 1922 3229 1923
rect 3254 1923 3255 1924
rect 3259 1923 3260 1927
rect 3254 1922 3260 1923
rect 3294 1927 3300 1928
rect 3294 1923 3295 1927
rect 3299 1926 3300 1927
rect 3383 1927 3389 1928
rect 3383 1926 3384 1927
rect 3299 1924 3384 1926
rect 3299 1923 3300 1924
rect 3294 1922 3300 1923
rect 3383 1923 3384 1924
rect 3388 1923 3389 1927
rect 3383 1922 3389 1923
rect 3391 1927 3397 1928
rect 3391 1923 3392 1927
rect 3396 1926 3397 1927
rect 3447 1927 3453 1928
rect 3447 1926 3448 1927
rect 3396 1924 3448 1926
rect 3396 1923 3397 1924
rect 3391 1922 3397 1923
rect 3447 1923 3448 1924
rect 3452 1923 3453 1927
rect 3447 1922 3453 1923
rect 3535 1927 3541 1928
rect 3535 1923 3536 1927
rect 3540 1926 3541 1927
rect 3608 1926 3610 1928
rect 3687 1927 3693 1928
rect 3687 1926 3688 1927
rect 3540 1924 3610 1926
rect 3679 1924 3688 1926
rect 3540 1923 3541 1924
rect 3535 1922 3541 1923
rect 2007 1918 2013 1919
rect 3446 1919 3452 1920
rect 1934 1915 1940 1916
rect 1934 1911 1935 1915
rect 1939 1911 1940 1915
rect 1934 1910 1940 1911
rect 2590 1915 2596 1916
rect 2590 1911 2591 1915
rect 2595 1914 2596 1915
rect 3446 1915 3447 1919
rect 3451 1918 3452 1919
rect 3679 1918 3681 1924
rect 3687 1923 3688 1924
rect 3692 1923 3693 1927
rect 3687 1922 3693 1923
rect 3774 1927 3780 1928
rect 3774 1923 3775 1927
rect 3779 1926 3780 1927
rect 3839 1927 3845 1928
rect 3839 1926 3840 1927
rect 3779 1924 3840 1926
rect 3779 1923 3780 1924
rect 3774 1922 3780 1923
rect 3839 1923 3840 1924
rect 3844 1923 3845 1927
rect 3839 1922 3845 1923
rect 3958 1927 3964 1928
rect 3958 1923 3959 1927
rect 3963 1926 3964 1927
rect 3967 1927 3973 1928
rect 3967 1926 3968 1927
rect 3963 1924 3968 1926
rect 3963 1923 3964 1924
rect 3958 1922 3964 1923
rect 3967 1923 3968 1924
rect 3972 1923 3973 1927
rect 3967 1922 3973 1923
rect 3451 1916 3681 1918
rect 3451 1915 3452 1916
rect 3446 1914 3452 1915
rect 2595 1912 2650 1914
rect 2595 1911 2596 1912
rect 2590 1910 2596 1911
rect 2006 1907 2012 1908
rect 2006 1906 2007 1907
rect 1801 1904 1874 1906
rect 1985 1904 2007 1906
rect 966 1902 972 1903
rect 2006 1903 2007 1904
rect 2011 1903 2012 1907
rect 2006 1902 2012 1903
rect 2479 1907 2485 1908
rect 2479 1903 2480 1907
rect 2484 1906 2485 1907
rect 2639 1907 2645 1908
rect 2639 1906 2640 1907
rect 2484 1904 2640 1906
rect 2484 1903 2485 1904
rect 2479 1902 2485 1903
rect 2639 1903 2640 1904
rect 2644 1903 2645 1907
rect 2648 1906 2650 1912
rect 2727 1907 2733 1908
rect 2727 1906 2728 1907
rect 2648 1904 2728 1906
rect 2639 1902 2645 1903
rect 2727 1903 2728 1904
rect 2732 1903 2733 1907
rect 2727 1902 2733 1903
rect 2862 1907 2868 1908
rect 2862 1903 2863 1907
rect 2867 1906 2868 1907
rect 2959 1907 2965 1908
rect 2959 1906 2960 1907
rect 2867 1904 2960 1906
rect 2867 1903 2868 1904
rect 2862 1902 2868 1903
rect 2959 1903 2960 1904
rect 2964 1903 2965 1907
rect 2959 1902 2965 1903
rect 3175 1907 3181 1908
rect 3175 1903 3176 1907
rect 3180 1906 3181 1907
rect 3295 1907 3301 1908
rect 3295 1906 3296 1907
rect 3180 1904 3296 1906
rect 3180 1903 3181 1904
rect 3175 1902 3181 1903
rect 3295 1903 3296 1904
rect 3300 1903 3301 1907
rect 3295 1902 3301 1903
rect 3383 1907 3389 1908
rect 3383 1903 3384 1907
rect 3388 1906 3389 1907
rect 3391 1907 3397 1908
rect 3391 1906 3392 1907
rect 3388 1904 3392 1906
rect 3388 1903 3389 1904
rect 3383 1902 3389 1903
rect 3391 1903 3392 1904
rect 3396 1903 3397 1907
rect 3391 1902 3397 1903
rect 3583 1907 3589 1908
rect 3583 1903 3584 1907
rect 3588 1906 3589 1907
rect 3606 1907 3612 1908
rect 3606 1906 3607 1907
rect 3588 1904 3607 1906
rect 3588 1903 3589 1904
rect 3583 1902 3589 1903
rect 3606 1903 3607 1904
rect 3611 1903 3612 1907
rect 3783 1907 3789 1908
rect 3783 1906 3784 1907
rect 3606 1902 3612 1903
rect 3679 1904 3784 1906
rect 2406 1899 2412 1900
rect 110 1896 116 1897
rect 110 1892 111 1896
rect 115 1892 116 1896
rect 110 1891 116 1892
rect 2030 1896 2036 1897
rect 2030 1892 2031 1896
rect 2035 1892 2036 1896
rect 2406 1895 2407 1899
rect 2411 1895 2412 1899
rect 2406 1894 2412 1895
rect 2654 1899 2660 1900
rect 2654 1895 2655 1899
rect 2659 1895 2660 1899
rect 2654 1894 2660 1895
rect 2886 1899 2892 1900
rect 2886 1895 2887 1899
rect 2891 1895 2892 1899
rect 2886 1894 2892 1895
rect 3102 1899 3108 1900
rect 3102 1895 3103 1899
rect 3107 1895 3108 1899
rect 3102 1894 3108 1895
rect 3310 1899 3316 1900
rect 3310 1895 3311 1899
rect 3315 1895 3316 1899
rect 3310 1894 3316 1895
rect 3510 1899 3516 1900
rect 3510 1895 3511 1899
rect 3515 1895 3516 1899
rect 3510 1894 3516 1895
rect 2030 1891 2036 1892
rect 2975 1891 2981 1892
rect 2975 1890 2976 1891
rect 2937 1888 2976 1890
rect 2430 1887 2436 1888
rect 2430 1883 2431 1887
rect 2435 1883 2436 1887
rect 2975 1887 2976 1888
rect 2980 1887 2981 1891
rect 3166 1891 3172 1892
rect 3166 1890 3167 1891
rect 3153 1888 3167 1890
rect 2975 1886 2981 1887
rect 3166 1887 3167 1888
rect 3171 1887 3172 1891
rect 3679 1890 3681 1904
rect 3783 1903 3784 1904
rect 3788 1903 3789 1907
rect 3783 1902 3789 1903
rect 3966 1907 3973 1908
rect 3966 1903 3967 1907
rect 3972 1903 3973 1907
rect 3966 1902 3973 1903
rect 3710 1899 3716 1900
rect 3710 1895 3711 1899
rect 3715 1895 3716 1899
rect 3710 1894 3716 1895
rect 3894 1899 3900 1900
rect 3894 1895 3895 1899
rect 3899 1895 3900 1899
rect 3894 1894 3900 1895
rect 3774 1891 3780 1892
rect 3774 1890 3775 1891
rect 3561 1888 3681 1890
rect 3761 1888 3775 1890
rect 3166 1886 3172 1887
rect 3774 1887 3775 1888
rect 3779 1887 3780 1891
rect 3774 1886 3780 1887
rect 3886 1887 3892 1888
rect 2430 1882 2436 1883
rect 3886 1883 3887 1887
rect 3891 1883 3892 1887
rect 3886 1882 3892 1883
rect 2070 1880 2076 1881
rect 110 1879 116 1880
rect 110 1875 111 1879
rect 115 1875 116 1879
rect 2030 1879 2036 1880
rect 2030 1875 2031 1879
rect 2035 1875 2036 1879
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 3990 1880 3996 1881
rect 3990 1876 3991 1880
rect 3995 1876 3996 1880
rect 3990 1875 3996 1876
rect 110 1874 116 1875
rect 150 1874 156 1875
rect 150 1870 151 1874
rect 155 1870 156 1874
rect 150 1869 156 1870
rect 270 1874 276 1875
rect 270 1870 271 1874
rect 275 1870 276 1874
rect 270 1869 276 1870
rect 406 1874 412 1875
rect 406 1870 407 1874
rect 411 1870 412 1874
rect 406 1869 412 1870
rect 542 1874 548 1875
rect 542 1870 543 1874
rect 547 1870 548 1874
rect 542 1869 548 1870
rect 678 1874 684 1875
rect 678 1870 679 1874
rect 683 1870 684 1874
rect 678 1869 684 1870
rect 822 1874 828 1875
rect 822 1870 823 1874
rect 827 1870 828 1874
rect 822 1869 828 1870
rect 982 1874 988 1875
rect 982 1870 983 1874
rect 987 1870 988 1874
rect 982 1869 988 1870
rect 1158 1874 1164 1875
rect 1158 1870 1159 1874
rect 1163 1870 1164 1874
rect 1158 1869 1164 1870
rect 1342 1874 1348 1875
rect 1342 1870 1343 1874
rect 1347 1870 1348 1874
rect 1342 1869 1348 1870
rect 1542 1874 1548 1875
rect 1542 1870 1543 1874
rect 1547 1870 1548 1874
rect 1542 1869 1548 1870
rect 1750 1874 1756 1875
rect 1750 1870 1751 1874
rect 1755 1870 1756 1874
rect 1750 1869 1756 1870
rect 1934 1874 1940 1875
rect 2030 1874 2036 1875
rect 1934 1870 1935 1874
rect 1939 1870 1940 1874
rect 1934 1869 1940 1870
rect 2070 1863 2076 1864
rect 2070 1859 2071 1863
rect 2075 1859 2076 1863
rect 3990 1863 3996 1864
rect 3990 1859 3991 1863
rect 3995 1859 3996 1863
rect 2070 1858 2076 1859
rect 2406 1858 2412 1859
rect 1042 1855 1048 1856
rect 1042 1851 1043 1855
rect 1047 1854 1048 1855
rect 1550 1855 1556 1856
rect 1550 1854 1551 1855
rect 1047 1852 1551 1854
rect 1047 1851 1048 1852
rect 1042 1850 1048 1851
rect 1550 1851 1551 1852
rect 1555 1851 1556 1855
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2654 1858 2660 1859
rect 2654 1854 2655 1858
rect 2659 1854 2660 1858
rect 2654 1853 2660 1854
rect 2886 1858 2892 1859
rect 2886 1854 2887 1858
rect 2891 1854 2892 1858
rect 2886 1853 2892 1854
rect 3102 1858 3108 1859
rect 3102 1854 3103 1858
rect 3107 1854 3108 1858
rect 3102 1853 3108 1854
rect 3310 1858 3316 1859
rect 3310 1854 3311 1858
rect 3315 1854 3316 1858
rect 3310 1853 3316 1854
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 3710 1858 3716 1859
rect 3710 1854 3711 1858
rect 3715 1854 3716 1858
rect 3710 1853 3716 1854
rect 3894 1858 3900 1859
rect 3990 1858 3996 1859
rect 3894 1854 3895 1858
rect 3899 1854 3900 1858
rect 3894 1853 3900 1854
rect 1550 1850 1556 1851
rect 150 1834 156 1835
rect 150 1830 151 1834
rect 155 1830 156 1834
rect 110 1829 116 1830
rect 150 1829 156 1830
rect 286 1834 292 1835
rect 286 1830 287 1834
rect 291 1830 292 1834
rect 286 1829 292 1830
rect 446 1834 452 1835
rect 446 1830 447 1834
rect 451 1830 452 1834
rect 446 1829 452 1830
rect 598 1834 604 1835
rect 598 1830 599 1834
rect 603 1830 604 1834
rect 598 1829 604 1830
rect 750 1834 756 1835
rect 750 1830 751 1834
rect 755 1830 756 1834
rect 750 1829 756 1830
rect 918 1834 924 1835
rect 918 1830 919 1834
rect 923 1830 924 1834
rect 918 1829 924 1830
rect 1102 1834 1108 1835
rect 1102 1830 1103 1834
rect 1107 1830 1108 1834
rect 1102 1829 1108 1830
rect 1302 1834 1308 1835
rect 1302 1830 1303 1834
rect 1307 1830 1308 1834
rect 1302 1829 1308 1830
rect 1510 1834 1516 1835
rect 1510 1830 1511 1834
rect 1515 1830 1516 1834
rect 1510 1829 1516 1830
rect 1734 1834 1740 1835
rect 1734 1830 1735 1834
rect 1739 1830 1740 1834
rect 1734 1829 1740 1830
rect 1934 1834 1940 1835
rect 1934 1830 1935 1834
rect 1939 1830 1940 1834
rect 1934 1829 1940 1830
rect 2030 1829 2036 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 2030 1825 2031 1829
rect 2035 1825 2036 1829
rect 2030 1824 2036 1825
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2070 1821 2076 1822
rect 2110 1821 2116 1822
rect 2382 1826 2388 1827
rect 2382 1822 2383 1826
rect 2387 1822 2388 1826
rect 2382 1821 2388 1822
rect 2646 1826 2652 1827
rect 2646 1822 2647 1826
rect 2651 1822 2652 1826
rect 2646 1821 2652 1822
rect 2886 1826 2892 1827
rect 2886 1822 2887 1826
rect 2891 1822 2892 1826
rect 2886 1821 2892 1822
rect 3094 1826 3100 1827
rect 3094 1822 3095 1826
rect 3099 1822 3100 1826
rect 3094 1821 3100 1822
rect 3286 1826 3292 1827
rect 3286 1822 3287 1826
rect 3291 1822 3292 1826
rect 3286 1821 3292 1822
rect 3454 1826 3460 1827
rect 3454 1822 3455 1826
rect 3459 1822 3460 1826
rect 3454 1821 3460 1822
rect 3614 1826 3620 1827
rect 3614 1822 3615 1826
rect 3619 1822 3620 1826
rect 3614 1821 3620 1822
rect 3766 1826 3772 1827
rect 3766 1822 3767 1826
rect 3771 1822 3772 1826
rect 3766 1821 3772 1822
rect 3894 1826 3900 1827
rect 3894 1822 3895 1826
rect 3899 1822 3900 1826
rect 3894 1821 3900 1822
rect 3990 1821 3996 1822
rect 2070 1817 2071 1821
rect 2075 1817 2076 1821
rect 2070 1816 2076 1817
rect 3990 1817 3991 1821
rect 3995 1817 3996 1821
rect 3990 1816 3996 1817
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 110 1807 116 1808
rect 2030 1812 2036 1813
rect 2030 1808 2031 1812
rect 2035 1808 2036 1812
rect 2030 1807 2036 1808
rect 2070 1804 2076 1805
rect 3990 1804 3996 1805
rect 231 1803 237 1804
rect 231 1802 232 1803
rect 201 1800 232 1802
rect 231 1799 232 1800
rect 236 1799 237 1803
rect 426 1803 432 1804
rect 426 1802 427 1803
rect 337 1800 427 1802
rect 231 1798 237 1799
rect 426 1799 427 1800
rect 431 1799 432 1803
rect 559 1803 565 1804
rect 559 1802 560 1803
rect 497 1800 560 1802
rect 426 1798 432 1799
rect 559 1799 560 1800
rect 564 1799 565 1803
rect 559 1798 565 1799
rect 614 1803 620 1804
rect 614 1799 615 1803
rect 619 1799 620 1803
rect 1042 1803 1048 1804
rect 1042 1802 1043 1803
rect 969 1800 1043 1802
rect 614 1798 620 1799
rect 1042 1799 1043 1800
rect 1047 1799 1048 1803
rect 2062 1803 2068 1804
rect 2062 1802 2063 1803
rect 1985 1800 2063 1802
rect 1042 1798 1048 1799
rect 2062 1799 2063 1800
rect 2067 1799 2068 1803
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 3902 1803 3908 1804
rect 3902 1802 3903 1803
rect 2070 1799 2076 1800
rect 3884 1800 3903 1802
rect 2062 1798 2068 1799
rect 2182 1795 2188 1796
rect 2182 1794 2183 1795
rect 150 1793 156 1794
rect 150 1789 151 1793
rect 155 1789 156 1793
rect 150 1788 156 1789
rect 286 1793 292 1794
rect 286 1789 287 1793
rect 291 1789 292 1793
rect 286 1788 292 1789
rect 446 1793 452 1794
rect 446 1789 447 1793
rect 451 1789 452 1793
rect 446 1788 452 1789
rect 598 1793 604 1794
rect 598 1789 599 1793
rect 603 1789 604 1793
rect 598 1788 604 1789
rect 750 1793 756 1794
rect 750 1789 751 1793
rect 755 1789 756 1793
rect 750 1788 756 1789
rect 918 1793 924 1794
rect 918 1789 919 1793
rect 923 1789 924 1793
rect 918 1788 924 1789
rect 1102 1793 1108 1794
rect 1102 1789 1103 1793
rect 1107 1789 1108 1793
rect 1102 1788 1108 1789
rect 1302 1793 1308 1794
rect 1302 1789 1303 1793
rect 1307 1789 1308 1793
rect 1302 1788 1308 1789
rect 1510 1793 1516 1794
rect 1510 1789 1511 1793
rect 1515 1789 1516 1793
rect 1510 1788 1516 1789
rect 1734 1793 1740 1794
rect 1734 1789 1735 1793
rect 1739 1789 1740 1793
rect 1734 1788 1740 1789
rect 1934 1793 1940 1794
rect 1934 1789 1935 1793
rect 1939 1789 1940 1793
rect 2161 1792 2183 1794
rect 2182 1791 2183 1792
rect 2187 1791 2188 1795
rect 2578 1795 2584 1796
rect 2578 1794 2579 1795
rect 2433 1792 2579 1794
rect 2182 1790 2188 1791
rect 2578 1791 2579 1792
rect 2583 1791 2584 1795
rect 2862 1795 2868 1796
rect 2862 1794 2863 1795
rect 2697 1792 2863 1794
rect 2578 1790 2584 1791
rect 2862 1791 2863 1792
rect 2867 1791 2868 1795
rect 3078 1795 3084 1796
rect 3078 1794 3079 1795
rect 2937 1792 3079 1794
rect 2862 1790 2868 1791
rect 3078 1791 3079 1792
rect 3083 1791 3084 1795
rect 3358 1795 3364 1796
rect 3358 1794 3359 1795
rect 3337 1792 3359 1794
rect 3078 1790 3084 1791
rect 3358 1791 3359 1792
rect 3363 1791 3364 1795
rect 3562 1795 3568 1796
rect 3562 1794 3563 1795
rect 3505 1792 3563 1794
rect 3358 1790 3364 1791
rect 3562 1791 3563 1792
rect 3567 1791 3568 1795
rect 3562 1790 3568 1791
rect 3606 1795 3612 1796
rect 3606 1791 3607 1795
rect 3611 1791 3612 1795
rect 3884 1794 3886 1800
rect 3902 1799 3903 1800
rect 3907 1799 3908 1803
rect 3990 1800 3991 1804
rect 3995 1800 3996 1804
rect 3990 1799 3996 1800
rect 3902 1798 3908 1799
rect 3966 1795 3972 1796
rect 3966 1794 3967 1795
rect 3817 1792 3886 1794
rect 3945 1792 3967 1794
rect 3606 1790 3612 1791
rect 3966 1791 3967 1792
rect 3971 1791 3972 1795
rect 3966 1790 3972 1791
rect 1934 1788 1940 1789
rect 2110 1785 2116 1786
rect 222 1783 229 1784
rect 222 1779 223 1783
rect 228 1779 229 1783
rect 222 1778 229 1779
rect 231 1783 237 1784
rect 231 1779 232 1783
rect 236 1782 237 1783
rect 359 1783 365 1784
rect 359 1782 360 1783
rect 236 1780 360 1782
rect 236 1779 237 1780
rect 231 1778 237 1779
rect 359 1779 360 1780
rect 364 1779 365 1783
rect 359 1778 365 1779
rect 426 1783 432 1784
rect 426 1779 427 1783
rect 431 1782 432 1783
rect 519 1783 525 1784
rect 519 1782 520 1783
rect 431 1780 520 1782
rect 431 1779 432 1780
rect 426 1778 432 1779
rect 519 1779 520 1780
rect 524 1779 525 1783
rect 519 1778 525 1779
rect 671 1783 677 1784
rect 671 1779 672 1783
rect 676 1782 677 1783
rect 735 1783 741 1784
rect 735 1782 736 1783
rect 676 1780 736 1782
rect 676 1779 677 1780
rect 671 1778 677 1779
rect 735 1779 736 1780
rect 740 1779 741 1783
rect 735 1778 741 1779
rect 814 1783 820 1784
rect 814 1779 815 1783
rect 819 1782 820 1783
rect 823 1783 829 1784
rect 823 1782 824 1783
rect 819 1780 824 1782
rect 819 1779 820 1780
rect 814 1778 820 1779
rect 823 1779 824 1780
rect 828 1779 829 1783
rect 823 1778 829 1779
rect 991 1783 997 1784
rect 991 1779 992 1783
rect 996 1782 997 1783
rect 1087 1783 1093 1784
rect 1087 1782 1088 1783
rect 996 1780 1088 1782
rect 996 1779 997 1780
rect 991 1778 997 1779
rect 1087 1779 1088 1780
rect 1092 1779 1093 1783
rect 1087 1778 1093 1779
rect 1175 1783 1181 1784
rect 1175 1779 1176 1783
rect 1180 1782 1181 1783
rect 1287 1783 1293 1784
rect 1287 1782 1288 1783
rect 1180 1780 1288 1782
rect 1180 1779 1181 1780
rect 1175 1778 1181 1779
rect 1287 1779 1288 1780
rect 1292 1779 1293 1783
rect 1287 1778 1293 1779
rect 1375 1783 1381 1784
rect 1375 1779 1376 1783
rect 1380 1782 1381 1783
rect 1495 1783 1501 1784
rect 1495 1782 1496 1783
rect 1380 1780 1496 1782
rect 1380 1779 1381 1780
rect 1375 1778 1381 1779
rect 1495 1779 1496 1780
rect 1500 1779 1501 1783
rect 1495 1778 1501 1779
rect 1583 1783 1589 1784
rect 1583 1779 1584 1783
rect 1588 1782 1589 1783
rect 1719 1783 1725 1784
rect 1719 1782 1720 1783
rect 1588 1780 1720 1782
rect 1588 1779 1589 1780
rect 1583 1778 1589 1779
rect 1719 1779 1720 1780
rect 1724 1779 1725 1783
rect 1719 1778 1725 1779
rect 1742 1783 1748 1784
rect 1742 1779 1743 1783
rect 1747 1782 1748 1783
rect 1807 1783 1813 1784
rect 1807 1782 1808 1783
rect 1747 1780 1808 1782
rect 1747 1779 1748 1780
rect 1742 1778 1748 1779
rect 1807 1779 1808 1780
rect 1812 1779 1813 1783
rect 1807 1778 1813 1779
rect 2006 1783 2013 1784
rect 2006 1779 2007 1783
rect 2012 1779 2013 1783
rect 2110 1781 2111 1785
rect 2115 1781 2116 1785
rect 2110 1780 2116 1781
rect 2382 1785 2388 1786
rect 2382 1781 2383 1785
rect 2387 1781 2388 1785
rect 2382 1780 2388 1781
rect 2646 1785 2652 1786
rect 2646 1781 2647 1785
rect 2651 1781 2652 1785
rect 2646 1780 2652 1781
rect 2886 1785 2892 1786
rect 2886 1781 2887 1785
rect 2891 1781 2892 1785
rect 2886 1780 2892 1781
rect 3094 1785 3100 1786
rect 3094 1781 3095 1785
rect 3099 1781 3100 1785
rect 3094 1780 3100 1781
rect 3286 1785 3292 1786
rect 3286 1781 3287 1785
rect 3291 1781 3292 1785
rect 3286 1780 3292 1781
rect 3454 1785 3460 1786
rect 3454 1781 3455 1785
rect 3459 1781 3460 1785
rect 3454 1780 3460 1781
rect 3614 1785 3620 1786
rect 3614 1781 3615 1785
rect 3619 1781 3620 1785
rect 3614 1780 3620 1781
rect 3766 1785 3772 1786
rect 3766 1781 3767 1785
rect 3771 1781 3772 1785
rect 3766 1780 3772 1781
rect 3894 1785 3900 1786
rect 3894 1781 3895 1785
rect 3899 1781 3900 1785
rect 3894 1780 3900 1781
rect 2006 1778 2013 1779
rect 2062 1775 2068 1776
rect 2062 1771 2063 1775
rect 2067 1774 2068 1775
rect 2183 1775 2189 1776
rect 2183 1774 2184 1775
rect 2067 1772 2184 1774
rect 2067 1771 2068 1772
rect 2062 1770 2068 1771
rect 2183 1771 2184 1772
rect 2188 1771 2189 1775
rect 2183 1770 2189 1771
rect 2430 1775 2436 1776
rect 2430 1771 2431 1775
rect 2435 1774 2436 1775
rect 2455 1775 2461 1776
rect 2455 1774 2456 1775
rect 2435 1772 2456 1774
rect 2435 1771 2436 1772
rect 2430 1770 2436 1771
rect 2455 1771 2456 1772
rect 2460 1771 2461 1775
rect 2455 1770 2461 1771
rect 2719 1775 2725 1776
rect 2719 1771 2720 1775
rect 2724 1774 2725 1775
rect 2959 1775 2965 1776
rect 2724 1772 2841 1774
rect 2724 1771 2725 1772
rect 2719 1770 2725 1771
rect 279 1763 285 1764
rect 279 1759 280 1763
rect 284 1762 285 1763
rect 367 1763 373 1764
rect 367 1762 368 1763
rect 284 1760 368 1762
rect 284 1759 285 1760
rect 279 1758 285 1759
rect 367 1759 368 1760
rect 372 1759 373 1763
rect 367 1758 373 1759
rect 455 1763 461 1764
rect 455 1759 456 1763
rect 460 1762 461 1763
rect 551 1763 557 1764
rect 551 1762 552 1763
rect 460 1760 552 1762
rect 460 1759 461 1760
rect 455 1758 461 1759
rect 551 1759 552 1760
rect 556 1759 557 1763
rect 551 1758 557 1759
rect 559 1763 565 1764
rect 559 1759 560 1763
rect 564 1762 565 1763
rect 639 1763 645 1764
rect 639 1762 640 1763
rect 564 1760 640 1762
rect 564 1759 565 1760
rect 559 1758 565 1759
rect 639 1759 640 1760
rect 644 1759 645 1763
rect 639 1758 645 1759
rect 823 1763 829 1764
rect 823 1759 824 1763
rect 828 1762 829 1763
rect 919 1763 925 1764
rect 919 1762 920 1763
rect 828 1760 920 1762
rect 828 1759 829 1760
rect 823 1758 829 1759
rect 919 1759 920 1760
rect 924 1759 925 1763
rect 919 1758 925 1759
rect 1006 1763 1013 1764
rect 1006 1759 1007 1763
rect 1012 1759 1013 1763
rect 1006 1758 1013 1759
rect 1183 1763 1189 1764
rect 1183 1759 1184 1763
rect 1188 1762 1189 1763
rect 1263 1763 1269 1764
rect 1263 1762 1264 1763
rect 1188 1760 1264 1762
rect 1188 1759 1189 1760
rect 1183 1758 1189 1759
rect 1263 1759 1264 1760
rect 1268 1759 1269 1763
rect 1263 1758 1269 1759
rect 1351 1763 1357 1764
rect 1351 1759 1352 1763
rect 1356 1762 1357 1763
rect 1439 1763 1445 1764
rect 1439 1762 1440 1763
rect 1356 1760 1440 1762
rect 1356 1759 1357 1760
rect 1351 1758 1357 1759
rect 1439 1759 1440 1760
rect 1444 1759 1445 1763
rect 1439 1758 1445 1759
rect 1527 1763 1533 1764
rect 1527 1759 1528 1763
rect 1532 1762 1533 1763
rect 1615 1763 1621 1764
rect 1615 1762 1616 1763
rect 1532 1760 1616 1762
rect 1532 1759 1533 1760
rect 1527 1758 1533 1759
rect 1615 1759 1616 1760
rect 1620 1759 1621 1763
rect 1615 1758 1621 1759
rect 1702 1763 1709 1764
rect 1702 1759 1703 1763
rect 1708 1759 1709 1763
rect 1702 1758 1709 1759
rect 2182 1763 2189 1764
rect 2182 1759 2183 1763
rect 2188 1759 2189 1763
rect 2359 1763 2365 1764
rect 2359 1762 2360 1763
rect 2182 1758 2189 1759
rect 2232 1760 2360 1762
rect 206 1755 212 1756
rect 206 1751 207 1755
rect 211 1751 212 1755
rect 206 1750 212 1751
rect 382 1755 388 1756
rect 382 1751 383 1755
rect 387 1751 388 1755
rect 382 1750 388 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 750 1755 756 1756
rect 750 1751 751 1755
rect 755 1751 756 1755
rect 750 1750 756 1751
rect 934 1755 940 1756
rect 934 1751 935 1755
rect 939 1751 940 1755
rect 934 1750 940 1751
rect 1110 1755 1116 1756
rect 1110 1751 1111 1755
rect 1115 1751 1116 1755
rect 1110 1750 1116 1751
rect 1278 1755 1284 1756
rect 1278 1751 1279 1755
rect 1283 1751 1284 1755
rect 1278 1750 1284 1751
rect 1454 1755 1460 1756
rect 1454 1751 1455 1755
rect 1459 1751 1460 1755
rect 1454 1750 1460 1751
rect 1630 1755 1636 1756
rect 1630 1751 1631 1755
rect 1635 1751 1636 1755
rect 1630 1750 1636 1751
rect 2110 1755 2116 1756
rect 2110 1751 2111 1755
rect 2115 1751 2116 1755
rect 2110 1750 2116 1751
rect 366 1747 372 1748
rect 366 1746 367 1747
rect 257 1744 367 1746
rect 366 1743 367 1744
rect 371 1743 372 1747
rect 814 1747 820 1748
rect 814 1746 815 1747
rect 801 1744 815 1746
rect 366 1742 372 1743
rect 814 1743 815 1744
rect 819 1743 820 1747
rect 1262 1747 1268 1748
rect 1262 1746 1263 1747
rect 1161 1744 1263 1746
rect 814 1742 820 1743
rect 1262 1743 1263 1744
rect 1267 1743 1268 1747
rect 2232 1746 2234 1760
rect 2359 1759 2360 1760
rect 2364 1759 2365 1763
rect 2567 1763 2573 1764
rect 2567 1762 2568 1763
rect 2359 1758 2365 1759
rect 2420 1760 2568 1762
rect 2286 1755 2292 1756
rect 2286 1751 2287 1755
rect 2291 1751 2292 1755
rect 2286 1750 2292 1751
rect 2420 1746 2422 1760
rect 2567 1759 2568 1760
rect 2572 1759 2573 1763
rect 2567 1758 2573 1759
rect 2578 1763 2584 1764
rect 2578 1759 2579 1763
rect 2583 1762 2584 1763
rect 2783 1763 2789 1764
rect 2783 1762 2784 1763
rect 2583 1760 2784 1762
rect 2583 1759 2584 1760
rect 2578 1758 2584 1759
rect 2783 1759 2784 1760
rect 2788 1759 2789 1763
rect 2839 1762 2841 1772
rect 2959 1771 2960 1775
rect 2964 1774 2965 1775
rect 3079 1775 3085 1776
rect 3079 1774 3080 1775
rect 2964 1772 3080 1774
rect 2964 1771 2965 1772
rect 2959 1770 2965 1771
rect 3079 1771 3080 1772
rect 3084 1771 3085 1775
rect 3079 1770 3085 1771
rect 3166 1775 3173 1776
rect 3166 1771 3167 1775
rect 3172 1771 3173 1775
rect 3359 1775 3365 1776
rect 3359 1774 3360 1775
rect 3166 1770 3173 1771
rect 3176 1772 3360 1774
rect 3078 1767 3084 1768
rect 2991 1764 2997 1765
rect 2903 1763 2909 1764
rect 2903 1762 2904 1763
rect 2839 1760 2904 1762
rect 2783 1758 2789 1759
rect 2903 1759 2904 1760
rect 2908 1759 2909 1763
rect 2903 1758 2909 1759
rect 2990 1763 2992 1764
rect 2990 1759 2991 1763
rect 2996 1760 2997 1764
rect 3078 1763 3079 1767
rect 3083 1766 3084 1767
rect 3176 1766 3178 1772
rect 3359 1771 3360 1772
rect 3364 1771 3365 1775
rect 3359 1770 3365 1771
rect 3526 1775 3533 1776
rect 3526 1771 3527 1775
rect 3532 1771 3533 1775
rect 3526 1770 3533 1771
rect 3562 1775 3568 1776
rect 3562 1771 3563 1775
rect 3567 1774 3568 1775
rect 3687 1775 3693 1776
rect 3687 1774 3688 1775
rect 3567 1772 3688 1774
rect 3567 1771 3568 1772
rect 3562 1770 3568 1771
rect 3687 1771 3688 1772
rect 3692 1771 3693 1775
rect 3687 1770 3693 1771
rect 3839 1775 3845 1776
rect 3839 1771 3840 1775
rect 3844 1774 3845 1775
rect 3886 1775 3892 1776
rect 3886 1774 3887 1775
rect 3844 1772 3887 1774
rect 3844 1771 3845 1772
rect 3839 1770 3845 1771
rect 3886 1771 3887 1772
rect 3891 1771 3892 1775
rect 3886 1770 3892 1771
rect 3902 1775 3908 1776
rect 3902 1771 3903 1775
rect 3907 1774 3908 1775
rect 3967 1775 3973 1776
rect 3967 1774 3968 1775
rect 3907 1772 3968 1774
rect 3907 1771 3908 1772
rect 3902 1770 3908 1771
rect 3967 1771 3968 1772
rect 3972 1771 3973 1775
rect 3967 1770 3973 1771
rect 3083 1764 3178 1766
rect 3083 1763 3084 1764
rect 3078 1762 3084 1763
rect 3191 1763 3197 1764
rect 2995 1759 2997 1760
rect 3191 1759 3192 1763
rect 3196 1762 3197 1763
rect 3303 1763 3309 1764
rect 3303 1762 3304 1763
rect 3196 1760 3304 1762
rect 3196 1759 3197 1760
rect 2990 1758 2996 1759
rect 3191 1758 3197 1759
rect 3303 1759 3304 1760
rect 3308 1759 3309 1763
rect 3303 1758 3309 1759
rect 3358 1763 3364 1764
rect 3358 1759 3359 1763
rect 3363 1762 3364 1763
rect 3391 1763 3397 1764
rect 3391 1762 3392 1763
rect 3363 1760 3392 1762
rect 3363 1759 3364 1760
rect 3358 1758 3364 1759
rect 3391 1759 3392 1760
rect 3396 1759 3397 1763
rect 3391 1758 3397 1759
rect 3583 1763 3589 1764
rect 3583 1759 3584 1763
rect 3588 1762 3589 1763
rect 3687 1763 3693 1764
rect 3687 1762 3688 1763
rect 3588 1760 3688 1762
rect 3588 1759 3589 1760
rect 3583 1758 3589 1759
rect 3687 1759 3688 1760
rect 3692 1759 3693 1763
rect 3687 1758 3693 1759
rect 3775 1763 3781 1764
rect 3775 1759 3776 1763
rect 3780 1762 3781 1763
rect 3879 1763 3885 1764
rect 3879 1762 3880 1763
rect 3780 1760 3880 1762
rect 3780 1759 3781 1760
rect 3775 1758 3781 1759
rect 3879 1759 3880 1760
rect 3884 1759 3885 1763
rect 3879 1758 3885 1759
rect 3966 1763 3973 1764
rect 3966 1759 3967 1763
rect 3972 1759 3973 1763
rect 3966 1758 3973 1759
rect 2494 1755 2500 1756
rect 2494 1751 2495 1755
rect 2499 1751 2500 1755
rect 2494 1750 2500 1751
rect 2710 1755 2716 1756
rect 2710 1751 2711 1755
rect 2715 1751 2716 1755
rect 2710 1750 2716 1751
rect 2918 1755 2924 1756
rect 2918 1751 2919 1755
rect 2923 1751 2924 1755
rect 2918 1750 2924 1751
rect 3118 1755 3124 1756
rect 3118 1751 3119 1755
rect 3123 1751 3124 1755
rect 3118 1750 3124 1751
rect 3318 1755 3324 1756
rect 3318 1751 3319 1755
rect 3323 1751 3324 1755
rect 3318 1750 3324 1751
rect 3510 1755 3516 1756
rect 3510 1751 3511 1755
rect 3515 1751 3516 1755
rect 3510 1750 3516 1751
rect 3702 1755 3708 1756
rect 3702 1751 3703 1755
rect 3707 1751 3708 1755
rect 3702 1750 3708 1751
rect 3894 1755 3900 1756
rect 3894 1751 3895 1755
rect 3899 1751 3900 1755
rect 3894 1750 3900 1751
rect 2161 1744 2234 1746
rect 2337 1744 2422 1746
rect 1262 1742 1268 1743
rect 2486 1743 2492 1744
rect 2486 1739 2487 1743
rect 2491 1739 2492 1743
rect 2486 1738 2492 1739
rect 2726 1743 2732 1744
rect 2726 1739 2727 1743
rect 2731 1739 2732 1743
rect 2726 1738 2732 1739
rect 3134 1743 3140 1744
rect 3134 1739 3135 1743
rect 3139 1739 3140 1743
rect 3134 1738 3140 1739
rect 3526 1743 3532 1744
rect 3526 1739 3527 1743
rect 3531 1739 3532 1743
rect 3526 1738 3532 1739
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 2030 1736 2036 1737
rect 2030 1732 2031 1736
rect 2035 1732 2036 1736
rect 2030 1731 2036 1732
rect 2070 1736 2076 1737
rect 2070 1732 2071 1736
rect 2075 1732 2076 1736
rect 2070 1731 2076 1732
rect 3990 1736 3996 1737
rect 3990 1732 3991 1736
rect 3995 1732 3996 1736
rect 3990 1731 3996 1732
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 2030 1719 2036 1720
rect 2030 1715 2031 1719
rect 2035 1715 2036 1719
rect 110 1714 116 1715
rect 206 1714 212 1715
rect 206 1710 207 1714
rect 211 1710 212 1714
rect 206 1709 212 1710
rect 382 1714 388 1715
rect 382 1710 383 1714
rect 387 1710 388 1714
rect 382 1709 388 1710
rect 566 1714 572 1715
rect 566 1710 567 1714
rect 571 1710 572 1714
rect 566 1709 572 1710
rect 750 1714 756 1715
rect 750 1710 751 1714
rect 755 1710 756 1714
rect 750 1709 756 1710
rect 934 1714 940 1715
rect 934 1710 935 1714
rect 939 1710 940 1714
rect 934 1709 940 1710
rect 1110 1714 1116 1715
rect 1110 1710 1111 1714
rect 1115 1710 1116 1714
rect 1110 1709 1116 1710
rect 1278 1714 1284 1715
rect 1278 1710 1279 1714
rect 1283 1710 1284 1714
rect 1278 1709 1284 1710
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1630 1714 1636 1715
rect 2030 1714 2036 1715
rect 2070 1719 2076 1720
rect 2070 1715 2071 1719
rect 2075 1715 2076 1719
rect 3990 1719 3996 1720
rect 3990 1715 3991 1719
rect 3995 1715 3996 1719
rect 2070 1714 2076 1715
rect 2110 1714 2116 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 2110 1710 2111 1714
rect 2115 1710 2116 1714
rect 2110 1709 2116 1710
rect 2286 1714 2292 1715
rect 2286 1710 2287 1714
rect 2291 1710 2292 1714
rect 2286 1709 2292 1710
rect 2494 1714 2500 1715
rect 2494 1710 2495 1714
rect 2499 1710 2500 1714
rect 2494 1709 2500 1710
rect 2710 1714 2716 1715
rect 2710 1710 2711 1714
rect 2715 1710 2716 1714
rect 2710 1709 2716 1710
rect 2918 1714 2924 1715
rect 2918 1710 2919 1714
rect 2923 1710 2924 1714
rect 2918 1709 2924 1710
rect 3118 1714 3124 1715
rect 3118 1710 3119 1714
rect 3123 1710 3124 1714
rect 3118 1709 3124 1710
rect 3318 1714 3324 1715
rect 3318 1710 3319 1714
rect 3323 1710 3324 1714
rect 3318 1709 3324 1710
rect 3510 1714 3516 1715
rect 3510 1710 3511 1714
rect 3515 1710 3516 1714
rect 3510 1709 3516 1710
rect 3702 1714 3708 1715
rect 3702 1710 3703 1714
rect 3707 1710 3708 1714
rect 3702 1709 3708 1710
rect 3894 1714 3900 1715
rect 3990 1714 3996 1715
rect 3894 1710 3895 1714
rect 3899 1710 3900 1714
rect 3894 1709 3900 1710
rect 302 1682 308 1683
rect 302 1678 303 1682
rect 307 1678 308 1682
rect 110 1677 116 1678
rect 302 1677 308 1678
rect 534 1682 540 1683
rect 534 1678 535 1682
rect 539 1678 540 1682
rect 534 1677 540 1678
rect 766 1682 772 1683
rect 766 1678 767 1682
rect 771 1678 772 1682
rect 766 1677 772 1678
rect 982 1682 988 1683
rect 982 1678 983 1682
rect 987 1678 988 1682
rect 982 1677 988 1678
rect 1190 1682 1196 1683
rect 1190 1678 1191 1682
rect 1195 1678 1196 1682
rect 1190 1677 1196 1678
rect 1382 1682 1388 1683
rect 1382 1678 1383 1682
rect 1387 1678 1388 1682
rect 1382 1677 1388 1678
rect 1566 1682 1572 1683
rect 1566 1678 1567 1682
rect 1571 1678 1572 1682
rect 1566 1677 1572 1678
rect 1742 1682 1748 1683
rect 1742 1678 1743 1682
rect 1747 1678 1748 1682
rect 1742 1677 1748 1678
rect 1926 1682 1932 1683
rect 1926 1678 1927 1682
rect 1931 1678 1932 1682
rect 1926 1677 1932 1678
rect 2030 1677 2036 1678
rect 110 1673 111 1677
rect 115 1673 116 1677
rect 110 1672 116 1673
rect 2030 1673 2031 1677
rect 2035 1673 2036 1677
rect 2030 1672 2036 1673
rect 2110 1674 2116 1675
rect 1367 1671 1373 1672
rect 1367 1667 1368 1671
rect 1372 1670 1373 1671
rect 1702 1671 1708 1672
rect 1702 1670 1703 1671
rect 1372 1668 1703 1670
rect 1372 1667 1373 1668
rect 1367 1666 1373 1667
rect 1702 1667 1703 1668
rect 1707 1667 1708 1671
rect 2110 1670 2111 1674
rect 2115 1670 2116 1674
rect 1702 1666 1708 1667
rect 2070 1669 2076 1670
rect 2110 1669 2116 1670
rect 2238 1674 2244 1675
rect 2238 1670 2239 1674
rect 2243 1670 2244 1674
rect 2238 1669 2244 1670
rect 2382 1674 2388 1675
rect 2382 1670 2383 1674
rect 2387 1670 2388 1674
rect 2382 1669 2388 1670
rect 2518 1674 2524 1675
rect 2518 1670 2519 1674
rect 2523 1670 2524 1674
rect 2518 1669 2524 1670
rect 2654 1674 2660 1675
rect 2654 1670 2655 1674
rect 2659 1670 2660 1674
rect 2654 1669 2660 1670
rect 2790 1674 2796 1675
rect 2790 1670 2791 1674
rect 2795 1670 2796 1674
rect 2790 1669 2796 1670
rect 2926 1674 2932 1675
rect 2926 1670 2927 1674
rect 2931 1670 2932 1674
rect 2926 1669 2932 1670
rect 3062 1674 3068 1675
rect 3062 1670 3063 1674
rect 3067 1670 3068 1674
rect 3062 1669 3068 1670
rect 3206 1674 3212 1675
rect 3206 1670 3207 1674
rect 3211 1670 3212 1674
rect 3206 1669 3212 1670
rect 3350 1674 3356 1675
rect 3350 1670 3351 1674
rect 3355 1670 3356 1674
rect 3350 1669 3356 1670
rect 3990 1669 3996 1670
rect 2070 1665 2071 1669
rect 2075 1665 2076 1669
rect 2070 1664 2076 1665
rect 3990 1665 3991 1669
rect 3995 1665 3996 1669
rect 3990 1664 3996 1665
rect 110 1660 116 1661
rect 110 1656 111 1660
rect 115 1656 116 1660
rect 110 1655 116 1656
rect 2030 1660 2036 1661
rect 2030 1656 2031 1660
rect 2035 1656 2036 1660
rect 2030 1655 2036 1656
rect 2070 1652 2076 1653
rect 386 1651 392 1652
rect 386 1650 387 1651
rect 353 1648 387 1650
rect 386 1647 387 1648
rect 391 1647 392 1651
rect 750 1651 756 1652
rect 750 1650 751 1651
rect 585 1648 751 1650
rect 386 1646 392 1647
rect 750 1647 751 1648
rect 755 1647 756 1651
rect 750 1646 756 1647
rect 790 1651 796 1652
rect 790 1647 791 1651
rect 795 1647 796 1651
rect 790 1646 796 1647
rect 1006 1651 1012 1652
rect 1006 1647 1007 1651
rect 1011 1647 1012 1651
rect 1367 1651 1373 1652
rect 1367 1650 1368 1651
rect 1241 1648 1368 1650
rect 1006 1646 1012 1647
rect 1367 1647 1368 1648
rect 1372 1647 1373 1651
rect 2070 1648 2071 1652
rect 2075 1648 2076 1652
rect 2070 1647 2076 1648
rect 3990 1652 3996 1653
rect 3990 1648 3991 1652
rect 3995 1648 3996 1652
rect 3990 1647 3996 1648
rect 1367 1646 1373 1647
rect 2182 1643 2188 1644
rect 2182 1642 2183 1643
rect 302 1641 308 1642
rect 302 1637 303 1641
rect 307 1637 308 1641
rect 302 1636 308 1637
rect 534 1641 540 1642
rect 534 1637 535 1641
rect 539 1637 540 1641
rect 534 1636 540 1637
rect 766 1641 772 1642
rect 766 1637 767 1641
rect 771 1637 772 1641
rect 766 1636 772 1637
rect 982 1641 988 1642
rect 982 1637 983 1641
rect 987 1637 988 1641
rect 982 1636 988 1637
rect 1190 1641 1196 1642
rect 1190 1637 1191 1641
rect 1195 1637 1196 1641
rect 1190 1636 1196 1637
rect 1382 1641 1388 1642
rect 1382 1637 1383 1641
rect 1387 1637 1388 1641
rect 1382 1636 1388 1637
rect 1566 1641 1572 1642
rect 1566 1637 1567 1641
rect 1571 1637 1572 1641
rect 1566 1636 1572 1637
rect 1742 1641 1748 1642
rect 1742 1637 1743 1641
rect 1747 1637 1748 1641
rect 1742 1636 1748 1637
rect 1926 1641 1932 1642
rect 1926 1637 1927 1641
rect 1931 1637 1932 1641
rect 2161 1640 2183 1642
rect 2182 1639 2183 1640
rect 2187 1639 2188 1643
rect 2614 1643 2620 1644
rect 2614 1642 2615 1643
rect 2569 1640 2615 1642
rect 2182 1638 2188 1639
rect 2614 1639 2615 1640
rect 2619 1639 2620 1643
rect 2910 1643 2916 1644
rect 2910 1642 2911 1643
rect 2841 1640 2911 1642
rect 2614 1638 2620 1639
rect 2910 1639 2911 1640
rect 2915 1639 2916 1643
rect 3190 1643 3196 1644
rect 3190 1642 3191 1643
rect 2977 1640 2994 1642
rect 3113 1640 3191 1642
rect 2910 1638 2916 1639
rect 2990 1639 2996 1640
rect 1926 1636 1932 1637
rect 2990 1635 2991 1639
rect 2995 1635 2996 1639
rect 3190 1639 3191 1640
rect 3195 1639 3196 1643
rect 3257 1640 3314 1642
rect 3190 1638 3196 1639
rect 2990 1634 2996 1635
rect 2110 1633 2116 1634
rect 366 1631 372 1632
rect 366 1627 367 1631
rect 371 1630 372 1631
rect 375 1631 381 1632
rect 375 1630 376 1631
rect 371 1628 376 1630
rect 371 1627 372 1628
rect 366 1626 372 1627
rect 375 1627 376 1628
rect 380 1627 381 1631
rect 375 1626 381 1627
rect 386 1631 392 1632
rect 386 1627 387 1631
rect 391 1630 392 1631
rect 607 1631 613 1632
rect 607 1630 608 1631
rect 391 1628 608 1630
rect 391 1627 392 1628
rect 386 1626 392 1627
rect 607 1627 608 1628
rect 612 1627 613 1631
rect 607 1626 613 1627
rect 750 1631 756 1632
rect 750 1627 751 1631
rect 755 1630 756 1631
rect 839 1631 845 1632
rect 839 1630 840 1631
rect 755 1628 840 1630
rect 755 1627 756 1628
rect 750 1626 756 1627
rect 839 1627 840 1628
rect 844 1627 845 1631
rect 839 1626 845 1627
rect 1055 1631 1061 1632
rect 1055 1627 1056 1631
rect 1060 1630 1061 1631
rect 1263 1631 1269 1632
rect 1060 1628 1082 1630
rect 1060 1627 1061 1628
rect 1055 1626 1061 1627
rect 471 1615 477 1616
rect 471 1611 472 1615
rect 476 1614 477 1615
rect 559 1615 565 1616
rect 559 1614 560 1615
rect 476 1612 560 1614
rect 476 1611 477 1612
rect 471 1610 477 1611
rect 559 1611 560 1612
rect 564 1611 565 1615
rect 559 1610 565 1611
rect 647 1615 653 1616
rect 647 1611 648 1615
rect 652 1614 653 1615
rect 735 1615 741 1616
rect 735 1614 736 1615
rect 652 1612 736 1614
rect 652 1611 653 1612
rect 647 1610 653 1611
rect 735 1611 736 1612
rect 740 1611 741 1615
rect 735 1610 741 1611
rect 790 1615 796 1616
rect 790 1611 791 1615
rect 795 1614 796 1615
rect 823 1615 829 1616
rect 823 1614 824 1615
rect 795 1612 824 1614
rect 795 1611 796 1612
rect 790 1610 796 1611
rect 823 1611 824 1612
rect 828 1611 829 1615
rect 823 1610 829 1611
rect 990 1615 996 1616
rect 990 1611 991 1615
rect 995 1614 996 1615
rect 1007 1615 1013 1616
rect 1007 1614 1008 1615
rect 995 1612 1008 1614
rect 995 1611 996 1612
rect 990 1610 996 1611
rect 1007 1611 1008 1612
rect 1012 1611 1013 1615
rect 1080 1614 1082 1628
rect 1263 1627 1264 1631
rect 1268 1630 1269 1631
rect 1367 1631 1373 1632
rect 1367 1630 1368 1631
rect 1268 1628 1368 1630
rect 1268 1627 1269 1628
rect 1263 1626 1269 1627
rect 1367 1627 1368 1628
rect 1372 1627 1373 1631
rect 1367 1626 1373 1627
rect 1455 1631 1461 1632
rect 1455 1627 1456 1631
rect 1460 1630 1461 1631
rect 1551 1631 1557 1632
rect 1551 1630 1552 1631
rect 1460 1628 1552 1630
rect 1460 1627 1461 1628
rect 1455 1626 1461 1627
rect 1551 1627 1552 1628
rect 1556 1627 1557 1631
rect 1551 1626 1557 1627
rect 1639 1631 1645 1632
rect 1639 1627 1640 1631
rect 1644 1630 1645 1631
rect 1727 1631 1733 1632
rect 1727 1630 1728 1631
rect 1644 1628 1728 1630
rect 1644 1627 1645 1628
rect 1639 1626 1645 1627
rect 1727 1627 1728 1628
rect 1732 1627 1733 1631
rect 1727 1626 1733 1627
rect 1815 1631 1821 1632
rect 1815 1627 1816 1631
rect 1820 1630 1821 1631
rect 1911 1631 1917 1632
rect 1911 1630 1912 1631
rect 1820 1628 1912 1630
rect 1820 1627 1821 1628
rect 1815 1626 1821 1627
rect 1911 1627 1912 1628
rect 1916 1627 1917 1631
rect 1911 1626 1917 1627
rect 1998 1631 2005 1632
rect 1998 1627 1999 1631
rect 2004 1627 2005 1631
rect 2110 1629 2111 1633
rect 2115 1629 2116 1633
rect 2110 1628 2116 1629
rect 2238 1633 2244 1634
rect 2238 1629 2239 1633
rect 2243 1629 2244 1633
rect 2238 1628 2244 1629
rect 2382 1633 2388 1634
rect 2382 1629 2383 1633
rect 2387 1629 2388 1633
rect 2382 1628 2388 1629
rect 2518 1633 2524 1634
rect 2518 1629 2519 1633
rect 2523 1629 2524 1633
rect 2518 1628 2524 1629
rect 2654 1633 2660 1634
rect 2654 1629 2655 1633
rect 2659 1629 2660 1633
rect 2654 1628 2660 1629
rect 2790 1633 2796 1634
rect 2790 1629 2791 1633
rect 2795 1629 2796 1633
rect 2790 1628 2796 1629
rect 2926 1633 2932 1634
rect 2926 1629 2927 1633
rect 2931 1629 2932 1633
rect 2926 1628 2932 1629
rect 3062 1633 3068 1634
rect 3062 1629 3063 1633
rect 3067 1629 3068 1633
rect 3062 1628 3068 1629
rect 3206 1633 3212 1634
rect 3206 1629 3207 1633
rect 3211 1629 3212 1633
rect 3206 1628 3212 1629
rect 3312 1630 3314 1640
rect 3350 1633 3356 1634
rect 3312 1628 3346 1630
rect 3350 1629 3351 1633
rect 3355 1629 3356 1633
rect 3350 1628 3356 1629
rect 1998 1626 2005 1627
rect 1430 1623 1436 1624
rect 1430 1619 1431 1623
rect 1435 1622 1436 1623
rect 2183 1623 2189 1624
rect 1435 1620 1562 1622
rect 1435 1619 1436 1620
rect 1430 1618 1436 1619
rect 1095 1615 1101 1616
rect 1095 1614 1096 1615
rect 1080 1612 1096 1614
rect 1007 1610 1013 1611
rect 1095 1611 1096 1612
rect 1100 1611 1101 1615
rect 1183 1615 1189 1616
rect 1183 1614 1184 1615
rect 1095 1610 1101 1611
rect 1104 1612 1184 1614
rect 398 1607 404 1608
rect 398 1603 399 1607
rect 403 1603 404 1607
rect 398 1602 404 1603
rect 574 1607 580 1608
rect 574 1603 575 1607
rect 579 1603 580 1607
rect 574 1602 580 1603
rect 750 1607 756 1608
rect 750 1603 751 1607
rect 755 1603 756 1607
rect 750 1602 756 1603
rect 934 1607 940 1608
rect 934 1603 935 1607
rect 939 1603 940 1607
rect 1104 1606 1106 1612
rect 1183 1611 1184 1612
rect 1188 1611 1189 1615
rect 1183 1610 1189 1611
rect 1351 1615 1357 1616
rect 1351 1611 1352 1615
rect 1356 1614 1357 1615
rect 1431 1615 1437 1616
rect 1431 1614 1432 1615
rect 1356 1612 1432 1614
rect 1356 1611 1357 1612
rect 1351 1610 1357 1611
rect 1431 1611 1432 1612
rect 1436 1611 1437 1615
rect 1431 1610 1437 1611
rect 1519 1615 1525 1616
rect 1519 1611 1520 1615
rect 1524 1614 1525 1615
rect 1550 1615 1556 1616
rect 1550 1614 1551 1615
rect 1524 1612 1551 1614
rect 1524 1611 1525 1612
rect 1519 1610 1525 1611
rect 1550 1611 1551 1612
rect 1555 1611 1556 1615
rect 1560 1614 1562 1620
rect 2183 1619 2184 1623
rect 2188 1622 2189 1623
rect 2223 1623 2229 1624
rect 2223 1622 2224 1623
rect 2188 1620 2224 1622
rect 2188 1619 2189 1620
rect 2183 1618 2189 1619
rect 2223 1619 2224 1620
rect 2228 1619 2229 1623
rect 2223 1618 2229 1619
rect 2311 1623 2317 1624
rect 2311 1619 2312 1623
rect 2316 1622 2317 1623
rect 2367 1623 2373 1624
rect 2367 1622 2368 1623
rect 2316 1620 2368 1622
rect 2316 1619 2317 1620
rect 2311 1618 2317 1619
rect 2367 1619 2368 1620
rect 2372 1619 2373 1623
rect 2367 1618 2373 1619
rect 2455 1623 2461 1624
rect 2455 1619 2456 1623
rect 2460 1622 2461 1623
rect 2486 1623 2492 1624
rect 2486 1622 2487 1623
rect 2460 1620 2487 1622
rect 2460 1619 2461 1620
rect 2455 1618 2461 1619
rect 2486 1619 2487 1620
rect 2491 1619 2492 1623
rect 2486 1618 2492 1619
rect 2591 1623 2597 1624
rect 2591 1619 2592 1623
rect 2596 1622 2597 1623
rect 2639 1623 2645 1624
rect 2639 1622 2640 1623
rect 2596 1620 2640 1622
rect 2596 1619 2597 1620
rect 2591 1618 2597 1619
rect 2639 1619 2640 1620
rect 2644 1619 2645 1623
rect 2639 1618 2645 1619
rect 2726 1623 2733 1624
rect 2726 1619 2727 1623
rect 2732 1619 2733 1623
rect 2726 1618 2733 1619
rect 2830 1623 2836 1624
rect 2830 1619 2831 1623
rect 2835 1622 2836 1623
rect 2863 1623 2869 1624
rect 2863 1622 2864 1623
rect 2835 1620 2864 1622
rect 2835 1619 2836 1620
rect 2830 1618 2836 1619
rect 2863 1619 2864 1620
rect 2868 1619 2869 1623
rect 2863 1618 2869 1619
rect 2910 1623 2916 1624
rect 2910 1619 2911 1623
rect 2915 1622 2916 1623
rect 2999 1623 3005 1624
rect 2999 1622 3000 1623
rect 2915 1620 3000 1622
rect 2915 1619 2916 1620
rect 2910 1618 2916 1619
rect 2999 1619 3000 1620
rect 3004 1619 3005 1623
rect 2999 1618 3005 1619
rect 3134 1623 3141 1624
rect 3134 1619 3135 1623
rect 3140 1619 3141 1623
rect 3134 1618 3141 1619
rect 3190 1623 3196 1624
rect 3190 1619 3191 1623
rect 3195 1622 3196 1623
rect 3279 1623 3285 1624
rect 3279 1622 3280 1623
rect 3195 1620 3280 1622
rect 3195 1619 3196 1620
rect 3190 1618 3196 1619
rect 3279 1619 3280 1620
rect 3284 1619 3285 1623
rect 3279 1618 3285 1619
rect 3330 1623 3341 1624
rect 3330 1619 3331 1623
rect 3335 1619 3336 1623
rect 3340 1619 3341 1623
rect 3344 1622 3346 1628
rect 3423 1623 3429 1624
rect 3423 1622 3424 1623
rect 3344 1620 3424 1622
rect 3330 1618 3341 1619
rect 3423 1619 3424 1620
rect 3428 1619 3429 1623
rect 3423 1618 3429 1619
rect 1679 1615 1685 1616
rect 1679 1614 1680 1615
rect 1560 1612 1680 1614
rect 1550 1610 1556 1611
rect 1679 1611 1680 1612
rect 1684 1611 1685 1615
rect 1839 1615 1845 1616
rect 1839 1614 1840 1615
rect 1679 1610 1685 1611
rect 1720 1612 1840 1614
rect 934 1602 940 1603
rect 1044 1604 1106 1606
rect 1110 1607 1116 1608
rect 558 1599 564 1600
rect 558 1598 559 1599
rect 449 1596 559 1598
rect 558 1595 559 1596
rect 563 1595 564 1599
rect 1044 1598 1046 1604
rect 1110 1603 1111 1607
rect 1115 1603 1116 1607
rect 1110 1602 1116 1603
rect 1278 1607 1284 1608
rect 1278 1603 1279 1607
rect 1283 1603 1284 1607
rect 1278 1602 1284 1603
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1603 1452 1607
rect 1446 1602 1452 1603
rect 1606 1607 1612 1608
rect 1606 1603 1607 1607
rect 1611 1603 1612 1607
rect 1606 1602 1612 1603
rect 1430 1599 1436 1600
rect 1430 1598 1431 1599
rect 985 1596 1046 1598
rect 1329 1596 1431 1598
rect 558 1594 564 1595
rect 1430 1595 1431 1596
rect 1435 1595 1436 1599
rect 1720 1598 1722 1612
rect 1839 1611 1840 1612
rect 1844 1611 1845 1615
rect 2007 1615 2013 1616
rect 2007 1614 2008 1615
rect 1839 1610 1845 1611
rect 1880 1612 2008 1614
rect 1766 1607 1772 1608
rect 1766 1603 1767 1607
rect 1771 1603 1772 1607
rect 1766 1602 1772 1603
rect 1880 1598 1882 1612
rect 2007 1611 2008 1612
rect 2012 1611 2013 1615
rect 2007 1610 2013 1611
rect 1934 1607 1940 1608
rect 1934 1603 1935 1607
rect 1939 1603 1940 1607
rect 1934 1602 1940 1603
rect 1998 1599 2004 1600
rect 1998 1598 1999 1599
rect 1657 1596 1722 1598
rect 1817 1596 1882 1598
rect 1985 1596 1999 1598
rect 1430 1594 1436 1595
rect 1998 1595 1999 1596
rect 2003 1595 2004 1599
rect 1998 1594 2004 1595
rect 2182 1599 2188 1600
rect 2182 1595 2183 1599
rect 2187 1598 2188 1599
rect 2239 1599 2245 1600
rect 2239 1598 2240 1599
rect 2187 1596 2240 1598
rect 2187 1595 2188 1596
rect 2182 1594 2188 1595
rect 2239 1595 2240 1596
rect 2244 1595 2245 1599
rect 2359 1599 2365 1600
rect 2359 1598 2360 1599
rect 2239 1594 2245 1595
rect 2260 1596 2360 1598
rect 2166 1591 2172 1592
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 110 1583 116 1584
rect 2030 1588 2036 1589
rect 2030 1584 2031 1588
rect 2035 1584 2036 1588
rect 2166 1587 2167 1591
rect 2171 1587 2172 1591
rect 2166 1586 2172 1587
rect 2030 1583 2036 1584
rect 2260 1582 2262 1596
rect 2359 1595 2360 1596
rect 2364 1595 2365 1599
rect 2479 1599 2485 1600
rect 2479 1598 2480 1599
rect 2359 1594 2365 1595
rect 2380 1596 2480 1598
rect 2286 1591 2292 1592
rect 2286 1587 2287 1591
rect 2291 1587 2292 1591
rect 2286 1586 2292 1587
rect 2380 1582 2382 1596
rect 2479 1595 2480 1596
rect 2484 1595 2485 1599
rect 2599 1599 2605 1600
rect 2599 1598 2600 1599
rect 2479 1594 2485 1595
rect 2500 1596 2600 1598
rect 2406 1591 2412 1592
rect 2406 1587 2407 1591
rect 2411 1587 2412 1591
rect 2406 1586 2412 1587
rect 2500 1582 2502 1596
rect 2599 1595 2600 1596
rect 2604 1595 2605 1599
rect 2599 1594 2605 1595
rect 2614 1599 2620 1600
rect 2614 1595 2615 1599
rect 2619 1598 2620 1599
rect 2719 1599 2725 1600
rect 2719 1598 2720 1599
rect 2619 1596 2720 1598
rect 2619 1595 2620 1596
rect 2614 1594 2620 1595
rect 2719 1595 2720 1596
rect 2724 1595 2725 1599
rect 2719 1594 2725 1595
rect 2839 1599 2845 1600
rect 2839 1595 2840 1599
rect 2844 1598 2845 1599
rect 2918 1599 2924 1600
rect 2918 1598 2919 1599
rect 2844 1596 2919 1598
rect 2844 1595 2845 1596
rect 2839 1594 2845 1595
rect 2918 1595 2919 1596
rect 2923 1595 2924 1599
rect 2918 1594 2924 1595
rect 2959 1599 2965 1600
rect 2959 1595 2960 1599
rect 2964 1598 2965 1599
rect 2991 1599 2997 1600
rect 2991 1598 2992 1599
rect 2964 1596 2992 1598
rect 2964 1595 2965 1596
rect 2959 1594 2965 1595
rect 2991 1595 2992 1596
rect 2996 1595 2997 1599
rect 2991 1594 2997 1595
rect 3079 1599 3085 1600
rect 3079 1595 3080 1599
rect 3084 1598 3085 1599
rect 3111 1599 3117 1600
rect 3111 1598 3112 1599
rect 3084 1596 3112 1598
rect 3084 1595 3085 1596
rect 3079 1594 3085 1595
rect 3111 1595 3112 1596
rect 3116 1595 3117 1599
rect 3111 1594 3117 1595
rect 3199 1599 3205 1600
rect 3199 1595 3200 1599
rect 3204 1598 3205 1599
rect 3239 1599 3245 1600
rect 3239 1598 3240 1599
rect 3204 1596 3240 1598
rect 3204 1595 3205 1596
rect 3199 1594 3205 1595
rect 3239 1595 3240 1596
rect 3244 1595 3245 1599
rect 3239 1594 3245 1595
rect 3327 1599 3336 1600
rect 3327 1595 3328 1599
rect 3335 1595 3336 1599
rect 3327 1594 3336 1595
rect 2526 1591 2532 1592
rect 2526 1587 2527 1591
rect 2531 1587 2532 1591
rect 2526 1586 2532 1587
rect 2646 1591 2652 1592
rect 2646 1587 2647 1591
rect 2651 1587 2652 1591
rect 2646 1586 2652 1587
rect 2766 1591 2772 1592
rect 2766 1587 2767 1591
rect 2771 1587 2772 1591
rect 2766 1586 2772 1587
rect 2886 1591 2892 1592
rect 2886 1587 2887 1591
rect 2891 1587 2892 1591
rect 2886 1586 2892 1587
rect 3006 1591 3012 1592
rect 3006 1587 3007 1591
rect 3011 1587 3012 1591
rect 3006 1586 3012 1587
rect 3126 1591 3132 1592
rect 3126 1587 3127 1591
rect 3131 1587 3132 1591
rect 3126 1586 3132 1587
rect 3254 1591 3260 1592
rect 3254 1587 3255 1591
rect 3259 1587 3260 1591
rect 3254 1586 3260 1587
rect 2746 1583 2752 1584
rect 2746 1582 2747 1583
rect 2217 1580 2262 1582
rect 2337 1580 2382 1582
rect 2457 1580 2502 1582
rect 2697 1580 2747 1582
rect 2534 1579 2540 1580
rect 2534 1575 2535 1579
rect 2539 1575 2540 1579
rect 2746 1579 2747 1580
rect 2751 1579 2752 1583
rect 2830 1583 2836 1584
rect 2830 1582 2831 1583
rect 2817 1580 2831 1582
rect 2746 1578 2752 1579
rect 2830 1579 2831 1580
rect 2835 1579 2836 1583
rect 2990 1583 2996 1584
rect 2990 1582 2991 1583
rect 2937 1580 2991 1582
rect 2830 1578 2836 1579
rect 2990 1579 2991 1580
rect 2995 1579 2996 1583
rect 2990 1578 2996 1579
rect 2534 1574 2540 1575
rect 2070 1572 2076 1573
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 2030 1571 2036 1572
rect 2030 1567 2031 1571
rect 2035 1567 2036 1571
rect 2070 1568 2071 1572
rect 2075 1568 2076 1572
rect 2070 1567 2076 1568
rect 3990 1572 3996 1573
rect 3990 1568 3991 1572
rect 3995 1568 3996 1572
rect 3990 1567 3996 1568
rect 110 1566 116 1567
rect 398 1566 404 1567
rect 398 1562 399 1566
rect 403 1562 404 1566
rect 398 1561 404 1562
rect 574 1566 580 1567
rect 574 1562 575 1566
rect 579 1562 580 1566
rect 574 1561 580 1562
rect 750 1566 756 1567
rect 750 1562 751 1566
rect 755 1562 756 1566
rect 750 1561 756 1562
rect 934 1566 940 1567
rect 934 1562 935 1566
rect 939 1562 940 1566
rect 934 1561 940 1562
rect 1110 1566 1116 1567
rect 1110 1562 1111 1566
rect 1115 1562 1116 1566
rect 1110 1561 1116 1562
rect 1278 1566 1284 1567
rect 1278 1562 1279 1566
rect 1283 1562 1284 1566
rect 1278 1561 1284 1562
rect 1446 1566 1452 1567
rect 1446 1562 1447 1566
rect 1451 1562 1452 1566
rect 1446 1561 1452 1562
rect 1606 1566 1612 1567
rect 1606 1562 1607 1566
rect 1611 1562 1612 1566
rect 1606 1561 1612 1562
rect 1766 1566 1772 1567
rect 1766 1562 1767 1566
rect 1771 1562 1772 1566
rect 1766 1561 1772 1562
rect 1934 1566 1940 1567
rect 2030 1566 2036 1567
rect 1934 1562 1935 1566
rect 1939 1562 1940 1566
rect 1934 1561 1940 1562
rect 2070 1555 2076 1556
rect 2070 1551 2071 1555
rect 2075 1551 2076 1555
rect 3990 1555 3996 1556
rect 3990 1551 3991 1555
rect 3995 1551 3996 1555
rect 2070 1550 2076 1551
rect 2166 1550 2172 1551
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2286 1550 2292 1551
rect 2286 1546 2287 1550
rect 2291 1546 2292 1550
rect 2286 1545 2292 1546
rect 2406 1550 2412 1551
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2526 1550 2532 1551
rect 2526 1546 2527 1550
rect 2531 1546 2532 1550
rect 2526 1545 2532 1546
rect 2646 1550 2652 1551
rect 2646 1546 2647 1550
rect 2651 1546 2652 1550
rect 2646 1545 2652 1546
rect 2766 1550 2772 1551
rect 2766 1546 2767 1550
rect 2771 1546 2772 1550
rect 2766 1545 2772 1546
rect 2886 1550 2892 1551
rect 2886 1546 2887 1550
rect 2891 1546 2892 1550
rect 2886 1545 2892 1546
rect 3006 1550 3012 1551
rect 3006 1546 3007 1550
rect 3011 1546 3012 1550
rect 3006 1545 3012 1546
rect 3126 1550 3132 1551
rect 3126 1546 3127 1550
rect 3131 1546 3132 1550
rect 3126 1545 3132 1546
rect 3254 1550 3260 1551
rect 3990 1550 3996 1551
rect 3254 1546 3255 1550
rect 3259 1546 3260 1550
rect 3254 1545 3260 1546
rect 502 1526 508 1527
rect 502 1522 503 1526
rect 507 1522 508 1526
rect 110 1521 116 1522
rect 502 1521 508 1522
rect 614 1526 620 1527
rect 614 1522 615 1526
rect 619 1522 620 1526
rect 614 1521 620 1522
rect 734 1526 740 1527
rect 734 1522 735 1526
rect 739 1522 740 1526
rect 734 1521 740 1522
rect 854 1526 860 1527
rect 854 1522 855 1526
rect 859 1522 860 1526
rect 854 1521 860 1522
rect 966 1526 972 1527
rect 966 1522 967 1526
rect 971 1522 972 1526
rect 966 1521 972 1522
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1198 1526 1204 1527
rect 1198 1522 1199 1526
rect 1203 1522 1204 1526
rect 1198 1521 1204 1522
rect 1318 1526 1324 1527
rect 1318 1522 1319 1526
rect 1323 1522 1324 1526
rect 1318 1521 1324 1522
rect 1438 1526 1444 1527
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1558 1526 1564 1527
rect 1558 1522 1559 1526
rect 1563 1522 1564 1526
rect 1558 1521 1564 1522
rect 2030 1521 2036 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 110 1516 116 1517
rect 2030 1517 2031 1521
rect 2035 1517 2036 1521
rect 2030 1516 2036 1517
rect 2350 1510 2356 1511
rect 2350 1506 2351 1510
rect 2355 1506 2356 1510
rect 2070 1505 2076 1506
rect 2350 1505 2356 1506
rect 2462 1510 2468 1511
rect 2462 1506 2463 1510
rect 2467 1506 2468 1510
rect 2462 1505 2468 1506
rect 2574 1510 2580 1511
rect 2574 1506 2575 1510
rect 2579 1506 2580 1510
rect 2574 1505 2580 1506
rect 2694 1510 2700 1511
rect 2694 1506 2695 1510
rect 2699 1506 2700 1510
rect 2694 1505 2700 1506
rect 2814 1510 2820 1511
rect 2814 1506 2815 1510
rect 2819 1506 2820 1510
rect 2814 1505 2820 1506
rect 2926 1510 2932 1511
rect 2926 1506 2927 1510
rect 2931 1506 2932 1510
rect 2926 1505 2932 1506
rect 3046 1510 3052 1511
rect 3046 1506 3047 1510
rect 3051 1506 3052 1510
rect 3046 1505 3052 1506
rect 3166 1510 3172 1511
rect 3166 1506 3167 1510
rect 3171 1506 3172 1510
rect 3166 1505 3172 1506
rect 3286 1510 3292 1511
rect 3286 1506 3287 1510
rect 3291 1506 3292 1510
rect 3286 1505 3292 1506
rect 3406 1510 3412 1511
rect 3406 1506 3407 1510
rect 3411 1506 3412 1510
rect 3406 1505 3412 1506
rect 3990 1505 3996 1506
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 110 1499 116 1500
rect 2030 1504 2036 1505
rect 2030 1500 2031 1504
rect 2035 1500 2036 1504
rect 2070 1501 2071 1505
rect 2075 1501 2076 1505
rect 2070 1500 2076 1501
rect 3990 1501 3991 1505
rect 3995 1501 3996 1505
rect 3990 1500 3996 1501
rect 2030 1499 2036 1500
rect 598 1495 604 1496
rect 598 1494 599 1495
rect 553 1492 599 1494
rect 598 1491 599 1492
rect 603 1491 604 1495
rect 718 1495 724 1496
rect 718 1494 719 1495
rect 665 1492 719 1494
rect 598 1490 604 1491
rect 718 1491 719 1492
rect 723 1491 724 1495
rect 718 1490 724 1491
rect 758 1495 764 1496
rect 758 1491 759 1495
rect 763 1491 764 1495
rect 950 1495 956 1496
rect 950 1494 951 1495
rect 905 1492 951 1494
rect 758 1490 764 1491
rect 950 1491 951 1492
rect 955 1491 956 1495
rect 950 1490 956 1491
rect 990 1495 996 1496
rect 990 1491 991 1495
rect 995 1491 996 1495
rect 1182 1495 1188 1496
rect 1182 1494 1183 1495
rect 1129 1492 1183 1494
rect 990 1490 996 1491
rect 1182 1491 1183 1492
rect 1187 1491 1188 1495
rect 1422 1495 1428 1496
rect 1422 1494 1423 1495
rect 1369 1492 1423 1494
rect 1182 1490 1188 1491
rect 1422 1491 1423 1492
rect 1427 1491 1428 1495
rect 1542 1495 1548 1496
rect 1542 1494 1543 1495
rect 1489 1492 1543 1494
rect 1422 1490 1428 1491
rect 1542 1491 1543 1492
rect 1547 1491 1548 1495
rect 1542 1490 1548 1491
rect 1550 1495 1556 1496
rect 1550 1491 1551 1495
rect 1555 1491 1556 1495
rect 1550 1490 1556 1491
rect 2070 1488 2076 1489
rect 502 1485 508 1486
rect 502 1481 503 1485
rect 507 1481 508 1485
rect 502 1480 508 1481
rect 614 1485 620 1486
rect 614 1481 615 1485
rect 619 1481 620 1485
rect 614 1480 620 1481
rect 734 1485 740 1486
rect 734 1481 735 1485
rect 739 1481 740 1485
rect 734 1480 740 1481
rect 854 1485 860 1486
rect 854 1481 855 1485
rect 859 1481 860 1485
rect 854 1480 860 1481
rect 966 1485 972 1486
rect 966 1481 967 1485
rect 971 1481 972 1485
rect 966 1480 972 1481
rect 1078 1485 1084 1486
rect 1078 1481 1079 1485
rect 1083 1481 1084 1485
rect 1078 1480 1084 1481
rect 1198 1485 1204 1486
rect 1198 1481 1199 1485
rect 1203 1481 1204 1485
rect 1198 1480 1204 1481
rect 1318 1485 1324 1486
rect 1318 1481 1319 1485
rect 1323 1481 1324 1485
rect 1318 1480 1324 1481
rect 1438 1485 1444 1486
rect 1438 1481 1439 1485
rect 1443 1481 1444 1485
rect 1438 1480 1444 1481
rect 1558 1485 1564 1486
rect 1558 1481 1559 1485
rect 1563 1481 1564 1485
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 3990 1488 3996 1489
rect 3990 1484 3991 1488
rect 3995 1484 3996 1488
rect 3990 1483 3996 1484
rect 1558 1480 1564 1481
rect 2446 1479 2452 1480
rect 2446 1478 2447 1479
rect 2401 1476 2447 1478
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1474 564 1475
rect 575 1475 581 1476
rect 575 1474 576 1475
rect 563 1472 576 1474
rect 563 1471 564 1472
rect 558 1470 564 1471
rect 575 1471 576 1472
rect 580 1471 581 1475
rect 575 1470 581 1471
rect 598 1475 604 1476
rect 598 1471 599 1475
rect 603 1474 604 1475
rect 687 1475 693 1476
rect 687 1474 688 1475
rect 603 1472 688 1474
rect 603 1471 604 1472
rect 598 1470 604 1471
rect 687 1471 688 1472
rect 692 1471 693 1475
rect 687 1470 693 1471
rect 718 1475 724 1476
rect 718 1471 719 1475
rect 723 1474 724 1475
rect 807 1475 813 1476
rect 807 1474 808 1475
rect 723 1472 808 1474
rect 723 1471 724 1472
rect 718 1470 724 1471
rect 807 1471 808 1472
rect 812 1471 813 1475
rect 807 1470 813 1471
rect 918 1475 924 1476
rect 918 1471 919 1475
rect 923 1474 924 1475
rect 927 1475 933 1476
rect 927 1474 928 1475
rect 923 1472 928 1474
rect 923 1471 924 1472
rect 918 1470 924 1471
rect 927 1471 928 1472
rect 932 1471 933 1475
rect 927 1470 933 1471
rect 950 1475 956 1476
rect 950 1471 951 1475
rect 955 1474 956 1475
rect 1039 1475 1045 1476
rect 1039 1474 1040 1475
rect 955 1472 1040 1474
rect 955 1471 956 1472
rect 950 1470 956 1471
rect 1039 1471 1040 1472
rect 1044 1471 1045 1475
rect 1039 1470 1045 1471
rect 1151 1475 1157 1476
rect 1151 1471 1152 1475
rect 1156 1474 1157 1475
rect 1183 1475 1189 1476
rect 1183 1474 1184 1475
rect 1156 1472 1184 1474
rect 1156 1471 1157 1472
rect 1151 1470 1157 1471
rect 1183 1471 1184 1472
rect 1188 1471 1189 1475
rect 1183 1470 1189 1471
rect 1270 1475 1277 1476
rect 1270 1471 1271 1475
rect 1276 1471 1277 1475
rect 1270 1470 1277 1471
rect 1391 1475 1397 1476
rect 1391 1471 1392 1475
rect 1396 1471 1397 1475
rect 1391 1470 1397 1471
rect 1422 1475 1428 1476
rect 1422 1471 1423 1475
rect 1427 1474 1428 1475
rect 1511 1475 1517 1476
rect 1511 1474 1512 1475
rect 1427 1472 1512 1474
rect 1427 1471 1428 1472
rect 1422 1470 1428 1471
rect 1511 1471 1512 1472
rect 1516 1471 1517 1475
rect 1511 1470 1517 1471
rect 1542 1475 1548 1476
rect 1542 1471 1543 1475
rect 1547 1474 1548 1475
rect 1631 1475 1637 1476
rect 1631 1474 1632 1475
rect 1547 1472 1632 1474
rect 1547 1471 1548 1472
rect 1542 1470 1548 1471
rect 1631 1471 1632 1472
rect 1636 1471 1637 1475
rect 2446 1475 2447 1476
rect 2451 1475 2452 1479
rect 2886 1479 2892 1480
rect 2886 1478 2887 1479
rect 2625 1476 2642 1478
rect 2865 1476 2887 1478
rect 2446 1474 2452 1475
rect 2638 1475 2644 1476
rect 1631 1470 1637 1471
rect 2638 1471 2639 1475
rect 2643 1471 2644 1475
rect 2886 1475 2887 1476
rect 2891 1475 2892 1479
rect 2886 1474 2892 1475
rect 2918 1479 2924 1480
rect 2918 1475 2919 1479
rect 2923 1475 2924 1479
rect 3150 1479 3156 1480
rect 3150 1478 3151 1479
rect 3097 1476 3151 1478
rect 2918 1474 2924 1475
rect 3150 1475 3151 1476
rect 3155 1475 3156 1479
rect 3270 1479 3276 1480
rect 3270 1478 3271 1479
rect 3217 1476 3271 1478
rect 3150 1474 3156 1475
rect 3270 1475 3271 1476
rect 3275 1475 3276 1479
rect 3337 1476 3398 1478
rect 3270 1474 3276 1475
rect 2638 1470 2644 1471
rect 1182 1467 1188 1468
rect 1182 1463 1183 1467
rect 1187 1466 1188 1467
rect 1393 1466 1395 1470
rect 1187 1464 1395 1466
rect 2350 1469 2356 1470
rect 2350 1465 2351 1469
rect 2355 1465 2356 1469
rect 2350 1464 2356 1465
rect 2462 1469 2468 1470
rect 2462 1465 2463 1469
rect 2467 1465 2468 1469
rect 2462 1464 2468 1465
rect 2574 1469 2580 1470
rect 2574 1465 2575 1469
rect 2579 1465 2580 1469
rect 2574 1464 2580 1465
rect 2694 1469 2700 1470
rect 2694 1465 2695 1469
rect 2699 1465 2700 1469
rect 2814 1469 2820 1470
rect 2694 1464 2700 1465
rect 2760 1464 2806 1466
rect 2814 1465 2815 1469
rect 2819 1465 2820 1469
rect 2814 1464 2820 1465
rect 2926 1469 2932 1470
rect 2926 1465 2927 1469
rect 2931 1465 2932 1469
rect 3046 1469 3052 1470
rect 2926 1464 2932 1465
rect 2990 1467 2996 1468
rect 1187 1463 1188 1464
rect 1182 1462 1188 1463
rect 2746 1463 2752 1464
rect 670 1459 676 1460
rect 670 1455 671 1459
rect 675 1458 676 1459
rect 1406 1459 1412 1460
rect 675 1456 770 1458
rect 675 1455 676 1456
rect 670 1454 676 1455
rect 655 1451 661 1452
rect 655 1447 656 1451
rect 660 1450 661 1451
rect 671 1451 677 1452
rect 671 1450 672 1451
rect 660 1448 672 1450
rect 660 1447 661 1448
rect 655 1446 661 1447
rect 671 1447 672 1448
rect 676 1447 677 1451
rect 671 1446 677 1447
rect 758 1451 765 1452
rect 758 1447 759 1451
rect 764 1447 765 1451
rect 768 1450 770 1456
rect 1406 1455 1407 1459
rect 1411 1458 1412 1459
rect 2423 1459 2429 1460
rect 1411 1456 1595 1458
rect 1411 1455 1412 1456
rect 1406 1454 1412 1455
rect 1593 1452 1595 1456
rect 2423 1455 2424 1459
rect 2428 1458 2429 1459
rect 2447 1459 2453 1460
rect 2447 1458 2448 1459
rect 2428 1456 2448 1458
rect 2428 1455 2429 1456
rect 2423 1454 2429 1455
rect 2447 1455 2448 1456
rect 2452 1455 2453 1459
rect 2447 1454 2453 1455
rect 2534 1459 2541 1460
rect 2534 1455 2535 1459
rect 2540 1455 2541 1459
rect 2534 1454 2541 1455
rect 2647 1459 2653 1460
rect 2647 1455 2648 1459
rect 2652 1458 2653 1459
rect 2679 1459 2685 1460
rect 2679 1458 2680 1459
rect 2652 1456 2680 1458
rect 2652 1455 2653 1456
rect 2647 1454 2653 1455
rect 2679 1455 2680 1456
rect 2684 1455 2685 1459
rect 2746 1459 2747 1463
rect 2751 1462 2752 1463
rect 2760 1462 2762 1464
rect 2751 1460 2762 1462
rect 2751 1459 2752 1460
rect 2746 1458 2752 1459
rect 2766 1459 2773 1460
rect 2679 1454 2685 1455
rect 2766 1455 2767 1459
rect 2772 1455 2773 1459
rect 2804 1458 2806 1464
rect 2990 1463 2991 1467
rect 2995 1466 2996 1467
rect 2995 1464 3010 1466
rect 3046 1465 3047 1469
rect 3051 1465 3052 1469
rect 3046 1464 3052 1465
rect 3166 1469 3172 1470
rect 3166 1465 3167 1469
rect 3171 1465 3172 1469
rect 3166 1464 3172 1465
rect 3286 1469 3292 1470
rect 3286 1465 3287 1469
rect 3291 1465 3292 1469
rect 3286 1464 3292 1465
rect 3396 1466 3398 1476
rect 3406 1469 3412 1470
rect 3396 1464 3402 1466
rect 3406 1465 3407 1469
rect 3411 1465 3412 1469
rect 3406 1464 3412 1465
rect 2995 1463 2996 1464
rect 2990 1462 2996 1463
rect 2887 1459 2893 1460
rect 2887 1458 2888 1459
rect 2804 1456 2888 1458
rect 2766 1454 2773 1455
rect 2887 1455 2888 1456
rect 2892 1455 2893 1459
rect 2887 1454 2893 1455
rect 2998 1459 3005 1460
rect 2998 1455 2999 1459
rect 3004 1455 3005 1459
rect 3008 1458 3010 1464
rect 3119 1459 3125 1460
rect 3119 1458 3120 1459
rect 3008 1456 3120 1458
rect 2998 1454 3005 1455
rect 3119 1455 3120 1456
rect 3124 1455 3125 1459
rect 3119 1454 3125 1455
rect 3150 1459 3156 1460
rect 3150 1455 3151 1459
rect 3155 1458 3156 1459
rect 3239 1459 3245 1460
rect 3239 1458 3240 1459
rect 3155 1456 3240 1458
rect 3155 1455 3156 1456
rect 3150 1454 3156 1455
rect 3239 1455 3240 1456
rect 3244 1455 3245 1459
rect 3239 1454 3245 1455
rect 3270 1459 3276 1460
rect 3270 1455 3271 1459
rect 3275 1458 3276 1459
rect 3359 1459 3365 1460
rect 3359 1458 3360 1459
rect 3275 1456 3360 1458
rect 3275 1455 3276 1456
rect 3270 1454 3276 1455
rect 3359 1455 3360 1456
rect 3364 1455 3365 1459
rect 3359 1454 3365 1455
rect 3378 1459 3384 1460
rect 3378 1455 3379 1459
rect 3383 1458 3384 1459
rect 3391 1459 3397 1460
rect 3391 1458 3392 1459
rect 3383 1456 3392 1458
rect 3383 1455 3384 1456
rect 3378 1454 3384 1455
rect 3391 1455 3392 1456
rect 3396 1455 3397 1459
rect 3400 1458 3402 1464
rect 3479 1459 3485 1460
rect 3479 1458 3480 1459
rect 3400 1456 3480 1458
rect 3391 1454 3397 1455
rect 3479 1455 3480 1456
rect 3484 1455 3485 1459
rect 3479 1454 3485 1455
rect 863 1451 869 1452
rect 863 1450 864 1451
rect 768 1448 864 1450
rect 758 1446 765 1447
rect 863 1447 864 1448
rect 868 1447 869 1451
rect 863 1446 869 1447
rect 967 1451 973 1452
rect 967 1447 968 1451
rect 972 1450 973 1451
rect 983 1451 989 1452
rect 983 1450 984 1451
rect 972 1448 984 1450
rect 972 1447 973 1448
rect 967 1446 973 1447
rect 983 1447 984 1448
rect 988 1447 989 1451
rect 983 1446 989 1447
rect 1071 1451 1077 1452
rect 1071 1447 1072 1451
rect 1076 1450 1077 1451
rect 1087 1451 1093 1452
rect 1087 1450 1088 1451
rect 1076 1448 1088 1450
rect 1076 1447 1077 1448
rect 1071 1446 1077 1447
rect 1087 1447 1088 1448
rect 1092 1447 1093 1451
rect 1087 1446 1093 1447
rect 1166 1451 1172 1452
rect 1166 1447 1167 1451
rect 1171 1450 1172 1451
rect 1175 1451 1181 1452
rect 1175 1450 1176 1451
rect 1171 1448 1176 1450
rect 1171 1447 1172 1448
rect 1166 1446 1172 1447
rect 1175 1447 1176 1448
rect 1180 1447 1181 1451
rect 1175 1446 1181 1447
rect 1279 1451 1285 1452
rect 1279 1447 1280 1451
rect 1284 1450 1285 1451
rect 1295 1451 1301 1452
rect 1295 1450 1296 1451
rect 1284 1448 1296 1450
rect 1284 1447 1285 1448
rect 1279 1446 1285 1447
rect 1295 1447 1296 1448
rect 1300 1447 1301 1451
rect 1295 1446 1301 1447
rect 1383 1451 1389 1452
rect 1383 1447 1384 1451
rect 1388 1450 1389 1451
rect 1399 1451 1405 1452
rect 1399 1450 1400 1451
rect 1388 1448 1400 1450
rect 1388 1447 1389 1448
rect 1383 1446 1389 1447
rect 1399 1447 1400 1448
rect 1404 1447 1405 1451
rect 1399 1446 1405 1447
rect 1487 1451 1493 1452
rect 1487 1447 1488 1451
rect 1492 1450 1493 1451
rect 1503 1451 1509 1452
rect 1503 1450 1504 1451
rect 1492 1448 1504 1450
rect 1492 1447 1493 1448
rect 1487 1446 1493 1447
rect 1503 1447 1504 1448
rect 1508 1447 1509 1451
rect 1503 1446 1509 1447
rect 1591 1451 1597 1452
rect 1591 1447 1592 1451
rect 1596 1447 1597 1451
rect 1591 1446 1597 1447
rect 582 1443 588 1444
rect 582 1439 583 1443
rect 587 1439 588 1443
rect 582 1438 588 1439
rect 686 1443 692 1444
rect 686 1439 687 1443
rect 691 1439 692 1443
rect 686 1438 692 1439
rect 790 1443 796 1444
rect 790 1439 791 1443
rect 795 1439 796 1443
rect 790 1438 796 1439
rect 894 1443 900 1444
rect 894 1439 895 1443
rect 899 1439 900 1443
rect 894 1438 900 1439
rect 998 1443 1004 1444
rect 998 1439 999 1443
rect 1003 1439 1004 1443
rect 998 1438 1004 1439
rect 1102 1443 1108 1444
rect 1102 1439 1103 1443
rect 1107 1439 1108 1443
rect 1102 1438 1108 1439
rect 1206 1443 1212 1444
rect 1206 1439 1207 1443
rect 1211 1439 1212 1443
rect 1206 1438 1212 1439
rect 1310 1443 1316 1444
rect 1310 1439 1311 1443
rect 1315 1439 1316 1443
rect 1310 1438 1316 1439
rect 1414 1443 1420 1444
rect 1414 1439 1415 1443
rect 1419 1439 1420 1443
rect 1414 1438 1420 1439
rect 1518 1443 1524 1444
rect 1518 1439 1519 1443
rect 1523 1439 1524 1443
rect 1518 1438 1524 1439
rect 670 1435 676 1436
rect 670 1434 671 1435
rect 633 1432 671 1434
rect 670 1431 671 1432
rect 675 1431 676 1435
rect 854 1435 860 1436
rect 854 1434 855 1435
rect 841 1432 855 1434
rect 670 1430 676 1431
rect 854 1431 855 1432
rect 859 1431 860 1435
rect 1270 1435 1276 1436
rect 1270 1434 1271 1435
rect 1257 1432 1271 1434
rect 854 1430 860 1431
rect 918 1431 924 1432
rect 918 1427 919 1431
rect 923 1427 924 1431
rect 1270 1431 1271 1432
rect 1275 1431 1276 1435
rect 1270 1430 1276 1431
rect 2415 1435 2421 1436
rect 2415 1431 2416 1435
rect 2420 1434 2421 1435
rect 2431 1435 2437 1436
rect 2431 1434 2432 1435
rect 2420 1432 2432 1434
rect 2420 1431 2421 1432
rect 2415 1430 2421 1431
rect 2431 1431 2432 1432
rect 2436 1431 2437 1435
rect 2431 1430 2437 1431
rect 2519 1435 2525 1436
rect 2519 1431 2520 1435
rect 2524 1434 2525 1435
rect 2551 1435 2557 1436
rect 2551 1434 2552 1435
rect 2524 1432 2552 1434
rect 2524 1431 2525 1432
rect 2519 1430 2525 1431
rect 2551 1431 2552 1432
rect 2556 1431 2557 1435
rect 2551 1430 2557 1431
rect 2638 1435 2645 1436
rect 2638 1431 2639 1435
rect 2644 1431 2645 1435
rect 2638 1430 2645 1431
rect 2767 1435 2773 1436
rect 2767 1431 2768 1435
rect 2772 1434 2773 1435
rect 2823 1435 2829 1436
rect 2823 1434 2824 1435
rect 2772 1432 2824 1434
rect 2772 1431 2773 1432
rect 2767 1430 2773 1431
rect 2823 1431 2824 1432
rect 2828 1431 2829 1435
rect 2823 1430 2829 1431
rect 2886 1435 2892 1436
rect 2886 1431 2887 1435
rect 2891 1434 2892 1435
rect 2911 1435 2917 1436
rect 2911 1434 2912 1435
rect 2891 1432 2912 1434
rect 2891 1431 2892 1432
rect 2886 1430 2892 1431
rect 2911 1431 2912 1432
rect 2916 1431 2917 1435
rect 2911 1430 2917 1431
rect 3063 1435 3069 1436
rect 3063 1431 3064 1435
rect 3068 1434 3069 1435
rect 3127 1435 3133 1436
rect 3127 1434 3128 1435
rect 3068 1432 3128 1434
rect 3068 1431 3069 1432
rect 3063 1430 3069 1431
rect 3127 1431 3128 1432
rect 3132 1431 3133 1435
rect 3127 1430 3133 1431
rect 3206 1435 3212 1436
rect 3206 1431 3207 1435
rect 3211 1434 3212 1435
rect 3215 1435 3221 1436
rect 3215 1434 3216 1435
rect 3211 1432 3216 1434
rect 3211 1431 3212 1432
rect 3206 1430 3212 1431
rect 3215 1431 3216 1432
rect 3220 1431 3221 1435
rect 3215 1430 3221 1431
rect 3375 1435 3384 1436
rect 3375 1431 3376 1435
rect 3383 1431 3384 1435
rect 3543 1435 3549 1436
rect 3543 1434 3544 1435
rect 3375 1430 3384 1431
rect 3420 1432 3544 1434
rect 918 1426 924 1427
rect 2342 1427 2348 1428
rect 110 1424 116 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 2030 1424 2036 1425
rect 2030 1420 2031 1424
rect 2035 1420 2036 1424
rect 2342 1423 2343 1427
rect 2347 1423 2348 1427
rect 2342 1422 2348 1423
rect 2446 1427 2452 1428
rect 2446 1423 2447 1427
rect 2451 1423 2452 1427
rect 2446 1422 2452 1423
rect 2566 1427 2572 1428
rect 2566 1423 2567 1427
rect 2571 1423 2572 1427
rect 2566 1422 2572 1423
rect 2694 1427 2700 1428
rect 2694 1423 2695 1427
rect 2699 1423 2700 1427
rect 2694 1422 2700 1423
rect 2838 1427 2844 1428
rect 2838 1423 2839 1427
rect 2843 1423 2844 1427
rect 2838 1422 2844 1423
rect 2990 1427 2996 1428
rect 2990 1423 2991 1427
rect 2995 1423 2996 1427
rect 2990 1422 2996 1423
rect 3142 1427 3148 1428
rect 3142 1423 3143 1427
rect 3147 1423 3148 1427
rect 3142 1422 3148 1423
rect 3302 1427 3308 1428
rect 3302 1423 3303 1427
rect 3307 1423 3308 1427
rect 3302 1422 3308 1423
rect 2030 1419 2036 1420
rect 2766 1419 2772 1420
rect 2766 1418 2767 1419
rect 2745 1416 2767 1418
rect 2358 1415 2364 1416
rect 2358 1411 2359 1415
rect 2363 1411 2364 1415
rect 2766 1415 2767 1416
rect 2771 1415 2772 1419
rect 3420 1418 3422 1432
rect 3543 1431 3544 1432
rect 3548 1431 3549 1435
rect 3719 1435 3725 1436
rect 3719 1434 3720 1435
rect 3543 1430 3549 1431
rect 3572 1432 3720 1434
rect 3470 1427 3476 1428
rect 3470 1423 3471 1427
rect 3475 1423 3476 1427
rect 3470 1422 3476 1423
rect 3572 1418 3574 1432
rect 3719 1431 3720 1432
rect 3724 1431 3725 1435
rect 3719 1430 3725 1431
rect 3814 1435 3820 1436
rect 3814 1431 3815 1435
rect 3819 1434 3820 1435
rect 3895 1435 3901 1436
rect 3895 1434 3896 1435
rect 3819 1432 3896 1434
rect 3819 1431 3820 1432
rect 3814 1430 3820 1431
rect 3895 1431 3896 1432
rect 3900 1431 3901 1435
rect 3895 1430 3901 1431
rect 3646 1427 3652 1428
rect 3646 1423 3647 1427
rect 3651 1423 3652 1427
rect 3646 1422 3652 1423
rect 3822 1427 3828 1428
rect 3822 1423 3823 1427
rect 3827 1423 3828 1427
rect 3822 1422 3828 1423
rect 3730 1419 3736 1420
rect 3730 1418 3731 1419
rect 3353 1416 3422 1418
rect 3521 1416 3574 1418
rect 3697 1416 3731 1418
rect 2766 1414 2772 1415
rect 2998 1415 3004 1416
rect 2358 1410 2364 1411
rect 2998 1411 2999 1415
rect 3003 1411 3004 1415
rect 3730 1415 3731 1416
rect 3735 1415 3736 1419
rect 3918 1419 3924 1420
rect 3918 1418 3919 1419
rect 3873 1416 3919 1418
rect 3730 1414 3736 1415
rect 3918 1415 3919 1416
rect 3923 1415 3924 1419
rect 3918 1414 3924 1415
rect 2998 1410 3004 1411
rect 2070 1408 2076 1409
rect 110 1407 116 1408
rect 110 1403 111 1407
rect 115 1403 116 1407
rect 2030 1407 2036 1408
rect 2030 1403 2031 1407
rect 2035 1403 2036 1407
rect 2070 1404 2071 1408
rect 2075 1404 2076 1408
rect 2070 1403 2076 1404
rect 3990 1408 3996 1409
rect 3990 1404 3991 1408
rect 3995 1404 3996 1408
rect 3990 1403 3996 1404
rect 110 1402 116 1403
rect 582 1402 588 1403
rect 582 1398 583 1402
rect 587 1398 588 1402
rect 582 1397 588 1398
rect 686 1402 692 1403
rect 686 1398 687 1402
rect 691 1398 692 1402
rect 686 1397 692 1398
rect 790 1402 796 1403
rect 790 1398 791 1402
rect 795 1398 796 1402
rect 790 1397 796 1398
rect 894 1402 900 1403
rect 894 1398 895 1402
rect 899 1398 900 1402
rect 894 1397 900 1398
rect 998 1402 1004 1403
rect 998 1398 999 1402
rect 1003 1398 1004 1402
rect 998 1397 1004 1398
rect 1102 1402 1108 1403
rect 1102 1398 1103 1402
rect 1107 1398 1108 1402
rect 1102 1397 1108 1398
rect 1206 1402 1212 1403
rect 1206 1398 1207 1402
rect 1211 1398 1212 1402
rect 1206 1397 1212 1398
rect 1310 1402 1316 1403
rect 1310 1398 1311 1402
rect 1315 1398 1316 1402
rect 1310 1397 1316 1398
rect 1414 1402 1420 1403
rect 1414 1398 1415 1402
rect 1419 1398 1420 1402
rect 1414 1397 1420 1398
rect 1518 1402 1524 1403
rect 2030 1402 2036 1403
rect 1518 1398 1519 1402
rect 1523 1398 1524 1402
rect 1518 1397 1524 1398
rect 2070 1391 2076 1392
rect 2070 1387 2071 1391
rect 2075 1387 2076 1391
rect 3990 1391 3996 1392
rect 3990 1387 3991 1391
rect 3995 1387 3996 1391
rect 2070 1386 2076 1387
rect 2342 1386 2348 1387
rect 2342 1382 2343 1386
rect 2347 1382 2348 1386
rect 2342 1381 2348 1382
rect 2446 1386 2452 1387
rect 2446 1382 2447 1386
rect 2451 1382 2452 1386
rect 2446 1381 2452 1382
rect 2566 1386 2572 1387
rect 2566 1382 2567 1386
rect 2571 1382 2572 1386
rect 2566 1381 2572 1382
rect 2694 1386 2700 1387
rect 2694 1382 2695 1386
rect 2699 1382 2700 1386
rect 2694 1381 2700 1382
rect 2838 1386 2844 1387
rect 2838 1382 2839 1386
rect 2843 1382 2844 1386
rect 2838 1381 2844 1382
rect 2990 1386 2996 1387
rect 2990 1382 2991 1386
rect 2995 1382 2996 1386
rect 2990 1381 2996 1382
rect 3142 1386 3148 1387
rect 3142 1382 3143 1386
rect 3147 1382 3148 1386
rect 3142 1381 3148 1382
rect 3302 1386 3308 1387
rect 3302 1382 3303 1386
rect 3307 1382 3308 1386
rect 3302 1381 3308 1382
rect 3470 1386 3476 1387
rect 3470 1382 3471 1386
rect 3475 1382 3476 1386
rect 3470 1381 3476 1382
rect 3646 1386 3652 1387
rect 3646 1382 3647 1386
rect 3651 1382 3652 1386
rect 3646 1381 3652 1382
rect 3822 1386 3828 1387
rect 3990 1386 3996 1387
rect 3822 1382 3823 1386
rect 3827 1382 3828 1386
rect 3822 1381 3828 1382
rect 550 1362 556 1363
rect 550 1358 551 1362
rect 555 1358 556 1362
rect 110 1357 116 1358
rect 550 1357 556 1358
rect 654 1362 660 1363
rect 654 1358 655 1362
rect 659 1358 660 1362
rect 654 1357 660 1358
rect 758 1362 764 1363
rect 758 1358 759 1362
rect 763 1358 764 1362
rect 758 1357 764 1358
rect 862 1362 868 1363
rect 862 1358 863 1362
rect 867 1358 868 1362
rect 862 1357 868 1358
rect 974 1362 980 1363
rect 974 1358 975 1362
rect 979 1358 980 1362
rect 974 1357 980 1358
rect 1086 1362 1092 1363
rect 1086 1358 1087 1362
rect 1091 1358 1092 1362
rect 1086 1357 1092 1358
rect 1198 1362 1204 1363
rect 1198 1358 1199 1362
rect 1203 1358 1204 1362
rect 1198 1357 1204 1358
rect 1310 1362 1316 1363
rect 1310 1358 1311 1362
rect 1315 1358 1316 1362
rect 1310 1357 1316 1358
rect 1430 1362 1436 1363
rect 1430 1358 1431 1362
rect 1435 1358 1436 1362
rect 1430 1357 1436 1358
rect 1550 1362 1556 1363
rect 1550 1358 1551 1362
rect 1555 1358 1556 1362
rect 1550 1357 1556 1358
rect 2030 1357 2036 1358
rect 110 1353 111 1357
rect 115 1353 116 1357
rect 110 1352 116 1353
rect 2030 1353 2031 1357
rect 2035 1353 2036 1357
rect 2030 1352 2036 1353
rect 2286 1346 2292 1347
rect 2286 1342 2287 1346
rect 2291 1342 2292 1346
rect 2070 1341 2076 1342
rect 2286 1341 2292 1342
rect 2406 1346 2412 1347
rect 2406 1342 2407 1346
rect 2411 1342 2412 1346
rect 2406 1341 2412 1342
rect 2542 1346 2548 1347
rect 2542 1342 2543 1346
rect 2547 1342 2548 1346
rect 2542 1341 2548 1342
rect 2694 1346 2700 1347
rect 2694 1342 2695 1346
rect 2699 1342 2700 1346
rect 2694 1341 2700 1342
rect 2854 1346 2860 1347
rect 2854 1342 2855 1346
rect 2859 1342 2860 1346
rect 2854 1341 2860 1342
rect 3014 1346 3020 1347
rect 3014 1342 3015 1346
rect 3019 1342 3020 1346
rect 3014 1341 3020 1342
rect 3182 1346 3188 1347
rect 3182 1342 3183 1346
rect 3187 1342 3188 1346
rect 3182 1341 3188 1342
rect 3350 1346 3356 1347
rect 3350 1342 3351 1346
rect 3355 1342 3356 1346
rect 3350 1341 3356 1342
rect 3518 1346 3524 1347
rect 3518 1342 3519 1346
rect 3523 1342 3524 1346
rect 3518 1341 3524 1342
rect 3686 1346 3692 1347
rect 3686 1342 3687 1346
rect 3691 1342 3692 1346
rect 3686 1341 3692 1342
rect 3854 1346 3860 1347
rect 3854 1342 3855 1346
rect 3859 1342 3860 1346
rect 3854 1341 3860 1342
rect 3990 1341 3996 1342
rect 110 1340 116 1341
rect 110 1336 111 1340
rect 115 1336 116 1340
rect 110 1335 116 1336
rect 2030 1340 2036 1341
rect 2030 1336 2031 1340
rect 2035 1336 2036 1340
rect 2070 1337 2071 1341
rect 2075 1337 2076 1341
rect 2070 1336 2076 1337
rect 3990 1337 3991 1341
rect 3995 1337 3996 1341
rect 3990 1336 3996 1337
rect 2030 1335 2036 1336
rect 638 1331 644 1332
rect 638 1330 639 1331
rect 601 1328 639 1330
rect 638 1327 639 1328
rect 643 1327 644 1331
rect 1166 1331 1172 1332
rect 1166 1330 1167 1331
rect 1137 1328 1167 1330
rect 638 1326 644 1327
rect 1166 1327 1167 1328
rect 1171 1327 1172 1331
rect 1406 1331 1412 1332
rect 1406 1330 1407 1331
rect 1361 1328 1407 1330
rect 1166 1326 1172 1327
rect 1406 1327 1407 1328
rect 1411 1327 1412 1331
rect 1406 1326 1412 1327
rect 2070 1324 2076 1325
rect 550 1321 556 1322
rect 550 1317 551 1321
rect 555 1317 556 1321
rect 550 1316 556 1317
rect 654 1321 660 1322
rect 654 1317 655 1321
rect 659 1317 660 1321
rect 654 1316 660 1317
rect 758 1321 764 1322
rect 758 1317 759 1321
rect 763 1317 764 1321
rect 758 1316 764 1317
rect 862 1321 868 1322
rect 862 1317 863 1321
rect 867 1317 868 1321
rect 862 1316 868 1317
rect 974 1321 980 1322
rect 974 1317 975 1321
rect 979 1317 980 1321
rect 974 1316 980 1317
rect 1086 1321 1092 1322
rect 1086 1317 1087 1321
rect 1091 1317 1092 1321
rect 1086 1316 1092 1317
rect 1198 1321 1204 1322
rect 1198 1317 1199 1321
rect 1203 1317 1204 1321
rect 1198 1316 1204 1317
rect 1310 1321 1316 1322
rect 1310 1317 1311 1321
rect 1315 1317 1316 1321
rect 1310 1316 1316 1317
rect 1430 1321 1436 1322
rect 1430 1317 1431 1321
rect 1435 1317 1436 1321
rect 1430 1316 1436 1317
rect 1550 1321 1556 1322
rect 1550 1317 1551 1321
rect 1555 1317 1556 1321
rect 2070 1320 2071 1324
rect 2075 1320 2076 1324
rect 2070 1319 2076 1320
rect 3990 1324 3996 1325
rect 3990 1320 3991 1324
rect 3995 1320 3996 1324
rect 3990 1319 3996 1320
rect 1550 1316 1556 1317
rect 2390 1315 2396 1316
rect 2390 1314 2391 1315
rect 2337 1312 2391 1314
rect 623 1311 629 1312
rect 623 1307 624 1311
rect 628 1310 629 1311
rect 639 1311 645 1312
rect 639 1310 640 1311
rect 628 1308 640 1310
rect 628 1307 629 1308
rect 623 1306 629 1307
rect 639 1307 640 1308
rect 644 1307 645 1311
rect 639 1306 645 1307
rect 727 1311 733 1312
rect 727 1307 728 1311
rect 732 1310 733 1311
rect 743 1311 749 1312
rect 743 1310 744 1311
rect 732 1308 744 1310
rect 732 1307 733 1308
rect 727 1306 733 1307
rect 743 1307 744 1308
rect 748 1307 749 1311
rect 743 1306 749 1307
rect 831 1311 837 1312
rect 831 1307 832 1311
rect 836 1310 837 1311
rect 847 1311 853 1312
rect 847 1310 848 1311
rect 836 1308 848 1310
rect 836 1307 837 1308
rect 831 1306 837 1307
rect 847 1307 848 1308
rect 852 1307 853 1311
rect 847 1306 853 1307
rect 935 1311 941 1312
rect 935 1307 936 1311
rect 940 1310 941 1311
rect 959 1311 965 1312
rect 959 1310 960 1311
rect 940 1308 960 1310
rect 940 1307 941 1308
rect 935 1306 941 1307
rect 959 1307 960 1308
rect 964 1307 965 1311
rect 1047 1311 1053 1312
rect 1047 1310 1048 1311
rect 959 1306 965 1307
rect 968 1308 1048 1310
rect 638 1303 644 1304
rect 638 1299 639 1303
rect 643 1302 644 1303
rect 854 1303 860 1304
rect 643 1300 806 1302
rect 643 1299 644 1300
rect 638 1298 644 1299
rect 415 1295 421 1296
rect 415 1291 416 1295
rect 420 1294 421 1295
rect 447 1295 453 1296
rect 447 1294 448 1295
rect 420 1292 448 1294
rect 420 1291 421 1292
rect 415 1290 421 1291
rect 447 1291 448 1292
rect 452 1291 453 1295
rect 447 1290 453 1291
rect 535 1295 541 1296
rect 535 1291 536 1295
rect 540 1294 541 1295
rect 583 1295 589 1296
rect 583 1294 584 1295
rect 540 1292 584 1294
rect 540 1291 541 1292
rect 535 1290 541 1291
rect 583 1291 584 1292
rect 588 1291 589 1295
rect 583 1290 589 1291
rect 671 1295 677 1296
rect 671 1291 672 1295
rect 676 1294 677 1295
rect 727 1295 733 1296
rect 727 1294 728 1295
rect 676 1292 728 1294
rect 676 1291 677 1292
rect 671 1290 677 1291
rect 727 1291 728 1292
rect 732 1291 733 1295
rect 727 1290 733 1291
rect 342 1287 348 1288
rect 342 1283 343 1287
rect 347 1283 348 1287
rect 342 1282 348 1283
rect 462 1287 468 1288
rect 462 1283 463 1287
rect 467 1283 468 1287
rect 462 1282 468 1283
rect 598 1287 604 1288
rect 598 1283 599 1287
rect 603 1283 604 1287
rect 598 1282 604 1283
rect 742 1287 748 1288
rect 742 1283 743 1287
rect 747 1283 748 1287
rect 804 1286 806 1300
rect 854 1299 855 1303
rect 859 1302 860 1303
rect 968 1302 970 1308
rect 1047 1307 1048 1308
rect 1052 1307 1053 1311
rect 1047 1306 1053 1307
rect 1159 1311 1165 1312
rect 1159 1307 1160 1311
rect 1164 1310 1165 1311
rect 1183 1311 1189 1312
rect 1183 1310 1184 1311
rect 1164 1308 1184 1310
rect 1164 1307 1165 1308
rect 1159 1306 1165 1307
rect 1183 1307 1184 1308
rect 1188 1307 1189 1311
rect 1183 1306 1189 1307
rect 1254 1311 1260 1312
rect 1254 1307 1255 1311
rect 1259 1310 1260 1311
rect 1271 1311 1277 1312
rect 1271 1310 1272 1311
rect 1259 1308 1272 1310
rect 1259 1307 1260 1308
rect 1254 1306 1260 1307
rect 1271 1307 1272 1308
rect 1276 1307 1277 1311
rect 1271 1306 1277 1307
rect 1383 1311 1389 1312
rect 1383 1307 1384 1311
rect 1388 1310 1389 1311
rect 1415 1311 1421 1312
rect 1415 1310 1416 1311
rect 1388 1308 1416 1310
rect 1388 1307 1389 1308
rect 1383 1306 1389 1307
rect 1415 1307 1416 1308
rect 1420 1307 1421 1311
rect 1415 1306 1421 1307
rect 1503 1311 1509 1312
rect 1503 1307 1504 1311
rect 1508 1310 1509 1311
rect 1535 1311 1541 1312
rect 1535 1310 1536 1311
rect 1508 1308 1536 1310
rect 1508 1307 1509 1308
rect 1503 1306 1509 1307
rect 1535 1307 1536 1308
rect 1540 1307 1541 1311
rect 1535 1306 1541 1307
rect 1606 1311 1612 1312
rect 1606 1307 1607 1311
rect 1611 1310 1612 1311
rect 1623 1311 1629 1312
rect 1623 1310 1624 1311
rect 1611 1308 1624 1310
rect 1611 1307 1612 1308
rect 1606 1306 1612 1307
rect 1623 1307 1624 1308
rect 1628 1307 1629 1311
rect 2390 1311 2391 1312
rect 2395 1311 2396 1315
rect 2526 1315 2532 1316
rect 2526 1314 2527 1315
rect 2457 1312 2527 1314
rect 2390 1310 2396 1311
rect 2526 1311 2527 1312
rect 2531 1311 2532 1315
rect 2671 1315 2677 1316
rect 2671 1314 2672 1315
rect 2593 1312 2672 1314
rect 2526 1310 2532 1311
rect 2671 1311 2672 1312
rect 2676 1311 2677 1315
rect 2838 1315 2844 1316
rect 2838 1314 2839 1315
rect 2745 1312 2839 1314
rect 2671 1310 2677 1311
rect 2838 1311 2839 1312
rect 2843 1311 2844 1315
rect 2926 1315 2932 1316
rect 2926 1314 2927 1315
rect 2905 1312 2927 1314
rect 2838 1310 2844 1311
rect 2926 1311 2927 1312
rect 2931 1311 2932 1315
rect 3166 1315 3172 1316
rect 3166 1314 3167 1315
rect 3065 1312 3167 1314
rect 2926 1310 2932 1311
rect 3166 1311 3167 1312
rect 3171 1311 3172 1315
rect 3166 1310 3172 1311
rect 3206 1315 3212 1316
rect 3206 1311 3207 1315
rect 3211 1311 3212 1315
rect 3926 1315 3932 1316
rect 3926 1314 3927 1315
rect 3905 1312 3927 1314
rect 3206 1310 3212 1311
rect 3926 1311 3927 1312
rect 3931 1311 3932 1315
rect 3926 1310 3932 1311
rect 1623 1306 1629 1307
rect 859 1300 970 1302
rect 2286 1305 2292 1306
rect 2286 1301 2287 1305
rect 2291 1301 2292 1305
rect 2286 1300 2292 1301
rect 2406 1305 2412 1306
rect 2406 1301 2407 1305
rect 2411 1301 2412 1305
rect 2406 1300 2412 1301
rect 2542 1305 2548 1306
rect 2542 1301 2543 1305
rect 2547 1301 2548 1305
rect 2542 1300 2548 1301
rect 2694 1305 2700 1306
rect 2694 1301 2695 1305
rect 2699 1301 2700 1305
rect 2694 1300 2700 1301
rect 2854 1305 2860 1306
rect 2854 1301 2855 1305
rect 2859 1301 2860 1305
rect 2854 1300 2860 1301
rect 3014 1305 3020 1306
rect 3014 1301 3015 1305
rect 3019 1301 3020 1305
rect 3014 1300 3020 1301
rect 3182 1305 3188 1306
rect 3182 1301 3183 1305
rect 3187 1301 3188 1305
rect 3182 1300 3188 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3518 1305 3524 1306
rect 3518 1301 3519 1305
rect 3523 1301 3524 1305
rect 3518 1300 3524 1301
rect 3686 1305 3692 1306
rect 3686 1301 3687 1305
rect 3691 1301 3692 1305
rect 3686 1300 3692 1301
rect 3854 1305 3860 1306
rect 3854 1301 3855 1305
rect 3859 1301 3860 1305
rect 3854 1300 3860 1301
rect 859 1299 860 1300
rect 854 1298 860 1299
rect 815 1295 821 1296
rect 815 1291 816 1295
rect 820 1294 821 1295
rect 887 1295 893 1296
rect 887 1294 888 1295
rect 820 1292 888 1294
rect 820 1291 821 1292
rect 815 1290 821 1291
rect 887 1291 888 1292
rect 892 1291 893 1295
rect 975 1295 981 1296
rect 975 1294 976 1295
rect 887 1290 893 1291
rect 896 1292 976 1294
rect 896 1286 898 1292
rect 975 1291 976 1292
rect 980 1291 981 1295
rect 975 1290 981 1291
rect 1126 1295 1132 1296
rect 1126 1291 1127 1295
rect 1131 1294 1132 1295
rect 1135 1295 1141 1296
rect 1135 1294 1136 1295
rect 1131 1292 1136 1294
rect 1131 1291 1132 1292
rect 1126 1290 1132 1291
rect 1135 1291 1136 1292
rect 1140 1291 1141 1295
rect 1303 1295 1309 1296
rect 1303 1294 1304 1295
rect 1135 1290 1141 1291
rect 1159 1292 1304 1294
rect 804 1284 898 1286
rect 902 1287 908 1288
rect 742 1282 748 1283
rect 902 1283 903 1287
rect 907 1283 908 1287
rect 902 1282 908 1283
rect 1062 1287 1068 1288
rect 1062 1283 1063 1287
rect 1067 1283 1068 1287
rect 1062 1282 1068 1283
rect 446 1279 452 1280
rect 446 1278 447 1279
rect 393 1276 447 1278
rect 446 1275 447 1276
rect 451 1275 452 1279
rect 1159 1278 1161 1292
rect 1303 1291 1304 1292
rect 1308 1291 1309 1295
rect 1303 1290 1309 1291
rect 1414 1295 1420 1296
rect 1414 1291 1415 1295
rect 1419 1294 1420 1295
rect 1479 1295 1485 1296
rect 1479 1294 1480 1295
rect 1419 1292 1480 1294
rect 1419 1291 1420 1292
rect 1414 1290 1420 1291
rect 1479 1291 1480 1292
rect 1484 1291 1485 1295
rect 1655 1295 1661 1296
rect 1655 1294 1656 1295
rect 1479 1290 1485 1291
rect 1528 1292 1656 1294
rect 1230 1287 1236 1288
rect 1230 1283 1231 1287
rect 1235 1283 1236 1287
rect 1230 1282 1236 1283
rect 1406 1287 1412 1288
rect 1406 1283 1407 1287
rect 1411 1283 1412 1287
rect 1406 1282 1412 1283
rect 1528 1278 1530 1292
rect 1655 1291 1656 1292
rect 1660 1291 1661 1295
rect 1655 1290 1661 1291
rect 2358 1295 2365 1296
rect 2358 1291 2359 1295
rect 2364 1291 2365 1295
rect 2358 1290 2365 1291
rect 2390 1295 2396 1296
rect 2390 1291 2391 1295
rect 2395 1294 2396 1295
rect 2479 1295 2485 1296
rect 2479 1294 2480 1295
rect 2395 1292 2480 1294
rect 2395 1291 2396 1292
rect 2390 1290 2396 1291
rect 2479 1291 2480 1292
rect 2484 1291 2485 1295
rect 2479 1290 2485 1291
rect 2526 1295 2532 1296
rect 2526 1291 2527 1295
rect 2531 1294 2532 1295
rect 2615 1295 2621 1296
rect 2615 1294 2616 1295
rect 2531 1292 2616 1294
rect 2531 1291 2532 1292
rect 2526 1290 2532 1291
rect 2615 1291 2616 1292
rect 2620 1291 2621 1295
rect 2615 1290 2621 1291
rect 2766 1295 2773 1296
rect 2766 1291 2767 1295
rect 2772 1291 2773 1295
rect 2766 1290 2773 1291
rect 2838 1295 2844 1296
rect 2838 1291 2839 1295
rect 2843 1294 2844 1295
rect 2927 1295 2933 1296
rect 2927 1294 2928 1295
rect 2843 1292 2928 1294
rect 2843 1291 2844 1292
rect 2838 1290 2844 1291
rect 2927 1291 2928 1292
rect 2932 1291 2933 1295
rect 2927 1290 2933 1291
rect 3086 1295 3093 1296
rect 3086 1291 3087 1295
rect 3092 1291 3093 1295
rect 3086 1290 3093 1291
rect 3166 1295 3172 1296
rect 3166 1291 3167 1295
rect 3171 1294 3172 1295
rect 3255 1295 3261 1296
rect 3255 1294 3256 1295
rect 3171 1292 3256 1294
rect 3171 1291 3172 1292
rect 3166 1290 3172 1291
rect 3255 1291 3256 1292
rect 3260 1291 3261 1295
rect 3255 1290 3261 1291
rect 3322 1295 3328 1296
rect 3322 1291 3323 1295
rect 3327 1294 3328 1295
rect 3335 1295 3341 1296
rect 3335 1294 3336 1295
rect 3327 1292 3336 1294
rect 3327 1291 3328 1292
rect 3322 1290 3328 1291
rect 3335 1291 3336 1292
rect 3340 1291 3341 1295
rect 3335 1290 3341 1291
rect 3423 1295 3429 1296
rect 3423 1291 3424 1295
rect 3428 1294 3429 1295
rect 3503 1295 3509 1296
rect 3503 1294 3504 1295
rect 3428 1292 3504 1294
rect 3428 1291 3429 1292
rect 3423 1290 3429 1291
rect 3503 1291 3504 1292
rect 3508 1291 3509 1295
rect 3503 1290 3509 1291
rect 3591 1295 3597 1296
rect 3591 1291 3592 1295
rect 3596 1294 3597 1295
rect 3671 1295 3677 1296
rect 3671 1294 3672 1295
rect 3596 1292 3672 1294
rect 3596 1291 3597 1292
rect 3591 1290 3597 1291
rect 3671 1291 3672 1292
rect 3676 1291 3677 1295
rect 3671 1290 3677 1291
rect 3730 1295 3736 1296
rect 3730 1291 3731 1295
rect 3735 1294 3736 1295
rect 3759 1295 3765 1296
rect 3759 1294 3760 1295
rect 3735 1292 3760 1294
rect 3735 1291 3736 1292
rect 3730 1290 3736 1291
rect 3759 1291 3760 1292
rect 3764 1291 3765 1295
rect 3759 1290 3765 1291
rect 3918 1295 3924 1296
rect 3918 1291 3919 1295
rect 3923 1294 3924 1295
rect 3927 1295 3933 1296
rect 3927 1294 3928 1295
rect 3923 1292 3928 1294
rect 3923 1291 3924 1292
rect 3918 1290 3924 1291
rect 3927 1291 3928 1292
rect 3932 1291 3933 1295
rect 3927 1290 3933 1291
rect 1582 1287 1588 1288
rect 1582 1283 1583 1287
rect 1587 1283 1588 1287
rect 1582 1282 1588 1283
rect 1113 1276 1161 1278
rect 1457 1276 1530 1278
rect 446 1274 452 1275
rect 1254 1275 1260 1276
rect 1254 1271 1255 1275
rect 1259 1271 1260 1275
rect 1254 1270 1260 1271
rect 1606 1275 1612 1276
rect 1606 1271 1607 1275
rect 1611 1271 1612 1275
rect 1606 1270 1612 1271
rect 2199 1275 2205 1276
rect 2199 1271 2200 1275
rect 2204 1274 2205 1275
rect 2279 1275 2285 1276
rect 2279 1274 2280 1275
rect 2204 1272 2280 1274
rect 2204 1271 2205 1272
rect 2199 1270 2205 1271
rect 2279 1271 2280 1272
rect 2284 1271 2285 1275
rect 2279 1270 2285 1271
rect 2367 1275 2373 1276
rect 2367 1271 2368 1275
rect 2372 1274 2373 1275
rect 2463 1275 2469 1276
rect 2463 1274 2464 1275
rect 2372 1272 2464 1274
rect 2372 1271 2373 1272
rect 2367 1270 2373 1271
rect 2463 1271 2464 1272
rect 2468 1271 2469 1275
rect 2463 1270 2469 1271
rect 2551 1275 2557 1276
rect 2551 1271 2552 1275
rect 2556 1274 2557 1275
rect 2663 1275 2669 1276
rect 2663 1274 2664 1275
rect 2556 1272 2664 1274
rect 2556 1271 2557 1272
rect 2551 1270 2557 1271
rect 2663 1271 2664 1272
rect 2668 1271 2669 1275
rect 2663 1270 2669 1271
rect 2671 1275 2677 1276
rect 2671 1271 2672 1275
rect 2676 1274 2677 1275
rect 2751 1275 2757 1276
rect 2751 1274 2752 1275
rect 2676 1272 2752 1274
rect 2676 1271 2677 1272
rect 2671 1270 2677 1271
rect 2751 1271 2752 1272
rect 2756 1271 2757 1275
rect 2751 1270 2757 1271
rect 2926 1275 2932 1276
rect 2926 1271 2927 1275
rect 2931 1274 2932 1275
rect 2951 1275 2957 1276
rect 2951 1274 2952 1275
rect 2931 1272 2952 1274
rect 2931 1271 2932 1272
rect 2926 1270 2932 1271
rect 2951 1271 2952 1272
rect 2956 1271 2957 1275
rect 2951 1270 2957 1271
rect 3006 1275 3012 1276
rect 3006 1271 3007 1275
rect 3011 1274 3012 1275
rect 3143 1275 3149 1276
rect 3143 1274 3144 1275
rect 3011 1272 3144 1274
rect 3011 1271 3012 1272
rect 3006 1270 3012 1271
rect 3143 1271 3144 1272
rect 3148 1271 3149 1275
rect 3143 1270 3149 1271
rect 3319 1275 3328 1276
rect 3319 1271 3320 1275
rect 3327 1271 3328 1275
rect 3487 1275 3493 1276
rect 3487 1274 3488 1275
rect 3319 1270 3328 1271
rect 3364 1272 3488 1274
rect 110 1268 116 1269
rect 110 1264 111 1268
rect 115 1264 116 1268
rect 110 1263 116 1264
rect 2030 1268 2036 1269
rect 2030 1264 2031 1268
rect 2035 1264 2036 1268
rect 2030 1263 2036 1264
rect 2126 1267 2132 1268
rect 2126 1263 2127 1267
rect 2131 1263 2132 1267
rect 2126 1262 2132 1263
rect 2294 1267 2300 1268
rect 2294 1263 2295 1267
rect 2299 1263 2300 1267
rect 2294 1262 2300 1263
rect 2478 1267 2484 1268
rect 2478 1263 2479 1267
rect 2483 1263 2484 1267
rect 2478 1262 2484 1263
rect 2678 1267 2684 1268
rect 2678 1263 2679 1267
rect 2683 1263 2684 1267
rect 2678 1262 2684 1263
rect 2878 1267 2884 1268
rect 2878 1263 2879 1267
rect 2883 1263 2884 1267
rect 2878 1262 2884 1263
rect 3070 1267 3076 1268
rect 3070 1263 3071 1267
rect 3075 1263 3076 1267
rect 3070 1262 3076 1263
rect 3246 1267 3252 1268
rect 3246 1263 3247 1267
rect 3251 1263 3252 1267
rect 3246 1262 3252 1263
rect 3364 1258 3366 1272
rect 3487 1271 3488 1272
rect 3492 1271 3493 1275
rect 3655 1275 3661 1276
rect 3655 1274 3656 1275
rect 3487 1270 3493 1271
rect 3529 1272 3656 1274
rect 3414 1267 3420 1268
rect 3414 1263 3415 1267
rect 3419 1263 3420 1267
rect 3414 1262 3420 1263
rect 3529 1258 3531 1272
rect 3655 1271 3656 1272
rect 3660 1271 3661 1275
rect 3823 1275 3829 1276
rect 3823 1274 3824 1275
rect 3655 1270 3661 1271
rect 3679 1272 3824 1274
rect 3582 1267 3588 1268
rect 3582 1263 3583 1267
rect 3587 1263 3588 1267
rect 3582 1262 3588 1263
rect 3679 1258 3681 1272
rect 3823 1271 3824 1272
rect 3828 1271 3829 1275
rect 3823 1270 3829 1271
rect 3926 1275 3932 1276
rect 3926 1271 3927 1275
rect 3931 1274 3932 1275
rect 3967 1275 3973 1276
rect 3967 1274 3968 1275
rect 3931 1272 3968 1274
rect 3931 1271 3932 1272
rect 3926 1270 3932 1271
rect 3967 1271 3968 1272
rect 3972 1271 3973 1275
rect 3967 1270 3973 1271
rect 3750 1267 3756 1268
rect 3750 1263 3751 1267
rect 3755 1263 3756 1267
rect 3750 1262 3756 1263
rect 3894 1267 3900 1268
rect 3894 1263 3895 1267
rect 3899 1263 3900 1267
rect 3894 1262 3900 1263
rect 3814 1259 3820 1260
rect 3814 1258 3815 1259
rect 3297 1256 3366 1258
rect 3465 1256 3531 1258
rect 3633 1256 3681 1258
rect 3801 1256 3815 1258
rect 2150 1255 2156 1256
rect 110 1251 116 1252
rect 110 1247 111 1251
rect 115 1247 116 1251
rect 2030 1251 2036 1252
rect 2030 1247 2031 1251
rect 2035 1247 2036 1251
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2870 1255 2876 1256
rect 2870 1251 2871 1255
rect 2875 1251 2876 1255
rect 2870 1250 2876 1251
rect 3086 1255 3092 1256
rect 3086 1251 3087 1255
rect 3091 1251 3092 1255
rect 3814 1255 3815 1256
rect 3819 1255 3820 1259
rect 3958 1259 3964 1260
rect 3958 1258 3959 1259
rect 3945 1256 3959 1258
rect 3814 1254 3820 1255
rect 3958 1255 3959 1256
rect 3963 1255 3964 1259
rect 3958 1254 3964 1255
rect 3086 1250 3092 1251
rect 110 1246 116 1247
rect 342 1246 348 1247
rect 342 1242 343 1246
rect 347 1242 348 1246
rect 342 1241 348 1242
rect 462 1246 468 1247
rect 462 1242 463 1246
rect 467 1242 468 1246
rect 462 1241 468 1242
rect 598 1246 604 1247
rect 598 1242 599 1246
rect 603 1242 604 1246
rect 598 1241 604 1242
rect 742 1246 748 1247
rect 742 1242 743 1246
rect 747 1242 748 1246
rect 742 1241 748 1242
rect 902 1246 908 1247
rect 902 1242 903 1246
rect 907 1242 908 1246
rect 902 1241 908 1242
rect 1062 1246 1068 1247
rect 1062 1242 1063 1246
rect 1067 1242 1068 1246
rect 1062 1241 1068 1242
rect 1230 1246 1236 1247
rect 1230 1242 1231 1246
rect 1235 1242 1236 1246
rect 1230 1241 1236 1242
rect 1406 1246 1412 1247
rect 1406 1242 1407 1246
rect 1411 1242 1412 1246
rect 1406 1241 1412 1242
rect 1582 1246 1588 1247
rect 2030 1246 2036 1247
rect 2070 1248 2076 1249
rect 1582 1242 1583 1246
rect 1587 1242 1588 1246
rect 2070 1244 2071 1248
rect 2075 1244 2076 1248
rect 2070 1243 2076 1244
rect 3990 1248 3996 1249
rect 3990 1244 3991 1248
rect 3995 1244 3996 1248
rect 3990 1243 3996 1244
rect 1582 1241 1588 1242
rect 446 1231 452 1232
rect 446 1227 447 1231
rect 451 1230 452 1231
rect 990 1231 996 1232
rect 990 1230 991 1231
rect 451 1228 991 1230
rect 451 1227 452 1228
rect 446 1226 452 1227
rect 990 1227 991 1228
rect 995 1227 996 1231
rect 990 1226 996 1227
rect 2070 1231 2076 1232
rect 2070 1227 2071 1231
rect 2075 1227 2076 1231
rect 3990 1231 3996 1232
rect 3990 1227 3991 1231
rect 3995 1227 3996 1231
rect 2070 1226 2076 1227
rect 2126 1226 2132 1227
rect 2126 1222 2127 1226
rect 2131 1222 2132 1226
rect 2126 1221 2132 1222
rect 2294 1226 2300 1227
rect 2294 1222 2295 1226
rect 2299 1222 2300 1226
rect 2294 1221 2300 1222
rect 2478 1226 2484 1227
rect 2478 1222 2479 1226
rect 2483 1222 2484 1226
rect 2478 1221 2484 1222
rect 2678 1226 2684 1227
rect 2678 1222 2679 1226
rect 2683 1222 2684 1226
rect 2678 1221 2684 1222
rect 2878 1226 2884 1227
rect 2878 1222 2879 1226
rect 2883 1222 2884 1226
rect 2878 1221 2884 1222
rect 3070 1226 3076 1227
rect 3070 1222 3071 1226
rect 3075 1222 3076 1226
rect 3070 1221 3076 1222
rect 3246 1226 3252 1227
rect 3246 1222 3247 1226
rect 3251 1222 3252 1226
rect 3246 1221 3252 1222
rect 3414 1226 3420 1227
rect 3414 1222 3415 1226
rect 3419 1222 3420 1226
rect 3414 1221 3420 1222
rect 3582 1226 3588 1227
rect 3582 1222 3583 1226
rect 3587 1222 3588 1226
rect 3582 1221 3588 1222
rect 3750 1226 3756 1227
rect 3750 1222 3751 1226
rect 3755 1222 3756 1226
rect 3750 1221 3756 1222
rect 3894 1226 3900 1227
rect 3990 1226 3996 1227
rect 3894 1222 3895 1226
rect 3899 1222 3900 1226
rect 3894 1221 3900 1222
rect 182 1214 188 1215
rect 182 1210 183 1214
rect 187 1210 188 1214
rect 110 1209 116 1210
rect 182 1209 188 1210
rect 350 1214 356 1215
rect 350 1210 351 1214
rect 355 1210 356 1214
rect 350 1209 356 1210
rect 534 1214 540 1215
rect 534 1210 535 1214
rect 539 1210 540 1214
rect 534 1209 540 1210
rect 726 1214 732 1215
rect 726 1210 727 1214
rect 731 1210 732 1214
rect 726 1209 732 1210
rect 918 1214 924 1215
rect 918 1210 919 1214
rect 923 1210 924 1214
rect 918 1209 924 1210
rect 1102 1214 1108 1215
rect 1102 1210 1103 1214
rect 1107 1210 1108 1214
rect 1102 1209 1108 1210
rect 1286 1214 1292 1215
rect 1286 1210 1287 1214
rect 1291 1210 1292 1214
rect 1286 1209 1292 1210
rect 1470 1214 1476 1215
rect 1470 1210 1471 1214
rect 1475 1210 1476 1214
rect 1470 1209 1476 1210
rect 1654 1214 1660 1215
rect 1654 1210 1655 1214
rect 1659 1210 1660 1214
rect 1654 1209 1660 1210
rect 1838 1214 1844 1215
rect 1838 1210 1839 1214
rect 1843 1210 1844 1214
rect 1838 1209 1844 1210
rect 2030 1209 2036 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 110 1204 116 1205
rect 2030 1205 2031 1209
rect 2035 1205 2036 1209
rect 2030 1204 2036 1205
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 110 1187 116 1188
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 334 1183 340 1184
rect 334 1182 335 1183
rect 233 1180 335 1182
rect 334 1179 335 1180
rect 339 1179 340 1183
rect 334 1178 340 1179
rect 1126 1183 1132 1184
rect 1126 1179 1127 1183
rect 1131 1179 1132 1183
rect 1414 1183 1420 1184
rect 1414 1182 1415 1183
rect 1337 1180 1415 1182
rect 1126 1178 1132 1179
rect 1414 1179 1415 1180
rect 1419 1179 1420 1183
rect 1414 1178 1420 1179
rect 2110 1182 2116 1183
rect 2110 1178 2111 1182
rect 2115 1178 2116 1182
rect 2070 1177 2076 1178
rect 2110 1177 2116 1178
rect 2246 1182 2252 1183
rect 2246 1178 2247 1182
rect 2251 1178 2252 1182
rect 2246 1177 2252 1178
rect 2406 1182 2412 1183
rect 2406 1178 2407 1182
rect 2411 1178 2412 1182
rect 2406 1177 2412 1178
rect 2558 1182 2564 1183
rect 2558 1178 2559 1182
rect 2563 1178 2564 1182
rect 2558 1177 2564 1178
rect 2702 1182 2708 1183
rect 2702 1178 2703 1182
rect 2707 1178 2708 1182
rect 2702 1177 2708 1178
rect 2862 1182 2868 1183
rect 2862 1178 2863 1182
rect 2867 1178 2868 1182
rect 2862 1177 2868 1178
rect 3038 1182 3044 1183
rect 3038 1178 3039 1182
rect 3043 1178 3044 1182
rect 3038 1177 3044 1178
rect 3238 1182 3244 1183
rect 3238 1178 3239 1182
rect 3243 1178 3244 1182
rect 3238 1177 3244 1178
rect 3454 1182 3460 1183
rect 3454 1178 3455 1182
rect 3459 1178 3460 1182
rect 3454 1177 3460 1178
rect 3686 1182 3692 1183
rect 3686 1178 3687 1182
rect 3691 1178 3692 1182
rect 3686 1177 3692 1178
rect 3894 1182 3900 1183
rect 3894 1178 3895 1182
rect 3899 1178 3900 1182
rect 3894 1177 3900 1178
rect 3990 1177 3996 1178
rect 182 1173 188 1174
rect 182 1169 183 1173
rect 187 1169 188 1173
rect 182 1168 188 1169
rect 350 1173 356 1174
rect 350 1169 351 1173
rect 355 1169 356 1173
rect 350 1168 356 1169
rect 534 1173 540 1174
rect 534 1169 535 1173
rect 539 1169 540 1173
rect 534 1168 540 1169
rect 726 1173 732 1174
rect 726 1169 727 1173
rect 731 1169 732 1173
rect 726 1168 732 1169
rect 918 1173 924 1174
rect 918 1169 919 1173
rect 923 1169 924 1173
rect 918 1168 924 1169
rect 1102 1173 1108 1174
rect 1102 1169 1103 1173
rect 1107 1169 1108 1173
rect 1102 1168 1108 1169
rect 1286 1173 1292 1174
rect 1286 1169 1287 1173
rect 1291 1169 1292 1173
rect 1286 1168 1292 1169
rect 1470 1173 1476 1174
rect 1470 1169 1471 1173
rect 1475 1169 1476 1173
rect 1470 1168 1476 1169
rect 1654 1173 1660 1174
rect 1654 1169 1655 1173
rect 1659 1169 1660 1173
rect 1654 1168 1660 1169
rect 1838 1173 1844 1174
rect 1838 1169 1839 1173
rect 1843 1169 1844 1173
rect 2070 1173 2071 1177
rect 2075 1173 2076 1177
rect 2070 1172 2076 1173
rect 3990 1173 3991 1177
rect 3995 1173 3996 1177
rect 3990 1172 3996 1173
rect 1838 1168 1844 1169
rect 255 1163 261 1164
rect 255 1159 256 1163
rect 260 1162 261 1163
rect 335 1163 341 1164
rect 335 1162 336 1163
rect 260 1160 336 1162
rect 260 1159 261 1160
rect 255 1158 261 1159
rect 335 1159 336 1160
rect 340 1159 341 1163
rect 335 1158 341 1159
rect 423 1163 429 1164
rect 423 1159 424 1163
rect 428 1162 429 1163
rect 519 1163 525 1164
rect 519 1162 520 1163
rect 428 1160 520 1162
rect 428 1159 429 1160
rect 423 1158 429 1159
rect 519 1159 520 1160
rect 524 1159 525 1163
rect 519 1158 525 1159
rect 607 1163 613 1164
rect 607 1159 608 1163
rect 612 1162 613 1163
rect 711 1163 717 1164
rect 711 1162 712 1163
rect 612 1160 712 1162
rect 612 1159 613 1160
rect 607 1158 613 1159
rect 711 1159 712 1160
rect 716 1159 717 1163
rect 711 1158 717 1159
rect 799 1163 805 1164
rect 799 1159 800 1163
rect 804 1162 805 1163
rect 903 1163 909 1164
rect 903 1162 904 1163
rect 804 1160 904 1162
rect 804 1159 805 1160
rect 799 1158 805 1159
rect 903 1159 904 1160
rect 908 1159 909 1163
rect 903 1158 909 1159
rect 990 1163 997 1164
rect 990 1159 991 1163
rect 996 1159 997 1163
rect 990 1158 997 1159
rect 1175 1163 1181 1164
rect 1175 1159 1176 1163
rect 1180 1162 1181 1163
rect 1186 1163 1192 1164
rect 1186 1162 1187 1163
rect 1180 1160 1187 1162
rect 1180 1159 1181 1160
rect 1175 1158 1181 1159
rect 1186 1159 1187 1160
rect 1191 1159 1192 1163
rect 1186 1158 1192 1159
rect 1359 1163 1365 1164
rect 1359 1159 1360 1163
rect 1364 1162 1365 1163
rect 1455 1163 1461 1164
rect 1455 1162 1456 1163
rect 1364 1160 1456 1162
rect 1364 1159 1365 1160
rect 1359 1158 1365 1159
rect 1455 1159 1456 1160
rect 1460 1159 1461 1163
rect 1455 1158 1461 1159
rect 1543 1163 1549 1164
rect 1543 1159 1544 1163
rect 1548 1162 1549 1163
rect 1639 1163 1645 1164
rect 1639 1162 1640 1163
rect 1548 1160 1640 1162
rect 1548 1159 1549 1160
rect 1543 1158 1549 1159
rect 1639 1159 1640 1160
rect 1644 1159 1645 1163
rect 1639 1158 1645 1159
rect 1727 1163 1733 1164
rect 1727 1159 1728 1163
rect 1732 1162 1733 1163
rect 1823 1163 1829 1164
rect 1823 1162 1824 1163
rect 1732 1160 1824 1162
rect 1732 1159 1733 1160
rect 1727 1158 1733 1159
rect 1823 1159 1824 1160
rect 1828 1159 1829 1163
rect 1823 1158 1829 1159
rect 1910 1163 1917 1164
rect 1910 1159 1911 1163
rect 1916 1159 1917 1163
rect 1910 1158 1917 1159
rect 2070 1160 2076 1161
rect 2070 1156 2071 1160
rect 2075 1156 2076 1160
rect 2070 1155 2076 1156
rect 3990 1160 3996 1161
rect 3990 1156 3991 1160
rect 3995 1156 3996 1160
rect 3990 1155 3996 1156
rect 334 1151 340 1152
rect 334 1147 335 1151
rect 339 1150 340 1151
rect 2230 1151 2236 1152
rect 2230 1150 2231 1151
rect 339 1148 906 1150
rect 2161 1148 2231 1150
rect 339 1147 340 1148
rect 334 1146 340 1147
rect 223 1143 229 1144
rect 223 1139 224 1143
rect 228 1142 229 1143
rect 287 1143 293 1144
rect 287 1142 288 1143
rect 228 1140 288 1142
rect 228 1139 229 1140
rect 223 1138 229 1139
rect 287 1139 288 1140
rect 292 1139 293 1143
rect 287 1138 293 1139
rect 375 1143 381 1144
rect 375 1139 376 1143
rect 380 1142 381 1143
rect 479 1143 485 1144
rect 479 1142 480 1143
rect 380 1140 480 1142
rect 380 1139 381 1140
rect 375 1138 381 1139
rect 479 1139 480 1140
rect 484 1139 485 1143
rect 479 1138 485 1139
rect 567 1143 573 1144
rect 567 1139 568 1143
rect 572 1142 573 1143
rect 687 1143 693 1144
rect 687 1142 688 1143
rect 572 1140 688 1142
rect 572 1139 573 1140
rect 567 1138 573 1139
rect 687 1139 688 1140
rect 692 1139 693 1143
rect 687 1138 693 1139
rect 775 1143 781 1144
rect 775 1139 776 1143
rect 780 1142 781 1143
rect 895 1143 901 1144
rect 895 1142 896 1143
rect 780 1140 896 1142
rect 780 1139 781 1140
rect 775 1138 781 1139
rect 895 1139 896 1140
rect 900 1139 901 1143
rect 904 1142 906 1148
rect 2230 1147 2231 1148
rect 2235 1147 2236 1151
rect 2390 1151 2396 1152
rect 2390 1150 2391 1151
rect 2297 1148 2391 1150
rect 2230 1146 2236 1147
rect 2390 1147 2391 1148
rect 2395 1147 2396 1151
rect 2503 1151 2509 1152
rect 2503 1150 2504 1151
rect 2457 1148 2504 1150
rect 2390 1146 2396 1147
rect 2503 1147 2504 1148
rect 2508 1147 2509 1151
rect 2662 1151 2668 1152
rect 2662 1150 2663 1151
rect 2609 1148 2663 1150
rect 2503 1146 2509 1147
rect 2662 1147 2663 1148
rect 2667 1147 2668 1151
rect 3006 1151 3012 1152
rect 3006 1150 3007 1151
rect 2913 1148 3007 1150
rect 2662 1146 2668 1147
rect 3006 1147 3007 1148
rect 3011 1147 3012 1151
rect 3966 1151 3972 1152
rect 3966 1150 3967 1151
rect 3945 1148 3967 1150
rect 3006 1146 3012 1147
rect 3966 1147 3967 1148
rect 3971 1147 3972 1151
rect 3966 1146 3972 1147
rect 983 1143 989 1144
rect 983 1142 984 1143
rect 904 1140 984 1142
rect 895 1138 901 1139
rect 983 1139 984 1140
rect 988 1139 989 1143
rect 983 1138 989 1139
rect 1082 1143 1088 1144
rect 1082 1139 1083 1143
rect 1087 1142 1088 1143
rect 1191 1143 1197 1144
rect 1191 1142 1192 1143
rect 1087 1140 1192 1142
rect 1087 1139 1088 1140
rect 1082 1138 1088 1139
rect 1191 1139 1192 1140
rect 1196 1139 1197 1143
rect 1191 1138 1197 1139
rect 1210 1143 1216 1144
rect 1210 1139 1211 1143
rect 1215 1142 1216 1143
rect 1391 1143 1397 1144
rect 1391 1142 1392 1143
rect 1215 1140 1392 1142
rect 1215 1139 1216 1140
rect 1210 1138 1216 1139
rect 1391 1139 1392 1140
rect 1396 1139 1397 1143
rect 1591 1143 1597 1144
rect 1591 1142 1592 1143
rect 1391 1138 1397 1139
rect 1452 1140 1592 1142
rect 150 1135 156 1136
rect 150 1131 151 1135
rect 155 1131 156 1135
rect 150 1130 156 1131
rect 302 1135 308 1136
rect 302 1131 303 1135
rect 307 1131 308 1135
rect 302 1130 308 1131
rect 494 1135 500 1136
rect 494 1131 495 1135
rect 499 1131 500 1135
rect 494 1130 500 1131
rect 702 1135 708 1136
rect 702 1131 703 1135
rect 707 1131 708 1135
rect 702 1130 708 1131
rect 910 1135 916 1136
rect 910 1131 911 1135
rect 915 1131 916 1135
rect 910 1130 916 1131
rect 1118 1135 1124 1136
rect 1118 1131 1119 1135
rect 1123 1131 1124 1135
rect 1118 1130 1124 1131
rect 1318 1135 1324 1136
rect 1318 1131 1319 1135
rect 1323 1131 1324 1135
rect 1318 1130 1324 1131
rect 231 1127 237 1128
rect 231 1126 232 1127
rect 201 1124 232 1126
rect 231 1123 232 1124
rect 236 1123 237 1127
rect 1186 1127 1192 1128
rect 1186 1126 1187 1127
rect 1169 1124 1187 1126
rect 231 1122 237 1123
rect 1186 1123 1187 1124
rect 1191 1123 1192 1127
rect 1452 1126 1454 1140
rect 1591 1139 1592 1140
rect 1596 1139 1597 1143
rect 1791 1143 1797 1144
rect 1791 1142 1792 1143
rect 1591 1138 1597 1139
rect 1652 1140 1792 1142
rect 1518 1135 1524 1136
rect 1518 1131 1519 1135
rect 1523 1131 1524 1135
rect 1518 1130 1524 1131
rect 1652 1126 1654 1140
rect 1791 1139 1792 1140
rect 1796 1139 1797 1143
rect 1991 1143 1997 1144
rect 1991 1142 1992 1143
rect 1791 1138 1797 1139
rect 1852 1140 1992 1142
rect 1718 1135 1724 1136
rect 1718 1131 1719 1135
rect 1723 1131 1724 1135
rect 1718 1130 1724 1131
rect 1852 1126 1854 1140
rect 1991 1139 1992 1140
rect 1996 1139 1997 1143
rect 1991 1138 1997 1139
rect 2110 1141 2116 1142
rect 2110 1137 2111 1141
rect 2115 1137 2116 1141
rect 2110 1136 2116 1137
rect 2246 1141 2252 1142
rect 2246 1137 2247 1141
rect 2251 1137 2252 1141
rect 2246 1136 2252 1137
rect 2406 1141 2412 1142
rect 2406 1137 2407 1141
rect 2411 1137 2412 1141
rect 2406 1136 2412 1137
rect 2558 1141 2564 1142
rect 2558 1137 2559 1141
rect 2563 1137 2564 1141
rect 2558 1136 2564 1137
rect 2702 1141 2708 1142
rect 2702 1137 2703 1141
rect 2707 1137 2708 1141
rect 2702 1136 2708 1137
rect 2862 1141 2868 1142
rect 2862 1137 2863 1141
rect 2867 1137 2868 1141
rect 2862 1136 2868 1137
rect 3038 1141 3044 1142
rect 3038 1137 3039 1141
rect 3043 1137 3044 1141
rect 3038 1136 3044 1137
rect 3238 1141 3244 1142
rect 3238 1137 3239 1141
rect 3243 1137 3244 1141
rect 3238 1136 3244 1137
rect 3454 1141 3460 1142
rect 3454 1137 3455 1141
rect 3459 1137 3460 1141
rect 3454 1136 3460 1137
rect 3686 1141 3692 1142
rect 3686 1137 3687 1141
rect 3691 1137 3692 1141
rect 3686 1136 3692 1137
rect 3894 1141 3900 1142
rect 3894 1137 3895 1141
rect 3899 1137 3900 1141
rect 3894 1136 3900 1137
rect 1918 1135 1924 1136
rect 1918 1131 1919 1135
rect 1923 1131 1924 1135
rect 1918 1130 1924 1131
rect 2150 1135 2156 1136
rect 2150 1131 2151 1135
rect 2155 1134 2156 1135
rect 2155 1133 2186 1134
rect 2155 1132 2189 1133
rect 2155 1131 2156 1132
rect 2150 1130 2156 1131
rect 2183 1128 2184 1132
rect 2188 1128 2189 1132
rect 1369 1124 1454 1126
rect 1569 1124 1654 1126
rect 1769 1124 1854 1126
rect 1910 1127 1916 1128
rect 2183 1127 2189 1128
rect 2230 1131 2236 1132
rect 2230 1127 2231 1131
rect 2235 1130 2236 1131
rect 2319 1131 2325 1132
rect 2319 1130 2320 1131
rect 2235 1128 2320 1130
rect 2235 1127 2236 1128
rect 1186 1122 1192 1123
rect 1910 1123 1911 1127
rect 1915 1123 1916 1127
rect 2230 1126 2236 1127
rect 2319 1127 2320 1128
rect 2324 1127 2325 1131
rect 2319 1126 2325 1127
rect 2390 1131 2396 1132
rect 2390 1127 2391 1131
rect 2395 1130 2396 1131
rect 2479 1131 2485 1132
rect 2479 1130 2480 1131
rect 2395 1128 2480 1130
rect 2395 1127 2396 1128
rect 2390 1126 2396 1127
rect 2479 1127 2480 1128
rect 2484 1127 2485 1131
rect 2479 1126 2485 1127
rect 2631 1131 2637 1132
rect 2631 1127 2632 1131
rect 2636 1130 2637 1131
rect 2687 1131 2693 1132
rect 2687 1130 2688 1131
rect 2636 1128 2688 1130
rect 2636 1127 2637 1128
rect 2631 1126 2637 1127
rect 2687 1127 2688 1128
rect 2692 1127 2693 1131
rect 2687 1126 2693 1127
rect 2775 1131 2781 1132
rect 2775 1127 2776 1131
rect 2780 1130 2781 1131
rect 2870 1131 2876 1132
rect 2870 1130 2871 1131
rect 2780 1128 2871 1130
rect 2780 1127 2781 1128
rect 2775 1126 2781 1127
rect 2870 1127 2871 1128
rect 2875 1127 2876 1131
rect 2870 1126 2876 1127
rect 2935 1131 2941 1132
rect 2935 1127 2936 1131
rect 2940 1130 2941 1131
rect 3023 1131 3029 1132
rect 3023 1130 3024 1131
rect 2940 1128 3024 1130
rect 2940 1127 2941 1128
rect 2935 1126 2941 1127
rect 3023 1127 3024 1128
rect 3028 1127 3029 1131
rect 3023 1126 3029 1127
rect 3111 1131 3117 1132
rect 3111 1127 3112 1131
rect 3116 1130 3117 1131
rect 3223 1131 3229 1132
rect 3223 1130 3224 1131
rect 3116 1128 3224 1130
rect 3116 1127 3117 1128
rect 3111 1126 3117 1127
rect 3223 1127 3224 1128
rect 3228 1127 3229 1131
rect 3223 1126 3229 1127
rect 3311 1131 3317 1132
rect 3311 1127 3312 1131
rect 3316 1130 3317 1131
rect 3439 1131 3445 1132
rect 3439 1130 3440 1131
rect 3316 1128 3440 1130
rect 3316 1127 3317 1128
rect 3311 1126 3317 1127
rect 3439 1127 3440 1128
rect 3444 1127 3445 1131
rect 3439 1126 3445 1127
rect 3527 1131 3533 1132
rect 3527 1127 3528 1131
rect 3532 1130 3533 1131
rect 3671 1131 3677 1132
rect 3671 1130 3672 1131
rect 3532 1128 3672 1130
rect 3532 1127 3533 1128
rect 3527 1126 3533 1127
rect 3671 1127 3672 1128
rect 3676 1127 3677 1131
rect 3759 1131 3765 1132
rect 3759 1130 3760 1131
rect 3671 1126 3677 1127
rect 3679 1128 3760 1130
rect 1910 1122 1916 1123
rect 3070 1123 3076 1124
rect 3070 1119 3071 1123
rect 3075 1122 3076 1123
rect 3679 1122 3681 1128
rect 3759 1127 3760 1128
rect 3764 1127 3765 1131
rect 3759 1126 3765 1127
rect 3958 1131 3964 1132
rect 3958 1127 3959 1131
rect 3963 1130 3964 1131
rect 3967 1131 3973 1132
rect 3967 1130 3968 1131
rect 3963 1128 3968 1130
rect 3963 1127 3964 1128
rect 3958 1126 3964 1127
rect 3967 1127 3968 1128
rect 3972 1127 3973 1131
rect 3967 1126 3973 1127
rect 3075 1120 3681 1122
rect 3075 1119 3076 1120
rect 3070 1118 3076 1119
rect 110 1116 116 1117
rect 110 1112 111 1116
rect 115 1112 116 1116
rect 110 1111 116 1112
rect 2030 1116 2036 1117
rect 2030 1112 2031 1116
rect 2035 1112 2036 1116
rect 2030 1111 2036 1112
rect 2183 1115 2189 1116
rect 2183 1111 2184 1115
rect 2188 1114 2189 1115
rect 2287 1115 2293 1116
rect 2287 1114 2288 1115
rect 2188 1112 2288 1114
rect 2188 1111 2189 1112
rect 2183 1110 2189 1111
rect 2287 1111 2288 1112
rect 2292 1111 2293 1115
rect 2287 1110 2293 1111
rect 2375 1115 2381 1116
rect 2375 1111 2376 1115
rect 2380 1114 2381 1115
rect 2495 1115 2501 1116
rect 2495 1114 2496 1115
rect 2380 1112 2496 1114
rect 2380 1111 2381 1112
rect 2375 1110 2381 1111
rect 2495 1111 2496 1112
rect 2500 1111 2501 1115
rect 2495 1110 2501 1111
rect 2503 1115 2509 1116
rect 2503 1111 2504 1115
rect 2508 1114 2509 1115
rect 2583 1115 2589 1116
rect 2583 1114 2584 1115
rect 2508 1112 2584 1114
rect 2508 1111 2509 1112
rect 2503 1110 2509 1111
rect 2583 1111 2584 1112
rect 2588 1111 2589 1115
rect 2583 1110 2589 1111
rect 2662 1115 2668 1116
rect 2662 1111 2663 1115
rect 2667 1114 2668 1115
rect 2775 1115 2781 1116
rect 2775 1114 2776 1115
rect 2667 1112 2776 1114
rect 2667 1111 2668 1112
rect 2662 1110 2668 1111
rect 2775 1111 2776 1112
rect 2780 1111 2781 1115
rect 2775 1110 2781 1111
rect 2967 1115 2973 1116
rect 2967 1111 2968 1115
rect 2972 1114 2973 1115
rect 3071 1115 3077 1116
rect 3071 1114 3072 1115
rect 2972 1112 3072 1114
rect 2972 1111 2973 1112
rect 2967 1110 2973 1111
rect 3071 1111 3072 1112
rect 3076 1111 3077 1115
rect 3071 1110 3077 1111
rect 3159 1115 3165 1116
rect 3159 1111 3160 1115
rect 3164 1114 3165 1115
rect 3271 1115 3277 1116
rect 3271 1114 3272 1115
rect 3164 1112 3272 1114
rect 3164 1111 3165 1112
rect 3159 1110 3165 1111
rect 3271 1111 3272 1112
rect 3276 1111 3277 1115
rect 3271 1110 3277 1111
rect 3359 1115 3365 1116
rect 3359 1111 3360 1115
rect 3364 1114 3365 1115
rect 3479 1115 3485 1116
rect 3479 1114 3480 1115
rect 3364 1112 3480 1114
rect 3364 1111 3365 1112
rect 3359 1110 3365 1111
rect 3479 1111 3480 1112
rect 3484 1111 3485 1115
rect 3479 1110 3485 1111
rect 3567 1115 3573 1116
rect 3567 1111 3568 1115
rect 3572 1114 3573 1115
rect 3687 1115 3693 1116
rect 3687 1114 3688 1115
rect 3572 1112 3688 1114
rect 3572 1111 3573 1112
rect 3567 1110 3573 1111
rect 3687 1111 3688 1112
rect 3692 1111 3693 1115
rect 3687 1110 3693 1111
rect 3758 1115 3764 1116
rect 3758 1111 3759 1115
rect 3763 1114 3764 1115
rect 3775 1115 3781 1116
rect 3775 1114 3776 1115
rect 3763 1112 3776 1114
rect 3763 1111 3764 1112
rect 3758 1110 3764 1111
rect 3775 1111 3776 1112
rect 3780 1111 3781 1115
rect 3775 1110 3781 1111
rect 3966 1115 3973 1116
rect 3966 1111 3967 1115
rect 3972 1111 3973 1115
rect 3966 1110 3973 1111
rect 2110 1107 2116 1108
rect 2110 1103 2111 1107
rect 2115 1103 2116 1107
rect 2110 1102 2116 1103
rect 2302 1107 2308 1108
rect 2302 1103 2303 1107
rect 2307 1103 2308 1107
rect 2302 1102 2308 1103
rect 2510 1107 2516 1108
rect 2510 1103 2511 1107
rect 2515 1103 2516 1107
rect 2510 1102 2516 1103
rect 2702 1107 2708 1108
rect 2702 1103 2703 1107
rect 2707 1103 2708 1107
rect 2702 1102 2708 1103
rect 2894 1107 2900 1108
rect 2894 1103 2895 1107
rect 2899 1103 2900 1107
rect 2894 1102 2900 1103
rect 3086 1107 3092 1108
rect 3086 1103 3087 1107
rect 3091 1103 3092 1107
rect 3086 1102 3092 1103
rect 3286 1107 3292 1108
rect 3286 1103 3287 1107
rect 3291 1103 3292 1107
rect 3286 1102 3292 1103
rect 3494 1107 3500 1108
rect 3494 1103 3495 1107
rect 3499 1103 3500 1107
rect 3494 1102 3500 1103
rect 3702 1107 3708 1108
rect 3702 1103 3703 1107
rect 3707 1103 3708 1107
rect 3702 1102 3708 1103
rect 3894 1107 3900 1108
rect 3894 1103 3895 1107
rect 3899 1103 3900 1107
rect 3894 1102 3900 1103
rect 110 1099 116 1100
rect 110 1095 111 1099
rect 115 1095 116 1099
rect 2030 1099 2036 1100
rect 2030 1095 2031 1099
rect 2035 1095 2036 1099
rect 2878 1099 2884 1100
rect 2878 1098 2879 1099
rect 2753 1096 2879 1098
rect 110 1094 116 1095
rect 150 1094 156 1095
rect 150 1090 151 1094
rect 155 1090 156 1094
rect 150 1089 156 1090
rect 302 1094 308 1095
rect 302 1090 303 1094
rect 307 1090 308 1094
rect 302 1089 308 1090
rect 494 1094 500 1095
rect 494 1090 495 1094
rect 499 1090 500 1094
rect 494 1089 500 1090
rect 702 1094 708 1095
rect 702 1090 703 1094
rect 707 1090 708 1094
rect 702 1089 708 1090
rect 910 1094 916 1095
rect 910 1090 911 1094
rect 915 1090 916 1094
rect 910 1089 916 1090
rect 1118 1094 1124 1095
rect 1118 1090 1119 1094
rect 1123 1090 1124 1094
rect 1118 1089 1124 1090
rect 1318 1094 1324 1095
rect 1318 1090 1319 1094
rect 1323 1090 1324 1094
rect 1318 1089 1324 1090
rect 1518 1094 1524 1095
rect 1518 1090 1519 1094
rect 1523 1090 1524 1094
rect 1518 1089 1524 1090
rect 1718 1094 1724 1095
rect 1718 1090 1719 1094
rect 1723 1090 1724 1094
rect 1718 1089 1724 1090
rect 1918 1094 1924 1095
rect 2030 1094 2036 1095
rect 2102 1095 2108 1096
rect 1918 1090 1919 1094
rect 1923 1090 1924 1094
rect 2102 1091 2103 1095
rect 2107 1091 2108 1095
rect 2878 1095 2879 1096
rect 2883 1095 2884 1099
rect 3070 1099 3076 1100
rect 3070 1098 3071 1099
rect 2945 1096 3071 1098
rect 2878 1094 2884 1095
rect 3070 1095 3071 1096
rect 3075 1095 3076 1099
rect 3958 1099 3964 1100
rect 3958 1098 3959 1099
rect 3945 1096 3959 1098
rect 3070 1094 3076 1095
rect 3958 1095 3959 1096
rect 3963 1095 3964 1099
rect 3958 1094 3964 1095
rect 2102 1090 2108 1091
rect 1918 1089 1924 1090
rect 2070 1088 2076 1089
rect 2070 1084 2071 1088
rect 2075 1084 2076 1088
rect 2070 1083 2076 1084
rect 3990 1088 3996 1089
rect 3990 1084 3991 1088
rect 3995 1084 3996 1088
rect 3990 1083 3996 1084
rect 2070 1071 2076 1072
rect 2070 1067 2071 1071
rect 2075 1067 2076 1071
rect 3990 1071 3996 1072
rect 3990 1067 3991 1071
rect 3995 1067 3996 1071
rect 2070 1066 2076 1067
rect 2110 1066 2116 1067
rect 2110 1062 2111 1066
rect 2115 1062 2116 1066
rect 2110 1061 2116 1062
rect 2302 1066 2308 1067
rect 2302 1062 2303 1066
rect 2307 1062 2308 1066
rect 2302 1061 2308 1062
rect 2510 1066 2516 1067
rect 2510 1062 2511 1066
rect 2515 1062 2516 1066
rect 2510 1061 2516 1062
rect 2702 1066 2708 1067
rect 2702 1062 2703 1066
rect 2707 1062 2708 1066
rect 2702 1061 2708 1062
rect 2894 1066 2900 1067
rect 2894 1062 2895 1066
rect 2899 1062 2900 1066
rect 2894 1061 2900 1062
rect 3086 1066 3092 1067
rect 3086 1062 3087 1066
rect 3091 1062 3092 1066
rect 3086 1061 3092 1062
rect 3286 1066 3292 1067
rect 3286 1062 3287 1066
rect 3291 1062 3292 1066
rect 3286 1061 3292 1062
rect 3494 1066 3500 1067
rect 3494 1062 3495 1066
rect 3499 1062 3500 1066
rect 3494 1061 3500 1062
rect 3702 1066 3708 1067
rect 3702 1062 3703 1066
rect 3707 1062 3708 1066
rect 3702 1061 3708 1062
rect 3894 1066 3900 1067
rect 3990 1066 3996 1067
rect 3894 1062 3895 1066
rect 3899 1062 3900 1066
rect 3894 1061 3900 1062
rect 150 1054 156 1055
rect 150 1050 151 1054
rect 155 1050 156 1054
rect 110 1049 116 1050
rect 150 1049 156 1050
rect 278 1054 284 1055
rect 278 1050 279 1054
rect 283 1050 284 1054
rect 278 1049 284 1050
rect 446 1054 452 1055
rect 446 1050 447 1054
rect 451 1050 452 1054
rect 446 1049 452 1050
rect 622 1054 628 1055
rect 622 1050 623 1054
rect 627 1050 628 1054
rect 622 1049 628 1050
rect 798 1054 804 1055
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 966 1054 972 1055
rect 966 1050 967 1054
rect 971 1050 972 1054
rect 966 1049 972 1050
rect 1126 1054 1132 1055
rect 1126 1050 1127 1054
rect 1131 1050 1132 1054
rect 1126 1049 1132 1050
rect 1278 1054 1284 1055
rect 1278 1050 1279 1054
rect 1283 1050 1284 1054
rect 1278 1049 1284 1050
rect 1422 1054 1428 1055
rect 1422 1050 1423 1054
rect 1427 1050 1428 1054
rect 1422 1049 1428 1050
rect 1558 1054 1564 1055
rect 1558 1050 1559 1054
rect 1563 1050 1564 1054
rect 1558 1049 1564 1050
rect 1694 1054 1700 1055
rect 1694 1050 1695 1054
rect 1699 1050 1700 1054
rect 1694 1049 1700 1050
rect 1822 1054 1828 1055
rect 1822 1050 1823 1054
rect 1827 1050 1828 1054
rect 1822 1049 1828 1050
rect 1934 1054 1940 1055
rect 1934 1050 1935 1054
rect 1939 1050 1940 1054
rect 1934 1049 1940 1050
rect 2030 1049 2036 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 2030 1045 2031 1049
rect 2035 1045 2036 1049
rect 2030 1044 2036 1045
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 2030 1032 2036 1033
rect 2030 1028 2031 1032
rect 2035 1028 2036 1032
rect 2030 1027 2036 1028
rect 222 1023 228 1024
rect 222 1022 223 1023
rect 201 1020 223 1022
rect 222 1019 223 1020
rect 227 1019 228 1023
rect 1082 1023 1088 1024
rect 1082 1022 1083 1023
rect 1017 1020 1083 1022
rect 222 1018 228 1019
rect 1082 1019 1083 1020
rect 1087 1019 1088 1023
rect 1210 1023 1216 1024
rect 1210 1022 1211 1023
rect 1177 1020 1211 1022
rect 1082 1018 1088 1019
rect 1210 1019 1211 1020
rect 1215 1019 1216 1023
rect 1406 1023 1412 1024
rect 1406 1022 1407 1023
rect 1329 1020 1407 1022
rect 1210 1018 1216 1019
rect 1406 1019 1407 1020
rect 1411 1019 1412 1023
rect 1406 1018 1412 1019
rect 2318 1018 2324 1019
rect 2318 1014 2319 1018
rect 2323 1014 2324 1018
rect 150 1013 156 1014
rect 150 1009 151 1013
rect 155 1009 156 1013
rect 150 1008 156 1009
rect 278 1013 284 1014
rect 278 1009 279 1013
rect 283 1009 284 1013
rect 278 1008 284 1009
rect 446 1013 452 1014
rect 446 1009 447 1013
rect 451 1009 452 1013
rect 446 1008 452 1009
rect 622 1013 628 1014
rect 622 1009 623 1013
rect 627 1009 628 1013
rect 622 1008 628 1009
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 966 1013 972 1014
rect 966 1009 967 1013
rect 971 1009 972 1013
rect 966 1008 972 1009
rect 1126 1013 1132 1014
rect 1126 1009 1127 1013
rect 1131 1009 1132 1013
rect 1126 1008 1132 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 1422 1013 1428 1014
rect 1422 1009 1423 1013
rect 1427 1009 1428 1013
rect 1422 1008 1428 1009
rect 1558 1013 1564 1014
rect 1558 1009 1559 1013
rect 1563 1009 1564 1013
rect 1558 1008 1564 1009
rect 1694 1013 1700 1014
rect 1694 1009 1695 1013
rect 1699 1009 1700 1013
rect 1694 1008 1700 1009
rect 1822 1013 1828 1014
rect 1822 1009 1823 1013
rect 1827 1009 1828 1013
rect 1822 1008 1828 1009
rect 1934 1013 1940 1014
rect 1934 1009 1935 1013
rect 1939 1009 1940 1013
rect 1934 1008 1940 1009
rect 2070 1013 2076 1014
rect 2318 1013 2324 1014
rect 2486 1018 2492 1019
rect 2486 1014 2487 1018
rect 2491 1014 2492 1018
rect 2486 1013 2492 1014
rect 2662 1018 2668 1019
rect 2662 1014 2663 1018
rect 2667 1014 2668 1018
rect 2662 1013 2668 1014
rect 2846 1018 2852 1019
rect 2846 1014 2847 1018
rect 2851 1014 2852 1018
rect 2846 1013 2852 1014
rect 3038 1018 3044 1019
rect 3038 1014 3039 1018
rect 3043 1014 3044 1018
rect 3038 1013 3044 1014
rect 3246 1018 3252 1019
rect 3246 1014 3247 1018
rect 3251 1014 3252 1018
rect 3246 1013 3252 1014
rect 3462 1018 3468 1019
rect 3462 1014 3463 1018
rect 3467 1014 3468 1018
rect 3462 1013 3468 1014
rect 3686 1018 3692 1019
rect 3686 1014 3687 1018
rect 3691 1014 3692 1018
rect 3686 1013 3692 1014
rect 3894 1018 3900 1019
rect 3894 1014 3895 1018
rect 3899 1014 3900 1018
rect 3894 1013 3900 1014
rect 3990 1013 3996 1014
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 3990 1009 3991 1013
rect 3995 1009 3996 1013
rect 3990 1008 3996 1009
rect 223 1003 229 1004
rect 223 999 224 1003
rect 228 1002 229 1003
rect 263 1003 269 1004
rect 263 1002 264 1003
rect 228 1000 264 1002
rect 228 999 229 1000
rect 223 998 229 999
rect 263 999 264 1000
rect 268 999 269 1003
rect 263 998 269 999
rect 351 1003 357 1004
rect 351 999 352 1003
rect 356 1002 357 1003
rect 431 1003 437 1004
rect 431 1002 432 1003
rect 356 1000 432 1002
rect 356 999 357 1000
rect 351 998 357 999
rect 431 999 432 1000
rect 436 999 437 1003
rect 431 998 437 999
rect 519 1003 525 1004
rect 519 999 520 1003
rect 524 1002 525 1003
rect 607 1003 613 1004
rect 607 1002 608 1003
rect 524 1000 608 1002
rect 524 999 525 1000
rect 519 998 525 999
rect 607 999 608 1000
rect 612 999 613 1003
rect 607 998 613 999
rect 695 1003 701 1004
rect 695 999 696 1003
rect 700 1002 701 1003
rect 783 1003 789 1004
rect 783 1002 784 1003
rect 700 1000 784 1002
rect 700 999 701 1000
rect 695 998 701 999
rect 783 999 784 1000
rect 788 999 789 1003
rect 871 1003 877 1004
rect 871 1002 872 1003
rect 783 998 789 999
rect 792 1000 872 1002
rect 231 995 237 996
rect 231 991 232 995
rect 236 994 237 995
rect 792 994 794 1000
rect 871 999 872 1000
rect 876 999 877 1003
rect 871 998 877 999
rect 1039 1003 1048 1004
rect 1039 999 1040 1003
rect 1047 999 1048 1003
rect 1039 998 1048 999
rect 1199 1003 1208 1004
rect 1199 999 1200 1003
rect 1207 999 1208 1003
rect 1199 998 1208 999
rect 1351 1003 1357 1004
rect 1351 999 1352 1003
rect 1356 1002 1357 1003
rect 1407 1003 1413 1004
rect 1407 1002 1408 1003
rect 1356 1000 1408 1002
rect 1356 999 1357 1000
rect 1351 998 1357 999
rect 1407 999 1408 1000
rect 1412 999 1413 1003
rect 1407 998 1413 999
rect 1495 1003 1501 1004
rect 1495 999 1496 1003
rect 1500 1002 1501 1003
rect 1543 1003 1549 1004
rect 1543 1002 1544 1003
rect 1500 1000 1544 1002
rect 1500 999 1501 1000
rect 1495 998 1501 999
rect 1543 999 1544 1000
rect 1548 999 1549 1003
rect 1543 998 1549 999
rect 1631 1003 1637 1004
rect 1631 999 1632 1003
rect 1636 1002 1637 1003
rect 1679 1003 1685 1004
rect 1679 1002 1680 1003
rect 1636 1000 1680 1002
rect 1636 999 1637 1000
rect 1631 998 1637 999
rect 1679 999 1680 1000
rect 1684 999 1685 1003
rect 1679 998 1685 999
rect 1767 1003 1773 1004
rect 1767 999 1768 1003
rect 1772 1002 1773 1003
rect 1807 1003 1813 1004
rect 1807 1002 1808 1003
rect 1772 1000 1808 1002
rect 1772 999 1773 1000
rect 1767 998 1773 999
rect 1807 999 1808 1000
rect 1812 999 1813 1003
rect 1807 998 1813 999
rect 1895 1003 1901 1004
rect 1895 999 1896 1003
rect 1900 1002 1901 1003
rect 1919 1003 1925 1004
rect 1919 1002 1920 1003
rect 1900 1000 1920 1002
rect 1900 999 1901 1000
rect 1895 998 1901 999
rect 1919 999 1920 1000
rect 1924 999 1925 1003
rect 1919 998 1925 999
rect 2007 1003 2013 1004
rect 2007 999 2008 1003
rect 2012 1002 2013 1003
rect 2102 1003 2108 1004
rect 2102 1002 2103 1003
rect 2012 1000 2103 1002
rect 2012 999 2013 1000
rect 2007 998 2013 999
rect 2102 999 2103 1000
rect 2107 999 2108 1003
rect 2102 998 2108 999
rect 236 992 794 994
rect 2070 996 2076 997
rect 2070 992 2071 996
rect 2075 992 2076 996
rect 236 991 237 992
rect 2070 991 2076 992
rect 3990 996 3996 997
rect 3990 992 3991 996
rect 3995 992 3996 996
rect 3990 991 3996 992
rect 231 990 237 991
rect 1406 987 1412 988
rect 1406 983 1407 987
rect 1411 986 1412 987
rect 2423 987 2429 988
rect 2423 986 2424 987
rect 1411 984 1578 986
rect 2369 984 2424 986
rect 1411 983 1412 984
rect 1406 982 1412 983
rect 222 979 229 980
rect 222 975 223 979
rect 228 975 229 979
rect 359 979 365 980
rect 359 978 360 979
rect 222 974 229 975
rect 268 976 360 978
rect 150 971 156 972
rect 150 967 151 971
rect 155 967 156 971
rect 150 966 156 967
rect 268 962 270 976
rect 359 975 360 976
rect 364 975 365 979
rect 543 979 549 980
rect 543 978 544 979
rect 359 974 365 975
rect 444 976 544 978
rect 286 971 292 972
rect 286 967 287 971
rect 291 967 292 971
rect 286 966 292 967
rect 444 962 446 976
rect 543 975 544 976
rect 548 975 549 979
rect 543 974 549 975
rect 743 979 749 980
rect 743 975 744 979
rect 748 978 749 979
rect 855 979 861 980
rect 855 978 856 979
rect 748 976 856 978
rect 748 975 749 976
rect 743 974 749 975
rect 855 975 856 976
rect 860 975 861 979
rect 943 979 949 980
rect 943 978 944 979
rect 936 976 944 978
rect 855 974 861 975
rect 934 975 940 976
rect 470 971 476 972
rect 470 967 471 971
rect 475 967 476 971
rect 470 966 476 967
rect 670 971 676 972
rect 670 967 671 971
rect 675 967 676 971
rect 670 966 676 967
rect 870 971 876 972
rect 870 967 871 971
rect 875 967 876 971
rect 934 971 935 975
rect 939 971 940 975
rect 943 975 944 976
rect 948 975 949 979
rect 943 974 949 975
rect 1042 979 1048 980
rect 1042 975 1043 979
rect 1047 978 1048 979
rect 1063 979 1069 980
rect 1063 978 1064 979
rect 1047 976 1064 978
rect 1047 975 1048 976
rect 1042 974 1048 975
rect 1063 975 1064 976
rect 1068 975 1069 979
rect 1151 979 1157 980
rect 1151 978 1152 979
rect 1063 974 1069 975
rect 1072 976 1152 978
rect 934 970 940 971
rect 998 971 1004 972
rect 870 966 876 967
rect 998 967 999 971
rect 1003 970 1004 971
rect 1072 970 1074 976
rect 1151 975 1152 976
rect 1156 975 1157 979
rect 1151 974 1157 975
rect 1202 979 1208 980
rect 1202 975 1203 979
rect 1207 978 1208 979
rect 1271 979 1277 980
rect 1271 978 1272 979
rect 1207 976 1272 978
rect 1207 975 1208 976
rect 1202 974 1208 975
rect 1271 975 1272 976
rect 1276 975 1277 979
rect 1271 974 1277 975
rect 1359 979 1365 980
rect 1359 975 1360 979
rect 1364 978 1365 979
rect 1479 979 1485 980
rect 1479 978 1480 979
rect 1364 976 1480 978
rect 1364 975 1365 976
rect 1359 974 1365 975
rect 1479 975 1480 976
rect 1484 975 1485 979
rect 1479 974 1485 975
rect 1502 979 1508 980
rect 1502 975 1503 979
rect 1507 978 1508 979
rect 1567 979 1573 980
rect 1567 978 1568 979
rect 1507 976 1568 978
rect 1507 975 1508 976
rect 1502 974 1508 975
rect 1567 975 1568 976
rect 1572 975 1573 979
rect 1576 978 1578 984
rect 2423 983 2424 984
rect 2428 983 2429 987
rect 3446 987 3452 988
rect 3446 986 3447 987
rect 2897 984 2970 986
rect 3297 984 3447 986
rect 2423 982 2429 983
rect 1775 979 1781 980
rect 1775 978 1776 979
rect 1576 976 1776 978
rect 1567 974 1573 975
rect 1775 975 1776 976
rect 1780 975 1781 979
rect 1983 979 1989 980
rect 1983 978 1984 979
rect 1775 974 1781 975
rect 1836 976 1984 978
rect 1003 968 1074 970
rect 1078 971 1084 972
rect 1003 967 1004 968
rect 998 966 1004 967
rect 1078 967 1079 971
rect 1083 967 1084 971
rect 1078 966 1084 967
rect 1286 971 1292 972
rect 1286 967 1287 971
rect 1291 967 1292 971
rect 1286 966 1292 967
rect 1494 971 1500 972
rect 1494 967 1495 971
rect 1499 967 1500 971
rect 1494 966 1500 967
rect 1702 971 1708 972
rect 1702 967 1703 971
rect 1707 967 1708 971
rect 1702 966 1708 967
rect 654 963 660 964
rect 654 962 655 963
rect 201 960 270 962
rect 337 960 446 962
rect 521 960 655 962
rect 654 959 655 960
rect 659 959 660 963
rect 1836 962 1838 976
rect 1983 975 1984 976
rect 1988 975 1989 979
rect 2968 978 2970 984
rect 3446 983 3447 984
rect 3451 983 3452 987
rect 3567 987 3573 988
rect 3567 986 3568 987
rect 3513 984 3568 986
rect 3446 982 3452 983
rect 3567 983 3568 984
rect 3572 983 3573 987
rect 3758 987 3764 988
rect 3758 986 3759 987
rect 3737 984 3759 986
rect 3567 982 3573 983
rect 3758 983 3759 984
rect 3763 983 3764 987
rect 3966 987 3972 988
rect 3966 986 3967 987
rect 3945 984 3967 986
rect 3758 982 3764 983
rect 3966 983 3967 984
rect 3971 983 3972 987
rect 3966 982 3972 983
rect 1983 974 1989 975
rect 2318 977 2324 978
rect 2318 973 2319 977
rect 2323 973 2324 977
rect 2318 972 2324 973
rect 2486 977 2492 978
rect 2486 973 2487 977
rect 2491 973 2492 977
rect 2486 972 2492 973
rect 2662 977 2668 978
rect 2662 973 2663 977
rect 2667 973 2668 977
rect 2662 972 2668 973
rect 2846 977 2852 978
rect 2846 973 2847 977
rect 2851 973 2852 977
rect 2968 976 3034 978
rect 2846 972 2852 973
rect 1910 971 1916 972
rect 1910 967 1911 971
rect 1915 967 1916 971
rect 1910 966 1916 967
rect 2391 967 2397 968
rect 1982 963 1988 964
rect 1982 962 1983 963
rect 1753 960 1838 962
rect 1961 960 1983 962
rect 654 958 660 959
rect 662 959 668 960
rect 662 955 663 959
rect 667 955 668 959
rect 1982 959 1983 960
rect 1987 959 1988 963
rect 2391 963 2392 967
rect 2396 966 2397 967
rect 2471 967 2477 968
rect 2471 966 2472 967
rect 2396 964 2472 966
rect 2396 963 2397 964
rect 2391 962 2397 963
rect 2471 963 2472 964
rect 2476 963 2477 967
rect 2471 962 2477 963
rect 2559 967 2565 968
rect 2559 963 2560 967
rect 2564 966 2565 967
rect 2647 967 2653 968
rect 2647 966 2648 967
rect 2564 964 2648 966
rect 2564 963 2565 964
rect 2559 962 2565 963
rect 2647 963 2648 964
rect 2652 963 2653 967
rect 2647 962 2653 963
rect 2670 967 2676 968
rect 2670 963 2671 967
rect 2675 966 2676 967
rect 2735 967 2741 968
rect 2735 966 2736 967
rect 2675 964 2736 966
rect 2675 963 2676 964
rect 2670 962 2676 963
rect 2735 963 2736 964
rect 2740 963 2741 967
rect 2735 962 2741 963
rect 2878 967 2884 968
rect 2878 963 2879 967
rect 2883 966 2884 967
rect 2919 967 2925 968
rect 2919 966 2920 967
rect 2883 964 2920 966
rect 2883 963 2884 964
rect 2878 962 2884 963
rect 2919 963 2920 964
rect 2924 963 2925 967
rect 2919 962 2925 963
rect 3023 967 3029 968
rect 3023 963 3024 967
rect 3028 963 3029 967
rect 3032 966 3034 976
rect 3038 977 3044 978
rect 3038 973 3039 977
rect 3043 973 3044 977
rect 3038 972 3044 973
rect 3246 977 3252 978
rect 3246 973 3247 977
rect 3251 973 3252 977
rect 3246 972 3252 973
rect 3462 977 3468 978
rect 3462 973 3463 977
rect 3467 973 3468 977
rect 3462 972 3468 973
rect 3686 977 3692 978
rect 3686 973 3687 977
rect 3691 973 3692 977
rect 3686 972 3692 973
rect 3894 977 3900 978
rect 3894 973 3895 977
rect 3899 973 3900 977
rect 3894 972 3900 973
rect 3111 967 3117 968
rect 3111 966 3112 967
rect 3032 964 3112 966
rect 3023 962 3029 963
rect 3111 963 3112 964
rect 3116 963 3117 967
rect 3111 962 3117 963
rect 3214 967 3220 968
rect 3214 963 3215 967
rect 3219 966 3220 967
rect 3319 967 3325 968
rect 3319 966 3320 967
rect 3219 964 3320 966
rect 3219 963 3220 964
rect 3214 962 3220 963
rect 3319 963 3320 964
rect 3324 963 3325 967
rect 3319 962 3325 963
rect 3446 967 3452 968
rect 3446 963 3447 967
rect 3451 966 3452 967
rect 3535 967 3541 968
rect 3535 966 3536 967
rect 3451 964 3536 966
rect 3451 963 3452 964
rect 3446 962 3452 963
rect 3535 963 3536 964
rect 3540 963 3541 967
rect 3535 962 3541 963
rect 3567 967 3573 968
rect 3567 963 3568 967
rect 3572 966 3573 967
rect 3759 967 3765 968
rect 3759 966 3760 967
rect 3572 964 3760 966
rect 3572 963 3573 964
rect 3567 962 3573 963
rect 3759 963 3760 964
rect 3764 963 3765 967
rect 3759 962 3765 963
rect 3958 967 3964 968
rect 3958 963 3959 967
rect 3963 966 3964 967
rect 3967 967 3973 968
rect 3967 966 3968 967
rect 3963 964 3968 966
rect 3963 963 3964 964
rect 3958 962 3964 963
rect 3967 963 3968 964
rect 3972 963 3973 967
rect 3967 962 3973 963
rect 1982 958 1988 959
rect 662 954 668 955
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 110 947 116 948
rect 2030 952 2036 953
rect 2030 948 2031 952
rect 2035 948 2036 952
rect 2030 947 2036 948
rect 2223 951 2229 952
rect 2223 947 2224 951
rect 2228 950 2229 951
rect 2271 951 2277 952
rect 2271 950 2272 951
rect 2228 948 2272 950
rect 2228 947 2229 948
rect 2223 946 2229 947
rect 2271 947 2272 948
rect 2276 947 2277 951
rect 2271 946 2277 947
rect 2359 951 2365 952
rect 2359 947 2360 951
rect 2364 950 2365 951
rect 2415 951 2421 952
rect 2415 950 2416 951
rect 2364 948 2416 950
rect 2364 947 2365 948
rect 2359 946 2365 947
rect 2415 947 2416 948
rect 2420 947 2421 951
rect 2415 946 2421 947
rect 2423 951 2429 952
rect 2423 947 2424 951
rect 2428 950 2429 951
rect 2503 951 2509 952
rect 2503 950 2504 951
rect 2428 948 2504 950
rect 2428 947 2429 948
rect 2423 946 2429 947
rect 2503 947 2504 948
rect 2508 947 2509 951
rect 2503 946 2509 947
rect 2663 951 2669 952
rect 2663 947 2664 951
rect 2668 950 2669 951
rect 2743 951 2749 952
rect 2743 950 2744 951
rect 2668 948 2744 950
rect 2668 947 2669 948
rect 2663 946 2669 947
rect 2743 947 2744 948
rect 2748 947 2749 951
rect 2743 946 2749 947
rect 2830 951 2837 952
rect 2830 947 2831 951
rect 2836 947 2837 951
rect 2830 946 2837 947
rect 3007 951 3013 952
rect 3007 947 3008 951
rect 3012 950 3013 951
rect 3024 950 3026 962
rect 3012 948 3026 950
rect 3191 951 3197 952
rect 3012 947 3013 948
rect 3007 946 3013 947
rect 3191 947 3192 951
rect 3196 950 3197 951
rect 3295 951 3301 952
rect 3295 950 3296 951
rect 3196 948 3296 950
rect 3196 947 3197 948
rect 3191 946 3197 947
rect 3295 947 3296 948
rect 3300 947 3301 951
rect 3295 946 3301 947
rect 3383 951 3389 952
rect 3383 947 3384 951
rect 3388 950 3389 951
rect 3495 951 3501 952
rect 3495 950 3496 951
rect 3388 948 3496 950
rect 3388 947 3389 948
rect 3383 946 3389 947
rect 3495 947 3496 948
rect 3500 947 3501 951
rect 3495 946 3501 947
rect 3583 951 3589 952
rect 3583 947 3584 951
rect 3588 950 3589 951
rect 3695 951 3701 952
rect 3695 950 3696 951
rect 3588 948 3696 950
rect 3588 947 3589 948
rect 3583 946 3589 947
rect 3695 947 3696 948
rect 3700 947 3701 951
rect 3695 946 3701 947
rect 3782 951 3789 952
rect 3782 947 3783 951
rect 3788 947 3789 951
rect 3782 946 3789 947
rect 3966 951 3973 952
rect 3966 947 3967 951
rect 3972 947 3973 951
rect 3966 946 3973 947
rect 2150 943 2156 944
rect 2150 939 2151 943
rect 2155 939 2156 943
rect 2150 938 2156 939
rect 2286 943 2292 944
rect 2286 939 2287 943
rect 2291 939 2292 943
rect 2286 938 2292 939
rect 2430 943 2436 944
rect 2430 939 2431 943
rect 2435 939 2436 943
rect 2430 938 2436 939
rect 2590 943 2596 944
rect 2590 939 2591 943
rect 2595 939 2596 943
rect 2590 938 2596 939
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2934 943 2940 944
rect 2934 939 2935 943
rect 2939 939 2940 943
rect 2934 938 2940 939
rect 3118 943 3124 944
rect 3118 939 3119 943
rect 3123 939 3124 943
rect 3118 938 3124 939
rect 3310 943 3316 944
rect 3310 939 3311 943
rect 3315 939 3316 943
rect 3310 938 3316 939
rect 3510 943 3516 944
rect 3510 939 3511 943
rect 3515 939 3516 943
rect 3510 938 3516 939
rect 3710 943 3716 944
rect 3710 939 3711 943
rect 3715 939 3716 943
rect 3710 938 3716 939
rect 3894 943 3900 944
rect 3894 939 3895 943
rect 3899 939 3900 943
rect 3894 938 3900 939
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 2030 935 2036 936
rect 2030 931 2031 935
rect 2035 931 2036 935
rect 2270 935 2276 936
rect 2270 934 2271 935
rect 2201 932 2271 934
rect 110 930 116 931
rect 150 930 156 931
rect 150 926 151 930
rect 155 926 156 930
rect 150 925 156 926
rect 286 930 292 931
rect 286 926 287 930
rect 291 926 292 930
rect 286 925 292 926
rect 470 930 476 931
rect 470 926 471 930
rect 475 926 476 930
rect 470 925 476 926
rect 670 930 676 931
rect 670 926 671 930
rect 675 926 676 930
rect 670 925 676 926
rect 870 930 876 931
rect 870 926 871 930
rect 875 926 876 930
rect 870 925 876 926
rect 1078 930 1084 931
rect 1078 926 1079 930
rect 1083 926 1084 930
rect 1078 925 1084 926
rect 1286 930 1292 931
rect 1286 926 1287 930
rect 1291 926 1292 930
rect 1286 925 1292 926
rect 1494 930 1500 931
rect 1494 926 1495 930
rect 1499 926 1500 930
rect 1494 925 1500 926
rect 1702 930 1708 931
rect 1702 926 1703 930
rect 1707 926 1708 930
rect 1702 925 1708 926
rect 1910 930 1916 931
rect 2030 930 2036 931
rect 2270 931 2271 932
rect 2275 931 2276 935
rect 2670 935 2676 936
rect 2670 934 2671 935
rect 2641 932 2671 934
rect 2270 930 2276 931
rect 2670 931 2671 932
rect 2675 931 2676 935
rect 3055 935 3061 936
rect 3055 934 3056 935
rect 2985 932 3056 934
rect 2670 930 2676 931
rect 3055 931 3056 932
rect 3060 931 3061 935
rect 3214 935 3220 936
rect 3214 934 3215 935
rect 3169 932 3215 934
rect 3055 930 3061 931
rect 3214 931 3215 932
rect 3219 931 3220 935
rect 3958 935 3964 936
rect 3958 934 3959 935
rect 3945 932 3959 934
rect 3214 930 3220 931
rect 3958 931 3959 932
rect 3963 931 3964 935
rect 3958 930 3964 931
rect 1910 926 1911 930
rect 1915 926 1916 930
rect 1910 925 1916 926
rect 2070 924 2076 925
rect 2070 920 2071 924
rect 2075 920 2076 924
rect 2070 919 2076 920
rect 3990 924 3996 925
rect 3990 920 3991 924
rect 3995 920 3996 924
rect 3990 919 3996 920
rect 1215 911 1221 912
rect 1215 907 1216 911
rect 1220 910 1221 911
rect 1502 911 1508 912
rect 1502 910 1503 911
rect 1220 908 1503 910
rect 1220 907 1221 908
rect 1215 906 1221 907
rect 1502 907 1503 908
rect 1507 907 1508 911
rect 1502 906 1508 907
rect 2070 907 2076 908
rect 2070 903 2071 907
rect 2075 903 2076 907
rect 3990 907 3996 908
rect 3990 903 3991 907
rect 3995 903 3996 907
rect 2070 902 2076 903
rect 2150 902 2156 903
rect 2150 898 2151 902
rect 2155 898 2156 902
rect 2150 897 2156 898
rect 2286 902 2292 903
rect 2286 898 2287 902
rect 2291 898 2292 902
rect 2286 897 2292 898
rect 2430 902 2436 903
rect 2430 898 2431 902
rect 2435 898 2436 902
rect 2430 897 2436 898
rect 2590 902 2596 903
rect 2590 898 2591 902
rect 2595 898 2596 902
rect 2590 897 2596 898
rect 2758 902 2764 903
rect 2758 898 2759 902
rect 2763 898 2764 902
rect 2758 897 2764 898
rect 2934 902 2940 903
rect 2934 898 2935 902
rect 2939 898 2940 902
rect 2934 897 2940 898
rect 3118 902 3124 903
rect 3118 898 3119 902
rect 3123 898 3124 902
rect 3118 897 3124 898
rect 3310 902 3316 903
rect 3310 898 3311 902
rect 3315 898 3316 902
rect 3310 897 3316 898
rect 3510 902 3516 903
rect 3510 898 3511 902
rect 3515 898 3516 902
rect 3510 897 3516 898
rect 3710 902 3716 903
rect 3710 898 3711 902
rect 3715 898 3716 902
rect 3710 897 3716 898
rect 3894 902 3900 903
rect 3990 902 3996 903
rect 3894 898 3895 902
rect 3899 898 3900 902
rect 3894 897 3900 898
rect 150 890 156 891
rect 150 886 151 890
rect 155 886 156 890
rect 110 885 116 886
rect 150 885 156 886
rect 318 890 324 891
rect 318 886 319 890
rect 323 886 324 890
rect 318 885 324 886
rect 518 890 524 891
rect 518 886 519 890
rect 523 886 524 890
rect 518 885 524 886
rect 726 890 732 891
rect 726 886 727 890
rect 731 886 732 890
rect 726 885 732 886
rect 934 890 940 891
rect 934 886 935 890
rect 939 886 940 890
rect 934 885 940 886
rect 1142 890 1148 891
rect 1142 886 1143 890
rect 1147 886 1148 890
rect 1142 885 1148 886
rect 1334 890 1340 891
rect 1334 886 1335 890
rect 1339 886 1340 890
rect 1334 885 1340 886
rect 1526 890 1532 891
rect 1526 886 1527 890
rect 1531 886 1532 890
rect 1526 885 1532 886
rect 1718 890 1724 891
rect 1718 886 1719 890
rect 1723 886 1724 890
rect 1718 885 1724 886
rect 1910 890 1916 891
rect 1910 886 1911 890
rect 1915 886 1916 890
rect 1910 885 1916 886
rect 2030 885 2036 886
rect 110 881 111 885
rect 115 881 116 885
rect 110 880 116 881
rect 2030 881 2031 885
rect 2035 881 2036 885
rect 2030 880 2036 881
rect 110 868 116 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 2030 868 2036 869
rect 2030 864 2031 868
rect 2035 864 2036 868
rect 2030 863 2036 864
rect 230 859 236 860
rect 230 858 231 859
rect 201 856 231 858
rect 230 855 231 856
rect 235 855 236 859
rect 230 854 236 855
rect 750 859 756 860
rect 750 855 751 859
rect 755 855 756 859
rect 1215 859 1221 860
rect 1215 858 1216 859
rect 1193 856 1216 858
rect 750 854 756 855
rect 1215 855 1216 856
rect 1220 855 1221 859
rect 1215 854 1221 855
rect 2110 858 2116 859
rect 2110 854 2111 858
rect 2115 854 2116 858
rect 2070 853 2076 854
rect 2110 853 2116 854
rect 2238 858 2244 859
rect 2238 854 2239 858
rect 2243 854 2244 858
rect 2238 853 2244 854
rect 2406 858 2412 859
rect 2406 854 2407 858
rect 2411 854 2412 858
rect 2406 853 2412 854
rect 2574 858 2580 859
rect 2574 854 2575 858
rect 2579 854 2580 858
rect 2574 853 2580 854
rect 2750 858 2756 859
rect 2750 854 2751 858
rect 2755 854 2756 858
rect 2750 853 2756 854
rect 2934 858 2940 859
rect 2934 854 2935 858
rect 2939 854 2940 858
rect 2934 853 2940 854
rect 3118 858 3124 859
rect 3118 854 3119 858
rect 3123 854 3124 858
rect 3118 853 3124 854
rect 3310 858 3316 859
rect 3310 854 3311 858
rect 3315 854 3316 858
rect 3310 853 3316 854
rect 3510 858 3516 859
rect 3510 854 3511 858
rect 3515 854 3516 858
rect 3510 853 3516 854
rect 3710 858 3716 859
rect 3710 854 3711 858
rect 3715 854 3716 858
rect 3710 853 3716 854
rect 3894 858 3900 859
rect 3894 854 3895 858
rect 3899 854 3900 858
rect 3894 853 3900 854
rect 3990 853 3996 854
rect 150 849 156 850
rect 150 845 151 849
rect 155 845 156 849
rect 150 844 156 845
rect 318 849 324 850
rect 318 845 319 849
rect 323 845 324 849
rect 318 844 324 845
rect 518 849 524 850
rect 518 845 519 849
rect 523 845 524 849
rect 518 844 524 845
rect 726 849 732 850
rect 726 845 727 849
rect 731 845 732 849
rect 726 844 732 845
rect 934 849 940 850
rect 934 845 935 849
rect 939 845 940 849
rect 934 844 940 845
rect 1142 849 1148 850
rect 1142 845 1143 849
rect 1147 845 1148 849
rect 1142 844 1148 845
rect 1334 849 1340 850
rect 1334 845 1335 849
rect 1339 845 1340 849
rect 1334 844 1340 845
rect 1526 849 1532 850
rect 1526 845 1527 849
rect 1531 845 1532 849
rect 1526 844 1532 845
rect 1718 849 1724 850
rect 1718 845 1719 849
rect 1723 845 1724 849
rect 1718 844 1724 845
rect 1910 849 1916 850
rect 1910 845 1911 849
rect 1915 845 1916 849
rect 2070 849 2071 853
rect 2075 849 2076 853
rect 2070 848 2076 849
rect 3990 849 3991 853
rect 3995 849 3996 853
rect 3990 848 3996 849
rect 1910 844 1916 845
rect 223 839 229 840
rect 223 835 224 839
rect 228 838 229 839
rect 303 839 309 840
rect 303 838 304 839
rect 228 836 304 838
rect 228 835 229 836
rect 223 834 229 835
rect 303 835 304 836
rect 308 835 309 839
rect 303 834 309 835
rect 391 839 397 840
rect 391 835 392 839
rect 396 838 397 839
rect 503 839 509 840
rect 503 838 504 839
rect 396 836 504 838
rect 396 835 397 836
rect 391 834 397 835
rect 503 835 504 836
rect 508 835 509 839
rect 503 834 509 835
rect 591 839 597 840
rect 591 835 592 839
rect 596 838 597 839
rect 662 839 668 840
rect 662 838 663 839
rect 596 836 663 838
rect 596 835 597 836
rect 591 834 597 835
rect 662 835 663 836
rect 667 835 668 839
rect 662 834 668 835
rect 799 839 805 840
rect 799 835 800 839
rect 804 838 805 839
rect 919 839 925 840
rect 919 838 920 839
rect 804 836 920 838
rect 804 835 805 836
rect 799 834 805 835
rect 919 835 920 836
rect 924 835 925 839
rect 1007 839 1013 840
rect 1007 838 1008 839
rect 919 834 925 835
rect 928 836 1008 838
rect 230 831 236 832
rect 230 827 231 831
rect 235 830 236 831
rect 928 830 930 836
rect 1007 835 1008 836
rect 1012 835 1013 839
rect 1007 834 1013 835
rect 1215 839 1221 840
rect 1215 835 1216 839
rect 1220 838 1221 839
rect 1319 839 1325 840
rect 1319 838 1320 839
rect 1220 836 1320 838
rect 1220 835 1221 836
rect 1215 834 1221 835
rect 1319 835 1320 836
rect 1324 835 1325 839
rect 1319 834 1325 835
rect 1407 839 1413 840
rect 1407 835 1408 839
rect 1412 838 1413 839
rect 1511 839 1517 840
rect 1511 838 1512 839
rect 1412 836 1512 838
rect 1412 835 1413 836
rect 1407 834 1413 835
rect 1511 835 1512 836
rect 1516 835 1517 839
rect 1511 834 1517 835
rect 1599 839 1605 840
rect 1599 835 1600 839
rect 1604 838 1605 839
rect 1703 839 1709 840
rect 1703 838 1704 839
rect 1604 836 1704 838
rect 1604 835 1605 836
rect 1599 834 1605 835
rect 1703 835 1704 836
rect 1708 835 1709 839
rect 1703 834 1709 835
rect 1791 839 1797 840
rect 1791 835 1792 839
rect 1796 838 1797 839
rect 1895 839 1901 840
rect 1895 838 1896 839
rect 1796 836 1896 838
rect 1796 835 1797 836
rect 1791 834 1797 835
rect 1895 835 1896 836
rect 1900 835 1901 839
rect 1895 834 1901 835
rect 1982 839 1989 840
rect 1982 835 1983 839
rect 1988 835 1989 839
rect 1982 834 1989 835
rect 2070 836 2076 837
rect 2070 832 2071 836
rect 2075 832 2076 836
rect 2070 831 2076 832
rect 3990 836 3996 837
rect 3990 832 3991 836
rect 3995 832 3996 836
rect 3990 831 3996 832
rect 235 828 930 830
rect 235 827 236 828
rect 230 826 236 827
rect 2182 827 2188 828
rect 2182 826 2183 827
rect 2161 824 2183 826
rect 2182 823 2183 824
rect 2187 823 2188 827
rect 2558 827 2564 828
rect 2558 826 2559 827
rect 2457 824 2559 826
rect 2182 822 2188 823
rect 2558 823 2559 824
rect 2563 823 2564 827
rect 2734 827 2740 828
rect 2734 826 2735 827
rect 2625 824 2735 826
rect 2558 822 2564 823
rect 2734 823 2735 824
rect 2739 823 2740 827
rect 2830 827 2836 828
rect 2830 826 2831 827
rect 2801 824 2831 826
rect 2734 822 2740 823
rect 2830 823 2831 824
rect 2835 823 2836 827
rect 3494 827 3500 828
rect 3494 826 3495 827
rect 3361 824 3495 826
rect 2830 822 2836 823
rect 3494 823 3495 824
rect 3499 823 3500 827
rect 3694 827 3700 828
rect 3694 826 3695 827
rect 3561 824 3695 826
rect 3494 822 3500 823
rect 3694 823 3695 824
rect 3699 823 3700 827
rect 3782 827 3788 828
rect 3782 826 3783 827
rect 3761 824 3783 826
rect 3694 822 3700 823
rect 3782 823 3783 824
rect 3787 823 3788 827
rect 3966 827 3972 828
rect 3966 826 3967 827
rect 3945 824 3967 826
rect 3782 822 3788 823
rect 3966 823 3967 824
rect 3971 823 3972 827
rect 3966 822 3972 823
rect 2110 817 2116 818
rect 335 815 341 816
rect 335 811 336 815
rect 340 814 341 815
rect 351 815 357 816
rect 351 814 352 815
rect 340 812 352 814
rect 340 811 341 812
rect 335 810 341 811
rect 351 811 352 812
rect 356 811 357 815
rect 351 810 357 811
rect 439 815 445 816
rect 439 811 440 815
rect 444 814 445 815
rect 463 815 469 816
rect 463 814 464 815
rect 444 812 464 814
rect 444 811 445 812
rect 439 810 445 811
rect 463 811 464 812
rect 468 811 469 815
rect 463 810 469 811
rect 551 815 557 816
rect 551 811 552 815
rect 556 814 557 815
rect 575 815 581 816
rect 575 814 576 815
rect 556 812 576 814
rect 556 811 557 812
rect 551 810 557 811
rect 575 811 576 812
rect 580 811 581 815
rect 575 810 581 811
rect 663 815 669 816
rect 663 811 664 815
rect 668 814 669 815
rect 695 815 701 816
rect 695 814 696 815
rect 668 812 696 814
rect 668 811 669 812
rect 663 810 669 811
rect 695 811 696 812
rect 700 811 701 815
rect 695 810 701 811
rect 750 815 756 816
rect 750 811 751 815
rect 755 814 756 815
rect 783 815 789 816
rect 783 814 784 815
rect 755 812 784 814
rect 755 811 756 812
rect 750 810 756 811
rect 783 811 784 812
rect 788 811 789 815
rect 783 810 789 811
rect 927 815 933 816
rect 927 811 928 815
rect 932 814 933 815
rect 1015 815 1021 816
rect 1015 814 1016 815
rect 932 812 1016 814
rect 932 811 933 812
rect 927 810 933 811
rect 1015 811 1016 812
rect 1020 811 1021 815
rect 1015 810 1021 811
rect 1103 815 1109 816
rect 1103 811 1104 815
rect 1108 814 1109 815
rect 1223 815 1229 816
rect 1223 814 1224 815
rect 1108 812 1224 814
rect 1108 811 1109 812
rect 1103 810 1109 811
rect 1223 811 1224 812
rect 1228 811 1229 815
rect 1223 810 1229 811
rect 1311 815 1317 816
rect 1311 811 1312 815
rect 1316 814 1317 815
rect 1455 815 1461 816
rect 1455 814 1456 815
rect 1316 812 1456 814
rect 1316 811 1317 812
rect 1311 810 1317 811
rect 1455 811 1456 812
rect 1460 811 1461 815
rect 1455 810 1461 811
rect 1543 815 1549 816
rect 1543 811 1544 815
rect 1548 814 1549 815
rect 1695 815 1701 816
rect 1695 814 1696 815
rect 1548 812 1696 814
rect 1548 811 1549 812
rect 1543 810 1549 811
rect 1695 811 1696 812
rect 1700 811 1701 815
rect 1695 810 1701 811
rect 1726 815 1732 816
rect 1726 811 1727 815
rect 1731 814 1732 815
rect 1783 815 1789 816
rect 1783 814 1784 815
rect 1731 812 1784 814
rect 1731 811 1732 812
rect 1726 810 1732 811
rect 1783 811 1784 812
rect 1788 811 1789 815
rect 1783 810 1789 811
rect 2007 815 2016 816
rect 2007 811 2008 815
rect 2015 811 2016 815
rect 2110 813 2111 817
rect 2115 813 2116 817
rect 2110 812 2116 813
rect 2238 817 2244 818
rect 2238 813 2239 817
rect 2243 813 2244 817
rect 2238 812 2244 813
rect 2406 817 2412 818
rect 2406 813 2407 817
rect 2411 813 2412 817
rect 2406 812 2412 813
rect 2574 817 2580 818
rect 2574 813 2575 817
rect 2579 813 2580 817
rect 2574 812 2580 813
rect 2750 817 2756 818
rect 2750 813 2751 817
rect 2755 813 2756 817
rect 2750 812 2756 813
rect 2934 817 2940 818
rect 2934 813 2935 817
rect 2939 813 2940 817
rect 3118 817 3124 818
rect 2934 812 2940 813
rect 3055 815 3061 816
rect 2007 810 2016 811
rect 3055 811 3056 815
rect 3060 814 3061 815
rect 3060 812 3114 814
rect 3118 813 3119 817
rect 3123 813 3124 817
rect 3118 812 3124 813
rect 3310 817 3316 818
rect 3310 813 3311 817
rect 3315 813 3316 817
rect 3310 812 3316 813
rect 3510 817 3516 818
rect 3510 813 3511 817
rect 3515 813 3516 817
rect 3510 812 3516 813
rect 3710 817 3716 818
rect 3710 813 3711 817
rect 3715 813 3716 817
rect 3710 812 3716 813
rect 3894 817 3900 818
rect 3894 813 3895 817
rect 3899 813 3900 817
rect 3894 812 3900 813
rect 3060 811 3061 812
rect 3055 810 3061 811
rect 262 807 268 808
rect 262 803 263 807
rect 267 803 268 807
rect 262 802 268 803
rect 366 807 372 808
rect 366 803 367 807
rect 371 803 372 807
rect 366 802 372 803
rect 478 807 484 808
rect 478 803 479 807
rect 483 803 484 807
rect 478 802 484 803
rect 590 807 596 808
rect 590 803 591 807
rect 595 803 596 807
rect 590 802 596 803
rect 710 807 716 808
rect 710 803 711 807
rect 715 803 716 807
rect 710 802 716 803
rect 854 807 860 808
rect 854 803 855 807
rect 859 803 860 807
rect 854 802 860 803
rect 1030 807 1036 808
rect 1030 803 1031 807
rect 1035 803 1036 807
rect 1030 802 1036 803
rect 1238 807 1244 808
rect 1238 803 1239 807
rect 1243 803 1244 807
rect 1238 802 1244 803
rect 1470 807 1476 808
rect 1470 803 1471 807
rect 1475 803 1476 807
rect 1470 802 1476 803
rect 1710 807 1716 808
rect 1710 803 1711 807
rect 1715 803 1716 807
rect 1710 802 1716 803
rect 1934 807 1940 808
rect 1934 803 1935 807
rect 1939 803 1940 807
rect 1934 802 1940 803
rect 2183 807 2189 808
rect 2183 803 2184 807
rect 2188 806 2189 807
rect 2223 807 2229 808
rect 2223 806 2224 807
rect 2188 804 2224 806
rect 2188 803 2189 804
rect 2183 802 2189 803
rect 2223 803 2224 804
rect 2228 803 2229 807
rect 2223 802 2229 803
rect 2270 807 2276 808
rect 2270 803 2271 807
rect 2275 806 2276 807
rect 2311 807 2317 808
rect 2311 806 2312 807
rect 2275 804 2312 806
rect 2275 803 2276 804
rect 2270 802 2276 803
rect 2311 803 2312 804
rect 2316 803 2317 807
rect 2311 802 2317 803
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 806 2460 807
rect 2479 807 2485 808
rect 2479 806 2480 807
rect 2459 804 2480 806
rect 2459 803 2460 804
rect 2454 802 2460 803
rect 2479 803 2480 804
rect 2484 803 2485 807
rect 2479 802 2485 803
rect 2558 807 2564 808
rect 2558 803 2559 807
rect 2563 806 2564 807
rect 2647 807 2653 808
rect 2647 806 2648 807
rect 2563 804 2648 806
rect 2563 803 2564 804
rect 2558 802 2564 803
rect 2647 803 2648 804
rect 2652 803 2653 807
rect 2647 802 2653 803
rect 2734 807 2740 808
rect 2734 803 2735 807
rect 2739 806 2740 807
rect 2823 807 2829 808
rect 2823 806 2824 807
rect 2739 804 2824 806
rect 2739 803 2740 804
rect 2734 802 2740 803
rect 2823 803 2824 804
rect 2828 803 2829 807
rect 2919 807 2925 808
rect 2919 806 2920 807
rect 2823 802 2829 803
rect 2839 804 2920 806
rect 350 799 356 800
rect 350 798 351 799
rect 313 796 351 798
rect 350 795 351 796
rect 355 795 356 799
rect 998 799 1004 800
rect 998 798 999 799
rect 905 796 999 798
rect 350 794 356 795
rect 998 795 999 796
rect 1003 795 1004 799
rect 998 794 1004 795
rect 1926 795 1932 796
rect 1926 791 1927 795
rect 1931 791 1932 795
rect 1926 790 1932 791
rect 2010 795 2016 796
rect 2010 791 2011 795
rect 2015 794 2016 795
rect 2095 795 2101 796
rect 2095 794 2096 795
rect 2015 792 2096 794
rect 2015 791 2016 792
rect 2010 790 2016 791
rect 2095 791 2096 792
rect 2100 791 2101 795
rect 2095 790 2101 791
rect 2182 795 2189 796
rect 2182 791 2183 795
rect 2188 791 2189 795
rect 2182 790 2189 791
rect 2462 795 2469 796
rect 2462 791 2463 795
rect 2468 791 2469 795
rect 2462 790 2469 791
rect 2751 795 2757 796
rect 2751 791 2752 795
rect 2756 794 2757 795
rect 2839 794 2841 804
rect 2919 803 2920 804
rect 2924 803 2925 807
rect 2919 802 2925 803
rect 3007 807 3013 808
rect 3007 803 3008 807
rect 3012 806 3013 807
rect 3103 807 3109 808
rect 3103 806 3104 807
rect 3012 804 3104 806
rect 3012 803 3013 804
rect 3007 802 3013 803
rect 3103 803 3104 804
rect 3108 803 3109 807
rect 3112 806 3114 812
rect 3191 807 3197 808
rect 3191 806 3192 807
rect 3112 804 3192 806
rect 3103 802 3109 803
rect 3191 803 3192 804
rect 3196 803 3197 807
rect 3191 802 3197 803
rect 3270 807 3276 808
rect 3270 803 3271 807
rect 3275 806 3276 807
rect 3383 807 3389 808
rect 3383 806 3384 807
rect 3275 804 3384 806
rect 3275 803 3276 804
rect 3270 802 3276 803
rect 3383 803 3384 804
rect 3388 803 3389 807
rect 3383 802 3389 803
rect 3494 807 3500 808
rect 3494 803 3495 807
rect 3499 806 3500 807
rect 3583 807 3589 808
rect 3583 806 3584 807
rect 3499 804 3584 806
rect 3499 803 3500 804
rect 3494 802 3500 803
rect 3583 803 3584 804
rect 3588 803 3589 807
rect 3583 802 3589 803
rect 3694 807 3700 808
rect 3694 803 3695 807
rect 3699 806 3700 807
rect 3783 807 3789 808
rect 3783 806 3784 807
rect 3699 804 3784 806
rect 3699 803 3700 804
rect 3694 802 3700 803
rect 3783 803 3784 804
rect 3788 803 3789 807
rect 3783 802 3789 803
rect 3958 807 3964 808
rect 3958 803 3959 807
rect 3963 806 3964 807
rect 3967 807 3973 808
rect 3967 806 3968 807
rect 3963 804 3968 806
rect 3963 803 3964 804
rect 3958 802 3964 803
rect 3967 803 3968 804
rect 3972 803 3973 807
rect 3967 802 3973 803
rect 3023 795 3029 796
rect 3023 794 3024 795
rect 2756 792 2841 794
rect 2932 792 3024 794
rect 2756 791 2757 792
rect 2751 790 2757 791
rect 110 788 116 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 2030 788 2036 789
rect 2030 784 2031 788
rect 2035 784 2036 788
rect 2030 783 2036 784
rect 2110 787 2116 788
rect 2110 783 2111 787
rect 2115 783 2116 787
rect 2110 782 2116 783
rect 2390 787 2396 788
rect 2390 783 2391 787
rect 2395 783 2396 787
rect 2390 782 2396 783
rect 2678 787 2684 788
rect 2678 783 2679 787
rect 2683 783 2684 787
rect 2678 782 2684 783
rect 2454 779 2460 780
rect 2454 778 2455 779
rect 2441 776 2455 778
rect 2454 775 2455 776
rect 2459 775 2460 779
rect 2932 778 2934 792
rect 3023 791 3024 792
rect 3028 791 3029 795
rect 3023 790 3029 791
rect 3271 795 3277 796
rect 3271 791 3272 795
rect 3276 794 3277 795
rect 3423 795 3429 796
rect 3423 794 3424 795
rect 3276 792 3424 794
rect 3276 791 3277 792
rect 3271 790 3277 791
rect 3423 791 3424 792
rect 3428 791 3429 795
rect 3423 790 3429 791
rect 3511 795 3517 796
rect 3511 791 3512 795
rect 3516 794 3517 795
rect 3655 795 3661 796
rect 3655 794 3656 795
rect 3516 792 3656 794
rect 3516 791 3517 792
rect 3511 790 3517 791
rect 3655 791 3656 792
rect 3660 791 3661 795
rect 3655 790 3661 791
rect 3743 795 3749 796
rect 3743 791 3744 795
rect 3748 794 3749 795
rect 3822 795 3828 796
rect 3822 794 3823 795
rect 3748 792 3823 794
rect 3748 791 3749 792
rect 3743 790 3749 791
rect 3822 791 3823 792
rect 3827 791 3828 795
rect 3822 790 3828 791
rect 3966 795 3973 796
rect 3966 791 3967 795
rect 3972 791 3973 795
rect 3966 790 3973 791
rect 2950 787 2956 788
rect 2950 783 2951 787
rect 2955 783 2956 787
rect 2950 782 2956 783
rect 3198 787 3204 788
rect 3198 783 3199 787
rect 3203 783 3204 787
rect 3198 782 3204 783
rect 3438 787 3444 788
rect 3438 783 3439 787
rect 3443 783 3444 787
rect 3438 782 3444 783
rect 3670 787 3676 788
rect 3670 783 3671 787
rect 3675 783 3676 787
rect 3670 782 3676 783
rect 3894 787 3900 788
rect 3894 783 3895 787
rect 3899 783 3900 787
rect 3894 782 3900 783
rect 3062 779 3068 780
rect 3062 778 3063 779
rect 2729 776 2934 778
rect 3001 776 3063 778
rect 2454 774 2460 775
rect 3062 775 3063 776
rect 3067 775 3068 779
rect 3270 779 3276 780
rect 3270 778 3271 779
rect 3249 776 3271 778
rect 3062 774 3068 775
rect 3270 775 3271 776
rect 3275 775 3276 779
rect 3270 774 3276 775
rect 3918 775 3924 776
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 2030 771 2036 772
rect 2030 767 2031 771
rect 2035 767 2036 771
rect 3918 771 3919 775
rect 3923 771 3924 775
rect 3918 770 3924 771
rect 110 766 116 767
rect 262 766 268 767
rect 262 762 263 766
rect 267 762 268 766
rect 262 761 268 762
rect 366 766 372 767
rect 366 762 367 766
rect 371 762 372 766
rect 366 761 372 762
rect 478 766 484 767
rect 478 762 479 766
rect 483 762 484 766
rect 478 761 484 762
rect 590 766 596 767
rect 590 762 591 766
rect 595 762 596 766
rect 590 761 596 762
rect 710 766 716 767
rect 710 762 711 766
rect 715 762 716 766
rect 710 761 716 762
rect 854 766 860 767
rect 854 762 855 766
rect 859 762 860 766
rect 854 761 860 762
rect 1030 766 1036 767
rect 1030 762 1031 766
rect 1035 762 1036 766
rect 1030 761 1036 762
rect 1238 766 1244 767
rect 1238 762 1239 766
rect 1243 762 1244 766
rect 1238 761 1244 762
rect 1470 766 1476 767
rect 1470 762 1471 766
rect 1475 762 1476 766
rect 1470 761 1476 762
rect 1710 766 1716 767
rect 1710 762 1711 766
rect 1715 762 1716 766
rect 1710 761 1716 762
rect 1934 766 1940 767
rect 2030 766 2036 767
rect 2070 768 2076 769
rect 1934 762 1935 766
rect 1939 762 1940 766
rect 2070 764 2071 768
rect 2075 764 2076 768
rect 2070 763 2076 764
rect 3990 768 3996 769
rect 3990 764 3991 768
rect 3995 764 3996 768
rect 3990 763 3996 764
rect 1934 761 1940 762
rect 2070 751 2076 752
rect 1078 747 1084 748
rect 1078 743 1079 747
rect 1083 746 1084 747
rect 1726 747 1732 748
rect 1726 746 1727 747
rect 1083 744 1727 746
rect 1083 743 1084 744
rect 1078 742 1084 743
rect 1726 743 1727 744
rect 1731 743 1732 747
rect 2070 747 2071 751
rect 2075 747 2076 751
rect 3990 751 3996 752
rect 3990 747 3991 751
rect 3995 747 3996 751
rect 2070 746 2076 747
rect 2110 746 2116 747
rect 1726 742 1732 743
rect 2110 742 2111 746
rect 2115 742 2116 746
rect 2110 741 2116 742
rect 2390 746 2396 747
rect 2390 742 2391 746
rect 2395 742 2396 746
rect 2390 741 2396 742
rect 2678 746 2684 747
rect 2678 742 2679 746
rect 2683 742 2684 746
rect 2678 741 2684 742
rect 2950 746 2956 747
rect 2950 742 2951 746
rect 2955 742 2956 746
rect 2950 741 2956 742
rect 3198 746 3204 747
rect 3198 742 3199 746
rect 3203 742 3204 746
rect 3198 741 3204 742
rect 3438 746 3444 747
rect 3438 742 3439 746
rect 3443 742 3444 746
rect 3438 741 3444 742
rect 3670 746 3676 747
rect 3670 742 3671 746
rect 3675 742 3676 746
rect 3670 741 3676 742
rect 3894 746 3900 747
rect 3990 746 3996 747
rect 3894 742 3895 746
rect 3899 742 3900 746
rect 3894 741 3900 742
rect 422 730 428 731
rect 422 726 423 730
rect 427 726 428 730
rect 110 725 116 726
rect 422 725 428 726
rect 526 730 532 731
rect 526 726 527 730
rect 531 726 532 730
rect 526 725 532 726
rect 638 730 644 731
rect 638 726 639 730
rect 643 726 644 730
rect 638 725 644 726
rect 758 730 764 731
rect 758 726 759 730
rect 763 726 764 730
rect 758 725 764 726
rect 878 730 884 731
rect 878 726 879 730
rect 883 726 884 730
rect 878 725 884 726
rect 1006 730 1012 731
rect 1006 726 1007 730
rect 1011 726 1012 730
rect 1006 725 1012 726
rect 1142 730 1148 731
rect 1142 726 1143 730
rect 1147 726 1148 730
rect 1142 725 1148 726
rect 1286 730 1292 731
rect 1286 726 1287 730
rect 1291 726 1292 730
rect 1286 725 1292 726
rect 1446 730 1452 731
rect 1446 726 1447 730
rect 1451 726 1452 730
rect 1446 725 1452 726
rect 1614 730 1620 731
rect 1614 726 1615 730
rect 1619 726 1620 730
rect 1614 725 1620 726
rect 1782 730 1788 731
rect 1782 726 1783 730
rect 1787 726 1788 730
rect 1782 725 1788 726
rect 1934 730 1940 731
rect 1934 726 1935 730
rect 1939 726 1940 730
rect 1934 725 1940 726
rect 2030 725 2036 726
rect 110 721 111 725
rect 115 721 116 725
rect 110 720 116 721
rect 2030 721 2031 725
rect 2035 721 2036 725
rect 2030 720 2036 721
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 110 703 116 704
rect 2030 708 2036 709
rect 2030 704 2031 708
rect 2035 704 2036 708
rect 2030 703 2036 704
rect 2110 706 2116 707
rect 2110 702 2111 706
rect 2115 702 2116 706
rect 2070 701 2076 702
rect 2110 701 2116 702
rect 2326 706 2332 707
rect 2326 702 2327 706
rect 2331 702 2332 706
rect 2326 701 2332 702
rect 2550 706 2556 707
rect 2550 702 2551 706
rect 2555 702 2556 706
rect 2550 701 2556 702
rect 2774 706 2780 707
rect 2774 702 2775 706
rect 2779 702 2780 706
rect 2774 701 2780 702
rect 2990 706 2996 707
rect 2990 702 2991 706
rect 2995 702 2996 706
rect 2990 701 2996 702
rect 3206 706 3212 707
rect 3206 702 3207 706
rect 3211 702 3212 706
rect 3206 701 3212 702
rect 3414 706 3420 707
rect 3414 702 3415 706
rect 3419 702 3420 706
rect 3414 701 3420 702
rect 3622 706 3628 707
rect 3622 702 3623 706
rect 3627 702 3628 706
rect 3622 701 3628 702
rect 3830 706 3836 707
rect 3830 702 3831 706
rect 3835 702 3836 706
rect 3830 701 3836 702
rect 3990 701 3996 702
rect 510 699 516 700
rect 510 698 511 699
rect 473 696 511 698
rect 510 695 511 696
rect 515 695 516 699
rect 622 699 628 700
rect 622 698 623 699
rect 577 696 623 698
rect 510 694 516 695
rect 622 695 623 696
rect 627 695 628 699
rect 742 699 748 700
rect 742 698 743 699
rect 689 696 743 698
rect 622 694 628 695
rect 742 695 743 696
rect 747 695 748 699
rect 862 699 868 700
rect 862 698 863 699
rect 809 696 863 698
rect 742 694 748 695
rect 862 695 863 696
rect 867 695 868 699
rect 862 694 868 695
rect 870 699 876 700
rect 870 695 871 699
rect 875 695 876 699
rect 1078 699 1084 700
rect 1078 698 1079 699
rect 1057 696 1079 698
rect 870 694 876 695
rect 1078 695 1079 696
rect 1083 695 1084 699
rect 1890 699 1896 700
rect 1890 698 1891 699
rect 1833 696 1891 698
rect 1078 694 1084 695
rect 1890 695 1891 696
rect 1895 695 1896 699
rect 2062 699 2068 700
rect 2062 698 2063 699
rect 1985 696 2063 698
rect 1890 694 1896 695
rect 2062 695 2063 696
rect 2067 695 2068 699
rect 2070 697 2071 701
rect 2075 697 2076 701
rect 2070 696 2076 697
rect 3990 697 3991 701
rect 3995 697 3996 701
rect 3990 696 3996 697
rect 2062 694 2068 695
rect 422 689 428 690
rect 422 685 423 689
rect 427 685 428 689
rect 422 684 428 685
rect 526 689 532 690
rect 526 685 527 689
rect 531 685 532 689
rect 526 684 532 685
rect 638 689 644 690
rect 638 685 639 689
rect 643 685 644 689
rect 638 684 644 685
rect 758 689 764 690
rect 758 685 759 689
rect 763 685 764 689
rect 758 684 764 685
rect 878 689 884 690
rect 878 685 879 689
rect 883 685 884 689
rect 878 684 884 685
rect 1006 689 1012 690
rect 1006 685 1007 689
rect 1011 685 1012 689
rect 1006 684 1012 685
rect 1142 689 1148 690
rect 1142 685 1143 689
rect 1147 685 1148 689
rect 1142 684 1148 685
rect 1286 689 1292 690
rect 1286 685 1287 689
rect 1291 685 1292 689
rect 1286 684 1292 685
rect 1446 689 1452 690
rect 1446 685 1447 689
rect 1451 685 1452 689
rect 1446 684 1452 685
rect 1614 689 1620 690
rect 1614 685 1615 689
rect 1619 685 1620 689
rect 1614 684 1620 685
rect 1782 689 1788 690
rect 1782 685 1783 689
rect 1787 685 1788 689
rect 1782 684 1788 685
rect 1934 689 1940 690
rect 1934 685 1935 689
rect 1939 685 1940 689
rect 1934 684 1940 685
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 350 679 356 680
rect 350 675 351 679
rect 355 678 356 679
rect 495 679 501 680
rect 495 678 496 679
rect 355 676 496 678
rect 355 675 356 676
rect 350 674 356 675
rect 495 675 496 676
rect 500 675 501 679
rect 495 674 501 675
rect 510 679 516 680
rect 510 675 511 679
rect 515 678 516 679
rect 599 679 605 680
rect 599 678 600 679
rect 515 676 600 678
rect 515 675 516 676
rect 510 674 516 675
rect 599 675 600 676
rect 604 675 605 679
rect 599 674 605 675
rect 622 679 628 680
rect 622 675 623 679
rect 627 678 628 679
rect 711 679 717 680
rect 711 678 712 679
rect 627 676 712 678
rect 627 675 628 676
rect 622 674 628 675
rect 711 675 712 676
rect 716 675 717 679
rect 711 674 717 675
rect 742 679 748 680
rect 742 675 743 679
rect 747 678 748 679
rect 831 679 837 680
rect 831 678 832 679
rect 747 676 832 678
rect 747 675 748 676
rect 742 674 748 675
rect 831 675 832 676
rect 836 675 837 679
rect 831 674 837 675
rect 862 679 868 680
rect 862 675 863 679
rect 867 678 868 679
rect 951 679 957 680
rect 951 678 952 679
rect 867 676 952 678
rect 867 675 868 676
rect 862 674 868 675
rect 951 675 952 676
rect 956 675 957 679
rect 951 674 957 675
rect 1079 679 1085 680
rect 1079 675 1080 679
rect 1084 678 1085 679
rect 1127 679 1133 680
rect 1127 678 1128 679
rect 1084 676 1128 678
rect 1084 675 1085 676
rect 1079 674 1085 675
rect 1127 675 1128 676
rect 1132 675 1133 679
rect 1127 674 1133 675
rect 1215 679 1221 680
rect 1215 675 1216 679
rect 1220 678 1221 679
rect 1271 679 1277 680
rect 1271 678 1272 679
rect 1220 676 1272 678
rect 1220 675 1221 676
rect 1215 674 1221 675
rect 1271 675 1272 676
rect 1276 675 1277 679
rect 1271 674 1277 675
rect 1359 679 1365 680
rect 1359 675 1360 679
rect 1364 678 1365 679
rect 1431 679 1437 680
rect 1431 678 1432 679
rect 1364 676 1432 678
rect 1364 675 1365 676
rect 1359 674 1365 675
rect 1431 675 1432 676
rect 1436 675 1437 679
rect 1431 674 1437 675
rect 1519 679 1525 680
rect 1519 675 1520 679
rect 1524 678 1525 679
rect 1599 679 1605 680
rect 1599 678 1600 679
rect 1524 676 1600 678
rect 1524 675 1525 676
rect 1519 674 1525 675
rect 1599 675 1600 676
rect 1604 675 1605 679
rect 1687 679 1693 680
rect 1687 678 1688 679
rect 1599 674 1605 675
rect 1608 676 1688 678
rect 1246 671 1252 672
rect 678 667 684 668
rect 678 663 679 667
rect 683 666 684 667
rect 1246 667 1247 671
rect 1251 670 1252 671
rect 1608 670 1610 676
rect 1687 675 1688 676
rect 1692 675 1693 679
rect 1687 674 1693 675
rect 1855 679 1861 680
rect 1855 675 1856 679
rect 1860 678 1861 679
rect 1926 679 1932 680
rect 1926 678 1927 679
rect 1860 676 1927 678
rect 1860 675 1861 676
rect 1855 674 1861 675
rect 1926 675 1927 676
rect 1931 675 1932 679
rect 2007 679 2013 680
rect 2070 679 2076 680
rect 3990 684 3996 685
rect 3990 680 3991 684
rect 3995 680 3996 684
rect 3990 679 3996 680
rect 2007 678 2008 679
rect 1926 674 1932 675
rect 1999 676 2008 678
rect 1251 668 1610 670
rect 1890 671 1896 672
rect 1251 667 1252 668
rect 1246 666 1252 667
rect 1890 667 1891 671
rect 1895 670 1896 671
rect 1999 670 2001 676
rect 2007 675 2008 676
rect 2012 675 2013 679
rect 2007 674 2013 675
rect 2182 675 2188 676
rect 2182 674 2183 675
rect 2161 672 2183 674
rect 2182 671 2183 672
rect 2187 671 2188 675
rect 2462 675 2468 676
rect 2462 674 2463 675
rect 2377 672 2463 674
rect 2182 670 2188 671
rect 2462 671 2463 672
rect 2467 671 2468 675
rect 3190 675 3196 676
rect 3190 674 3191 675
rect 3041 672 3191 674
rect 2462 670 2468 671
rect 3190 671 3191 672
rect 3195 671 3196 675
rect 3190 670 3196 671
rect 3198 675 3204 676
rect 3198 671 3199 675
rect 3203 671 3204 675
rect 3546 675 3552 676
rect 3546 674 3547 675
rect 3465 672 3547 674
rect 3198 670 3204 671
rect 3546 671 3547 672
rect 3551 671 3552 675
rect 3546 670 3552 671
rect 3822 675 3828 676
rect 3822 671 3823 675
rect 3827 671 3828 675
rect 3822 670 3828 671
rect 1895 668 2001 670
rect 1895 667 1896 668
rect 1890 666 1896 667
rect 683 664 1026 666
rect 683 663 684 664
rect 678 662 684 663
rect 870 659 876 660
rect 663 655 669 656
rect 663 651 664 655
rect 668 654 669 655
rect 679 655 685 656
rect 679 654 680 655
rect 668 652 680 654
rect 668 651 669 652
rect 663 650 669 651
rect 679 651 680 652
rect 684 651 685 655
rect 679 650 685 651
rect 767 655 773 656
rect 767 651 768 655
rect 772 654 773 655
rect 791 655 797 656
rect 791 654 792 655
rect 772 652 792 654
rect 772 651 773 652
rect 767 650 773 651
rect 791 651 792 652
rect 796 651 797 655
rect 870 655 871 659
rect 875 658 876 659
rect 875 657 885 658
rect 875 656 880 657
rect 875 655 876 656
rect 870 654 876 655
rect 879 653 880 656
rect 884 653 885 657
rect 879 652 885 653
rect 991 655 997 656
rect 791 650 797 651
rect 991 651 992 655
rect 996 654 997 655
rect 1015 655 1021 656
rect 1015 654 1016 655
rect 996 652 1016 654
rect 996 651 997 652
rect 991 650 997 651
rect 1015 651 1016 652
rect 1020 651 1021 655
rect 1024 654 1026 664
rect 2110 665 2116 666
rect 2110 661 2111 665
rect 2115 661 2116 665
rect 2110 660 2116 661
rect 2326 665 2332 666
rect 2326 661 2327 665
rect 2331 661 2332 665
rect 2326 660 2332 661
rect 2550 665 2556 666
rect 2550 661 2551 665
rect 2555 661 2556 665
rect 2550 660 2556 661
rect 2774 665 2780 666
rect 2774 661 2775 665
rect 2779 661 2780 665
rect 2774 660 2780 661
rect 2990 665 2996 666
rect 2990 661 2991 665
rect 2995 661 2996 665
rect 2990 660 2996 661
rect 3206 665 3212 666
rect 3206 661 3207 665
rect 3211 661 3212 665
rect 3206 660 3212 661
rect 3414 665 3420 666
rect 3414 661 3415 665
rect 3419 661 3420 665
rect 3414 660 3420 661
rect 3622 665 3628 666
rect 3622 661 3623 665
rect 3627 661 3628 665
rect 3622 660 3628 661
rect 3830 665 3836 666
rect 3830 661 3831 665
rect 3835 661 3836 665
rect 3830 660 3836 661
rect 1103 655 1109 656
rect 1103 654 1104 655
rect 1024 652 1104 654
rect 1015 650 1021 651
rect 1103 651 1104 652
rect 1108 651 1109 655
rect 1103 650 1109 651
rect 1215 655 1221 656
rect 1215 651 1216 655
rect 1220 654 1221 655
rect 1247 655 1253 656
rect 1247 654 1248 655
rect 1220 652 1248 654
rect 1220 651 1221 652
rect 1215 650 1221 651
rect 1247 651 1248 652
rect 1252 651 1253 655
rect 1247 650 1253 651
rect 1335 655 1341 656
rect 1335 651 1336 655
rect 1340 654 1341 655
rect 1367 655 1373 656
rect 1367 654 1368 655
rect 1340 652 1368 654
rect 1340 651 1341 652
rect 1335 650 1341 651
rect 1367 651 1368 652
rect 1372 651 1373 655
rect 1367 650 1373 651
rect 1455 655 1461 656
rect 1455 651 1456 655
rect 1460 654 1461 655
rect 1487 655 1493 656
rect 1487 654 1488 655
rect 1460 652 1488 654
rect 1460 651 1461 652
rect 1455 650 1461 651
rect 1487 651 1488 652
rect 1492 651 1493 655
rect 1487 650 1493 651
rect 1575 655 1581 656
rect 1575 651 1576 655
rect 1580 654 1581 655
rect 1607 655 1613 656
rect 1607 654 1608 655
rect 1580 652 1608 654
rect 1580 651 1581 652
rect 1575 650 1581 651
rect 1607 651 1608 652
rect 1612 651 1613 655
rect 1695 655 1701 656
rect 1695 654 1696 655
rect 1607 650 1613 651
rect 1616 652 1696 654
rect 590 647 596 648
rect 590 643 591 647
rect 595 643 596 647
rect 590 642 596 643
rect 694 647 700 648
rect 694 643 695 647
rect 699 643 700 647
rect 694 642 700 643
rect 806 647 812 648
rect 806 643 807 647
rect 811 643 812 647
rect 806 642 812 643
rect 918 647 924 648
rect 918 643 919 647
rect 923 643 924 647
rect 918 642 924 643
rect 1030 647 1036 648
rect 1030 643 1031 647
rect 1035 643 1036 647
rect 1030 642 1036 643
rect 1142 647 1148 648
rect 1142 643 1143 647
rect 1147 643 1148 647
rect 1142 642 1148 643
rect 1262 647 1268 648
rect 1262 643 1263 647
rect 1267 643 1268 647
rect 1262 642 1268 643
rect 1382 647 1388 648
rect 1382 643 1383 647
rect 1387 643 1388 647
rect 1382 642 1388 643
rect 1502 647 1508 648
rect 1502 643 1503 647
rect 1507 643 1508 647
rect 1502 642 1508 643
rect 1566 647 1572 648
rect 1566 643 1567 647
rect 1571 646 1572 647
rect 1616 646 1618 652
rect 1695 651 1696 652
rect 1700 651 1701 655
rect 1695 650 1701 651
rect 2062 655 2068 656
rect 2062 651 2063 655
rect 2067 654 2068 655
rect 2183 655 2189 656
rect 2183 654 2184 655
rect 2067 652 2184 654
rect 2067 651 2068 652
rect 2062 650 2068 651
rect 2183 651 2184 652
rect 2188 651 2189 655
rect 2183 650 2189 651
rect 2399 655 2405 656
rect 2399 651 2400 655
rect 2404 654 2405 655
rect 2535 655 2541 656
rect 2535 654 2536 655
rect 2404 652 2536 654
rect 2404 651 2405 652
rect 2399 650 2405 651
rect 2535 651 2536 652
rect 2540 651 2541 655
rect 2535 650 2541 651
rect 2623 655 2629 656
rect 2623 651 2624 655
rect 2628 654 2629 655
rect 2759 655 2765 656
rect 2759 654 2760 655
rect 2628 652 2760 654
rect 2628 651 2629 652
rect 2623 650 2629 651
rect 2759 651 2760 652
rect 2764 651 2765 655
rect 2847 655 2853 656
rect 2847 654 2848 655
rect 2759 650 2765 651
rect 2839 652 2848 654
rect 1571 644 1618 646
rect 1622 647 1628 648
rect 1571 643 1572 644
rect 1566 642 1572 643
rect 1622 643 1623 647
rect 1627 643 1628 647
rect 1622 642 1628 643
rect 2722 647 2728 648
rect 2722 643 2723 647
rect 2727 646 2728 647
rect 2839 646 2841 652
rect 2847 651 2848 652
rect 2852 651 2853 655
rect 2847 650 2853 651
rect 3062 655 3069 656
rect 3062 651 3063 655
rect 3068 651 3069 655
rect 3062 650 3069 651
rect 3190 655 3196 656
rect 3190 651 3191 655
rect 3195 654 3196 655
rect 3279 655 3285 656
rect 3279 654 3280 655
rect 3195 652 3280 654
rect 3195 651 3196 652
rect 3190 650 3196 651
rect 3279 651 3280 652
rect 3284 651 3285 655
rect 3279 650 3285 651
rect 3487 655 3493 656
rect 3487 651 3488 655
rect 3492 654 3493 655
rect 3607 655 3613 656
rect 3607 654 3608 655
rect 3492 652 3608 654
rect 3492 651 3493 652
rect 3487 650 3493 651
rect 3607 651 3608 652
rect 3612 651 3613 655
rect 3607 650 3613 651
rect 3694 655 3701 656
rect 3694 651 3695 655
rect 3700 651 3701 655
rect 3903 655 3909 656
rect 3903 654 3904 655
rect 3694 650 3701 651
rect 3792 652 3904 654
rect 2727 644 2841 646
rect 3110 647 3116 648
rect 2727 643 2728 644
rect 2722 642 2728 643
rect 3110 643 3111 647
rect 3115 646 3116 647
rect 3546 647 3552 648
rect 3115 644 3210 646
rect 3115 643 3116 644
rect 3110 642 3116 643
rect 678 639 684 640
rect 678 638 679 639
rect 641 636 679 638
rect 678 635 679 636
rect 683 635 684 639
rect 1246 639 1252 640
rect 1246 638 1247 639
rect 1193 636 1247 638
rect 678 634 684 635
rect 942 635 948 636
rect 942 631 943 635
rect 947 631 948 635
rect 1246 635 1247 636
rect 1251 635 1252 639
rect 1246 634 1252 635
rect 2182 639 2188 640
rect 2182 635 2183 639
rect 2187 638 2188 639
rect 2199 639 2205 640
rect 2199 638 2200 639
rect 2187 636 2200 638
rect 2187 635 2188 636
rect 2182 634 2188 635
rect 2199 635 2200 636
rect 2204 635 2205 639
rect 2367 639 2373 640
rect 2367 638 2368 639
rect 2199 634 2205 635
rect 2244 636 2368 638
rect 942 630 948 631
rect 2126 631 2132 632
rect 110 628 116 629
rect 110 624 111 628
rect 115 624 116 628
rect 110 623 116 624
rect 2030 628 2036 629
rect 2030 624 2031 628
rect 2035 624 2036 628
rect 2126 627 2127 631
rect 2131 627 2132 631
rect 2126 626 2132 627
rect 2030 623 2036 624
rect 2244 622 2246 636
rect 2367 635 2368 636
rect 2372 635 2373 639
rect 2527 639 2533 640
rect 2527 638 2528 639
rect 2367 634 2373 635
rect 2408 636 2528 638
rect 2294 631 2300 632
rect 2294 627 2295 631
rect 2299 627 2300 631
rect 2294 626 2300 627
rect 2408 622 2410 636
rect 2527 635 2528 636
rect 2532 635 2533 639
rect 2527 634 2533 635
rect 2687 639 2693 640
rect 2687 635 2688 639
rect 2692 638 2693 639
rect 2767 639 2773 640
rect 2767 638 2768 639
rect 2692 636 2768 638
rect 2692 635 2693 636
rect 2687 634 2693 635
rect 2767 635 2768 636
rect 2772 635 2773 639
rect 2767 634 2773 635
rect 2855 639 2861 640
rect 2855 635 2856 639
rect 2860 638 2861 639
rect 2870 639 2876 640
rect 2870 638 2871 639
rect 2860 636 2871 638
rect 2860 635 2861 636
rect 2855 634 2861 635
rect 2870 635 2871 636
rect 2875 635 2876 639
rect 2870 634 2876 635
rect 3023 639 3029 640
rect 3023 635 3024 639
rect 3028 638 3029 639
rect 3111 639 3117 640
rect 3111 638 3112 639
rect 3028 636 3112 638
rect 3028 635 3029 636
rect 3023 634 3029 635
rect 3111 635 3112 636
rect 3116 635 3117 639
rect 3111 634 3117 635
rect 3198 639 3205 640
rect 3198 635 3199 639
rect 3204 635 3205 639
rect 3208 638 3210 644
rect 3546 643 3547 647
rect 3551 646 3552 647
rect 3792 646 3794 652
rect 3903 651 3904 652
rect 3908 651 3909 655
rect 3903 650 3909 651
rect 3551 644 3794 646
rect 3551 643 3552 644
rect 3546 642 3552 643
rect 3918 643 3924 644
rect 3375 639 3381 640
rect 3375 638 3376 639
rect 3208 636 3376 638
rect 3198 634 3205 635
rect 3375 635 3376 636
rect 3380 635 3381 639
rect 3559 639 3565 640
rect 3559 638 3560 639
rect 3375 634 3381 635
rect 3428 636 3560 638
rect 2454 631 2460 632
rect 2454 627 2455 631
rect 2459 627 2460 631
rect 2454 626 2460 627
rect 2614 631 2620 632
rect 2614 627 2615 631
rect 2619 627 2620 631
rect 2614 626 2620 627
rect 2782 631 2788 632
rect 2782 627 2783 631
rect 2787 627 2788 631
rect 2782 626 2788 627
rect 2950 631 2956 632
rect 2950 627 2951 631
rect 2955 627 2956 631
rect 2950 626 2956 627
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 2518 623 2524 624
rect 2518 622 2519 623
rect 2177 620 2246 622
rect 2345 620 2410 622
rect 2505 620 2519 622
rect 2518 619 2519 620
rect 2523 619 2524 623
rect 2722 623 2728 624
rect 2722 622 2723 623
rect 2665 620 2723 622
rect 2518 618 2524 619
rect 2722 619 2723 620
rect 2727 619 2728 623
rect 3110 623 3116 624
rect 3110 622 3111 623
rect 3001 620 3111 622
rect 2722 618 2728 619
rect 3110 619 3111 620
rect 3115 619 3116 623
rect 3428 622 3430 636
rect 3559 635 3560 636
rect 3564 635 3565 639
rect 3559 634 3565 635
rect 3751 639 3757 640
rect 3751 635 3752 639
rect 3756 638 3757 639
rect 3814 639 3820 640
rect 3814 638 3815 639
rect 3756 636 3815 638
rect 3756 635 3757 636
rect 3751 634 3757 635
rect 3814 635 3815 636
rect 3819 635 3820 639
rect 3918 639 3919 643
rect 3923 642 3924 643
rect 3923 641 3954 642
rect 3923 640 3957 641
rect 3923 639 3924 640
rect 3918 638 3924 639
rect 3951 636 3952 640
rect 3956 636 3957 640
rect 3951 635 3957 636
rect 3814 634 3820 635
rect 3486 631 3492 632
rect 3486 627 3487 631
rect 3491 627 3492 631
rect 3486 626 3492 627
rect 3678 631 3684 632
rect 3678 627 3679 631
rect 3683 627 3684 631
rect 3678 626 3684 627
rect 3878 631 3884 632
rect 3878 627 3879 631
rect 3883 627 3884 631
rect 3878 626 3884 627
rect 3353 620 3430 622
rect 3110 618 3116 619
rect 3478 619 3484 620
rect 3478 615 3479 619
rect 3483 615 3484 619
rect 3478 614 3484 615
rect 3694 619 3700 620
rect 3694 615 3695 619
rect 3699 615 3700 619
rect 3694 614 3700 615
rect 3894 619 3900 620
rect 3894 615 3895 619
rect 3899 615 3900 619
rect 3894 614 3900 615
rect 2070 612 2076 613
rect 110 611 116 612
rect 110 607 111 611
rect 115 607 116 611
rect 2030 611 2036 612
rect 2030 607 2031 611
rect 2035 607 2036 611
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 3990 612 3996 613
rect 3990 608 3991 612
rect 3995 608 3996 612
rect 3990 607 3996 608
rect 110 606 116 607
rect 590 606 596 607
rect 590 602 591 606
rect 595 602 596 606
rect 590 601 596 602
rect 694 606 700 607
rect 694 602 695 606
rect 699 602 700 606
rect 694 601 700 602
rect 806 606 812 607
rect 806 602 807 606
rect 811 602 812 606
rect 806 601 812 602
rect 918 606 924 607
rect 918 602 919 606
rect 923 602 924 606
rect 918 601 924 602
rect 1030 606 1036 607
rect 1030 602 1031 606
rect 1035 602 1036 606
rect 1030 601 1036 602
rect 1142 606 1148 607
rect 1142 602 1143 606
rect 1147 602 1148 606
rect 1142 601 1148 602
rect 1262 606 1268 607
rect 1262 602 1263 606
rect 1267 602 1268 606
rect 1262 601 1268 602
rect 1382 606 1388 607
rect 1382 602 1383 606
rect 1387 602 1388 606
rect 1382 601 1388 602
rect 1502 606 1508 607
rect 1502 602 1503 606
rect 1507 602 1508 606
rect 1502 601 1508 602
rect 1622 606 1628 607
rect 2030 606 2036 607
rect 1622 602 1623 606
rect 1627 602 1628 606
rect 1622 601 1628 602
rect 2070 595 2076 596
rect 2070 591 2071 595
rect 2075 591 2076 595
rect 3990 595 3996 596
rect 3990 591 3991 595
rect 3995 591 3996 595
rect 2070 590 2076 591
rect 2126 590 2132 591
rect 2126 586 2127 590
rect 2131 586 2132 590
rect 2126 585 2132 586
rect 2294 590 2300 591
rect 2294 586 2295 590
rect 2299 586 2300 590
rect 2294 585 2300 586
rect 2454 590 2460 591
rect 2454 586 2455 590
rect 2459 586 2460 590
rect 2454 585 2460 586
rect 2614 590 2620 591
rect 2614 586 2615 590
rect 2619 586 2620 590
rect 2614 585 2620 586
rect 2782 590 2788 591
rect 2782 586 2783 590
rect 2787 586 2788 590
rect 2782 585 2788 586
rect 2950 590 2956 591
rect 2950 586 2951 590
rect 2955 586 2956 590
rect 2950 585 2956 586
rect 3126 590 3132 591
rect 3126 586 3127 590
rect 3131 586 3132 590
rect 3126 585 3132 586
rect 3302 590 3308 591
rect 3302 586 3303 590
rect 3307 586 3308 590
rect 3302 585 3308 586
rect 3486 590 3492 591
rect 3486 586 3487 590
rect 3491 586 3492 590
rect 3486 585 3492 586
rect 3678 590 3684 591
rect 3678 586 3679 590
rect 3683 586 3684 590
rect 3678 585 3684 586
rect 3878 590 3884 591
rect 3990 590 3996 591
rect 3878 586 3879 590
rect 3883 586 3884 590
rect 3878 585 3884 586
rect 662 566 668 567
rect 662 562 663 566
rect 667 562 668 566
rect 110 561 116 562
rect 662 561 668 562
rect 774 566 780 567
rect 774 562 775 566
rect 779 562 780 566
rect 774 561 780 562
rect 894 566 900 567
rect 894 562 895 566
rect 899 562 900 566
rect 894 561 900 562
rect 1022 566 1028 567
rect 1022 562 1023 566
rect 1027 562 1028 566
rect 1022 561 1028 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 1302 566 1308 567
rect 1302 562 1303 566
rect 1307 562 1308 566
rect 1302 561 1308 562
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1590 566 1596 567
rect 1590 562 1591 566
rect 1595 562 1596 566
rect 1590 561 1596 562
rect 1734 566 1740 567
rect 1734 562 1735 566
rect 1739 562 1740 566
rect 1734 561 1740 562
rect 1878 566 1884 567
rect 1878 562 1879 566
rect 1883 562 1884 566
rect 1878 561 1884 562
rect 2030 561 2036 562
rect 110 557 111 561
rect 115 557 116 561
rect 110 556 116 557
rect 2030 557 2031 561
rect 2035 557 2036 561
rect 2030 556 2036 557
rect 2302 550 2308 551
rect 2302 546 2303 550
rect 2307 546 2308 550
rect 2070 545 2076 546
rect 2302 545 2308 546
rect 2446 550 2452 551
rect 2446 546 2447 550
rect 2451 546 2452 550
rect 2446 545 2452 546
rect 2590 550 2596 551
rect 2590 546 2591 550
rect 2595 546 2596 550
rect 2590 545 2596 546
rect 2734 550 2740 551
rect 2734 546 2735 550
rect 2739 546 2740 550
rect 2734 545 2740 546
rect 2878 550 2884 551
rect 2878 546 2879 550
rect 2883 546 2884 550
rect 2878 545 2884 546
rect 3030 550 3036 551
rect 3030 546 3031 550
rect 3035 546 3036 550
rect 3030 545 3036 546
rect 3182 550 3188 551
rect 3182 546 3183 550
rect 3187 546 3188 550
rect 3182 545 3188 546
rect 3334 550 3340 551
rect 3334 546 3335 550
rect 3339 546 3340 550
rect 3334 545 3340 546
rect 3494 550 3500 551
rect 3494 546 3495 550
rect 3499 546 3500 550
rect 3494 545 3500 546
rect 3654 550 3660 551
rect 3654 546 3655 550
rect 3659 546 3660 550
rect 3654 545 3660 546
rect 3822 550 3828 551
rect 3822 546 3823 550
rect 3827 546 3828 550
rect 3822 545 3828 546
rect 3990 545 3996 546
rect 110 544 116 545
rect 110 540 111 544
rect 115 540 116 544
rect 110 539 116 540
rect 2030 544 2036 545
rect 2030 540 2031 544
rect 2035 540 2036 544
rect 2070 541 2071 545
rect 2075 541 2076 545
rect 2070 540 2076 541
rect 3990 541 3991 545
rect 3995 541 3996 545
rect 3990 540 3996 541
rect 2030 539 2036 540
rect 743 535 749 536
rect 743 534 744 535
rect 713 532 744 534
rect 743 531 744 532
rect 748 531 749 535
rect 878 535 884 536
rect 878 534 879 535
rect 825 532 879 534
rect 743 530 749 531
rect 878 531 879 532
rect 883 531 884 535
rect 1103 535 1109 536
rect 1103 534 1104 535
rect 1073 532 1104 534
rect 878 530 884 531
rect 1103 531 1104 532
rect 1108 531 1109 535
rect 1266 535 1272 536
rect 1266 534 1267 535
rect 1209 532 1267 534
rect 1103 530 1109 531
rect 1266 531 1267 532
rect 1271 531 1272 535
rect 1266 530 1272 531
rect 1326 535 1332 536
rect 1326 531 1327 535
rect 1331 531 1332 535
rect 1566 535 1572 536
rect 1566 534 1567 535
rect 1497 532 1567 534
rect 1326 530 1332 531
rect 1566 531 1567 532
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 2070 528 2076 529
rect 662 525 668 526
rect 662 521 663 525
rect 667 521 668 525
rect 662 520 668 521
rect 774 525 780 526
rect 774 521 775 525
rect 779 521 780 525
rect 774 520 780 521
rect 894 525 900 526
rect 894 521 895 525
rect 899 521 900 525
rect 894 520 900 521
rect 1022 525 1028 526
rect 1022 521 1023 525
rect 1027 521 1028 525
rect 1022 520 1028 521
rect 1158 525 1164 526
rect 1158 521 1159 525
rect 1163 521 1164 525
rect 1158 520 1164 521
rect 1302 525 1308 526
rect 1302 521 1303 525
rect 1307 521 1308 525
rect 1302 520 1308 521
rect 1446 525 1452 526
rect 1446 521 1447 525
rect 1451 521 1452 525
rect 1446 520 1452 521
rect 1590 525 1596 526
rect 1590 521 1591 525
rect 1595 521 1596 525
rect 1590 520 1596 521
rect 1734 525 1740 526
rect 1734 521 1735 525
rect 1739 521 1740 525
rect 1734 520 1740 521
rect 1878 525 1884 526
rect 1878 521 1879 525
rect 1883 521 1884 525
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2070 523 2076 524
rect 3990 528 3996 529
rect 3990 524 3991 528
rect 3995 524 3996 528
rect 3990 523 3996 524
rect 1878 520 1884 521
rect 2430 519 2436 520
rect 2430 518 2431 519
rect 2353 516 2431 518
rect 735 515 741 516
rect 735 511 736 515
rect 740 514 741 515
rect 823 515 829 516
rect 823 514 824 515
rect 740 512 824 514
rect 740 511 741 512
rect 735 510 741 511
rect 823 511 824 512
rect 828 511 829 515
rect 823 510 829 511
rect 847 515 853 516
rect 847 511 848 515
rect 852 514 853 515
rect 879 515 885 516
rect 879 514 880 515
rect 852 512 880 514
rect 852 511 853 512
rect 847 510 853 511
rect 879 511 880 512
rect 884 511 885 515
rect 879 510 885 511
rect 942 515 948 516
rect 942 511 943 515
rect 947 514 948 515
rect 967 515 973 516
rect 967 514 968 515
rect 947 512 968 514
rect 947 511 948 512
rect 942 510 948 511
rect 967 511 968 512
rect 972 511 973 515
rect 1095 515 1101 516
rect 1095 514 1096 515
rect 967 510 973 511
rect 976 512 1096 514
rect 878 507 884 508
rect 878 503 879 507
rect 883 506 884 507
rect 976 506 978 512
rect 1095 511 1096 512
rect 1100 511 1101 515
rect 1095 510 1101 511
rect 1103 515 1109 516
rect 1103 511 1104 515
rect 1108 514 1109 515
rect 1231 515 1237 516
rect 1231 514 1232 515
rect 1108 512 1232 514
rect 1108 511 1109 512
rect 1103 510 1109 511
rect 1231 511 1232 512
rect 1236 511 1237 515
rect 1231 510 1237 511
rect 1266 515 1272 516
rect 1266 511 1267 515
rect 1271 514 1272 515
rect 1375 515 1381 516
rect 1375 514 1376 515
rect 1271 512 1376 514
rect 1271 511 1272 512
rect 1266 510 1272 511
rect 1375 511 1376 512
rect 1380 511 1381 515
rect 1375 510 1381 511
rect 1519 515 1525 516
rect 1519 511 1520 515
rect 1524 514 1525 515
rect 1575 515 1581 516
rect 1575 514 1576 515
rect 1524 512 1576 514
rect 1524 511 1525 512
rect 1519 510 1525 511
rect 1575 511 1576 512
rect 1580 511 1581 515
rect 1575 510 1581 511
rect 1663 515 1669 516
rect 1663 511 1664 515
rect 1668 514 1669 515
rect 1719 515 1725 516
rect 1719 514 1720 515
rect 1668 512 1720 514
rect 1668 511 1669 512
rect 1663 510 1669 511
rect 1719 511 1720 512
rect 1724 511 1725 515
rect 1719 510 1725 511
rect 1807 515 1813 516
rect 1807 511 1808 515
rect 1812 514 1813 515
rect 1863 515 1869 516
rect 1863 514 1864 515
rect 1812 512 1864 514
rect 1812 511 1813 512
rect 1807 510 1813 511
rect 1863 511 1864 512
rect 1868 511 1869 515
rect 1863 510 1869 511
rect 1950 515 1957 516
rect 1950 511 1951 515
rect 1956 511 1957 515
rect 2430 515 2431 516
rect 2435 515 2436 519
rect 2718 519 2724 520
rect 2718 518 2719 519
rect 2641 516 2719 518
rect 2430 514 2436 515
rect 2718 515 2719 516
rect 2723 515 2724 519
rect 2806 519 2812 520
rect 2806 518 2807 519
rect 2785 516 2807 518
rect 2718 514 2724 515
rect 2806 515 2807 516
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 2870 519 2876 520
rect 2870 515 2871 519
rect 2875 515 2876 519
rect 3166 519 3172 520
rect 3166 518 3167 519
rect 3081 516 3167 518
rect 2870 514 2876 515
rect 3166 515 3167 516
rect 3171 515 3172 519
rect 3583 519 3589 520
rect 3583 518 3584 519
rect 3545 516 3584 518
rect 3166 514 3172 515
rect 3583 515 3584 516
rect 3588 515 3589 519
rect 3814 519 3820 520
rect 3705 516 3722 518
rect 3583 514 3589 515
rect 3718 515 3724 516
rect 1950 510 1957 511
rect 3718 511 3719 515
rect 3723 511 3724 515
rect 3814 515 3815 519
rect 3819 515 3820 519
rect 3814 514 3820 515
rect 3718 510 3724 511
rect 883 504 978 506
rect 2302 509 2308 510
rect 2302 505 2303 509
rect 2307 505 2308 509
rect 2302 504 2308 505
rect 2446 509 2452 510
rect 2446 505 2447 509
rect 2451 505 2452 509
rect 2446 504 2452 505
rect 2590 509 2596 510
rect 2590 505 2591 509
rect 2595 505 2596 509
rect 2590 504 2596 505
rect 2734 509 2740 510
rect 2734 505 2735 509
rect 2739 505 2740 509
rect 2734 504 2740 505
rect 2878 509 2884 510
rect 2878 505 2879 509
rect 2883 505 2884 509
rect 2878 504 2884 505
rect 3030 509 3036 510
rect 3030 505 3031 509
rect 3035 505 3036 509
rect 3030 504 3036 505
rect 3182 509 3188 510
rect 3182 505 3183 509
rect 3187 505 3188 509
rect 3182 504 3188 505
rect 3334 509 3340 510
rect 3334 505 3335 509
rect 3339 505 3340 509
rect 3334 504 3340 505
rect 3494 509 3500 510
rect 3494 505 3495 509
rect 3499 505 3500 509
rect 3494 504 3500 505
rect 3654 509 3660 510
rect 3654 505 3655 509
rect 3659 505 3660 509
rect 3654 504 3660 505
rect 3822 509 3828 510
rect 3822 505 3823 509
rect 3827 505 3828 509
rect 3822 504 3828 505
rect 883 503 884 504
rect 878 502 884 503
rect 2375 499 2381 500
rect 2375 495 2376 499
rect 2380 498 2381 499
rect 2431 499 2437 500
rect 2431 498 2432 499
rect 2380 496 2432 498
rect 2380 495 2381 496
rect 2375 494 2381 495
rect 2431 495 2432 496
rect 2436 495 2437 499
rect 2431 494 2437 495
rect 2518 499 2525 500
rect 2518 495 2519 499
rect 2524 495 2525 499
rect 2663 499 2669 500
rect 2663 498 2664 499
rect 2518 494 2525 495
rect 2528 496 2664 498
rect 2430 491 2436 492
rect 607 487 613 488
rect 607 483 608 487
rect 612 486 613 487
rect 623 487 629 488
rect 623 486 624 487
rect 612 484 624 486
rect 612 483 613 484
rect 607 482 613 483
rect 623 483 624 484
rect 628 483 629 487
rect 623 482 629 483
rect 711 487 717 488
rect 711 483 712 487
rect 716 486 717 487
rect 727 487 733 488
rect 727 486 728 487
rect 716 484 728 486
rect 716 483 717 484
rect 711 482 717 483
rect 727 483 728 484
rect 732 483 733 487
rect 727 482 733 483
rect 743 487 749 488
rect 743 483 744 487
rect 748 486 749 487
rect 815 487 821 488
rect 815 486 816 487
rect 748 484 816 486
rect 748 483 749 484
rect 743 482 749 483
rect 815 483 816 484
rect 820 483 821 487
rect 815 482 821 483
rect 823 487 829 488
rect 823 483 824 487
rect 828 486 829 487
rect 831 487 837 488
rect 831 486 832 487
rect 828 484 832 486
rect 828 483 829 484
rect 823 482 829 483
rect 831 483 832 484
rect 836 483 837 487
rect 831 482 837 483
rect 919 487 925 488
rect 919 483 920 487
rect 924 486 925 487
rect 951 487 957 488
rect 951 486 952 487
rect 924 484 952 486
rect 924 483 925 484
rect 919 482 925 483
rect 951 483 952 484
rect 956 483 957 487
rect 951 482 957 483
rect 1038 487 1045 488
rect 1038 483 1039 487
rect 1044 483 1045 487
rect 1038 482 1045 483
rect 1175 487 1181 488
rect 1175 483 1176 487
rect 1180 486 1181 487
rect 1239 487 1245 488
rect 1239 486 1240 487
rect 1180 484 1240 486
rect 1180 483 1181 484
rect 1175 482 1181 483
rect 1239 483 1240 484
rect 1244 483 1245 487
rect 1239 482 1245 483
rect 1326 487 1333 488
rect 1326 483 1327 487
rect 1332 483 1333 487
rect 1326 482 1333 483
rect 1487 487 1493 488
rect 1487 483 1488 487
rect 1492 486 1493 487
rect 1575 487 1581 488
rect 1575 486 1576 487
rect 1492 484 1576 486
rect 1492 483 1493 484
rect 1487 482 1493 483
rect 1575 483 1576 484
rect 1580 483 1581 487
rect 1575 482 1581 483
rect 1598 487 1604 488
rect 1598 483 1599 487
rect 1603 486 1604 487
rect 1663 487 1669 488
rect 1663 486 1664 487
rect 1603 484 1664 486
rect 1603 483 1604 484
rect 1598 482 1604 483
rect 1663 483 1664 484
rect 1668 483 1669 487
rect 1663 482 1669 483
rect 1846 487 1853 488
rect 1846 483 1847 487
rect 1852 483 1853 487
rect 2007 487 2013 488
rect 2007 486 2008 487
rect 1846 482 1853 483
rect 1884 484 2008 486
rect 534 479 540 480
rect 534 475 535 479
rect 539 475 540 479
rect 534 474 540 475
rect 638 479 644 480
rect 638 475 639 479
rect 643 475 644 479
rect 638 474 644 475
rect 742 479 748 480
rect 742 475 743 479
rect 747 475 748 479
rect 742 474 748 475
rect 846 479 852 480
rect 846 475 847 479
rect 851 475 852 479
rect 846 474 852 475
rect 966 479 972 480
rect 966 475 967 479
rect 971 475 972 479
rect 966 474 972 475
rect 1102 479 1108 480
rect 1102 475 1103 479
rect 1107 475 1108 479
rect 1102 474 1108 475
rect 1254 479 1260 480
rect 1254 475 1255 479
rect 1259 475 1260 479
rect 1254 474 1260 475
rect 1414 479 1420 480
rect 1414 475 1415 479
rect 1419 475 1420 479
rect 1414 474 1420 475
rect 1590 479 1596 480
rect 1590 475 1591 479
rect 1595 475 1596 479
rect 1590 474 1596 475
rect 1774 479 1780 480
rect 1774 475 1775 479
rect 1779 475 1780 479
rect 1774 474 1780 475
rect 1238 471 1244 472
rect 1238 470 1239 471
rect 1153 468 1239 470
rect 558 467 564 468
rect 558 463 559 467
rect 563 463 564 467
rect 1238 467 1239 468
rect 1243 467 1244 471
rect 1884 470 1886 484
rect 2007 483 2008 484
rect 2012 483 2013 487
rect 2430 487 2431 491
rect 2435 490 2436 491
rect 2528 490 2530 496
rect 2663 495 2664 496
rect 2668 495 2669 499
rect 2663 494 2669 495
rect 2718 499 2724 500
rect 2718 495 2719 499
rect 2723 498 2724 499
rect 2807 499 2813 500
rect 2807 498 2808 499
rect 2723 496 2808 498
rect 2723 495 2724 496
rect 2718 494 2724 495
rect 2807 495 2808 496
rect 2812 495 2813 499
rect 2807 494 2813 495
rect 2951 499 2960 500
rect 2951 495 2952 499
rect 2959 495 2960 499
rect 2951 494 2960 495
rect 3103 499 3109 500
rect 3103 495 3104 499
rect 3108 498 3109 499
rect 3167 499 3173 500
rect 3167 498 3168 499
rect 3108 496 3168 498
rect 3108 495 3109 496
rect 3103 494 3109 495
rect 3167 495 3168 496
rect 3172 495 3173 499
rect 3167 494 3173 495
rect 3255 499 3261 500
rect 3255 495 3256 499
rect 3260 498 3261 499
rect 3319 499 3325 500
rect 3319 498 3320 499
rect 3260 496 3320 498
rect 3260 495 3261 496
rect 3255 494 3261 495
rect 3319 495 3320 496
rect 3324 495 3325 499
rect 3319 494 3325 495
rect 3407 499 3413 500
rect 3407 495 3408 499
rect 3412 498 3413 499
rect 3478 499 3484 500
rect 3478 498 3479 499
rect 3412 496 3479 498
rect 3412 495 3413 496
rect 3407 494 3413 495
rect 3478 495 3479 496
rect 3483 495 3484 499
rect 3478 494 3484 495
rect 3566 499 3573 500
rect 3566 495 3567 499
rect 3572 495 3573 499
rect 3566 494 3573 495
rect 3583 499 3589 500
rect 3583 495 3584 499
rect 3588 498 3589 499
rect 3727 499 3733 500
rect 3727 498 3728 499
rect 3588 496 3728 498
rect 3588 495 3589 496
rect 3583 494 3589 495
rect 3727 495 3728 496
rect 3732 495 3733 499
rect 3727 494 3733 495
rect 3894 499 3901 500
rect 3894 495 3895 499
rect 3900 495 3901 499
rect 3894 494 3901 495
rect 2435 488 2530 490
rect 2435 487 2436 488
rect 2430 486 2436 487
rect 2598 487 2604 488
rect 2007 482 2013 483
rect 2598 483 2599 487
rect 2603 486 2604 487
rect 2603 484 2841 486
rect 2603 483 2604 484
rect 2598 482 2604 483
rect 1934 479 1940 480
rect 1934 475 1935 479
rect 1939 475 1940 479
rect 1934 474 1940 475
rect 2583 479 2589 480
rect 2583 475 2584 479
rect 2588 478 2589 479
rect 2599 479 2605 480
rect 2599 478 2600 479
rect 2588 476 2600 478
rect 2588 475 2589 476
rect 2583 474 2589 475
rect 2599 475 2600 476
rect 2604 475 2605 479
rect 2599 474 2605 475
rect 2687 479 2693 480
rect 2687 475 2688 479
rect 2692 478 2693 479
rect 2719 479 2725 480
rect 2719 478 2720 479
rect 2692 476 2720 478
rect 2692 475 2693 476
rect 2687 474 2693 475
rect 2719 475 2720 476
rect 2724 475 2725 479
rect 2719 474 2725 475
rect 2806 479 2813 480
rect 2806 475 2807 479
rect 2812 475 2813 479
rect 2839 478 2841 484
rect 2935 479 2941 480
rect 2935 478 2936 479
rect 2839 476 2936 478
rect 2806 474 2813 475
rect 2935 475 2936 476
rect 2940 475 2941 479
rect 2935 474 2941 475
rect 2954 479 2960 480
rect 2954 475 2955 479
rect 2959 478 2960 479
rect 2991 479 2997 480
rect 2991 478 2992 479
rect 2959 476 2992 478
rect 2959 475 2960 476
rect 2954 474 2960 475
rect 2991 475 2992 476
rect 2996 475 2997 479
rect 2991 474 2997 475
rect 3079 479 3085 480
rect 3079 475 3080 479
rect 3084 478 3085 479
rect 3143 479 3149 480
rect 3143 478 3144 479
rect 3084 476 3144 478
rect 3084 475 3085 476
rect 3079 474 3085 475
rect 3143 475 3144 476
rect 3148 475 3149 479
rect 3143 474 3149 475
rect 3231 479 3237 480
rect 3231 475 3232 479
rect 3236 478 3237 479
rect 3303 479 3309 480
rect 3303 478 3304 479
rect 3236 476 3304 478
rect 3236 475 3237 476
rect 3231 474 3237 475
rect 3303 475 3304 476
rect 3308 475 3309 479
rect 3303 474 3309 475
rect 3390 479 3397 480
rect 3390 475 3391 479
rect 3396 475 3397 479
rect 3390 474 3397 475
rect 3551 479 3557 480
rect 3551 475 3552 479
rect 3556 478 3557 479
rect 3631 479 3637 480
rect 3631 478 3632 479
rect 3556 476 3632 478
rect 3556 475 3557 476
rect 3551 474 3557 475
rect 3631 475 3632 476
rect 3636 475 3637 479
rect 3631 474 3637 475
rect 3718 479 3725 480
rect 3718 475 3719 479
rect 3724 475 3725 479
rect 3718 474 3725 475
rect 3838 479 3844 480
rect 3838 475 3839 479
rect 3843 478 3844 479
rect 3895 479 3901 480
rect 3895 478 3896 479
rect 3843 476 3896 478
rect 3843 475 3844 476
rect 3838 474 3844 475
rect 3895 475 3896 476
rect 3900 475 3901 479
rect 3895 474 3901 475
rect 1825 468 1886 470
rect 2510 471 2516 472
rect 1238 466 1244 467
rect 1406 467 1412 468
rect 558 462 564 463
rect 1406 463 1407 467
rect 1411 463 1412 467
rect 1406 462 1412 463
rect 1950 467 1956 468
rect 1950 463 1951 467
rect 1955 463 1956 467
rect 2510 467 2511 471
rect 2515 467 2516 471
rect 2510 466 2516 467
rect 2614 471 2620 472
rect 2614 467 2615 471
rect 2619 467 2620 471
rect 2614 466 2620 467
rect 2734 471 2740 472
rect 2734 467 2735 471
rect 2739 467 2740 471
rect 2734 466 2740 467
rect 2862 471 2868 472
rect 2862 467 2863 471
rect 2867 467 2868 471
rect 2862 466 2868 467
rect 3006 471 3012 472
rect 3006 467 3007 471
rect 3011 467 3012 471
rect 3006 466 3012 467
rect 3158 471 3164 472
rect 3158 467 3159 471
rect 3163 467 3164 471
rect 3158 466 3164 467
rect 3318 471 3324 472
rect 3318 467 3319 471
rect 3323 467 3324 471
rect 3318 466 3324 467
rect 3478 471 3484 472
rect 3478 467 3479 471
rect 3483 467 3484 471
rect 3478 466 3484 467
rect 3646 471 3652 472
rect 3646 467 3647 471
rect 3651 467 3652 471
rect 3646 466 3652 467
rect 3822 471 3828 472
rect 3822 467 3823 471
rect 3827 467 3828 471
rect 3822 466 3828 467
rect 1950 462 1956 463
rect 2598 463 2604 464
rect 2598 462 2599 463
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 110 455 116 456
rect 2030 460 2036 461
rect 2561 460 2599 462
rect 2030 456 2031 460
rect 2035 456 2036 460
rect 2598 459 2599 460
rect 2603 459 2604 463
rect 3586 463 3592 464
rect 3586 462 3587 463
rect 3529 460 3587 462
rect 2598 458 2604 459
rect 2886 459 2892 460
rect 2030 455 2036 456
rect 2886 455 2887 459
rect 2891 455 2892 459
rect 3586 459 3587 460
rect 3591 459 3592 463
rect 3958 463 3964 464
rect 3958 462 3959 463
rect 3873 460 3959 462
rect 3586 458 3592 459
rect 3958 459 3959 460
rect 3963 459 3964 463
rect 3958 458 3964 459
rect 2886 454 2892 455
rect 2070 452 2076 453
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 3990 452 3996 453
rect 3990 448 3991 452
rect 3995 448 3996 452
rect 3990 447 3996 448
rect 110 443 116 444
rect 110 439 111 443
rect 115 439 116 443
rect 2030 443 2036 444
rect 2030 439 2031 443
rect 2035 439 2036 443
rect 110 438 116 439
rect 534 438 540 439
rect 534 434 535 438
rect 539 434 540 438
rect 534 433 540 434
rect 638 438 644 439
rect 638 434 639 438
rect 643 434 644 438
rect 638 433 644 434
rect 742 438 748 439
rect 742 434 743 438
rect 747 434 748 438
rect 742 433 748 434
rect 846 438 852 439
rect 846 434 847 438
rect 851 434 852 438
rect 846 433 852 434
rect 966 438 972 439
rect 966 434 967 438
rect 971 434 972 438
rect 966 433 972 434
rect 1102 438 1108 439
rect 1102 434 1103 438
rect 1107 434 1108 438
rect 1102 433 1108 434
rect 1254 438 1260 439
rect 1254 434 1255 438
rect 1259 434 1260 438
rect 1254 433 1260 434
rect 1414 438 1420 439
rect 1414 434 1415 438
rect 1419 434 1420 438
rect 1414 433 1420 434
rect 1590 438 1596 439
rect 1590 434 1591 438
rect 1595 434 1596 438
rect 1590 433 1596 434
rect 1774 438 1780 439
rect 1774 434 1775 438
rect 1779 434 1780 438
rect 1774 433 1780 434
rect 1934 438 1940 439
rect 2030 438 2036 439
rect 1934 434 1935 438
rect 1939 434 1940 438
rect 1934 433 1940 434
rect 2070 435 2076 436
rect 2070 431 2071 435
rect 2075 431 2076 435
rect 3990 435 3996 436
rect 3990 431 3991 435
rect 3995 431 3996 435
rect 2070 430 2076 431
rect 2510 430 2516 431
rect 2510 426 2511 430
rect 2515 426 2516 430
rect 2510 425 2516 426
rect 2614 430 2620 431
rect 2614 426 2615 430
rect 2619 426 2620 430
rect 2614 425 2620 426
rect 2734 430 2740 431
rect 2734 426 2735 430
rect 2739 426 2740 430
rect 2734 425 2740 426
rect 2862 430 2868 431
rect 2862 426 2863 430
rect 2867 426 2868 430
rect 2862 425 2868 426
rect 3006 430 3012 431
rect 3006 426 3007 430
rect 3011 426 3012 430
rect 3006 425 3012 426
rect 3158 430 3164 431
rect 3158 426 3159 430
rect 3163 426 3164 430
rect 3158 425 3164 426
rect 3318 430 3324 431
rect 3318 426 3319 430
rect 3323 426 3324 430
rect 3318 425 3324 426
rect 3478 430 3484 431
rect 3478 426 3479 430
rect 3483 426 3484 430
rect 3478 425 3484 426
rect 3646 430 3652 431
rect 3646 426 3647 430
rect 3651 426 3652 430
rect 3646 425 3652 426
rect 3822 430 3828 431
rect 3990 430 3996 431
rect 3822 426 3823 430
rect 3827 426 3828 430
rect 3822 425 3828 426
rect 3103 415 3109 416
rect 3103 411 3104 415
rect 3108 414 3109 415
rect 3390 415 3396 416
rect 3390 414 3391 415
rect 3108 412 3391 414
rect 3108 411 3109 412
rect 3103 410 3109 411
rect 3390 411 3391 412
rect 3395 411 3396 415
rect 3390 410 3396 411
rect 3586 403 3592 404
rect 494 402 500 403
rect 494 398 495 402
rect 499 398 500 402
rect 110 397 116 398
rect 494 397 500 398
rect 630 402 636 403
rect 630 398 631 402
rect 635 398 636 402
rect 630 397 636 398
rect 766 402 772 403
rect 766 398 767 402
rect 771 398 772 402
rect 766 397 772 398
rect 910 402 916 403
rect 910 398 911 402
rect 915 398 916 402
rect 910 397 916 398
rect 1046 402 1052 403
rect 1046 398 1047 402
rect 1051 398 1052 402
rect 1046 397 1052 398
rect 1182 402 1188 403
rect 1182 398 1183 402
rect 1187 398 1188 402
rect 1182 397 1188 398
rect 1318 402 1324 403
rect 1318 398 1319 402
rect 1323 398 1324 402
rect 1318 397 1324 398
rect 1446 402 1452 403
rect 1446 398 1447 402
rect 1451 398 1452 402
rect 1446 397 1452 398
rect 1574 402 1580 403
rect 1574 398 1575 402
rect 1579 398 1580 402
rect 1574 397 1580 398
rect 1702 402 1708 403
rect 1702 398 1703 402
rect 1707 398 1708 402
rect 1702 397 1708 398
rect 1830 402 1836 403
rect 1830 398 1831 402
rect 1835 398 1836 402
rect 1830 397 1836 398
rect 1934 402 1940 403
rect 1934 398 1935 402
rect 1939 398 1940 402
rect 3586 399 3587 403
rect 3591 402 3592 403
rect 3782 403 3788 404
rect 3782 402 3783 403
rect 3591 400 3783 402
rect 3591 399 3592 400
rect 3586 398 3592 399
rect 3782 399 3783 400
rect 3787 399 3788 403
rect 3782 398 3788 399
rect 1934 397 1940 398
rect 2030 397 2036 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2590 386 2596 387
rect 2590 382 2591 386
rect 2595 382 2596 386
rect 2070 381 2076 382
rect 2590 381 2596 382
rect 2694 386 2700 387
rect 2694 382 2695 386
rect 2699 382 2700 386
rect 2694 381 2700 382
rect 2814 386 2820 387
rect 2814 382 2815 386
rect 2819 382 2820 386
rect 2814 381 2820 382
rect 2958 386 2964 387
rect 2958 382 2959 386
rect 2963 382 2964 386
rect 2958 381 2964 382
rect 3118 386 3124 387
rect 3118 382 3119 386
rect 3123 382 3124 386
rect 3118 381 3124 382
rect 3302 386 3308 387
rect 3302 382 3303 386
rect 3307 382 3308 386
rect 3302 381 3308 382
rect 3502 386 3508 387
rect 3502 382 3503 386
rect 3507 382 3508 386
rect 3502 381 3508 382
rect 3710 386 3716 387
rect 3710 382 3711 386
rect 3715 382 3716 386
rect 3710 381 3716 382
rect 3894 386 3900 387
rect 3894 382 3895 386
rect 3899 382 3900 386
rect 3894 381 3900 382
rect 3990 381 3996 382
rect 110 380 116 381
rect 110 376 111 380
rect 115 376 116 380
rect 110 375 116 376
rect 2030 380 2036 381
rect 2030 376 2031 380
rect 2035 376 2036 380
rect 2070 377 2071 381
rect 2075 377 2076 381
rect 2070 376 2076 377
rect 3990 377 3991 381
rect 3995 377 3996 381
rect 3990 376 3996 377
rect 2030 375 2036 376
rect 614 371 620 372
rect 614 370 615 371
rect 545 368 615 370
rect 614 367 615 368
rect 619 367 620 371
rect 750 371 756 372
rect 750 370 751 371
rect 681 368 751 370
rect 614 366 620 367
rect 750 367 751 368
rect 755 367 756 371
rect 838 371 844 372
rect 838 370 839 371
rect 817 368 839 370
rect 750 366 756 367
rect 838 367 839 368
rect 843 367 844 371
rect 1030 371 1036 372
rect 1030 370 1031 371
rect 961 368 1031 370
rect 838 366 844 367
rect 1030 367 1031 368
rect 1035 367 1036 371
rect 1030 366 1036 367
rect 1038 371 1044 372
rect 1038 367 1039 371
rect 1043 367 1044 371
rect 1302 371 1308 372
rect 1302 370 1303 371
rect 1233 368 1303 370
rect 1038 366 1044 367
rect 1302 367 1303 368
rect 1307 367 1308 371
rect 1558 371 1564 372
rect 1558 370 1559 371
rect 1497 368 1559 370
rect 1302 366 1308 367
rect 1558 367 1559 368
rect 1563 367 1564 371
rect 1686 371 1692 372
rect 1686 370 1687 371
rect 1625 368 1687 370
rect 1558 366 1564 367
rect 1686 367 1687 368
rect 1691 367 1692 371
rect 1774 371 1780 372
rect 1774 370 1775 371
rect 1753 368 1775 370
rect 1686 366 1692 367
rect 1774 367 1775 368
rect 1779 367 1780 371
rect 1774 366 1780 367
rect 1846 371 1852 372
rect 1846 367 1847 371
rect 1851 367 1852 371
rect 1846 366 1852 367
rect 2070 364 2076 365
rect 494 361 500 362
rect 494 357 495 361
rect 499 357 500 361
rect 494 356 500 357
rect 630 361 636 362
rect 630 357 631 361
rect 635 357 636 361
rect 630 356 636 357
rect 766 361 772 362
rect 766 357 767 361
rect 771 357 772 361
rect 766 356 772 357
rect 910 361 916 362
rect 910 357 911 361
rect 915 357 916 361
rect 910 356 916 357
rect 1046 361 1052 362
rect 1046 357 1047 361
rect 1051 357 1052 361
rect 1046 356 1052 357
rect 1182 361 1188 362
rect 1182 357 1183 361
rect 1187 357 1188 361
rect 1182 356 1188 357
rect 1318 361 1324 362
rect 1318 357 1319 361
rect 1323 357 1324 361
rect 1318 356 1324 357
rect 1446 361 1452 362
rect 1446 357 1447 361
rect 1451 357 1452 361
rect 1446 356 1452 357
rect 1574 361 1580 362
rect 1574 357 1575 361
rect 1579 357 1580 361
rect 1574 356 1580 357
rect 1702 361 1708 362
rect 1702 357 1703 361
rect 1707 357 1708 361
rect 1702 356 1708 357
rect 1830 361 1836 362
rect 1830 357 1831 361
rect 1835 357 1836 361
rect 1830 356 1836 357
rect 1934 361 1940 362
rect 1934 357 1935 361
rect 1939 357 1940 361
rect 2070 360 2071 364
rect 2075 360 2076 364
rect 2070 359 2076 360
rect 3990 364 3996 365
rect 3990 360 3991 364
rect 3995 360 3996 364
rect 3990 359 3996 360
rect 1934 356 1940 357
rect 3103 355 3109 356
rect 3103 354 3104 355
rect 3009 352 3104 354
rect 558 351 564 352
rect 558 347 559 351
rect 563 350 564 351
rect 567 351 573 352
rect 567 350 568 351
rect 563 348 568 350
rect 563 347 564 348
rect 558 346 564 347
rect 567 347 568 348
rect 572 347 573 351
rect 567 346 573 347
rect 614 351 620 352
rect 614 347 615 351
rect 619 350 620 351
rect 703 351 709 352
rect 703 350 704 351
rect 619 348 704 350
rect 619 347 620 348
rect 614 346 620 347
rect 703 347 704 348
rect 708 347 709 351
rect 703 346 709 347
rect 750 351 756 352
rect 750 347 751 351
rect 755 350 756 351
rect 839 351 845 352
rect 839 350 840 351
rect 755 348 840 350
rect 755 347 756 348
rect 750 346 756 347
rect 839 347 840 348
rect 844 347 845 351
rect 839 346 845 347
rect 966 351 972 352
rect 966 347 967 351
rect 971 350 972 351
rect 983 351 989 352
rect 983 350 984 351
rect 971 348 984 350
rect 971 347 972 348
rect 966 346 972 347
rect 983 347 984 348
rect 988 347 989 351
rect 983 346 989 347
rect 1030 351 1036 352
rect 1030 347 1031 351
rect 1035 350 1036 351
rect 1119 351 1125 352
rect 1119 350 1120 351
rect 1035 348 1120 350
rect 1035 347 1036 348
rect 1030 346 1036 347
rect 1119 347 1120 348
rect 1124 347 1125 351
rect 1119 346 1125 347
rect 1255 351 1261 352
rect 1255 347 1256 351
rect 1260 350 1261 351
rect 1303 351 1309 352
rect 1303 350 1304 351
rect 1260 348 1304 350
rect 1260 347 1261 348
rect 1255 346 1261 347
rect 1303 347 1304 348
rect 1308 347 1309 351
rect 1303 346 1309 347
rect 1391 351 1397 352
rect 1391 347 1392 351
rect 1396 350 1397 351
rect 1406 351 1412 352
rect 1406 350 1407 351
rect 1396 348 1407 350
rect 1396 347 1397 348
rect 1391 346 1397 347
rect 1406 347 1407 348
rect 1411 347 1412 351
rect 1519 351 1525 352
rect 1519 350 1520 351
rect 1406 346 1412 347
rect 1416 348 1520 350
rect 1302 343 1308 344
rect 1302 339 1303 343
rect 1307 342 1308 343
rect 1416 342 1418 348
rect 1519 347 1520 348
rect 1524 347 1525 351
rect 1519 346 1525 347
rect 1558 351 1564 352
rect 1558 347 1559 351
rect 1563 350 1564 351
rect 1647 351 1653 352
rect 1647 350 1648 351
rect 1563 348 1648 350
rect 1563 347 1564 348
rect 1558 346 1564 347
rect 1647 347 1648 348
rect 1652 347 1653 351
rect 1647 346 1653 347
rect 1686 351 1692 352
rect 1686 347 1687 351
rect 1691 350 1692 351
rect 1775 351 1781 352
rect 1775 350 1776 351
rect 1691 348 1776 350
rect 1691 347 1692 348
rect 1686 346 1692 347
rect 1775 347 1776 348
rect 1780 347 1781 351
rect 1775 346 1781 347
rect 1903 351 1909 352
rect 1903 347 1904 351
rect 1908 350 1909 351
rect 1919 351 1925 352
rect 1919 350 1920 351
rect 1908 348 1920 350
rect 1908 347 1909 348
rect 1903 346 1909 347
rect 1919 347 1920 348
rect 1924 347 1925 351
rect 1919 346 1925 347
rect 2007 351 2013 352
rect 2007 347 2008 351
rect 2012 350 2013 351
rect 2094 351 2100 352
rect 2094 350 2095 351
rect 2012 348 2095 350
rect 2012 347 2013 348
rect 2007 346 2013 347
rect 2094 347 2095 348
rect 2099 347 2100 351
rect 3103 351 3104 352
rect 3108 351 3109 355
rect 3838 355 3844 356
rect 3838 354 3839 355
rect 3761 352 3839 354
rect 3103 350 3109 351
rect 3838 351 3839 352
rect 3843 351 3844 355
rect 3966 355 3972 356
rect 3966 354 3967 355
rect 3945 352 3967 354
rect 3838 350 3844 351
rect 3966 351 3967 352
rect 3971 351 3972 355
rect 3966 350 3972 351
rect 2094 346 2100 347
rect 1307 340 1418 342
rect 2590 345 2596 346
rect 2590 341 2591 345
rect 2595 341 2596 345
rect 2590 340 2596 341
rect 2694 345 2700 346
rect 2694 341 2695 345
rect 2699 341 2700 345
rect 2694 340 2700 341
rect 2814 345 2820 346
rect 2814 341 2815 345
rect 2819 341 2820 345
rect 2814 340 2820 341
rect 2958 345 2964 346
rect 2958 341 2959 345
rect 2963 341 2964 345
rect 2958 340 2964 341
rect 3118 345 3124 346
rect 3118 341 3119 345
rect 3123 341 3124 345
rect 3118 340 3124 341
rect 3302 345 3308 346
rect 3302 341 3303 345
rect 3307 341 3308 345
rect 3302 340 3308 341
rect 3502 345 3508 346
rect 3502 341 3503 345
rect 3507 341 3508 345
rect 3502 340 3508 341
rect 3710 345 3716 346
rect 3710 341 3711 345
rect 3715 341 3716 345
rect 3710 340 3716 341
rect 3894 345 3900 346
rect 3894 341 3895 345
rect 3899 341 3900 345
rect 3894 340 3900 341
rect 1307 339 1308 340
rect 1302 338 1308 339
rect 446 335 452 336
rect 446 331 447 335
rect 451 334 452 335
rect 854 335 860 336
rect 854 334 855 335
rect 451 332 855 334
rect 451 331 452 332
rect 446 330 452 331
rect 854 331 855 332
rect 859 331 860 335
rect 854 330 860 331
rect 1686 335 1692 336
rect 1686 331 1687 335
rect 1691 334 1692 335
rect 2575 335 2581 336
rect 2575 334 2576 335
rect 1691 332 1786 334
rect 1691 331 1692 332
rect 1686 330 1692 331
rect 407 327 413 328
rect 407 323 408 327
rect 412 326 413 327
rect 447 327 453 328
rect 447 326 448 327
rect 412 324 448 326
rect 412 323 413 324
rect 407 322 413 323
rect 447 323 448 324
rect 452 323 453 327
rect 447 322 453 323
rect 535 327 541 328
rect 535 323 536 327
rect 540 326 541 327
rect 591 327 597 328
rect 591 326 592 327
rect 540 324 592 326
rect 540 323 541 324
rect 535 322 541 323
rect 591 323 592 324
rect 596 323 597 327
rect 591 322 597 323
rect 679 327 685 328
rect 679 323 680 327
rect 684 326 685 327
rect 751 327 757 328
rect 751 326 752 327
rect 684 324 752 326
rect 684 323 685 324
rect 679 322 685 323
rect 751 323 752 324
rect 756 323 757 327
rect 751 322 757 323
rect 838 327 845 328
rect 838 323 839 327
rect 844 323 845 327
rect 838 322 845 323
rect 1015 327 1021 328
rect 1015 323 1016 327
rect 1020 326 1021 327
rect 1111 327 1117 328
rect 1111 326 1112 327
rect 1020 324 1112 326
rect 1020 323 1021 324
rect 1015 322 1021 323
rect 1111 323 1112 324
rect 1116 323 1117 327
rect 1111 322 1117 323
rect 1199 327 1205 328
rect 1199 323 1200 327
rect 1204 326 1205 327
rect 1295 327 1301 328
rect 1295 326 1296 327
rect 1204 324 1296 326
rect 1204 323 1205 324
rect 1199 322 1205 323
rect 1295 323 1296 324
rect 1300 323 1301 327
rect 1295 322 1301 323
rect 1382 327 1389 328
rect 1382 323 1383 327
rect 1388 323 1389 327
rect 1382 322 1389 323
rect 1575 327 1581 328
rect 1575 323 1576 327
rect 1580 326 1581 327
rect 1687 327 1693 328
rect 1687 326 1688 327
rect 1580 324 1688 326
rect 1580 323 1581 324
rect 1575 322 1581 323
rect 1687 323 1688 324
rect 1692 323 1693 327
rect 1687 322 1693 323
rect 1774 327 1781 328
rect 1774 323 1775 327
rect 1780 323 1781 327
rect 1784 326 1786 332
rect 2556 332 2576 334
rect 1975 327 1981 328
rect 1975 326 1976 327
rect 1784 324 1976 326
rect 1774 322 1781 323
rect 1975 323 1976 324
rect 1980 323 1981 327
rect 1975 322 1981 323
rect 2094 323 2101 324
rect 334 319 340 320
rect 334 315 335 319
rect 339 315 340 319
rect 334 314 340 315
rect 462 319 468 320
rect 462 315 463 319
rect 467 315 468 319
rect 462 314 468 315
rect 606 319 612 320
rect 606 315 607 319
rect 611 315 612 319
rect 606 314 612 315
rect 766 319 772 320
rect 766 315 767 319
rect 771 315 772 319
rect 766 314 772 315
rect 942 319 948 320
rect 942 315 943 319
rect 947 315 948 319
rect 942 314 948 315
rect 1126 319 1132 320
rect 1126 315 1127 319
rect 1131 315 1132 319
rect 1126 314 1132 315
rect 1310 319 1316 320
rect 1310 315 1311 319
rect 1315 315 1316 319
rect 1310 314 1316 315
rect 1502 319 1508 320
rect 1502 315 1503 319
rect 1507 315 1508 319
rect 1502 314 1508 315
rect 1702 319 1708 320
rect 1702 315 1703 319
rect 1707 315 1708 319
rect 1702 314 1708 315
rect 1902 319 1908 320
rect 1902 315 1903 319
rect 1907 315 1908 319
rect 2094 319 2095 323
rect 2100 319 2101 323
rect 2094 318 2101 319
rect 2183 323 2189 324
rect 2183 319 2184 323
rect 2188 322 2189 323
rect 2255 323 2261 324
rect 2255 322 2256 323
rect 2188 320 2256 322
rect 2188 319 2189 320
rect 2183 318 2189 319
rect 2255 319 2256 320
rect 2260 319 2261 323
rect 2255 318 2261 319
rect 2343 323 2349 324
rect 2343 319 2344 323
rect 2348 322 2349 323
rect 2462 323 2468 324
rect 2462 322 2463 323
rect 2348 320 2463 322
rect 2348 319 2349 320
rect 2343 318 2349 319
rect 2462 319 2463 320
rect 2467 319 2468 323
rect 2462 318 2468 319
rect 2527 323 2533 324
rect 2527 319 2528 323
rect 2532 322 2533 323
rect 2556 322 2558 332
rect 2575 331 2576 332
rect 2580 331 2581 335
rect 2575 330 2581 331
rect 2663 335 2669 336
rect 2663 331 2664 335
rect 2668 334 2669 335
rect 2679 335 2685 336
rect 2679 334 2680 335
rect 2668 332 2680 334
rect 2668 331 2669 332
rect 2663 330 2669 331
rect 2679 331 2680 332
rect 2684 331 2685 335
rect 2679 330 2685 331
rect 2767 335 2773 336
rect 2767 331 2768 335
rect 2772 334 2773 335
rect 2799 335 2805 336
rect 2799 334 2800 335
rect 2772 332 2800 334
rect 2772 331 2773 332
rect 2767 330 2773 331
rect 2799 331 2800 332
rect 2804 331 2805 335
rect 2799 330 2805 331
rect 2886 335 2893 336
rect 2886 331 2887 335
rect 2892 331 2893 335
rect 2886 330 2893 331
rect 3031 335 3037 336
rect 3031 331 3032 335
rect 3036 334 3037 335
rect 3103 335 3109 336
rect 3103 334 3104 335
rect 3036 332 3104 334
rect 3036 331 3037 332
rect 3031 330 3037 331
rect 3103 331 3104 332
rect 3108 331 3109 335
rect 3103 330 3109 331
rect 3191 335 3197 336
rect 3191 331 3192 335
rect 3196 334 3197 335
rect 3287 335 3293 336
rect 3287 334 3288 335
rect 3196 332 3288 334
rect 3196 331 3197 332
rect 3191 330 3197 331
rect 3287 331 3288 332
rect 3292 331 3293 335
rect 3287 330 3293 331
rect 3375 335 3381 336
rect 3375 331 3376 335
rect 3380 334 3381 335
rect 3487 335 3493 336
rect 3487 334 3488 335
rect 3380 332 3488 334
rect 3380 331 3381 332
rect 3375 330 3381 331
rect 3487 331 3488 332
rect 3492 331 3493 335
rect 3487 330 3493 331
rect 3510 335 3516 336
rect 3510 331 3511 335
rect 3515 334 3516 335
rect 3575 335 3581 336
rect 3575 334 3576 335
rect 3515 332 3576 334
rect 3515 331 3516 332
rect 3510 330 3516 331
rect 3575 331 3576 332
rect 3580 331 3581 335
rect 3575 330 3581 331
rect 3782 335 3789 336
rect 3782 331 3783 335
rect 3788 331 3789 335
rect 3782 330 3789 331
rect 3958 335 3964 336
rect 3958 331 3959 335
rect 3963 334 3964 335
rect 3967 335 3973 336
rect 3967 334 3968 335
rect 3963 332 3968 334
rect 3963 331 3964 332
rect 3958 330 3964 331
rect 3967 331 3968 332
rect 3972 331 3973 335
rect 3967 330 3973 331
rect 2703 323 2709 324
rect 2703 322 2704 323
rect 2532 320 2558 322
rect 2576 320 2704 322
rect 2532 319 2533 320
rect 2527 318 2533 319
rect 1902 314 1908 315
rect 2110 315 2116 316
rect 446 311 452 312
rect 446 310 447 311
rect 385 308 447 310
rect 446 307 447 308
rect 451 307 452 311
rect 1686 311 1692 312
rect 1686 310 1687 311
rect 1553 308 1687 310
rect 446 306 452 307
rect 966 307 972 308
rect 966 303 967 307
rect 971 303 972 307
rect 1686 307 1687 308
rect 1691 307 1692 311
rect 2110 311 2111 315
rect 2115 311 2116 315
rect 2110 310 2116 311
rect 2270 315 2276 316
rect 2270 311 2271 315
rect 2275 311 2276 315
rect 2270 310 2276 311
rect 2454 315 2460 316
rect 2454 311 2455 315
rect 2459 311 2460 315
rect 2454 310 2460 311
rect 1686 306 1692 307
rect 1894 307 1900 308
rect 966 302 972 303
rect 1894 303 1895 307
rect 1899 303 1900 307
rect 2576 306 2578 320
rect 2703 319 2704 320
rect 2708 319 2709 323
rect 2703 318 2709 319
rect 2879 323 2885 324
rect 2879 319 2880 323
rect 2884 322 2885 323
rect 2983 323 2989 324
rect 2983 322 2984 323
rect 2884 320 2984 322
rect 2884 319 2885 320
rect 2879 318 2885 319
rect 2983 319 2984 320
rect 2988 319 2989 323
rect 2983 318 2989 319
rect 3071 323 3077 324
rect 3071 319 3072 323
rect 3076 322 3077 323
rect 3199 323 3205 324
rect 3199 322 3200 323
rect 3076 320 3200 322
rect 3076 319 3077 320
rect 3071 318 3077 319
rect 3199 319 3200 320
rect 3204 319 3205 323
rect 3199 318 3205 319
rect 3287 323 3293 324
rect 3287 319 3288 323
rect 3292 322 3293 323
rect 3423 323 3429 324
rect 3423 322 3424 323
rect 3292 320 3424 322
rect 3292 319 3293 320
rect 3287 318 3293 319
rect 3423 319 3424 320
rect 3428 319 3429 323
rect 3423 318 3429 319
rect 3511 323 3517 324
rect 3511 319 3512 323
rect 3516 322 3517 323
rect 3663 323 3669 324
rect 3663 322 3664 323
rect 3516 320 3664 322
rect 3516 319 3517 320
rect 3511 318 3517 319
rect 3663 319 3664 320
rect 3668 319 3669 323
rect 3663 318 3669 319
rect 3686 323 3692 324
rect 3686 319 3687 323
rect 3691 322 3692 323
rect 3751 323 3757 324
rect 3751 322 3752 323
rect 3691 320 3752 322
rect 3691 319 3692 320
rect 3686 318 3692 319
rect 3751 319 3752 320
rect 3756 319 3757 323
rect 3751 318 3757 319
rect 3966 323 3973 324
rect 3966 319 3967 323
rect 3972 319 3973 323
rect 3966 318 3973 319
rect 2630 315 2636 316
rect 2630 311 2631 315
rect 2635 311 2636 315
rect 2630 310 2636 311
rect 2806 315 2812 316
rect 2806 311 2807 315
rect 2811 311 2812 315
rect 2806 310 2812 311
rect 2998 315 3004 316
rect 2998 311 2999 315
rect 3003 311 3004 315
rect 2998 310 3004 311
rect 3214 315 3220 316
rect 3214 311 3215 315
rect 3219 311 3220 315
rect 3214 310 3220 311
rect 3438 315 3444 316
rect 3438 311 3439 315
rect 3443 311 3444 315
rect 3438 310 3444 311
rect 3678 315 3684 316
rect 3678 311 3679 315
rect 3683 311 3684 315
rect 3678 310 3684 311
rect 3894 315 3900 316
rect 3894 311 3895 315
rect 3899 311 3900 315
rect 3894 310 3900 311
rect 2758 307 2764 308
rect 2758 306 2759 307
rect 2505 304 2578 306
rect 2681 304 2759 306
rect 1894 302 1900 303
rect 2758 303 2759 304
rect 2763 303 2764 307
rect 2982 307 2988 308
rect 2982 306 2983 307
rect 2857 304 2983 306
rect 2758 302 2764 303
rect 2982 303 2983 304
rect 2987 303 2988 307
rect 3958 307 3964 308
rect 3958 306 3959 307
rect 3945 304 3959 306
rect 2982 302 2988 303
rect 3958 303 3959 304
rect 3963 303 3964 307
rect 3958 302 3964 303
rect 110 300 116 301
rect 110 296 111 300
rect 115 296 116 300
rect 110 295 116 296
rect 2030 300 2036 301
rect 2030 296 2031 300
rect 2035 296 2036 300
rect 2030 295 2036 296
rect 2070 296 2076 297
rect 2070 292 2071 296
rect 2075 292 2076 296
rect 2070 291 2076 292
rect 3990 296 3996 297
rect 3990 292 3991 296
rect 3995 292 3996 296
rect 3990 291 3996 292
rect 110 283 116 284
rect 110 279 111 283
rect 115 279 116 283
rect 2030 283 2036 284
rect 2030 279 2031 283
rect 2035 279 2036 283
rect 110 278 116 279
rect 334 278 340 279
rect 334 274 335 278
rect 339 274 340 278
rect 334 273 340 274
rect 462 278 468 279
rect 462 274 463 278
rect 467 274 468 278
rect 462 273 468 274
rect 606 278 612 279
rect 606 274 607 278
rect 611 274 612 278
rect 606 273 612 274
rect 766 278 772 279
rect 766 274 767 278
rect 771 274 772 278
rect 766 273 772 274
rect 942 278 948 279
rect 942 274 943 278
rect 947 274 948 278
rect 942 273 948 274
rect 1126 278 1132 279
rect 1126 274 1127 278
rect 1131 274 1132 278
rect 1126 273 1132 274
rect 1310 278 1316 279
rect 1310 274 1311 278
rect 1315 274 1316 278
rect 1310 273 1316 274
rect 1502 278 1508 279
rect 1502 274 1503 278
rect 1507 274 1508 278
rect 1502 273 1508 274
rect 1702 278 1708 279
rect 1702 274 1703 278
rect 1707 274 1708 278
rect 1702 273 1708 274
rect 1902 278 1908 279
rect 2030 278 2036 279
rect 2070 279 2076 280
rect 1902 274 1903 278
rect 1907 274 1908 278
rect 2070 275 2071 279
rect 2075 275 2076 279
rect 3990 279 3996 280
rect 3990 275 3991 279
rect 3995 275 3996 279
rect 2070 274 2076 275
rect 2110 274 2116 275
rect 1902 273 1908 274
rect 2110 270 2111 274
rect 2115 270 2116 274
rect 2110 269 2116 270
rect 2270 274 2276 275
rect 2270 270 2271 274
rect 2275 270 2276 274
rect 2270 269 2276 270
rect 2454 274 2460 275
rect 2454 270 2455 274
rect 2459 270 2460 274
rect 2454 269 2460 270
rect 2630 274 2636 275
rect 2630 270 2631 274
rect 2635 270 2636 274
rect 2630 269 2636 270
rect 2806 274 2812 275
rect 2806 270 2807 274
rect 2811 270 2812 274
rect 2806 269 2812 270
rect 2998 274 3004 275
rect 2998 270 2999 274
rect 3003 270 3004 274
rect 2998 269 3004 270
rect 3214 274 3220 275
rect 3214 270 3215 274
rect 3219 270 3220 274
rect 3214 269 3220 270
rect 3438 274 3444 275
rect 3438 270 3439 274
rect 3443 270 3444 274
rect 3438 269 3444 270
rect 3678 274 3684 275
rect 3678 270 3679 274
rect 3683 270 3684 274
rect 3678 269 3684 270
rect 3894 274 3900 275
rect 3990 274 3996 275
rect 3894 270 3895 274
rect 3899 270 3900 274
rect 3894 269 3900 270
rect 2110 242 2116 243
rect 150 238 156 239
rect 150 234 151 238
rect 155 234 156 238
rect 110 233 116 234
rect 150 233 156 234
rect 278 238 284 239
rect 278 234 279 238
rect 283 234 284 238
rect 278 233 284 234
rect 430 238 436 239
rect 430 234 431 238
rect 435 234 436 238
rect 430 233 436 234
rect 598 238 604 239
rect 598 234 599 238
rect 603 234 604 238
rect 598 233 604 234
rect 782 238 788 239
rect 782 234 783 238
rect 787 234 788 238
rect 782 233 788 234
rect 974 238 980 239
rect 974 234 975 238
rect 979 234 980 238
rect 974 233 980 234
rect 1174 238 1180 239
rect 1174 234 1175 238
rect 1179 234 1180 238
rect 1174 233 1180 234
rect 1374 238 1380 239
rect 1374 234 1375 238
rect 1379 234 1380 238
rect 1374 233 1380 234
rect 1582 238 1588 239
rect 1582 234 1583 238
rect 1587 234 1588 238
rect 1582 233 1588 234
rect 1798 238 1804 239
rect 2110 238 2111 242
rect 2115 238 2116 242
rect 1798 234 1799 238
rect 1803 234 1804 238
rect 2070 237 2076 238
rect 2110 237 2116 238
rect 2270 242 2276 243
rect 2270 238 2271 242
rect 2275 238 2276 242
rect 2270 237 2276 238
rect 2470 242 2476 243
rect 2470 238 2471 242
rect 2475 238 2476 242
rect 2470 237 2476 238
rect 2686 242 2692 243
rect 2686 238 2687 242
rect 2691 238 2692 242
rect 2686 237 2692 238
rect 2902 242 2908 243
rect 2902 238 2903 242
rect 2907 238 2908 242
rect 2902 237 2908 238
rect 3110 242 3116 243
rect 3110 238 3111 242
rect 3115 238 3116 242
rect 3110 237 3116 238
rect 3318 242 3324 243
rect 3318 238 3319 242
rect 3323 238 3324 242
rect 3318 237 3324 238
rect 3518 242 3524 243
rect 3518 238 3519 242
rect 3523 238 3524 242
rect 3518 237 3524 238
rect 3718 242 3724 243
rect 3718 238 3719 242
rect 3723 238 3724 242
rect 3718 237 3724 238
rect 3894 242 3900 243
rect 3894 238 3895 242
rect 3899 238 3900 242
rect 3894 237 3900 238
rect 3990 237 3996 238
rect 1798 233 1804 234
rect 2030 233 2036 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 2030 229 2031 233
rect 2035 229 2036 233
rect 2070 233 2071 237
rect 2075 233 2076 237
rect 2070 232 2076 233
rect 3990 233 3991 237
rect 3995 233 3996 237
rect 3990 232 3996 233
rect 2030 228 2036 229
rect 3302 231 3308 232
rect 3302 227 3303 231
rect 3307 230 3308 231
rect 3686 231 3692 232
rect 3686 230 3687 231
rect 3307 228 3687 230
rect 3307 227 3308 228
rect 3302 226 3308 227
rect 3686 227 3687 228
rect 3691 227 3692 231
rect 3686 226 3692 227
rect 2070 220 2076 221
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 110 211 116 212
rect 2030 216 2036 217
rect 2030 212 2031 216
rect 2035 212 2036 216
rect 2070 216 2071 220
rect 2075 216 2076 220
rect 2070 215 2076 216
rect 3990 220 3996 221
rect 3990 216 3991 220
rect 3995 216 3996 220
rect 3990 215 3996 216
rect 2030 211 2036 212
rect 2254 211 2260 212
rect 2254 210 2255 211
rect 2161 208 2255 210
rect 230 207 236 208
rect 230 206 231 207
rect 201 204 231 206
rect 230 203 231 204
rect 235 203 236 207
rect 1158 207 1164 208
rect 1158 206 1159 207
rect 1025 204 1159 206
rect 230 202 236 203
rect 1158 203 1159 204
rect 1163 203 1164 207
rect 1358 207 1364 208
rect 1358 206 1359 207
rect 1225 204 1359 206
rect 1158 202 1164 203
rect 1358 203 1359 204
rect 1363 203 1364 207
rect 1358 202 1364 203
rect 1382 207 1388 208
rect 1382 203 1383 207
rect 1387 203 1388 207
rect 1767 207 1773 208
rect 1767 206 1768 207
rect 1633 204 1768 206
rect 1382 202 1388 203
rect 1767 203 1768 204
rect 1772 203 1773 207
rect 2254 207 2255 208
rect 2259 207 2260 211
rect 2454 211 2460 212
rect 2454 210 2455 211
rect 2321 208 2455 210
rect 2254 206 2260 207
rect 2454 207 2455 208
rect 2459 207 2460 211
rect 2454 206 2460 207
rect 2462 211 2468 212
rect 2462 207 2463 211
rect 2467 207 2468 211
rect 2767 211 2773 212
rect 2767 210 2768 211
rect 2737 208 2768 210
rect 2462 206 2468 207
rect 2767 207 2768 208
rect 2772 207 2773 211
rect 3302 211 3308 212
rect 3302 210 3303 211
rect 3161 208 3303 210
rect 2767 206 2773 207
rect 3302 207 3303 208
rect 3307 207 3308 211
rect 3495 211 3501 212
rect 3495 210 3496 211
rect 3369 208 3496 210
rect 3302 206 3308 207
rect 3495 207 3496 208
rect 3500 207 3501 211
rect 3966 211 3972 212
rect 3966 210 3967 211
rect 3945 208 3967 210
rect 3495 206 3501 207
rect 3966 207 3967 208
rect 3971 207 3972 211
rect 3966 206 3972 207
rect 1767 202 1773 203
rect 2110 201 2116 202
rect 150 197 156 198
rect 150 193 151 197
rect 155 193 156 197
rect 150 192 156 193
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 430 197 436 198
rect 430 193 431 197
rect 435 193 436 197
rect 430 192 436 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 782 197 788 198
rect 782 193 783 197
rect 787 193 788 197
rect 782 192 788 193
rect 974 197 980 198
rect 974 193 975 197
rect 979 193 980 197
rect 974 192 980 193
rect 1174 197 1180 198
rect 1174 193 1175 197
rect 1179 193 1180 197
rect 1174 192 1180 193
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1582 197 1588 198
rect 1582 193 1583 197
rect 1587 193 1588 197
rect 1582 192 1588 193
rect 1798 197 1804 198
rect 1798 193 1799 197
rect 1803 193 1804 197
rect 2110 197 2111 201
rect 2115 197 2116 201
rect 2110 196 2116 197
rect 2270 201 2276 202
rect 2270 197 2271 201
rect 2275 197 2276 201
rect 2270 196 2276 197
rect 2470 201 2476 202
rect 2470 197 2471 201
rect 2475 197 2476 201
rect 2470 196 2476 197
rect 2686 201 2692 202
rect 2686 197 2687 201
rect 2691 197 2692 201
rect 2902 201 2908 202
rect 2686 196 2692 197
rect 2855 199 2861 200
rect 2855 195 2856 199
rect 2860 198 2861 199
rect 2887 199 2893 200
rect 2887 198 2888 199
rect 2860 196 2888 198
rect 2860 195 2861 196
rect 2855 194 2861 195
rect 2887 195 2888 196
rect 2892 195 2893 199
rect 2902 197 2903 201
rect 2907 197 2908 201
rect 2902 196 2908 197
rect 3110 201 3116 202
rect 3110 197 3111 201
rect 3115 197 3116 201
rect 3110 196 3116 197
rect 3318 201 3324 202
rect 3318 197 3319 201
rect 3323 197 3324 201
rect 3318 196 3324 197
rect 3518 201 3524 202
rect 3518 197 3519 201
rect 3523 197 3524 201
rect 3518 196 3524 197
rect 3718 201 3724 202
rect 3718 197 3719 201
rect 3723 197 3724 201
rect 3718 196 3724 197
rect 3894 201 3900 202
rect 3894 197 3895 201
rect 3899 197 3900 201
rect 3894 196 3900 197
rect 2887 194 2893 195
rect 1798 192 1804 193
rect 2174 191 2180 192
rect 223 187 229 188
rect 223 183 224 187
rect 228 186 229 187
rect 263 187 269 188
rect 263 186 264 187
rect 228 184 264 186
rect 228 183 229 184
rect 223 182 229 183
rect 263 183 264 184
rect 268 183 269 187
rect 263 182 269 183
rect 351 187 357 188
rect 351 183 352 187
rect 356 186 357 187
rect 415 187 421 188
rect 415 186 416 187
rect 356 184 416 186
rect 356 183 357 184
rect 351 182 357 183
rect 415 183 416 184
rect 420 183 421 187
rect 415 182 421 183
rect 503 187 509 188
rect 503 183 504 187
rect 508 186 509 187
rect 583 187 589 188
rect 583 186 584 187
rect 508 184 584 186
rect 508 183 509 184
rect 503 182 509 183
rect 583 183 584 184
rect 588 183 589 187
rect 583 182 589 183
rect 671 187 677 188
rect 671 183 672 187
rect 676 186 677 187
rect 767 187 773 188
rect 767 186 768 187
rect 676 184 768 186
rect 676 183 677 184
rect 671 182 677 183
rect 767 183 768 184
rect 772 183 773 187
rect 767 182 773 183
rect 854 187 861 188
rect 854 183 855 187
rect 860 183 861 187
rect 854 182 861 183
rect 1038 187 1044 188
rect 1038 183 1039 187
rect 1043 186 1044 187
rect 1047 187 1053 188
rect 1047 186 1048 187
rect 1043 184 1048 186
rect 1043 183 1044 184
rect 1038 182 1044 183
rect 1047 183 1048 184
rect 1052 183 1053 187
rect 1047 182 1053 183
rect 1158 187 1164 188
rect 1158 183 1159 187
rect 1163 186 1164 187
rect 1247 187 1253 188
rect 1247 186 1248 187
rect 1163 184 1248 186
rect 1163 183 1164 184
rect 1158 182 1164 183
rect 1247 183 1248 184
rect 1252 183 1253 187
rect 1247 182 1253 183
rect 1358 187 1364 188
rect 1358 183 1359 187
rect 1363 186 1364 187
rect 1447 187 1453 188
rect 1447 186 1448 187
rect 1363 184 1448 186
rect 1363 183 1364 184
rect 1358 182 1364 183
rect 1447 183 1448 184
rect 1452 183 1453 187
rect 1447 182 1453 183
rect 1655 187 1661 188
rect 1655 183 1656 187
rect 1660 186 1661 187
rect 1783 187 1789 188
rect 1783 186 1784 187
rect 1660 184 1784 186
rect 1660 183 1661 184
rect 1655 182 1661 183
rect 1783 183 1784 184
rect 1788 183 1789 187
rect 1783 182 1789 183
rect 1871 187 1877 188
rect 1871 183 1872 187
rect 1876 186 1877 187
rect 1894 187 1900 188
rect 1894 186 1895 187
rect 1876 184 1895 186
rect 1876 183 1877 184
rect 1871 182 1877 183
rect 1894 183 1895 184
rect 1899 183 1900 187
rect 2174 187 2175 191
rect 2179 190 2180 191
rect 2183 191 2189 192
rect 2183 190 2184 191
rect 2179 188 2184 190
rect 2179 187 2180 188
rect 2174 186 2180 187
rect 2183 187 2184 188
rect 2188 187 2189 191
rect 2183 186 2189 187
rect 2254 191 2260 192
rect 2254 187 2255 191
rect 2259 190 2260 191
rect 2343 191 2349 192
rect 2343 190 2344 191
rect 2259 188 2344 190
rect 2259 187 2260 188
rect 2254 186 2260 187
rect 2343 187 2344 188
rect 2348 187 2349 191
rect 2343 186 2349 187
rect 2454 191 2460 192
rect 2454 187 2455 191
rect 2459 190 2460 191
rect 2543 191 2549 192
rect 2543 190 2544 191
rect 2459 188 2544 190
rect 2459 187 2460 188
rect 2454 186 2460 187
rect 2543 187 2544 188
rect 2548 187 2549 191
rect 2543 186 2549 187
rect 2758 191 2765 192
rect 2758 187 2759 191
rect 2764 187 2765 191
rect 2758 186 2765 187
rect 2767 191 2773 192
rect 2767 187 2768 191
rect 2772 190 2773 191
rect 2975 191 2981 192
rect 2975 190 2976 191
rect 2772 188 2976 190
rect 2772 187 2773 188
rect 2767 186 2773 187
rect 2975 187 2976 188
rect 2980 187 2981 191
rect 2975 186 2981 187
rect 2998 191 3004 192
rect 2998 187 2999 191
rect 3003 190 3004 191
rect 3183 191 3189 192
rect 3183 190 3184 191
rect 3003 188 3184 190
rect 3003 187 3004 188
rect 2998 186 3004 187
rect 3183 187 3184 188
rect 3188 187 3189 191
rect 3183 186 3189 187
rect 3391 191 3397 192
rect 3391 187 3392 191
rect 3396 190 3397 191
rect 3503 191 3509 192
rect 3503 190 3504 191
rect 3396 188 3504 190
rect 3396 187 3397 188
rect 3391 186 3397 187
rect 3503 187 3504 188
rect 3508 187 3509 191
rect 3503 186 3509 187
rect 3591 191 3597 192
rect 3591 187 3592 191
rect 3596 190 3597 191
rect 3703 191 3709 192
rect 3703 190 3704 191
rect 3596 188 3704 190
rect 3596 187 3597 188
rect 3591 186 3597 187
rect 3703 187 3704 188
rect 3708 187 3709 191
rect 3703 186 3709 187
rect 3782 191 3788 192
rect 3782 187 3783 191
rect 3787 190 3788 191
rect 3791 191 3797 192
rect 3791 190 3792 191
rect 3787 188 3792 190
rect 3787 187 3788 188
rect 3782 186 3788 187
rect 3791 187 3792 188
rect 3796 187 3797 191
rect 3791 186 3797 187
rect 3958 191 3964 192
rect 3958 187 3959 191
rect 3963 190 3964 191
rect 3967 191 3973 192
rect 3967 190 3968 191
rect 3963 188 3968 190
rect 3963 187 3964 188
rect 3958 186 3964 187
rect 3967 187 3968 188
rect 3972 187 3973 191
rect 3967 186 3973 187
rect 1894 182 1900 183
rect 230 159 236 160
rect 230 155 231 159
rect 235 158 236 159
rect 3495 159 3501 160
rect 235 156 874 158
rect 235 155 236 156
rect 230 154 236 155
rect 223 151 229 152
rect 223 147 224 151
rect 228 150 229 151
rect 239 151 245 152
rect 239 150 240 151
rect 228 148 240 150
rect 228 147 229 148
rect 223 146 229 147
rect 239 147 240 148
rect 244 147 245 151
rect 239 146 245 147
rect 327 151 333 152
rect 327 147 328 151
rect 332 150 333 151
rect 343 151 349 152
rect 343 150 344 151
rect 332 148 344 150
rect 332 147 333 148
rect 327 146 333 147
rect 343 147 344 148
rect 348 147 349 151
rect 343 146 349 147
rect 431 151 437 152
rect 431 147 432 151
rect 436 150 437 151
rect 455 151 461 152
rect 455 150 456 151
rect 436 148 456 150
rect 436 147 437 148
rect 431 146 437 147
rect 455 147 456 148
rect 460 147 461 151
rect 455 146 461 147
rect 543 151 549 152
rect 543 147 544 151
rect 548 150 549 151
rect 591 151 597 152
rect 591 150 592 151
rect 548 148 592 150
rect 548 147 549 148
rect 543 146 549 147
rect 591 147 592 148
rect 596 147 597 151
rect 591 146 597 147
rect 679 151 685 152
rect 679 147 680 151
rect 684 150 685 151
rect 727 151 733 152
rect 727 150 728 151
rect 684 148 728 150
rect 684 147 685 148
rect 679 146 685 147
rect 727 147 728 148
rect 732 147 733 151
rect 727 146 733 147
rect 815 151 821 152
rect 815 147 816 151
rect 820 150 821 151
rect 863 151 869 152
rect 863 150 864 151
rect 820 148 864 150
rect 820 147 821 148
rect 815 146 821 147
rect 863 147 864 148
rect 868 147 869 151
rect 872 150 874 156
rect 3495 155 3496 159
rect 3500 158 3501 159
rect 3500 156 3681 158
rect 3500 155 3501 156
rect 3495 154 3501 155
rect 951 151 957 152
rect 951 150 952 151
rect 872 148 952 150
rect 863 146 869 147
rect 951 147 952 148
rect 956 147 957 151
rect 951 146 957 147
rect 1087 151 1093 152
rect 1087 147 1088 151
rect 1092 150 1093 151
rect 1135 151 1141 152
rect 1135 150 1136 151
rect 1092 148 1136 150
rect 1092 147 1093 148
rect 1087 146 1093 147
rect 1135 147 1136 148
rect 1140 147 1141 151
rect 1135 146 1141 147
rect 1223 151 1229 152
rect 1223 147 1224 151
rect 1228 150 1229 151
rect 1263 151 1269 152
rect 1263 150 1264 151
rect 1228 148 1264 150
rect 1228 147 1229 148
rect 1223 146 1229 147
rect 1263 147 1264 148
rect 1268 147 1269 151
rect 1263 146 1269 147
rect 1351 151 1357 152
rect 1351 147 1352 151
rect 1356 150 1357 151
rect 1383 151 1389 152
rect 1383 150 1384 151
rect 1356 148 1384 150
rect 1356 147 1357 148
rect 1351 146 1357 147
rect 1383 147 1384 148
rect 1388 147 1389 151
rect 1383 146 1389 147
rect 1471 151 1477 152
rect 1471 147 1472 151
rect 1476 150 1477 151
rect 1503 151 1509 152
rect 1503 150 1504 151
rect 1476 148 1504 150
rect 1476 147 1477 148
rect 1471 146 1477 147
rect 1503 147 1504 148
rect 1508 147 1509 151
rect 1503 146 1509 147
rect 1591 151 1597 152
rect 1591 147 1592 151
rect 1596 150 1597 151
rect 1631 151 1637 152
rect 1631 150 1632 151
rect 1596 148 1632 150
rect 1596 147 1597 148
rect 1591 146 1597 147
rect 1631 147 1632 148
rect 1636 147 1637 151
rect 1631 146 1637 147
rect 1719 151 1725 152
rect 1719 147 1720 151
rect 1724 150 1725 151
rect 1759 151 1765 152
rect 1759 150 1760 151
rect 1724 148 1760 150
rect 1724 147 1725 148
rect 1719 146 1725 147
rect 1759 147 1760 148
rect 1764 147 1765 151
rect 1759 146 1765 147
rect 1767 151 1773 152
rect 1767 147 1768 151
rect 1772 150 1773 151
rect 1847 151 1853 152
rect 1847 150 1848 151
rect 1772 148 1848 150
rect 1772 147 1773 148
rect 1767 146 1773 147
rect 1847 147 1848 148
rect 1852 147 1853 151
rect 1847 146 1853 147
rect 2183 151 2189 152
rect 2183 147 2184 151
rect 2188 150 2189 151
rect 2199 151 2205 152
rect 2199 150 2200 151
rect 2188 148 2200 150
rect 2188 147 2189 148
rect 2183 146 2189 147
rect 2199 147 2200 148
rect 2204 147 2205 151
rect 2199 146 2205 147
rect 2287 151 2293 152
rect 2287 147 2288 151
rect 2292 150 2293 151
rect 2303 151 2309 152
rect 2303 150 2304 151
rect 2292 148 2304 150
rect 2292 147 2293 148
rect 2287 146 2293 147
rect 2303 147 2304 148
rect 2308 147 2309 151
rect 2303 146 2309 147
rect 2391 151 2397 152
rect 2391 147 2392 151
rect 2396 150 2397 151
rect 2407 151 2413 152
rect 2407 150 2408 151
rect 2396 148 2408 150
rect 2396 147 2397 148
rect 2391 146 2397 147
rect 2407 147 2408 148
rect 2412 147 2413 151
rect 2407 146 2413 147
rect 2495 151 2501 152
rect 2495 147 2496 151
rect 2500 150 2501 151
rect 2511 151 2517 152
rect 2511 150 2512 151
rect 2500 148 2512 150
rect 2500 147 2501 148
rect 2495 146 2501 147
rect 2511 147 2512 148
rect 2516 147 2517 151
rect 2511 146 2517 147
rect 2599 151 2605 152
rect 2599 147 2600 151
rect 2604 150 2605 151
rect 2639 151 2645 152
rect 2639 150 2640 151
rect 2604 148 2640 150
rect 2604 147 2605 148
rect 2599 146 2605 147
rect 2639 147 2640 148
rect 2644 147 2645 151
rect 2639 146 2645 147
rect 2727 151 2733 152
rect 2727 147 2728 151
rect 2732 150 2733 151
rect 2759 151 2765 152
rect 2759 150 2760 151
rect 2732 148 2760 150
rect 2732 147 2733 148
rect 2727 146 2733 147
rect 2759 147 2760 148
rect 2764 147 2765 151
rect 2759 146 2765 147
rect 2847 151 2853 152
rect 2847 147 2848 151
rect 2852 150 2853 151
rect 2855 151 2861 152
rect 2855 150 2856 151
rect 2852 148 2856 150
rect 2852 147 2853 148
rect 2847 146 2853 147
rect 2855 147 2856 148
rect 2860 147 2861 151
rect 2855 146 2861 147
rect 2967 151 2973 152
rect 2967 147 2968 151
rect 2972 150 2973 151
rect 2999 151 3005 152
rect 2999 150 3000 151
rect 2972 148 3000 150
rect 2972 147 2973 148
rect 2967 146 2973 147
rect 2999 147 3000 148
rect 3004 147 3005 151
rect 2999 146 3005 147
rect 3087 151 3093 152
rect 3087 147 3088 151
rect 3092 150 3093 151
rect 3119 151 3125 152
rect 3119 150 3120 151
rect 3092 148 3120 150
rect 3092 147 3093 148
rect 3087 146 3093 147
rect 3119 147 3120 148
rect 3124 147 3125 151
rect 3119 146 3125 147
rect 3207 151 3213 152
rect 3207 147 3208 151
rect 3212 150 3213 151
rect 3231 151 3237 152
rect 3231 150 3232 151
rect 3212 148 3232 150
rect 3212 147 3213 148
rect 3207 146 3213 147
rect 3231 147 3232 148
rect 3236 147 3237 151
rect 3231 146 3237 147
rect 3319 151 3325 152
rect 3319 147 3320 151
rect 3324 150 3325 151
rect 3343 151 3349 152
rect 3343 150 3344 151
rect 3324 148 3344 150
rect 3324 147 3325 148
rect 3319 146 3325 147
rect 3343 147 3344 148
rect 3348 147 3349 151
rect 3343 146 3349 147
rect 3431 151 3437 152
rect 3431 147 3432 151
rect 3436 150 3437 151
rect 3455 151 3461 152
rect 3455 150 3456 151
rect 3436 148 3456 150
rect 3436 147 3437 148
rect 3431 146 3437 147
rect 3455 147 3456 148
rect 3460 147 3461 151
rect 3455 146 3461 147
rect 3543 151 3549 152
rect 3543 147 3544 151
rect 3548 150 3549 151
rect 3567 151 3573 152
rect 3567 150 3568 151
rect 3548 148 3568 150
rect 3548 147 3549 148
rect 3543 146 3549 147
rect 3567 147 3568 148
rect 3572 147 3573 151
rect 3567 146 3573 147
rect 3655 151 3661 152
rect 3655 147 3656 151
rect 3660 150 3661 151
rect 3671 151 3677 152
rect 3671 150 3672 151
rect 3660 148 3672 150
rect 3660 147 3661 148
rect 3655 146 3661 147
rect 3671 147 3672 148
rect 3676 147 3677 151
rect 3679 150 3681 156
rect 3759 151 3765 152
rect 3759 150 3760 151
rect 3679 148 3760 150
rect 3671 146 3677 147
rect 3759 147 3760 148
rect 3764 147 3765 151
rect 3759 146 3765 147
rect 3863 151 3869 152
rect 3863 147 3864 151
rect 3868 150 3869 151
rect 3879 151 3885 152
rect 3879 150 3880 151
rect 3868 148 3880 150
rect 3868 147 3869 148
rect 3863 146 3869 147
rect 3879 147 3880 148
rect 3884 147 3885 151
rect 3879 146 3885 147
rect 3966 151 3973 152
rect 3966 147 3967 151
rect 3972 147 3973 151
rect 3966 146 3973 147
rect 150 143 156 144
rect 150 139 151 143
rect 155 139 156 143
rect 150 138 156 139
rect 254 143 260 144
rect 254 139 255 143
rect 259 139 260 143
rect 254 138 260 139
rect 358 143 364 144
rect 358 139 359 143
rect 363 139 364 143
rect 358 138 364 139
rect 470 143 476 144
rect 470 139 471 143
rect 475 139 476 143
rect 470 138 476 139
rect 606 143 612 144
rect 606 139 607 143
rect 611 139 612 143
rect 606 138 612 139
rect 742 143 748 144
rect 742 139 743 143
rect 747 139 748 143
rect 742 138 748 139
rect 878 143 884 144
rect 878 139 879 143
rect 883 139 884 143
rect 878 138 884 139
rect 1014 143 1020 144
rect 1014 139 1015 143
rect 1019 139 1020 143
rect 1014 138 1020 139
rect 1150 143 1156 144
rect 1150 139 1151 143
rect 1155 139 1156 143
rect 1150 138 1156 139
rect 1278 143 1284 144
rect 1278 139 1279 143
rect 1283 139 1284 143
rect 1278 138 1284 139
rect 1398 143 1404 144
rect 1398 139 1399 143
rect 1403 139 1404 143
rect 1398 138 1404 139
rect 1518 143 1524 144
rect 1518 139 1519 143
rect 1523 139 1524 143
rect 1518 138 1524 139
rect 1646 143 1652 144
rect 1646 139 1647 143
rect 1651 139 1652 143
rect 1646 138 1652 139
rect 1774 143 1780 144
rect 1774 139 1775 143
rect 1779 139 1780 143
rect 1774 138 1780 139
rect 2110 143 2116 144
rect 2110 139 2111 143
rect 2115 139 2116 143
rect 2110 138 2116 139
rect 2214 143 2220 144
rect 2214 139 2215 143
rect 2219 139 2220 143
rect 2214 138 2220 139
rect 2318 143 2324 144
rect 2318 139 2319 143
rect 2323 139 2324 143
rect 2318 138 2324 139
rect 2422 143 2428 144
rect 2422 139 2423 143
rect 2427 139 2428 143
rect 2422 138 2428 139
rect 2526 143 2532 144
rect 2526 139 2527 143
rect 2531 139 2532 143
rect 2526 138 2532 139
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2774 143 2780 144
rect 2774 139 2775 143
rect 2779 139 2780 143
rect 2774 138 2780 139
rect 2894 143 2900 144
rect 2894 139 2895 143
rect 2899 139 2900 143
rect 2894 138 2900 139
rect 3014 143 3020 144
rect 3014 139 3015 143
rect 3019 139 3020 143
rect 3014 138 3020 139
rect 3134 143 3140 144
rect 3134 139 3135 143
rect 3139 139 3140 143
rect 3134 138 3140 139
rect 3246 143 3252 144
rect 3246 139 3247 143
rect 3251 139 3252 143
rect 3246 138 3252 139
rect 3358 143 3364 144
rect 3358 139 3359 143
rect 3363 139 3364 143
rect 3358 138 3364 139
rect 3470 143 3476 144
rect 3470 139 3471 143
rect 3475 139 3476 143
rect 3470 138 3476 139
rect 3582 143 3588 144
rect 3582 139 3583 143
rect 3587 139 3588 143
rect 3582 138 3588 139
rect 3686 143 3692 144
rect 3686 139 3687 143
rect 3691 139 3692 143
rect 3686 138 3692 139
rect 3790 143 3796 144
rect 3790 139 3791 143
rect 3795 139 3796 143
rect 3790 138 3796 139
rect 3894 143 3900 144
rect 3894 139 3895 143
rect 3899 139 3900 143
rect 3894 138 3900 139
rect 2174 135 2180 136
rect 2174 134 2175 135
rect 2161 132 2175 134
rect 1038 131 1044 132
rect 1038 127 1039 131
rect 1043 127 1044 131
rect 2174 131 2175 132
rect 2179 131 2180 135
rect 2998 135 3004 136
rect 2998 134 2999 135
rect 2945 132 2999 134
rect 2174 130 2180 131
rect 2998 131 2999 132
rect 3003 131 3004 135
rect 2998 130 3004 131
rect 3782 135 3788 136
rect 3782 131 3783 135
rect 3787 131 3788 135
rect 3782 130 3788 131
rect 1038 126 1044 127
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 110 119 116 120
rect 2030 124 2036 125
rect 2030 120 2031 124
rect 2035 120 2036 124
rect 2030 119 2036 120
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 3990 124 3996 125
rect 3990 120 3991 124
rect 3995 120 3996 124
rect 3990 119 3996 120
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 2030 107 2036 108
rect 2030 103 2031 107
rect 2035 103 2036 107
rect 110 102 116 103
rect 150 102 156 103
rect 150 98 151 102
rect 155 98 156 102
rect 150 97 156 98
rect 254 102 260 103
rect 254 98 255 102
rect 259 98 260 102
rect 254 97 260 98
rect 358 102 364 103
rect 358 98 359 102
rect 363 98 364 102
rect 358 97 364 98
rect 470 102 476 103
rect 470 98 471 102
rect 475 98 476 102
rect 470 97 476 98
rect 606 102 612 103
rect 606 98 607 102
rect 611 98 612 102
rect 606 97 612 98
rect 742 102 748 103
rect 742 98 743 102
rect 747 98 748 102
rect 742 97 748 98
rect 878 102 884 103
rect 878 98 879 102
rect 883 98 884 102
rect 878 97 884 98
rect 1014 102 1020 103
rect 1014 98 1015 102
rect 1019 98 1020 102
rect 1014 97 1020 98
rect 1150 102 1156 103
rect 1150 98 1151 102
rect 1155 98 1156 102
rect 1150 97 1156 98
rect 1278 102 1284 103
rect 1278 98 1279 102
rect 1283 98 1284 102
rect 1278 97 1284 98
rect 1398 102 1404 103
rect 1398 98 1399 102
rect 1403 98 1404 102
rect 1398 97 1404 98
rect 1518 102 1524 103
rect 1518 98 1519 102
rect 1523 98 1524 102
rect 1518 97 1524 98
rect 1646 102 1652 103
rect 1646 98 1647 102
rect 1651 98 1652 102
rect 1646 97 1652 98
rect 1774 102 1780 103
rect 2030 102 2036 103
rect 2070 107 2076 108
rect 2070 103 2071 107
rect 2075 103 2076 107
rect 3990 107 3996 108
rect 3990 103 3991 107
rect 3995 103 3996 107
rect 2070 102 2076 103
rect 2110 102 2116 103
rect 1774 98 1775 102
rect 1779 98 1780 102
rect 1774 97 1780 98
rect 2110 98 2111 102
rect 2115 98 2116 102
rect 2110 97 2116 98
rect 2214 102 2220 103
rect 2214 98 2215 102
rect 2219 98 2220 102
rect 2214 97 2220 98
rect 2318 102 2324 103
rect 2318 98 2319 102
rect 2323 98 2324 102
rect 2318 97 2324 98
rect 2422 102 2428 103
rect 2422 98 2423 102
rect 2427 98 2428 102
rect 2422 97 2428 98
rect 2526 102 2532 103
rect 2526 98 2527 102
rect 2531 98 2532 102
rect 2526 97 2532 98
rect 2654 102 2660 103
rect 2654 98 2655 102
rect 2659 98 2660 102
rect 2654 97 2660 98
rect 2774 102 2780 103
rect 2774 98 2775 102
rect 2779 98 2780 102
rect 2774 97 2780 98
rect 2894 102 2900 103
rect 2894 98 2895 102
rect 2899 98 2900 102
rect 2894 97 2900 98
rect 3014 102 3020 103
rect 3014 98 3015 102
rect 3019 98 3020 102
rect 3014 97 3020 98
rect 3134 102 3140 103
rect 3134 98 3135 102
rect 3139 98 3140 102
rect 3134 97 3140 98
rect 3246 102 3252 103
rect 3246 98 3247 102
rect 3251 98 3252 102
rect 3246 97 3252 98
rect 3358 102 3364 103
rect 3358 98 3359 102
rect 3363 98 3364 102
rect 3358 97 3364 98
rect 3470 102 3476 103
rect 3470 98 3471 102
rect 3475 98 3476 102
rect 3470 97 3476 98
rect 3582 102 3588 103
rect 3582 98 3583 102
rect 3587 98 3588 102
rect 3582 97 3588 98
rect 3686 102 3692 103
rect 3686 98 3687 102
rect 3691 98 3692 102
rect 3686 97 3692 98
rect 3790 102 3796 103
rect 3790 98 3791 102
rect 3795 98 3796 102
rect 3790 97 3796 98
rect 3894 102 3900 103
rect 3990 102 3996 103
rect 3894 98 3895 102
rect 3899 98 3900 102
rect 3894 97 3900 98
<< m3c >>
rect 327 4046 331 4050
rect 431 4046 435 4050
rect 535 4046 539 4050
rect 639 4046 643 4050
rect 743 4046 747 4050
rect 847 4046 851 4050
rect 951 4046 955 4050
rect 1055 4046 1059 4050
rect 1159 4046 1163 4050
rect 1263 4046 1267 4050
rect 1367 4046 1371 4050
rect 1471 4046 1475 4050
rect 2263 4046 2267 4050
rect 111 4041 115 4045
rect 2031 4041 2035 4045
rect 2367 4046 2371 4050
rect 2471 4046 2475 4050
rect 2575 4046 2579 4050
rect 2679 4046 2683 4050
rect 2071 4041 2075 4045
rect 3991 4041 3995 4045
rect 111 4024 115 4028
rect 2031 4024 2035 4028
rect 2071 4024 2075 4028
rect 3991 4024 3995 4028
rect 411 4015 415 4019
rect 519 4015 523 4019
rect 623 4015 627 4019
rect 727 4015 731 4019
rect 831 4015 835 4019
rect 935 4015 939 4019
rect 1039 4015 1043 4019
rect 1247 4015 1251 4019
rect 2335 4015 2339 4019
rect 327 4005 331 4009
rect 431 4005 435 4009
rect 535 4005 539 4009
rect 639 4005 643 4009
rect 743 4005 747 4009
rect 847 4005 851 4009
rect 951 4005 955 4009
rect 1055 4005 1059 4009
rect 1159 4005 1163 4009
rect 1263 4005 1267 4009
rect 1367 4005 1371 4009
rect 1471 4005 1475 4009
rect 2263 4005 2267 4009
rect 2367 4005 2371 4009
rect 2471 4005 2475 4009
rect 2599 4015 2603 4019
rect 2575 4005 2579 4009
rect 2679 4005 2683 4009
rect 411 3995 415 3999
rect 519 3995 523 3999
rect 623 3995 627 3999
rect 727 3995 731 3999
rect 831 3995 835 3999
rect 935 3995 939 3999
rect 1039 3995 1043 3999
rect 863 3979 864 3983
rect 864 3979 867 3983
rect 1255 3987 1259 3991
rect 2415 3995 2419 3999
rect 1287 3979 1291 3983
rect 1775 3979 1776 3983
rect 1776 3979 1779 3983
rect 2295 3983 2299 3987
rect 2335 3987 2339 3991
rect 175 3971 179 3975
rect 383 3971 387 3975
rect 591 3971 595 3975
rect 791 3971 795 3975
rect 983 3971 987 3975
rect 1167 3971 1171 3975
rect 1343 3971 1347 3975
rect 1519 3971 1523 3975
rect 1703 3971 1707 3975
rect 2231 3975 2235 3979
rect 2599 3983 2603 3987
rect 2391 3975 2395 3979
rect 2551 3975 2555 3979
rect 3883 3983 3887 3987
rect 2703 3975 2707 3979
rect 2847 3975 2851 3979
rect 2983 3975 2987 3979
rect 3119 3975 3123 3979
rect 3247 3975 3251 3979
rect 3367 3975 3371 3979
rect 3479 3975 3483 3979
rect 3599 3975 3603 3979
rect 3719 3975 3723 3979
rect 3839 3975 3843 3979
rect 1075 3963 1079 3967
rect 1503 3963 1507 3967
rect 1511 3959 1515 3963
rect 2415 3963 2419 3967
rect 2727 3963 2731 3967
rect 2951 3967 2955 3971
rect 111 3952 115 3956
rect 2031 3952 2035 3956
rect 2071 3956 2075 3960
rect 3991 3956 3995 3960
rect 111 3935 115 3939
rect 2031 3935 2035 3939
rect 2071 3939 2075 3943
rect 3991 3939 3995 3943
rect 175 3930 179 3934
rect 383 3930 387 3934
rect 591 3930 595 3934
rect 791 3930 795 3934
rect 983 3930 987 3934
rect 1167 3930 1171 3934
rect 1343 3930 1347 3934
rect 1519 3930 1523 3934
rect 2231 3934 2235 3938
rect 1703 3930 1707 3934
rect 2391 3934 2395 3938
rect 2551 3934 2555 3938
rect 2703 3934 2707 3938
rect 2847 3934 2851 3938
rect 2983 3934 2987 3938
rect 3119 3934 3123 3938
rect 3247 3934 3251 3938
rect 3367 3934 3371 3938
rect 3479 3934 3483 3938
rect 3599 3934 3603 3938
rect 3719 3934 3723 3938
rect 3839 3934 3843 3938
rect 359 3898 363 3902
rect 551 3898 555 3902
rect 735 3898 739 3902
rect 919 3898 923 3902
rect 1087 3898 1091 3902
rect 1247 3898 1251 3902
rect 1399 3898 1403 3902
rect 1543 3898 1547 3902
rect 1679 3898 1683 3902
rect 1815 3898 1819 3902
rect 2223 3902 2227 3906
rect 1935 3898 1939 3902
rect 2455 3902 2459 3906
rect 2671 3902 2675 3906
rect 2879 3902 2883 3906
rect 3071 3902 3075 3906
rect 3247 3902 3251 3906
rect 3415 3902 3419 3906
rect 3583 3902 3587 3906
rect 3751 3902 3755 3906
rect 111 3893 115 3897
rect 2031 3893 2035 3897
rect 2071 3897 2075 3901
rect 3991 3897 3995 3901
rect 111 3876 115 3880
rect 2031 3876 2035 3880
rect 2071 3880 2075 3884
rect 3991 3880 3995 3884
rect 535 3867 539 3871
rect 359 3857 363 3861
rect 551 3857 555 3861
rect 719 3855 723 3859
rect 735 3857 739 3861
rect 919 3857 923 3861
rect 1087 3857 1091 3861
rect 1663 3867 1667 3871
rect 1799 3867 1803 3871
rect 1903 3867 1907 3871
rect 2007 3867 2011 3871
rect 2295 3871 2299 3875
rect 2527 3871 2531 3875
rect 3055 3871 3059 3875
rect 3735 3871 3739 3875
rect 3883 3871 3887 3875
rect 1247 3857 1251 3861
rect 1399 3857 1403 3861
rect 1543 3857 1547 3861
rect 1679 3857 1683 3861
rect 1815 3857 1819 3861
rect 1935 3857 1939 3861
rect 2223 3861 2227 3865
rect 2455 3861 2459 3865
rect 2671 3861 2675 3865
rect 2879 3861 2883 3865
rect 3071 3861 3075 3865
rect 3247 3861 3251 3865
rect 3415 3861 3419 3865
rect 3583 3861 3587 3865
rect 3751 3861 3755 3865
rect 1511 3847 1515 3851
rect 1663 3847 1667 3851
rect 1799 3847 1803 3851
rect 1903 3847 1907 3851
rect 2255 3851 2259 3855
rect 2727 3851 2731 3855
rect 2951 3851 2952 3855
rect 2952 3851 2955 3855
rect 3487 3851 3488 3855
rect 3488 3851 3491 3855
rect 3511 3851 3515 3855
rect 3735 3851 3739 3855
rect 1103 3835 1104 3839
rect 1104 3835 1107 3839
rect 2007 3835 2008 3839
rect 2008 3835 2011 3839
rect 2263 3839 2264 3843
rect 2264 3839 2267 3843
rect 2527 3839 2531 3843
rect 583 3827 587 3831
rect 735 3827 739 3831
rect 887 3827 891 3831
rect 1031 3827 1035 3831
rect 1175 3827 1179 3831
rect 1311 3827 1315 3831
rect 1447 3827 1451 3831
rect 1575 3827 1579 3831
rect 1703 3827 1707 3831
rect 1831 3827 1835 3831
rect 1935 3827 1939 3831
rect 2191 3831 2195 3835
rect 2487 3831 2491 3835
rect 2759 3831 2763 3835
rect 719 3819 723 3823
rect 1295 3819 1299 3823
rect 2255 3823 2259 3827
rect 2631 3823 2635 3827
rect 2999 3831 3003 3835
rect 3647 3839 3651 3843
rect 3215 3831 3219 3835
rect 3407 3831 3411 3835
rect 3583 3831 3587 3835
rect 3751 3831 3755 3835
rect 3391 3823 3395 3827
rect 3511 3823 3515 3827
rect 3895 3831 3899 3835
rect 3967 3823 3971 3827
rect 111 3808 115 3812
rect 2031 3808 2035 3812
rect 2071 3812 2075 3816
rect 3991 3812 3995 3816
rect 111 3791 115 3795
rect 2031 3791 2035 3795
rect 2071 3795 2075 3799
rect 3991 3795 3995 3799
rect 583 3786 587 3790
rect 735 3786 739 3790
rect 887 3786 891 3790
rect 1031 3786 1035 3790
rect 1175 3786 1179 3790
rect 1311 3786 1315 3790
rect 1447 3786 1451 3790
rect 1575 3786 1579 3790
rect 1703 3786 1707 3790
rect 1831 3786 1835 3790
rect 2191 3790 2195 3794
rect 1935 3786 1939 3790
rect 2487 3790 2491 3794
rect 2759 3790 2763 3794
rect 2999 3790 3003 3794
rect 3215 3790 3219 3794
rect 3407 3790 3411 3794
rect 3583 3790 3587 3794
rect 3751 3790 3755 3794
rect 3895 3790 3899 3794
rect 3391 3775 3395 3779
rect 3551 3775 3555 3779
rect 1295 3759 1299 3763
rect 1839 3759 1843 3763
rect 2111 3758 2115 3762
rect 2335 3758 2339 3762
rect 2559 3758 2563 3762
rect 2775 3758 2779 3762
rect 2975 3758 2979 3762
rect 3159 3758 3163 3762
rect 3327 3758 3331 3762
rect 3479 3758 3483 3762
rect 3623 3758 3627 3762
rect 3767 3758 3771 3762
rect 3895 3758 3899 3762
rect 2071 3753 2075 3757
rect 3991 3753 3995 3757
rect 599 3742 603 3746
rect 719 3742 723 3746
rect 847 3742 851 3746
rect 983 3742 987 3746
rect 1111 3742 1115 3746
rect 1239 3742 1243 3746
rect 1367 3742 1371 3746
rect 1495 3742 1499 3746
rect 1631 3742 1635 3746
rect 1767 3742 1771 3746
rect 111 3737 115 3741
rect 2031 3737 2035 3741
rect 2071 3736 2075 3740
rect 3991 3736 3995 3740
rect 2263 3727 2267 3731
rect 2699 3727 2703 3731
rect 2887 3727 2891 3731
rect 3143 3727 3147 3731
rect 3647 3727 3651 3731
rect 111 3720 115 3724
rect 2031 3720 2035 3724
rect 2111 3717 2115 3721
rect 2335 3717 2339 3721
rect 2559 3717 2563 3721
rect 2775 3717 2779 3721
rect 2975 3717 2979 3721
rect 3159 3717 3163 3721
rect 3327 3717 3331 3721
rect 3479 3717 3483 3721
rect 3623 3717 3627 3721
rect 3767 3717 3771 3721
rect 3895 3717 3899 3721
rect 703 3711 707 3715
rect 967 3711 971 3715
rect 1103 3711 1107 3715
rect 1351 3711 1355 3715
rect 2631 3707 2632 3711
rect 2632 3707 2635 3711
rect 2699 3707 2703 3711
rect 3551 3707 3552 3711
rect 3552 3707 3555 3711
rect 3967 3707 3968 3711
rect 3968 3707 3971 3711
rect 599 3701 603 3705
rect 719 3701 723 3705
rect 847 3701 851 3705
rect 983 3701 987 3705
rect 1111 3701 1115 3705
rect 1239 3701 1243 3705
rect 1367 3701 1371 3705
rect 1495 3701 1499 3705
rect 1631 3701 1635 3705
rect 1767 3701 1771 3705
rect 783 3691 787 3695
rect 703 3683 707 3687
rect 967 3691 971 3695
rect 1839 3691 1840 3695
rect 1840 3691 1843 3695
rect 3143 3691 3147 3695
rect 1351 3683 1355 3687
rect 687 3675 688 3679
rect 688 3675 691 3679
rect 911 3675 915 3679
rect 2051 3683 2055 3687
rect 2111 3675 2115 3679
rect 471 3667 475 3671
rect 615 3667 619 3671
rect 759 3667 763 3671
rect 903 3667 907 3671
rect 1047 3667 1051 3671
rect 1191 3667 1195 3671
rect 1335 3667 1339 3671
rect 1479 3667 1483 3671
rect 2887 3683 2888 3687
rect 2888 3683 2891 3687
rect 2255 3675 2259 3679
rect 2439 3675 2443 3679
rect 2623 3675 2627 3679
rect 2815 3675 2819 3679
rect 3007 3675 3011 3679
rect 3199 3675 3203 3679
rect 3391 3675 3395 3679
rect 3583 3675 3587 3679
rect 599 3659 603 3663
rect 783 3655 787 3659
rect 1175 3659 1179 3663
rect 2431 3663 2435 3667
rect 3183 3667 3187 3671
rect 2071 3656 2075 3660
rect 3991 3656 3995 3660
rect 111 3648 115 3652
rect 2031 3648 2035 3652
rect 2071 3639 2075 3643
rect 3991 3639 3995 3643
rect 111 3631 115 3635
rect 2031 3631 2035 3635
rect 2111 3634 2115 3638
rect 2255 3634 2259 3638
rect 2439 3634 2443 3638
rect 2623 3634 2627 3638
rect 2815 3634 2819 3638
rect 3007 3634 3011 3638
rect 3199 3634 3203 3638
rect 3391 3634 3395 3638
rect 3583 3634 3587 3638
rect 471 3626 475 3630
rect 615 3626 619 3630
rect 759 3626 763 3630
rect 903 3626 907 3630
rect 1047 3626 1051 3630
rect 1191 3626 1195 3630
rect 1335 3626 1339 3630
rect 1479 3626 1483 3630
rect 247 3594 251 3598
rect 375 3594 379 3598
rect 519 3594 523 3598
rect 679 3594 683 3598
rect 847 3594 851 3598
rect 1023 3594 1027 3598
rect 1207 3594 1211 3598
rect 1391 3594 1395 3598
rect 1575 3594 1579 3598
rect 1767 3594 1771 3598
rect 1935 3594 1939 3598
rect 111 3589 115 3593
rect 2031 3589 2035 3593
rect 2359 3590 2363 3594
rect 2583 3590 2587 3594
rect 2799 3590 2803 3594
rect 3007 3590 3011 3594
rect 3215 3590 3219 3594
rect 3431 3590 3435 3594
rect 2071 3585 2075 3589
rect 3991 3585 3995 3589
rect 3183 3579 3187 3583
rect 3503 3579 3507 3583
rect 111 3572 115 3576
rect 2031 3572 2035 3576
rect 2071 3568 2075 3572
rect 359 3563 363 3567
rect 663 3563 667 3567
rect 687 3563 691 3567
rect 1039 3563 1043 3567
rect 1751 3563 1755 3567
rect 1879 3563 1883 3567
rect 3991 3568 3995 3572
rect 2051 3563 2055 3567
rect 2567 3559 2571 3563
rect 247 3553 251 3557
rect 375 3553 379 3557
rect 519 3553 523 3557
rect 679 3553 683 3557
rect 847 3553 851 3557
rect 1023 3553 1027 3557
rect 1207 3553 1211 3557
rect 1391 3553 1395 3557
rect 1575 3553 1579 3557
rect 1767 3553 1771 3557
rect 1935 3553 1939 3557
rect 2647 3555 2651 3559
rect 2991 3559 2995 3563
rect 2359 3549 2363 3553
rect 2583 3549 2587 3553
rect 2799 3549 2803 3553
rect 3007 3549 3011 3553
rect 3215 3549 3219 3553
rect 3431 3549 3435 3553
rect 423 3543 427 3547
rect 359 3535 363 3539
rect 1463 3543 1464 3547
rect 1464 3543 1467 3547
rect 1647 3543 1648 3547
rect 1648 3543 1651 3547
rect 1751 3543 1755 3547
rect 1879 3543 1883 3547
rect 663 3535 667 3539
rect 2431 3539 2432 3543
rect 2432 3539 2435 3543
rect 2567 3539 2571 3543
rect 3503 3539 3504 3543
rect 3504 3539 3507 3543
rect 231 3527 235 3531
rect 415 3519 419 3523
rect 951 3527 955 3531
rect 1039 3519 1040 3523
rect 1040 3519 1043 3523
rect 1567 3527 1571 3531
rect 2991 3531 2995 3535
rect 151 3511 155 3515
rect 263 3511 267 3515
rect 399 3511 403 3515
rect 543 3511 547 3515
rect 687 3511 691 3515
rect 831 3511 835 3515
rect 967 3511 971 3515
rect 1095 3511 1099 3515
rect 231 3503 235 3507
rect 423 3499 427 3503
rect 951 3503 955 3507
rect 1223 3511 1227 3515
rect 1535 3519 1536 3523
rect 1536 3519 1539 3523
rect 2647 3523 2648 3527
rect 2648 3523 2651 3527
rect 1343 3511 1347 3515
rect 1463 3511 1467 3515
rect 1583 3511 1587 3515
rect 1711 3511 1715 3515
rect 2439 3515 2443 3519
rect 2575 3515 2579 3519
rect 2703 3515 2707 3519
rect 2831 3515 2835 3519
rect 2951 3515 2955 3519
rect 3071 3515 3075 3519
rect 3199 3515 3203 3519
rect 3327 3515 3331 3519
rect 1447 3503 1451 3507
rect 1567 3503 1571 3507
rect 1647 3503 1651 3507
rect 2431 3503 2435 3507
rect 2787 3507 2791 3511
rect 111 3492 115 3496
rect 2031 3492 2035 3496
rect 2071 3496 2075 3500
rect 3991 3496 3995 3500
rect 111 3475 115 3479
rect 2031 3475 2035 3479
rect 2071 3479 2075 3483
rect 3991 3479 3995 3483
rect 151 3470 155 3474
rect 263 3470 267 3474
rect 399 3470 403 3474
rect 543 3470 547 3474
rect 687 3470 691 3474
rect 831 3470 835 3474
rect 967 3470 971 3474
rect 1095 3470 1099 3474
rect 1223 3470 1227 3474
rect 1343 3470 1347 3474
rect 1463 3470 1467 3474
rect 1583 3470 1587 3474
rect 2439 3474 2443 3478
rect 1711 3470 1715 3474
rect 2575 3474 2579 3478
rect 2703 3474 2707 3478
rect 2831 3474 2835 3478
rect 2951 3474 2955 3478
rect 3071 3474 3075 3478
rect 3199 3474 3203 3478
rect 3327 3474 3331 3478
rect 151 3438 155 3442
rect 423 3438 427 3442
rect 743 3438 747 3442
rect 1071 3438 1075 3442
rect 2359 3442 2363 3446
rect 1399 3438 1403 3442
rect 2463 3442 2467 3446
rect 2567 3442 2571 3446
rect 2671 3442 2675 3446
rect 2775 3442 2779 3446
rect 2879 3442 2883 3446
rect 2983 3442 2987 3446
rect 3087 3442 3091 3446
rect 3191 3442 3195 3446
rect 111 3433 115 3437
rect 2031 3433 2035 3437
rect 2071 3437 2075 3441
rect 3991 3437 3995 3441
rect 111 3416 115 3420
rect 2031 3416 2035 3420
rect 2071 3420 2075 3424
rect 3991 3420 3995 3424
rect 407 3407 411 3411
rect 415 3407 419 3411
rect 1535 3407 1539 3411
rect 2447 3411 2451 3415
rect 2487 3411 2491 3415
rect 2639 3411 2643 3415
rect 151 3397 155 3401
rect 423 3397 427 3401
rect 743 3397 747 3401
rect 1071 3397 1075 3401
rect 1399 3397 1403 3401
rect 2359 3401 2363 3405
rect 2463 3401 2467 3405
rect 2567 3401 2571 3405
rect 2671 3401 2675 3405
rect 2775 3401 2779 3405
rect 2879 3401 2883 3405
rect 2983 3401 2987 3405
rect 3087 3401 3091 3405
rect 3191 3401 3195 3405
rect 215 3387 219 3391
rect 407 3379 411 3383
rect 1447 3387 1451 3391
rect 2431 3391 2432 3395
rect 2432 3391 2435 3395
rect 2447 3391 2451 3395
rect 2787 3383 2791 3387
rect 2839 3359 2843 3363
rect 995 3351 999 3355
rect 2003 3351 2007 3355
rect 2487 3351 2491 3355
rect 151 3343 155 3347
rect 319 3343 323 3347
rect 527 3343 531 3347
rect 743 3343 747 3347
rect 959 3343 963 3347
rect 1167 3343 1171 3347
rect 1367 3343 1371 3347
rect 1559 3343 1563 3347
rect 1751 3343 1755 3347
rect 1935 3343 1939 3347
rect 2439 3343 2443 3347
rect 215 3335 219 3339
rect 2639 3351 2643 3355
rect 2543 3343 2547 3347
rect 2647 3343 2651 3347
rect 2607 3335 2611 3339
rect 2751 3343 2755 3347
rect 2855 3343 2859 3347
rect 2959 3343 2963 3347
rect 2839 3335 2843 3339
rect 2919 3335 2923 3339
rect 111 3324 115 3328
rect 2031 3324 2035 3328
rect 2071 3324 2075 3328
rect 3991 3324 3995 3328
rect 111 3307 115 3311
rect 2031 3307 2035 3311
rect 151 3302 155 3306
rect 319 3302 323 3306
rect 527 3302 531 3306
rect 743 3302 747 3306
rect 959 3302 963 3306
rect 1167 3302 1171 3306
rect 1367 3302 1371 3306
rect 1559 3302 1563 3306
rect 1751 3302 1755 3306
rect 2071 3307 2075 3311
rect 3991 3307 3995 3311
rect 1935 3302 1939 3306
rect 2439 3302 2443 3306
rect 2543 3302 2547 3306
rect 2647 3302 2651 3306
rect 2751 3302 2755 3306
rect 2855 3302 2859 3306
rect 2959 3302 2963 3306
rect 995 3287 999 3291
rect 2527 3270 2531 3274
rect 2631 3270 2635 3274
rect 2735 3270 2739 3274
rect 2839 3270 2843 3274
rect 2943 3270 2947 3274
rect 3047 3270 3051 3274
rect 3151 3270 3155 3274
rect 3255 3270 3259 3274
rect 311 3262 315 3266
rect 479 3262 483 3266
rect 655 3262 659 3266
rect 847 3262 851 3266
rect 1039 3262 1043 3266
rect 1231 3262 1235 3266
rect 1431 3262 1435 3266
rect 1631 3262 1635 3266
rect 1831 3262 1835 3266
rect 2071 3265 2075 3269
rect 3991 3265 3995 3269
rect 111 3257 115 3261
rect 2031 3257 2035 3261
rect 2071 3248 2075 3252
rect 3991 3248 3995 3252
rect 111 3240 115 3244
rect 2031 3240 2035 3244
rect 2615 3239 2619 3243
rect 2719 3239 2723 3243
rect 3031 3239 3035 3243
rect 1255 3231 1259 3235
rect 2003 3231 2007 3235
rect 2527 3229 2531 3233
rect 2631 3229 2635 3233
rect 2735 3229 2739 3233
rect 2839 3229 2843 3233
rect 2943 3229 2947 3233
rect 3047 3229 3051 3233
rect 3175 3239 3179 3243
rect 3151 3229 3155 3233
rect 3255 3229 3259 3233
rect 311 3221 315 3225
rect 479 3221 483 3225
rect 655 3221 659 3225
rect 847 3221 851 3225
rect 1039 3221 1043 3225
rect 1231 3221 1235 3225
rect 1431 3221 1435 3225
rect 1631 3221 1635 3225
rect 1831 3221 1835 3225
rect 2600 3219 2604 3223
rect 1047 3211 1051 3215
rect 1775 3211 1779 3215
rect 2615 3215 2619 3219
rect 2912 3219 2916 3223
rect 3015 3219 3016 3223
rect 3016 3219 3019 3223
rect 3031 3219 3035 3223
rect 3175 3207 3179 3211
rect 3399 3207 3403 3211
rect 1127 3195 1128 3199
rect 1128 3195 1131 3199
rect 1255 3195 1259 3199
rect 623 3187 627 3191
rect 759 3187 763 3191
rect 903 3187 907 3191
rect 1055 3187 1059 3191
rect 1207 3187 1211 3191
rect 743 3179 747 3183
rect 1351 3187 1355 3191
rect 2007 3195 2008 3199
rect 2008 3195 2011 3199
rect 2399 3199 2403 3203
rect 2551 3199 2555 3203
rect 2695 3199 2699 3203
rect 2839 3199 2843 3203
rect 2975 3199 2979 3203
rect 3111 3199 3115 3203
rect 3247 3199 3251 3203
rect 3391 3199 3395 3203
rect 1503 3187 1507 3191
rect 1655 3187 1659 3191
rect 1807 3187 1811 3191
rect 1935 3187 1939 3191
rect 2415 3187 2419 3191
rect 2959 3191 2963 3195
rect 3263 3187 3267 3191
rect 1639 3179 1643 3183
rect 1775 3179 1779 3183
rect 2071 3180 2075 3184
rect 3991 3180 3995 3184
rect 111 3168 115 3172
rect 2031 3168 2035 3172
rect 2071 3163 2075 3167
rect 3991 3163 3995 3167
rect 2399 3158 2403 3162
rect 2551 3158 2555 3162
rect 2695 3158 2699 3162
rect 2839 3158 2843 3162
rect 2975 3158 2979 3162
rect 3111 3158 3115 3162
rect 3247 3158 3251 3162
rect 3391 3158 3395 3162
rect 111 3151 115 3155
rect 2031 3151 2035 3155
rect 623 3146 627 3150
rect 759 3146 763 3150
rect 903 3146 907 3150
rect 1055 3146 1059 3150
rect 1207 3146 1211 3150
rect 1351 3146 1355 3150
rect 1503 3146 1507 3150
rect 1655 3146 1659 3150
rect 1807 3146 1811 3150
rect 1935 3146 1939 3150
rect 599 3114 603 3118
rect 703 3114 707 3118
rect 807 3114 811 3118
rect 911 3114 915 3118
rect 1039 3114 1043 3118
rect 1183 3114 1187 3118
rect 1359 3114 1363 3118
rect 1551 3114 1555 3118
rect 1751 3114 1755 3118
rect 1935 3114 1939 3118
rect 2111 3114 2115 3118
rect 111 3109 115 3113
rect 2031 3109 2035 3113
rect 2343 3114 2347 3118
rect 2583 3114 2587 3118
rect 2799 3114 2803 3118
rect 2999 3114 3003 3118
rect 3191 3114 3195 3118
rect 3375 3114 3379 3118
rect 3567 3114 3571 3118
rect 2071 3109 2075 3113
rect 3991 3109 3995 3113
rect 111 3092 115 3096
rect 2031 3092 2035 3096
rect 2071 3092 2075 3096
rect 3991 3092 3995 3096
rect 687 3083 691 3087
rect 791 3083 795 3087
rect 895 3083 899 3087
rect 1023 3083 1027 3087
rect 1127 3083 1131 3087
rect 2007 3083 2011 3087
rect 2567 3083 2571 3087
rect 2663 3083 2667 3087
rect 2983 3083 2987 3087
rect 3551 3083 3555 3087
rect 3663 3083 3667 3087
rect 599 3073 603 3077
rect 703 3073 707 3077
rect 807 3073 811 3077
rect 911 3073 915 3077
rect 1039 3073 1043 3077
rect 1183 3073 1187 3077
rect 1359 3073 1363 3077
rect 1551 3073 1555 3077
rect 1639 3071 1643 3075
rect 1751 3073 1755 3077
rect 1935 3073 1939 3077
rect 2111 3073 2115 3077
rect 2343 3073 2347 3077
rect 2583 3073 2587 3077
rect 2799 3073 2803 3077
rect 2999 3073 3003 3077
rect 3191 3073 3195 3077
rect 3375 3073 3379 3077
rect 3567 3073 3571 3077
rect 663 3063 667 3067
rect 687 3063 691 3067
rect 791 3063 795 3067
rect 895 3063 899 3067
rect 1023 3063 1027 3067
rect 1167 3063 1168 3067
rect 1168 3063 1171 3067
rect 2175 3063 2179 3067
rect 2415 3063 2416 3067
rect 2416 3063 2419 3067
rect 2567 3063 2571 3067
rect 3263 3063 3264 3067
rect 3264 3063 3267 3067
rect 399 3051 403 3055
rect 311 3035 315 3039
rect 415 3035 419 3039
rect 527 3035 531 3039
rect 599 3039 603 3043
rect 959 3051 963 3055
rect 2983 3055 2987 3059
rect 3551 3063 3555 3067
rect 1167 3043 1168 3047
rect 1168 3043 1171 3047
rect 2527 3047 2528 3051
rect 2528 3047 2531 3051
rect 2663 3047 2667 3051
rect 639 3035 643 3039
rect 751 3035 755 3039
rect 863 3035 867 3039
rect 975 3035 979 3039
rect 1095 3035 1099 3039
rect 1215 3035 1219 3039
rect 1335 3035 1339 3039
rect 2111 3039 2115 3043
rect 2263 3039 2267 3043
rect 2455 3039 2459 3043
rect 2655 3039 2659 3043
rect 399 3027 403 3031
rect 663 3023 667 3027
rect 959 3027 963 3031
rect 2175 3031 2179 3035
rect 3663 3047 3667 3051
rect 2855 3039 2859 3043
rect 3055 3039 3059 3043
rect 3255 3039 3259 3043
rect 3455 3039 3459 3043
rect 3655 3039 3659 3043
rect 2919 3031 2923 3035
rect 3151 3031 3155 3035
rect 1207 3023 1211 3027
rect 111 3016 115 3020
rect 2031 3016 2035 3020
rect 2071 3020 2075 3024
rect 3991 3020 3995 3024
rect 111 2999 115 3003
rect 2031 2999 2035 3003
rect 2071 3003 2075 3007
rect 3991 3003 3995 3007
rect 311 2994 315 2998
rect 415 2994 419 2998
rect 527 2994 531 2998
rect 639 2994 643 2998
rect 751 2994 755 2998
rect 863 2994 867 2998
rect 975 2994 979 2998
rect 1095 2994 1099 2998
rect 1215 2994 1219 2998
rect 2111 2998 2115 3002
rect 1335 2994 1339 2998
rect 2263 2998 2267 3002
rect 2455 2998 2459 3002
rect 2655 2998 2659 3002
rect 2855 2998 2859 3002
rect 3055 2998 3059 3002
rect 3255 2998 3259 3002
rect 3455 2998 3459 3002
rect 3655 2998 3659 3002
rect 2339 2983 2343 2987
rect 2527 2983 2531 2987
rect 2111 2966 2115 2970
rect 2359 2966 2363 2970
rect 2607 2966 2611 2970
rect 2847 2966 2851 2970
rect 3079 2966 3083 2970
rect 3303 2966 3307 2970
rect 3535 2966 3539 2970
rect 3767 2966 3771 2970
rect 2071 2961 2075 2965
rect 3991 2961 3995 2965
rect 151 2954 155 2958
rect 271 2954 275 2958
rect 431 2954 435 2958
rect 607 2954 611 2958
rect 783 2954 787 2958
rect 959 2954 963 2958
rect 1135 2954 1139 2958
rect 1303 2954 1307 2958
rect 1471 2954 1475 2958
rect 1647 2954 1651 2958
rect 111 2949 115 2953
rect 2031 2949 2035 2953
rect 2071 2944 2075 2948
rect 3991 2944 3995 2948
rect 111 2932 115 2936
rect 2031 2932 2035 2936
rect 2339 2935 2343 2939
rect 3287 2935 3291 2939
rect 3519 2935 3523 2939
rect 3751 2935 3755 2939
rect 231 2923 235 2927
rect 599 2923 603 2927
rect 983 2923 987 2927
rect 1267 2923 1271 2927
rect 1455 2923 1459 2927
rect 1631 2923 1635 2927
rect 1719 2923 1723 2927
rect 2111 2925 2115 2929
rect 2359 2925 2363 2929
rect 2423 2923 2427 2927
rect 2607 2925 2611 2929
rect 2847 2925 2851 2929
rect 3079 2925 3083 2929
rect 3303 2925 3307 2929
rect 3535 2925 3539 2929
rect 3767 2925 3771 2929
rect 151 2913 155 2917
rect 271 2913 275 2917
rect 431 2913 435 2917
rect 607 2913 611 2917
rect 783 2913 787 2917
rect 959 2913 963 2917
rect 1135 2913 1139 2917
rect 1303 2913 1307 2917
rect 1471 2913 1475 2917
rect 1647 2913 1651 2917
rect 2435 2915 2436 2919
rect 2436 2915 2439 2919
rect 2919 2915 2920 2919
rect 2920 2915 2923 2919
rect 3151 2915 3152 2919
rect 3152 2915 3155 2919
rect 3287 2915 3291 2919
rect 3519 2915 3523 2919
rect 3751 2915 3755 2919
rect 515 2903 519 2907
rect 231 2895 235 2899
rect 1035 2903 1036 2907
rect 1036 2903 1039 2907
rect 1207 2903 1208 2907
rect 1208 2903 1211 2907
rect 1267 2903 1271 2907
rect 1455 2903 1459 2907
rect 1631 2903 1635 2907
rect 2423 2895 2427 2899
rect 2435 2895 2439 2899
rect 2975 2895 2976 2899
rect 2976 2895 2979 2899
rect 2111 2887 2115 2891
rect 2279 2887 2283 2891
rect 2487 2887 2491 2891
rect 2695 2887 2699 2891
rect 2903 2887 2907 2891
rect 3111 2887 3115 2891
rect 3303 2887 3307 2891
rect 3495 2887 3499 2891
rect 3687 2887 3691 2891
rect 3879 2887 3883 2891
rect 223 2879 224 2883
rect 224 2879 227 2883
rect 151 2871 155 2875
rect 287 2871 291 2875
rect 983 2879 987 2883
rect 1035 2879 1039 2883
rect 1535 2879 1539 2883
rect 1719 2879 1723 2883
rect 2231 2879 2235 2883
rect 3287 2879 3291 2883
rect 447 2871 451 2875
rect 599 2871 603 2875
rect 759 2871 763 2875
rect 927 2871 931 2875
rect 1103 2871 1107 2875
rect 1287 2871 1291 2875
rect 1479 2871 1483 2875
rect 1671 2871 1675 2875
rect 2071 2868 2075 2872
rect 3991 2868 3995 2872
rect 515 2863 519 2867
rect 591 2859 595 2863
rect 1695 2859 1699 2863
rect 111 2852 115 2856
rect 2031 2852 2035 2856
rect 2071 2851 2075 2855
rect 3991 2851 3995 2855
rect 2111 2846 2115 2850
rect 2279 2846 2283 2850
rect 2487 2846 2491 2850
rect 2695 2846 2699 2850
rect 2903 2846 2907 2850
rect 3111 2846 3115 2850
rect 3303 2846 3307 2850
rect 3495 2846 3499 2850
rect 3687 2846 3691 2850
rect 3879 2846 3883 2850
rect 111 2835 115 2839
rect 2031 2835 2035 2839
rect 151 2830 155 2834
rect 287 2830 291 2834
rect 447 2830 451 2834
rect 599 2830 603 2834
rect 759 2830 763 2834
rect 927 2830 931 2834
rect 1103 2830 1107 2834
rect 1287 2830 1291 2834
rect 1479 2830 1483 2834
rect 1671 2830 1675 2834
rect 3287 2819 3291 2823
rect 3839 2819 3843 2823
rect 2143 2802 2147 2806
rect 2319 2802 2323 2806
rect 2503 2802 2507 2806
rect 2695 2802 2699 2806
rect 2887 2802 2891 2806
rect 3079 2802 3083 2806
rect 3263 2802 3267 2806
rect 3439 2802 3443 2806
rect 3615 2802 3619 2806
rect 3791 2802 3795 2806
rect 2071 2797 2075 2801
rect 3991 2797 3995 2801
rect 151 2786 155 2790
rect 319 2786 323 2790
rect 503 2786 507 2790
rect 687 2786 691 2790
rect 871 2786 875 2790
rect 1055 2786 1059 2790
rect 1239 2786 1243 2790
rect 1431 2786 1435 2790
rect 1631 2786 1635 2790
rect 1831 2786 1835 2790
rect 111 2781 115 2785
rect 2031 2781 2035 2785
rect 2071 2780 2075 2784
rect 3991 2780 3995 2784
rect 2167 2771 2171 2775
rect 2679 2771 2683 2775
rect 2871 2771 2875 2775
rect 2975 2771 2979 2775
rect 3247 2771 3251 2775
rect 111 2764 115 2768
rect 2031 2764 2035 2768
rect 2143 2761 2147 2765
rect 223 2755 227 2759
rect 671 2755 675 2759
rect 151 2745 155 2749
rect 319 2745 323 2749
rect 503 2745 507 2749
rect 687 2745 691 2749
rect 1223 2755 1227 2759
rect 1415 2755 1419 2759
rect 1535 2755 1539 2759
rect 1815 2755 1819 2759
rect 1903 2755 1907 2759
rect 2231 2759 2235 2763
rect 2319 2761 2323 2765
rect 2503 2761 2507 2765
rect 2695 2761 2699 2765
rect 2887 2761 2891 2765
rect 3079 2761 3083 2765
rect 3263 2761 3267 2765
rect 3439 2761 3443 2765
rect 3615 2761 3619 2765
rect 3791 2761 3795 2765
rect 2519 2751 2523 2755
rect 2679 2751 2683 2755
rect 2871 2751 2875 2755
rect 3839 2751 3843 2755
rect 871 2745 875 2749
rect 1055 2745 1059 2749
rect 1239 2745 1243 2749
rect 1431 2745 1435 2749
rect 1631 2745 1635 2749
rect 1831 2745 1835 2749
rect 391 2735 392 2739
rect 392 2735 395 2739
rect 591 2735 595 2739
rect 671 2735 675 2739
rect 1047 2735 1051 2739
rect 1223 2735 1227 2739
rect 1415 2735 1419 2739
rect 1695 2735 1699 2739
rect 1815 2735 1819 2739
rect 3247 2735 3251 2739
rect 2167 2727 2171 2731
rect 247 2719 251 2723
rect 183 2711 187 2715
rect 1647 2719 1651 2723
rect 1903 2719 1907 2723
rect 2111 2719 2115 2723
rect 383 2711 387 2715
rect 583 2711 587 2715
rect 783 2711 787 2715
rect 983 2711 987 2715
rect 1199 2711 1203 2715
rect 1415 2711 1419 2715
rect 1639 2711 1643 2715
rect 1871 2711 1875 2715
rect 2863 2727 2867 2731
rect 2279 2719 2283 2723
rect 2455 2719 2459 2723
rect 2639 2719 2643 2723
rect 2815 2719 2819 2723
rect 2983 2719 2987 2723
rect 3143 2719 3147 2723
rect 3303 2719 3307 2723
rect 3463 2719 3467 2723
rect 3623 2719 3627 2723
rect 2343 2711 2347 2715
rect 2519 2711 2523 2715
rect 3127 2711 3131 2715
rect 391 2699 395 2703
rect 671 2703 675 2707
rect 1047 2703 1051 2707
rect 1999 2703 2003 2707
rect 2071 2700 2075 2704
rect 3991 2700 3995 2704
rect 111 2692 115 2696
rect 2031 2692 2035 2696
rect 2071 2683 2075 2687
rect 3991 2683 3995 2687
rect 111 2675 115 2679
rect 2031 2675 2035 2679
rect 2111 2678 2115 2682
rect 2279 2678 2283 2682
rect 2455 2678 2459 2682
rect 2639 2678 2643 2682
rect 2815 2678 2819 2682
rect 2983 2678 2987 2682
rect 3143 2678 3147 2682
rect 3303 2678 3307 2682
rect 3463 2678 3467 2682
rect 3623 2678 3627 2682
rect 183 2670 187 2674
rect 383 2670 387 2674
rect 583 2670 587 2674
rect 783 2670 787 2674
rect 983 2670 987 2674
rect 1199 2670 1203 2674
rect 1415 2670 1419 2674
rect 1639 2670 1643 2674
rect 1871 2670 1875 2674
rect 255 2630 259 2634
rect 423 2630 427 2634
rect 599 2630 603 2634
rect 775 2630 779 2634
rect 959 2630 963 2634
rect 1151 2630 1155 2634
rect 1343 2630 1347 2634
rect 1535 2630 1539 2634
rect 1727 2630 1731 2634
rect 2111 2634 2115 2638
rect 1927 2630 1931 2634
rect 2263 2634 2267 2638
rect 2431 2634 2435 2638
rect 2599 2634 2603 2638
rect 2751 2634 2755 2638
rect 2895 2634 2899 2638
rect 3039 2634 3043 2638
rect 3175 2634 3179 2638
rect 3311 2634 3315 2638
rect 3455 2634 3459 2638
rect 111 2625 115 2629
rect 2031 2625 2035 2629
rect 2071 2629 2075 2633
rect 3991 2629 3995 2633
rect 1223 2619 1227 2623
rect 1647 2619 1651 2623
rect 111 2608 115 2612
rect 2031 2608 2035 2612
rect 2071 2612 2075 2616
rect 3991 2612 3995 2616
rect 247 2599 251 2603
rect 255 2589 259 2593
rect 423 2589 427 2593
rect 599 2589 603 2593
rect 799 2599 803 2603
rect 1223 2599 1227 2603
rect 1799 2599 1803 2603
rect 2183 2603 2187 2607
rect 2583 2603 2587 2607
rect 2863 2603 2867 2607
rect 3023 2603 3027 2607
rect 775 2589 779 2593
rect 959 2589 963 2593
rect 1151 2589 1155 2593
rect 1343 2589 1347 2593
rect 1535 2589 1539 2593
rect 1727 2589 1731 2593
rect 1927 2589 1931 2593
rect 2111 2593 2115 2597
rect 2263 2593 2267 2597
rect 2431 2593 2435 2597
rect 2599 2593 2603 2597
rect 2751 2593 2755 2597
rect 2895 2593 2899 2597
rect 3039 2593 3043 2597
rect 3175 2593 3179 2597
rect 3311 2593 3315 2597
rect 3455 2593 3459 2597
rect 431 2563 435 2567
rect 671 2579 672 2583
rect 672 2579 675 2583
rect 1583 2579 1587 2583
rect 1999 2579 2000 2583
rect 2000 2579 2003 2583
rect 2336 2583 2340 2587
rect 2683 2583 2687 2587
rect 319 2555 323 2559
rect 799 2563 803 2567
rect 535 2555 539 2559
rect 743 2555 747 2559
rect 1455 2563 1459 2567
rect 2583 2575 2587 2579
rect 3527 2583 3528 2587
rect 3528 2583 3531 2587
rect 1799 2563 1803 2567
rect 2183 2563 2184 2567
rect 2184 2563 2187 2567
rect 2539 2563 2543 2567
rect 3023 2571 3027 2575
rect 951 2555 955 2559
rect 1159 2555 1163 2559
rect 1359 2555 1363 2559
rect 1559 2555 1563 2559
rect 1759 2555 1763 2559
rect 1935 2555 1939 2559
rect 2111 2555 2115 2559
rect 2271 2555 2275 2559
rect 2447 2555 2451 2559
rect 2615 2555 2619 2559
rect 2767 2555 2771 2559
rect 2911 2555 2915 2559
rect 3047 2555 3051 2559
rect 3183 2555 3187 2559
rect 3319 2555 3323 2559
rect 1031 2547 1035 2551
rect 1583 2543 1587 2547
rect 1859 2547 1863 2551
rect 2007 2547 2011 2551
rect 2683 2547 2687 2551
rect 2895 2547 2899 2551
rect 111 2536 115 2540
rect 2031 2536 2035 2540
rect 2071 2536 2075 2540
rect 3991 2536 3995 2540
rect 111 2519 115 2523
rect 2031 2519 2035 2523
rect 319 2514 323 2518
rect 535 2514 539 2518
rect 743 2514 747 2518
rect 951 2514 955 2518
rect 1159 2514 1163 2518
rect 1359 2514 1363 2518
rect 1559 2514 1563 2518
rect 1759 2514 1763 2518
rect 2071 2519 2075 2523
rect 3991 2519 3995 2523
rect 1935 2514 1939 2518
rect 2111 2514 2115 2518
rect 2271 2514 2275 2518
rect 2447 2514 2451 2518
rect 2615 2514 2619 2518
rect 2767 2514 2771 2518
rect 2911 2514 2915 2518
rect 3047 2514 3051 2518
rect 3183 2514 3187 2518
rect 3319 2514 3323 2518
rect 279 2482 283 2486
rect 439 2482 443 2486
rect 607 2482 611 2486
rect 783 2482 787 2486
rect 959 2482 963 2486
rect 1127 2482 1131 2486
rect 1295 2482 1299 2486
rect 1463 2482 1467 2486
rect 1623 2482 1627 2486
rect 1791 2482 1795 2486
rect 1935 2482 1939 2486
rect 111 2477 115 2481
rect 2031 2477 2035 2481
rect 2623 2470 2627 2474
rect 2743 2470 2747 2474
rect 2871 2470 2875 2474
rect 3015 2470 3019 2474
rect 3159 2470 3163 2474
rect 3311 2470 3315 2474
rect 3463 2470 3467 2474
rect 3615 2470 3619 2474
rect 3767 2470 3771 2474
rect 3895 2470 3899 2474
rect 2071 2465 2075 2469
rect 111 2460 115 2464
rect 3991 2465 3995 2469
rect 2031 2460 2035 2464
rect 419 2451 423 2455
rect 431 2451 435 2455
rect 679 2451 683 2455
rect 1279 2451 1283 2455
rect 1455 2451 1459 2455
rect 1695 2451 1699 2455
rect 2071 2448 2075 2452
rect 3991 2448 3995 2452
rect 279 2441 283 2445
rect 439 2441 443 2445
rect 607 2441 611 2445
rect 783 2441 787 2445
rect 959 2441 963 2445
rect 1127 2441 1131 2445
rect 1295 2441 1299 2445
rect 1463 2441 1467 2445
rect 1623 2441 1627 2445
rect 1791 2441 1795 2445
rect 1935 2441 1939 2445
rect 2539 2439 2543 2443
rect 2943 2439 2947 2443
rect 3567 2439 3571 2443
rect 3879 2439 3883 2443
rect 3967 2439 3971 2443
rect 351 2431 352 2435
rect 352 2431 355 2435
rect 419 2431 423 2435
rect 1031 2431 1032 2435
rect 1032 2431 1035 2435
rect 1371 2431 1372 2435
rect 1372 2431 1375 2435
rect 1279 2423 1283 2427
rect 1859 2431 1863 2435
rect 1891 2431 1895 2435
rect 2007 2431 2008 2435
rect 2008 2431 2011 2435
rect 2623 2429 2627 2433
rect 2743 2429 2747 2433
rect 2871 2429 2875 2433
rect 3015 2429 3019 2433
rect 3159 2429 3163 2433
rect 3311 2429 3315 2433
rect 3463 2429 3467 2433
rect 3615 2429 3619 2433
rect 3767 2429 3771 2433
rect 3895 2429 3899 2433
rect 2791 2419 2795 2423
rect 679 2411 683 2415
rect 1007 2411 1011 2415
rect 327 2403 331 2407
rect 471 2403 475 2407
rect 623 2403 627 2407
rect 783 2403 787 2407
rect 943 2403 947 2407
rect 1095 2403 1099 2407
rect 1371 2411 1375 2415
rect 351 2391 355 2395
rect 687 2395 691 2399
rect 1247 2403 1251 2407
rect 1695 2411 1699 2415
rect 1891 2411 1892 2415
rect 1892 2411 1895 2415
rect 1391 2403 1395 2407
rect 1535 2403 1539 2407
rect 1671 2403 1675 2407
rect 1815 2403 1819 2407
rect 2895 2411 2899 2415
rect 3687 2419 3688 2423
rect 3688 2419 3691 2423
rect 3567 2411 3571 2415
rect 3879 2419 3883 2423
rect 1935 2403 1939 2407
rect 2583 2403 2587 2407
rect 1527 2391 1531 2395
rect 2007 2395 2011 2399
rect 2663 2395 2667 2399
rect 3039 2403 3043 2407
rect 2943 2395 2947 2399
rect 3967 2395 3968 2399
rect 3968 2395 3971 2399
rect 111 2384 115 2388
rect 2031 2384 2035 2388
rect 2487 2387 2491 2391
rect 2599 2387 2603 2391
rect 2727 2387 2731 2391
rect 2879 2387 2883 2391
rect 3055 2387 3059 2391
rect 3247 2387 3251 2391
rect 3455 2387 3459 2391
rect 3679 2387 3683 2391
rect 3895 2387 3899 2391
rect 2583 2379 2587 2383
rect 2791 2379 2795 2383
rect 3039 2379 3043 2383
rect 3119 2379 3123 2383
rect 3687 2375 3691 2379
rect 3959 2379 3963 2383
rect 111 2367 115 2371
rect 2031 2367 2035 2371
rect 2071 2368 2075 2372
rect 3991 2368 3995 2372
rect 327 2362 331 2366
rect 471 2362 475 2366
rect 623 2362 627 2366
rect 783 2362 787 2366
rect 943 2362 947 2366
rect 1095 2362 1099 2366
rect 1247 2362 1251 2366
rect 1391 2362 1395 2366
rect 1535 2362 1539 2366
rect 1671 2362 1675 2366
rect 1815 2362 1819 2366
rect 1935 2362 1939 2366
rect 2071 2351 2075 2355
rect 3991 2351 3995 2355
rect 2487 2346 2491 2350
rect 2599 2346 2603 2350
rect 2727 2346 2731 2350
rect 2879 2346 2883 2350
rect 3055 2346 3059 2350
rect 3247 2346 3251 2350
rect 3455 2346 3459 2350
rect 3679 2346 3683 2350
rect 3895 2346 3899 2350
rect 359 2322 363 2326
rect 495 2322 499 2326
rect 639 2322 643 2326
rect 783 2322 787 2326
rect 935 2322 939 2326
rect 1087 2322 1091 2326
rect 1247 2322 1251 2326
rect 1415 2322 1419 2326
rect 1591 2322 1595 2326
rect 1775 2322 1779 2326
rect 1935 2322 1939 2326
rect 111 2317 115 2321
rect 2031 2317 2035 2321
rect 111 2300 115 2304
rect 2031 2300 2035 2304
rect 2111 2302 2115 2306
rect 2223 2302 2227 2306
rect 2359 2302 2363 2306
rect 2511 2302 2515 2306
rect 2671 2302 2675 2306
rect 2847 2302 2851 2306
rect 3039 2302 3043 2306
rect 3247 2302 3251 2306
rect 3463 2302 3467 2306
rect 3687 2302 3691 2306
rect 3895 2302 3899 2306
rect 2071 2297 2075 2301
rect 3991 2297 3995 2301
rect 479 2291 483 2295
rect 767 2291 771 2295
rect 919 2291 923 2295
rect 1007 2291 1011 2295
rect 1575 2291 1579 2295
rect 1759 2291 1763 2295
rect 1767 2291 1771 2295
rect 2183 2291 2187 2295
rect 359 2281 363 2285
rect 495 2281 499 2285
rect 639 2281 643 2285
rect 783 2281 787 2285
rect 935 2281 939 2285
rect 1087 2281 1091 2285
rect 1247 2281 1251 2285
rect 1415 2281 1419 2285
rect 1591 2281 1595 2285
rect 1775 2281 1779 2285
rect 1935 2281 1939 2285
rect 2071 2280 2075 2284
rect 3991 2280 3995 2284
rect 687 2271 691 2275
rect 703 2271 707 2275
rect 767 2271 771 2275
rect 919 2271 923 2275
rect 1095 2271 1099 2275
rect 1527 2271 1531 2275
rect 1575 2271 1579 2275
rect 1759 2271 1763 2275
rect 2007 2271 2008 2275
rect 2008 2271 2011 2275
rect 2111 2261 2115 2265
rect 2495 2271 2499 2275
rect 2655 2271 2659 2275
rect 2663 2271 2667 2275
rect 3023 2271 3027 2275
rect 3967 2271 3971 2275
rect 2223 2261 2227 2265
rect 2359 2261 2363 2265
rect 2511 2261 2515 2265
rect 2671 2261 2675 2265
rect 2847 2261 2851 2265
rect 3039 2261 3043 2265
rect 3247 2261 3251 2265
rect 3463 2261 3467 2265
rect 3687 2261 3691 2265
rect 3895 2261 3899 2265
rect 479 2255 483 2259
rect 919 2247 923 2251
rect 1407 2247 1411 2251
rect 1767 2247 1768 2251
rect 1768 2247 1771 2251
rect 2183 2251 2184 2255
rect 2184 2251 2187 2255
rect 2435 2251 2436 2255
rect 2436 2251 2439 2255
rect 2495 2251 2499 2255
rect 2655 2251 2659 2255
rect 3112 2251 3116 2255
rect 3155 2251 3159 2255
rect 239 2239 243 2243
rect 391 2239 395 2243
rect 551 2239 555 2243
rect 711 2239 715 2243
rect 871 2239 875 2243
rect 1031 2239 1035 2243
rect 1191 2239 1195 2243
rect 1359 2239 1363 2243
rect 1527 2239 1531 2243
rect 1695 2239 1699 2243
rect 3023 2243 3027 2247
rect 3771 2251 3775 2255
rect 3959 2251 3963 2255
rect 223 2231 227 2235
rect 703 2231 707 2235
rect 1095 2231 1099 2235
rect 1535 2227 1539 2231
rect 111 2220 115 2224
rect 2031 2220 2035 2224
rect 2111 2223 2115 2227
rect 2435 2231 2439 2235
rect 2687 2231 2691 2235
rect 3155 2231 3156 2235
rect 3156 2231 3159 2235
rect 2279 2223 2283 2227
rect 2479 2223 2483 2227
rect 2679 2223 2683 2227
rect 2879 2223 2883 2227
rect 3079 2223 3083 2227
rect 3259 2227 3263 2231
rect 3279 2223 3283 2227
rect 2391 2215 2395 2219
rect 3063 2215 3067 2219
rect 3719 2231 3723 2235
rect 3967 2231 3968 2235
rect 3968 2231 3971 2235
rect 3487 2223 3491 2227
rect 3703 2223 3707 2227
rect 3895 2223 3899 2227
rect 3479 2211 3483 2215
rect 3771 2215 3775 2219
rect 3959 2215 3963 2219
rect 111 2203 115 2207
rect 2031 2203 2035 2207
rect 2071 2204 2075 2208
rect 3991 2204 3995 2208
rect 239 2198 243 2202
rect 391 2198 395 2202
rect 551 2198 555 2202
rect 711 2198 715 2202
rect 871 2198 875 2202
rect 1031 2198 1035 2202
rect 1191 2198 1195 2202
rect 1359 2198 1363 2202
rect 1527 2198 1531 2202
rect 1695 2198 1699 2202
rect 2071 2187 2075 2191
rect 3991 2187 3995 2191
rect 2111 2182 2115 2186
rect 2279 2182 2283 2186
rect 2479 2182 2483 2186
rect 2679 2182 2683 2186
rect 2879 2182 2883 2186
rect 3079 2182 3083 2186
rect 3279 2182 3283 2186
rect 3487 2182 3491 2186
rect 3703 2182 3707 2186
rect 3895 2182 3899 2186
rect 151 2154 155 2158
rect 319 2154 323 2158
rect 511 2154 515 2158
rect 703 2154 707 2158
rect 895 2154 899 2158
rect 1087 2154 1091 2158
rect 1279 2154 1283 2158
rect 1463 2154 1467 2158
rect 1655 2154 1659 2158
rect 1847 2154 1851 2158
rect 111 2149 115 2153
rect 2031 2149 2035 2153
rect 2143 2142 2147 2146
rect 2319 2142 2323 2146
rect 2495 2142 2499 2146
rect 2679 2142 2683 2146
rect 2863 2142 2867 2146
rect 3039 2142 3043 2146
rect 3215 2142 3219 2146
rect 3391 2142 3395 2146
rect 3567 2142 3571 2146
rect 3743 2142 3747 2146
rect 3895 2142 3899 2146
rect 2071 2137 2075 2141
rect 111 2132 115 2136
rect 3991 2137 3995 2141
rect 2031 2132 2035 2136
rect 239 2123 243 2127
rect 451 2123 455 2127
rect 535 2123 539 2127
rect 879 2123 883 2127
rect 919 2123 923 2127
rect 1407 2123 1411 2127
rect 1639 2123 1643 2127
rect 151 2113 155 2117
rect 319 2113 323 2117
rect 511 2113 515 2117
rect 703 2113 707 2117
rect 895 2113 899 2117
rect 1087 2113 1091 2117
rect 1279 2113 1283 2117
rect 1463 2113 1467 2117
rect 1655 2113 1659 2117
rect 2071 2120 2075 2124
rect 1847 2113 1851 2117
rect 223 2103 224 2107
rect 224 2103 227 2107
rect 239 2103 243 2107
rect 451 2103 455 2107
rect 727 2103 731 2107
rect 879 2103 883 2107
rect 1115 2103 1119 2107
rect 1535 2103 1536 2107
rect 1536 2103 1539 2107
rect 1639 2103 1643 2107
rect 1739 2103 1743 2107
rect 2215 2111 2219 2115
rect 2687 2119 2691 2123
rect 3991 2120 3995 2124
rect 3111 2111 3115 2115
rect 3719 2111 3723 2115
rect 3967 2111 3971 2115
rect 2143 2101 2147 2105
rect 2319 2101 2323 2105
rect 2495 2101 2499 2105
rect 2679 2101 2683 2105
rect 2863 2101 2867 2105
rect 3039 2101 3043 2105
rect 3215 2101 3219 2105
rect 3391 2101 3395 2105
rect 3567 2101 3571 2105
rect 3743 2101 3747 2105
rect 3895 2101 3899 2105
rect 2391 2091 2392 2095
rect 2392 2091 2395 2095
rect 2927 2091 2931 2095
rect 3479 2091 3483 2095
rect 3815 2091 3816 2095
rect 3816 2091 3819 2095
rect 3959 2091 3963 2095
rect 535 2083 539 2087
rect 919 2083 920 2087
rect 920 2083 923 2087
rect 1455 2083 1459 2087
rect 1739 2083 1740 2087
rect 1740 2083 1743 2087
rect 151 2075 155 2079
rect 303 2075 307 2079
rect 479 2075 483 2079
rect 663 2075 667 2079
rect 847 2075 851 2079
rect 1039 2075 1043 2079
rect 1239 2075 1243 2079
rect 1447 2075 1451 2079
rect 1663 2075 1667 2079
rect 223 2067 227 2071
rect 727 2067 731 2071
rect 1115 2067 1119 2071
rect 1879 2075 1883 2079
rect 3247 2075 3251 2079
rect 2007 2067 2011 2071
rect 2215 2067 2219 2071
rect 111 2056 115 2060
rect 2031 2056 2035 2060
rect 2207 2059 2211 2063
rect 2647 2067 2648 2071
rect 2648 2067 2651 2071
rect 2391 2059 2395 2063
rect 2575 2059 2579 2063
rect 2759 2059 2763 2063
rect 3111 2067 3115 2071
rect 3639 2067 3643 2071
rect 2935 2059 2939 2063
rect 3103 2059 3107 2063
rect 3263 2059 3267 2063
rect 3423 2059 3427 2063
rect 3583 2059 3587 2063
rect 2383 2047 2387 2051
rect 2927 2051 2931 2055
rect 3247 2051 3251 2055
rect 3967 2067 3968 2071
rect 3968 2067 3971 2071
rect 3751 2059 3755 2063
rect 3895 2059 3899 2063
rect 3255 2047 3259 2051
rect 3815 2051 3819 2055
rect 3959 2051 3963 2055
rect 111 2039 115 2043
rect 2031 2039 2035 2043
rect 2071 2040 2075 2044
rect 3991 2040 3995 2044
rect 151 2034 155 2038
rect 303 2034 307 2038
rect 479 2034 483 2038
rect 663 2034 667 2038
rect 847 2034 851 2038
rect 1039 2034 1043 2038
rect 1239 2034 1243 2038
rect 1447 2034 1451 2038
rect 1663 2034 1667 2038
rect 1879 2034 1883 2038
rect 2071 2023 2075 2027
rect 3991 2023 3995 2027
rect 2207 2018 2211 2022
rect 2391 2018 2395 2022
rect 2575 2018 2579 2022
rect 2759 2018 2763 2022
rect 2935 2018 2939 2022
rect 3103 2018 3107 2022
rect 3263 2018 3267 2022
rect 3423 2018 3427 2022
rect 3583 2018 3587 2022
rect 3751 2018 3755 2022
rect 3895 2018 3899 2022
rect 151 1994 155 1998
rect 303 1994 307 1998
rect 487 1994 491 1998
rect 687 1994 691 1998
rect 895 1994 899 1998
rect 1103 1994 1107 1998
rect 1311 1994 1315 1998
rect 1527 1994 1531 1998
rect 1743 1994 1747 1998
rect 1935 1994 1939 1998
rect 111 1989 115 1993
rect 2031 1989 2035 1993
rect 111 1972 115 1976
rect 2031 1972 2035 1976
rect 2279 1974 2283 1978
rect 2463 1974 2467 1978
rect 2639 1974 2643 1978
rect 2815 1974 2819 1978
rect 2983 1974 2987 1978
rect 3151 1974 3155 1978
rect 3311 1974 3315 1978
rect 3463 1974 3467 1978
rect 3615 1974 3619 1978
rect 3767 1974 3771 1978
rect 3895 1974 3899 1978
rect 2071 1969 2075 1973
rect 3991 1969 3995 1973
rect 439 1963 443 1967
rect 479 1963 483 1967
rect 879 1963 883 1967
rect 919 1963 923 1967
rect 1295 1963 1299 1967
rect 1455 1963 1459 1967
rect 1671 1963 1675 1967
rect 151 1953 155 1957
rect 303 1953 307 1957
rect 487 1953 491 1957
rect 687 1953 691 1957
rect 895 1953 899 1957
rect 1103 1953 1107 1957
rect 1311 1953 1315 1957
rect 1527 1953 1531 1957
rect 1743 1953 1747 1957
rect 1935 1953 1939 1957
rect 2071 1952 2075 1956
rect 3991 1952 3995 1956
rect 223 1943 224 1947
rect 224 1943 227 1947
rect 439 1943 443 1947
rect 743 1943 747 1947
rect 879 1943 883 1947
rect 967 1935 971 1939
rect 1295 1943 1299 1947
rect 2007 1943 2008 1947
rect 2008 1943 2011 1947
rect 2447 1943 2451 1947
rect 2591 1943 2595 1947
rect 2647 1943 2651 1947
rect 3295 1943 3299 1947
rect 3447 1943 3451 1947
rect 3639 1943 3643 1947
rect 3967 1943 3971 1947
rect 2279 1933 2283 1937
rect 2463 1933 2467 1937
rect 2639 1933 2643 1937
rect 2815 1933 2819 1937
rect 2983 1933 2987 1937
rect 3151 1933 3155 1937
rect 3311 1933 3315 1937
rect 3463 1933 3467 1937
rect 3615 1933 3619 1937
rect 3767 1933 3771 1937
rect 3895 1933 3899 1937
rect 479 1919 480 1923
rect 480 1919 483 1923
rect 615 1919 616 1923
rect 616 1919 619 1923
rect 151 1911 155 1915
rect 271 1911 275 1915
rect 407 1911 411 1915
rect 543 1911 547 1915
rect 223 1903 227 1907
rect 1551 1919 1555 1923
rect 1671 1919 1675 1923
rect 679 1911 683 1915
rect 823 1911 827 1915
rect 983 1911 987 1915
rect 1159 1911 1163 1915
rect 1343 1911 1347 1915
rect 1543 1911 1547 1915
rect 1751 1911 1755 1915
rect 743 1903 747 1907
rect 967 1903 971 1907
rect 2383 1923 2387 1927
rect 2447 1923 2451 1927
rect 3255 1923 3259 1927
rect 3295 1923 3299 1927
rect 1935 1911 1939 1915
rect 2591 1911 2595 1915
rect 3447 1915 3451 1919
rect 3775 1923 3779 1927
rect 3959 1923 3963 1927
rect 2007 1903 2011 1907
rect 2863 1903 2867 1907
rect 3607 1903 3611 1907
rect 111 1892 115 1896
rect 2031 1892 2035 1896
rect 2407 1895 2411 1899
rect 2655 1895 2659 1899
rect 2887 1895 2891 1899
rect 3103 1895 3107 1899
rect 3311 1895 3315 1899
rect 3511 1895 3515 1899
rect 2431 1883 2435 1887
rect 3167 1887 3171 1891
rect 3967 1903 3968 1907
rect 3968 1903 3971 1907
rect 3711 1895 3715 1899
rect 3895 1895 3899 1899
rect 3775 1887 3779 1891
rect 3887 1883 3891 1887
rect 111 1875 115 1879
rect 2031 1875 2035 1879
rect 2071 1876 2075 1880
rect 3991 1876 3995 1880
rect 151 1870 155 1874
rect 271 1870 275 1874
rect 407 1870 411 1874
rect 543 1870 547 1874
rect 679 1870 683 1874
rect 823 1870 827 1874
rect 983 1870 987 1874
rect 1159 1870 1163 1874
rect 1343 1870 1347 1874
rect 1543 1870 1547 1874
rect 1751 1870 1755 1874
rect 1935 1870 1939 1874
rect 2071 1859 2075 1863
rect 3991 1859 3995 1863
rect 1043 1851 1047 1855
rect 1551 1851 1555 1855
rect 2407 1854 2411 1858
rect 2655 1854 2659 1858
rect 2887 1854 2891 1858
rect 3103 1854 3107 1858
rect 3311 1854 3315 1858
rect 3511 1854 3515 1858
rect 3711 1854 3715 1858
rect 3895 1854 3899 1858
rect 151 1830 155 1834
rect 287 1830 291 1834
rect 447 1830 451 1834
rect 599 1830 603 1834
rect 751 1830 755 1834
rect 919 1830 923 1834
rect 1103 1830 1107 1834
rect 1303 1830 1307 1834
rect 1511 1830 1515 1834
rect 1735 1830 1739 1834
rect 1935 1830 1939 1834
rect 111 1825 115 1829
rect 2031 1825 2035 1829
rect 2111 1822 2115 1826
rect 2383 1822 2387 1826
rect 2647 1822 2651 1826
rect 2887 1822 2891 1826
rect 3095 1822 3099 1826
rect 3287 1822 3291 1826
rect 3455 1822 3459 1826
rect 3615 1822 3619 1826
rect 3767 1822 3771 1826
rect 3895 1822 3899 1826
rect 2071 1817 2075 1821
rect 3991 1817 3995 1821
rect 111 1808 115 1812
rect 2031 1808 2035 1812
rect 427 1799 431 1803
rect 615 1799 619 1803
rect 1043 1799 1047 1803
rect 2063 1799 2067 1803
rect 2071 1800 2075 1804
rect 151 1789 155 1793
rect 287 1789 291 1793
rect 447 1789 451 1793
rect 599 1789 603 1793
rect 751 1789 755 1793
rect 919 1789 923 1793
rect 1103 1789 1107 1793
rect 1303 1789 1307 1793
rect 1511 1789 1515 1793
rect 1735 1789 1739 1793
rect 1935 1789 1939 1793
rect 2183 1791 2187 1795
rect 2579 1791 2583 1795
rect 2863 1791 2867 1795
rect 3079 1791 3083 1795
rect 3359 1791 3363 1795
rect 3563 1791 3567 1795
rect 3607 1791 3611 1795
rect 3903 1799 3907 1803
rect 3991 1800 3995 1804
rect 3967 1791 3971 1795
rect 223 1779 224 1783
rect 224 1779 227 1783
rect 427 1779 431 1783
rect 815 1779 819 1783
rect 1743 1779 1747 1783
rect 2007 1779 2008 1783
rect 2008 1779 2011 1783
rect 2111 1781 2115 1785
rect 2383 1781 2387 1785
rect 2647 1781 2651 1785
rect 2887 1781 2891 1785
rect 3095 1781 3099 1785
rect 3287 1781 3291 1785
rect 3455 1781 3459 1785
rect 3615 1781 3619 1785
rect 3767 1781 3771 1785
rect 3895 1781 3899 1785
rect 2063 1771 2067 1775
rect 2431 1771 2435 1775
rect 1007 1759 1008 1763
rect 1008 1759 1011 1763
rect 1703 1759 1704 1763
rect 1704 1759 1707 1763
rect 2183 1759 2184 1763
rect 2184 1759 2187 1763
rect 207 1751 211 1755
rect 383 1751 387 1755
rect 567 1751 571 1755
rect 751 1751 755 1755
rect 935 1751 939 1755
rect 1111 1751 1115 1755
rect 1279 1751 1283 1755
rect 1455 1751 1459 1755
rect 1631 1751 1635 1755
rect 2111 1751 2115 1755
rect 367 1743 371 1747
rect 815 1743 819 1747
rect 1263 1743 1267 1747
rect 2287 1751 2291 1755
rect 2579 1759 2583 1763
rect 3167 1771 3168 1775
rect 3168 1771 3171 1775
rect 2991 1760 2992 1763
rect 2992 1760 2995 1763
rect 3079 1763 3083 1767
rect 3527 1771 3528 1775
rect 3528 1771 3531 1775
rect 3563 1771 3567 1775
rect 3887 1771 3891 1775
rect 3903 1771 3907 1775
rect 2991 1759 2995 1760
rect 3359 1759 3363 1763
rect 3967 1759 3968 1763
rect 3968 1759 3971 1763
rect 2495 1751 2499 1755
rect 2711 1751 2715 1755
rect 2919 1751 2923 1755
rect 3119 1751 3123 1755
rect 3319 1751 3323 1755
rect 3511 1751 3515 1755
rect 3703 1751 3707 1755
rect 3895 1751 3899 1755
rect 2487 1739 2491 1743
rect 2727 1739 2731 1743
rect 3135 1739 3139 1743
rect 3527 1739 3531 1743
rect 111 1732 115 1736
rect 2031 1732 2035 1736
rect 2071 1732 2075 1736
rect 3991 1732 3995 1736
rect 111 1715 115 1719
rect 2031 1715 2035 1719
rect 207 1710 211 1714
rect 383 1710 387 1714
rect 567 1710 571 1714
rect 751 1710 755 1714
rect 935 1710 939 1714
rect 1111 1710 1115 1714
rect 1279 1710 1283 1714
rect 1455 1710 1459 1714
rect 2071 1715 2075 1719
rect 3991 1715 3995 1719
rect 1631 1710 1635 1714
rect 2111 1710 2115 1714
rect 2287 1710 2291 1714
rect 2495 1710 2499 1714
rect 2711 1710 2715 1714
rect 2919 1710 2923 1714
rect 3119 1710 3123 1714
rect 3319 1710 3323 1714
rect 3511 1710 3515 1714
rect 3703 1710 3707 1714
rect 3895 1710 3899 1714
rect 303 1678 307 1682
rect 535 1678 539 1682
rect 767 1678 771 1682
rect 983 1678 987 1682
rect 1191 1678 1195 1682
rect 1383 1678 1387 1682
rect 1567 1678 1571 1682
rect 1743 1678 1747 1682
rect 1927 1678 1931 1682
rect 111 1673 115 1677
rect 2031 1673 2035 1677
rect 1703 1667 1707 1671
rect 2111 1670 2115 1674
rect 2239 1670 2243 1674
rect 2383 1670 2387 1674
rect 2519 1670 2523 1674
rect 2655 1670 2659 1674
rect 2791 1670 2795 1674
rect 2927 1670 2931 1674
rect 3063 1670 3067 1674
rect 3207 1670 3211 1674
rect 3351 1670 3355 1674
rect 2071 1665 2075 1669
rect 3991 1665 3995 1669
rect 111 1656 115 1660
rect 2031 1656 2035 1660
rect 387 1647 391 1651
rect 751 1647 755 1651
rect 791 1647 795 1651
rect 1007 1647 1011 1651
rect 2071 1648 2075 1652
rect 3991 1648 3995 1652
rect 303 1637 307 1641
rect 535 1637 539 1641
rect 767 1637 771 1641
rect 983 1637 987 1641
rect 1191 1637 1195 1641
rect 1383 1637 1387 1641
rect 1567 1637 1571 1641
rect 1743 1637 1747 1641
rect 1927 1637 1931 1641
rect 2183 1639 2187 1643
rect 2615 1639 2619 1643
rect 2911 1639 2915 1643
rect 2991 1635 2995 1639
rect 3191 1639 3195 1643
rect 367 1627 371 1631
rect 387 1627 391 1631
rect 751 1627 755 1631
rect 791 1611 795 1615
rect 991 1611 995 1615
rect 1999 1627 2000 1631
rect 2000 1627 2003 1631
rect 2111 1629 2115 1633
rect 2239 1629 2243 1633
rect 2383 1629 2387 1633
rect 2519 1629 2523 1633
rect 2655 1629 2659 1633
rect 2791 1629 2795 1633
rect 2927 1629 2931 1633
rect 3063 1629 3067 1633
rect 3207 1629 3211 1633
rect 3351 1629 3355 1633
rect 1431 1619 1435 1623
rect 399 1603 403 1607
rect 575 1603 579 1607
rect 751 1603 755 1607
rect 935 1603 939 1607
rect 1551 1611 1555 1615
rect 2487 1619 2491 1623
rect 2727 1619 2728 1623
rect 2728 1619 2731 1623
rect 2831 1619 2835 1623
rect 2911 1619 2915 1623
rect 3135 1619 3136 1623
rect 3136 1619 3139 1623
rect 3191 1619 3195 1623
rect 3331 1619 3335 1623
rect 559 1595 563 1599
rect 1111 1603 1115 1607
rect 1279 1603 1283 1607
rect 1447 1603 1451 1607
rect 1607 1603 1611 1607
rect 1431 1595 1435 1599
rect 1767 1603 1771 1607
rect 1935 1603 1939 1607
rect 1999 1595 2003 1599
rect 2183 1595 2187 1599
rect 111 1584 115 1588
rect 2031 1584 2035 1588
rect 2167 1587 2171 1591
rect 2287 1587 2291 1591
rect 2407 1587 2411 1591
rect 2615 1595 2619 1599
rect 2919 1595 2923 1599
rect 3331 1595 3332 1599
rect 3332 1595 3335 1599
rect 2527 1587 2531 1591
rect 2647 1587 2651 1591
rect 2767 1587 2771 1591
rect 2887 1587 2891 1591
rect 3007 1587 3011 1591
rect 3127 1587 3131 1591
rect 3255 1587 3259 1591
rect 2535 1575 2539 1579
rect 2747 1579 2751 1583
rect 2831 1579 2835 1583
rect 2991 1579 2995 1583
rect 111 1567 115 1571
rect 2031 1567 2035 1571
rect 2071 1568 2075 1572
rect 3991 1568 3995 1572
rect 399 1562 403 1566
rect 575 1562 579 1566
rect 751 1562 755 1566
rect 935 1562 939 1566
rect 1111 1562 1115 1566
rect 1279 1562 1283 1566
rect 1447 1562 1451 1566
rect 1607 1562 1611 1566
rect 1767 1562 1771 1566
rect 1935 1562 1939 1566
rect 2071 1551 2075 1555
rect 3991 1551 3995 1555
rect 2167 1546 2171 1550
rect 2287 1546 2291 1550
rect 2407 1546 2411 1550
rect 2527 1546 2531 1550
rect 2647 1546 2651 1550
rect 2767 1546 2771 1550
rect 2887 1546 2891 1550
rect 3007 1546 3011 1550
rect 3127 1546 3131 1550
rect 3255 1546 3259 1550
rect 503 1522 507 1526
rect 615 1522 619 1526
rect 735 1522 739 1526
rect 855 1522 859 1526
rect 967 1522 971 1526
rect 1079 1522 1083 1526
rect 1199 1522 1203 1526
rect 1319 1522 1323 1526
rect 1439 1522 1443 1526
rect 1559 1522 1563 1526
rect 111 1517 115 1521
rect 2031 1517 2035 1521
rect 2351 1506 2355 1510
rect 2463 1506 2467 1510
rect 2575 1506 2579 1510
rect 2695 1506 2699 1510
rect 2815 1506 2819 1510
rect 2927 1506 2931 1510
rect 3047 1506 3051 1510
rect 3167 1506 3171 1510
rect 3287 1506 3291 1510
rect 3407 1506 3411 1510
rect 111 1500 115 1504
rect 2031 1500 2035 1504
rect 2071 1501 2075 1505
rect 3991 1501 3995 1505
rect 599 1491 603 1495
rect 719 1491 723 1495
rect 759 1491 763 1495
rect 951 1491 955 1495
rect 991 1491 995 1495
rect 1183 1491 1187 1495
rect 1423 1491 1427 1495
rect 1543 1491 1547 1495
rect 1551 1491 1555 1495
rect 503 1481 507 1485
rect 615 1481 619 1485
rect 735 1481 739 1485
rect 855 1481 859 1485
rect 967 1481 971 1485
rect 1079 1481 1083 1485
rect 1199 1481 1203 1485
rect 1319 1481 1323 1485
rect 1439 1481 1443 1485
rect 1559 1481 1563 1485
rect 2071 1484 2075 1488
rect 3991 1484 3995 1488
rect 559 1471 563 1475
rect 599 1471 603 1475
rect 719 1471 723 1475
rect 919 1471 923 1475
rect 951 1471 955 1475
rect 1271 1471 1272 1475
rect 1272 1471 1275 1475
rect 1423 1471 1427 1475
rect 1543 1471 1547 1475
rect 2447 1475 2451 1479
rect 2639 1471 2643 1475
rect 2887 1475 2891 1479
rect 2919 1475 2923 1479
rect 3151 1475 3155 1479
rect 3271 1475 3275 1479
rect 1183 1463 1187 1467
rect 2351 1465 2355 1469
rect 2463 1465 2467 1469
rect 2575 1465 2579 1469
rect 2695 1465 2699 1469
rect 2815 1465 2819 1469
rect 2927 1465 2931 1469
rect 671 1455 675 1459
rect 759 1447 760 1451
rect 760 1447 763 1451
rect 1407 1455 1411 1459
rect 2535 1455 2536 1459
rect 2536 1455 2539 1459
rect 2747 1459 2751 1463
rect 2767 1455 2768 1459
rect 2768 1455 2771 1459
rect 2991 1463 2995 1467
rect 3047 1465 3051 1469
rect 3167 1465 3171 1469
rect 3287 1465 3291 1469
rect 3407 1465 3411 1469
rect 2999 1455 3000 1459
rect 3000 1455 3003 1459
rect 3151 1455 3155 1459
rect 3271 1455 3275 1459
rect 3379 1455 3383 1459
rect 1167 1447 1171 1451
rect 583 1439 587 1443
rect 687 1439 691 1443
rect 791 1439 795 1443
rect 895 1439 899 1443
rect 999 1439 1003 1443
rect 1103 1439 1107 1443
rect 1207 1439 1211 1443
rect 1311 1439 1315 1443
rect 1415 1439 1419 1443
rect 1519 1439 1523 1443
rect 671 1431 675 1435
rect 855 1431 859 1435
rect 919 1427 923 1431
rect 1271 1431 1275 1435
rect 2639 1431 2640 1435
rect 2640 1431 2643 1435
rect 2887 1431 2891 1435
rect 3207 1431 3211 1435
rect 3379 1431 3380 1435
rect 3380 1431 3383 1435
rect 111 1420 115 1424
rect 2031 1420 2035 1424
rect 2343 1423 2347 1427
rect 2447 1423 2451 1427
rect 2567 1423 2571 1427
rect 2695 1423 2699 1427
rect 2839 1423 2843 1427
rect 2991 1423 2995 1427
rect 3143 1423 3147 1427
rect 3303 1423 3307 1427
rect 2359 1411 2363 1415
rect 2767 1415 2771 1419
rect 3471 1423 3475 1427
rect 3815 1431 3819 1435
rect 3647 1423 3651 1427
rect 3823 1423 3827 1427
rect 2999 1411 3003 1415
rect 3731 1415 3735 1419
rect 3919 1415 3923 1419
rect 111 1403 115 1407
rect 2031 1403 2035 1407
rect 2071 1404 2075 1408
rect 3991 1404 3995 1408
rect 583 1398 587 1402
rect 687 1398 691 1402
rect 791 1398 795 1402
rect 895 1398 899 1402
rect 999 1398 1003 1402
rect 1103 1398 1107 1402
rect 1207 1398 1211 1402
rect 1311 1398 1315 1402
rect 1415 1398 1419 1402
rect 1519 1398 1523 1402
rect 2071 1387 2075 1391
rect 3991 1387 3995 1391
rect 2343 1382 2347 1386
rect 2447 1382 2451 1386
rect 2567 1382 2571 1386
rect 2695 1382 2699 1386
rect 2839 1382 2843 1386
rect 2991 1382 2995 1386
rect 3143 1382 3147 1386
rect 3303 1382 3307 1386
rect 3471 1382 3475 1386
rect 3647 1382 3651 1386
rect 3823 1382 3827 1386
rect 551 1358 555 1362
rect 655 1358 659 1362
rect 759 1358 763 1362
rect 863 1358 867 1362
rect 975 1358 979 1362
rect 1087 1358 1091 1362
rect 1199 1358 1203 1362
rect 1311 1358 1315 1362
rect 1431 1358 1435 1362
rect 1551 1358 1555 1362
rect 111 1353 115 1357
rect 2031 1353 2035 1357
rect 2287 1342 2291 1346
rect 2407 1342 2411 1346
rect 2543 1342 2547 1346
rect 2695 1342 2699 1346
rect 2855 1342 2859 1346
rect 3015 1342 3019 1346
rect 3183 1342 3187 1346
rect 3351 1342 3355 1346
rect 3519 1342 3523 1346
rect 3687 1342 3691 1346
rect 3855 1342 3859 1346
rect 111 1336 115 1340
rect 2031 1336 2035 1340
rect 2071 1337 2075 1341
rect 3991 1337 3995 1341
rect 639 1327 643 1331
rect 1167 1327 1171 1331
rect 1407 1327 1411 1331
rect 551 1317 555 1321
rect 655 1317 659 1321
rect 759 1317 763 1321
rect 863 1317 867 1321
rect 975 1317 979 1321
rect 1087 1317 1091 1321
rect 1199 1317 1203 1321
rect 1311 1317 1315 1321
rect 1431 1317 1435 1321
rect 1551 1317 1555 1321
rect 2071 1320 2075 1324
rect 3991 1320 3995 1324
rect 639 1299 643 1303
rect 343 1283 347 1287
rect 463 1283 467 1287
rect 599 1283 603 1287
rect 743 1283 747 1287
rect 855 1299 859 1303
rect 1255 1307 1259 1311
rect 1607 1307 1611 1311
rect 2391 1311 2395 1315
rect 2527 1311 2531 1315
rect 2839 1311 2843 1315
rect 2927 1311 2931 1315
rect 3167 1311 3171 1315
rect 3207 1311 3211 1315
rect 3927 1311 3931 1315
rect 2287 1301 2291 1305
rect 2407 1301 2411 1305
rect 2543 1301 2547 1305
rect 2695 1301 2699 1305
rect 2855 1301 2859 1305
rect 3015 1301 3019 1305
rect 3183 1301 3187 1305
rect 3351 1301 3355 1305
rect 3519 1301 3523 1305
rect 3687 1301 3691 1305
rect 3855 1301 3859 1305
rect 1127 1291 1131 1295
rect 903 1283 907 1287
rect 1063 1283 1067 1287
rect 447 1275 451 1279
rect 1415 1291 1419 1295
rect 1231 1283 1235 1287
rect 1407 1283 1411 1287
rect 2359 1291 2360 1295
rect 2360 1291 2363 1295
rect 2391 1291 2395 1295
rect 2527 1291 2531 1295
rect 2767 1291 2768 1295
rect 2768 1291 2771 1295
rect 2839 1291 2843 1295
rect 3087 1291 3088 1295
rect 3088 1291 3091 1295
rect 3167 1291 3171 1295
rect 3323 1291 3327 1295
rect 3731 1291 3735 1295
rect 3919 1291 3923 1295
rect 1583 1283 1587 1287
rect 1255 1271 1259 1275
rect 1607 1271 1611 1275
rect 2927 1271 2931 1275
rect 3007 1271 3011 1275
rect 3323 1271 3324 1275
rect 3324 1271 3327 1275
rect 111 1264 115 1268
rect 2031 1264 2035 1268
rect 2127 1263 2131 1267
rect 2295 1263 2299 1267
rect 2479 1263 2483 1267
rect 2679 1263 2683 1267
rect 2879 1263 2883 1267
rect 3071 1263 3075 1267
rect 3247 1263 3251 1267
rect 3415 1263 3419 1267
rect 3583 1263 3587 1267
rect 3927 1271 3931 1275
rect 3751 1263 3755 1267
rect 3895 1263 3899 1267
rect 111 1247 115 1251
rect 2031 1247 2035 1251
rect 2151 1251 2155 1255
rect 2871 1251 2875 1255
rect 3087 1251 3091 1255
rect 3815 1255 3819 1259
rect 3959 1255 3963 1259
rect 343 1242 347 1246
rect 463 1242 467 1246
rect 599 1242 603 1246
rect 743 1242 747 1246
rect 903 1242 907 1246
rect 1063 1242 1067 1246
rect 1231 1242 1235 1246
rect 1407 1242 1411 1246
rect 1583 1242 1587 1246
rect 2071 1244 2075 1248
rect 3991 1244 3995 1248
rect 447 1227 451 1231
rect 991 1227 995 1231
rect 2071 1227 2075 1231
rect 3991 1227 3995 1231
rect 2127 1222 2131 1226
rect 2295 1222 2299 1226
rect 2479 1222 2483 1226
rect 2679 1222 2683 1226
rect 2879 1222 2883 1226
rect 3071 1222 3075 1226
rect 3247 1222 3251 1226
rect 3415 1222 3419 1226
rect 3583 1222 3587 1226
rect 3751 1222 3755 1226
rect 3895 1222 3899 1226
rect 183 1210 187 1214
rect 351 1210 355 1214
rect 535 1210 539 1214
rect 727 1210 731 1214
rect 919 1210 923 1214
rect 1103 1210 1107 1214
rect 1287 1210 1291 1214
rect 1471 1210 1475 1214
rect 1655 1210 1659 1214
rect 1839 1210 1843 1214
rect 111 1205 115 1209
rect 2031 1205 2035 1209
rect 111 1188 115 1192
rect 2031 1188 2035 1192
rect 335 1179 339 1183
rect 1127 1179 1131 1183
rect 1415 1179 1419 1183
rect 2111 1178 2115 1182
rect 2247 1178 2251 1182
rect 2407 1178 2411 1182
rect 2559 1178 2563 1182
rect 2703 1178 2707 1182
rect 2863 1178 2867 1182
rect 3039 1178 3043 1182
rect 3239 1178 3243 1182
rect 3455 1178 3459 1182
rect 3687 1178 3691 1182
rect 3895 1178 3899 1182
rect 183 1169 187 1173
rect 351 1169 355 1173
rect 535 1169 539 1173
rect 727 1169 731 1173
rect 919 1169 923 1173
rect 1103 1169 1107 1173
rect 1287 1169 1291 1173
rect 1471 1169 1475 1173
rect 1655 1169 1659 1173
rect 1839 1169 1843 1173
rect 2071 1173 2075 1177
rect 3991 1173 3995 1177
rect 991 1159 992 1163
rect 992 1159 995 1163
rect 1187 1159 1191 1163
rect 1911 1159 1912 1163
rect 1912 1159 1915 1163
rect 2071 1156 2075 1160
rect 3991 1156 3995 1160
rect 335 1147 339 1151
rect 2231 1147 2235 1151
rect 2391 1147 2395 1151
rect 2663 1147 2667 1151
rect 3007 1147 3011 1151
rect 3967 1147 3971 1151
rect 1083 1139 1087 1143
rect 1211 1139 1215 1143
rect 151 1131 155 1135
rect 303 1131 307 1135
rect 495 1131 499 1135
rect 703 1131 707 1135
rect 911 1131 915 1135
rect 1119 1131 1123 1135
rect 1319 1131 1323 1135
rect 1187 1123 1191 1127
rect 1519 1131 1523 1135
rect 1719 1131 1723 1135
rect 2111 1137 2115 1141
rect 2247 1137 2251 1141
rect 2407 1137 2411 1141
rect 2559 1137 2563 1141
rect 2703 1137 2707 1141
rect 2863 1137 2867 1141
rect 3039 1137 3043 1141
rect 3239 1137 3243 1141
rect 3455 1137 3459 1141
rect 3687 1137 3691 1141
rect 3895 1137 3899 1141
rect 1919 1131 1923 1135
rect 2151 1131 2155 1135
rect 2231 1127 2235 1131
rect 1911 1123 1915 1127
rect 2391 1127 2395 1131
rect 2871 1127 2875 1131
rect 3071 1119 3075 1123
rect 3959 1127 3963 1131
rect 111 1112 115 1116
rect 2031 1112 2035 1116
rect 2663 1111 2667 1115
rect 3759 1111 3763 1115
rect 3967 1111 3968 1115
rect 3968 1111 3971 1115
rect 2111 1103 2115 1107
rect 2303 1103 2307 1107
rect 2511 1103 2515 1107
rect 2703 1103 2707 1107
rect 2895 1103 2899 1107
rect 3087 1103 3091 1107
rect 3287 1103 3291 1107
rect 3495 1103 3499 1107
rect 3703 1103 3707 1107
rect 3895 1103 3899 1107
rect 111 1095 115 1099
rect 2031 1095 2035 1099
rect 151 1090 155 1094
rect 303 1090 307 1094
rect 495 1090 499 1094
rect 703 1090 707 1094
rect 911 1090 915 1094
rect 1119 1090 1123 1094
rect 1319 1090 1323 1094
rect 1519 1090 1523 1094
rect 1719 1090 1723 1094
rect 1919 1090 1923 1094
rect 2103 1091 2107 1095
rect 2879 1095 2883 1099
rect 3071 1095 3075 1099
rect 3959 1095 3963 1099
rect 2071 1084 2075 1088
rect 3991 1084 3995 1088
rect 2071 1067 2075 1071
rect 3991 1067 3995 1071
rect 2111 1062 2115 1066
rect 2303 1062 2307 1066
rect 2511 1062 2515 1066
rect 2703 1062 2707 1066
rect 2895 1062 2899 1066
rect 3087 1062 3091 1066
rect 3287 1062 3291 1066
rect 3495 1062 3499 1066
rect 3703 1062 3707 1066
rect 3895 1062 3899 1066
rect 151 1050 155 1054
rect 279 1050 283 1054
rect 447 1050 451 1054
rect 623 1050 627 1054
rect 799 1050 803 1054
rect 967 1050 971 1054
rect 1127 1050 1131 1054
rect 1279 1050 1283 1054
rect 1423 1050 1427 1054
rect 1559 1050 1563 1054
rect 1695 1050 1699 1054
rect 1823 1050 1827 1054
rect 1935 1050 1939 1054
rect 111 1045 115 1049
rect 2031 1045 2035 1049
rect 111 1028 115 1032
rect 2031 1028 2035 1032
rect 223 1019 227 1023
rect 1083 1019 1087 1023
rect 1211 1019 1215 1023
rect 1407 1019 1411 1023
rect 2319 1014 2323 1018
rect 151 1009 155 1013
rect 279 1009 283 1013
rect 447 1009 451 1013
rect 623 1009 627 1013
rect 799 1009 803 1013
rect 967 1009 971 1013
rect 1127 1009 1131 1013
rect 1279 1009 1283 1013
rect 1423 1009 1427 1013
rect 1559 1009 1563 1013
rect 1695 1009 1699 1013
rect 1823 1009 1827 1013
rect 1935 1009 1939 1013
rect 2487 1014 2491 1018
rect 2663 1014 2667 1018
rect 2847 1014 2851 1018
rect 3039 1014 3043 1018
rect 3247 1014 3251 1018
rect 3463 1014 3467 1018
rect 3687 1014 3691 1018
rect 3895 1014 3899 1018
rect 2071 1009 2075 1013
rect 3991 1009 3995 1013
rect 1043 999 1044 1003
rect 1044 999 1047 1003
rect 1203 999 1204 1003
rect 1204 999 1207 1003
rect 2103 999 2107 1003
rect 2071 992 2075 996
rect 3991 992 3995 996
rect 1407 983 1411 987
rect 223 975 224 979
rect 224 975 227 979
rect 151 967 155 971
rect 287 967 291 971
rect 471 967 475 971
rect 671 967 675 971
rect 871 967 875 971
rect 935 971 939 975
rect 1043 975 1047 979
rect 999 967 1003 971
rect 1203 975 1207 979
rect 1503 975 1507 979
rect 1079 967 1083 971
rect 1287 967 1291 971
rect 1495 967 1499 971
rect 1703 967 1707 971
rect 655 959 659 963
rect 3447 983 3451 987
rect 3759 983 3763 987
rect 3967 983 3971 987
rect 2319 973 2323 977
rect 2487 973 2491 977
rect 2663 973 2667 977
rect 2847 973 2851 977
rect 1911 967 1915 971
rect 663 955 667 959
rect 1983 959 1987 963
rect 2671 963 2675 967
rect 2879 963 2883 967
rect 3039 973 3043 977
rect 3247 973 3251 977
rect 3463 973 3467 977
rect 3687 973 3691 977
rect 3895 973 3899 977
rect 3215 963 3219 967
rect 3447 963 3451 967
rect 3959 963 3963 967
rect 111 948 115 952
rect 2031 948 2035 952
rect 2831 947 2832 951
rect 2832 947 2835 951
rect 3783 947 3784 951
rect 3784 947 3787 951
rect 3967 947 3968 951
rect 3968 947 3971 951
rect 2151 939 2155 943
rect 2287 939 2291 943
rect 2431 939 2435 943
rect 2591 939 2595 943
rect 2759 939 2763 943
rect 2935 939 2939 943
rect 3119 939 3123 943
rect 3311 939 3315 943
rect 3511 939 3515 943
rect 3711 939 3715 943
rect 3895 939 3899 943
rect 111 931 115 935
rect 2031 931 2035 935
rect 151 926 155 930
rect 287 926 291 930
rect 471 926 475 930
rect 671 926 675 930
rect 871 926 875 930
rect 1079 926 1083 930
rect 1287 926 1291 930
rect 1495 926 1499 930
rect 1703 926 1707 930
rect 2271 931 2275 935
rect 2671 931 2675 935
rect 3215 931 3219 935
rect 3959 931 3963 935
rect 1911 926 1915 930
rect 2071 920 2075 924
rect 3991 920 3995 924
rect 1503 907 1507 911
rect 2071 903 2075 907
rect 3991 903 3995 907
rect 2151 898 2155 902
rect 2287 898 2291 902
rect 2431 898 2435 902
rect 2591 898 2595 902
rect 2759 898 2763 902
rect 2935 898 2939 902
rect 3119 898 3123 902
rect 3311 898 3315 902
rect 3511 898 3515 902
rect 3711 898 3715 902
rect 3895 898 3899 902
rect 151 886 155 890
rect 319 886 323 890
rect 519 886 523 890
rect 727 886 731 890
rect 935 886 939 890
rect 1143 886 1147 890
rect 1335 886 1339 890
rect 1527 886 1531 890
rect 1719 886 1723 890
rect 1911 886 1915 890
rect 111 881 115 885
rect 2031 881 2035 885
rect 111 864 115 868
rect 2031 864 2035 868
rect 231 855 235 859
rect 751 855 755 859
rect 2111 854 2115 858
rect 2239 854 2243 858
rect 2407 854 2411 858
rect 2575 854 2579 858
rect 2751 854 2755 858
rect 2935 854 2939 858
rect 3119 854 3123 858
rect 3311 854 3315 858
rect 3511 854 3515 858
rect 3711 854 3715 858
rect 3895 854 3899 858
rect 151 845 155 849
rect 319 845 323 849
rect 519 845 523 849
rect 727 845 731 849
rect 935 845 939 849
rect 1143 845 1147 849
rect 1335 845 1339 849
rect 1527 845 1531 849
rect 1719 845 1723 849
rect 1911 845 1915 849
rect 2071 849 2075 853
rect 3991 849 3995 853
rect 663 835 667 839
rect 231 827 235 831
rect 1983 835 1984 839
rect 1984 835 1987 839
rect 2071 832 2075 836
rect 3991 832 3995 836
rect 2183 823 2187 827
rect 2559 823 2563 827
rect 2735 823 2739 827
rect 2831 823 2835 827
rect 3495 823 3499 827
rect 3695 823 3699 827
rect 3783 823 3787 827
rect 3967 823 3971 827
rect 751 811 755 815
rect 1727 811 1731 815
rect 2011 811 2012 815
rect 2012 811 2015 815
rect 2111 813 2115 817
rect 2239 813 2243 817
rect 2407 813 2411 817
rect 2575 813 2579 817
rect 2751 813 2755 817
rect 2935 813 2939 817
rect 3119 813 3123 817
rect 3311 813 3315 817
rect 3511 813 3515 817
rect 3711 813 3715 817
rect 3895 813 3899 817
rect 263 803 267 807
rect 367 803 371 807
rect 479 803 483 807
rect 591 803 595 807
rect 711 803 715 807
rect 855 803 859 807
rect 1031 803 1035 807
rect 1239 803 1243 807
rect 1471 803 1475 807
rect 1711 803 1715 807
rect 1935 803 1939 807
rect 2271 803 2275 807
rect 2455 803 2459 807
rect 2559 803 2563 807
rect 2735 803 2739 807
rect 351 795 355 799
rect 999 795 1003 799
rect 1927 791 1931 795
rect 2011 791 2015 795
rect 2183 791 2184 795
rect 2184 791 2187 795
rect 2463 791 2464 795
rect 2464 791 2467 795
rect 3271 803 3275 807
rect 3495 803 3499 807
rect 3695 803 3699 807
rect 3959 803 3963 807
rect 111 784 115 788
rect 2031 784 2035 788
rect 2111 783 2115 787
rect 2391 783 2395 787
rect 2679 783 2683 787
rect 2455 775 2459 779
rect 3823 791 3827 795
rect 3967 791 3968 795
rect 3968 791 3971 795
rect 2951 783 2955 787
rect 3199 783 3203 787
rect 3439 783 3443 787
rect 3671 783 3675 787
rect 3895 783 3899 787
rect 3063 775 3067 779
rect 3271 775 3275 779
rect 111 767 115 771
rect 2031 767 2035 771
rect 3919 771 3923 775
rect 263 762 267 766
rect 367 762 371 766
rect 479 762 483 766
rect 591 762 595 766
rect 711 762 715 766
rect 855 762 859 766
rect 1031 762 1035 766
rect 1239 762 1243 766
rect 1471 762 1475 766
rect 1711 762 1715 766
rect 1935 762 1939 766
rect 2071 764 2075 768
rect 3991 764 3995 768
rect 1079 743 1083 747
rect 1727 743 1731 747
rect 2071 747 2075 751
rect 3991 747 3995 751
rect 2111 742 2115 746
rect 2391 742 2395 746
rect 2679 742 2683 746
rect 2951 742 2955 746
rect 3199 742 3203 746
rect 3439 742 3443 746
rect 3671 742 3675 746
rect 3895 742 3899 746
rect 423 726 427 730
rect 527 726 531 730
rect 639 726 643 730
rect 759 726 763 730
rect 879 726 883 730
rect 1007 726 1011 730
rect 1143 726 1147 730
rect 1287 726 1291 730
rect 1447 726 1451 730
rect 1615 726 1619 730
rect 1783 726 1787 730
rect 1935 726 1939 730
rect 111 721 115 725
rect 2031 721 2035 725
rect 111 704 115 708
rect 2031 704 2035 708
rect 2111 702 2115 706
rect 2327 702 2331 706
rect 2551 702 2555 706
rect 2775 702 2779 706
rect 2991 702 2995 706
rect 3207 702 3211 706
rect 3415 702 3419 706
rect 3623 702 3627 706
rect 3831 702 3835 706
rect 511 695 515 699
rect 623 695 627 699
rect 743 695 747 699
rect 863 695 867 699
rect 871 695 875 699
rect 1079 695 1083 699
rect 1891 695 1895 699
rect 2063 695 2067 699
rect 2071 697 2075 701
rect 3991 697 3995 701
rect 423 685 427 689
rect 527 685 531 689
rect 639 685 643 689
rect 759 685 763 689
rect 879 685 883 689
rect 1007 685 1011 689
rect 1143 685 1147 689
rect 1287 685 1291 689
rect 1447 685 1451 689
rect 1615 685 1619 689
rect 1783 685 1787 689
rect 1935 685 1939 689
rect 2071 680 2075 684
rect 351 675 355 679
rect 511 675 515 679
rect 623 675 627 679
rect 743 675 747 679
rect 863 675 867 679
rect 679 663 683 667
rect 1247 667 1251 671
rect 1927 675 1931 679
rect 3991 680 3995 684
rect 1891 667 1895 671
rect 2183 671 2187 675
rect 2463 671 2467 675
rect 3191 671 3195 675
rect 3199 671 3203 675
rect 3547 671 3551 675
rect 3823 671 3827 675
rect 871 655 875 659
rect 2111 661 2115 665
rect 2327 661 2331 665
rect 2551 661 2555 665
rect 2775 661 2779 665
rect 2991 661 2995 665
rect 3207 661 3211 665
rect 3415 661 3419 665
rect 3623 661 3627 665
rect 3831 661 3835 665
rect 591 643 595 647
rect 695 643 699 647
rect 807 643 811 647
rect 919 643 923 647
rect 1031 643 1035 647
rect 1143 643 1147 647
rect 1263 643 1267 647
rect 1383 643 1387 647
rect 1503 643 1507 647
rect 1567 643 1571 647
rect 2063 651 2067 655
rect 1623 643 1627 647
rect 2723 643 2727 647
rect 3063 651 3064 655
rect 3064 651 3067 655
rect 3191 651 3195 655
rect 3695 651 3696 655
rect 3696 651 3699 655
rect 3111 643 3115 647
rect 679 635 683 639
rect 943 631 947 635
rect 1247 635 1251 639
rect 2183 635 2187 639
rect 111 624 115 628
rect 2031 624 2035 628
rect 2127 627 2131 631
rect 2295 627 2299 631
rect 2871 635 2875 639
rect 3199 635 3200 639
rect 3200 635 3203 639
rect 3547 643 3551 647
rect 2455 627 2459 631
rect 2615 627 2619 631
rect 2783 627 2787 631
rect 2951 627 2955 631
rect 3127 627 3131 631
rect 3303 627 3307 631
rect 2519 619 2523 623
rect 2723 619 2727 623
rect 3111 619 3115 623
rect 3815 635 3819 639
rect 3919 639 3923 643
rect 3487 627 3491 631
rect 3679 627 3683 631
rect 3879 627 3883 631
rect 3479 615 3483 619
rect 3695 615 3699 619
rect 3895 615 3899 619
rect 111 607 115 611
rect 2031 607 2035 611
rect 2071 608 2075 612
rect 3991 608 3995 612
rect 591 602 595 606
rect 695 602 699 606
rect 807 602 811 606
rect 919 602 923 606
rect 1031 602 1035 606
rect 1143 602 1147 606
rect 1263 602 1267 606
rect 1383 602 1387 606
rect 1503 602 1507 606
rect 1623 602 1627 606
rect 2071 591 2075 595
rect 3991 591 3995 595
rect 2127 586 2131 590
rect 2295 586 2299 590
rect 2455 586 2459 590
rect 2615 586 2619 590
rect 2783 586 2787 590
rect 2951 586 2955 590
rect 3127 586 3131 590
rect 3303 586 3307 590
rect 3487 586 3491 590
rect 3679 586 3683 590
rect 3879 586 3883 590
rect 663 562 667 566
rect 775 562 779 566
rect 895 562 899 566
rect 1023 562 1027 566
rect 1159 562 1163 566
rect 1303 562 1307 566
rect 1447 562 1451 566
rect 1591 562 1595 566
rect 1735 562 1739 566
rect 1879 562 1883 566
rect 111 557 115 561
rect 2031 557 2035 561
rect 2303 546 2307 550
rect 2447 546 2451 550
rect 2591 546 2595 550
rect 2735 546 2739 550
rect 2879 546 2883 550
rect 3031 546 3035 550
rect 3183 546 3187 550
rect 3335 546 3339 550
rect 3495 546 3499 550
rect 3655 546 3659 550
rect 3823 546 3827 550
rect 111 540 115 544
rect 2031 540 2035 544
rect 2071 541 2075 545
rect 3991 541 3995 545
rect 879 531 883 535
rect 1267 531 1271 535
rect 1327 531 1331 535
rect 1567 531 1571 535
rect 663 521 667 525
rect 775 521 779 525
rect 895 521 899 525
rect 1023 521 1027 525
rect 1159 521 1163 525
rect 1303 521 1307 525
rect 1447 521 1451 525
rect 1591 521 1595 525
rect 1735 521 1739 525
rect 1879 521 1883 525
rect 2071 524 2075 528
rect 3991 524 3995 528
rect 943 511 947 515
rect 879 503 883 507
rect 1267 511 1271 515
rect 1951 511 1952 515
rect 1952 511 1955 515
rect 2431 515 2435 519
rect 2719 515 2723 519
rect 2807 515 2811 519
rect 2871 515 2875 519
rect 3167 515 3171 519
rect 3719 511 3723 515
rect 3815 515 3819 519
rect 2303 505 2307 509
rect 2447 505 2451 509
rect 2591 505 2595 509
rect 2735 505 2739 509
rect 2879 505 2883 509
rect 3031 505 3035 509
rect 3183 505 3187 509
rect 3335 505 3339 509
rect 3495 505 3499 509
rect 3655 505 3659 509
rect 3823 505 3827 509
rect 2519 495 2520 499
rect 2520 495 2523 499
rect 1039 483 1040 487
rect 1040 483 1043 487
rect 1327 483 1328 487
rect 1328 483 1331 487
rect 1599 483 1603 487
rect 1847 483 1848 487
rect 1848 483 1851 487
rect 535 475 539 479
rect 639 475 643 479
rect 743 475 747 479
rect 847 475 851 479
rect 967 475 971 479
rect 1103 475 1107 479
rect 1255 475 1259 479
rect 1415 475 1419 479
rect 1591 475 1595 479
rect 1775 475 1779 479
rect 559 463 563 467
rect 1239 467 1243 471
rect 2431 487 2435 491
rect 2719 495 2723 499
rect 2955 495 2956 499
rect 2956 495 2959 499
rect 3479 495 3483 499
rect 3567 495 3568 499
rect 3568 495 3571 499
rect 3895 495 3896 499
rect 3896 495 3899 499
rect 2599 483 2603 487
rect 1935 475 1939 479
rect 2807 475 2808 479
rect 2808 475 2811 479
rect 2955 475 2959 479
rect 3391 475 3392 479
rect 3392 475 3395 479
rect 3719 475 3720 479
rect 3720 475 3723 479
rect 3839 475 3843 479
rect 1407 463 1411 467
rect 1951 463 1955 467
rect 2511 467 2515 471
rect 2615 467 2619 471
rect 2735 467 2739 471
rect 2863 467 2867 471
rect 3007 467 3011 471
rect 3159 467 3163 471
rect 3319 467 3323 471
rect 3479 467 3483 471
rect 3647 467 3651 471
rect 3823 467 3827 471
rect 111 456 115 460
rect 2031 456 2035 460
rect 2599 459 2603 463
rect 2887 455 2891 459
rect 3587 459 3591 463
rect 3959 459 3963 463
rect 2071 448 2075 452
rect 3991 448 3995 452
rect 111 439 115 443
rect 2031 439 2035 443
rect 535 434 539 438
rect 639 434 643 438
rect 743 434 747 438
rect 847 434 851 438
rect 967 434 971 438
rect 1103 434 1107 438
rect 1255 434 1259 438
rect 1415 434 1419 438
rect 1591 434 1595 438
rect 1775 434 1779 438
rect 1935 434 1939 438
rect 2071 431 2075 435
rect 3991 431 3995 435
rect 2511 426 2515 430
rect 2615 426 2619 430
rect 2735 426 2739 430
rect 2863 426 2867 430
rect 3007 426 3011 430
rect 3159 426 3163 430
rect 3319 426 3323 430
rect 3479 426 3483 430
rect 3647 426 3651 430
rect 3823 426 3827 430
rect 3391 411 3395 415
rect 495 398 499 402
rect 631 398 635 402
rect 767 398 771 402
rect 911 398 915 402
rect 1047 398 1051 402
rect 1183 398 1187 402
rect 1319 398 1323 402
rect 1447 398 1451 402
rect 1575 398 1579 402
rect 1703 398 1707 402
rect 1831 398 1835 402
rect 1935 398 1939 402
rect 3587 399 3591 403
rect 3783 399 3787 403
rect 111 393 115 397
rect 2031 393 2035 397
rect 2591 382 2595 386
rect 2695 382 2699 386
rect 2815 382 2819 386
rect 2959 382 2963 386
rect 3119 382 3123 386
rect 3303 382 3307 386
rect 3503 382 3507 386
rect 3711 382 3715 386
rect 3895 382 3899 386
rect 111 376 115 380
rect 2031 376 2035 380
rect 2071 377 2075 381
rect 3991 377 3995 381
rect 615 367 619 371
rect 751 367 755 371
rect 839 367 843 371
rect 1031 367 1035 371
rect 1039 367 1043 371
rect 1303 367 1307 371
rect 1559 367 1563 371
rect 1687 367 1691 371
rect 1775 367 1779 371
rect 1847 367 1851 371
rect 495 357 499 361
rect 631 357 635 361
rect 767 357 771 361
rect 911 357 915 361
rect 1047 357 1051 361
rect 1183 357 1187 361
rect 1319 357 1323 361
rect 1447 357 1451 361
rect 1575 357 1579 361
rect 1703 357 1707 361
rect 1831 357 1835 361
rect 1935 357 1939 361
rect 2071 360 2075 364
rect 3991 360 3995 364
rect 559 347 563 351
rect 615 347 619 351
rect 751 347 755 351
rect 967 347 971 351
rect 1031 347 1035 351
rect 1407 347 1411 351
rect 1303 339 1307 343
rect 1559 347 1563 351
rect 1687 347 1691 351
rect 2095 347 2099 351
rect 3839 351 3843 355
rect 3967 351 3971 355
rect 2591 341 2595 345
rect 2695 341 2699 345
rect 2815 341 2819 345
rect 2959 341 2963 345
rect 3119 341 3123 345
rect 3303 341 3307 345
rect 3503 341 3507 345
rect 3711 341 3715 345
rect 3895 341 3899 345
rect 447 331 451 335
rect 855 331 859 335
rect 1687 331 1691 335
rect 839 323 840 327
rect 840 323 843 327
rect 1383 323 1384 327
rect 1384 323 1387 327
rect 1775 323 1776 327
rect 1776 323 1779 327
rect 335 315 339 319
rect 463 315 467 319
rect 607 315 611 319
rect 767 315 771 319
rect 943 315 947 319
rect 1127 315 1131 319
rect 1311 315 1315 319
rect 1503 315 1507 319
rect 1703 315 1707 319
rect 1903 315 1907 319
rect 2095 319 2096 323
rect 2096 319 2099 323
rect 2463 319 2467 323
rect 2887 331 2888 335
rect 2888 331 2891 335
rect 3511 331 3515 335
rect 3783 331 3784 335
rect 3784 331 3787 335
rect 3959 331 3963 335
rect 447 307 451 311
rect 967 303 971 307
rect 1687 307 1691 311
rect 2111 311 2115 315
rect 2271 311 2275 315
rect 2455 311 2459 315
rect 1895 303 1899 307
rect 3687 319 3691 323
rect 3967 319 3968 323
rect 3968 319 3971 323
rect 2631 311 2635 315
rect 2807 311 2811 315
rect 2999 311 3003 315
rect 3215 311 3219 315
rect 3439 311 3443 315
rect 3679 311 3683 315
rect 3895 311 3899 315
rect 2759 303 2763 307
rect 2983 303 2987 307
rect 3959 303 3963 307
rect 111 296 115 300
rect 2031 296 2035 300
rect 2071 292 2075 296
rect 3991 292 3995 296
rect 111 279 115 283
rect 2031 279 2035 283
rect 335 274 339 278
rect 463 274 467 278
rect 607 274 611 278
rect 767 274 771 278
rect 943 274 947 278
rect 1127 274 1131 278
rect 1311 274 1315 278
rect 1503 274 1507 278
rect 1703 274 1707 278
rect 1903 274 1907 278
rect 2071 275 2075 279
rect 3991 275 3995 279
rect 2111 270 2115 274
rect 2271 270 2275 274
rect 2455 270 2459 274
rect 2631 270 2635 274
rect 2807 270 2811 274
rect 2999 270 3003 274
rect 3215 270 3219 274
rect 3439 270 3443 274
rect 3679 270 3683 274
rect 3895 270 3899 274
rect 151 234 155 238
rect 279 234 283 238
rect 431 234 435 238
rect 599 234 603 238
rect 783 234 787 238
rect 975 234 979 238
rect 1175 234 1179 238
rect 1375 234 1379 238
rect 1583 234 1587 238
rect 2111 238 2115 242
rect 1799 234 1803 238
rect 2271 238 2275 242
rect 2471 238 2475 242
rect 2687 238 2691 242
rect 2903 238 2907 242
rect 3111 238 3115 242
rect 3319 238 3323 242
rect 3519 238 3523 242
rect 3719 238 3723 242
rect 3895 238 3899 242
rect 111 229 115 233
rect 2031 229 2035 233
rect 2071 233 2075 237
rect 3991 233 3995 237
rect 3303 227 3307 231
rect 3687 227 3691 231
rect 111 212 115 216
rect 2031 212 2035 216
rect 2071 216 2075 220
rect 3991 216 3995 220
rect 231 203 235 207
rect 1159 203 1163 207
rect 1359 203 1363 207
rect 1383 203 1387 207
rect 2255 207 2259 211
rect 2455 207 2459 211
rect 2463 207 2467 211
rect 3303 207 3307 211
rect 3967 207 3971 211
rect 151 193 155 197
rect 279 193 283 197
rect 431 193 435 197
rect 599 193 603 197
rect 783 193 787 197
rect 975 193 979 197
rect 1175 193 1179 197
rect 1375 193 1379 197
rect 1583 193 1587 197
rect 1799 193 1803 197
rect 2111 197 2115 201
rect 2271 197 2275 201
rect 2471 197 2475 201
rect 2687 197 2691 201
rect 2903 197 2907 201
rect 3111 197 3115 201
rect 3319 197 3323 201
rect 3519 197 3523 201
rect 3719 197 3723 201
rect 3895 197 3899 201
rect 855 183 856 187
rect 856 183 859 187
rect 1039 183 1043 187
rect 1159 183 1163 187
rect 1359 183 1363 187
rect 1895 183 1899 187
rect 2175 187 2179 191
rect 2255 187 2259 191
rect 2455 187 2459 191
rect 2759 187 2760 191
rect 2760 187 2763 191
rect 2999 187 3003 191
rect 3783 187 3787 191
rect 3959 187 3963 191
rect 231 155 235 159
rect 3967 147 3968 151
rect 3968 147 3971 151
rect 151 139 155 143
rect 255 139 259 143
rect 359 139 363 143
rect 471 139 475 143
rect 607 139 611 143
rect 743 139 747 143
rect 879 139 883 143
rect 1015 139 1019 143
rect 1151 139 1155 143
rect 1279 139 1283 143
rect 1399 139 1403 143
rect 1519 139 1523 143
rect 1647 139 1651 143
rect 1775 139 1779 143
rect 2111 139 2115 143
rect 2215 139 2219 143
rect 2319 139 2323 143
rect 2423 139 2427 143
rect 2527 139 2531 143
rect 2655 139 2659 143
rect 2775 139 2779 143
rect 2895 139 2899 143
rect 3015 139 3019 143
rect 3135 139 3139 143
rect 3247 139 3251 143
rect 3359 139 3363 143
rect 3471 139 3475 143
rect 3583 139 3587 143
rect 3687 139 3691 143
rect 3791 139 3795 143
rect 3895 139 3899 143
rect 1039 127 1043 131
rect 2175 131 2179 135
rect 2999 131 3003 135
rect 3783 131 3787 135
rect 111 120 115 124
rect 2031 120 2035 124
rect 2071 120 2075 124
rect 3991 120 3995 124
rect 111 103 115 107
rect 2031 103 2035 107
rect 151 98 155 102
rect 255 98 259 102
rect 359 98 363 102
rect 471 98 475 102
rect 607 98 611 102
rect 743 98 747 102
rect 879 98 883 102
rect 1015 98 1019 102
rect 1151 98 1155 102
rect 1279 98 1283 102
rect 1399 98 1403 102
rect 1519 98 1523 102
rect 1647 98 1651 102
rect 2071 103 2075 107
rect 3991 103 3995 107
rect 1775 98 1779 102
rect 2111 98 2115 102
rect 2215 98 2219 102
rect 2319 98 2323 102
rect 2423 98 2427 102
rect 2527 98 2531 102
rect 2655 98 2659 102
rect 2775 98 2779 102
rect 2895 98 2899 102
rect 3015 98 3019 102
rect 3135 98 3139 102
rect 3247 98 3251 102
rect 3359 98 3363 102
rect 3471 98 3475 102
rect 3583 98 3587 102
rect 3687 98 3691 102
rect 3791 98 3795 102
rect 3895 98 3899 102
<< m3 >>
rect 111 4066 115 4067
rect 111 4061 115 4062
rect 327 4066 331 4067
rect 327 4061 331 4062
rect 431 4066 435 4067
rect 431 4061 435 4062
rect 535 4066 539 4067
rect 535 4061 539 4062
rect 639 4066 643 4067
rect 639 4061 643 4062
rect 743 4066 747 4067
rect 743 4061 747 4062
rect 847 4066 851 4067
rect 847 4061 851 4062
rect 951 4066 955 4067
rect 951 4061 955 4062
rect 1055 4066 1059 4067
rect 1055 4061 1059 4062
rect 1159 4066 1163 4067
rect 1159 4061 1163 4062
rect 1263 4066 1267 4067
rect 1263 4061 1267 4062
rect 1367 4066 1371 4067
rect 1367 4061 1371 4062
rect 1471 4066 1475 4067
rect 1471 4061 1475 4062
rect 2031 4066 2035 4067
rect 2031 4061 2035 4062
rect 2071 4066 2075 4067
rect 2071 4061 2075 4062
rect 2263 4066 2267 4067
rect 2263 4061 2267 4062
rect 2367 4066 2371 4067
rect 2367 4061 2371 4062
rect 2471 4066 2475 4067
rect 2471 4061 2475 4062
rect 2575 4066 2579 4067
rect 2575 4061 2579 4062
rect 2679 4066 2683 4067
rect 2679 4061 2683 4062
rect 3991 4066 3995 4067
rect 3991 4061 3995 4062
rect 112 4046 114 4061
rect 328 4051 330 4061
rect 432 4051 434 4061
rect 536 4051 538 4061
rect 640 4051 642 4061
rect 744 4051 746 4061
rect 848 4051 850 4061
rect 952 4051 954 4061
rect 1056 4051 1058 4061
rect 1160 4051 1162 4061
rect 1264 4051 1266 4061
rect 1368 4051 1370 4061
rect 1472 4051 1474 4061
rect 326 4050 332 4051
rect 326 4046 327 4050
rect 331 4046 332 4050
rect 110 4045 116 4046
rect 326 4045 332 4046
rect 430 4050 436 4051
rect 430 4046 431 4050
rect 435 4046 436 4050
rect 430 4045 436 4046
rect 534 4050 540 4051
rect 534 4046 535 4050
rect 539 4046 540 4050
rect 534 4045 540 4046
rect 638 4050 644 4051
rect 638 4046 639 4050
rect 643 4046 644 4050
rect 638 4045 644 4046
rect 742 4050 748 4051
rect 742 4046 743 4050
rect 747 4046 748 4050
rect 742 4045 748 4046
rect 846 4050 852 4051
rect 846 4046 847 4050
rect 851 4046 852 4050
rect 846 4045 852 4046
rect 950 4050 956 4051
rect 950 4046 951 4050
rect 955 4046 956 4050
rect 950 4045 956 4046
rect 1054 4050 1060 4051
rect 1054 4046 1055 4050
rect 1059 4046 1060 4050
rect 1054 4045 1060 4046
rect 1158 4050 1164 4051
rect 1158 4046 1159 4050
rect 1163 4046 1164 4050
rect 1158 4045 1164 4046
rect 1262 4050 1268 4051
rect 1262 4046 1263 4050
rect 1267 4046 1268 4050
rect 1262 4045 1268 4046
rect 1366 4050 1372 4051
rect 1366 4046 1367 4050
rect 1371 4046 1372 4050
rect 1366 4045 1372 4046
rect 1470 4050 1476 4051
rect 1470 4046 1471 4050
rect 1475 4046 1476 4050
rect 2032 4046 2034 4061
rect 2072 4046 2074 4061
rect 2264 4051 2266 4061
rect 2368 4051 2370 4061
rect 2472 4051 2474 4061
rect 2576 4051 2578 4061
rect 2680 4051 2682 4061
rect 2262 4050 2268 4051
rect 2262 4046 2263 4050
rect 2267 4046 2268 4050
rect 1470 4045 1476 4046
rect 2030 4045 2036 4046
rect 110 4041 111 4045
rect 115 4041 116 4045
rect 110 4040 116 4041
rect 2030 4041 2031 4045
rect 2035 4041 2036 4045
rect 2030 4040 2036 4041
rect 2070 4045 2076 4046
rect 2262 4045 2268 4046
rect 2366 4050 2372 4051
rect 2366 4046 2367 4050
rect 2371 4046 2372 4050
rect 2366 4045 2372 4046
rect 2470 4050 2476 4051
rect 2470 4046 2471 4050
rect 2475 4046 2476 4050
rect 2470 4045 2476 4046
rect 2574 4050 2580 4051
rect 2574 4046 2575 4050
rect 2579 4046 2580 4050
rect 2574 4045 2580 4046
rect 2678 4050 2684 4051
rect 2678 4046 2679 4050
rect 2683 4046 2684 4050
rect 3992 4046 3994 4061
rect 2678 4045 2684 4046
rect 3990 4045 3996 4046
rect 2070 4041 2071 4045
rect 2075 4041 2076 4045
rect 2070 4040 2076 4041
rect 3990 4041 3991 4045
rect 3995 4041 3996 4045
rect 3990 4040 3996 4041
rect 110 4028 116 4029
rect 110 4024 111 4028
rect 115 4024 116 4028
rect 110 4023 116 4024
rect 2030 4028 2036 4029
rect 2030 4024 2031 4028
rect 2035 4024 2036 4028
rect 2030 4023 2036 4024
rect 2070 4028 2076 4029
rect 2070 4024 2071 4028
rect 2075 4024 2076 4028
rect 2070 4023 2076 4024
rect 3990 4028 3996 4029
rect 3990 4024 3991 4028
rect 3995 4024 3996 4028
rect 3990 4023 3996 4024
rect 112 3991 114 4023
rect 410 4019 416 4020
rect 410 4015 411 4019
rect 415 4015 416 4019
rect 410 4014 416 4015
rect 518 4019 524 4020
rect 518 4015 519 4019
rect 523 4015 524 4019
rect 518 4014 524 4015
rect 622 4019 628 4020
rect 622 4015 623 4019
rect 627 4015 628 4019
rect 622 4014 628 4015
rect 726 4019 732 4020
rect 726 4015 727 4019
rect 731 4015 732 4019
rect 726 4014 732 4015
rect 830 4019 836 4020
rect 830 4015 831 4019
rect 835 4015 836 4019
rect 830 4014 836 4015
rect 934 4019 940 4020
rect 934 4015 935 4019
rect 939 4015 940 4019
rect 934 4014 940 4015
rect 1038 4019 1044 4020
rect 1038 4015 1039 4019
rect 1043 4015 1044 4019
rect 1038 4014 1044 4015
rect 1246 4019 1252 4020
rect 1246 4015 1247 4019
rect 1251 4018 1252 4019
rect 1251 4016 1258 4018
rect 1251 4015 1252 4016
rect 1246 4014 1252 4015
rect 326 4009 332 4010
rect 326 4005 327 4009
rect 331 4005 332 4009
rect 326 4004 332 4005
rect 328 3991 330 4004
rect 412 4000 414 4014
rect 430 4009 436 4010
rect 430 4005 431 4009
rect 435 4005 436 4009
rect 430 4004 436 4005
rect 410 3999 416 4000
rect 410 3995 411 3999
rect 415 3995 416 3999
rect 410 3994 416 3995
rect 432 3991 434 4004
rect 520 4000 522 4014
rect 534 4009 540 4010
rect 534 4005 535 4009
rect 539 4005 540 4009
rect 534 4004 540 4005
rect 518 3999 524 4000
rect 518 3995 519 3999
rect 523 3995 524 3999
rect 518 3994 524 3995
rect 536 3991 538 4004
rect 624 4000 626 4014
rect 638 4009 644 4010
rect 638 4005 639 4009
rect 643 4005 644 4009
rect 638 4004 644 4005
rect 622 3999 628 4000
rect 622 3995 623 3999
rect 627 3995 628 3999
rect 622 3994 628 3995
rect 640 3991 642 4004
rect 728 4000 730 4014
rect 742 4009 748 4010
rect 742 4005 743 4009
rect 747 4005 748 4009
rect 742 4004 748 4005
rect 726 3999 732 4000
rect 726 3995 727 3999
rect 731 3995 732 3999
rect 726 3994 732 3995
rect 744 3991 746 4004
rect 832 4000 834 4014
rect 846 4009 852 4010
rect 846 4005 847 4009
rect 851 4005 852 4009
rect 846 4004 852 4005
rect 830 3999 836 4000
rect 830 3995 831 3999
rect 835 3995 836 3999
rect 830 3994 836 3995
rect 848 3991 850 4004
rect 936 4000 938 4014
rect 950 4009 956 4010
rect 950 4005 951 4009
rect 955 4005 956 4009
rect 950 4004 956 4005
rect 934 3999 940 4000
rect 934 3995 935 3999
rect 939 3995 940 3999
rect 934 3994 940 3995
rect 952 3991 954 4004
rect 1040 4000 1042 4014
rect 1054 4009 1060 4010
rect 1054 4005 1055 4009
rect 1059 4005 1060 4009
rect 1054 4004 1060 4005
rect 1158 4009 1164 4010
rect 1158 4005 1159 4009
rect 1163 4005 1164 4009
rect 1158 4004 1164 4005
rect 1038 3999 1044 4000
rect 1038 3995 1039 3999
rect 1043 3995 1044 3999
rect 1038 3994 1044 3995
rect 1056 3991 1058 4004
rect 1160 3991 1162 4004
rect 1256 3992 1258 4016
rect 1262 4009 1268 4010
rect 1262 4005 1263 4009
rect 1267 4005 1268 4009
rect 1262 4004 1268 4005
rect 1366 4009 1372 4010
rect 1366 4005 1367 4009
rect 1371 4005 1372 4009
rect 1366 4004 1372 4005
rect 1470 4009 1476 4010
rect 1470 4005 1471 4009
rect 1475 4005 1476 4009
rect 1470 4004 1476 4005
rect 1254 3991 1260 3992
rect 1264 3991 1266 4004
rect 1368 3991 1370 4004
rect 1472 3991 1474 4004
rect 2032 3991 2034 4023
rect 2072 3995 2074 4023
rect 2334 4019 2340 4020
rect 2334 4015 2335 4019
rect 2339 4015 2340 4019
rect 2334 4014 2340 4015
rect 2598 4019 2604 4020
rect 2598 4015 2599 4019
rect 2603 4015 2604 4019
rect 2598 4014 2604 4015
rect 2262 4009 2268 4010
rect 2262 4005 2263 4009
rect 2267 4005 2268 4009
rect 2262 4004 2268 4005
rect 2264 3995 2266 4004
rect 2071 3994 2075 3995
rect 111 3990 115 3991
rect 111 3985 115 3986
rect 175 3990 179 3991
rect 175 3985 179 3986
rect 327 3990 331 3991
rect 327 3985 331 3986
rect 383 3990 387 3991
rect 383 3985 387 3986
rect 431 3990 435 3991
rect 431 3985 435 3986
rect 535 3990 539 3991
rect 535 3985 539 3986
rect 591 3990 595 3991
rect 591 3985 595 3986
rect 639 3990 643 3991
rect 639 3985 643 3986
rect 743 3990 747 3991
rect 743 3985 747 3986
rect 791 3990 795 3991
rect 791 3985 795 3986
rect 847 3990 851 3991
rect 847 3985 851 3986
rect 951 3990 955 3991
rect 951 3985 955 3986
rect 983 3990 987 3991
rect 983 3985 987 3986
rect 1055 3990 1059 3991
rect 1055 3985 1059 3986
rect 1159 3990 1163 3991
rect 1159 3985 1163 3986
rect 1167 3990 1171 3991
rect 1254 3987 1255 3991
rect 1259 3987 1260 3991
rect 1254 3986 1260 3987
rect 1263 3990 1267 3991
rect 1167 3985 1171 3986
rect 1263 3985 1267 3986
rect 1343 3990 1347 3991
rect 1343 3985 1347 3986
rect 1367 3990 1371 3991
rect 1367 3985 1371 3986
rect 1471 3990 1475 3991
rect 1471 3985 1475 3986
rect 1519 3990 1523 3991
rect 1519 3985 1523 3986
rect 1703 3990 1707 3991
rect 1703 3985 1707 3986
rect 2031 3990 2035 3991
rect 2071 3989 2075 3990
rect 2231 3994 2235 3995
rect 2231 3989 2235 3990
rect 2263 3994 2267 3995
rect 2336 3992 2338 4014
rect 2366 4009 2372 4010
rect 2366 4005 2367 4009
rect 2371 4005 2372 4009
rect 2366 4004 2372 4005
rect 2470 4009 2476 4010
rect 2470 4005 2471 4009
rect 2475 4005 2476 4009
rect 2470 4004 2476 4005
rect 2574 4009 2580 4010
rect 2574 4005 2575 4009
rect 2579 4005 2580 4009
rect 2574 4004 2580 4005
rect 2368 3995 2370 4004
rect 2414 3999 2420 4000
rect 2414 3995 2415 3999
rect 2419 3995 2420 3999
rect 2472 3995 2474 4004
rect 2576 3995 2578 4004
rect 2367 3994 2371 3995
rect 2263 3989 2267 3990
rect 2334 3991 2340 3992
rect 2031 3985 2035 3986
rect 112 3957 114 3985
rect 176 3976 178 3985
rect 384 3976 386 3985
rect 592 3976 594 3985
rect 792 3976 794 3985
rect 862 3983 868 3984
rect 862 3979 863 3983
rect 867 3979 868 3983
rect 862 3978 868 3979
rect 174 3975 180 3976
rect 174 3971 175 3975
rect 179 3971 180 3975
rect 174 3970 180 3971
rect 382 3975 388 3976
rect 382 3971 383 3975
rect 387 3971 388 3975
rect 382 3970 388 3971
rect 590 3975 596 3976
rect 590 3971 591 3975
rect 595 3971 596 3975
rect 590 3970 596 3971
rect 790 3975 796 3976
rect 790 3971 791 3975
rect 795 3971 796 3975
rect 790 3970 796 3971
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 110 3951 116 3952
rect 110 3939 116 3940
rect 110 3935 111 3939
rect 115 3935 116 3939
rect 110 3934 116 3935
rect 174 3934 180 3935
rect 112 3919 114 3934
rect 174 3930 175 3934
rect 179 3930 180 3934
rect 174 3929 180 3930
rect 382 3934 388 3935
rect 382 3930 383 3934
rect 387 3930 388 3934
rect 382 3929 388 3930
rect 590 3934 596 3935
rect 590 3930 591 3934
rect 595 3930 596 3934
rect 590 3929 596 3930
rect 790 3934 796 3935
rect 790 3930 791 3934
rect 795 3930 796 3934
rect 790 3929 796 3930
rect 176 3919 178 3929
rect 384 3919 386 3929
rect 592 3919 594 3929
rect 792 3919 794 3929
rect 111 3918 115 3919
rect 111 3913 115 3914
rect 175 3918 179 3919
rect 175 3913 179 3914
rect 359 3918 363 3919
rect 359 3913 363 3914
rect 383 3918 387 3919
rect 383 3913 387 3914
rect 551 3918 555 3919
rect 551 3913 555 3914
rect 591 3918 595 3919
rect 591 3913 595 3914
rect 735 3918 739 3919
rect 735 3913 739 3914
rect 791 3918 795 3919
rect 791 3913 795 3914
rect 112 3898 114 3913
rect 360 3903 362 3913
rect 535 3908 539 3909
rect 535 3903 539 3904
rect 552 3903 554 3913
rect 736 3903 738 3913
rect 864 3909 866 3978
rect 984 3976 986 3985
rect 1075 3980 1079 3981
rect 1168 3976 1170 3985
rect 1286 3983 1292 3984
rect 1286 3978 1287 3983
rect 1291 3978 1292 3983
rect 1344 3976 1346 3985
rect 1503 3980 1507 3981
rect 1520 3976 1522 3985
rect 1704 3976 1706 3985
rect 1774 3983 1780 3984
rect 1774 3978 1775 3983
rect 1779 3978 1780 3983
rect 982 3975 988 3976
rect 1075 3975 1079 3976
rect 1166 3975 1172 3976
rect 1287 3975 1291 3976
rect 1342 3975 1348 3976
rect 1503 3975 1507 3976
rect 1518 3975 1524 3976
rect 982 3971 983 3975
rect 987 3971 988 3975
rect 982 3970 988 3971
rect 1076 3968 1078 3975
rect 1166 3971 1167 3975
rect 1171 3971 1172 3975
rect 1166 3970 1172 3971
rect 1342 3971 1343 3975
rect 1347 3971 1348 3975
rect 1342 3970 1348 3971
rect 1504 3968 1506 3975
rect 1518 3971 1519 3975
rect 1523 3971 1524 3975
rect 1518 3970 1524 3971
rect 1702 3975 1708 3976
rect 1775 3975 1779 3976
rect 1702 3971 1703 3975
rect 1707 3971 1708 3975
rect 1702 3970 1708 3971
rect 1074 3967 1080 3968
rect 1074 3963 1075 3967
rect 1079 3963 1080 3967
rect 1074 3962 1080 3963
rect 1502 3967 1508 3968
rect 1502 3963 1503 3967
rect 1507 3963 1508 3967
rect 1502 3962 1508 3963
rect 1510 3963 1516 3964
rect 1510 3959 1511 3963
rect 1515 3959 1516 3963
rect 1510 3958 1516 3959
rect 982 3934 988 3935
rect 982 3930 983 3934
rect 987 3930 988 3934
rect 982 3929 988 3930
rect 1166 3934 1172 3935
rect 1166 3930 1167 3934
rect 1171 3930 1172 3934
rect 1166 3929 1172 3930
rect 1342 3934 1348 3935
rect 1342 3930 1343 3934
rect 1347 3930 1348 3934
rect 1342 3929 1348 3930
rect 984 3919 986 3929
rect 1168 3919 1170 3929
rect 1344 3919 1346 3929
rect 919 3918 923 3919
rect 919 3913 923 3914
rect 983 3918 987 3919
rect 983 3913 987 3914
rect 1087 3918 1091 3919
rect 1087 3913 1091 3914
rect 1167 3918 1171 3919
rect 1167 3913 1171 3914
rect 1247 3918 1251 3919
rect 1247 3913 1251 3914
rect 1343 3918 1347 3919
rect 1343 3913 1347 3914
rect 1399 3918 1403 3919
rect 1399 3913 1403 3914
rect 863 3908 867 3909
rect 863 3903 867 3904
rect 920 3903 922 3913
rect 1088 3903 1090 3913
rect 1248 3903 1250 3913
rect 1400 3903 1402 3913
rect 358 3902 364 3903
rect 358 3898 359 3902
rect 363 3898 364 3902
rect 110 3897 116 3898
rect 358 3897 364 3898
rect 110 3893 111 3897
rect 115 3893 116 3897
rect 110 3892 116 3893
rect 110 3880 116 3881
rect 110 3876 111 3880
rect 115 3876 116 3880
rect 110 3875 116 3876
rect 112 3847 114 3875
rect 536 3872 538 3903
rect 550 3902 556 3903
rect 550 3898 551 3902
rect 555 3898 556 3902
rect 550 3897 556 3898
rect 734 3902 740 3903
rect 734 3898 735 3902
rect 739 3898 740 3902
rect 734 3897 740 3898
rect 918 3902 924 3903
rect 918 3898 919 3902
rect 923 3898 924 3902
rect 918 3897 924 3898
rect 1086 3902 1092 3903
rect 1086 3898 1087 3902
rect 1091 3898 1092 3902
rect 1086 3897 1092 3898
rect 1246 3902 1252 3903
rect 1246 3898 1247 3902
rect 1251 3898 1252 3902
rect 1246 3897 1252 3898
rect 1398 3902 1404 3903
rect 1398 3898 1399 3902
rect 1403 3898 1404 3902
rect 1398 3897 1404 3898
rect 534 3871 540 3872
rect 534 3867 535 3871
rect 539 3867 540 3871
rect 534 3866 540 3867
rect 358 3861 364 3862
rect 358 3857 359 3861
rect 363 3857 364 3861
rect 358 3856 364 3857
rect 550 3861 556 3862
rect 550 3857 551 3861
rect 555 3857 556 3861
rect 734 3861 740 3862
rect 550 3856 556 3857
rect 718 3859 724 3860
rect 360 3847 362 3856
rect 552 3847 554 3856
rect 718 3855 719 3859
rect 723 3855 724 3859
rect 734 3857 735 3861
rect 739 3857 740 3861
rect 734 3856 740 3857
rect 918 3861 924 3862
rect 918 3857 919 3861
rect 923 3857 924 3861
rect 918 3856 924 3857
rect 1086 3861 1092 3862
rect 1086 3857 1087 3861
rect 1091 3857 1092 3861
rect 1086 3856 1092 3857
rect 1246 3861 1252 3862
rect 1246 3857 1247 3861
rect 1251 3857 1252 3861
rect 1246 3856 1252 3857
rect 1398 3861 1404 3862
rect 1398 3857 1399 3861
rect 1403 3857 1404 3861
rect 1398 3856 1404 3857
rect 718 3854 724 3855
rect 111 3846 115 3847
rect 111 3841 115 3842
rect 359 3846 363 3847
rect 359 3841 363 3842
rect 551 3846 555 3847
rect 551 3841 555 3842
rect 583 3846 587 3847
rect 583 3841 587 3842
rect 112 3813 114 3841
rect 584 3832 586 3841
rect 582 3831 588 3832
rect 582 3827 583 3831
rect 587 3827 588 3831
rect 582 3826 588 3827
rect 720 3824 722 3854
rect 736 3847 738 3856
rect 920 3847 922 3856
rect 1088 3847 1090 3856
rect 1248 3847 1250 3856
rect 1400 3847 1402 3856
rect 1512 3852 1514 3958
rect 2032 3957 2034 3985
rect 2072 3961 2074 3989
rect 2232 3980 2234 3989
rect 2294 3987 2300 3988
rect 2294 3983 2295 3987
rect 2299 3983 2300 3987
rect 2334 3987 2335 3991
rect 2339 3987 2340 3991
rect 2367 3989 2371 3990
rect 2391 3994 2395 3995
rect 2414 3994 2420 3995
rect 2471 3994 2475 3995
rect 2391 3989 2395 3990
rect 2334 3986 2340 3987
rect 2294 3982 2300 3983
rect 2230 3979 2236 3980
rect 2230 3975 2231 3979
rect 2235 3975 2236 3979
rect 2230 3974 2236 3975
rect 2070 3960 2076 3961
rect 2030 3956 2036 3957
rect 2030 3952 2031 3956
rect 2035 3952 2036 3956
rect 2070 3956 2071 3960
rect 2075 3956 2076 3960
rect 2070 3955 2076 3956
rect 2030 3951 2036 3952
rect 2070 3943 2076 3944
rect 2030 3939 2036 3940
rect 2030 3935 2031 3939
rect 2035 3935 2036 3939
rect 2070 3939 2071 3943
rect 2075 3939 2076 3943
rect 2070 3938 2076 3939
rect 2230 3938 2236 3939
rect 1518 3934 1524 3935
rect 1518 3930 1519 3934
rect 1523 3930 1524 3934
rect 1518 3929 1524 3930
rect 1702 3934 1708 3935
rect 2030 3934 2036 3935
rect 1702 3930 1703 3934
rect 1707 3930 1708 3934
rect 1702 3929 1708 3930
rect 1520 3919 1522 3929
rect 1704 3919 1706 3929
rect 2032 3919 2034 3934
rect 2072 3923 2074 3938
rect 2230 3934 2231 3938
rect 2235 3934 2236 3938
rect 2230 3933 2236 3934
rect 2232 3923 2234 3933
rect 2071 3922 2075 3923
rect 1519 3918 1523 3919
rect 1519 3913 1523 3914
rect 1543 3918 1547 3919
rect 1543 3913 1547 3914
rect 1679 3918 1683 3919
rect 1679 3913 1683 3914
rect 1703 3918 1707 3919
rect 1703 3913 1707 3914
rect 1815 3918 1819 3919
rect 1815 3913 1819 3914
rect 1935 3918 1939 3919
rect 1935 3913 1939 3914
rect 2031 3918 2035 3919
rect 2071 3917 2075 3918
rect 2223 3922 2227 3923
rect 2223 3917 2227 3918
rect 2231 3922 2235 3923
rect 2231 3917 2235 3918
rect 2031 3913 2035 3914
rect 1544 3903 1546 3913
rect 1680 3903 1682 3913
rect 1816 3903 1818 3913
rect 1936 3903 1938 3913
rect 1542 3902 1548 3903
rect 1542 3898 1543 3902
rect 1547 3898 1548 3902
rect 1542 3897 1548 3898
rect 1678 3902 1684 3903
rect 1678 3898 1679 3902
rect 1683 3898 1684 3902
rect 1678 3897 1684 3898
rect 1814 3902 1820 3903
rect 1814 3898 1815 3902
rect 1819 3898 1820 3902
rect 1814 3897 1820 3898
rect 1934 3902 1940 3903
rect 1934 3898 1935 3902
rect 1939 3898 1940 3902
rect 2032 3898 2034 3913
rect 2072 3902 2074 3917
rect 2224 3907 2226 3917
rect 2222 3906 2228 3907
rect 2222 3902 2223 3906
rect 2227 3902 2228 3906
rect 2070 3901 2076 3902
rect 2222 3901 2228 3902
rect 1934 3897 1940 3898
rect 2030 3897 2036 3898
rect 2030 3893 2031 3897
rect 2035 3893 2036 3897
rect 2070 3897 2071 3901
rect 2075 3897 2076 3901
rect 2070 3896 2076 3897
rect 2030 3892 2036 3893
rect 2070 3884 2076 3885
rect 2030 3880 2036 3881
rect 2030 3876 2031 3880
rect 2035 3876 2036 3880
rect 2070 3880 2071 3884
rect 2075 3880 2076 3884
rect 2070 3879 2076 3880
rect 2030 3875 2036 3876
rect 1662 3871 1668 3872
rect 1662 3867 1663 3871
rect 1667 3867 1668 3871
rect 1662 3866 1668 3867
rect 1798 3871 1804 3872
rect 1798 3867 1799 3871
rect 1803 3867 1804 3871
rect 1798 3866 1804 3867
rect 1902 3871 1908 3872
rect 1902 3867 1903 3871
rect 1907 3867 1908 3871
rect 1902 3866 1908 3867
rect 2006 3871 2012 3872
rect 2006 3867 2007 3871
rect 2011 3867 2012 3871
rect 2006 3866 2012 3867
rect 1542 3861 1548 3862
rect 1542 3857 1543 3861
rect 1547 3857 1548 3861
rect 1542 3856 1548 3857
rect 1510 3851 1516 3852
rect 1510 3847 1511 3851
rect 1515 3847 1516 3851
rect 1544 3847 1546 3856
rect 1664 3852 1666 3866
rect 1678 3861 1684 3862
rect 1678 3857 1679 3861
rect 1683 3857 1684 3861
rect 1678 3856 1684 3857
rect 1662 3851 1668 3852
rect 1662 3847 1663 3851
rect 1667 3847 1668 3851
rect 1680 3847 1682 3856
rect 1800 3852 1802 3866
rect 1814 3861 1820 3862
rect 1814 3857 1815 3861
rect 1819 3857 1820 3861
rect 1814 3856 1820 3857
rect 1798 3851 1804 3852
rect 1798 3847 1799 3851
rect 1803 3847 1804 3851
rect 1816 3847 1818 3856
rect 1904 3852 1906 3866
rect 1934 3861 1940 3862
rect 1934 3857 1935 3861
rect 1939 3857 1940 3861
rect 1934 3856 1940 3857
rect 1902 3851 1908 3852
rect 1902 3847 1903 3851
rect 1907 3847 1908 3851
rect 1936 3847 1938 3856
rect 735 3846 739 3847
rect 735 3841 739 3842
rect 887 3846 891 3847
rect 887 3841 891 3842
rect 919 3846 923 3847
rect 919 3841 923 3842
rect 1031 3846 1035 3847
rect 1031 3841 1035 3842
rect 1087 3846 1091 3847
rect 1087 3841 1091 3842
rect 1175 3846 1179 3847
rect 1175 3841 1179 3842
rect 1247 3846 1251 3847
rect 1247 3841 1251 3842
rect 1311 3846 1315 3847
rect 1311 3841 1315 3842
rect 1399 3846 1403 3847
rect 1399 3841 1403 3842
rect 1447 3846 1451 3847
rect 1510 3846 1516 3847
rect 1543 3846 1547 3847
rect 1447 3841 1451 3842
rect 1543 3841 1547 3842
rect 1575 3846 1579 3847
rect 1662 3846 1668 3847
rect 1679 3846 1683 3847
rect 1575 3841 1579 3842
rect 1679 3841 1683 3842
rect 1703 3846 1707 3847
rect 1798 3846 1804 3847
rect 1815 3846 1819 3847
rect 1703 3841 1707 3842
rect 1815 3841 1819 3842
rect 1831 3846 1835 3847
rect 1902 3846 1908 3847
rect 1935 3846 1939 3847
rect 1831 3841 1835 3842
rect 1935 3841 1939 3842
rect 736 3832 738 3841
rect 888 3832 890 3841
rect 1032 3832 1034 3841
rect 1102 3839 1108 3840
rect 1102 3835 1103 3839
rect 1107 3835 1108 3839
rect 1102 3834 1108 3835
rect 734 3831 740 3832
rect 734 3827 735 3831
rect 739 3827 740 3831
rect 734 3826 740 3827
rect 886 3831 892 3832
rect 886 3827 887 3831
rect 891 3827 892 3831
rect 886 3826 892 3827
rect 1030 3831 1036 3832
rect 1030 3827 1031 3831
rect 1035 3827 1036 3831
rect 1030 3826 1036 3827
rect 718 3823 724 3824
rect 718 3819 719 3823
rect 723 3819 724 3823
rect 718 3818 724 3819
rect 110 3812 116 3813
rect 110 3808 111 3812
rect 115 3808 116 3812
rect 110 3807 116 3808
rect 110 3795 116 3796
rect 110 3791 111 3795
rect 115 3791 116 3795
rect 110 3790 116 3791
rect 582 3790 588 3791
rect 112 3763 114 3790
rect 582 3786 583 3790
rect 587 3786 588 3790
rect 582 3785 588 3786
rect 734 3790 740 3791
rect 734 3786 735 3790
rect 739 3786 740 3790
rect 734 3785 740 3786
rect 886 3790 892 3791
rect 886 3786 887 3790
rect 891 3786 892 3790
rect 886 3785 892 3786
rect 1030 3790 1036 3791
rect 1030 3786 1031 3790
rect 1035 3786 1036 3790
rect 1030 3785 1036 3786
rect 584 3763 586 3785
rect 736 3763 738 3785
rect 888 3763 890 3785
rect 1032 3763 1034 3785
rect 111 3762 115 3763
rect 111 3757 115 3758
rect 583 3762 587 3763
rect 583 3757 587 3758
rect 599 3762 603 3763
rect 599 3757 603 3758
rect 719 3762 723 3763
rect 719 3757 723 3758
rect 735 3762 739 3763
rect 735 3757 739 3758
rect 847 3762 851 3763
rect 847 3757 851 3758
rect 887 3762 891 3763
rect 887 3757 891 3758
rect 983 3762 987 3763
rect 983 3757 987 3758
rect 1031 3762 1035 3763
rect 1031 3757 1035 3758
rect 112 3742 114 3757
rect 600 3747 602 3757
rect 720 3747 722 3757
rect 848 3747 850 3757
rect 984 3747 986 3757
rect 598 3746 604 3747
rect 598 3742 599 3746
rect 603 3742 604 3746
rect 110 3741 116 3742
rect 598 3741 604 3742
rect 718 3746 724 3747
rect 718 3742 719 3746
rect 723 3742 724 3746
rect 718 3741 724 3742
rect 846 3746 852 3747
rect 846 3742 847 3746
rect 851 3742 852 3746
rect 846 3741 852 3742
rect 982 3746 988 3747
rect 982 3742 983 3746
rect 987 3742 988 3746
rect 982 3741 988 3742
rect 110 3737 111 3741
rect 115 3737 116 3741
rect 110 3736 116 3737
rect 110 3724 116 3725
rect 110 3720 111 3724
rect 115 3720 116 3724
rect 110 3719 116 3720
rect 112 3687 114 3719
rect 1104 3716 1106 3834
rect 1176 3832 1178 3841
rect 1312 3832 1314 3841
rect 1448 3832 1450 3841
rect 1576 3832 1578 3841
rect 1704 3832 1706 3841
rect 1832 3832 1834 3841
rect 1936 3832 1938 3841
rect 2008 3840 2010 3866
rect 2032 3847 2034 3875
rect 2072 3851 2074 3879
rect 2296 3876 2298 3982
rect 2392 3980 2394 3989
rect 2390 3979 2396 3980
rect 2390 3975 2391 3979
rect 2395 3975 2396 3979
rect 2390 3974 2396 3975
rect 2416 3968 2418 3994
rect 2471 3989 2475 3990
rect 2551 3994 2555 3995
rect 2551 3989 2555 3990
rect 2575 3994 2579 3995
rect 2575 3989 2579 3990
rect 2552 3980 2554 3989
rect 2600 3988 2602 4014
rect 2678 4009 2684 4010
rect 2678 4005 2679 4009
rect 2683 4005 2684 4009
rect 2678 4004 2684 4005
rect 2680 3995 2682 4004
rect 3992 3995 3994 4023
rect 2679 3994 2683 3995
rect 2679 3989 2683 3990
rect 2703 3994 2707 3995
rect 2703 3989 2707 3990
rect 2847 3994 2851 3995
rect 2847 3989 2851 3990
rect 2983 3994 2987 3995
rect 2983 3989 2987 3990
rect 3119 3994 3123 3995
rect 3119 3989 3123 3990
rect 3247 3994 3251 3995
rect 3247 3989 3251 3990
rect 3367 3994 3371 3995
rect 3367 3989 3371 3990
rect 3479 3994 3483 3995
rect 3479 3989 3483 3990
rect 3599 3994 3603 3995
rect 3599 3989 3603 3990
rect 3719 3994 3723 3995
rect 3719 3989 3723 3990
rect 3839 3994 3843 3995
rect 3839 3989 3843 3990
rect 3991 3994 3995 3995
rect 3991 3989 3995 3990
rect 2598 3987 2604 3988
rect 2598 3983 2599 3987
rect 2603 3983 2604 3987
rect 2598 3982 2604 3983
rect 2704 3980 2706 3989
rect 2848 3980 2850 3989
rect 2984 3980 2986 3989
rect 3120 3980 3122 3989
rect 3248 3980 3250 3989
rect 3368 3980 3370 3989
rect 3480 3980 3482 3989
rect 3600 3980 3602 3989
rect 3720 3980 3722 3989
rect 3840 3980 3842 3989
rect 3882 3987 3888 3988
rect 3882 3983 3883 3987
rect 3887 3983 3888 3987
rect 3882 3982 3888 3983
rect 2550 3979 2556 3980
rect 2550 3975 2551 3979
rect 2555 3975 2556 3979
rect 2550 3974 2556 3975
rect 2702 3979 2708 3980
rect 2702 3975 2703 3979
rect 2707 3975 2708 3979
rect 2702 3974 2708 3975
rect 2846 3979 2852 3980
rect 2846 3975 2847 3979
rect 2851 3975 2852 3979
rect 2846 3974 2852 3975
rect 2982 3979 2988 3980
rect 2982 3975 2983 3979
rect 2987 3975 2988 3979
rect 2982 3974 2988 3975
rect 3118 3979 3124 3980
rect 3118 3975 3119 3979
rect 3123 3975 3124 3979
rect 3118 3974 3124 3975
rect 3246 3979 3252 3980
rect 3246 3975 3247 3979
rect 3251 3975 3252 3979
rect 3246 3974 3252 3975
rect 3366 3979 3372 3980
rect 3366 3975 3367 3979
rect 3371 3975 3372 3979
rect 3366 3974 3372 3975
rect 3478 3979 3484 3980
rect 3478 3975 3479 3979
rect 3483 3975 3484 3979
rect 3478 3974 3484 3975
rect 3598 3979 3604 3980
rect 3598 3975 3599 3979
rect 3603 3975 3604 3979
rect 3598 3974 3604 3975
rect 3718 3979 3724 3980
rect 3718 3975 3719 3979
rect 3723 3975 3724 3979
rect 3718 3974 3724 3975
rect 3838 3979 3844 3980
rect 3838 3975 3839 3979
rect 3843 3975 3844 3979
rect 3838 3974 3844 3975
rect 2950 3971 2956 3972
rect 2414 3967 2420 3968
rect 2414 3963 2415 3967
rect 2419 3963 2420 3967
rect 2414 3962 2420 3963
rect 2726 3967 2732 3968
rect 2726 3963 2727 3967
rect 2731 3963 2732 3967
rect 2950 3967 2951 3971
rect 2955 3967 2956 3971
rect 2950 3966 2956 3967
rect 2726 3962 2732 3963
rect 2390 3938 2396 3939
rect 2390 3934 2391 3938
rect 2395 3934 2396 3938
rect 2390 3933 2396 3934
rect 2550 3938 2556 3939
rect 2550 3934 2551 3938
rect 2555 3934 2556 3938
rect 2550 3933 2556 3934
rect 2702 3938 2708 3939
rect 2702 3934 2703 3938
rect 2707 3934 2708 3938
rect 2702 3933 2708 3934
rect 2392 3923 2394 3933
rect 2552 3923 2554 3933
rect 2704 3923 2706 3933
rect 2391 3922 2395 3923
rect 2391 3917 2395 3918
rect 2455 3922 2459 3923
rect 2455 3917 2459 3918
rect 2551 3922 2555 3923
rect 2551 3917 2555 3918
rect 2671 3922 2675 3923
rect 2671 3917 2675 3918
rect 2703 3922 2707 3923
rect 2703 3917 2707 3918
rect 2456 3907 2458 3917
rect 2672 3907 2674 3917
rect 2454 3906 2460 3907
rect 2454 3902 2455 3906
rect 2459 3902 2460 3906
rect 2454 3901 2460 3902
rect 2670 3906 2676 3907
rect 2670 3902 2671 3906
rect 2675 3902 2676 3906
rect 2670 3901 2676 3902
rect 2294 3875 2300 3876
rect 2294 3871 2295 3875
rect 2299 3871 2300 3875
rect 2294 3870 2300 3871
rect 2526 3875 2532 3876
rect 2526 3871 2527 3875
rect 2531 3871 2532 3875
rect 2526 3870 2532 3871
rect 2222 3865 2228 3866
rect 2222 3861 2223 3865
rect 2227 3861 2228 3865
rect 2222 3860 2228 3861
rect 2454 3865 2460 3866
rect 2454 3861 2455 3865
rect 2459 3861 2460 3865
rect 2454 3860 2460 3861
rect 2224 3851 2226 3860
rect 2254 3855 2260 3856
rect 2254 3851 2255 3855
rect 2259 3851 2260 3855
rect 2456 3851 2458 3860
rect 2071 3850 2075 3851
rect 2031 3846 2035 3847
rect 2071 3845 2075 3846
rect 2191 3850 2195 3851
rect 2191 3845 2195 3846
rect 2223 3850 2227 3851
rect 2254 3850 2260 3851
rect 2455 3850 2459 3851
rect 2223 3845 2227 3846
rect 2031 3841 2035 3842
rect 2006 3839 2012 3840
rect 2006 3835 2007 3839
rect 2011 3835 2012 3839
rect 2006 3834 2012 3835
rect 1174 3831 1180 3832
rect 1174 3827 1175 3831
rect 1179 3827 1180 3831
rect 1174 3826 1180 3827
rect 1310 3831 1316 3832
rect 1310 3827 1311 3831
rect 1315 3827 1316 3831
rect 1310 3826 1316 3827
rect 1446 3831 1452 3832
rect 1446 3827 1447 3831
rect 1451 3827 1452 3831
rect 1446 3826 1452 3827
rect 1574 3831 1580 3832
rect 1574 3827 1575 3831
rect 1579 3827 1580 3831
rect 1574 3826 1580 3827
rect 1702 3831 1708 3832
rect 1702 3827 1703 3831
rect 1707 3827 1708 3831
rect 1702 3826 1708 3827
rect 1830 3831 1836 3832
rect 1830 3827 1831 3831
rect 1835 3827 1836 3831
rect 1830 3826 1836 3827
rect 1934 3831 1940 3832
rect 1934 3827 1935 3831
rect 1939 3827 1940 3831
rect 1934 3826 1940 3827
rect 1294 3823 1300 3824
rect 1294 3819 1295 3823
rect 1299 3819 1300 3823
rect 1294 3818 1300 3819
rect 1174 3790 1180 3791
rect 1174 3786 1175 3790
rect 1179 3786 1180 3790
rect 1174 3785 1180 3786
rect 1176 3763 1178 3785
rect 1296 3764 1298 3818
rect 2032 3813 2034 3841
rect 2072 3817 2074 3845
rect 2192 3836 2194 3845
rect 2190 3835 2196 3836
rect 2190 3831 2191 3835
rect 2195 3831 2196 3835
rect 2190 3830 2196 3831
rect 2256 3828 2258 3850
rect 2455 3845 2459 3846
rect 2487 3850 2491 3851
rect 2487 3845 2491 3846
rect 2262 3843 2268 3844
rect 2262 3839 2263 3843
rect 2267 3839 2268 3843
rect 2262 3838 2268 3839
rect 2254 3827 2260 3828
rect 2254 3823 2255 3827
rect 2259 3823 2260 3827
rect 2254 3822 2260 3823
rect 2070 3816 2076 3817
rect 2030 3812 2036 3813
rect 2030 3808 2031 3812
rect 2035 3808 2036 3812
rect 2070 3812 2071 3816
rect 2075 3812 2076 3816
rect 2070 3811 2076 3812
rect 2030 3807 2036 3808
rect 2070 3799 2076 3800
rect 2030 3795 2036 3796
rect 2030 3791 2031 3795
rect 2035 3791 2036 3795
rect 2070 3795 2071 3799
rect 2075 3795 2076 3799
rect 2070 3794 2076 3795
rect 2190 3794 2196 3795
rect 1310 3790 1316 3791
rect 1310 3786 1311 3790
rect 1315 3786 1316 3790
rect 1310 3785 1316 3786
rect 1446 3790 1452 3791
rect 1446 3786 1447 3790
rect 1451 3786 1452 3790
rect 1446 3785 1452 3786
rect 1574 3790 1580 3791
rect 1574 3786 1575 3790
rect 1579 3786 1580 3790
rect 1574 3785 1580 3786
rect 1702 3790 1708 3791
rect 1702 3786 1703 3790
rect 1707 3786 1708 3790
rect 1702 3785 1708 3786
rect 1830 3790 1836 3791
rect 1830 3786 1831 3790
rect 1835 3786 1836 3790
rect 1830 3785 1836 3786
rect 1934 3790 1940 3791
rect 2030 3790 2036 3791
rect 1934 3786 1935 3790
rect 1939 3786 1940 3790
rect 1934 3785 1940 3786
rect 1294 3763 1300 3764
rect 1312 3763 1314 3785
rect 1448 3763 1450 3785
rect 1576 3763 1578 3785
rect 1704 3763 1706 3785
rect 1832 3763 1834 3785
rect 1838 3763 1844 3764
rect 1936 3763 1938 3785
rect 2032 3763 2034 3790
rect 2072 3779 2074 3794
rect 2190 3790 2191 3794
rect 2195 3790 2196 3794
rect 2190 3789 2196 3790
rect 2192 3779 2194 3789
rect 2071 3778 2075 3779
rect 2071 3773 2075 3774
rect 2111 3778 2115 3779
rect 2111 3773 2115 3774
rect 2191 3778 2195 3779
rect 2191 3773 2195 3774
rect 1111 3762 1115 3763
rect 1111 3757 1115 3758
rect 1175 3762 1179 3763
rect 1175 3757 1179 3758
rect 1239 3762 1243 3763
rect 1294 3759 1295 3763
rect 1299 3759 1300 3763
rect 1294 3758 1300 3759
rect 1311 3762 1315 3763
rect 1239 3757 1243 3758
rect 1311 3757 1315 3758
rect 1367 3762 1371 3763
rect 1367 3757 1371 3758
rect 1447 3762 1451 3763
rect 1447 3757 1451 3758
rect 1495 3762 1499 3763
rect 1495 3757 1499 3758
rect 1575 3762 1579 3763
rect 1575 3757 1579 3758
rect 1631 3762 1635 3763
rect 1631 3757 1635 3758
rect 1703 3762 1707 3763
rect 1703 3757 1707 3758
rect 1767 3762 1771 3763
rect 1767 3757 1771 3758
rect 1831 3762 1835 3763
rect 1838 3759 1839 3763
rect 1843 3759 1844 3763
rect 1838 3758 1844 3759
rect 1935 3762 1939 3763
rect 1831 3757 1835 3758
rect 1112 3747 1114 3757
rect 1240 3747 1242 3757
rect 1368 3747 1370 3757
rect 1496 3747 1498 3757
rect 1632 3747 1634 3757
rect 1768 3747 1770 3757
rect 1110 3746 1116 3747
rect 1110 3742 1111 3746
rect 1115 3742 1116 3746
rect 1110 3741 1116 3742
rect 1238 3746 1244 3747
rect 1238 3742 1239 3746
rect 1243 3742 1244 3746
rect 1238 3741 1244 3742
rect 1366 3746 1372 3747
rect 1366 3742 1367 3746
rect 1371 3742 1372 3746
rect 1366 3741 1372 3742
rect 1494 3746 1500 3747
rect 1494 3742 1495 3746
rect 1499 3742 1500 3746
rect 1494 3741 1500 3742
rect 1630 3746 1636 3747
rect 1630 3742 1631 3746
rect 1635 3742 1636 3746
rect 1630 3741 1636 3742
rect 1766 3746 1772 3747
rect 1766 3742 1767 3746
rect 1771 3742 1772 3746
rect 1766 3741 1772 3742
rect 702 3715 708 3716
rect 702 3711 703 3715
rect 707 3711 708 3715
rect 702 3710 708 3711
rect 966 3715 972 3716
rect 966 3711 967 3715
rect 971 3711 972 3715
rect 966 3710 972 3711
rect 1102 3715 1108 3716
rect 1102 3711 1103 3715
rect 1107 3711 1108 3715
rect 1102 3710 1108 3711
rect 1350 3715 1356 3716
rect 1350 3711 1351 3715
rect 1355 3711 1356 3715
rect 1350 3710 1356 3711
rect 598 3705 604 3706
rect 598 3701 599 3705
rect 603 3701 604 3705
rect 598 3700 604 3701
rect 600 3687 602 3700
rect 704 3688 706 3710
rect 718 3705 724 3706
rect 718 3701 719 3705
rect 723 3701 724 3705
rect 718 3700 724 3701
rect 846 3705 852 3706
rect 846 3701 847 3705
rect 851 3701 852 3705
rect 846 3700 852 3701
rect 702 3687 708 3688
rect 720 3687 722 3700
rect 782 3695 788 3696
rect 782 3691 783 3695
rect 787 3691 788 3695
rect 782 3690 788 3691
rect 111 3686 115 3687
rect 111 3681 115 3682
rect 471 3686 475 3687
rect 471 3681 475 3682
rect 599 3686 603 3687
rect 599 3681 603 3682
rect 615 3686 619 3687
rect 702 3683 703 3687
rect 707 3683 708 3687
rect 702 3682 708 3683
rect 719 3686 723 3687
rect 615 3681 619 3682
rect 719 3681 723 3682
rect 759 3686 763 3687
rect 759 3681 763 3682
rect 112 3653 114 3681
rect 472 3672 474 3681
rect 616 3672 618 3681
rect 686 3679 692 3680
rect 686 3675 687 3679
rect 691 3675 692 3679
rect 686 3674 692 3675
rect 470 3671 476 3672
rect 470 3667 471 3671
rect 475 3667 476 3671
rect 614 3671 620 3672
rect 470 3666 476 3667
rect 599 3668 603 3669
rect 614 3667 615 3671
rect 619 3667 620 3671
rect 614 3666 620 3667
rect 598 3663 604 3664
rect 598 3659 599 3663
rect 603 3659 604 3663
rect 598 3658 604 3659
rect 110 3652 116 3653
rect 110 3648 111 3652
rect 115 3648 116 3652
rect 110 3647 116 3648
rect 110 3635 116 3636
rect 110 3631 111 3635
rect 115 3631 116 3635
rect 110 3630 116 3631
rect 470 3630 476 3631
rect 112 3615 114 3630
rect 470 3626 471 3630
rect 475 3626 476 3630
rect 470 3625 476 3626
rect 614 3630 620 3631
rect 614 3626 615 3630
rect 619 3626 620 3630
rect 614 3625 620 3626
rect 472 3615 474 3625
rect 616 3615 618 3625
rect 111 3614 115 3615
rect 111 3609 115 3610
rect 247 3614 251 3615
rect 247 3609 251 3610
rect 375 3614 379 3615
rect 375 3609 379 3610
rect 471 3614 475 3615
rect 471 3609 475 3610
rect 519 3614 523 3615
rect 519 3609 523 3610
rect 615 3614 619 3615
rect 615 3609 619 3610
rect 679 3614 683 3615
rect 679 3609 683 3610
rect 112 3594 114 3609
rect 248 3599 250 3609
rect 376 3599 378 3609
rect 520 3599 522 3609
rect 680 3599 682 3609
rect 246 3598 252 3599
rect 246 3594 247 3598
rect 251 3594 252 3598
rect 110 3593 116 3594
rect 246 3593 252 3594
rect 374 3598 380 3599
rect 374 3594 375 3598
rect 379 3594 380 3598
rect 374 3593 380 3594
rect 518 3598 524 3599
rect 518 3594 519 3598
rect 523 3594 524 3598
rect 518 3593 524 3594
rect 678 3598 684 3599
rect 678 3594 679 3598
rect 683 3594 684 3598
rect 678 3593 684 3594
rect 110 3589 111 3593
rect 115 3589 116 3593
rect 110 3588 116 3589
rect 110 3576 116 3577
rect 110 3572 111 3576
rect 115 3572 116 3576
rect 110 3571 116 3572
rect 112 3531 114 3571
rect 688 3568 690 3674
rect 760 3672 762 3681
rect 758 3671 764 3672
rect 758 3667 759 3671
rect 763 3667 764 3671
rect 758 3666 764 3667
rect 784 3660 786 3690
rect 848 3687 850 3700
rect 968 3696 970 3710
rect 982 3705 988 3706
rect 982 3701 983 3705
rect 987 3701 988 3705
rect 982 3700 988 3701
rect 1110 3705 1116 3706
rect 1110 3701 1111 3705
rect 1115 3701 1116 3705
rect 1110 3700 1116 3701
rect 1238 3705 1244 3706
rect 1238 3701 1239 3705
rect 1243 3701 1244 3705
rect 1238 3700 1244 3701
rect 966 3695 972 3696
rect 966 3691 967 3695
rect 971 3691 972 3695
rect 966 3690 972 3691
rect 984 3687 986 3700
rect 1112 3687 1114 3700
rect 1240 3687 1242 3700
rect 1352 3688 1354 3710
rect 1366 3705 1372 3706
rect 1366 3701 1367 3705
rect 1371 3701 1372 3705
rect 1366 3700 1372 3701
rect 1494 3705 1500 3706
rect 1494 3701 1495 3705
rect 1499 3701 1500 3705
rect 1494 3700 1500 3701
rect 1630 3705 1636 3706
rect 1630 3701 1631 3705
rect 1635 3701 1636 3705
rect 1630 3700 1636 3701
rect 1766 3705 1772 3706
rect 1766 3701 1767 3705
rect 1771 3701 1772 3705
rect 1766 3700 1772 3701
rect 1350 3687 1356 3688
rect 1368 3687 1370 3700
rect 1496 3687 1498 3700
rect 1632 3687 1634 3700
rect 1768 3687 1770 3700
rect 1840 3696 1842 3758
rect 1935 3757 1939 3758
rect 2031 3762 2035 3763
rect 2072 3758 2074 3773
rect 2112 3763 2114 3773
rect 2110 3762 2116 3763
rect 2110 3758 2111 3762
rect 2115 3758 2116 3762
rect 2031 3757 2035 3758
rect 2070 3757 2076 3758
rect 2110 3757 2116 3758
rect 2032 3742 2034 3757
rect 2070 3753 2071 3757
rect 2075 3753 2076 3757
rect 2070 3752 2076 3753
rect 2030 3741 2036 3742
rect 2030 3737 2031 3741
rect 2035 3737 2036 3741
rect 2030 3736 2036 3737
rect 2070 3740 2076 3741
rect 2070 3736 2071 3740
rect 2075 3736 2076 3740
rect 2070 3735 2076 3736
rect 2030 3724 2036 3725
rect 2030 3720 2031 3724
rect 2035 3720 2036 3724
rect 2030 3719 2036 3720
rect 1838 3695 1844 3696
rect 1838 3691 1839 3695
rect 1843 3691 1844 3695
rect 1838 3690 1844 3691
rect 2032 3687 2034 3719
rect 2072 3695 2074 3735
rect 2264 3732 2266 3838
rect 2488 3836 2490 3845
rect 2528 3844 2530 3870
rect 2670 3865 2676 3866
rect 2670 3861 2671 3865
rect 2675 3861 2676 3865
rect 2670 3860 2676 3861
rect 2672 3851 2674 3860
rect 2728 3856 2730 3962
rect 2846 3938 2852 3939
rect 2846 3934 2847 3938
rect 2851 3934 2852 3938
rect 2846 3933 2852 3934
rect 2848 3923 2850 3933
rect 2847 3922 2851 3923
rect 2847 3917 2851 3918
rect 2879 3922 2883 3923
rect 2879 3917 2883 3918
rect 2880 3907 2882 3917
rect 2878 3906 2884 3907
rect 2878 3902 2879 3906
rect 2883 3902 2884 3906
rect 2878 3901 2884 3902
rect 2878 3865 2884 3866
rect 2878 3861 2879 3865
rect 2883 3861 2884 3865
rect 2878 3860 2884 3861
rect 2726 3855 2732 3856
rect 2726 3851 2727 3855
rect 2731 3851 2732 3855
rect 2880 3851 2882 3860
rect 2952 3856 2954 3966
rect 2982 3938 2988 3939
rect 2982 3934 2983 3938
rect 2987 3934 2988 3938
rect 2982 3933 2988 3934
rect 3118 3938 3124 3939
rect 3118 3934 3119 3938
rect 3123 3934 3124 3938
rect 3118 3933 3124 3934
rect 3246 3938 3252 3939
rect 3246 3934 3247 3938
rect 3251 3934 3252 3938
rect 3246 3933 3252 3934
rect 3366 3938 3372 3939
rect 3366 3934 3367 3938
rect 3371 3934 3372 3938
rect 3366 3933 3372 3934
rect 3478 3938 3484 3939
rect 3478 3934 3479 3938
rect 3483 3934 3484 3938
rect 3478 3933 3484 3934
rect 3598 3938 3604 3939
rect 3598 3934 3599 3938
rect 3603 3934 3604 3938
rect 3598 3933 3604 3934
rect 3718 3938 3724 3939
rect 3718 3934 3719 3938
rect 3723 3934 3724 3938
rect 3718 3933 3724 3934
rect 3838 3938 3844 3939
rect 3838 3934 3839 3938
rect 3843 3934 3844 3938
rect 3838 3933 3844 3934
rect 2984 3923 2986 3933
rect 3120 3923 3122 3933
rect 3248 3923 3250 3933
rect 3368 3923 3370 3933
rect 3480 3923 3482 3933
rect 3600 3923 3602 3933
rect 3720 3923 3722 3933
rect 3840 3923 3842 3933
rect 2983 3922 2987 3923
rect 2983 3917 2987 3918
rect 3071 3922 3075 3923
rect 3071 3917 3075 3918
rect 3119 3922 3123 3923
rect 3119 3917 3123 3918
rect 3247 3922 3251 3923
rect 3247 3917 3251 3918
rect 3367 3922 3371 3923
rect 3367 3917 3371 3918
rect 3415 3922 3419 3923
rect 3415 3917 3419 3918
rect 3479 3922 3483 3923
rect 3479 3917 3483 3918
rect 3583 3922 3587 3923
rect 3583 3917 3587 3918
rect 3599 3922 3603 3923
rect 3599 3917 3603 3918
rect 3719 3922 3723 3923
rect 3719 3917 3723 3918
rect 3751 3922 3755 3923
rect 3751 3917 3755 3918
rect 3839 3922 3843 3923
rect 3839 3917 3843 3918
rect 3072 3907 3074 3917
rect 3248 3907 3250 3917
rect 3416 3907 3418 3917
rect 3584 3907 3586 3917
rect 3752 3907 3754 3917
rect 3070 3906 3076 3907
rect 3070 3902 3071 3906
rect 3075 3902 3076 3906
rect 3070 3901 3076 3902
rect 3246 3906 3252 3907
rect 3246 3902 3247 3906
rect 3251 3902 3252 3906
rect 3246 3901 3252 3902
rect 3414 3906 3420 3907
rect 3414 3902 3415 3906
rect 3419 3902 3420 3906
rect 3414 3901 3420 3902
rect 3582 3906 3588 3907
rect 3582 3902 3583 3906
rect 3587 3902 3588 3906
rect 3582 3901 3588 3902
rect 3750 3906 3756 3907
rect 3750 3902 3751 3906
rect 3755 3902 3756 3906
rect 3750 3901 3756 3902
rect 3884 3876 3886 3982
rect 3992 3961 3994 3989
rect 3990 3960 3996 3961
rect 3990 3956 3991 3960
rect 3995 3956 3996 3960
rect 3990 3955 3996 3956
rect 3990 3943 3996 3944
rect 3990 3939 3991 3943
rect 3995 3939 3996 3943
rect 3990 3938 3996 3939
rect 3992 3923 3994 3938
rect 3991 3922 3995 3923
rect 3991 3917 3995 3918
rect 3992 3902 3994 3917
rect 3990 3901 3996 3902
rect 3990 3897 3991 3901
rect 3995 3897 3996 3901
rect 3990 3896 3996 3897
rect 3990 3884 3996 3885
rect 3990 3880 3991 3884
rect 3995 3880 3996 3884
rect 3990 3879 3996 3880
rect 3054 3875 3060 3876
rect 3054 3871 3055 3875
rect 3059 3871 3060 3875
rect 3054 3870 3060 3871
rect 3734 3875 3740 3876
rect 3734 3871 3735 3875
rect 3739 3871 3740 3875
rect 3734 3870 3740 3871
rect 3882 3875 3888 3876
rect 3882 3871 3883 3875
rect 3887 3871 3888 3875
rect 3882 3870 3888 3871
rect 3056 3861 3058 3870
rect 3070 3865 3076 3866
rect 3070 3861 3071 3865
rect 3075 3861 3076 3865
rect 3055 3860 3059 3861
rect 3070 3860 3076 3861
rect 3246 3865 3252 3866
rect 3246 3861 3247 3865
rect 3251 3861 3252 3865
rect 3246 3860 3252 3861
rect 3414 3865 3420 3866
rect 3414 3861 3415 3865
rect 3419 3861 3420 3865
rect 3582 3865 3588 3866
rect 3582 3861 3583 3865
rect 3587 3861 3588 3865
rect 3414 3860 3420 3861
rect 3487 3860 3491 3861
rect 3582 3860 3588 3861
rect 2950 3855 2956 3856
rect 3055 3855 3059 3856
rect 2950 3851 2951 3855
rect 2955 3851 2956 3855
rect 3072 3851 3074 3860
rect 3248 3851 3250 3860
rect 3416 3851 3418 3860
rect 3486 3855 3492 3856
rect 3486 3851 3487 3855
rect 3491 3851 3492 3855
rect 2671 3850 2675 3851
rect 2726 3850 2732 3851
rect 2759 3850 2763 3851
rect 2671 3845 2675 3846
rect 2759 3845 2763 3846
rect 2879 3850 2883 3851
rect 2950 3850 2956 3851
rect 2999 3850 3003 3851
rect 2879 3845 2883 3846
rect 2999 3845 3003 3846
rect 3071 3850 3075 3851
rect 3071 3845 3075 3846
rect 3215 3850 3219 3851
rect 3215 3845 3219 3846
rect 3247 3850 3251 3851
rect 3247 3845 3251 3846
rect 3407 3850 3411 3851
rect 3407 3845 3411 3846
rect 3415 3850 3419 3851
rect 3486 3850 3492 3851
rect 3510 3855 3516 3856
rect 3510 3851 3511 3855
rect 3515 3851 3516 3855
rect 3584 3851 3586 3860
rect 3736 3856 3738 3870
rect 3750 3865 3756 3866
rect 3750 3861 3751 3865
rect 3755 3861 3756 3865
rect 3750 3860 3756 3861
rect 3734 3855 3740 3856
rect 3734 3851 3735 3855
rect 3739 3851 3740 3855
rect 3752 3851 3754 3860
rect 3992 3851 3994 3879
rect 3510 3850 3516 3851
rect 3583 3850 3587 3851
rect 3734 3850 3740 3851
rect 3751 3850 3755 3851
rect 3415 3845 3419 3846
rect 2526 3843 2532 3844
rect 2526 3839 2527 3843
rect 2531 3839 2532 3843
rect 2526 3838 2532 3839
rect 2760 3836 2762 3845
rect 3000 3836 3002 3845
rect 3216 3836 3218 3845
rect 3408 3836 3410 3845
rect 2486 3835 2492 3836
rect 2486 3831 2487 3835
rect 2491 3831 2492 3835
rect 2486 3830 2492 3831
rect 2758 3835 2764 3836
rect 2758 3831 2759 3835
rect 2763 3831 2764 3835
rect 2758 3830 2764 3831
rect 2998 3835 3004 3836
rect 2998 3831 2999 3835
rect 3003 3831 3004 3835
rect 2998 3830 3004 3831
rect 3214 3835 3220 3836
rect 3214 3831 3215 3835
rect 3219 3831 3220 3835
rect 3214 3830 3220 3831
rect 3406 3835 3412 3836
rect 3406 3831 3407 3835
rect 3411 3831 3412 3835
rect 3406 3830 3412 3831
rect 3512 3828 3514 3850
rect 3583 3845 3587 3846
rect 3751 3845 3755 3846
rect 3895 3850 3899 3851
rect 3895 3845 3899 3846
rect 3991 3850 3995 3851
rect 3991 3845 3995 3846
rect 3584 3836 3586 3845
rect 3646 3843 3652 3844
rect 3646 3839 3647 3843
rect 3651 3839 3652 3843
rect 3646 3838 3652 3839
rect 3582 3835 3588 3836
rect 3582 3831 3583 3835
rect 3587 3831 3588 3835
rect 3582 3830 3588 3831
rect 2630 3827 2636 3828
rect 2630 3823 2631 3827
rect 2635 3823 2636 3827
rect 2630 3822 2636 3823
rect 3390 3827 3396 3828
rect 3390 3823 3391 3827
rect 3395 3823 3396 3827
rect 3390 3822 3396 3823
rect 3510 3827 3516 3828
rect 3510 3823 3511 3827
rect 3515 3823 3516 3827
rect 3510 3822 3516 3823
rect 2486 3794 2492 3795
rect 2486 3790 2487 3794
rect 2491 3790 2492 3794
rect 2486 3789 2492 3790
rect 2488 3779 2490 3789
rect 2335 3778 2339 3779
rect 2335 3773 2339 3774
rect 2487 3778 2491 3779
rect 2487 3773 2491 3774
rect 2559 3778 2563 3779
rect 2559 3773 2563 3774
rect 2336 3763 2338 3773
rect 2560 3763 2562 3773
rect 2334 3762 2340 3763
rect 2334 3758 2335 3762
rect 2339 3758 2340 3762
rect 2334 3757 2340 3758
rect 2558 3762 2564 3763
rect 2558 3758 2559 3762
rect 2563 3758 2564 3762
rect 2558 3757 2564 3758
rect 2262 3731 2268 3732
rect 2262 3727 2263 3731
rect 2267 3727 2268 3731
rect 2262 3726 2268 3727
rect 2110 3721 2116 3722
rect 2110 3717 2111 3721
rect 2115 3717 2116 3721
rect 2110 3716 2116 3717
rect 2334 3721 2340 3722
rect 2334 3717 2335 3721
rect 2339 3717 2340 3721
rect 2334 3716 2340 3717
rect 2558 3721 2564 3722
rect 2558 3717 2559 3721
rect 2563 3717 2564 3721
rect 2558 3716 2564 3717
rect 2112 3695 2114 3716
rect 2336 3695 2338 3716
rect 2560 3695 2562 3716
rect 2632 3712 2634 3822
rect 2758 3794 2764 3795
rect 2758 3790 2759 3794
rect 2763 3790 2764 3794
rect 2758 3789 2764 3790
rect 2998 3794 3004 3795
rect 2998 3790 2999 3794
rect 3003 3790 3004 3794
rect 2998 3789 3004 3790
rect 3214 3794 3220 3795
rect 3214 3790 3215 3794
rect 3219 3790 3220 3794
rect 3214 3789 3220 3790
rect 2760 3779 2762 3789
rect 3000 3779 3002 3789
rect 3216 3779 3218 3789
rect 3392 3780 3394 3822
rect 3406 3794 3412 3795
rect 3406 3790 3407 3794
rect 3411 3790 3412 3794
rect 3406 3789 3412 3790
rect 3582 3794 3588 3795
rect 3582 3790 3583 3794
rect 3587 3790 3588 3794
rect 3582 3789 3588 3790
rect 3390 3779 3396 3780
rect 3408 3779 3410 3789
rect 3550 3779 3556 3780
rect 3584 3779 3586 3789
rect 2759 3778 2763 3779
rect 2759 3773 2763 3774
rect 2775 3778 2779 3779
rect 2775 3773 2779 3774
rect 2975 3778 2979 3779
rect 2975 3773 2979 3774
rect 2999 3778 3003 3779
rect 2999 3773 3003 3774
rect 3159 3778 3163 3779
rect 3159 3773 3163 3774
rect 3215 3778 3219 3779
rect 3215 3773 3219 3774
rect 3327 3778 3331 3779
rect 3390 3775 3391 3779
rect 3395 3775 3396 3779
rect 3390 3774 3396 3775
rect 3407 3778 3411 3779
rect 3327 3773 3331 3774
rect 3407 3773 3411 3774
rect 3479 3778 3483 3779
rect 3550 3775 3551 3779
rect 3555 3775 3556 3779
rect 3550 3774 3556 3775
rect 3583 3778 3587 3779
rect 3479 3773 3483 3774
rect 2776 3763 2778 3773
rect 2976 3763 2978 3773
rect 3160 3763 3162 3773
rect 3328 3763 3330 3773
rect 3480 3763 3482 3773
rect 2774 3762 2780 3763
rect 2774 3758 2775 3762
rect 2779 3758 2780 3762
rect 2774 3757 2780 3758
rect 2974 3762 2980 3763
rect 2974 3758 2975 3762
rect 2979 3758 2980 3762
rect 2974 3757 2980 3758
rect 3158 3762 3164 3763
rect 3158 3758 3159 3762
rect 3163 3758 3164 3762
rect 3158 3757 3164 3758
rect 3326 3762 3332 3763
rect 3326 3758 3327 3762
rect 3331 3758 3332 3762
rect 3326 3757 3332 3758
rect 3478 3762 3484 3763
rect 3478 3758 3479 3762
rect 3483 3758 3484 3762
rect 3478 3757 3484 3758
rect 2698 3731 2704 3732
rect 2698 3727 2699 3731
rect 2703 3727 2704 3731
rect 2698 3726 2704 3727
rect 2886 3731 2892 3732
rect 2886 3727 2887 3731
rect 2891 3727 2892 3731
rect 2886 3726 2892 3727
rect 3142 3731 3148 3732
rect 3142 3727 3143 3731
rect 3147 3727 3148 3731
rect 3142 3726 3148 3727
rect 2700 3712 2702 3726
rect 2774 3721 2780 3722
rect 2774 3717 2775 3721
rect 2779 3717 2780 3721
rect 2774 3716 2780 3717
rect 2630 3711 2636 3712
rect 2630 3707 2631 3711
rect 2635 3707 2636 3711
rect 2630 3706 2636 3707
rect 2698 3711 2704 3712
rect 2698 3707 2699 3711
rect 2703 3707 2704 3711
rect 2698 3706 2704 3707
rect 2776 3695 2778 3716
rect 2071 3694 2075 3695
rect 2071 3689 2075 3690
rect 2111 3694 2115 3695
rect 2111 3689 2115 3690
rect 2255 3694 2259 3695
rect 2255 3689 2259 3690
rect 2335 3694 2339 3695
rect 2335 3689 2339 3690
rect 2439 3694 2443 3695
rect 2439 3689 2443 3690
rect 2559 3694 2563 3695
rect 2559 3689 2563 3690
rect 2623 3694 2627 3695
rect 2623 3689 2627 3690
rect 2775 3694 2779 3695
rect 2775 3689 2779 3690
rect 2815 3694 2819 3695
rect 2815 3689 2819 3690
rect 2050 3687 2056 3688
rect 847 3686 851 3687
rect 847 3681 851 3682
rect 903 3686 907 3687
rect 903 3681 907 3682
rect 983 3686 987 3687
rect 983 3681 987 3682
rect 1047 3686 1051 3687
rect 1047 3681 1051 3682
rect 1111 3686 1115 3687
rect 1111 3681 1115 3682
rect 1191 3686 1195 3687
rect 1191 3681 1195 3682
rect 1239 3686 1243 3687
rect 1239 3681 1243 3682
rect 1335 3686 1339 3687
rect 1350 3683 1351 3687
rect 1355 3683 1356 3687
rect 1350 3682 1356 3683
rect 1367 3686 1371 3687
rect 1335 3681 1339 3682
rect 1367 3681 1371 3682
rect 1479 3686 1483 3687
rect 1479 3681 1483 3682
rect 1495 3686 1499 3687
rect 1495 3681 1499 3682
rect 1631 3686 1635 3687
rect 1631 3681 1635 3682
rect 1767 3686 1771 3687
rect 1767 3681 1771 3682
rect 2031 3686 2035 3687
rect 2050 3683 2051 3687
rect 2055 3683 2056 3687
rect 2050 3682 2056 3683
rect 2031 3681 2035 3682
rect 904 3672 906 3681
rect 910 3679 916 3680
rect 910 3675 911 3679
rect 915 3675 916 3679
rect 910 3674 916 3675
rect 902 3671 908 3672
rect 902 3667 903 3671
rect 907 3667 908 3671
rect 912 3669 914 3674
rect 1048 3672 1050 3681
rect 1192 3672 1194 3681
rect 1336 3672 1338 3681
rect 1480 3672 1482 3681
rect 1046 3671 1052 3672
rect 902 3666 908 3667
rect 911 3668 915 3669
rect 1046 3667 1047 3671
rect 1051 3667 1052 3671
rect 1046 3666 1052 3667
rect 1190 3671 1196 3672
rect 1190 3667 1191 3671
rect 1195 3667 1196 3671
rect 1190 3666 1196 3667
rect 1334 3671 1340 3672
rect 1334 3667 1335 3671
rect 1339 3667 1340 3671
rect 1334 3666 1340 3667
rect 1478 3671 1484 3672
rect 1478 3667 1479 3671
rect 1483 3667 1484 3671
rect 1478 3666 1484 3667
rect 911 3663 915 3664
rect 1174 3663 1180 3664
rect 782 3659 788 3660
rect 782 3655 783 3659
rect 787 3655 788 3659
rect 1174 3659 1175 3663
rect 1179 3659 1180 3663
rect 1174 3658 1180 3659
rect 782 3654 788 3655
rect 758 3630 764 3631
rect 758 3626 759 3630
rect 763 3626 764 3630
rect 758 3625 764 3626
rect 902 3630 908 3631
rect 902 3626 903 3630
rect 907 3626 908 3630
rect 902 3625 908 3626
rect 1046 3630 1052 3631
rect 1046 3626 1047 3630
rect 1051 3626 1052 3630
rect 1046 3625 1052 3626
rect 760 3615 762 3625
rect 904 3615 906 3625
rect 1048 3615 1050 3625
rect 759 3614 763 3615
rect 759 3609 763 3610
rect 847 3614 851 3615
rect 847 3609 851 3610
rect 903 3614 907 3615
rect 903 3609 907 3610
rect 1023 3614 1027 3615
rect 1023 3609 1027 3610
rect 1047 3614 1051 3615
rect 1047 3609 1051 3610
rect 848 3599 850 3609
rect 1024 3599 1026 3609
rect 846 3598 852 3599
rect 846 3594 847 3598
rect 851 3594 852 3598
rect 846 3593 852 3594
rect 1022 3598 1028 3599
rect 1022 3594 1023 3598
rect 1027 3594 1028 3598
rect 1022 3593 1028 3594
rect 358 3567 364 3568
rect 358 3563 359 3567
rect 363 3563 364 3567
rect 358 3562 364 3563
rect 662 3567 668 3568
rect 662 3563 663 3567
rect 667 3563 668 3567
rect 662 3562 668 3563
rect 686 3567 692 3568
rect 686 3563 687 3567
rect 691 3563 692 3567
rect 686 3562 692 3563
rect 1038 3567 1044 3568
rect 1038 3563 1039 3567
rect 1043 3563 1044 3567
rect 1038 3562 1044 3563
rect 246 3557 252 3558
rect 246 3553 247 3557
rect 251 3553 252 3557
rect 246 3552 252 3553
rect 230 3531 236 3532
rect 248 3531 250 3552
rect 360 3540 362 3562
rect 374 3557 380 3558
rect 374 3553 375 3557
rect 379 3553 380 3557
rect 374 3552 380 3553
rect 518 3557 524 3558
rect 518 3553 519 3557
rect 523 3553 524 3557
rect 518 3552 524 3553
rect 358 3539 364 3540
rect 358 3535 359 3539
rect 363 3535 364 3539
rect 358 3534 364 3535
rect 376 3531 378 3552
rect 422 3547 428 3548
rect 422 3543 423 3547
rect 427 3543 428 3547
rect 422 3542 428 3543
rect 111 3530 115 3531
rect 111 3525 115 3526
rect 151 3530 155 3531
rect 230 3527 231 3531
rect 235 3527 236 3531
rect 230 3526 236 3527
rect 247 3530 251 3531
rect 151 3525 155 3526
rect 112 3497 114 3525
rect 152 3516 154 3525
rect 150 3515 156 3516
rect 150 3511 151 3515
rect 155 3511 156 3515
rect 150 3510 156 3511
rect 232 3508 234 3526
rect 247 3525 251 3526
rect 263 3530 267 3531
rect 263 3525 267 3526
rect 375 3530 379 3531
rect 375 3525 379 3526
rect 399 3530 403 3531
rect 399 3525 403 3526
rect 264 3516 266 3525
rect 400 3516 402 3525
rect 414 3523 420 3524
rect 414 3519 415 3523
rect 419 3519 420 3523
rect 414 3518 420 3519
rect 262 3515 268 3516
rect 262 3511 263 3515
rect 267 3511 268 3515
rect 262 3510 268 3511
rect 398 3515 404 3516
rect 398 3511 399 3515
rect 403 3511 404 3515
rect 398 3510 404 3511
rect 230 3507 236 3508
rect 230 3503 231 3507
rect 235 3503 236 3507
rect 230 3502 236 3503
rect 110 3496 116 3497
rect 110 3492 111 3496
rect 115 3492 116 3496
rect 110 3491 116 3492
rect 110 3479 116 3480
rect 110 3475 111 3479
rect 115 3475 116 3479
rect 110 3474 116 3475
rect 150 3474 156 3475
rect 112 3459 114 3474
rect 150 3470 151 3474
rect 155 3470 156 3474
rect 150 3469 156 3470
rect 262 3474 268 3475
rect 262 3470 263 3474
rect 267 3470 268 3474
rect 262 3469 268 3470
rect 398 3474 404 3475
rect 398 3470 399 3474
rect 403 3470 404 3474
rect 398 3469 404 3470
rect 152 3459 154 3469
rect 264 3459 266 3469
rect 400 3459 402 3469
rect 111 3458 115 3459
rect 111 3453 115 3454
rect 151 3458 155 3459
rect 151 3453 155 3454
rect 263 3458 267 3459
rect 263 3453 267 3454
rect 399 3458 403 3459
rect 399 3453 403 3454
rect 112 3438 114 3453
rect 152 3443 154 3453
rect 150 3442 156 3443
rect 150 3438 151 3442
rect 155 3438 156 3442
rect 110 3437 116 3438
rect 150 3437 156 3438
rect 110 3433 111 3437
rect 115 3433 116 3437
rect 110 3432 116 3433
rect 110 3420 116 3421
rect 110 3416 111 3420
rect 115 3416 116 3420
rect 110 3415 116 3416
rect 112 3363 114 3415
rect 416 3412 418 3518
rect 424 3504 426 3542
rect 520 3531 522 3552
rect 664 3540 666 3562
rect 678 3557 684 3558
rect 678 3553 679 3557
rect 683 3553 684 3557
rect 678 3552 684 3553
rect 846 3557 852 3558
rect 846 3553 847 3557
rect 851 3553 852 3557
rect 846 3552 852 3553
rect 1022 3557 1028 3558
rect 1022 3553 1023 3557
rect 1027 3553 1028 3557
rect 1022 3552 1028 3553
rect 662 3539 668 3540
rect 662 3535 663 3539
rect 667 3535 668 3539
rect 662 3534 668 3535
rect 680 3531 682 3552
rect 848 3531 850 3552
rect 950 3531 956 3532
rect 1024 3531 1026 3552
rect 519 3530 523 3531
rect 519 3525 523 3526
rect 543 3530 547 3531
rect 543 3525 547 3526
rect 679 3530 683 3531
rect 679 3525 683 3526
rect 687 3530 691 3531
rect 687 3525 691 3526
rect 831 3530 835 3531
rect 831 3525 835 3526
rect 847 3530 851 3531
rect 950 3527 951 3531
rect 955 3527 956 3531
rect 950 3526 956 3527
rect 967 3530 971 3531
rect 847 3525 851 3526
rect 544 3516 546 3525
rect 688 3516 690 3525
rect 832 3516 834 3525
rect 542 3515 548 3516
rect 542 3511 543 3515
rect 547 3511 548 3515
rect 542 3510 548 3511
rect 686 3515 692 3516
rect 686 3511 687 3515
rect 691 3511 692 3515
rect 686 3510 692 3511
rect 830 3515 836 3516
rect 830 3511 831 3515
rect 835 3511 836 3515
rect 830 3510 836 3511
rect 952 3508 954 3526
rect 967 3525 971 3526
rect 1023 3530 1027 3531
rect 1023 3525 1027 3526
rect 968 3516 970 3525
rect 1040 3524 1042 3562
rect 1176 3557 1178 3658
rect 2032 3653 2034 3681
rect 2030 3652 2036 3653
rect 2030 3648 2031 3652
rect 2035 3648 2036 3652
rect 2030 3647 2036 3648
rect 2030 3635 2036 3636
rect 2030 3631 2031 3635
rect 2035 3631 2036 3635
rect 1190 3630 1196 3631
rect 1190 3626 1191 3630
rect 1195 3626 1196 3630
rect 1190 3625 1196 3626
rect 1334 3630 1340 3631
rect 1334 3626 1335 3630
rect 1339 3626 1340 3630
rect 1334 3625 1340 3626
rect 1478 3630 1484 3631
rect 2030 3630 2036 3631
rect 1478 3626 1479 3630
rect 1483 3626 1484 3630
rect 1478 3625 1484 3626
rect 1192 3615 1194 3625
rect 1336 3615 1338 3625
rect 1480 3615 1482 3625
rect 2032 3615 2034 3630
rect 1191 3614 1195 3615
rect 1191 3609 1195 3610
rect 1207 3614 1211 3615
rect 1207 3609 1211 3610
rect 1335 3614 1339 3615
rect 1335 3609 1339 3610
rect 1391 3614 1395 3615
rect 1391 3609 1395 3610
rect 1479 3614 1483 3615
rect 1479 3609 1483 3610
rect 1575 3614 1579 3615
rect 1575 3609 1579 3610
rect 1767 3614 1771 3615
rect 1767 3609 1771 3610
rect 1935 3614 1939 3615
rect 1935 3609 1939 3610
rect 2031 3614 2035 3615
rect 2031 3609 2035 3610
rect 1208 3599 1210 3609
rect 1392 3599 1394 3609
rect 1576 3599 1578 3609
rect 1768 3599 1770 3609
rect 1936 3599 1938 3609
rect 1206 3598 1212 3599
rect 1206 3594 1207 3598
rect 1211 3594 1212 3598
rect 1206 3593 1212 3594
rect 1390 3598 1396 3599
rect 1390 3594 1391 3598
rect 1395 3594 1396 3598
rect 1390 3593 1396 3594
rect 1574 3598 1580 3599
rect 1574 3594 1575 3598
rect 1579 3594 1580 3598
rect 1574 3593 1580 3594
rect 1766 3598 1772 3599
rect 1766 3594 1767 3598
rect 1771 3594 1772 3598
rect 1766 3593 1772 3594
rect 1934 3598 1940 3599
rect 1934 3594 1935 3598
rect 1939 3594 1940 3598
rect 2032 3594 2034 3609
rect 1934 3593 1940 3594
rect 2030 3593 2036 3594
rect 2030 3589 2031 3593
rect 2035 3589 2036 3593
rect 2030 3588 2036 3589
rect 2030 3576 2036 3577
rect 2030 3572 2031 3576
rect 2035 3572 2036 3576
rect 2030 3571 2036 3572
rect 1750 3567 1756 3568
rect 1750 3563 1751 3567
rect 1755 3563 1756 3567
rect 1750 3562 1756 3563
rect 1878 3567 1884 3568
rect 1878 3563 1879 3567
rect 1883 3563 1884 3567
rect 1878 3562 1884 3563
rect 1206 3557 1212 3558
rect 1175 3556 1179 3557
rect 1206 3553 1207 3557
rect 1211 3553 1212 3557
rect 1206 3552 1212 3553
rect 1390 3557 1396 3558
rect 1574 3557 1580 3558
rect 1390 3553 1391 3557
rect 1395 3553 1396 3557
rect 1390 3552 1396 3553
rect 1463 3556 1467 3557
rect 1574 3553 1575 3557
rect 1579 3553 1580 3557
rect 1574 3552 1580 3553
rect 1175 3551 1179 3552
rect 1208 3531 1210 3552
rect 1392 3531 1394 3552
rect 1463 3551 1467 3552
rect 1464 3548 1466 3551
rect 1462 3547 1468 3548
rect 1462 3543 1463 3547
rect 1467 3543 1468 3547
rect 1462 3542 1468 3543
rect 1566 3531 1572 3532
rect 1576 3531 1578 3552
rect 1752 3548 1754 3562
rect 1766 3557 1772 3558
rect 1766 3553 1767 3557
rect 1771 3553 1772 3557
rect 1766 3552 1772 3553
rect 1646 3547 1652 3548
rect 1646 3543 1647 3547
rect 1651 3543 1652 3547
rect 1646 3542 1652 3543
rect 1750 3547 1756 3548
rect 1750 3543 1751 3547
rect 1755 3543 1756 3547
rect 1750 3542 1756 3543
rect 1095 3530 1099 3531
rect 1095 3525 1099 3526
rect 1207 3530 1211 3531
rect 1207 3525 1211 3526
rect 1223 3530 1227 3531
rect 1223 3525 1227 3526
rect 1343 3530 1347 3531
rect 1343 3525 1347 3526
rect 1391 3530 1395 3531
rect 1391 3525 1395 3526
rect 1463 3530 1467 3531
rect 1566 3527 1567 3531
rect 1571 3527 1572 3531
rect 1566 3526 1572 3527
rect 1575 3530 1579 3531
rect 1463 3525 1467 3526
rect 1038 3523 1044 3524
rect 1038 3519 1039 3523
rect 1043 3519 1044 3523
rect 1038 3518 1044 3519
rect 1096 3516 1098 3525
rect 1224 3516 1226 3525
rect 1344 3516 1346 3525
rect 1464 3516 1466 3525
rect 1534 3523 1540 3524
rect 1534 3519 1535 3523
rect 1539 3519 1540 3523
rect 1534 3518 1540 3519
rect 966 3515 972 3516
rect 966 3511 967 3515
rect 971 3511 972 3515
rect 966 3510 972 3511
rect 1094 3515 1100 3516
rect 1094 3511 1095 3515
rect 1099 3511 1100 3515
rect 1094 3510 1100 3511
rect 1222 3515 1228 3516
rect 1222 3511 1223 3515
rect 1227 3511 1228 3515
rect 1222 3510 1228 3511
rect 1342 3515 1348 3516
rect 1342 3511 1343 3515
rect 1347 3511 1348 3515
rect 1342 3510 1348 3511
rect 1462 3515 1468 3516
rect 1462 3511 1463 3515
rect 1467 3511 1468 3515
rect 1462 3510 1468 3511
rect 950 3507 956 3508
rect 422 3503 428 3504
rect 422 3499 423 3503
rect 427 3499 428 3503
rect 950 3503 951 3507
rect 955 3503 956 3507
rect 950 3502 956 3503
rect 1446 3507 1452 3508
rect 1446 3503 1447 3507
rect 1451 3503 1452 3507
rect 1446 3502 1452 3503
rect 422 3498 428 3499
rect 542 3474 548 3475
rect 542 3470 543 3474
rect 547 3470 548 3474
rect 542 3469 548 3470
rect 686 3474 692 3475
rect 686 3470 687 3474
rect 691 3470 692 3474
rect 686 3469 692 3470
rect 830 3474 836 3475
rect 830 3470 831 3474
rect 835 3470 836 3474
rect 830 3469 836 3470
rect 966 3474 972 3475
rect 966 3470 967 3474
rect 971 3470 972 3474
rect 966 3469 972 3470
rect 1094 3474 1100 3475
rect 1094 3470 1095 3474
rect 1099 3470 1100 3474
rect 1094 3469 1100 3470
rect 1222 3474 1228 3475
rect 1222 3470 1223 3474
rect 1227 3470 1228 3474
rect 1222 3469 1228 3470
rect 1342 3474 1348 3475
rect 1342 3470 1343 3474
rect 1347 3470 1348 3474
rect 1342 3469 1348 3470
rect 544 3459 546 3469
rect 688 3459 690 3469
rect 832 3459 834 3469
rect 968 3459 970 3469
rect 1096 3459 1098 3469
rect 1224 3459 1226 3469
rect 1344 3459 1346 3469
rect 423 3458 427 3459
rect 423 3453 427 3454
rect 543 3458 547 3459
rect 543 3453 547 3454
rect 687 3458 691 3459
rect 687 3453 691 3454
rect 743 3458 747 3459
rect 743 3453 747 3454
rect 831 3458 835 3459
rect 831 3453 835 3454
rect 967 3458 971 3459
rect 967 3453 971 3454
rect 1071 3458 1075 3459
rect 1071 3453 1075 3454
rect 1095 3458 1099 3459
rect 1095 3453 1099 3454
rect 1223 3458 1227 3459
rect 1223 3453 1227 3454
rect 1343 3458 1347 3459
rect 1343 3453 1347 3454
rect 1399 3458 1403 3459
rect 1399 3453 1403 3454
rect 424 3443 426 3453
rect 744 3443 746 3453
rect 1072 3443 1074 3453
rect 1400 3443 1402 3453
rect 422 3442 428 3443
rect 422 3438 423 3442
rect 427 3438 428 3442
rect 422 3437 428 3438
rect 742 3442 748 3443
rect 742 3438 743 3442
rect 747 3438 748 3442
rect 742 3437 748 3438
rect 1070 3442 1076 3443
rect 1070 3438 1071 3442
rect 1075 3438 1076 3442
rect 1070 3437 1076 3438
rect 1398 3442 1404 3443
rect 1398 3438 1399 3442
rect 1403 3438 1404 3442
rect 1398 3437 1404 3438
rect 406 3411 412 3412
rect 406 3407 407 3411
rect 411 3407 412 3411
rect 406 3406 412 3407
rect 414 3411 420 3412
rect 414 3407 415 3411
rect 419 3407 420 3411
rect 414 3406 420 3407
rect 150 3401 156 3402
rect 150 3397 151 3401
rect 155 3397 156 3401
rect 150 3396 156 3397
rect 152 3363 154 3396
rect 214 3391 220 3392
rect 214 3387 215 3391
rect 219 3387 220 3391
rect 214 3386 220 3387
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 151 3362 155 3363
rect 151 3357 155 3358
rect 112 3329 114 3357
rect 152 3348 154 3357
rect 150 3347 156 3348
rect 150 3343 151 3347
rect 155 3343 156 3347
rect 150 3342 156 3343
rect 216 3340 218 3386
rect 408 3384 410 3406
rect 422 3401 428 3402
rect 422 3397 423 3401
rect 427 3397 428 3401
rect 422 3396 428 3397
rect 742 3401 748 3402
rect 742 3397 743 3401
rect 747 3397 748 3401
rect 742 3396 748 3397
rect 1070 3401 1076 3402
rect 1070 3397 1071 3401
rect 1075 3397 1076 3401
rect 1070 3396 1076 3397
rect 1398 3401 1404 3402
rect 1398 3397 1399 3401
rect 1403 3397 1404 3401
rect 1398 3396 1404 3397
rect 406 3383 412 3384
rect 406 3379 407 3383
rect 411 3379 412 3383
rect 406 3378 412 3379
rect 424 3363 426 3396
rect 744 3363 746 3396
rect 1072 3363 1074 3396
rect 1400 3363 1402 3396
rect 1448 3392 1450 3502
rect 1462 3474 1468 3475
rect 1462 3470 1463 3474
rect 1467 3470 1468 3474
rect 1462 3469 1468 3470
rect 1464 3459 1466 3469
rect 1463 3458 1467 3459
rect 1463 3453 1467 3454
rect 1536 3412 1538 3518
rect 1568 3508 1570 3526
rect 1575 3525 1579 3526
rect 1583 3530 1587 3531
rect 1583 3525 1587 3526
rect 1584 3516 1586 3525
rect 1582 3515 1588 3516
rect 1582 3511 1583 3515
rect 1587 3511 1588 3515
rect 1582 3510 1588 3511
rect 1648 3508 1650 3542
rect 1768 3531 1770 3552
rect 1880 3548 1882 3562
rect 1934 3557 1940 3558
rect 1934 3553 1935 3557
rect 1939 3553 1940 3557
rect 1934 3552 1940 3553
rect 1878 3547 1884 3548
rect 1878 3543 1879 3547
rect 1883 3543 1884 3547
rect 1878 3542 1884 3543
rect 1936 3531 1938 3552
rect 2032 3531 2034 3571
rect 2052 3568 2054 3682
rect 2072 3661 2074 3689
rect 2112 3680 2114 3689
rect 2256 3680 2258 3689
rect 2440 3680 2442 3689
rect 2624 3680 2626 3689
rect 2816 3680 2818 3689
rect 2888 3688 2890 3726
rect 2974 3721 2980 3722
rect 2974 3717 2975 3721
rect 2979 3717 2980 3721
rect 2974 3716 2980 3717
rect 2976 3695 2978 3716
rect 3144 3696 3146 3726
rect 3158 3721 3164 3722
rect 3158 3717 3159 3721
rect 3163 3717 3164 3721
rect 3158 3716 3164 3717
rect 3326 3721 3332 3722
rect 3326 3717 3327 3721
rect 3331 3717 3332 3721
rect 3326 3716 3332 3717
rect 3478 3721 3484 3722
rect 3478 3717 3479 3721
rect 3483 3717 3484 3721
rect 3478 3716 3484 3717
rect 3142 3695 3148 3696
rect 3160 3695 3162 3716
rect 3328 3695 3330 3716
rect 3480 3695 3482 3716
rect 3552 3712 3554 3774
rect 3583 3773 3587 3774
rect 3623 3778 3627 3779
rect 3623 3773 3627 3774
rect 3624 3763 3626 3773
rect 3622 3762 3628 3763
rect 3622 3758 3623 3762
rect 3627 3758 3628 3762
rect 3622 3757 3628 3758
rect 3648 3732 3650 3838
rect 3752 3836 3754 3845
rect 3896 3836 3898 3845
rect 3750 3835 3756 3836
rect 3750 3831 3751 3835
rect 3755 3831 3756 3835
rect 3750 3830 3756 3831
rect 3894 3835 3900 3836
rect 3894 3831 3895 3835
rect 3899 3831 3900 3835
rect 3894 3830 3900 3831
rect 3966 3827 3972 3828
rect 3966 3823 3967 3827
rect 3971 3823 3972 3827
rect 3966 3822 3972 3823
rect 3750 3794 3756 3795
rect 3750 3790 3751 3794
rect 3755 3790 3756 3794
rect 3750 3789 3756 3790
rect 3894 3794 3900 3795
rect 3894 3790 3895 3794
rect 3899 3790 3900 3794
rect 3894 3789 3900 3790
rect 3752 3779 3754 3789
rect 3896 3779 3898 3789
rect 3751 3778 3755 3779
rect 3751 3773 3755 3774
rect 3767 3778 3771 3779
rect 3767 3773 3771 3774
rect 3895 3778 3899 3779
rect 3895 3773 3899 3774
rect 3768 3763 3770 3773
rect 3896 3763 3898 3773
rect 3766 3762 3772 3763
rect 3766 3758 3767 3762
rect 3771 3758 3772 3762
rect 3766 3757 3772 3758
rect 3894 3762 3900 3763
rect 3894 3758 3895 3762
rect 3899 3758 3900 3762
rect 3894 3757 3900 3758
rect 3646 3731 3652 3732
rect 3646 3727 3647 3731
rect 3651 3727 3652 3731
rect 3646 3726 3652 3727
rect 3622 3721 3628 3722
rect 3622 3717 3623 3721
rect 3627 3717 3628 3721
rect 3622 3716 3628 3717
rect 3766 3721 3772 3722
rect 3766 3717 3767 3721
rect 3771 3717 3772 3721
rect 3766 3716 3772 3717
rect 3894 3721 3900 3722
rect 3894 3717 3895 3721
rect 3899 3717 3900 3721
rect 3894 3716 3900 3717
rect 3550 3711 3556 3712
rect 3550 3707 3551 3711
rect 3555 3707 3556 3711
rect 3550 3706 3556 3707
rect 3624 3695 3626 3716
rect 3768 3695 3770 3716
rect 3896 3695 3898 3716
rect 3968 3712 3970 3822
rect 3992 3817 3994 3845
rect 3990 3816 3996 3817
rect 3990 3812 3991 3816
rect 3995 3812 3996 3816
rect 3990 3811 3996 3812
rect 3990 3799 3996 3800
rect 3990 3795 3991 3799
rect 3995 3795 3996 3799
rect 3990 3794 3996 3795
rect 3992 3779 3994 3794
rect 3991 3778 3995 3779
rect 3991 3773 3995 3774
rect 3992 3758 3994 3773
rect 3990 3757 3996 3758
rect 3990 3753 3991 3757
rect 3995 3753 3996 3757
rect 3990 3752 3996 3753
rect 3990 3740 3996 3741
rect 3990 3736 3991 3740
rect 3995 3736 3996 3740
rect 3990 3735 3996 3736
rect 3966 3711 3972 3712
rect 3966 3707 3967 3711
rect 3971 3707 3972 3711
rect 3966 3706 3972 3707
rect 3992 3695 3994 3735
rect 2975 3694 2979 3695
rect 2975 3689 2979 3690
rect 3007 3694 3011 3695
rect 3142 3691 3143 3695
rect 3147 3691 3148 3695
rect 3142 3690 3148 3691
rect 3159 3694 3163 3695
rect 3007 3689 3011 3690
rect 3159 3689 3163 3690
rect 3199 3694 3203 3695
rect 3199 3689 3203 3690
rect 3327 3694 3331 3695
rect 3327 3689 3331 3690
rect 3391 3694 3395 3695
rect 3391 3689 3395 3690
rect 3479 3694 3483 3695
rect 3479 3689 3483 3690
rect 3583 3694 3587 3695
rect 3583 3689 3587 3690
rect 3623 3694 3627 3695
rect 3623 3689 3627 3690
rect 3767 3694 3771 3695
rect 3767 3689 3771 3690
rect 3895 3694 3899 3695
rect 3895 3689 3899 3690
rect 3991 3694 3995 3695
rect 3991 3689 3995 3690
rect 2886 3687 2892 3688
rect 2886 3683 2887 3687
rect 2891 3683 2892 3687
rect 2886 3682 2892 3683
rect 3008 3680 3010 3689
rect 3200 3680 3202 3689
rect 3392 3680 3394 3689
rect 3584 3680 3586 3689
rect 2110 3679 2116 3680
rect 2110 3675 2111 3679
rect 2115 3675 2116 3679
rect 2110 3674 2116 3675
rect 2254 3679 2260 3680
rect 2254 3675 2255 3679
rect 2259 3675 2260 3679
rect 2254 3674 2260 3675
rect 2438 3679 2444 3680
rect 2438 3675 2439 3679
rect 2443 3675 2444 3679
rect 2438 3674 2444 3675
rect 2622 3679 2628 3680
rect 2622 3675 2623 3679
rect 2627 3675 2628 3679
rect 2622 3674 2628 3675
rect 2814 3679 2820 3680
rect 2814 3675 2815 3679
rect 2819 3675 2820 3679
rect 2814 3674 2820 3675
rect 3006 3679 3012 3680
rect 3006 3675 3007 3679
rect 3011 3675 3012 3679
rect 3006 3674 3012 3675
rect 3198 3679 3204 3680
rect 3198 3675 3199 3679
rect 3203 3675 3204 3679
rect 3198 3674 3204 3675
rect 3390 3679 3396 3680
rect 3390 3675 3391 3679
rect 3395 3675 3396 3679
rect 3390 3674 3396 3675
rect 3582 3679 3588 3680
rect 3582 3675 3583 3679
rect 3587 3675 3588 3679
rect 3582 3674 3588 3675
rect 3182 3671 3188 3672
rect 2430 3667 2436 3668
rect 2430 3663 2431 3667
rect 2435 3663 2436 3667
rect 3182 3667 3183 3671
rect 3187 3667 3188 3671
rect 3182 3666 3188 3667
rect 2430 3662 2436 3663
rect 2070 3660 2076 3661
rect 2070 3656 2071 3660
rect 2075 3656 2076 3660
rect 2070 3655 2076 3656
rect 2070 3643 2076 3644
rect 2070 3639 2071 3643
rect 2075 3639 2076 3643
rect 2070 3638 2076 3639
rect 2110 3638 2116 3639
rect 2072 3611 2074 3638
rect 2110 3634 2111 3638
rect 2115 3634 2116 3638
rect 2110 3633 2116 3634
rect 2254 3638 2260 3639
rect 2254 3634 2255 3638
rect 2259 3634 2260 3638
rect 2254 3633 2260 3634
rect 2112 3611 2114 3633
rect 2256 3611 2258 3633
rect 2071 3610 2075 3611
rect 2071 3605 2075 3606
rect 2111 3610 2115 3611
rect 2111 3605 2115 3606
rect 2255 3610 2259 3611
rect 2255 3605 2259 3606
rect 2359 3610 2363 3611
rect 2359 3605 2363 3606
rect 2072 3590 2074 3605
rect 2360 3595 2362 3605
rect 2358 3594 2364 3595
rect 2358 3590 2359 3594
rect 2363 3590 2364 3594
rect 2070 3589 2076 3590
rect 2358 3589 2364 3590
rect 2070 3585 2071 3589
rect 2075 3585 2076 3589
rect 2070 3584 2076 3585
rect 2070 3572 2076 3573
rect 2070 3568 2071 3572
rect 2075 3568 2076 3572
rect 2050 3567 2056 3568
rect 2070 3567 2076 3568
rect 2050 3563 2051 3567
rect 2055 3563 2056 3567
rect 2050 3562 2056 3563
rect 2072 3535 2074 3567
rect 2358 3553 2364 3554
rect 2358 3549 2359 3553
rect 2363 3549 2364 3553
rect 2358 3548 2364 3549
rect 2360 3535 2362 3548
rect 2432 3544 2434 3662
rect 2438 3638 2444 3639
rect 2438 3634 2439 3638
rect 2443 3634 2444 3638
rect 2438 3633 2444 3634
rect 2622 3638 2628 3639
rect 2622 3634 2623 3638
rect 2627 3634 2628 3638
rect 2622 3633 2628 3634
rect 2814 3638 2820 3639
rect 2814 3634 2815 3638
rect 2819 3634 2820 3638
rect 2814 3633 2820 3634
rect 3006 3638 3012 3639
rect 3006 3634 3007 3638
rect 3011 3634 3012 3638
rect 3006 3633 3012 3634
rect 2440 3611 2442 3633
rect 2624 3611 2626 3633
rect 2816 3611 2818 3633
rect 3008 3611 3010 3633
rect 2439 3610 2443 3611
rect 2439 3605 2443 3606
rect 2583 3610 2587 3611
rect 2583 3605 2587 3606
rect 2623 3610 2627 3611
rect 2623 3605 2627 3606
rect 2799 3610 2803 3611
rect 2799 3605 2803 3606
rect 2815 3610 2819 3611
rect 2815 3605 2819 3606
rect 3007 3610 3011 3611
rect 3007 3605 3011 3606
rect 2584 3595 2586 3605
rect 2800 3595 2802 3605
rect 3008 3595 3010 3605
rect 2582 3594 2588 3595
rect 2582 3590 2583 3594
rect 2587 3590 2588 3594
rect 2582 3589 2588 3590
rect 2798 3594 2804 3595
rect 2798 3590 2799 3594
rect 2803 3590 2804 3594
rect 2798 3589 2804 3590
rect 3006 3594 3012 3595
rect 3006 3590 3007 3594
rect 3011 3590 3012 3594
rect 3006 3589 3012 3590
rect 3184 3584 3186 3666
rect 3992 3661 3994 3689
rect 3990 3660 3996 3661
rect 3990 3656 3991 3660
rect 3995 3656 3996 3660
rect 3990 3655 3996 3656
rect 3990 3643 3996 3644
rect 3990 3639 3991 3643
rect 3995 3639 3996 3643
rect 3198 3638 3204 3639
rect 3198 3634 3199 3638
rect 3203 3634 3204 3638
rect 3198 3633 3204 3634
rect 3390 3638 3396 3639
rect 3390 3634 3391 3638
rect 3395 3634 3396 3638
rect 3390 3633 3396 3634
rect 3582 3638 3588 3639
rect 3990 3638 3996 3639
rect 3582 3634 3583 3638
rect 3587 3634 3588 3638
rect 3582 3633 3588 3634
rect 3200 3611 3202 3633
rect 3392 3611 3394 3633
rect 3584 3611 3586 3633
rect 3992 3611 3994 3638
rect 3199 3610 3203 3611
rect 3199 3605 3203 3606
rect 3215 3610 3219 3611
rect 3215 3605 3219 3606
rect 3391 3610 3395 3611
rect 3391 3605 3395 3606
rect 3431 3610 3435 3611
rect 3431 3605 3435 3606
rect 3583 3610 3587 3611
rect 3583 3605 3587 3606
rect 3991 3610 3995 3611
rect 3991 3605 3995 3606
rect 3216 3595 3218 3605
rect 3432 3595 3434 3605
rect 3214 3594 3220 3595
rect 3214 3590 3215 3594
rect 3219 3590 3220 3594
rect 3214 3589 3220 3590
rect 3430 3594 3436 3595
rect 3430 3590 3431 3594
rect 3435 3590 3436 3594
rect 3992 3590 3994 3605
rect 3430 3589 3436 3590
rect 3990 3589 3996 3590
rect 3990 3585 3991 3589
rect 3995 3585 3996 3589
rect 3990 3584 3996 3585
rect 3182 3583 3188 3584
rect 3182 3579 3183 3583
rect 3187 3579 3188 3583
rect 3182 3578 3188 3579
rect 3502 3583 3508 3584
rect 3502 3579 3503 3583
rect 3507 3579 3508 3583
rect 3502 3578 3508 3579
rect 2566 3563 2572 3564
rect 2566 3559 2567 3563
rect 2571 3559 2572 3563
rect 2990 3563 2996 3564
rect 2566 3558 2572 3559
rect 2646 3559 2652 3560
rect 2568 3544 2570 3558
rect 2646 3555 2647 3559
rect 2651 3555 2652 3559
rect 2990 3559 2991 3563
rect 2995 3559 2996 3563
rect 2990 3558 2996 3559
rect 2646 3554 2652 3555
rect 2582 3553 2588 3554
rect 2582 3549 2583 3553
rect 2587 3549 2588 3553
rect 2582 3548 2588 3549
rect 2430 3543 2436 3544
rect 2430 3539 2431 3543
rect 2435 3539 2436 3543
rect 2430 3538 2436 3539
rect 2566 3543 2572 3544
rect 2566 3539 2567 3543
rect 2571 3539 2572 3543
rect 2566 3538 2572 3539
rect 2584 3535 2586 3548
rect 2071 3534 2075 3535
rect 1711 3530 1715 3531
rect 1711 3525 1715 3526
rect 1767 3530 1771 3531
rect 1767 3525 1771 3526
rect 1935 3530 1939 3531
rect 1935 3525 1939 3526
rect 2031 3530 2035 3531
rect 2071 3529 2075 3530
rect 2359 3534 2363 3535
rect 2359 3529 2363 3530
rect 2439 3534 2443 3535
rect 2439 3529 2443 3530
rect 2575 3534 2579 3535
rect 2575 3529 2579 3530
rect 2583 3534 2587 3535
rect 2583 3529 2587 3530
rect 2031 3525 2035 3526
rect 1712 3516 1714 3525
rect 1710 3515 1716 3516
rect 1710 3511 1711 3515
rect 1715 3511 1716 3515
rect 1710 3510 1716 3511
rect 1566 3507 1572 3508
rect 1566 3503 1567 3507
rect 1571 3503 1572 3507
rect 1566 3502 1572 3503
rect 1646 3507 1652 3508
rect 1646 3503 1647 3507
rect 1651 3503 1652 3507
rect 1646 3502 1652 3503
rect 2032 3497 2034 3525
rect 2072 3501 2074 3529
rect 2440 3520 2442 3529
rect 2576 3520 2578 3529
rect 2648 3528 2650 3554
rect 2798 3553 2804 3554
rect 2798 3549 2799 3553
rect 2803 3549 2804 3553
rect 2798 3548 2804 3549
rect 2800 3535 2802 3548
rect 2992 3536 2994 3558
rect 3006 3553 3012 3554
rect 3006 3549 3007 3553
rect 3011 3549 3012 3553
rect 3006 3548 3012 3549
rect 3214 3553 3220 3554
rect 3214 3549 3215 3553
rect 3219 3549 3220 3553
rect 3214 3548 3220 3549
rect 3430 3553 3436 3554
rect 3430 3549 3431 3553
rect 3435 3549 3436 3553
rect 3430 3548 3436 3549
rect 2990 3535 2996 3536
rect 3008 3535 3010 3548
rect 3216 3535 3218 3548
rect 3432 3535 3434 3548
rect 3504 3544 3506 3578
rect 3990 3572 3996 3573
rect 3990 3568 3991 3572
rect 3995 3568 3996 3572
rect 3990 3567 3996 3568
rect 3502 3543 3508 3544
rect 3502 3539 3503 3543
rect 3507 3539 3508 3543
rect 3502 3538 3508 3539
rect 3992 3535 3994 3567
rect 2703 3534 2707 3535
rect 2703 3529 2707 3530
rect 2799 3534 2803 3535
rect 2799 3529 2803 3530
rect 2831 3534 2835 3535
rect 2831 3529 2835 3530
rect 2951 3534 2955 3535
rect 2990 3531 2991 3535
rect 2995 3531 2996 3535
rect 2990 3530 2996 3531
rect 3007 3534 3011 3535
rect 2951 3529 2955 3530
rect 3007 3529 3011 3530
rect 3071 3534 3075 3535
rect 3071 3529 3075 3530
rect 3199 3534 3203 3535
rect 3199 3529 3203 3530
rect 3215 3534 3219 3535
rect 3215 3529 3219 3530
rect 3327 3534 3331 3535
rect 3327 3529 3331 3530
rect 3431 3534 3435 3535
rect 3431 3529 3435 3530
rect 3991 3534 3995 3535
rect 3991 3529 3995 3530
rect 2646 3527 2652 3528
rect 2646 3523 2647 3527
rect 2651 3523 2652 3527
rect 2646 3522 2652 3523
rect 2704 3520 2706 3529
rect 2832 3520 2834 3529
rect 2952 3520 2954 3529
rect 3072 3520 3074 3529
rect 3200 3520 3202 3529
rect 3328 3520 3330 3529
rect 2438 3519 2444 3520
rect 2438 3515 2439 3519
rect 2443 3515 2444 3519
rect 2438 3514 2444 3515
rect 2574 3519 2580 3520
rect 2574 3515 2575 3519
rect 2579 3515 2580 3519
rect 2574 3514 2580 3515
rect 2702 3519 2708 3520
rect 2702 3515 2703 3519
rect 2707 3515 2708 3519
rect 2702 3514 2708 3515
rect 2830 3519 2836 3520
rect 2830 3515 2831 3519
rect 2835 3515 2836 3519
rect 2830 3514 2836 3515
rect 2950 3519 2956 3520
rect 2950 3515 2951 3519
rect 2955 3515 2956 3519
rect 2950 3514 2956 3515
rect 3070 3519 3076 3520
rect 3070 3515 3071 3519
rect 3075 3515 3076 3519
rect 3070 3514 3076 3515
rect 3198 3519 3204 3520
rect 3198 3515 3199 3519
rect 3203 3515 3204 3519
rect 3198 3514 3204 3515
rect 3326 3519 3332 3520
rect 3326 3515 3327 3519
rect 3331 3515 3332 3519
rect 3326 3514 3332 3515
rect 2786 3511 2792 3512
rect 2430 3507 2436 3508
rect 2430 3503 2431 3507
rect 2435 3503 2436 3507
rect 2786 3507 2787 3511
rect 2791 3507 2792 3511
rect 2786 3506 2792 3507
rect 2430 3502 2436 3503
rect 2070 3500 2076 3501
rect 2030 3496 2036 3497
rect 2030 3492 2031 3496
rect 2035 3492 2036 3496
rect 2070 3496 2071 3500
rect 2075 3496 2076 3500
rect 2070 3495 2076 3496
rect 2030 3491 2036 3492
rect 2070 3483 2076 3484
rect 2030 3479 2036 3480
rect 2030 3475 2031 3479
rect 2035 3475 2036 3479
rect 2070 3479 2071 3483
rect 2075 3479 2076 3483
rect 2070 3478 2076 3479
rect 1582 3474 1588 3475
rect 1582 3470 1583 3474
rect 1587 3470 1588 3474
rect 1582 3469 1588 3470
rect 1710 3474 1716 3475
rect 2030 3474 2036 3475
rect 1710 3470 1711 3474
rect 1715 3470 1716 3474
rect 1710 3469 1716 3470
rect 1584 3459 1586 3469
rect 1712 3459 1714 3469
rect 2032 3459 2034 3474
rect 2072 3463 2074 3478
rect 2071 3462 2075 3463
rect 1583 3458 1587 3459
rect 1583 3453 1587 3454
rect 1711 3458 1715 3459
rect 1711 3453 1715 3454
rect 2031 3458 2035 3459
rect 2071 3457 2075 3458
rect 2359 3462 2363 3463
rect 2359 3457 2363 3458
rect 2031 3453 2035 3454
rect 2032 3438 2034 3453
rect 2072 3442 2074 3457
rect 2360 3447 2362 3457
rect 2358 3446 2364 3447
rect 2358 3442 2359 3446
rect 2363 3442 2364 3446
rect 2070 3441 2076 3442
rect 2358 3441 2364 3442
rect 2030 3437 2036 3438
rect 2030 3433 2031 3437
rect 2035 3433 2036 3437
rect 2070 3437 2071 3441
rect 2075 3437 2076 3441
rect 2070 3436 2076 3437
rect 2030 3432 2036 3433
rect 2070 3424 2076 3425
rect 2030 3420 2036 3421
rect 2030 3416 2031 3420
rect 2035 3416 2036 3420
rect 2070 3420 2071 3424
rect 2075 3420 2076 3424
rect 2070 3419 2076 3420
rect 2030 3415 2036 3416
rect 1534 3411 1540 3412
rect 1534 3407 1535 3411
rect 1539 3407 1540 3411
rect 1534 3406 1540 3407
rect 1446 3391 1452 3392
rect 1446 3387 1447 3391
rect 1451 3387 1452 3391
rect 1446 3386 1452 3387
rect 2032 3363 2034 3415
rect 2072 3363 2074 3419
rect 2358 3405 2364 3406
rect 2358 3401 2359 3405
rect 2363 3401 2364 3405
rect 2358 3400 2364 3401
rect 2360 3363 2362 3400
rect 2432 3396 2434 3502
rect 2438 3478 2444 3479
rect 2438 3474 2439 3478
rect 2443 3474 2444 3478
rect 2438 3473 2444 3474
rect 2574 3478 2580 3479
rect 2574 3474 2575 3478
rect 2579 3474 2580 3478
rect 2574 3473 2580 3474
rect 2702 3478 2708 3479
rect 2702 3474 2703 3478
rect 2707 3474 2708 3478
rect 2702 3473 2708 3474
rect 2440 3463 2442 3473
rect 2576 3463 2578 3473
rect 2704 3463 2706 3473
rect 2439 3462 2443 3463
rect 2439 3457 2443 3458
rect 2463 3462 2467 3463
rect 2463 3457 2467 3458
rect 2567 3462 2571 3463
rect 2567 3457 2571 3458
rect 2575 3462 2579 3463
rect 2575 3457 2579 3458
rect 2671 3462 2675 3463
rect 2671 3457 2675 3458
rect 2703 3462 2707 3463
rect 2703 3457 2707 3458
rect 2775 3462 2779 3463
rect 2775 3457 2779 3458
rect 2464 3447 2466 3457
rect 2568 3447 2570 3457
rect 2672 3447 2674 3457
rect 2776 3447 2778 3457
rect 2462 3446 2468 3447
rect 2462 3442 2463 3446
rect 2467 3442 2468 3446
rect 2462 3441 2468 3442
rect 2566 3446 2572 3447
rect 2566 3442 2567 3446
rect 2571 3442 2572 3446
rect 2566 3441 2572 3442
rect 2670 3446 2676 3447
rect 2670 3442 2671 3446
rect 2675 3442 2676 3446
rect 2670 3441 2676 3442
rect 2774 3446 2780 3447
rect 2774 3442 2775 3446
rect 2779 3442 2780 3446
rect 2774 3441 2780 3442
rect 2446 3415 2452 3416
rect 2446 3411 2447 3415
rect 2451 3411 2452 3415
rect 2446 3410 2452 3411
rect 2486 3415 2492 3416
rect 2486 3411 2487 3415
rect 2491 3411 2492 3415
rect 2486 3410 2492 3411
rect 2638 3415 2644 3416
rect 2638 3411 2639 3415
rect 2643 3411 2644 3415
rect 2638 3410 2644 3411
rect 2448 3396 2450 3410
rect 2462 3405 2468 3406
rect 2462 3401 2463 3405
rect 2467 3401 2468 3405
rect 2462 3400 2468 3401
rect 2430 3395 2436 3396
rect 2430 3391 2431 3395
rect 2435 3391 2436 3395
rect 2430 3390 2436 3391
rect 2446 3395 2452 3396
rect 2446 3391 2447 3395
rect 2451 3391 2452 3395
rect 2446 3390 2452 3391
rect 2464 3363 2466 3400
rect 319 3362 323 3363
rect 319 3357 323 3358
rect 423 3362 427 3363
rect 423 3357 427 3358
rect 527 3362 531 3363
rect 527 3357 531 3358
rect 743 3362 747 3363
rect 743 3357 747 3358
rect 959 3362 963 3363
rect 959 3357 963 3358
rect 1071 3362 1075 3363
rect 1071 3357 1075 3358
rect 1167 3362 1171 3363
rect 1167 3357 1171 3358
rect 1367 3362 1371 3363
rect 1367 3357 1371 3358
rect 1399 3362 1403 3363
rect 1399 3357 1403 3358
rect 1559 3362 1563 3363
rect 1559 3357 1563 3358
rect 1751 3362 1755 3363
rect 1751 3357 1755 3358
rect 1935 3362 1939 3363
rect 1935 3357 1939 3358
rect 2031 3362 2035 3363
rect 2031 3357 2035 3358
rect 2071 3362 2075 3363
rect 2071 3357 2075 3358
rect 2359 3362 2363 3363
rect 2359 3357 2363 3358
rect 2439 3362 2443 3363
rect 2439 3357 2443 3358
rect 2463 3362 2467 3363
rect 2463 3357 2467 3358
rect 320 3348 322 3357
rect 528 3348 530 3357
rect 744 3348 746 3357
rect 960 3348 962 3357
rect 994 3355 1000 3356
rect 994 3351 995 3355
rect 999 3351 1000 3355
rect 994 3350 1000 3351
rect 318 3347 324 3348
rect 318 3343 319 3347
rect 323 3343 324 3347
rect 318 3342 324 3343
rect 526 3347 532 3348
rect 526 3343 527 3347
rect 531 3343 532 3347
rect 526 3342 532 3343
rect 742 3347 748 3348
rect 742 3343 743 3347
rect 747 3343 748 3347
rect 742 3342 748 3343
rect 958 3347 964 3348
rect 958 3343 959 3347
rect 963 3343 964 3347
rect 958 3342 964 3343
rect 214 3339 220 3340
rect 214 3335 215 3339
rect 219 3335 220 3339
rect 214 3334 220 3335
rect 110 3328 116 3329
rect 110 3324 111 3328
rect 115 3324 116 3328
rect 110 3323 116 3324
rect 110 3311 116 3312
rect 110 3307 111 3311
rect 115 3307 116 3311
rect 110 3306 116 3307
rect 150 3306 156 3307
rect 112 3283 114 3306
rect 150 3302 151 3306
rect 155 3302 156 3306
rect 150 3301 156 3302
rect 318 3306 324 3307
rect 318 3302 319 3306
rect 323 3302 324 3306
rect 318 3301 324 3302
rect 526 3306 532 3307
rect 526 3302 527 3306
rect 531 3302 532 3306
rect 526 3301 532 3302
rect 742 3306 748 3307
rect 742 3302 743 3306
rect 747 3302 748 3306
rect 742 3301 748 3302
rect 958 3306 964 3307
rect 958 3302 959 3306
rect 963 3302 964 3306
rect 958 3301 964 3302
rect 152 3283 154 3301
rect 320 3283 322 3301
rect 528 3283 530 3301
rect 744 3283 746 3301
rect 960 3283 962 3301
rect 996 3292 998 3350
rect 1168 3348 1170 3357
rect 1368 3348 1370 3357
rect 1560 3348 1562 3357
rect 1752 3348 1754 3357
rect 1936 3348 1938 3357
rect 2002 3355 2008 3356
rect 2002 3351 2003 3355
rect 2007 3351 2008 3355
rect 2002 3350 2008 3351
rect 1166 3347 1172 3348
rect 1166 3343 1167 3347
rect 1171 3343 1172 3347
rect 1166 3342 1172 3343
rect 1366 3347 1372 3348
rect 1366 3343 1367 3347
rect 1371 3343 1372 3347
rect 1366 3342 1372 3343
rect 1558 3347 1564 3348
rect 1558 3343 1559 3347
rect 1563 3343 1564 3347
rect 1558 3342 1564 3343
rect 1750 3347 1756 3348
rect 1750 3343 1751 3347
rect 1755 3343 1756 3347
rect 1750 3342 1756 3343
rect 1934 3347 1940 3348
rect 1934 3343 1935 3347
rect 1939 3343 1940 3347
rect 1934 3342 1940 3343
rect 1166 3306 1172 3307
rect 1166 3302 1167 3306
rect 1171 3302 1172 3306
rect 1166 3301 1172 3302
rect 1366 3306 1372 3307
rect 1366 3302 1367 3306
rect 1371 3302 1372 3306
rect 1366 3301 1372 3302
rect 1558 3306 1564 3307
rect 1558 3302 1559 3306
rect 1563 3302 1564 3306
rect 1558 3301 1564 3302
rect 1750 3306 1756 3307
rect 1750 3302 1751 3306
rect 1755 3302 1756 3306
rect 1750 3301 1756 3302
rect 1934 3306 1940 3307
rect 1934 3302 1935 3306
rect 1939 3302 1940 3306
rect 1934 3301 1940 3302
rect 994 3291 1000 3292
rect 994 3287 995 3291
rect 999 3287 1000 3291
rect 994 3286 1000 3287
rect 1168 3283 1170 3301
rect 1368 3283 1370 3301
rect 1560 3283 1562 3301
rect 1752 3283 1754 3301
rect 1936 3283 1938 3301
rect 111 3282 115 3283
rect 111 3277 115 3278
rect 151 3282 155 3283
rect 151 3277 155 3278
rect 311 3282 315 3283
rect 311 3277 315 3278
rect 319 3282 323 3283
rect 319 3277 323 3278
rect 479 3282 483 3283
rect 479 3277 483 3278
rect 527 3282 531 3283
rect 527 3277 531 3278
rect 655 3282 659 3283
rect 655 3277 659 3278
rect 743 3282 747 3283
rect 743 3277 747 3278
rect 847 3282 851 3283
rect 847 3277 851 3278
rect 959 3282 963 3283
rect 959 3277 963 3278
rect 1039 3282 1043 3283
rect 1039 3277 1043 3278
rect 1167 3282 1171 3283
rect 1167 3277 1171 3278
rect 1231 3282 1235 3283
rect 1231 3277 1235 3278
rect 1367 3282 1371 3283
rect 1367 3277 1371 3278
rect 1431 3282 1435 3283
rect 1431 3277 1435 3278
rect 1559 3282 1563 3283
rect 1559 3277 1563 3278
rect 1631 3282 1635 3283
rect 1631 3277 1635 3278
rect 1751 3282 1755 3283
rect 1751 3277 1755 3278
rect 1831 3282 1835 3283
rect 1831 3277 1835 3278
rect 1935 3282 1939 3283
rect 1935 3277 1939 3278
rect 112 3262 114 3277
rect 312 3267 314 3277
rect 480 3267 482 3277
rect 656 3267 658 3277
rect 848 3267 850 3277
rect 1040 3267 1042 3277
rect 1232 3267 1234 3277
rect 1432 3267 1434 3277
rect 1632 3267 1634 3277
rect 1832 3267 1834 3277
rect 310 3266 316 3267
rect 310 3262 311 3266
rect 315 3262 316 3266
rect 110 3261 116 3262
rect 310 3261 316 3262
rect 478 3266 484 3267
rect 478 3262 479 3266
rect 483 3262 484 3266
rect 478 3261 484 3262
rect 654 3266 660 3267
rect 654 3262 655 3266
rect 659 3262 660 3266
rect 654 3261 660 3262
rect 846 3266 852 3267
rect 846 3262 847 3266
rect 851 3262 852 3266
rect 846 3261 852 3262
rect 1038 3266 1044 3267
rect 1038 3262 1039 3266
rect 1043 3262 1044 3266
rect 1038 3261 1044 3262
rect 1230 3266 1236 3267
rect 1230 3262 1231 3266
rect 1235 3262 1236 3266
rect 1230 3261 1236 3262
rect 1430 3266 1436 3267
rect 1430 3262 1431 3266
rect 1435 3262 1436 3266
rect 1430 3261 1436 3262
rect 1630 3266 1636 3267
rect 1630 3262 1631 3266
rect 1635 3262 1636 3266
rect 1630 3261 1636 3262
rect 1830 3266 1836 3267
rect 1830 3262 1831 3266
rect 1835 3262 1836 3266
rect 1830 3261 1836 3262
rect 110 3257 111 3261
rect 115 3257 116 3261
rect 110 3256 116 3257
rect 110 3244 116 3245
rect 110 3240 111 3244
rect 115 3240 116 3244
rect 110 3239 116 3240
rect 112 3207 114 3239
rect 2004 3236 2006 3350
rect 2032 3329 2034 3357
rect 2072 3329 2074 3357
rect 2440 3348 2442 3357
rect 2488 3356 2490 3410
rect 2566 3405 2572 3406
rect 2566 3401 2567 3405
rect 2571 3401 2572 3405
rect 2566 3400 2572 3401
rect 2568 3363 2570 3400
rect 2543 3362 2547 3363
rect 2543 3357 2547 3358
rect 2567 3362 2571 3363
rect 2567 3357 2571 3358
rect 2486 3355 2492 3356
rect 2486 3351 2487 3355
rect 2491 3351 2492 3355
rect 2486 3350 2492 3351
rect 2544 3348 2546 3357
rect 2640 3356 2642 3410
rect 2670 3405 2676 3406
rect 2670 3401 2671 3405
rect 2675 3401 2676 3405
rect 2670 3400 2676 3401
rect 2774 3405 2780 3406
rect 2774 3401 2775 3405
rect 2779 3401 2780 3405
rect 2774 3400 2780 3401
rect 2672 3363 2674 3400
rect 2776 3363 2778 3400
rect 2788 3388 2790 3506
rect 3992 3501 3994 3529
rect 3990 3500 3996 3501
rect 3990 3496 3991 3500
rect 3995 3496 3996 3500
rect 3990 3495 3996 3496
rect 3990 3483 3996 3484
rect 3990 3479 3991 3483
rect 3995 3479 3996 3483
rect 2830 3478 2836 3479
rect 2830 3474 2831 3478
rect 2835 3474 2836 3478
rect 2830 3473 2836 3474
rect 2950 3478 2956 3479
rect 2950 3474 2951 3478
rect 2955 3474 2956 3478
rect 2950 3473 2956 3474
rect 3070 3478 3076 3479
rect 3070 3474 3071 3478
rect 3075 3474 3076 3478
rect 3070 3473 3076 3474
rect 3198 3478 3204 3479
rect 3198 3474 3199 3478
rect 3203 3474 3204 3478
rect 3198 3473 3204 3474
rect 3326 3478 3332 3479
rect 3990 3478 3996 3479
rect 3326 3474 3327 3478
rect 3331 3474 3332 3478
rect 3326 3473 3332 3474
rect 2832 3463 2834 3473
rect 2952 3463 2954 3473
rect 3072 3463 3074 3473
rect 3200 3463 3202 3473
rect 3328 3463 3330 3473
rect 3992 3463 3994 3478
rect 2831 3462 2835 3463
rect 2831 3457 2835 3458
rect 2879 3462 2883 3463
rect 2879 3457 2883 3458
rect 2951 3462 2955 3463
rect 2951 3457 2955 3458
rect 2983 3462 2987 3463
rect 2983 3457 2987 3458
rect 3071 3462 3075 3463
rect 3071 3457 3075 3458
rect 3087 3462 3091 3463
rect 3087 3457 3091 3458
rect 3191 3462 3195 3463
rect 3191 3457 3195 3458
rect 3199 3462 3203 3463
rect 3199 3457 3203 3458
rect 3327 3462 3331 3463
rect 3327 3457 3331 3458
rect 3991 3462 3995 3463
rect 3991 3457 3995 3458
rect 2880 3447 2882 3457
rect 2984 3447 2986 3457
rect 3088 3447 3090 3457
rect 3192 3447 3194 3457
rect 2878 3446 2884 3447
rect 2878 3442 2879 3446
rect 2883 3442 2884 3446
rect 2878 3441 2884 3442
rect 2982 3446 2988 3447
rect 2982 3442 2983 3446
rect 2987 3442 2988 3446
rect 2982 3441 2988 3442
rect 3086 3446 3092 3447
rect 3086 3442 3087 3446
rect 3091 3442 3092 3446
rect 3086 3441 3092 3442
rect 3190 3446 3196 3447
rect 3190 3442 3191 3446
rect 3195 3442 3196 3446
rect 3992 3442 3994 3457
rect 3190 3441 3196 3442
rect 3990 3441 3996 3442
rect 3990 3437 3991 3441
rect 3995 3437 3996 3441
rect 3990 3436 3996 3437
rect 3990 3424 3996 3425
rect 3990 3420 3991 3424
rect 3995 3420 3996 3424
rect 3990 3419 3996 3420
rect 2878 3405 2884 3406
rect 2878 3401 2879 3405
rect 2883 3401 2884 3405
rect 2878 3400 2884 3401
rect 2982 3405 2988 3406
rect 2982 3401 2983 3405
rect 2987 3401 2988 3405
rect 2982 3400 2988 3401
rect 3086 3405 3092 3406
rect 3086 3401 3087 3405
rect 3091 3401 3092 3405
rect 3086 3400 3092 3401
rect 3190 3405 3196 3406
rect 3190 3401 3191 3405
rect 3195 3401 3196 3405
rect 3190 3400 3196 3401
rect 2786 3387 2792 3388
rect 2786 3383 2787 3387
rect 2791 3383 2792 3387
rect 2786 3382 2792 3383
rect 2838 3363 2844 3364
rect 2880 3363 2882 3400
rect 2984 3363 2986 3400
rect 3088 3363 3090 3400
rect 3192 3363 3194 3400
rect 3992 3363 3994 3419
rect 2647 3362 2651 3363
rect 2647 3357 2651 3358
rect 2671 3362 2675 3363
rect 2671 3357 2675 3358
rect 2751 3362 2755 3363
rect 2751 3357 2755 3358
rect 2775 3362 2779 3363
rect 2838 3359 2839 3363
rect 2843 3359 2844 3363
rect 2838 3358 2844 3359
rect 2855 3362 2859 3363
rect 2775 3357 2779 3358
rect 2638 3355 2644 3356
rect 2638 3351 2639 3355
rect 2643 3351 2644 3355
rect 2638 3350 2644 3351
rect 2648 3348 2650 3357
rect 2752 3348 2754 3357
rect 2438 3347 2444 3348
rect 2438 3343 2439 3347
rect 2443 3343 2444 3347
rect 2438 3342 2444 3343
rect 2542 3347 2548 3348
rect 2542 3343 2543 3347
rect 2547 3343 2548 3347
rect 2542 3342 2548 3343
rect 2646 3347 2652 3348
rect 2646 3343 2647 3347
rect 2651 3343 2652 3347
rect 2646 3342 2652 3343
rect 2750 3347 2756 3348
rect 2750 3343 2751 3347
rect 2755 3343 2756 3347
rect 2750 3342 2756 3343
rect 2840 3340 2842 3358
rect 2855 3357 2859 3358
rect 2879 3362 2883 3363
rect 2879 3357 2883 3358
rect 2959 3362 2963 3363
rect 2959 3357 2963 3358
rect 2983 3362 2987 3363
rect 2983 3357 2987 3358
rect 3087 3362 3091 3363
rect 3087 3357 3091 3358
rect 3191 3362 3195 3363
rect 3191 3357 3195 3358
rect 3991 3362 3995 3363
rect 3991 3357 3995 3358
rect 2856 3348 2858 3357
rect 2960 3348 2962 3357
rect 2854 3347 2860 3348
rect 2854 3343 2855 3347
rect 2859 3343 2860 3347
rect 2854 3342 2860 3343
rect 2958 3347 2964 3348
rect 2958 3343 2959 3347
rect 2963 3343 2964 3347
rect 2958 3342 2964 3343
rect 2606 3339 2612 3340
rect 2606 3335 2607 3339
rect 2611 3335 2612 3339
rect 2606 3334 2612 3335
rect 2838 3339 2844 3340
rect 2838 3335 2839 3339
rect 2843 3335 2844 3339
rect 2838 3334 2844 3335
rect 2918 3339 2924 3340
rect 2918 3335 2919 3339
rect 2923 3335 2924 3339
rect 2918 3334 2924 3335
rect 2030 3328 2036 3329
rect 2030 3324 2031 3328
rect 2035 3324 2036 3328
rect 2030 3323 2036 3324
rect 2070 3328 2076 3329
rect 2070 3324 2071 3328
rect 2075 3324 2076 3328
rect 2070 3323 2076 3324
rect 2030 3311 2036 3312
rect 2030 3307 2031 3311
rect 2035 3307 2036 3311
rect 2030 3306 2036 3307
rect 2070 3311 2076 3312
rect 2070 3307 2071 3311
rect 2075 3307 2076 3311
rect 2070 3306 2076 3307
rect 2438 3306 2444 3307
rect 2032 3283 2034 3306
rect 2072 3291 2074 3306
rect 2438 3302 2439 3306
rect 2443 3302 2444 3306
rect 2438 3301 2444 3302
rect 2542 3306 2548 3307
rect 2542 3302 2543 3306
rect 2547 3302 2548 3306
rect 2542 3301 2548 3302
rect 2440 3291 2442 3301
rect 2544 3291 2546 3301
rect 2071 3290 2075 3291
rect 2071 3285 2075 3286
rect 2439 3290 2443 3291
rect 2439 3285 2443 3286
rect 2527 3290 2531 3291
rect 2527 3285 2531 3286
rect 2543 3290 2547 3291
rect 2543 3285 2547 3286
rect 2031 3282 2035 3283
rect 2031 3277 2035 3278
rect 2032 3262 2034 3277
rect 2072 3270 2074 3285
rect 2528 3275 2530 3285
rect 2526 3274 2532 3275
rect 2526 3270 2527 3274
rect 2531 3270 2532 3274
rect 2070 3269 2076 3270
rect 2526 3269 2532 3270
rect 2070 3265 2071 3269
rect 2075 3265 2076 3269
rect 2070 3264 2076 3265
rect 2030 3261 2036 3262
rect 2030 3257 2031 3261
rect 2035 3257 2036 3261
rect 2030 3256 2036 3257
rect 2070 3252 2076 3253
rect 2070 3248 2071 3252
rect 2075 3248 2076 3252
rect 2070 3247 2076 3248
rect 2030 3244 2036 3245
rect 2030 3240 2031 3244
rect 2035 3240 2036 3244
rect 2030 3239 2036 3240
rect 1254 3235 1260 3236
rect 1254 3231 1255 3235
rect 1259 3231 1260 3235
rect 1254 3230 1260 3231
rect 2002 3235 2008 3236
rect 2002 3231 2003 3235
rect 2007 3231 2008 3235
rect 2002 3230 2008 3231
rect 310 3225 316 3226
rect 310 3221 311 3225
rect 315 3221 316 3225
rect 310 3220 316 3221
rect 478 3225 484 3226
rect 478 3221 479 3225
rect 483 3221 484 3225
rect 478 3220 484 3221
rect 654 3225 660 3226
rect 654 3221 655 3225
rect 659 3221 660 3225
rect 654 3220 660 3221
rect 846 3225 852 3226
rect 846 3221 847 3225
rect 851 3221 852 3225
rect 846 3220 852 3221
rect 1038 3225 1044 3226
rect 1038 3221 1039 3225
rect 1043 3221 1044 3225
rect 1038 3220 1044 3221
rect 1230 3225 1236 3226
rect 1230 3221 1231 3225
rect 1235 3221 1236 3225
rect 1230 3220 1236 3221
rect 312 3207 314 3220
rect 480 3207 482 3220
rect 656 3207 658 3220
rect 848 3207 850 3220
rect 1040 3207 1042 3220
rect 1046 3215 1052 3216
rect 1046 3211 1047 3215
rect 1051 3211 1052 3215
rect 1046 3210 1052 3211
rect 111 3206 115 3207
rect 111 3201 115 3202
rect 311 3206 315 3207
rect 311 3201 315 3202
rect 479 3206 483 3207
rect 479 3201 483 3202
rect 623 3206 627 3207
rect 623 3201 627 3202
rect 655 3206 659 3207
rect 655 3201 659 3202
rect 759 3206 763 3207
rect 759 3201 763 3202
rect 847 3206 851 3207
rect 847 3201 851 3202
rect 903 3206 907 3207
rect 903 3201 907 3202
rect 1039 3206 1043 3207
rect 1039 3201 1043 3202
rect 112 3173 114 3201
rect 624 3192 626 3201
rect 743 3196 747 3197
rect 760 3192 762 3201
rect 904 3192 906 3201
rect 1048 3197 1050 3210
rect 1232 3207 1234 3220
rect 1055 3206 1059 3207
rect 1055 3201 1059 3202
rect 1207 3206 1211 3207
rect 1207 3201 1211 3202
rect 1231 3206 1235 3207
rect 1231 3201 1235 3202
rect 1047 3196 1051 3197
rect 1056 3192 1058 3201
rect 1126 3199 1132 3200
rect 1126 3195 1127 3199
rect 1131 3195 1132 3199
rect 1126 3194 1132 3195
rect 622 3191 628 3192
rect 743 3191 747 3192
rect 758 3191 764 3192
rect 622 3187 623 3191
rect 627 3187 628 3191
rect 622 3186 628 3187
rect 744 3184 746 3191
rect 758 3187 759 3191
rect 763 3187 764 3191
rect 758 3186 764 3187
rect 902 3191 908 3192
rect 1047 3191 1051 3192
rect 1054 3191 1060 3192
rect 902 3187 903 3191
rect 907 3187 908 3191
rect 902 3186 908 3187
rect 1054 3187 1055 3191
rect 1059 3187 1060 3191
rect 1054 3186 1060 3187
rect 742 3183 748 3184
rect 742 3179 743 3183
rect 747 3179 748 3183
rect 742 3178 748 3179
rect 110 3172 116 3173
rect 110 3168 111 3172
rect 115 3168 116 3172
rect 110 3167 116 3168
rect 110 3155 116 3156
rect 110 3151 111 3155
rect 115 3151 116 3155
rect 110 3150 116 3151
rect 622 3150 628 3151
rect 112 3135 114 3150
rect 622 3146 623 3150
rect 627 3146 628 3150
rect 622 3145 628 3146
rect 758 3150 764 3151
rect 758 3146 759 3150
rect 763 3146 764 3150
rect 758 3145 764 3146
rect 902 3150 908 3151
rect 902 3146 903 3150
rect 907 3146 908 3150
rect 902 3145 908 3146
rect 1054 3150 1060 3151
rect 1054 3146 1055 3150
rect 1059 3146 1060 3150
rect 1054 3145 1060 3146
rect 624 3135 626 3145
rect 760 3135 762 3145
rect 904 3135 906 3145
rect 1056 3135 1058 3145
rect 111 3134 115 3135
rect 111 3129 115 3130
rect 599 3134 603 3135
rect 599 3129 603 3130
rect 623 3134 627 3135
rect 623 3129 627 3130
rect 703 3134 707 3135
rect 703 3129 707 3130
rect 759 3134 763 3135
rect 759 3129 763 3130
rect 807 3134 811 3135
rect 807 3129 811 3130
rect 903 3134 907 3135
rect 903 3129 907 3130
rect 911 3134 915 3135
rect 911 3129 915 3130
rect 1039 3134 1043 3135
rect 1039 3129 1043 3130
rect 1055 3134 1059 3135
rect 1055 3129 1059 3130
rect 112 3114 114 3129
rect 600 3119 602 3129
rect 704 3119 706 3129
rect 808 3119 810 3129
rect 912 3119 914 3129
rect 1040 3119 1042 3129
rect 598 3118 604 3119
rect 598 3114 599 3118
rect 603 3114 604 3118
rect 110 3113 116 3114
rect 598 3113 604 3114
rect 702 3118 708 3119
rect 702 3114 703 3118
rect 707 3114 708 3118
rect 702 3113 708 3114
rect 806 3118 812 3119
rect 806 3114 807 3118
rect 811 3114 812 3118
rect 806 3113 812 3114
rect 910 3118 916 3119
rect 910 3114 911 3118
rect 915 3114 916 3118
rect 910 3113 916 3114
rect 1038 3118 1044 3119
rect 1038 3114 1039 3118
rect 1043 3114 1044 3118
rect 1038 3113 1044 3114
rect 110 3109 111 3113
rect 115 3109 116 3113
rect 110 3108 116 3109
rect 110 3096 116 3097
rect 110 3092 111 3096
rect 115 3092 116 3096
rect 110 3091 116 3092
rect 112 3055 114 3091
rect 1128 3088 1130 3194
rect 1208 3192 1210 3201
rect 1256 3200 1258 3230
rect 1430 3225 1436 3226
rect 1430 3221 1431 3225
rect 1435 3221 1436 3225
rect 1430 3220 1436 3221
rect 1630 3225 1636 3226
rect 1630 3221 1631 3225
rect 1635 3221 1636 3225
rect 1630 3220 1636 3221
rect 1830 3225 1836 3226
rect 1830 3221 1831 3225
rect 1835 3221 1836 3225
rect 1830 3220 1836 3221
rect 1432 3207 1434 3220
rect 1632 3207 1634 3220
rect 1774 3215 1780 3216
rect 1774 3211 1775 3215
rect 1779 3211 1780 3215
rect 1774 3210 1780 3211
rect 1351 3206 1355 3207
rect 1351 3201 1355 3202
rect 1431 3206 1435 3207
rect 1431 3201 1435 3202
rect 1503 3206 1507 3207
rect 1503 3201 1507 3202
rect 1631 3206 1635 3207
rect 1631 3201 1635 3202
rect 1655 3206 1659 3207
rect 1655 3201 1659 3202
rect 1254 3199 1260 3200
rect 1254 3195 1255 3199
rect 1259 3195 1260 3199
rect 1254 3194 1260 3195
rect 1352 3192 1354 3201
rect 1504 3192 1506 3201
rect 1656 3192 1658 3201
rect 1206 3191 1212 3192
rect 1206 3187 1207 3191
rect 1211 3187 1212 3191
rect 1206 3186 1212 3187
rect 1350 3191 1356 3192
rect 1350 3187 1351 3191
rect 1355 3187 1356 3191
rect 1350 3186 1356 3187
rect 1502 3191 1508 3192
rect 1502 3187 1503 3191
rect 1507 3187 1508 3191
rect 1502 3186 1508 3187
rect 1654 3191 1660 3192
rect 1654 3187 1655 3191
rect 1659 3187 1660 3191
rect 1654 3186 1660 3187
rect 1776 3184 1778 3210
rect 1832 3207 1834 3220
rect 2032 3207 2034 3239
rect 2072 3219 2074 3247
rect 2526 3233 2532 3234
rect 2526 3229 2527 3233
rect 2531 3229 2532 3233
rect 2526 3228 2532 3229
rect 2528 3219 2530 3228
rect 2599 3223 2605 3224
rect 2599 3219 2600 3223
rect 2604 3222 2605 3223
rect 2608 3222 2610 3334
rect 2646 3306 2652 3307
rect 2646 3302 2647 3306
rect 2651 3302 2652 3306
rect 2646 3301 2652 3302
rect 2750 3306 2756 3307
rect 2750 3302 2751 3306
rect 2755 3302 2756 3306
rect 2750 3301 2756 3302
rect 2854 3306 2860 3307
rect 2854 3302 2855 3306
rect 2859 3302 2860 3306
rect 2854 3301 2860 3302
rect 2648 3291 2650 3301
rect 2752 3291 2754 3301
rect 2856 3291 2858 3301
rect 2631 3290 2635 3291
rect 2631 3285 2635 3286
rect 2647 3290 2651 3291
rect 2647 3285 2651 3286
rect 2735 3290 2739 3291
rect 2735 3285 2739 3286
rect 2751 3290 2755 3291
rect 2751 3285 2755 3286
rect 2839 3290 2843 3291
rect 2839 3285 2843 3286
rect 2855 3290 2859 3291
rect 2855 3285 2859 3286
rect 2632 3275 2634 3285
rect 2736 3275 2738 3285
rect 2840 3275 2842 3285
rect 2630 3274 2636 3275
rect 2630 3270 2631 3274
rect 2635 3270 2636 3274
rect 2630 3269 2636 3270
rect 2734 3274 2740 3275
rect 2734 3270 2735 3274
rect 2739 3270 2740 3274
rect 2734 3269 2740 3270
rect 2838 3274 2844 3275
rect 2838 3270 2839 3274
rect 2843 3270 2844 3274
rect 2838 3269 2844 3270
rect 2614 3243 2620 3244
rect 2614 3239 2615 3243
rect 2619 3239 2620 3243
rect 2614 3238 2620 3239
rect 2718 3243 2724 3244
rect 2718 3239 2719 3243
rect 2723 3239 2724 3243
rect 2718 3238 2724 3239
rect 2604 3220 2610 3222
rect 2616 3220 2618 3238
rect 2630 3233 2636 3234
rect 2630 3229 2631 3233
rect 2635 3229 2636 3233
rect 2720 3229 2722 3238
rect 2734 3233 2740 3234
rect 2734 3229 2735 3233
rect 2739 3229 2740 3233
rect 2630 3228 2636 3229
rect 2719 3228 2723 3229
rect 2734 3228 2740 3229
rect 2838 3233 2844 3234
rect 2838 3229 2839 3233
rect 2843 3229 2844 3233
rect 2838 3228 2844 3229
rect 2604 3219 2605 3220
rect 2071 3218 2075 3219
rect 2071 3213 2075 3214
rect 2399 3218 2403 3219
rect 2399 3213 2403 3214
rect 2527 3218 2531 3219
rect 2527 3213 2531 3214
rect 2551 3218 2555 3219
rect 2599 3218 2605 3219
rect 2614 3219 2620 3220
rect 2632 3219 2634 3228
rect 2719 3223 2723 3224
rect 2736 3219 2738 3228
rect 2840 3219 2842 3228
rect 2911 3223 2917 3224
rect 2911 3219 2912 3223
rect 2916 3222 2917 3223
rect 2920 3222 2922 3334
rect 3992 3329 3994 3357
rect 3990 3328 3996 3329
rect 3990 3324 3991 3328
rect 3995 3324 3996 3328
rect 3990 3323 3996 3324
rect 3990 3311 3996 3312
rect 3990 3307 3991 3311
rect 3995 3307 3996 3311
rect 2958 3306 2964 3307
rect 3990 3306 3996 3307
rect 2958 3302 2959 3306
rect 2963 3302 2964 3306
rect 2958 3301 2964 3302
rect 2960 3291 2962 3301
rect 3992 3291 3994 3306
rect 2943 3290 2947 3291
rect 2943 3285 2947 3286
rect 2959 3290 2963 3291
rect 2959 3285 2963 3286
rect 3047 3290 3051 3291
rect 3047 3285 3051 3286
rect 3151 3290 3155 3291
rect 3151 3285 3155 3286
rect 3255 3290 3259 3291
rect 3255 3285 3259 3286
rect 3991 3290 3995 3291
rect 3991 3285 3995 3286
rect 2944 3275 2946 3285
rect 3048 3275 3050 3285
rect 3152 3275 3154 3285
rect 3256 3275 3258 3285
rect 2942 3274 2948 3275
rect 2942 3270 2943 3274
rect 2947 3270 2948 3274
rect 2942 3269 2948 3270
rect 3046 3274 3052 3275
rect 3046 3270 3047 3274
rect 3051 3270 3052 3274
rect 3046 3269 3052 3270
rect 3150 3274 3156 3275
rect 3150 3270 3151 3274
rect 3155 3270 3156 3274
rect 3150 3269 3156 3270
rect 3254 3274 3260 3275
rect 3254 3270 3255 3274
rect 3259 3270 3260 3274
rect 3992 3270 3994 3285
rect 3254 3269 3260 3270
rect 3990 3269 3996 3270
rect 3990 3265 3991 3269
rect 3995 3265 3996 3269
rect 3990 3264 3996 3265
rect 3990 3252 3996 3253
rect 3990 3248 3991 3252
rect 3995 3248 3996 3252
rect 3990 3247 3996 3248
rect 3030 3243 3036 3244
rect 3030 3239 3031 3243
rect 3035 3239 3036 3243
rect 3030 3238 3036 3239
rect 3174 3243 3180 3244
rect 3174 3239 3175 3243
rect 3179 3239 3180 3243
rect 3174 3238 3180 3239
rect 2942 3233 2948 3234
rect 2942 3229 2943 3233
rect 2947 3229 2948 3233
rect 2942 3228 2948 3229
rect 3015 3228 3019 3229
rect 2916 3220 2922 3222
rect 2916 3219 2917 3220
rect 2944 3219 2946 3228
rect 3032 3224 3034 3238
rect 3046 3233 3052 3234
rect 3046 3229 3047 3233
rect 3051 3229 3052 3233
rect 3046 3228 3052 3229
rect 3150 3233 3156 3234
rect 3150 3229 3151 3233
rect 3155 3229 3156 3233
rect 3150 3228 3156 3229
rect 3014 3223 3020 3224
rect 3014 3219 3015 3223
rect 3019 3219 3020 3223
rect 2614 3215 2615 3219
rect 2619 3215 2620 3219
rect 2614 3214 2620 3215
rect 2631 3218 2635 3219
rect 2551 3213 2555 3214
rect 2631 3213 2635 3214
rect 2695 3218 2699 3219
rect 2695 3213 2699 3214
rect 2735 3218 2739 3219
rect 2735 3213 2739 3214
rect 2839 3218 2843 3219
rect 2911 3218 2917 3219
rect 2943 3218 2947 3219
rect 2839 3213 2843 3214
rect 2943 3213 2947 3214
rect 2975 3218 2979 3219
rect 3014 3218 3020 3219
rect 3030 3223 3036 3224
rect 3030 3219 3031 3223
rect 3035 3219 3036 3223
rect 3048 3219 3050 3228
rect 3152 3219 3154 3228
rect 3030 3218 3036 3219
rect 3047 3218 3051 3219
rect 2975 3213 2979 3214
rect 3047 3213 3051 3214
rect 3111 3218 3115 3219
rect 3111 3213 3115 3214
rect 3151 3218 3155 3219
rect 3151 3213 3155 3214
rect 1807 3206 1811 3207
rect 1807 3201 1811 3202
rect 1831 3206 1835 3207
rect 1831 3201 1835 3202
rect 1935 3206 1939 3207
rect 1935 3201 1939 3202
rect 2031 3206 2035 3207
rect 2031 3201 2035 3202
rect 1808 3192 1810 3201
rect 1936 3192 1938 3201
rect 2006 3199 2012 3200
rect 2006 3195 2007 3199
rect 2011 3195 2012 3199
rect 2006 3194 2012 3195
rect 1806 3191 1812 3192
rect 1806 3187 1807 3191
rect 1811 3187 1812 3191
rect 1806 3186 1812 3187
rect 1934 3191 1940 3192
rect 1934 3187 1935 3191
rect 1939 3187 1940 3191
rect 1934 3186 1940 3187
rect 1638 3183 1644 3184
rect 1638 3179 1639 3183
rect 1643 3179 1644 3183
rect 1638 3178 1644 3179
rect 1774 3183 1780 3184
rect 1774 3179 1775 3183
rect 1779 3179 1780 3183
rect 1774 3178 1780 3179
rect 1206 3150 1212 3151
rect 1206 3146 1207 3150
rect 1211 3146 1212 3150
rect 1206 3145 1212 3146
rect 1350 3150 1356 3151
rect 1350 3146 1351 3150
rect 1355 3146 1356 3150
rect 1350 3145 1356 3146
rect 1502 3150 1508 3151
rect 1502 3146 1503 3150
rect 1507 3146 1508 3150
rect 1502 3145 1508 3146
rect 1208 3135 1210 3145
rect 1352 3135 1354 3145
rect 1504 3135 1506 3145
rect 1183 3134 1187 3135
rect 1183 3129 1187 3130
rect 1207 3134 1211 3135
rect 1207 3129 1211 3130
rect 1351 3134 1355 3135
rect 1351 3129 1355 3130
rect 1359 3134 1363 3135
rect 1359 3129 1363 3130
rect 1503 3134 1507 3135
rect 1503 3129 1507 3130
rect 1551 3134 1555 3135
rect 1551 3129 1555 3130
rect 1184 3119 1186 3129
rect 1360 3119 1362 3129
rect 1552 3119 1554 3129
rect 1182 3118 1188 3119
rect 1182 3114 1183 3118
rect 1187 3114 1188 3118
rect 1182 3113 1188 3114
rect 1358 3118 1364 3119
rect 1358 3114 1359 3118
rect 1363 3114 1364 3118
rect 1358 3113 1364 3114
rect 1550 3118 1556 3119
rect 1550 3114 1551 3118
rect 1555 3114 1556 3118
rect 1550 3113 1556 3114
rect 686 3087 692 3088
rect 686 3083 687 3087
rect 691 3083 692 3087
rect 686 3082 692 3083
rect 790 3087 796 3088
rect 790 3083 791 3087
rect 795 3083 796 3087
rect 790 3082 796 3083
rect 894 3087 900 3088
rect 894 3083 895 3087
rect 899 3083 900 3087
rect 894 3082 900 3083
rect 1022 3087 1028 3088
rect 1022 3083 1023 3087
rect 1027 3083 1028 3087
rect 1022 3082 1028 3083
rect 1126 3087 1132 3088
rect 1126 3083 1127 3087
rect 1131 3083 1132 3087
rect 1126 3082 1132 3083
rect 598 3077 604 3078
rect 598 3073 599 3077
rect 603 3073 604 3077
rect 598 3072 604 3073
rect 398 3055 404 3056
rect 600 3055 602 3072
rect 688 3068 690 3082
rect 702 3077 708 3078
rect 702 3073 703 3077
rect 707 3073 708 3077
rect 702 3072 708 3073
rect 662 3067 668 3068
rect 662 3063 663 3067
rect 667 3063 668 3067
rect 662 3062 668 3063
rect 686 3067 692 3068
rect 686 3063 687 3067
rect 691 3063 692 3067
rect 686 3062 692 3063
rect 111 3054 115 3055
rect 111 3049 115 3050
rect 311 3054 315 3055
rect 398 3051 399 3055
rect 403 3051 404 3055
rect 398 3050 404 3051
rect 415 3054 419 3055
rect 311 3049 315 3050
rect 112 3021 114 3049
rect 312 3040 314 3049
rect 310 3039 316 3040
rect 310 3035 311 3039
rect 315 3035 316 3039
rect 310 3034 316 3035
rect 400 3032 402 3050
rect 415 3049 419 3050
rect 527 3054 531 3055
rect 527 3049 531 3050
rect 599 3054 603 3055
rect 599 3049 603 3050
rect 639 3054 643 3055
rect 639 3049 643 3050
rect 416 3040 418 3049
rect 528 3040 530 3049
rect 598 3043 604 3044
rect 414 3039 420 3040
rect 414 3035 415 3039
rect 419 3035 420 3039
rect 414 3034 420 3035
rect 526 3039 532 3040
rect 526 3035 527 3039
rect 531 3035 532 3039
rect 598 3039 599 3043
rect 603 3039 604 3043
rect 640 3040 642 3049
rect 598 3038 604 3039
rect 638 3039 644 3040
rect 526 3034 532 3035
rect 398 3031 404 3032
rect 398 3027 399 3031
rect 403 3027 404 3031
rect 398 3026 404 3027
rect 110 3020 116 3021
rect 110 3016 111 3020
rect 115 3016 116 3020
rect 110 3015 116 3016
rect 110 3003 116 3004
rect 110 2999 111 3003
rect 115 2999 116 3003
rect 110 2998 116 2999
rect 310 2998 316 2999
rect 112 2975 114 2998
rect 310 2994 311 2998
rect 315 2994 316 2998
rect 310 2993 316 2994
rect 414 2998 420 2999
rect 414 2994 415 2998
rect 419 2994 420 2998
rect 414 2993 420 2994
rect 526 2998 532 2999
rect 526 2994 527 2998
rect 531 2994 532 2998
rect 526 2993 532 2994
rect 312 2975 314 2993
rect 416 2975 418 2993
rect 528 2975 530 2993
rect 111 2974 115 2975
rect 111 2969 115 2970
rect 151 2974 155 2975
rect 151 2969 155 2970
rect 271 2974 275 2975
rect 271 2969 275 2970
rect 311 2974 315 2975
rect 311 2969 315 2970
rect 415 2974 419 2975
rect 415 2969 419 2970
rect 431 2974 435 2975
rect 431 2969 435 2970
rect 527 2974 531 2975
rect 527 2969 531 2970
rect 112 2954 114 2969
rect 152 2959 154 2969
rect 272 2959 274 2969
rect 432 2959 434 2969
rect 150 2958 156 2959
rect 150 2954 151 2958
rect 155 2954 156 2958
rect 110 2953 116 2954
rect 150 2953 156 2954
rect 270 2958 276 2959
rect 270 2954 271 2958
rect 275 2954 276 2958
rect 270 2953 276 2954
rect 430 2958 436 2959
rect 430 2954 431 2958
rect 435 2954 436 2958
rect 430 2953 436 2954
rect 110 2949 111 2953
rect 115 2949 116 2953
rect 110 2948 116 2949
rect 110 2936 116 2937
rect 110 2932 111 2936
rect 115 2932 116 2936
rect 110 2931 116 2932
rect 112 2891 114 2931
rect 600 2928 602 3038
rect 638 3035 639 3039
rect 643 3035 644 3039
rect 638 3034 644 3035
rect 664 3028 666 3062
rect 704 3055 706 3072
rect 792 3068 794 3082
rect 806 3077 812 3078
rect 806 3073 807 3077
rect 811 3073 812 3077
rect 806 3072 812 3073
rect 790 3067 796 3068
rect 790 3063 791 3067
rect 795 3063 796 3067
rect 790 3062 796 3063
rect 808 3055 810 3072
rect 896 3068 898 3082
rect 910 3077 916 3078
rect 910 3073 911 3077
rect 915 3073 916 3077
rect 910 3072 916 3073
rect 894 3067 900 3068
rect 894 3063 895 3067
rect 899 3063 900 3067
rect 894 3062 900 3063
rect 912 3055 914 3072
rect 1024 3068 1026 3082
rect 1038 3077 1044 3078
rect 1038 3073 1039 3077
rect 1043 3073 1044 3077
rect 1038 3072 1044 3073
rect 1182 3077 1188 3078
rect 1182 3073 1183 3077
rect 1187 3073 1188 3077
rect 1182 3072 1188 3073
rect 1358 3077 1364 3078
rect 1358 3073 1359 3077
rect 1363 3073 1364 3077
rect 1358 3072 1364 3073
rect 1550 3077 1556 3078
rect 1550 3073 1551 3077
rect 1555 3073 1556 3077
rect 1640 3076 1642 3178
rect 1654 3150 1660 3151
rect 1654 3146 1655 3150
rect 1659 3146 1660 3150
rect 1654 3145 1660 3146
rect 1806 3150 1812 3151
rect 1806 3146 1807 3150
rect 1811 3146 1812 3150
rect 1806 3145 1812 3146
rect 1934 3150 1940 3151
rect 1934 3146 1935 3150
rect 1939 3146 1940 3150
rect 1934 3145 1940 3146
rect 1656 3135 1658 3145
rect 1808 3135 1810 3145
rect 1936 3135 1938 3145
rect 1655 3134 1659 3135
rect 1655 3129 1659 3130
rect 1751 3134 1755 3135
rect 1751 3129 1755 3130
rect 1807 3134 1811 3135
rect 1807 3129 1811 3130
rect 1935 3134 1939 3135
rect 1935 3129 1939 3130
rect 1752 3119 1754 3129
rect 1936 3119 1938 3129
rect 1750 3118 1756 3119
rect 1750 3114 1751 3118
rect 1755 3114 1756 3118
rect 1750 3113 1756 3114
rect 1934 3118 1940 3119
rect 1934 3114 1935 3118
rect 1939 3114 1940 3118
rect 1934 3113 1940 3114
rect 2008 3088 2010 3194
rect 2032 3173 2034 3201
rect 2072 3185 2074 3213
rect 2400 3204 2402 3213
rect 2552 3204 2554 3213
rect 2696 3204 2698 3213
rect 2840 3204 2842 3213
rect 2976 3204 2978 3213
rect 3112 3204 3114 3213
rect 3176 3212 3178 3238
rect 3254 3233 3260 3234
rect 3254 3229 3255 3233
rect 3259 3229 3260 3233
rect 3254 3228 3260 3229
rect 3256 3219 3258 3228
rect 3992 3219 3994 3247
rect 3247 3218 3251 3219
rect 3247 3213 3251 3214
rect 3255 3218 3259 3219
rect 3255 3213 3259 3214
rect 3391 3218 3395 3219
rect 3391 3213 3395 3214
rect 3991 3218 3995 3219
rect 3991 3213 3995 3214
rect 3174 3211 3180 3212
rect 3174 3207 3175 3211
rect 3179 3207 3180 3211
rect 3174 3206 3180 3207
rect 3248 3204 3250 3213
rect 3392 3204 3394 3213
rect 3398 3211 3404 3212
rect 3398 3207 3399 3211
rect 3403 3207 3404 3211
rect 3398 3206 3404 3207
rect 2398 3203 2404 3204
rect 2398 3199 2399 3203
rect 2403 3199 2404 3203
rect 2398 3198 2404 3199
rect 2550 3203 2556 3204
rect 2550 3199 2551 3203
rect 2555 3199 2556 3203
rect 2550 3198 2556 3199
rect 2694 3203 2700 3204
rect 2694 3199 2695 3203
rect 2699 3199 2700 3203
rect 2694 3198 2700 3199
rect 2838 3203 2844 3204
rect 2838 3199 2839 3203
rect 2843 3199 2844 3203
rect 2838 3198 2844 3199
rect 2974 3203 2980 3204
rect 2974 3199 2975 3203
rect 2979 3199 2980 3203
rect 2974 3198 2980 3199
rect 3110 3203 3116 3204
rect 3110 3199 3111 3203
rect 3115 3199 3116 3203
rect 3110 3198 3116 3199
rect 3246 3203 3252 3204
rect 3246 3199 3247 3203
rect 3251 3199 3252 3203
rect 3246 3198 3252 3199
rect 3390 3203 3396 3204
rect 3390 3199 3391 3203
rect 3395 3199 3396 3203
rect 3390 3198 3396 3199
rect 3400 3197 3402 3206
rect 2959 3196 2963 3197
rect 3399 3196 3403 3197
rect 2414 3191 2420 3192
rect 2414 3187 2415 3191
rect 2419 3187 2420 3191
rect 2958 3191 2959 3196
rect 2963 3191 2964 3196
rect 2958 3190 2964 3191
rect 3262 3191 3268 3192
rect 3399 3191 3403 3192
rect 2414 3186 2420 3187
rect 3262 3187 3263 3191
rect 3267 3187 3268 3191
rect 3262 3186 3268 3187
rect 2070 3184 2076 3185
rect 2070 3180 2071 3184
rect 2075 3180 2076 3184
rect 2070 3179 2076 3180
rect 2030 3172 2036 3173
rect 2030 3168 2031 3172
rect 2035 3168 2036 3172
rect 2030 3167 2036 3168
rect 2070 3167 2076 3168
rect 2070 3163 2071 3167
rect 2075 3163 2076 3167
rect 2070 3162 2076 3163
rect 2398 3162 2404 3163
rect 2030 3155 2036 3156
rect 2030 3151 2031 3155
rect 2035 3151 2036 3155
rect 2030 3150 2036 3151
rect 2032 3135 2034 3150
rect 2072 3135 2074 3162
rect 2398 3158 2399 3162
rect 2403 3158 2404 3162
rect 2398 3157 2404 3158
rect 2400 3135 2402 3157
rect 2031 3134 2035 3135
rect 2031 3129 2035 3130
rect 2071 3134 2075 3135
rect 2071 3129 2075 3130
rect 2111 3134 2115 3135
rect 2111 3129 2115 3130
rect 2343 3134 2347 3135
rect 2343 3129 2347 3130
rect 2399 3134 2403 3135
rect 2399 3129 2403 3130
rect 2032 3114 2034 3129
rect 2072 3114 2074 3129
rect 2112 3119 2114 3129
rect 2344 3119 2346 3129
rect 2110 3118 2116 3119
rect 2110 3114 2111 3118
rect 2115 3114 2116 3118
rect 2030 3113 2036 3114
rect 2030 3109 2031 3113
rect 2035 3109 2036 3113
rect 2030 3108 2036 3109
rect 2070 3113 2076 3114
rect 2110 3113 2116 3114
rect 2342 3118 2348 3119
rect 2342 3114 2343 3118
rect 2347 3114 2348 3118
rect 2342 3113 2348 3114
rect 2070 3109 2071 3113
rect 2075 3109 2076 3113
rect 2070 3108 2076 3109
rect 2030 3096 2036 3097
rect 2030 3092 2031 3096
rect 2035 3092 2036 3096
rect 2030 3091 2036 3092
rect 2070 3096 2076 3097
rect 2070 3092 2071 3096
rect 2075 3092 2076 3096
rect 2070 3091 2076 3092
rect 2006 3087 2012 3088
rect 2006 3083 2007 3087
rect 2011 3083 2012 3087
rect 2006 3082 2012 3083
rect 1750 3077 1756 3078
rect 1550 3072 1556 3073
rect 1638 3075 1644 3076
rect 1022 3067 1028 3068
rect 1022 3063 1023 3067
rect 1027 3063 1028 3067
rect 1022 3062 1028 3063
rect 958 3055 964 3056
rect 1040 3055 1042 3072
rect 1166 3067 1172 3068
rect 1166 3063 1167 3067
rect 1171 3063 1172 3067
rect 1166 3062 1172 3063
rect 703 3054 707 3055
rect 703 3049 707 3050
rect 751 3054 755 3055
rect 751 3049 755 3050
rect 807 3054 811 3055
rect 807 3049 811 3050
rect 863 3054 867 3055
rect 863 3049 867 3050
rect 911 3054 915 3055
rect 958 3051 959 3055
rect 963 3051 964 3055
rect 958 3050 964 3051
rect 975 3054 979 3055
rect 911 3049 915 3050
rect 752 3040 754 3049
rect 864 3040 866 3049
rect 750 3039 756 3040
rect 750 3035 751 3039
rect 755 3035 756 3039
rect 750 3034 756 3035
rect 862 3039 868 3040
rect 862 3035 863 3039
rect 867 3035 868 3039
rect 862 3034 868 3035
rect 960 3032 962 3050
rect 975 3049 979 3050
rect 1039 3054 1043 3055
rect 1039 3049 1043 3050
rect 1095 3054 1099 3055
rect 1095 3049 1099 3050
rect 976 3040 978 3049
rect 1096 3040 1098 3049
rect 1168 3048 1170 3062
rect 1184 3055 1186 3072
rect 1360 3055 1362 3072
rect 1552 3055 1554 3072
rect 1638 3071 1639 3075
rect 1643 3071 1644 3075
rect 1750 3073 1751 3077
rect 1755 3073 1756 3077
rect 1750 3072 1756 3073
rect 1934 3077 1940 3078
rect 1934 3073 1935 3077
rect 1939 3073 1940 3077
rect 1934 3072 1940 3073
rect 1638 3070 1644 3071
rect 1752 3055 1754 3072
rect 1936 3055 1938 3072
rect 2032 3055 2034 3091
rect 2072 3059 2074 3091
rect 2110 3077 2116 3078
rect 2110 3073 2111 3077
rect 2115 3073 2116 3077
rect 2110 3072 2116 3073
rect 2342 3077 2348 3078
rect 2342 3073 2343 3077
rect 2347 3073 2348 3077
rect 2342 3072 2348 3073
rect 2112 3059 2114 3072
rect 2174 3067 2180 3068
rect 2174 3063 2175 3067
rect 2179 3063 2180 3067
rect 2174 3062 2180 3063
rect 2071 3058 2075 3059
rect 1183 3054 1187 3055
rect 1183 3049 1187 3050
rect 1215 3054 1219 3055
rect 1215 3049 1219 3050
rect 1335 3054 1339 3055
rect 1335 3049 1339 3050
rect 1359 3054 1363 3055
rect 1359 3049 1363 3050
rect 1551 3054 1555 3055
rect 1551 3049 1555 3050
rect 1751 3054 1755 3055
rect 1751 3049 1755 3050
rect 1935 3054 1939 3055
rect 1935 3049 1939 3050
rect 2031 3054 2035 3055
rect 2071 3053 2075 3054
rect 2111 3058 2115 3059
rect 2111 3053 2115 3054
rect 2031 3049 2035 3050
rect 1166 3047 1172 3048
rect 1166 3043 1167 3047
rect 1171 3043 1172 3047
rect 1166 3042 1172 3043
rect 1216 3040 1218 3049
rect 1336 3040 1338 3049
rect 974 3039 980 3040
rect 974 3035 975 3039
rect 979 3035 980 3039
rect 974 3034 980 3035
rect 1094 3039 1100 3040
rect 1094 3035 1095 3039
rect 1099 3035 1100 3039
rect 1094 3034 1100 3035
rect 1214 3039 1220 3040
rect 1214 3035 1215 3039
rect 1219 3035 1220 3039
rect 1214 3034 1220 3035
rect 1334 3039 1340 3040
rect 1334 3035 1335 3039
rect 1339 3035 1340 3039
rect 1334 3034 1340 3035
rect 958 3031 964 3032
rect 662 3027 668 3028
rect 662 3023 663 3027
rect 667 3023 668 3027
rect 958 3027 959 3031
rect 963 3027 964 3031
rect 958 3026 964 3027
rect 1206 3027 1212 3028
rect 662 3022 668 3023
rect 1206 3023 1207 3027
rect 1211 3023 1212 3027
rect 1206 3022 1212 3023
rect 638 2998 644 2999
rect 638 2994 639 2998
rect 643 2994 644 2998
rect 638 2993 644 2994
rect 750 2998 756 2999
rect 750 2994 751 2998
rect 755 2994 756 2998
rect 750 2993 756 2994
rect 862 2998 868 2999
rect 862 2994 863 2998
rect 867 2994 868 2998
rect 862 2993 868 2994
rect 974 2998 980 2999
rect 974 2994 975 2998
rect 979 2994 980 2998
rect 974 2993 980 2994
rect 1094 2998 1100 2999
rect 1094 2994 1095 2998
rect 1099 2994 1100 2998
rect 1094 2993 1100 2994
rect 640 2975 642 2993
rect 752 2975 754 2993
rect 864 2975 866 2993
rect 976 2975 978 2993
rect 1096 2975 1098 2993
rect 607 2974 611 2975
rect 607 2969 611 2970
rect 639 2974 643 2975
rect 639 2969 643 2970
rect 751 2974 755 2975
rect 751 2969 755 2970
rect 783 2974 787 2975
rect 783 2969 787 2970
rect 863 2974 867 2975
rect 863 2969 867 2970
rect 959 2974 963 2975
rect 959 2969 963 2970
rect 975 2974 979 2975
rect 975 2969 979 2970
rect 1095 2974 1099 2975
rect 1095 2969 1099 2970
rect 1135 2974 1139 2975
rect 1135 2969 1139 2970
rect 608 2959 610 2969
rect 784 2959 786 2969
rect 960 2959 962 2969
rect 1136 2959 1138 2969
rect 606 2958 612 2959
rect 606 2954 607 2958
rect 611 2954 612 2958
rect 606 2953 612 2954
rect 782 2958 788 2959
rect 782 2954 783 2958
rect 787 2954 788 2958
rect 782 2953 788 2954
rect 958 2958 964 2959
rect 958 2954 959 2958
rect 963 2954 964 2958
rect 958 2953 964 2954
rect 1134 2958 1140 2959
rect 1134 2954 1135 2958
rect 1139 2954 1140 2958
rect 1134 2953 1140 2954
rect 230 2927 236 2928
rect 230 2923 231 2927
rect 235 2923 236 2927
rect 230 2922 236 2923
rect 598 2927 604 2928
rect 598 2923 599 2927
rect 603 2923 604 2927
rect 598 2922 604 2923
rect 982 2927 988 2928
rect 982 2923 983 2927
rect 987 2923 988 2927
rect 982 2922 988 2923
rect 150 2917 156 2918
rect 150 2913 151 2917
rect 155 2913 156 2917
rect 150 2912 156 2913
rect 152 2891 154 2912
rect 232 2900 234 2922
rect 270 2917 276 2918
rect 270 2913 271 2917
rect 275 2913 276 2917
rect 270 2912 276 2913
rect 430 2917 436 2918
rect 430 2913 431 2917
rect 435 2913 436 2917
rect 430 2912 436 2913
rect 606 2917 612 2918
rect 606 2913 607 2917
rect 611 2913 612 2917
rect 606 2912 612 2913
rect 782 2917 788 2918
rect 782 2913 783 2917
rect 787 2913 788 2917
rect 782 2912 788 2913
rect 958 2917 964 2918
rect 958 2913 959 2917
rect 963 2913 964 2917
rect 958 2912 964 2913
rect 230 2899 236 2900
rect 230 2895 231 2899
rect 235 2895 236 2899
rect 230 2894 236 2895
rect 272 2891 274 2912
rect 432 2891 434 2912
rect 514 2907 520 2908
rect 514 2903 515 2907
rect 519 2903 520 2907
rect 514 2902 520 2903
rect 111 2890 115 2891
rect 111 2885 115 2886
rect 151 2890 155 2891
rect 151 2885 155 2886
rect 271 2890 275 2891
rect 271 2885 275 2886
rect 287 2890 291 2891
rect 287 2885 291 2886
rect 431 2890 435 2891
rect 431 2885 435 2886
rect 447 2890 451 2891
rect 447 2885 451 2886
rect 112 2857 114 2885
rect 152 2876 154 2885
rect 222 2883 228 2884
rect 222 2879 223 2883
rect 227 2879 228 2883
rect 222 2878 228 2879
rect 150 2875 156 2876
rect 150 2871 151 2875
rect 155 2871 156 2875
rect 150 2870 156 2871
rect 110 2856 116 2857
rect 110 2852 111 2856
rect 115 2852 116 2856
rect 110 2851 116 2852
rect 110 2839 116 2840
rect 110 2835 111 2839
rect 115 2835 116 2839
rect 110 2834 116 2835
rect 150 2834 156 2835
rect 112 2807 114 2834
rect 150 2830 151 2834
rect 155 2830 156 2834
rect 150 2829 156 2830
rect 152 2807 154 2829
rect 111 2806 115 2807
rect 111 2801 115 2802
rect 151 2806 155 2807
rect 151 2801 155 2802
rect 112 2786 114 2801
rect 152 2791 154 2801
rect 150 2790 156 2791
rect 150 2786 151 2790
rect 155 2786 156 2790
rect 110 2785 116 2786
rect 150 2785 156 2786
rect 110 2781 111 2785
rect 115 2781 116 2785
rect 110 2780 116 2781
rect 110 2768 116 2769
rect 110 2764 111 2768
rect 115 2764 116 2768
rect 110 2763 116 2764
rect 112 2731 114 2763
rect 224 2760 226 2878
rect 288 2876 290 2885
rect 448 2876 450 2885
rect 286 2875 292 2876
rect 286 2871 287 2875
rect 291 2871 292 2875
rect 286 2870 292 2871
rect 446 2875 452 2876
rect 446 2871 447 2875
rect 451 2871 452 2875
rect 446 2870 452 2871
rect 516 2868 518 2902
rect 608 2891 610 2912
rect 784 2891 786 2912
rect 960 2891 962 2912
rect 599 2890 603 2891
rect 599 2885 603 2886
rect 607 2890 611 2891
rect 607 2885 611 2886
rect 759 2890 763 2891
rect 759 2885 763 2886
rect 783 2890 787 2891
rect 783 2885 787 2886
rect 927 2890 931 2891
rect 927 2885 931 2886
rect 959 2890 963 2891
rect 959 2885 963 2886
rect 600 2876 602 2885
rect 760 2876 762 2885
rect 928 2876 930 2885
rect 984 2884 986 2922
rect 1134 2917 1140 2918
rect 1134 2913 1135 2917
rect 1139 2913 1140 2917
rect 1134 2912 1140 2913
rect 1034 2907 1040 2908
rect 1034 2903 1035 2907
rect 1039 2903 1040 2907
rect 1034 2902 1040 2903
rect 1036 2884 1038 2902
rect 1136 2891 1138 2912
rect 1208 2908 1210 3022
rect 2032 3021 2034 3049
rect 2072 3025 2074 3053
rect 2112 3044 2114 3053
rect 2110 3043 2116 3044
rect 2110 3039 2111 3043
rect 2115 3039 2116 3043
rect 2110 3038 2116 3039
rect 2176 3036 2178 3062
rect 2344 3059 2346 3072
rect 2416 3068 2418 3186
rect 2550 3162 2556 3163
rect 2550 3158 2551 3162
rect 2555 3158 2556 3162
rect 2550 3157 2556 3158
rect 2694 3162 2700 3163
rect 2694 3158 2695 3162
rect 2699 3158 2700 3162
rect 2694 3157 2700 3158
rect 2838 3162 2844 3163
rect 2838 3158 2839 3162
rect 2843 3158 2844 3162
rect 2838 3157 2844 3158
rect 2974 3162 2980 3163
rect 2974 3158 2975 3162
rect 2979 3158 2980 3162
rect 2974 3157 2980 3158
rect 3110 3162 3116 3163
rect 3110 3158 3111 3162
rect 3115 3158 3116 3162
rect 3110 3157 3116 3158
rect 3246 3162 3252 3163
rect 3246 3158 3247 3162
rect 3251 3158 3252 3162
rect 3246 3157 3252 3158
rect 2552 3135 2554 3157
rect 2696 3135 2698 3157
rect 2840 3135 2842 3157
rect 2976 3135 2978 3157
rect 3112 3135 3114 3157
rect 3248 3135 3250 3157
rect 2551 3134 2555 3135
rect 2551 3129 2555 3130
rect 2583 3134 2587 3135
rect 2583 3129 2587 3130
rect 2695 3134 2699 3135
rect 2695 3129 2699 3130
rect 2799 3134 2803 3135
rect 2799 3129 2803 3130
rect 2839 3134 2843 3135
rect 2839 3129 2843 3130
rect 2975 3134 2979 3135
rect 2975 3129 2979 3130
rect 2999 3134 3003 3135
rect 2999 3129 3003 3130
rect 3111 3134 3115 3135
rect 3111 3129 3115 3130
rect 3191 3134 3195 3135
rect 3191 3129 3195 3130
rect 3247 3134 3251 3135
rect 3247 3129 3251 3130
rect 2584 3119 2586 3129
rect 2800 3119 2802 3129
rect 3000 3119 3002 3129
rect 3192 3119 3194 3129
rect 2582 3118 2588 3119
rect 2582 3114 2583 3118
rect 2587 3114 2588 3118
rect 2582 3113 2588 3114
rect 2798 3118 2804 3119
rect 2798 3114 2799 3118
rect 2803 3114 2804 3118
rect 2798 3113 2804 3114
rect 2998 3118 3004 3119
rect 2998 3114 2999 3118
rect 3003 3114 3004 3118
rect 2998 3113 3004 3114
rect 3190 3118 3196 3119
rect 3190 3114 3191 3118
rect 3195 3114 3196 3118
rect 3190 3113 3196 3114
rect 2566 3087 2572 3088
rect 2566 3083 2567 3087
rect 2571 3083 2572 3087
rect 2566 3082 2572 3083
rect 2662 3087 2668 3088
rect 2662 3083 2663 3087
rect 2667 3083 2668 3087
rect 2662 3082 2668 3083
rect 2982 3087 2988 3088
rect 2982 3083 2983 3087
rect 2987 3083 2988 3087
rect 2982 3082 2988 3083
rect 2568 3068 2570 3082
rect 2582 3077 2588 3078
rect 2582 3073 2583 3077
rect 2587 3073 2588 3077
rect 2582 3072 2588 3073
rect 2414 3067 2420 3068
rect 2414 3063 2415 3067
rect 2419 3063 2420 3067
rect 2414 3062 2420 3063
rect 2566 3067 2572 3068
rect 2566 3063 2567 3067
rect 2571 3063 2572 3067
rect 2566 3062 2572 3063
rect 2584 3059 2586 3072
rect 2263 3058 2267 3059
rect 2263 3053 2267 3054
rect 2343 3058 2347 3059
rect 2343 3053 2347 3054
rect 2455 3058 2459 3059
rect 2455 3053 2459 3054
rect 2583 3058 2587 3059
rect 2583 3053 2587 3054
rect 2655 3058 2659 3059
rect 2655 3053 2659 3054
rect 2264 3044 2266 3053
rect 2456 3044 2458 3053
rect 2526 3051 2532 3052
rect 2526 3047 2527 3051
rect 2531 3047 2532 3051
rect 2526 3046 2532 3047
rect 2262 3043 2268 3044
rect 2262 3039 2263 3043
rect 2267 3039 2268 3043
rect 2262 3038 2268 3039
rect 2454 3043 2460 3044
rect 2454 3039 2455 3043
rect 2459 3039 2460 3043
rect 2454 3038 2460 3039
rect 2174 3035 2180 3036
rect 2174 3031 2175 3035
rect 2179 3031 2180 3035
rect 2174 3030 2180 3031
rect 2070 3024 2076 3025
rect 2030 3020 2036 3021
rect 2030 3016 2031 3020
rect 2035 3016 2036 3020
rect 2070 3020 2071 3024
rect 2075 3020 2076 3024
rect 2070 3019 2076 3020
rect 2030 3015 2036 3016
rect 2070 3007 2076 3008
rect 2030 3003 2036 3004
rect 2030 2999 2031 3003
rect 2035 2999 2036 3003
rect 2070 3003 2071 3007
rect 2075 3003 2076 3007
rect 2070 3002 2076 3003
rect 2110 3002 2116 3003
rect 1214 2998 1220 2999
rect 1214 2994 1215 2998
rect 1219 2994 1220 2998
rect 1214 2993 1220 2994
rect 1334 2998 1340 2999
rect 2030 2998 2036 2999
rect 1334 2994 1335 2998
rect 1339 2994 1340 2998
rect 1334 2993 1340 2994
rect 1216 2975 1218 2993
rect 1336 2975 1338 2993
rect 2032 2975 2034 2998
rect 2072 2987 2074 3002
rect 2110 2998 2111 3002
rect 2115 2998 2116 3002
rect 2110 2997 2116 2998
rect 2262 3002 2268 3003
rect 2262 2998 2263 3002
rect 2267 2998 2268 3002
rect 2262 2997 2268 2998
rect 2454 3002 2460 3003
rect 2454 2998 2455 3002
rect 2459 2998 2460 3002
rect 2454 2997 2460 2998
rect 2112 2987 2114 2997
rect 2264 2987 2266 2997
rect 2338 2987 2344 2988
rect 2456 2987 2458 2997
rect 2528 2988 2530 3046
rect 2656 3044 2658 3053
rect 2664 3052 2666 3082
rect 2798 3077 2804 3078
rect 2798 3073 2799 3077
rect 2803 3073 2804 3077
rect 2798 3072 2804 3073
rect 2800 3059 2802 3072
rect 2984 3060 2986 3082
rect 2998 3077 3004 3078
rect 2998 3073 2999 3077
rect 3003 3073 3004 3077
rect 2998 3072 3004 3073
rect 3190 3077 3196 3078
rect 3190 3073 3191 3077
rect 3195 3073 3196 3077
rect 3190 3072 3196 3073
rect 2982 3059 2988 3060
rect 3000 3059 3002 3072
rect 3192 3059 3194 3072
rect 3264 3068 3266 3186
rect 3992 3185 3994 3213
rect 3990 3184 3996 3185
rect 3990 3180 3991 3184
rect 3995 3180 3996 3184
rect 3990 3179 3996 3180
rect 3990 3167 3996 3168
rect 3990 3163 3991 3167
rect 3995 3163 3996 3167
rect 3390 3162 3396 3163
rect 3990 3162 3996 3163
rect 3390 3158 3391 3162
rect 3395 3158 3396 3162
rect 3390 3157 3396 3158
rect 3392 3135 3394 3157
rect 3992 3135 3994 3162
rect 3375 3134 3379 3135
rect 3375 3129 3379 3130
rect 3391 3134 3395 3135
rect 3391 3129 3395 3130
rect 3567 3134 3571 3135
rect 3567 3129 3571 3130
rect 3991 3134 3995 3135
rect 3991 3129 3995 3130
rect 3376 3119 3378 3129
rect 3568 3119 3570 3129
rect 3374 3118 3380 3119
rect 3374 3114 3375 3118
rect 3379 3114 3380 3118
rect 3374 3113 3380 3114
rect 3566 3118 3572 3119
rect 3566 3114 3567 3118
rect 3571 3114 3572 3118
rect 3992 3114 3994 3129
rect 3566 3113 3572 3114
rect 3990 3113 3996 3114
rect 3990 3109 3991 3113
rect 3995 3109 3996 3113
rect 3990 3108 3996 3109
rect 3990 3096 3996 3097
rect 3990 3092 3991 3096
rect 3995 3092 3996 3096
rect 3990 3091 3996 3092
rect 3550 3087 3556 3088
rect 3550 3083 3551 3087
rect 3555 3083 3556 3087
rect 3550 3082 3556 3083
rect 3662 3087 3668 3088
rect 3662 3083 3663 3087
rect 3667 3083 3668 3087
rect 3662 3082 3668 3083
rect 3374 3077 3380 3078
rect 3374 3073 3375 3077
rect 3379 3073 3380 3077
rect 3374 3072 3380 3073
rect 3262 3067 3268 3068
rect 3262 3063 3263 3067
rect 3267 3063 3268 3067
rect 3262 3062 3268 3063
rect 3376 3059 3378 3072
rect 3552 3068 3554 3082
rect 3566 3077 3572 3078
rect 3566 3073 3567 3077
rect 3571 3073 3572 3077
rect 3566 3072 3572 3073
rect 3550 3067 3556 3068
rect 3550 3063 3551 3067
rect 3555 3063 3556 3067
rect 3550 3062 3556 3063
rect 3568 3059 3570 3072
rect 2799 3058 2803 3059
rect 2799 3053 2803 3054
rect 2855 3058 2859 3059
rect 2982 3055 2983 3059
rect 2987 3055 2988 3059
rect 2982 3054 2988 3055
rect 2999 3058 3003 3059
rect 2855 3053 2859 3054
rect 2999 3053 3003 3054
rect 3055 3058 3059 3059
rect 3055 3053 3059 3054
rect 3191 3058 3195 3059
rect 3191 3053 3195 3054
rect 3255 3058 3259 3059
rect 3255 3053 3259 3054
rect 3375 3058 3379 3059
rect 3375 3053 3379 3054
rect 3455 3058 3459 3059
rect 3455 3053 3459 3054
rect 3567 3058 3571 3059
rect 3567 3053 3571 3054
rect 3655 3058 3659 3059
rect 3655 3053 3659 3054
rect 2662 3051 2668 3052
rect 2662 3047 2663 3051
rect 2667 3047 2668 3051
rect 2662 3046 2668 3047
rect 2856 3044 2858 3053
rect 3056 3044 3058 3053
rect 3256 3044 3258 3053
rect 3456 3044 3458 3053
rect 3656 3044 3658 3053
rect 3664 3052 3666 3082
rect 3992 3059 3994 3091
rect 3991 3058 3995 3059
rect 3991 3053 3995 3054
rect 3662 3051 3668 3052
rect 3662 3047 3663 3051
rect 3667 3047 3668 3051
rect 3662 3046 3668 3047
rect 2654 3043 2660 3044
rect 2654 3039 2655 3043
rect 2659 3039 2660 3043
rect 2654 3038 2660 3039
rect 2854 3043 2860 3044
rect 2854 3039 2855 3043
rect 2859 3039 2860 3043
rect 2854 3038 2860 3039
rect 3054 3043 3060 3044
rect 3054 3039 3055 3043
rect 3059 3039 3060 3043
rect 3054 3038 3060 3039
rect 3254 3043 3260 3044
rect 3254 3039 3255 3043
rect 3259 3039 3260 3043
rect 3254 3038 3260 3039
rect 3454 3043 3460 3044
rect 3454 3039 3455 3043
rect 3459 3039 3460 3043
rect 3454 3038 3460 3039
rect 3654 3043 3660 3044
rect 3654 3039 3655 3043
rect 3659 3039 3660 3043
rect 3654 3038 3660 3039
rect 2918 3035 2924 3036
rect 2918 3031 2919 3035
rect 2923 3031 2924 3035
rect 2918 3030 2924 3031
rect 3150 3035 3156 3036
rect 3150 3031 3151 3035
rect 3155 3031 3156 3035
rect 3150 3030 3156 3031
rect 2654 3002 2660 3003
rect 2654 2998 2655 3002
rect 2659 2998 2660 3002
rect 2654 2997 2660 2998
rect 2854 3002 2860 3003
rect 2854 2998 2855 3002
rect 2859 2998 2860 3002
rect 2854 2997 2860 2998
rect 2526 2987 2532 2988
rect 2656 2987 2658 2997
rect 2856 2987 2858 2997
rect 2071 2986 2075 2987
rect 2071 2981 2075 2982
rect 2111 2986 2115 2987
rect 2111 2981 2115 2982
rect 2263 2986 2267 2987
rect 2338 2983 2339 2987
rect 2343 2983 2344 2987
rect 2338 2982 2344 2983
rect 2359 2986 2363 2987
rect 2263 2981 2267 2982
rect 1215 2974 1219 2975
rect 1215 2969 1219 2970
rect 1303 2974 1307 2975
rect 1303 2969 1307 2970
rect 1335 2974 1339 2975
rect 1335 2969 1339 2970
rect 1471 2974 1475 2975
rect 1471 2969 1475 2970
rect 1647 2974 1651 2975
rect 1647 2969 1651 2970
rect 2031 2974 2035 2975
rect 2031 2969 2035 2970
rect 1304 2959 1306 2969
rect 1472 2959 1474 2969
rect 1648 2959 1650 2969
rect 1302 2958 1308 2959
rect 1302 2954 1303 2958
rect 1307 2954 1308 2958
rect 1302 2953 1308 2954
rect 1470 2958 1476 2959
rect 1470 2954 1471 2958
rect 1475 2954 1476 2958
rect 1470 2953 1476 2954
rect 1646 2958 1652 2959
rect 1646 2954 1647 2958
rect 1651 2954 1652 2958
rect 2032 2954 2034 2969
rect 2072 2966 2074 2981
rect 2112 2971 2114 2981
rect 2110 2970 2116 2971
rect 2110 2966 2111 2970
rect 2115 2966 2116 2970
rect 2070 2965 2076 2966
rect 2110 2965 2116 2966
rect 2070 2961 2071 2965
rect 2075 2961 2076 2965
rect 2070 2960 2076 2961
rect 1646 2953 1652 2954
rect 2030 2953 2036 2954
rect 2030 2949 2031 2953
rect 2035 2949 2036 2953
rect 2030 2948 2036 2949
rect 2070 2948 2076 2949
rect 2070 2944 2071 2948
rect 2075 2944 2076 2948
rect 2070 2943 2076 2944
rect 2030 2936 2036 2937
rect 2030 2932 2031 2936
rect 2035 2932 2036 2936
rect 2030 2931 2036 2932
rect 1266 2927 1272 2928
rect 1266 2923 1267 2927
rect 1271 2923 1272 2927
rect 1266 2922 1272 2923
rect 1454 2927 1460 2928
rect 1454 2923 1455 2927
rect 1459 2923 1460 2927
rect 1454 2922 1460 2923
rect 1630 2927 1636 2928
rect 1630 2923 1631 2927
rect 1635 2923 1636 2927
rect 1630 2922 1636 2923
rect 1718 2927 1724 2928
rect 1718 2923 1719 2927
rect 1723 2923 1724 2927
rect 1718 2922 1724 2923
rect 1268 2908 1270 2922
rect 1302 2917 1308 2918
rect 1302 2913 1303 2917
rect 1307 2913 1308 2917
rect 1302 2912 1308 2913
rect 1206 2907 1212 2908
rect 1206 2903 1207 2907
rect 1211 2903 1212 2907
rect 1206 2902 1212 2903
rect 1266 2907 1272 2908
rect 1266 2903 1267 2907
rect 1271 2903 1272 2907
rect 1266 2902 1272 2903
rect 1304 2891 1306 2912
rect 1456 2908 1458 2922
rect 1470 2917 1476 2918
rect 1470 2913 1471 2917
rect 1475 2913 1476 2917
rect 1470 2912 1476 2913
rect 1454 2907 1460 2908
rect 1454 2903 1455 2907
rect 1459 2903 1460 2907
rect 1454 2902 1460 2903
rect 1472 2891 1474 2912
rect 1632 2908 1634 2922
rect 1646 2917 1652 2918
rect 1646 2913 1647 2917
rect 1651 2913 1652 2917
rect 1646 2912 1652 2913
rect 1630 2907 1636 2908
rect 1630 2903 1631 2907
rect 1635 2903 1636 2907
rect 1630 2902 1636 2903
rect 1648 2891 1650 2912
rect 1103 2890 1107 2891
rect 1103 2885 1107 2886
rect 1135 2890 1139 2891
rect 1135 2885 1139 2886
rect 1287 2890 1291 2891
rect 1287 2885 1291 2886
rect 1303 2890 1307 2891
rect 1303 2885 1307 2886
rect 1471 2890 1475 2891
rect 1471 2885 1475 2886
rect 1479 2890 1483 2891
rect 1479 2885 1483 2886
rect 1647 2890 1651 2891
rect 1647 2885 1651 2886
rect 1671 2890 1675 2891
rect 1671 2885 1675 2886
rect 982 2883 988 2884
rect 982 2879 983 2883
rect 987 2879 988 2883
rect 982 2878 988 2879
rect 1034 2883 1040 2884
rect 1034 2879 1035 2883
rect 1039 2879 1040 2883
rect 1034 2878 1040 2879
rect 1104 2876 1106 2885
rect 1288 2876 1290 2885
rect 1480 2876 1482 2885
rect 1534 2883 1540 2884
rect 1534 2879 1535 2883
rect 1539 2879 1540 2883
rect 1534 2878 1540 2879
rect 598 2875 604 2876
rect 598 2871 599 2875
rect 603 2871 604 2875
rect 598 2870 604 2871
rect 758 2875 764 2876
rect 758 2871 759 2875
rect 763 2871 764 2875
rect 758 2870 764 2871
rect 926 2875 932 2876
rect 926 2871 927 2875
rect 931 2871 932 2875
rect 926 2870 932 2871
rect 1102 2875 1108 2876
rect 1102 2871 1103 2875
rect 1107 2871 1108 2875
rect 1102 2870 1108 2871
rect 1286 2875 1292 2876
rect 1286 2871 1287 2875
rect 1291 2871 1292 2875
rect 1286 2870 1292 2871
rect 1478 2875 1484 2876
rect 1478 2871 1479 2875
rect 1483 2871 1484 2875
rect 1478 2870 1484 2871
rect 514 2867 520 2868
rect 514 2863 515 2867
rect 519 2863 520 2867
rect 514 2862 520 2863
rect 590 2863 596 2864
rect 590 2859 591 2863
rect 595 2859 596 2863
rect 590 2858 596 2859
rect 286 2834 292 2835
rect 286 2830 287 2834
rect 291 2830 292 2834
rect 286 2829 292 2830
rect 446 2834 452 2835
rect 446 2830 447 2834
rect 451 2830 452 2834
rect 446 2829 452 2830
rect 288 2807 290 2829
rect 448 2807 450 2829
rect 287 2806 291 2807
rect 287 2801 291 2802
rect 319 2806 323 2807
rect 319 2801 323 2802
rect 447 2806 451 2807
rect 447 2801 451 2802
rect 503 2806 507 2807
rect 503 2801 507 2802
rect 320 2791 322 2801
rect 504 2791 506 2801
rect 318 2790 324 2791
rect 318 2786 319 2790
rect 323 2786 324 2790
rect 318 2785 324 2786
rect 502 2790 508 2791
rect 502 2786 503 2790
rect 507 2786 508 2790
rect 502 2785 508 2786
rect 222 2759 228 2760
rect 222 2755 223 2759
rect 227 2755 228 2759
rect 222 2754 228 2755
rect 150 2749 156 2750
rect 150 2745 151 2749
rect 155 2745 156 2749
rect 150 2744 156 2745
rect 318 2749 324 2750
rect 318 2745 319 2749
rect 323 2745 324 2749
rect 318 2744 324 2745
rect 502 2749 508 2750
rect 502 2745 503 2749
rect 507 2745 508 2749
rect 502 2744 508 2745
rect 152 2731 154 2744
rect 320 2731 322 2744
rect 390 2739 396 2740
rect 390 2735 391 2739
rect 395 2735 396 2739
rect 390 2734 396 2735
rect 111 2730 115 2731
rect 111 2725 115 2726
rect 151 2730 155 2731
rect 151 2725 155 2726
rect 183 2730 187 2731
rect 183 2725 187 2726
rect 319 2730 323 2731
rect 319 2725 323 2726
rect 383 2730 387 2731
rect 383 2725 387 2726
rect 112 2697 114 2725
rect 184 2716 186 2725
rect 246 2723 252 2724
rect 246 2719 247 2723
rect 251 2719 252 2723
rect 246 2718 252 2719
rect 182 2715 188 2716
rect 182 2711 183 2715
rect 187 2711 188 2715
rect 182 2710 188 2711
rect 110 2696 116 2697
rect 110 2692 111 2696
rect 115 2692 116 2696
rect 110 2691 116 2692
rect 110 2679 116 2680
rect 110 2675 111 2679
rect 115 2675 116 2679
rect 110 2674 116 2675
rect 182 2674 188 2675
rect 112 2651 114 2674
rect 182 2670 183 2674
rect 187 2670 188 2674
rect 182 2669 188 2670
rect 184 2651 186 2669
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 183 2650 187 2651
rect 183 2645 187 2646
rect 112 2630 114 2645
rect 110 2629 116 2630
rect 110 2625 111 2629
rect 115 2625 116 2629
rect 110 2624 116 2625
rect 110 2612 116 2613
rect 110 2608 111 2612
rect 115 2608 116 2612
rect 110 2607 116 2608
rect 112 2575 114 2607
rect 248 2604 250 2718
rect 384 2716 386 2725
rect 382 2715 388 2716
rect 382 2711 383 2715
rect 387 2711 388 2715
rect 382 2710 388 2711
rect 392 2704 394 2734
rect 504 2731 506 2744
rect 592 2740 594 2858
rect 598 2834 604 2835
rect 598 2830 599 2834
rect 603 2830 604 2834
rect 598 2829 604 2830
rect 758 2834 764 2835
rect 758 2830 759 2834
rect 763 2830 764 2834
rect 758 2829 764 2830
rect 926 2834 932 2835
rect 926 2830 927 2834
rect 931 2830 932 2834
rect 926 2829 932 2830
rect 1102 2834 1108 2835
rect 1102 2830 1103 2834
rect 1107 2830 1108 2834
rect 1102 2829 1108 2830
rect 1286 2834 1292 2835
rect 1286 2830 1287 2834
rect 1291 2830 1292 2834
rect 1286 2829 1292 2830
rect 1478 2834 1484 2835
rect 1478 2830 1479 2834
rect 1483 2830 1484 2834
rect 1478 2829 1484 2830
rect 600 2807 602 2829
rect 760 2807 762 2829
rect 928 2807 930 2829
rect 1104 2807 1106 2829
rect 1288 2807 1290 2829
rect 1480 2807 1482 2829
rect 599 2806 603 2807
rect 599 2801 603 2802
rect 687 2806 691 2807
rect 687 2801 691 2802
rect 759 2806 763 2807
rect 759 2801 763 2802
rect 871 2806 875 2807
rect 871 2801 875 2802
rect 927 2806 931 2807
rect 927 2801 931 2802
rect 1055 2806 1059 2807
rect 1055 2801 1059 2802
rect 1103 2806 1107 2807
rect 1103 2801 1107 2802
rect 1239 2806 1243 2807
rect 1239 2801 1243 2802
rect 1287 2806 1291 2807
rect 1287 2801 1291 2802
rect 1431 2806 1435 2807
rect 1431 2801 1435 2802
rect 1479 2806 1483 2807
rect 1479 2801 1483 2802
rect 688 2791 690 2801
rect 872 2791 874 2801
rect 1056 2791 1058 2801
rect 1240 2791 1242 2801
rect 1432 2791 1434 2801
rect 686 2790 692 2791
rect 686 2786 687 2790
rect 691 2786 692 2790
rect 686 2785 692 2786
rect 870 2790 876 2791
rect 870 2786 871 2790
rect 875 2786 876 2790
rect 870 2785 876 2786
rect 1054 2790 1060 2791
rect 1054 2786 1055 2790
rect 1059 2786 1060 2790
rect 1054 2785 1060 2786
rect 1238 2790 1244 2791
rect 1238 2786 1239 2790
rect 1243 2786 1244 2790
rect 1238 2785 1244 2786
rect 1430 2790 1436 2791
rect 1430 2786 1431 2790
rect 1435 2786 1436 2790
rect 1430 2785 1436 2786
rect 1536 2760 1538 2878
rect 1672 2876 1674 2885
rect 1720 2884 1722 2922
rect 2032 2891 2034 2931
rect 2072 2907 2074 2943
rect 2340 2940 2342 2982
rect 2359 2981 2363 2982
rect 2455 2986 2459 2987
rect 2526 2983 2527 2987
rect 2531 2983 2532 2987
rect 2526 2982 2532 2983
rect 2607 2986 2611 2987
rect 2455 2981 2459 2982
rect 2607 2981 2611 2982
rect 2655 2986 2659 2987
rect 2655 2981 2659 2982
rect 2847 2986 2851 2987
rect 2847 2981 2851 2982
rect 2855 2986 2859 2987
rect 2855 2981 2859 2982
rect 2360 2971 2362 2981
rect 2608 2971 2610 2981
rect 2848 2971 2850 2981
rect 2358 2970 2364 2971
rect 2358 2966 2359 2970
rect 2363 2966 2364 2970
rect 2358 2965 2364 2966
rect 2606 2970 2612 2971
rect 2606 2966 2607 2970
rect 2611 2966 2612 2970
rect 2606 2965 2612 2966
rect 2846 2970 2852 2971
rect 2846 2966 2847 2970
rect 2851 2966 2852 2970
rect 2846 2965 2852 2966
rect 2338 2939 2344 2940
rect 2338 2935 2339 2939
rect 2343 2935 2344 2939
rect 2338 2934 2344 2935
rect 2110 2929 2116 2930
rect 2110 2925 2111 2929
rect 2115 2925 2116 2929
rect 2110 2924 2116 2925
rect 2358 2929 2364 2930
rect 2358 2925 2359 2929
rect 2363 2925 2364 2929
rect 2606 2929 2612 2930
rect 2358 2924 2364 2925
rect 2422 2927 2428 2928
rect 2112 2907 2114 2924
rect 2360 2907 2362 2924
rect 2422 2923 2423 2927
rect 2427 2923 2428 2927
rect 2606 2925 2607 2929
rect 2611 2925 2612 2929
rect 2606 2924 2612 2925
rect 2846 2929 2852 2930
rect 2846 2925 2847 2929
rect 2851 2925 2852 2929
rect 2846 2924 2852 2925
rect 2422 2922 2428 2923
rect 2071 2906 2075 2907
rect 2071 2901 2075 2902
rect 2111 2906 2115 2907
rect 2111 2901 2115 2902
rect 2279 2906 2283 2907
rect 2279 2901 2283 2902
rect 2359 2906 2363 2907
rect 2359 2901 2363 2902
rect 2031 2890 2035 2891
rect 2031 2885 2035 2886
rect 1718 2883 1724 2884
rect 1718 2879 1719 2883
rect 1723 2879 1724 2883
rect 1718 2878 1724 2879
rect 1670 2875 1676 2876
rect 1670 2871 1671 2875
rect 1675 2871 1676 2875
rect 1670 2870 1676 2871
rect 1694 2863 1700 2864
rect 1694 2859 1695 2863
rect 1699 2859 1700 2863
rect 1694 2858 1700 2859
rect 1670 2834 1676 2835
rect 1670 2830 1671 2834
rect 1675 2830 1676 2834
rect 1670 2829 1676 2830
rect 1672 2807 1674 2829
rect 1631 2806 1635 2807
rect 1631 2801 1635 2802
rect 1671 2806 1675 2807
rect 1671 2801 1675 2802
rect 1632 2791 1634 2801
rect 1630 2790 1636 2791
rect 1630 2786 1631 2790
rect 1635 2786 1636 2790
rect 1630 2785 1636 2786
rect 670 2759 676 2760
rect 670 2755 671 2759
rect 675 2755 676 2759
rect 670 2754 676 2755
rect 1222 2759 1228 2760
rect 1222 2755 1223 2759
rect 1227 2755 1228 2759
rect 1222 2754 1228 2755
rect 1414 2759 1420 2760
rect 1414 2755 1415 2759
rect 1419 2755 1420 2759
rect 1414 2754 1420 2755
rect 1534 2759 1540 2760
rect 1534 2755 1535 2759
rect 1539 2755 1540 2759
rect 1534 2754 1540 2755
rect 672 2740 674 2754
rect 686 2749 692 2750
rect 686 2745 687 2749
rect 691 2745 692 2749
rect 686 2744 692 2745
rect 870 2749 876 2750
rect 870 2745 871 2749
rect 875 2745 876 2749
rect 870 2744 876 2745
rect 1054 2749 1060 2750
rect 1054 2745 1055 2749
rect 1059 2745 1060 2749
rect 1054 2744 1060 2745
rect 590 2739 596 2740
rect 590 2735 591 2739
rect 595 2735 596 2739
rect 590 2734 596 2735
rect 670 2739 676 2740
rect 670 2735 671 2739
rect 675 2735 676 2739
rect 670 2734 676 2735
rect 688 2731 690 2744
rect 872 2731 874 2744
rect 1046 2739 1052 2740
rect 1046 2735 1047 2739
rect 1051 2735 1052 2739
rect 1046 2734 1052 2735
rect 503 2730 507 2731
rect 503 2725 507 2726
rect 583 2730 587 2731
rect 583 2725 587 2726
rect 687 2730 691 2731
rect 687 2725 691 2726
rect 783 2730 787 2731
rect 783 2725 787 2726
rect 871 2730 875 2731
rect 871 2725 875 2726
rect 983 2730 987 2731
rect 983 2725 987 2726
rect 584 2716 586 2725
rect 784 2716 786 2725
rect 984 2716 986 2725
rect 582 2715 588 2716
rect 582 2711 583 2715
rect 587 2711 588 2715
rect 582 2710 588 2711
rect 782 2715 788 2716
rect 782 2711 783 2715
rect 787 2711 788 2715
rect 782 2710 788 2711
rect 982 2715 988 2716
rect 982 2711 983 2715
rect 987 2711 988 2715
rect 982 2710 988 2711
rect 1048 2708 1050 2734
rect 1056 2731 1058 2744
rect 1224 2740 1226 2754
rect 1238 2749 1244 2750
rect 1238 2745 1239 2749
rect 1243 2745 1244 2749
rect 1238 2744 1244 2745
rect 1222 2739 1228 2740
rect 1222 2735 1223 2739
rect 1227 2735 1228 2739
rect 1222 2734 1228 2735
rect 1240 2731 1242 2744
rect 1416 2740 1418 2754
rect 1430 2749 1436 2750
rect 1430 2745 1431 2749
rect 1435 2745 1436 2749
rect 1430 2744 1436 2745
rect 1630 2749 1636 2750
rect 1630 2745 1631 2749
rect 1635 2745 1636 2749
rect 1630 2744 1636 2745
rect 1414 2739 1420 2740
rect 1414 2735 1415 2739
rect 1419 2735 1420 2739
rect 1414 2734 1420 2735
rect 1432 2731 1434 2744
rect 1632 2731 1634 2744
rect 1696 2740 1698 2858
rect 2032 2857 2034 2885
rect 2072 2873 2074 2901
rect 2112 2892 2114 2901
rect 2280 2892 2282 2901
rect 2424 2900 2426 2922
rect 2434 2919 2440 2920
rect 2434 2915 2435 2919
rect 2439 2915 2440 2919
rect 2434 2914 2440 2915
rect 2436 2900 2438 2914
rect 2608 2907 2610 2924
rect 2848 2907 2850 2924
rect 2920 2920 2922 3030
rect 3054 3002 3060 3003
rect 3054 2998 3055 3002
rect 3059 2998 3060 3002
rect 3054 2997 3060 2998
rect 3056 2987 3058 2997
rect 3055 2986 3059 2987
rect 3055 2981 3059 2982
rect 3079 2986 3083 2987
rect 3079 2981 3083 2982
rect 3080 2971 3082 2981
rect 3078 2970 3084 2971
rect 3078 2966 3079 2970
rect 3083 2966 3084 2970
rect 3078 2965 3084 2966
rect 3078 2929 3084 2930
rect 3078 2925 3079 2929
rect 3083 2925 3084 2929
rect 3078 2924 3084 2925
rect 2918 2919 2924 2920
rect 2918 2915 2919 2919
rect 2923 2915 2924 2919
rect 2918 2914 2924 2915
rect 3080 2907 3082 2924
rect 3152 2920 3154 3030
rect 3992 3025 3994 3053
rect 3990 3024 3996 3025
rect 3990 3020 3991 3024
rect 3995 3020 3996 3024
rect 3990 3019 3996 3020
rect 3990 3007 3996 3008
rect 3990 3003 3991 3007
rect 3995 3003 3996 3007
rect 3254 3002 3260 3003
rect 3254 2998 3255 3002
rect 3259 2998 3260 3002
rect 3254 2997 3260 2998
rect 3454 3002 3460 3003
rect 3454 2998 3455 3002
rect 3459 2998 3460 3002
rect 3454 2997 3460 2998
rect 3654 3002 3660 3003
rect 3990 3002 3996 3003
rect 3654 2998 3655 3002
rect 3659 2998 3660 3002
rect 3654 2997 3660 2998
rect 3256 2987 3258 2997
rect 3456 2987 3458 2997
rect 3656 2987 3658 2997
rect 3992 2987 3994 3002
rect 3255 2986 3259 2987
rect 3255 2981 3259 2982
rect 3303 2986 3307 2987
rect 3303 2981 3307 2982
rect 3455 2986 3459 2987
rect 3455 2981 3459 2982
rect 3535 2986 3539 2987
rect 3535 2981 3539 2982
rect 3655 2986 3659 2987
rect 3655 2981 3659 2982
rect 3767 2986 3771 2987
rect 3767 2981 3771 2982
rect 3991 2986 3995 2987
rect 3991 2981 3995 2982
rect 3304 2971 3306 2981
rect 3536 2971 3538 2981
rect 3768 2971 3770 2981
rect 3302 2970 3308 2971
rect 3302 2966 3303 2970
rect 3307 2966 3308 2970
rect 3302 2965 3308 2966
rect 3534 2970 3540 2971
rect 3534 2966 3535 2970
rect 3539 2966 3540 2970
rect 3534 2965 3540 2966
rect 3766 2970 3772 2971
rect 3766 2966 3767 2970
rect 3771 2966 3772 2970
rect 3992 2966 3994 2981
rect 3766 2965 3772 2966
rect 3990 2965 3996 2966
rect 3990 2961 3991 2965
rect 3995 2961 3996 2965
rect 3990 2960 3996 2961
rect 3990 2948 3996 2949
rect 3990 2944 3991 2948
rect 3995 2944 3996 2948
rect 3990 2943 3996 2944
rect 3286 2939 3292 2940
rect 3286 2935 3287 2939
rect 3291 2935 3292 2939
rect 3286 2934 3292 2935
rect 3518 2939 3524 2940
rect 3518 2935 3519 2939
rect 3523 2935 3524 2939
rect 3518 2934 3524 2935
rect 3750 2939 3756 2940
rect 3750 2935 3751 2939
rect 3755 2935 3756 2939
rect 3750 2934 3756 2935
rect 3288 2920 3290 2934
rect 3302 2929 3308 2930
rect 3302 2925 3303 2929
rect 3307 2925 3308 2929
rect 3302 2924 3308 2925
rect 3150 2919 3156 2920
rect 3150 2915 3151 2919
rect 3155 2915 3156 2919
rect 3150 2914 3156 2915
rect 3286 2919 3292 2920
rect 3286 2915 3287 2919
rect 3291 2915 3292 2919
rect 3286 2914 3292 2915
rect 3304 2907 3306 2924
rect 3520 2920 3522 2934
rect 3534 2929 3540 2930
rect 3534 2925 3535 2929
rect 3539 2925 3540 2929
rect 3534 2924 3540 2925
rect 3518 2919 3524 2920
rect 3518 2915 3519 2919
rect 3523 2915 3524 2919
rect 3518 2914 3524 2915
rect 3536 2907 3538 2924
rect 3752 2920 3754 2934
rect 3766 2929 3772 2930
rect 3766 2925 3767 2929
rect 3771 2925 3772 2929
rect 3766 2924 3772 2925
rect 3750 2919 3756 2920
rect 3750 2915 3751 2919
rect 3755 2915 3756 2919
rect 3750 2914 3756 2915
rect 3768 2907 3770 2924
rect 3992 2907 3994 2943
rect 2487 2906 2491 2907
rect 2487 2901 2491 2902
rect 2607 2906 2611 2907
rect 2607 2901 2611 2902
rect 2695 2906 2699 2907
rect 2695 2901 2699 2902
rect 2847 2906 2851 2907
rect 2847 2901 2851 2902
rect 2903 2906 2907 2907
rect 2903 2901 2907 2902
rect 3079 2906 3083 2907
rect 3079 2901 3083 2902
rect 3111 2906 3115 2907
rect 3111 2901 3115 2902
rect 3303 2906 3307 2907
rect 3303 2901 3307 2902
rect 3495 2906 3499 2907
rect 3495 2901 3499 2902
rect 3535 2906 3539 2907
rect 3535 2901 3539 2902
rect 3687 2906 3691 2907
rect 3687 2901 3691 2902
rect 3767 2906 3771 2907
rect 3767 2901 3771 2902
rect 3879 2906 3883 2907
rect 3879 2901 3883 2902
rect 3991 2906 3995 2907
rect 3991 2901 3995 2902
rect 2422 2899 2428 2900
rect 2422 2895 2423 2899
rect 2427 2895 2428 2899
rect 2422 2894 2428 2895
rect 2434 2899 2440 2900
rect 2434 2895 2435 2899
rect 2439 2895 2440 2899
rect 2434 2894 2440 2895
rect 2488 2892 2490 2901
rect 2696 2892 2698 2901
rect 2904 2892 2906 2901
rect 2974 2899 2980 2900
rect 2974 2895 2975 2899
rect 2979 2895 2980 2899
rect 2974 2894 2980 2895
rect 2110 2891 2116 2892
rect 2110 2887 2111 2891
rect 2115 2887 2116 2891
rect 2110 2886 2116 2887
rect 2278 2891 2284 2892
rect 2278 2887 2279 2891
rect 2283 2887 2284 2891
rect 2278 2886 2284 2887
rect 2486 2891 2492 2892
rect 2486 2887 2487 2891
rect 2491 2887 2492 2891
rect 2486 2886 2492 2887
rect 2694 2891 2700 2892
rect 2694 2887 2695 2891
rect 2699 2887 2700 2891
rect 2694 2886 2700 2887
rect 2902 2891 2908 2892
rect 2902 2887 2903 2891
rect 2907 2887 2908 2891
rect 2902 2886 2908 2887
rect 2230 2883 2236 2884
rect 2230 2879 2231 2883
rect 2235 2879 2236 2883
rect 2230 2878 2236 2879
rect 2070 2872 2076 2873
rect 2070 2868 2071 2872
rect 2075 2868 2076 2872
rect 2070 2867 2076 2868
rect 2030 2856 2036 2857
rect 2030 2852 2031 2856
rect 2035 2852 2036 2856
rect 2030 2851 2036 2852
rect 2070 2855 2076 2856
rect 2070 2851 2071 2855
rect 2075 2851 2076 2855
rect 2070 2850 2076 2851
rect 2110 2850 2116 2851
rect 2030 2839 2036 2840
rect 2030 2835 2031 2839
rect 2035 2835 2036 2839
rect 2030 2834 2036 2835
rect 2032 2807 2034 2834
rect 2072 2823 2074 2850
rect 2110 2846 2111 2850
rect 2115 2846 2116 2850
rect 2110 2845 2116 2846
rect 2112 2823 2114 2845
rect 2071 2822 2075 2823
rect 2071 2817 2075 2818
rect 2111 2822 2115 2823
rect 2111 2817 2115 2818
rect 2143 2822 2147 2823
rect 2143 2817 2147 2818
rect 1831 2806 1835 2807
rect 1831 2801 1835 2802
rect 2031 2806 2035 2807
rect 2072 2802 2074 2817
rect 2144 2807 2146 2817
rect 2142 2806 2148 2807
rect 2142 2802 2143 2806
rect 2147 2802 2148 2806
rect 2031 2801 2035 2802
rect 2070 2801 2076 2802
rect 2142 2801 2148 2802
rect 1832 2791 1834 2801
rect 1830 2790 1836 2791
rect 1830 2786 1831 2790
rect 1835 2786 1836 2790
rect 2032 2786 2034 2801
rect 2070 2797 2071 2801
rect 2075 2797 2076 2801
rect 2070 2796 2076 2797
rect 1830 2785 1836 2786
rect 2030 2785 2036 2786
rect 2030 2781 2031 2785
rect 2035 2781 2036 2785
rect 2030 2780 2036 2781
rect 2070 2784 2076 2785
rect 2070 2780 2071 2784
rect 2075 2780 2076 2784
rect 2070 2779 2076 2780
rect 2030 2768 2036 2769
rect 2030 2764 2031 2768
rect 2035 2764 2036 2768
rect 2030 2763 2036 2764
rect 1814 2759 1820 2760
rect 1814 2755 1815 2759
rect 1819 2755 1820 2759
rect 1814 2754 1820 2755
rect 1902 2759 1908 2760
rect 1902 2755 1903 2759
rect 1907 2755 1908 2759
rect 1902 2754 1908 2755
rect 1816 2740 1818 2754
rect 1830 2749 1836 2750
rect 1830 2745 1831 2749
rect 1835 2745 1836 2749
rect 1830 2744 1836 2745
rect 1694 2739 1700 2740
rect 1694 2735 1695 2739
rect 1699 2735 1700 2739
rect 1694 2734 1700 2735
rect 1814 2739 1820 2740
rect 1814 2735 1815 2739
rect 1819 2735 1820 2739
rect 1814 2734 1820 2735
rect 1832 2731 1834 2744
rect 1055 2730 1059 2731
rect 1055 2725 1059 2726
rect 1199 2730 1203 2731
rect 1199 2725 1203 2726
rect 1239 2730 1243 2731
rect 1239 2725 1243 2726
rect 1415 2730 1419 2731
rect 1415 2725 1419 2726
rect 1431 2730 1435 2731
rect 1431 2725 1435 2726
rect 1631 2730 1635 2731
rect 1631 2725 1635 2726
rect 1639 2730 1643 2731
rect 1639 2725 1643 2726
rect 1831 2730 1835 2731
rect 1831 2725 1835 2726
rect 1871 2730 1875 2731
rect 1871 2725 1875 2726
rect 1200 2716 1202 2725
rect 1416 2716 1418 2725
rect 1640 2716 1642 2725
rect 1646 2723 1652 2724
rect 1646 2719 1647 2723
rect 1651 2719 1652 2723
rect 1646 2718 1652 2719
rect 1198 2715 1204 2716
rect 1198 2711 1199 2715
rect 1203 2711 1204 2715
rect 1198 2710 1204 2711
rect 1414 2715 1420 2716
rect 1414 2711 1415 2715
rect 1419 2711 1420 2715
rect 1414 2710 1420 2711
rect 1638 2715 1644 2716
rect 1638 2711 1639 2715
rect 1643 2711 1644 2715
rect 1638 2710 1644 2711
rect 670 2707 676 2708
rect 390 2703 396 2704
rect 390 2699 391 2703
rect 395 2699 396 2703
rect 670 2703 671 2707
rect 675 2703 676 2707
rect 670 2702 676 2703
rect 1046 2707 1052 2708
rect 1046 2703 1047 2707
rect 1051 2703 1052 2707
rect 1046 2702 1052 2703
rect 390 2698 396 2699
rect 382 2674 388 2675
rect 382 2670 383 2674
rect 387 2670 388 2674
rect 382 2669 388 2670
rect 582 2674 588 2675
rect 582 2670 583 2674
rect 587 2670 588 2674
rect 582 2669 588 2670
rect 384 2651 386 2669
rect 584 2651 586 2669
rect 255 2650 259 2651
rect 255 2645 259 2646
rect 383 2650 387 2651
rect 383 2645 387 2646
rect 423 2650 427 2651
rect 423 2645 427 2646
rect 583 2650 587 2651
rect 583 2645 587 2646
rect 599 2650 603 2651
rect 599 2645 603 2646
rect 256 2635 258 2645
rect 424 2635 426 2645
rect 600 2635 602 2645
rect 254 2634 260 2635
rect 254 2630 255 2634
rect 259 2630 260 2634
rect 254 2629 260 2630
rect 422 2634 428 2635
rect 422 2630 423 2634
rect 427 2630 428 2634
rect 422 2629 428 2630
rect 598 2634 604 2635
rect 598 2630 599 2634
rect 603 2630 604 2634
rect 598 2629 604 2630
rect 246 2603 252 2604
rect 246 2599 247 2603
rect 251 2599 252 2603
rect 246 2598 252 2599
rect 254 2593 260 2594
rect 254 2589 255 2593
rect 259 2589 260 2593
rect 254 2588 260 2589
rect 422 2593 428 2594
rect 422 2589 423 2593
rect 427 2589 428 2593
rect 422 2588 428 2589
rect 598 2593 604 2594
rect 598 2589 599 2593
rect 603 2589 604 2593
rect 598 2588 604 2589
rect 256 2575 258 2588
rect 424 2575 426 2588
rect 600 2575 602 2588
rect 672 2584 674 2702
rect 782 2674 788 2675
rect 782 2670 783 2674
rect 787 2670 788 2674
rect 782 2669 788 2670
rect 982 2674 988 2675
rect 982 2670 983 2674
rect 987 2670 988 2674
rect 982 2669 988 2670
rect 1198 2674 1204 2675
rect 1198 2670 1199 2674
rect 1203 2670 1204 2674
rect 1198 2669 1204 2670
rect 1414 2674 1420 2675
rect 1414 2670 1415 2674
rect 1419 2670 1420 2674
rect 1414 2669 1420 2670
rect 1638 2674 1644 2675
rect 1638 2670 1639 2674
rect 1643 2670 1644 2674
rect 1638 2669 1644 2670
rect 784 2651 786 2669
rect 984 2651 986 2669
rect 1200 2651 1202 2669
rect 1416 2651 1418 2669
rect 1640 2651 1642 2669
rect 775 2650 779 2651
rect 775 2645 779 2646
rect 783 2650 787 2651
rect 783 2645 787 2646
rect 959 2650 963 2651
rect 959 2645 963 2646
rect 983 2650 987 2651
rect 983 2645 987 2646
rect 1151 2650 1155 2651
rect 1151 2645 1155 2646
rect 1199 2650 1203 2651
rect 1199 2645 1203 2646
rect 1343 2650 1347 2651
rect 1343 2645 1347 2646
rect 1415 2650 1419 2651
rect 1415 2645 1419 2646
rect 1535 2650 1539 2651
rect 1535 2645 1539 2646
rect 1639 2650 1643 2651
rect 1639 2645 1643 2646
rect 776 2635 778 2645
rect 960 2635 962 2645
rect 1152 2635 1154 2645
rect 1344 2635 1346 2645
rect 1536 2635 1538 2645
rect 774 2634 780 2635
rect 774 2630 775 2634
rect 779 2630 780 2634
rect 774 2629 780 2630
rect 958 2634 964 2635
rect 958 2630 959 2634
rect 963 2630 964 2634
rect 958 2629 964 2630
rect 1150 2634 1156 2635
rect 1150 2630 1151 2634
rect 1155 2630 1156 2634
rect 1150 2629 1156 2630
rect 1342 2634 1348 2635
rect 1342 2630 1343 2634
rect 1347 2630 1348 2634
rect 1342 2629 1348 2630
rect 1534 2634 1540 2635
rect 1534 2630 1535 2634
rect 1539 2630 1540 2634
rect 1534 2629 1540 2630
rect 1648 2624 1650 2718
rect 1872 2716 1874 2725
rect 1904 2724 1906 2754
rect 2032 2731 2034 2763
rect 2072 2739 2074 2779
rect 2166 2775 2172 2776
rect 2166 2771 2167 2775
rect 2171 2771 2172 2775
rect 2166 2770 2172 2771
rect 2142 2765 2148 2766
rect 2142 2761 2143 2765
rect 2147 2761 2148 2765
rect 2142 2760 2148 2761
rect 2144 2739 2146 2760
rect 2071 2738 2075 2739
rect 2071 2733 2075 2734
rect 2111 2738 2115 2739
rect 2111 2733 2115 2734
rect 2143 2738 2147 2739
rect 2143 2733 2147 2734
rect 2031 2730 2035 2731
rect 2031 2725 2035 2726
rect 1902 2723 1908 2724
rect 1902 2719 1903 2723
rect 1907 2719 1908 2723
rect 1902 2718 1908 2719
rect 1870 2715 1876 2716
rect 1870 2711 1871 2715
rect 1875 2711 1876 2715
rect 1870 2710 1876 2711
rect 1998 2707 2004 2708
rect 1998 2703 1999 2707
rect 2003 2703 2004 2707
rect 1998 2702 2004 2703
rect 1870 2674 1876 2675
rect 1870 2670 1871 2674
rect 1875 2670 1876 2674
rect 1870 2669 1876 2670
rect 1872 2651 1874 2669
rect 1727 2650 1731 2651
rect 1727 2645 1731 2646
rect 1871 2650 1875 2651
rect 1871 2645 1875 2646
rect 1927 2650 1931 2651
rect 1927 2645 1931 2646
rect 1728 2635 1730 2645
rect 1928 2635 1930 2645
rect 1726 2634 1732 2635
rect 1726 2630 1727 2634
rect 1731 2630 1732 2634
rect 1726 2629 1732 2630
rect 1926 2634 1932 2635
rect 1926 2630 1927 2634
rect 1931 2630 1932 2634
rect 1926 2629 1932 2630
rect 1222 2623 1228 2624
rect 1222 2619 1223 2623
rect 1227 2619 1228 2623
rect 1222 2618 1228 2619
rect 1646 2623 1652 2624
rect 1646 2619 1647 2623
rect 1651 2619 1652 2623
rect 1646 2618 1652 2619
rect 1224 2604 1226 2618
rect 798 2603 804 2604
rect 798 2599 799 2603
rect 803 2599 804 2603
rect 798 2598 804 2599
rect 1222 2603 1228 2604
rect 1222 2599 1223 2603
rect 1227 2599 1228 2603
rect 1222 2598 1228 2599
rect 1798 2603 1804 2604
rect 1798 2599 1799 2603
rect 1803 2599 1804 2603
rect 1798 2598 1804 2599
rect 774 2593 780 2594
rect 774 2589 775 2593
rect 779 2589 780 2593
rect 774 2588 780 2589
rect 670 2583 676 2584
rect 670 2579 671 2583
rect 675 2579 676 2583
rect 670 2578 676 2579
rect 776 2575 778 2588
rect 111 2574 115 2575
rect 111 2569 115 2570
rect 255 2574 259 2575
rect 255 2569 259 2570
rect 319 2574 323 2575
rect 319 2569 323 2570
rect 423 2574 427 2575
rect 423 2569 427 2570
rect 535 2574 539 2575
rect 535 2569 539 2570
rect 599 2574 603 2575
rect 599 2569 603 2570
rect 743 2574 747 2575
rect 743 2569 747 2570
rect 775 2574 779 2575
rect 775 2569 779 2570
rect 112 2541 114 2569
rect 320 2560 322 2569
rect 430 2567 436 2568
rect 430 2563 431 2567
rect 435 2563 436 2567
rect 430 2562 436 2563
rect 318 2559 324 2560
rect 318 2555 319 2559
rect 323 2555 324 2559
rect 318 2554 324 2555
rect 110 2540 116 2541
rect 110 2536 111 2540
rect 115 2536 116 2540
rect 110 2535 116 2536
rect 110 2523 116 2524
rect 110 2519 111 2523
rect 115 2519 116 2523
rect 110 2518 116 2519
rect 318 2518 324 2519
rect 112 2503 114 2518
rect 318 2514 319 2518
rect 323 2514 324 2518
rect 318 2513 324 2514
rect 320 2503 322 2513
rect 111 2502 115 2503
rect 111 2497 115 2498
rect 279 2502 283 2503
rect 279 2497 283 2498
rect 319 2502 323 2503
rect 319 2497 323 2498
rect 112 2482 114 2497
rect 280 2487 282 2497
rect 278 2486 284 2487
rect 278 2482 279 2486
rect 283 2482 284 2486
rect 110 2481 116 2482
rect 278 2481 284 2482
rect 110 2477 111 2481
rect 115 2477 116 2481
rect 110 2476 116 2477
rect 110 2464 116 2465
rect 110 2460 111 2464
rect 115 2460 116 2464
rect 110 2459 116 2460
rect 112 2423 114 2459
rect 432 2456 434 2562
rect 536 2560 538 2569
rect 744 2560 746 2569
rect 800 2568 802 2598
rect 958 2593 964 2594
rect 958 2589 959 2593
rect 963 2589 964 2593
rect 958 2588 964 2589
rect 1150 2593 1156 2594
rect 1150 2589 1151 2593
rect 1155 2589 1156 2593
rect 1150 2588 1156 2589
rect 1342 2593 1348 2594
rect 1342 2589 1343 2593
rect 1347 2589 1348 2593
rect 1342 2588 1348 2589
rect 1534 2593 1540 2594
rect 1534 2589 1535 2593
rect 1539 2589 1540 2593
rect 1534 2588 1540 2589
rect 1726 2593 1732 2594
rect 1726 2589 1727 2593
rect 1731 2589 1732 2593
rect 1726 2588 1732 2589
rect 960 2575 962 2588
rect 1152 2575 1154 2588
rect 1344 2575 1346 2588
rect 1536 2575 1538 2588
rect 1582 2583 1588 2584
rect 1582 2579 1583 2583
rect 1587 2579 1588 2583
rect 1582 2578 1588 2579
rect 951 2574 955 2575
rect 951 2569 955 2570
rect 959 2574 963 2575
rect 959 2569 963 2570
rect 1151 2574 1155 2575
rect 1151 2569 1155 2570
rect 1159 2574 1163 2575
rect 1159 2569 1163 2570
rect 1343 2574 1347 2575
rect 1343 2569 1347 2570
rect 1359 2574 1363 2575
rect 1359 2569 1363 2570
rect 1535 2574 1539 2575
rect 1535 2569 1539 2570
rect 1559 2574 1563 2575
rect 1559 2569 1563 2570
rect 798 2567 804 2568
rect 798 2563 799 2567
rect 803 2563 804 2567
rect 798 2562 804 2563
rect 952 2560 954 2569
rect 1160 2560 1162 2569
rect 1360 2560 1362 2569
rect 1454 2567 1460 2568
rect 1454 2563 1455 2567
rect 1459 2563 1460 2567
rect 1454 2562 1460 2563
rect 534 2559 540 2560
rect 534 2555 535 2559
rect 539 2555 540 2559
rect 534 2554 540 2555
rect 742 2559 748 2560
rect 742 2555 743 2559
rect 747 2555 748 2559
rect 742 2554 748 2555
rect 950 2559 956 2560
rect 950 2555 951 2559
rect 955 2555 956 2559
rect 950 2554 956 2555
rect 1158 2559 1164 2560
rect 1158 2555 1159 2559
rect 1163 2555 1164 2559
rect 1158 2554 1164 2555
rect 1358 2559 1364 2560
rect 1358 2555 1359 2559
rect 1363 2555 1364 2559
rect 1358 2554 1364 2555
rect 1030 2551 1036 2552
rect 1030 2547 1031 2551
rect 1035 2547 1036 2551
rect 1030 2546 1036 2547
rect 534 2518 540 2519
rect 534 2514 535 2518
rect 539 2514 540 2518
rect 534 2513 540 2514
rect 742 2518 748 2519
rect 742 2514 743 2518
rect 747 2514 748 2518
rect 742 2513 748 2514
rect 950 2518 956 2519
rect 950 2514 951 2518
rect 955 2514 956 2518
rect 950 2513 956 2514
rect 536 2503 538 2513
rect 744 2503 746 2513
rect 952 2503 954 2513
rect 439 2502 443 2503
rect 439 2497 443 2498
rect 535 2502 539 2503
rect 535 2497 539 2498
rect 607 2502 611 2503
rect 607 2497 611 2498
rect 743 2502 747 2503
rect 743 2497 747 2498
rect 783 2502 787 2503
rect 783 2497 787 2498
rect 951 2502 955 2503
rect 951 2497 955 2498
rect 959 2502 963 2503
rect 959 2497 963 2498
rect 440 2487 442 2497
rect 608 2487 610 2497
rect 784 2487 786 2497
rect 960 2487 962 2497
rect 438 2486 444 2487
rect 438 2482 439 2486
rect 443 2482 444 2486
rect 438 2481 444 2482
rect 606 2486 612 2487
rect 606 2482 607 2486
rect 611 2482 612 2486
rect 606 2481 612 2482
rect 782 2486 788 2487
rect 782 2482 783 2486
rect 787 2482 788 2486
rect 782 2481 788 2482
rect 958 2486 964 2487
rect 958 2482 959 2486
rect 963 2482 964 2486
rect 958 2481 964 2482
rect 418 2455 424 2456
rect 418 2451 419 2455
rect 423 2451 424 2455
rect 418 2450 424 2451
rect 430 2455 436 2456
rect 430 2451 431 2455
rect 435 2451 436 2455
rect 430 2450 436 2451
rect 678 2455 684 2456
rect 678 2451 679 2455
rect 683 2451 684 2455
rect 678 2450 684 2451
rect 278 2445 284 2446
rect 278 2441 279 2445
rect 283 2441 284 2445
rect 278 2440 284 2441
rect 280 2423 282 2440
rect 420 2436 422 2450
rect 438 2445 444 2446
rect 438 2441 439 2445
rect 443 2441 444 2445
rect 438 2440 444 2441
rect 606 2445 612 2446
rect 606 2441 607 2445
rect 611 2441 612 2445
rect 606 2440 612 2441
rect 350 2435 356 2436
rect 350 2431 351 2435
rect 355 2431 356 2435
rect 350 2430 356 2431
rect 418 2435 424 2436
rect 418 2431 419 2435
rect 423 2431 424 2435
rect 418 2430 424 2431
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 279 2422 283 2423
rect 279 2417 283 2418
rect 327 2422 331 2423
rect 327 2417 331 2418
rect 112 2389 114 2417
rect 328 2408 330 2417
rect 326 2407 332 2408
rect 326 2403 327 2407
rect 331 2403 332 2407
rect 326 2402 332 2403
rect 352 2396 354 2430
rect 440 2423 442 2440
rect 608 2423 610 2440
rect 439 2422 443 2423
rect 439 2417 443 2418
rect 471 2422 475 2423
rect 471 2417 475 2418
rect 607 2422 611 2423
rect 607 2417 611 2418
rect 623 2422 627 2423
rect 623 2417 627 2418
rect 472 2408 474 2417
rect 624 2408 626 2417
rect 680 2416 682 2450
rect 782 2445 788 2446
rect 782 2441 783 2445
rect 787 2441 788 2445
rect 782 2440 788 2441
rect 958 2445 964 2446
rect 958 2441 959 2445
rect 963 2441 964 2445
rect 958 2440 964 2441
rect 784 2423 786 2440
rect 960 2423 962 2440
rect 1032 2436 1034 2546
rect 1158 2518 1164 2519
rect 1158 2514 1159 2518
rect 1163 2514 1164 2518
rect 1158 2513 1164 2514
rect 1358 2518 1364 2519
rect 1358 2514 1359 2518
rect 1363 2514 1364 2518
rect 1358 2513 1364 2514
rect 1160 2503 1162 2513
rect 1360 2503 1362 2513
rect 1127 2502 1131 2503
rect 1127 2497 1131 2498
rect 1159 2502 1163 2503
rect 1159 2497 1163 2498
rect 1295 2502 1299 2503
rect 1295 2497 1299 2498
rect 1359 2502 1363 2503
rect 1359 2497 1363 2498
rect 1128 2487 1130 2497
rect 1296 2487 1298 2497
rect 1126 2486 1132 2487
rect 1126 2482 1127 2486
rect 1131 2482 1132 2486
rect 1126 2481 1132 2482
rect 1294 2486 1300 2487
rect 1294 2482 1295 2486
rect 1299 2482 1300 2486
rect 1294 2481 1300 2482
rect 1456 2456 1458 2562
rect 1560 2560 1562 2569
rect 1558 2559 1564 2560
rect 1558 2555 1559 2559
rect 1563 2555 1564 2559
rect 1558 2554 1564 2555
rect 1584 2548 1586 2578
rect 1728 2575 1730 2588
rect 1727 2574 1731 2575
rect 1727 2569 1731 2570
rect 1759 2574 1763 2575
rect 1759 2569 1763 2570
rect 1760 2560 1762 2569
rect 1800 2568 1802 2598
rect 1926 2593 1932 2594
rect 1926 2589 1927 2593
rect 1931 2589 1932 2593
rect 1926 2588 1932 2589
rect 1928 2575 1930 2588
rect 2000 2584 2002 2702
rect 2032 2697 2034 2725
rect 2072 2705 2074 2733
rect 2112 2724 2114 2733
rect 2168 2732 2170 2770
rect 2232 2764 2234 2878
rect 2278 2850 2284 2851
rect 2278 2846 2279 2850
rect 2283 2846 2284 2850
rect 2278 2845 2284 2846
rect 2486 2850 2492 2851
rect 2486 2846 2487 2850
rect 2491 2846 2492 2850
rect 2486 2845 2492 2846
rect 2694 2850 2700 2851
rect 2694 2846 2695 2850
rect 2699 2846 2700 2850
rect 2694 2845 2700 2846
rect 2902 2850 2908 2851
rect 2902 2846 2903 2850
rect 2907 2846 2908 2850
rect 2902 2845 2908 2846
rect 2280 2823 2282 2845
rect 2488 2823 2490 2845
rect 2696 2823 2698 2845
rect 2904 2823 2906 2845
rect 2279 2822 2283 2823
rect 2279 2817 2283 2818
rect 2319 2822 2323 2823
rect 2319 2817 2323 2818
rect 2487 2822 2491 2823
rect 2487 2817 2491 2818
rect 2503 2822 2507 2823
rect 2503 2817 2507 2818
rect 2695 2822 2699 2823
rect 2695 2817 2699 2818
rect 2887 2822 2891 2823
rect 2887 2817 2891 2818
rect 2903 2822 2907 2823
rect 2903 2817 2907 2818
rect 2320 2807 2322 2817
rect 2504 2807 2506 2817
rect 2696 2807 2698 2817
rect 2888 2807 2890 2817
rect 2318 2806 2324 2807
rect 2318 2802 2319 2806
rect 2323 2802 2324 2806
rect 2318 2801 2324 2802
rect 2502 2806 2508 2807
rect 2502 2802 2503 2806
rect 2507 2802 2508 2806
rect 2502 2801 2508 2802
rect 2694 2806 2700 2807
rect 2694 2802 2695 2806
rect 2699 2802 2700 2806
rect 2694 2801 2700 2802
rect 2886 2806 2892 2807
rect 2886 2802 2887 2806
rect 2891 2802 2892 2806
rect 2886 2801 2892 2802
rect 2976 2776 2978 2894
rect 3112 2892 3114 2901
rect 3304 2892 3306 2901
rect 3496 2892 3498 2901
rect 3688 2892 3690 2901
rect 3880 2892 3882 2901
rect 3110 2891 3116 2892
rect 3110 2887 3111 2891
rect 3115 2887 3116 2891
rect 3110 2886 3116 2887
rect 3302 2891 3308 2892
rect 3302 2887 3303 2891
rect 3307 2887 3308 2891
rect 3302 2886 3308 2887
rect 3494 2891 3500 2892
rect 3494 2887 3495 2891
rect 3499 2887 3500 2891
rect 3494 2886 3500 2887
rect 3686 2891 3692 2892
rect 3686 2887 3687 2891
rect 3691 2887 3692 2891
rect 3686 2886 3692 2887
rect 3878 2891 3884 2892
rect 3878 2887 3879 2891
rect 3883 2887 3884 2891
rect 3878 2886 3884 2887
rect 3286 2883 3292 2884
rect 3286 2879 3287 2883
rect 3291 2879 3292 2883
rect 3286 2878 3292 2879
rect 3110 2850 3116 2851
rect 3110 2846 3111 2850
rect 3115 2846 3116 2850
rect 3110 2845 3116 2846
rect 3112 2823 3114 2845
rect 3288 2824 3290 2878
rect 3992 2873 3994 2901
rect 3990 2872 3996 2873
rect 3990 2868 3991 2872
rect 3995 2868 3996 2872
rect 3990 2867 3996 2868
rect 3990 2855 3996 2856
rect 3990 2851 3991 2855
rect 3995 2851 3996 2855
rect 3302 2850 3308 2851
rect 3302 2846 3303 2850
rect 3307 2846 3308 2850
rect 3302 2845 3308 2846
rect 3494 2850 3500 2851
rect 3494 2846 3495 2850
rect 3499 2846 3500 2850
rect 3494 2845 3500 2846
rect 3686 2850 3692 2851
rect 3686 2846 3687 2850
rect 3691 2846 3692 2850
rect 3686 2845 3692 2846
rect 3878 2850 3884 2851
rect 3990 2850 3996 2851
rect 3878 2846 3879 2850
rect 3883 2846 3884 2850
rect 3878 2845 3884 2846
rect 3286 2823 3292 2824
rect 3304 2823 3306 2845
rect 3496 2823 3498 2845
rect 3688 2823 3690 2845
rect 3838 2823 3844 2824
rect 3880 2823 3882 2845
rect 3992 2823 3994 2850
rect 3079 2822 3083 2823
rect 3079 2817 3083 2818
rect 3111 2822 3115 2823
rect 3111 2817 3115 2818
rect 3263 2822 3267 2823
rect 3286 2819 3287 2823
rect 3291 2819 3292 2823
rect 3286 2818 3292 2819
rect 3303 2822 3307 2823
rect 3263 2817 3267 2818
rect 3303 2817 3307 2818
rect 3439 2822 3443 2823
rect 3439 2817 3443 2818
rect 3495 2822 3499 2823
rect 3495 2817 3499 2818
rect 3615 2822 3619 2823
rect 3615 2817 3619 2818
rect 3687 2822 3691 2823
rect 3687 2817 3691 2818
rect 3791 2822 3795 2823
rect 3838 2819 3839 2823
rect 3843 2819 3844 2823
rect 3838 2818 3844 2819
rect 3879 2822 3883 2823
rect 3791 2817 3795 2818
rect 3080 2807 3082 2817
rect 3264 2807 3266 2817
rect 3440 2807 3442 2817
rect 3616 2807 3618 2817
rect 3792 2807 3794 2817
rect 3078 2806 3084 2807
rect 3078 2802 3079 2806
rect 3083 2802 3084 2806
rect 3078 2801 3084 2802
rect 3262 2806 3268 2807
rect 3262 2802 3263 2806
rect 3267 2802 3268 2806
rect 3262 2801 3268 2802
rect 3438 2806 3444 2807
rect 3438 2802 3439 2806
rect 3443 2802 3444 2806
rect 3438 2801 3444 2802
rect 3614 2806 3620 2807
rect 3614 2802 3615 2806
rect 3619 2802 3620 2806
rect 3614 2801 3620 2802
rect 3790 2806 3796 2807
rect 3790 2802 3791 2806
rect 3795 2802 3796 2806
rect 3790 2801 3796 2802
rect 2678 2775 2684 2776
rect 2678 2771 2679 2775
rect 2683 2771 2684 2775
rect 2678 2770 2684 2771
rect 2870 2775 2876 2776
rect 2870 2771 2871 2775
rect 2875 2771 2876 2775
rect 2870 2770 2876 2771
rect 2974 2775 2980 2776
rect 2974 2771 2975 2775
rect 2979 2771 2980 2775
rect 2974 2770 2980 2771
rect 3246 2775 3252 2776
rect 3246 2771 3247 2775
rect 3251 2771 3252 2775
rect 3246 2770 3252 2771
rect 2318 2765 2324 2766
rect 2230 2763 2236 2764
rect 2230 2759 2231 2763
rect 2235 2759 2236 2763
rect 2318 2761 2319 2765
rect 2323 2761 2324 2765
rect 2318 2760 2324 2761
rect 2502 2765 2508 2766
rect 2502 2761 2503 2765
rect 2507 2761 2508 2765
rect 2502 2760 2508 2761
rect 2230 2758 2236 2759
rect 2320 2739 2322 2760
rect 2504 2739 2506 2760
rect 2680 2756 2682 2770
rect 2694 2765 2700 2766
rect 2694 2761 2695 2765
rect 2699 2761 2700 2765
rect 2694 2760 2700 2761
rect 2518 2755 2524 2756
rect 2518 2751 2519 2755
rect 2523 2751 2524 2755
rect 2518 2750 2524 2751
rect 2678 2755 2684 2756
rect 2678 2751 2679 2755
rect 2683 2751 2684 2755
rect 2678 2750 2684 2751
rect 2279 2738 2283 2739
rect 2279 2733 2283 2734
rect 2319 2738 2323 2739
rect 2319 2733 2323 2734
rect 2455 2738 2459 2739
rect 2455 2733 2459 2734
rect 2503 2738 2507 2739
rect 2503 2733 2507 2734
rect 2166 2731 2172 2732
rect 2166 2727 2167 2731
rect 2171 2727 2172 2731
rect 2166 2726 2172 2727
rect 2280 2724 2282 2733
rect 2456 2724 2458 2733
rect 2110 2723 2116 2724
rect 2110 2719 2111 2723
rect 2115 2719 2116 2723
rect 2110 2718 2116 2719
rect 2278 2723 2284 2724
rect 2278 2719 2279 2723
rect 2283 2719 2284 2723
rect 2278 2718 2284 2719
rect 2454 2723 2460 2724
rect 2454 2719 2455 2723
rect 2459 2719 2460 2723
rect 2454 2718 2460 2719
rect 2520 2716 2522 2750
rect 2696 2739 2698 2760
rect 2872 2756 2874 2770
rect 2886 2765 2892 2766
rect 2886 2761 2887 2765
rect 2891 2761 2892 2765
rect 2886 2760 2892 2761
rect 3078 2765 3084 2766
rect 3078 2761 3079 2765
rect 3083 2761 3084 2765
rect 3078 2760 3084 2761
rect 2870 2755 2876 2756
rect 2870 2751 2871 2755
rect 2875 2751 2876 2755
rect 2870 2750 2876 2751
rect 2888 2739 2890 2760
rect 3080 2739 3082 2760
rect 3248 2740 3250 2770
rect 3262 2765 3268 2766
rect 3262 2761 3263 2765
rect 3267 2761 3268 2765
rect 3262 2760 3268 2761
rect 3438 2765 3444 2766
rect 3438 2761 3439 2765
rect 3443 2761 3444 2765
rect 3438 2760 3444 2761
rect 3614 2765 3620 2766
rect 3614 2761 3615 2765
rect 3619 2761 3620 2765
rect 3614 2760 3620 2761
rect 3790 2765 3796 2766
rect 3790 2761 3791 2765
rect 3795 2761 3796 2765
rect 3790 2760 3796 2761
rect 3246 2739 3252 2740
rect 3264 2739 3266 2760
rect 3440 2739 3442 2760
rect 3616 2739 3618 2760
rect 3792 2739 3794 2760
rect 3840 2756 3842 2818
rect 3879 2817 3883 2818
rect 3991 2822 3995 2823
rect 3991 2817 3995 2818
rect 3992 2802 3994 2817
rect 3990 2801 3996 2802
rect 3990 2797 3991 2801
rect 3995 2797 3996 2801
rect 3990 2796 3996 2797
rect 3990 2784 3996 2785
rect 3990 2780 3991 2784
rect 3995 2780 3996 2784
rect 3990 2779 3996 2780
rect 3838 2755 3844 2756
rect 3838 2751 3839 2755
rect 3843 2751 3844 2755
rect 3838 2750 3844 2751
rect 3992 2739 3994 2779
rect 2639 2738 2643 2739
rect 2639 2733 2643 2734
rect 2695 2738 2699 2739
rect 2695 2733 2699 2734
rect 2815 2738 2819 2739
rect 2815 2733 2819 2734
rect 2887 2738 2891 2739
rect 2887 2733 2891 2734
rect 2983 2738 2987 2739
rect 2983 2733 2987 2734
rect 3079 2738 3083 2739
rect 3079 2733 3083 2734
rect 3143 2738 3147 2739
rect 3246 2735 3247 2739
rect 3251 2735 3252 2739
rect 3246 2734 3252 2735
rect 3263 2738 3267 2739
rect 3143 2733 3147 2734
rect 3263 2733 3267 2734
rect 3303 2738 3307 2739
rect 3303 2733 3307 2734
rect 3439 2738 3443 2739
rect 3439 2733 3443 2734
rect 3463 2738 3467 2739
rect 3463 2733 3467 2734
rect 3615 2738 3619 2739
rect 3615 2733 3619 2734
rect 3623 2738 3627 2739
rect 3623 2733 3627 2734
rect 3791 2738 3795 2739
rect 3791 2733 3795 2734
rect 3991 2738 3995 2739
rect 3991 2733 3995 2734
rect 2640 2724 2642 2733
rect 2816 2724 2818 2733
rect 2862 2731 2868 2732
rect 2862 2727 2863 2731
rect 2867 2727 2868 2731
rect 2862 2726 2868 2727
rect 2638 2723 2644 2724
rect 2638 2719 2639 2723
rect 2643 2719 2644 2723
rect 2638 2718 2644 2719
rect 2814 2723 2820 2724
rect 2814 2719 2815 2723
rect 2819 2719 2820 2723
rect 2814 2718 2820 2719
rect 2342 2715 2348 2716
rect 2342 2711 2343 2715
rect 2347 2711 2348 2715
rect 2342 2710 2348 2711
rect 2518 2715 2524 2716
rect 2518 2711 2519 2715
rect 2523 2711 2524 2715
rect 2518 2710 2524 2711
rect 2070 2704 2076 2705
rect 2070 2700 2071 2704
rect 2075 2700 2076 2704
rect 2070 2699 2076 2700
rect 2030 2696 2036 2697
rect 2030 2692 2031 2696
rect 2035 2692 2036 2696
rect 2030 2691 2036 2692
rect 2070 2687 2076 2688
rect 2070 2683 2071 2687
rect 2075 2683 2076 2687
rect 2070 2682 2076 2683
rect 2110 2682 2116 2683
rect 2030 2679 2036 2680
rect 2030 2675 2031 2679
rect 2035 2675 2036 2679
rect 2030 2674 2036 2675
rect 2032 2651 2034 2674
rect 2072 2655 2074 2682
rect 2110 2678 2111 2682
rect 2115 2678 2116 2682
rect 2110 2677 2116 2678
rect 2278 2682 2284 2683
rect 2278 2678 2279 2682
rect 2283 2678 2284 2682
rect 2278 2677 2284 2678
rect 2112 2655 2114 2677
rect 2280 2655 2282 2677
rect 2071 2654 2075 2655
rect 2031 2650 2035 2651
rect 2071 2649 2075 2650
rect 2111 2654 2115 2655
rect 2111 2649 2115 2650
rect 2263 2654 2267 2655
rect 2263 2649 2267 2650
rect 2279 2654 2283 2655
rect 2279 2649 2283 2650
rect 2031 2645 2035 2646
rect 2032 2630 2034 2645
rect 2072 2634 2074 2649
rect 2112 2639 2114 2649
rect 2264 2639 2266 2649
rect 2110 2638 2116 2639
rect 2110 2634 2111 2638
rect 2115 2634 2116 2638
rect 2070 2633 2076 2634
rect 2110 2633 2116 2634
rect 2262 2638 2268 2639
rect 2262 2634 2263 2638
rect 2267 2634 2268 2638
rect 2262 2633 2268 2634
rect 2030 2629 2036 2630
rect 2030 2625 2031 2629
rect 2035 2625 2036 2629
rect 2070 2629 2071 2633
rect 2075 2629 2076 2633
rect 2070 2628 2076 2629
rect 2030 2624 2036 2625
rect 2070 2616 2076 2617
rect 2030 2612 2036 2613
rect 2030 2608 2031 2612
rect 2035 2608 2036 2612
rect 2070 2612 2071 2616
rect 2075 2612 2076 2616
rect 2070 2611 2076 2612
rect 2030 2607 2036 2608
rect 1998 2583 2004 2584
rect 1998 2579 1999 2583
rect 2003 2579 2004 2583
rect 1998 2578 2004 2579
rect 2032 2575 2034 2607
rect 2072 2575 2074 2611
rect 2182 2607 2188 2608
rect 2182 2603 2183 2607
rect 2187 2603 2188 2607
rect 2182 2602 2188 2603
rect 2110 2597 2116 2598
rect 2110 2593 2111 2597
rect 2115 2593 2116 2597
rect 2110 2592 2116 2593
rect 2112 2575 2114 2592
rect 1927 2574 1931 2575
rect 1927 2569 1931 2570
rect 1935 2574 1939 2575
rect 1935 2569 1939 2570
rect 2031 2574 2035 2575
rect 2031 2569 2035 2570
rect 2071 2574 2075 2575
rect 2071 2569 2075 2570
rect 2111 2574 2115 2575
rect 2111 2569 2115 2570
rect 1798 2567 1804 2568
rect 1798 2563 1799 2567
rect 1803 2563 1804 2567
rect 1798 2562 1804 2563
rect 1936 2560 1938 2569
rect 1758 2559 1764 2560
rect 1758 2555 1759 2559
rect 1763 2555 1764 2559
rect 1758 2554 1764 2555
rect 1934 2559 1940 2560
rect 1934 2555 1935 2559
rect 1939 2555 1940 2559
rect 1934 2554 1940 2555
rect 1858 2551 1864 2552
rect 1582 2547 1588 2548
rect 1582 2543 1583 2547
rect 1587 2543 1588 2547
rect 1858 2547 1859 2551
rect 1863 2547 1864 2551
rect 1858 2546 1864 2547
rect 2006 2551 2012 2552
rect 2006 2547 2007 2551
rect 2011 2547 2012 2551
rect 2006 2546 2012 2547
rect 1582 2542 1588 2543
rect 1558 2518 1564 2519
rect 1558 2514 1559 2518
rect 1563 2514 1564 2518
rect 1558 2513 1564 2514
rect 1758 2518 1764 2519
rect 1758 2514 1759 2518
rect 1763 2514 1764 2518
rect 1758 2513 1764 2514
rect 1560 2503 1562 2513
rect 1760 2503 1762 2513
rect 1463 2502 1467 2503
rect 1463 2497 1467 2498
rect 1559 2502 1563 2503
rect 1559 2497 1563 2498
rect 1623 2502 1627 2503
rect 1623 2497 1627 2498
rect 1759 2502 1763 2503
rect 1759 2497 1763 2498
rect 1791 2502 1795 2503
rect 1791 2497 1795 2498
rect 1464 2487 1466 2497
rect 1624 2487 1626 2497
rect 1792 2487 1794 2497
rect 1462 2486 1468 2487
rect 1462 2482 1463 2486
rect 1467 2482 1468 2486
rect 1462 2481 1468 2482
rect 1622 2486 1628 2487
rect 1622 2482 1623 2486
rect 1627 2482 1628 2486
rect 1622 2481 1628 2482
rect 1790 2486 1796 2487
rect 1790 2482 1791 2486
rect 1795 2482 1796 2486
rect 1790 2481 1796 2482
rect 1278 2455 1284 2456
rect 1278 2451 1279 2455
rect 1283 2451 1284 2455
rect 1278 2450 1284 2451
rect 1454 2455 1460 2456
rect 1454 2451 1455 2455
rect 1459 2451 1460 2455
rect 1454 2450 1460 2451
rect 1694 2455 1700 2456
rect 1694 2451 1695 2455
rect 1699 2451 1700 2455
rect 1694 2450 1700 2451
rect 1126 2445 1132 2446
rect 1126 2441 1127 2445
rect 1131 2441 1132 2445
rect 1126 2440 1132 2441
rect 1030 2435 1036 2436
rect 1030 2431 1031 2435
rect 1035 2431 1036 2435
rect 1030 2430 1036 2431
rect 1128 2423 1130 2440
rect 1280 2428 1282 2450
rect 1294 2445 1300 2446
rect 1294 2441 1295 2445
rect 1299 2441 1300 2445
rect 1294 2440 1300 2441
rect 1462 2445 1468 2446
rect 1462 2441 1463 2445
rect 1467 2441 1468 2445
rect 1462 2440 1468 2441
rect 1622 2445 1628 2446
rect 1622 2441 1623 2445
rect 1627 2441 1628 2445
rect 1622 2440 1628 2441
rect 1278 2427 1284 2428
rect 1278 2423 1279 2427
rect 1283 2423 1284 2427
rect 1296 2423 1298 2440
rect 1370 2435 1376 2436
rect 1370 2431 1371 2435
rect 1375 2431 1376 2435
rect 1370 2430 1376 2431
rect 783 2422 787 2423
rect 783 2417 787 2418
rect 943 2422 947 2423
rect 943 2417 947 2418
rect 959 2422 963 2423
rect 959 2417 963 2418
rect 1095 2422 1099 2423
rect 1095 2417 1099 2418
rect 1127 2422 1131 2423
rect 1127 2417 1131 2418
rect 1247 2422 1251 2423
rect 1278 2422 1284 2423
rect 1295 2422 1299 2423
rect 1247 2417 1251 2418
rect 1295 2417 1299 2418
rect 678 2415 684 2416
rect 678 2411 679 2415
rect 683 2411 684 2415
rect 678 2410 684 2411
rect 784 2408 786 2417
rect 944 2408 946 2417
rect 1006 2415 1012 2416
rect 1006 2411 1007 2415
rect 1011 2411 1012 2415
rect 1006 2410 1012 2411
rect 470 2407 476 2408
rect 470 2403 471 2407
rect 475 2403 476 2407
rect 470 2402 476 2403
rect 622 2407 628 2408
rect 622 2403 623 2407
rect 627 2403 628 2407
rect 622 2402 628 2403
rect 782 2407 788 2408
rect 782 2403 783 2407
rect 787 2403 788 2407
rect 782 2402 788 2403
rect 942 2407 948 2408
rect 942 2403 943 2407
rect 947 2403 948 2407
rect 942 2402 948 2403
rect 686 2399 692 2400
rect 350 2395 356 2396
rect 350 2391 351 2395
rect 355 2391 356 2395
rect 686 2395 687 2399
rect 691 2395 692 2399
rect 686 2394 692 2395
rect 350 2390 356 2391
rect 110 2388 116 2389
rect 110 2384 111 2388
rect 115 2384 116 2388
rect 110 2383 116 2384
rect 110 2371 116 2372
rect 110 2367 111 2371
rect 115 2367 116 2371
rect 110 2366 116 2367
rect 326 2366 332 2367
rect 112 2343 114 2366
rect 326 2362 327 2366
rect 331 2362 332 2366
rect 326 2361 332 2362
rect 470 2366 476 2367
rect 470 2362 471 2366
rect 475 2362 476 2366
rect 470 2361 476 2362
rect 622 2366 628 2367
rect 622 2362 623 2366
rect 627 2362 628 2366
rect 622 2361 628 2362
rect 328 2343 330 2361
rect 472 2343 474 2361
rect 624 2343 626 2361
rect 111 2342 115 2343
rect 111 2337 115 2338
rect 327 2342 331 2343
rect 327 2337 331 2338
rect 359 2342 363 2343
rect 359 2337 363 2338
rect 471 2342 475 2343
rect 471 2337 475 2338
rect 495 2342 499 2343
rect 495 2337 499 2338
rect 623 2342 627 2343
rect 623 2337 627 2338
rect 639 2342 643 2343
rect 639 2337 643 2338
rect 112 2322 114 2337
rect 360 2327 362 2337
rect 496 2327 498 2337
rect 640 2327 642 2337
rect 358 2326 364 2327
rect 358 2322 359 2326
rect 363 2322 364 2326
rect 110 2321 116 2322
rect 358 2321 364 2322
rect 494 2326 500 2327
rect 494 2322 495 2326
rect 499 2322 500 2326
rect 494 2321 500 2322
rect 638 2326 644 2327
rect 638 2322 639 2326
rect 643 2322 644 2326
rect 638 2321 644 2322
rect 110 2317 111 2321
rect 115 2317 116 2321
rect 110 2316 116 2317
rect 110 2304 116 2305
rect 110 2300 111 2304
rect 115 2300 116 2304
rect 110 2299 116 2300
rect 112 2259 114 2299
rect 478 2295 484 2296
rect 478 2291 479 2295
rect 483 2291 484 2295
rect 478 2290 484 2291
rect 358 2285 364 2286
rect 358 2281 359 2285
rect 363 2281 364 2285
rect 358 2280 364 2281
rect 360 2259 362 2280
rect 480 2260 482 2290
rect 494 2285 500 2286
rect 494 2281 495 2285
rect 499 2281 500 2285
rect 494 2280 500 2281
rect 638 2285 644 2286
rect 638 2281 639 2285
rect 643 2281 644 2285
rect 638 2280 644 2281
rect 478 2259 484 2260
rect 496 2259 498 2280
rect 640 2259 642 2280
rect 688 2276 690 2394
rect 782 2366 788 2367
rect 782 2362 783 2366
rect 787 2362 788 2366
rect 782 2361 788 2362
rect 942 2366 948 2367
rect 942 2362 943 2366
rect 947 2362 948 2366
rect 942 2361 948 2362
rect 784 2343 786 2361
rect 944 2343 946 2361
rect 783 2342 787 2343
rect 783 2337 787 2338
rect 935 2342 939 2343
rect 935 2337 939 2338
rect 943 2342 947 2343
rect 943 2337 947 2338
rect 784 2327 786 2337
rect 936 2327 938 2337
rect 782 2326 788 2327
rect 782 2322 783 2326
rect 787 2322 788 2326
rect 782 2321 788 2322
rect 934 2326 940 2327
rect 934 2322 935 2326
rect 939 2322 940 2326
rect 934 2321 940 2322
rect 1008 2296 1010 2410
rect 1096 2408 1098 2417
rect 1248 2408 1250 2417
rect 1372 2416 1374 2430
rect 1464 2423 1466 2440
rect 1624 2423 1626 2440
rect 1391 2422 1395 2423
rect 1391 2417 1395 2418
rect 1463 2422 1467 2423
rect 1463 2417 1467 2418
rect 1535 2422 1539 2423
rect 1535 2417 1539 2418
rect 1623 2422 1627 2423
rect 1623 2417 1627 2418
rect 1671 2422 1675 2423
rect 1671 2417 1675 2418
rect 1370 2415 1376 2416
rect 1370 2411 1371 2415
rect 1375 2411 1376 2415
rect 1370 2410 1376 2411
rect 1392 2408 1394 2417
rect 1536 2408 1538 2417
rect 1672 2408 1674 2417
rect 1696 2416 1698 2450
rect 1790 2445 1796 2446
rect 1790 2441 1791 2445
rect 1795 2441 1796 2445
rect 1790 2440 1796 2441
rect 1792 2423 1794 2440
rect 1860 2436 1862 2546
rect 1934 2518 1940 2519
rect 1934 2514 1935 2518
rect 1939 2514 1940 2518
rect 1934 2513 1940 2514
rect 1936 2503 1938 2513
rect 1935 2502 1939 2503
rect 1935 2497 1939 2498
rect 1936 2487 1938 2497
rect 1934 2486 1940 2487
rect 1934 2482 1935 2486
rect 1939 2482 1940 2486
rect 1934 2481 1940 2482
rect 1934 2445 1940 2446
rect 1934 2441 1935 2445
rect 1939 2441 1940 2445
rect 1934 2440 1940 2441
rect 1858 2435 1864 2436
rect 1858 2431 1859 2435
rect 1863 2431 1864 2435
rect 1858 2430 1864 2431
rect 1890 2435 1896 2436
rect 1890 2431 1891 2435
rect 1895 2431 1896 2435
rect 1890 2430 1896 2431
rect 1791 2422 1795 2423
rect 1791 2417 1795 2418
rect 1815 2422 1819 2423
rect 1815 2417 1819 2418
rect 1694 2415 1700 2416
rect 1694 2411 1695 2415
rect 1699 2411 1700 2415
rect 1694 2410 1700 2411
rect 1816 2408 1818 2417
rect 1892 2416 1894 2430
rect 1936 2423 1938 2440
rect 2008 2436 2010 2546
rect 2032 2541 2034 2569
rect 2072 2541 2074 2569
rect 2112 2560 2114 2569
rect 2184 2568 2186 2602
rect 2262 2597 2268 2598
rect 2262 2593 2263 2597
rect 2267 2593 2268 2597
rect 2262 2592 2268 2593
rect 2264 2575 2266 2592
rect 2335 2587 2341 2588
rect 2335 2583 2336 2587
rect 2340 2586 2341 2587
rect 2344 2586 2346 2710
rect 2454 2682 2460 2683
rect 2454 2678 2455 2682
rect 2459 2678 2460 2682
rect 2454 2677 2460 2678
rect 2638 2682 2644 2683
rect 2638 2678 2639 2682
rect 2643 2678 2644 2682
rect 2638 2677 2644 2678
rect 2814 2682 2820 2683
rect 2814 2678 2815 2682
rect 2819 2678 2820 2682
rect 2814 2677 2820 2678
rect 2456 2655 2458 2677
rect 2640 2655 2642 2677
rect 2816 2655 2818 2677
rect 2431 2654 2435 2655
rect 2431 2649 2435 2650
rect 2455 2654 2459 2655
rect 2455 2649 2459 2650
rect 2599 2654 2603 2655
rect 2599 2649 2603 2650
rect 2639 2654 2643 2655
rect 2639 2649 2643 2650
rect 2751 2654 2755 2655
rect 2751 2649 2755 2650
rect 2815 2654 2819 2655
rect 2815 2649 2819 2650
rect 2432 2639 2434 2649
rect 2600 2639 2602 2649
rect 2752 2639 2754 2649
rect 2430 2638 2436 2639
rect 2430 2634 2431 2638
rect 2435 2634 2436 2638
rect 2430 2633 2436 2634
rect 2598 2638 2604 2639
rect 2598 2634 2599 2638
rect 2603 2634 2604 2638
rect 2598 2633 2604 2634
rect 2750 2638 2756 2639
rect 2750 2634 2751 2638
rect 2755 2634 2756 2638
rect 2750 2633 2756 2634
rect 2864 2608 2866 2726
rect 2984 2724 2986 2733
rect 3144 2724 3146 2733
rect 3304 2724 3306 2733
rect 3464 2724 3466 2733
rect 3624 2724 3626 2733
rect 2982 2723 2988 2724
rect 2982 2719 2983 2723
rect 2987 2719 2988 2723
rect 2982 2718 2988 2719
rect 3142 2723 3148 2724
rect 3142 2719 3143 2723
rect 3147 2719 3148 2723
rect 3142 2718 3148 2719
rect 3302 2723 3308 2724
rect 3302 2719 3303 2723
rect 3307 2719 3308 2723
rect 3302 2718 3308 2719
rect 3462 2723 3468 2724
rect 3462 2719 3463 2723
rect 3467 2719 3468 2723
rect 3462 2718 3468 2719
rect 3622 2723 3628 2724
rect 3622 2719 3623 2723
rect 3627 2719 3628 2723
rect 3622 2718 3628 2719
rect 3126 2715 3132 2716
rect 3126 2711 3127 2715
rect 3131 2711 3132 2715
rect 3126 2710 3132 2711
rect 2982 2682 2988 2683
rect 2982 2678 2983 2682
rect 2987 2678 2988 2682
rect 2982 2677 2988 2678
rect 2984 2655 2986 2677
rect 2895 2654 2899 2655
rect 2895 2649 2899 2650
rect 2983 2654 2987 2655
rect 2983 2649 2987 2650
rect 3039 2654 3043 2655
rect 3039 2649 3043 2650
rect 2896 2639 2898 2649
rect 3040 2639 3042 2649
rect 2894 2638 2900 2639
rect 2894 2634 2895 2638
rect 2899 2634 2900 2638
rect 2894 2633 2900 2634
rect 3038 2638 3044 2639
rect 3038 2634 3039 2638
rect 3043 2634 3044 2638
rect 3038 2633 3044 2634
rect 2582 2607 2588 2608
rect 2582 2603 2583 2607
rect 2587 2603 2588 2607
rect 2582 2602 2588 2603
rect 2862 2607 2868 2608
rect 2862 2603 2863 2607
rect 2867 2603 2868 2607
rect 2862 2602 2868 2603
rect 3022 2607 3028 2608
rect 3022 2603 3023 2607
rect 3027 2603 3028 2607
rect 3022 2602 3028 2603
rect 2430 2597 2436 2598
rect 2430 2593 2431 2597
rect 2435 2593 2436 2597
rect 2430 2592 2436 2593
rect 2340 2584 2346 2586
rect 2340 2583 2341 2584
rect 2335 2582 2341 2583
rect 2432 2575 2434 2592
rect 2584 2580 2586 2602
rect 2598 2597 2604 2598
rect 2598 2593 2599 2597
rect 2603 2593 2604 2597
rect 2598 2592 2604 2593
rect 2750 2597 2756 2598
rect 2750 2593 2751 2597
rect 2755 2593 2756 2597
rect 2750 2592 2756 2593
rect 2894 2597 2900 2598
rect 2894 2593 2895 2597
rect 2899 2593 2900 2597
rect 2894 2592 2900 2593
rect 2582 2579 2588 2580
rect 2582 2575 2583 2579
rect 2587 2575 2588 2579
rect 2600 2575 2602 2592
rect 2682 2587 2688 2588
rect 2682 2583 2683 2587
rect 2687 2583 2688 2587
rect 2682 2582 2688 2583
rect 2263 2574 2267 2575
rect 2263 2569 2267 2570
rect 2271 2574 2275 2575
rect 2271 2569 2275 2570
rect 2431 2574 2435 2575
rect 2431 2569 2435 2570
rect 2447 2574 2451 2575
rect 2582 2574 2588 2575
rect 2599 2574 2603 2575
rect 2447 2569 2451 2570
rect 2599 2569 2603 2570
rect 2615 2574 2619 2575
rect 2615 2569 2619 2570
rect 2182 2567 2188 2568
rect 2182 2563 2183 2567
rect 2187 2563 2188 2567
rect 2182 2562 2188 2563
rect 2272 2560 2274 2569
rect 2448 2560 2450 2569
rect 2538 2567 2544 2568
rect 2538 2563 2539 2567
rect 2543 2563 2544 2567
rect 2538 2562 2544 2563
rect 2110 2559 2116 2560
rect 2110 2555 2111 2559
rect 2115 2555 2116 2559
rect 2110 2554 2116 2555
rect 2270 2559 2276 2560
rect 2270 2555 2271 2559
rect 2275 2555 2276 2559
rect 2270 2554 2276 2555
rect 2446 2559 2452 2560
rect 2446 2555 2447 2559
rect 2451 2555 2452 2559
rect 2446 2554 2452 2555
rect 2030 2540 2036 2541
rect 2030 2536 2031 2540
rect 2035 2536 2036 2540
rect 2030 2535 2036 2536
rect 2070 2540 2076 2541
rect 2070 2536 2071 2540
rect 2075 2536 2076 2540
rect 2070 2535 2076 2536
rect 2030 2523 2036 2524
rect 2030 2519 2031 2523
rect 2035 2519 2036 2523
rect 2030 2518 2036 2519
rect 2070 2523 2076 2524
rect 2070 2519 2071 2523
rect 2075 2519 2076 2523
rect 2070 2518 2076 2519
rect 2110 2518 2116 2519
rect 2032 2503 2034 2518
rect 2031 2502 2035 2503
rect 2031 2497 2035 2498
rect 2032 2482 2034 2497
rect 2072 2491 2074 2518
rect 2110 2514 2111 2518
rect 2115 2514 2116 2518
rect 2110 2513 2116 2514
rect 2270 2518 2276 2519
rect 2270 2514 2271 2518
rect 2275 2514 2276 2518
rect 2270 2513 2276 2514
rect 2446 2518 2452 2519
rect 2446 2514 2447 2518
rect 2451 2514 2452 2518
rect 2446 2513 2452 2514
rect 2112 2491 2114 2513
rect 2272 2491 2274 2513
rect 2448 2491 2450 2513
rect 2071 2490 2075 2491
rect 2071 2485 2075 2486
rect 2111 2490 2115 2491
rect 2111 2485 2115 2486
rect 2271 2490 2275 2491
rect 2271 2485 2275 2486
rect 2447 2490 2451 2491
rect 2447 2485 2451 2486
rect 2030 2481 2036 2482
rect 2030 2477 2031 2481
rect 2035 2477 2036 2481
rect 2030 2476 2036 2477
rect 2072 2470 2074 2485
rect 2070 2469 2076 2470
rect 2070 2465 2071 2469
rect 2075 2465 2076 2469
rect 2030 2464 2036 2465
rect 2070 2464 2076 2465
rect 2030 2460 2031 2464
rect 2035 2460 2036 2464
rect 2030 2459 2036 2460
rect 2006 2435 2012 2436
rect 2006 2431 2007 2435
rect 2011 2431 2012 2435
rect 2006 2430 2012 2431
rect 2032 2423 2034 2459
rect 2070 2452 2076 2453
rect 2070 2448 2071 2452
rect 2075 2448 2076 2452
rect 2070 2447 2076 2448
rect 1935 2422 1939 2423
rect 1935 2417 1939 2418
rect 2031 2422 2035 2423
rect 2031 2417 2035 2418
rect 1890 2415 1896 2416
rect 1890 2411 1891 2415
rect 1895 2411 1896 2415
rect 1890 2410 1896 2411
rect 1936 2408 1938 2417
rect 1094 2407 1100 2408
rect 1094 2403 1095 2407
rect 1099 2403 1100 2407
rect 1094 2402 1100 2403
rect 1246 2407 1252 2408
rect 1246 2403 1247 2407
rect 1251 2403 1252 2407
rect 1246 2402 1252 2403
rect 1390 2407 1396 2408
rect 1390 2403 1391 2407
rect 1395 2403 1396 2407
rect 1390 2402 1396 2403
rect 1534 2407 1540 2408
rect 1534 2403 1535 2407
rect 1539 2403 1540 2407
rect 1534 2402 1540 2403
rect 1670 2407 1676 2408
rect 1670 2403 1671 2407
rect 1675 2403 1676 2407
rect 1670 2402 1676 2403
rect 1814 2407 1820 2408
rect 1814 2403 1815 2407
rect 1819 2403 1820 2407
rect 1814 2402 1820 2403
rect 1934 2407 1940 2408
rect 1934 2403 1935 2407
rect 1939 2403 1940 2407
rect 1934 2402 1940 2403
rect 2006 2399 2012 2400
rect 1526 2395 1532 2396
rect 1526 2391 1527 2395
rect 1531 2391 1532 2395
rect 2006 2395 2007 2399
rect 2011 2395 2012 2399
rect 2006 2394 2012 2395
rect 1526 2390 1532 2391
rect 1094 2366 1100 2367
rect 1094 2362 1095 2366
rect 1099 2362 1100 2366
rect 1094 2361 1100 2362
rect 1246 2366 1252 2367
rect 1246 2362 1247 2366
rect 1251 2362 1252 2366
rect 1246 2361 1252 2362
rect 1390 2366 1396 2367
rect 1390 2362 1391 2366
rect 1395 2362 1396 2366
rect 1390 2361 1396 2362
rect 1096 2343 1098 2361
rect 1248 2343 1250 2361
rect 1392 2343 1394 2361
rect 1087 2342 1091 2343
rect 1087 2337 1091 2338
rect 1095 2342 1099 2343
rect 1095 2337 1099 2338
rect 1247 2342 1251 2343
rect 1247 2337 1251 2338
rect 1391 2342 1395 2343
rect 1391 2337 1395 2338
rect 1415 2342 1419 2343
rect 1415 2337 1419 2338
rect 1088 2327 1090 2337
rect 1248 2327 1250 2337
rect 1416 2327 1418 2337
rect 1086 2326 1092 2327
rect 1086 2322 1087 2326
rect 1091 2322 1092 2326
rect 1086 2321 1092 2322
rect 1246 2326 1252 2327
rect 1246 2322 1247 2326
rect 1251 2322 1252 2326
rect 1246 2321 1252 2322
rect 1414 2326 1420 2327
rect 1414 2322 1415 2326
rect 1419 2322 1420 2326
rect 1414 2321 1420 2322
rect 766 2295 772 2296
rect 766 2291 767 2295
rect 771 2291 772 2295
rect 766 2290 772 2291
rect 918 2295 924 2296
rect 918 2291 919 2295
rect 923 2291 924 2295
rect 918 2290 924 2291
rect 1006 2295 1012 2296
rect 1006 2291 1007 2295
rect 1011 2291 1012 2295
rect 1006 2290 1012 2291
rect 768 2276 770 2290
rect 782 2285 788 2286
rect 782 2281 783 2285
rect 787 2281 788 2285
rect 782 2280 788 2281
rect 686 2275 692 2276
rect 686 2271 687 2275
rect 691 2271 692 2275
rect 686 2270 692 2271
rect 702 2275 708 2276
rect 702 2271 703 2275
rect 707 2271 708 2275
rect 702 2270 708 2271
rect 766 2275 772 2276
rect 766 2271 767 2275
rect 771 2271 772 2275
rect 766 2270 772 2271
rect 111 2258 115 2259
rect 111 2253 115 2254
rect 239 2258 243 2259
rect 239 2253 243 2254
rect 359 2258 363 2259
rect 359 2253 363 2254
rect 391 2258 395 2259
rect 478 2255 479 2259
rect 483 2255 484 2259
rect 478 2254 484 2255
rect 495 2258 499 2259
rect 391 2253 395 2254
rect 495 2253 499 2254
rect 551 2258 555 2259
rect 551 2253 555 2254
rect 639 2258 643 2259
rect 639 2253 643 2254
rect 112 2225 114 2253
rect 240 2244 242 2253
rect 392 2244 394 2253
rect 552 2244 554 2253
rect 238 2243 244 2244
rect 238 2239 239 2243
rect 243 2239 244 2243
rect 238 2238 244 2239
rect 390 2243 396 2244
rect 390 2239 391 2243
rect 395 2239 396 2243
rect 390 2238 396 2239
rect 550 2243 556 2244
rect 550 2239 551 2243
rect 555 2239 556 2243
rect 550 2238 556 2239
rect 704 2236 706 2270
rect 784 2259 786 2280
rect 920 2276 922 2290
rect 934 2285 940 2286
rect 934 2281 935 2285
rect 939 2281 940 2285
rect 934 2280 940 2281
rect 1086 2285 1092 2286
rect 1086 2281 1087 2285
rect 1091 2281 1092 2285
rect 1086 2280 1092 2281
rect 1246 2285 1252 2286
rect 1246 2281 1247 2285
rect 1251 2281 1252 2285
rect 1246 2280 1252 2281
rect 1414 2285 1420 2286
rect 1414 2281 1415 2285
rect 1419 2281 1420 2285
rect 1414 2280 1420 2281
rect 918 2275 924 2276
rect 918 2271 919 2275
rect 923 2271 924 2275
rect 918 2270 924 2271
rect 936 2259 938 2280
rect 1088 2259 1090 2280
rect 1094 2275 1100 2276
rect 1094 2271 1095 2275
rect 1099 2271 1100 2275
rect 1094 2270 1100 2271
rect 711 2258 715 2259
rect 711 2253 715 2254
rect 783 2258 787 2259
rect 783 2253 787 2254
rect 871 2258 875 2259
rect 871 2253 875 2254
rect 935 2258 939 2259
rect 935 2253 939 2254
rect 1031 2258 1035 2259
rect 1031 2253 1035 2254
rect 1087 2258 1091 2259
rect 1087 2253 1091 2254
rect 712 2244 714 2253
rect 872 2244 874 2253
rect 918 2251 924 2252
rect 918 2247 919 2251
rect 923 2247 924 2251
rect 918 2246 924 2247
rect 710 2243 716 2244
rect 710 2239 711 2243
rect 715 2239 716 2243
rect 710 2238 716 2239
rect 870 2243 876 2244
rect 870 2239 871 2243
rect 875 2239 876 2243
rect 870 2238 876 2239
rect 222 2235 228 2236
rect 222 2231 223 2235
rect 227 2231 228 2235
rect 222 2230 228 2231
rect 702 2235 708 2236
rect 702 2231 703 2235
rect 707 2231 708 2235
rect 702 2230 708 2231
rect 110 2224 116 2225
rect 110 2220 111 2224
rect 115 2220 116 2224
rect 110 2219 116 2220
rect 110 2207 116 2208
rect 110 2203 111 2207
rect 115 2203 116 2207
rect 110 2202 116 2203
rect 112 2175 114 2202
rect 111 2174 115 2175
rect 111 2169 115 2170
rect 151 2174 155 2175
rect 151 2169 155 2170
rect 112 2154 114 2169
rect 152 2159 154 2169
rect 150 2158 156 2159
rect 150 2154 151 2158
rect 155 2154 156 2158
rect 110 2153 116 2154
rect 150 2153 156 2154
rect 110 2149 111 2153
rect 115 2149 116 2153
rect 110 2148 116 2149
rect 110 2136 116 2137
rect 110 2132 111 2136
rect 115 2132 116 2136
rect 110 2131 116 2132
rect 112 2095 114 2131
rect 150 2117 156 2118
rect 150 2113 151 2117
rect 155 2113 156 2117
rect 150 2112 156 2113
rect 152 2095 154 2112
rect 224 2108 226 2230
rect 238 2202 244 2203
rect 238 2198 239 2202
rect 243 2198 244 2202
rect 238 2197 244 2198
rect 390 2202 396 2203
rect 390 2198 391 2202
rect 395 2198 396 2202
rect 390 2197 396 2198
rect 550 2202 556 2203
rect 550 2198 551 2202
rect 555 2198 556 2202
rect 550 2197 556 2198
rect 710 2202 716 2203
rect 710 2198 711 2202
rect 715 2198 716 2202
rect 710 2197 716 2198
rect 870 2202 876 2203
rect 870 2198 871 2202
rect 875 2198 876 2202
rect 870 2197 876 2198
rect 240 2175 242 2197
rect 392 2175 394 2197
rect 552 2175 554 2197
rect 712 2175 714 2197
rect 872 2175 874 2197
rect 239 2174 243 2175
rect 239 2169 243 2170
rect 319 2174 323 2175
rect 319 2169 323 2170
rect 391 2174 395 2175
rect 391 2169 395 2170
rect 511 2174 515 2175
rect 511 2169 515 2170
rect 551 2174 555 2175
rect 551 2169 555 2170
rect 703 2174 707 2175
rect 703 2169 707 2170
rect 711 2174 715 2175
rect 711 2169 715 2170
rect 871 2174 875 2175
rect 871 2169 875 2170
rect 895 2174 899 2175
rect 895 2169 899 2170
rect 320 2159 322 2169
rect 512 2159 514 2169
rect 704 2159 706 2169
rect 896 2159 898 2169
rect 318 2158 324 2159
rect 318 2154 319 2158
rect 323 2154 324 2158
rect 318 2153 324 2154
rect 510 2158 516 2159
rect 510 2154 511 2158
rect 515 2154 516 2158
rect 510 2153 516 2154
rect 702 2158 708 2159
rect 702 2154 703 2158
rect 707 2154 708 2158
rect 702 2153 708 2154
rect 894 2158 900 2159
rect 894 2154 895 2158
rect 899 2154 900 2158
rect 894 2153 900 2154
rect 920 2128 922 2246
rect 1032 2244 1034 2253
rect 1030 2243 1036 2244
rect 1030 2239 1031 2243
rect 1035 2239 1036 2243
rect 1030 2238 1036 2239
rect 1096 2236 1098 2270
rect 1248 2259 1250 2280
rect 1416 2259 1418 2280
rect 1528 2276 1530 2390
rect 1534 2366 1540 2367
rect 1534 2362 1535 2366
rect 1539 2362 1540 2366
rect 1534 2361 1540 2362
rect 1670 2366 1676 2367
rect 1670 2362 1671 2366
rect 1675 2362 1676 2366
rect 1670 2361 1676 2362
rect 1814 2366 1820 2367
rect 1814 2362 1815 2366
rect 1819 2362 1820 2366
rect 1814 2361 1820 2362
rect 1934 2366 1940 2367
rect 1934 2362 1935 2366
rect 1939 2362 1940 2366
rect 1934 2361 1940 2362
rect 1536 2343 1538 2361
rect 1672 2343 1674 2361
rect 1816 2343 1818 2361
rect 1936 2343 1938 2361
rect 1535 2342 1539 2343
rect 1535 2337 1539 2338
rect 1591 2342 1595 2343
rect 1591 2337 1595 2338
rect 1671 2342 1675 2343
rect 1671 2337 1675 2338
rect 1775 2342 1779 2343
rect 1775 2337 1779 2338
rect 1815 2342 1819 2343
rect 1815 2337 1819 2338
rect 1935 2342 1939 2343
rect 1935 2337 1939 2338
rect 1592 2327 1594 2337
rect 1776 2327 1778 2337
rect 1936 2327 1938 2337
rect 1590 2326 1596 2327
rect 1590 2322 1591 2326
rect 1595 2322 1596 2326
rect 1590 2321 1596 2322
rect 1774 2326 1780 2327
rect 1774 2322 1775 2326
rect 1779 2322 1780 2326
rect 1774 2321 1780 2322
rect 1934 2326 1940 2327
rect 1934 2322 1935 2326
rect 1939 2322 1940 2326
rect 1934 2321 1940 2322
rect 1574 2295 1580 2296
rect 1574 2291 1575 2295
rect 1579 2291 1580 2295
rect 1574 2290 1580 2291
rect 1758 2295 1764 2296
rect 1758 2291 1759 2295
rect 1763 2291 1764 2295
rect 1758 2290 1764 2291
rect 1766 2295 1772 2296
rect 1766 2291 1767 2295
rect 1771 2291 1772 2295
rect 1766 2290 1772 2291
rect 1576 2276 1578 2290
rect 1590 2285 1596 2286
rect 1590 2281 1591 2285
rect 1595 2281 1596 2285
rect 1590 2280 1596 2281
rect 1526 2275 1532 2276
rect 1526 2271 1527 2275
rect 1531 2271 1532 2275
rect 1526 2270 1532 2271
rect 1574 2275 1580 2276
rect 1574 2271 1575 2275
rect 1579 2271 1580 2275
rect 1574 2270 1580 2271
rect 1592 2259 1594 2280
rect 1760 2276 1762 2290
rect 1758 2275 1764 2276
rect 1758 2271 1759 2275
rect 1763 2271 1764 2275
rect 1758 2270 1764 2271
rect 1191 2258 1195 2259
rect 1191 2253 1195 2254
rect 1247 2258 1251 2259
rect 1247 2253 1251 2254
rect 1359 2258 1363 2259
rect 1359 2253 1363 2254
rect 1415 2258 1419 2259
rect 1415 2253 1419 2254
rect 1527 2258 1531 2259
rect 1527 2253 1531 2254
rect 1591 2258 1595 2259
rect 1591 2253 1595 2254
rect 1695 2258 1699 2259
rect 1695 2253 1699 2254
rect 1192 2244 1194 2253
rect 1360 2244 1362 2253
rect 1406 2251 1412 2252
rect 1406 2247 1407 2251
rect 1411 2247 1412 2251
rect 1406 2246 1412 2247
rect 1190 2243 1196 2244
rect 1190 2239 1191 2243
rect 1195 2239 1196 2243
rect 1190 2238 1196 2239
rect 1358 2243 1364 2244
rect 1358 2239 1359 2243
rect 1363 2239 1364 2243
rect 1358 2238 1364 2239
rect 1094 2235 1100 2236
rect 1094 2231 1095 2235
rect 1099 2231 1100 2235
rect 1094 2230 1100 2231
rect 1030 2202 1036 2203
rect 1030 2198 1031 2202
rect 1035 2198 1036 2202
rect 1030 2197 1036 2198
rect 1190 2202 1196 2203
rect 1190 2198 1191 2202
rect 1195 2198 1196 2202
rect 1190 2197 1196 2198
rect 1358 2202 1364 2203
rect 1358 2198 1359 2202
rect 1363 2198 1364 2202
rect 1358 2197 1364 2198
rect 1032 2175 1034 2197
rect 1192 2175 1194 2197
rect 1360 2175 1362 2197
rect 1031 2174 1035 2175
rect 1031 2169 1035 2170
rect 1087 2174 1091 2175
rect 1087 2169 1091 2170
rect 1191 2174 1195 2175
rect 1191 2169 1195 2170
rect 1279 2174 1283 2175
rect 1279 2169 1283 2170
rect 1359 2174 1363 2175
rect 1359 2169 1363 2170
rect 1088 2159 1090 2169
rect 1280 2159 1282 2169
rect 1086 2158 1092 2159
rect 1086 2154 1087 2158
rect 1091 2154 1092 2158
rect 1086 2153 1092 2154
rect 1278 2158 1284 2159
rect 1278 2154 1279 2158
rect 1283 2154 1284 2158
rect 1278 2153 1284 2154
rect 1408 2128 1410 2246
rect 1528 2244 1530 2253
rect 1696 2244 1698 2253
rect 1768 2252 1770 2290
rect 1774 2285 1780 2286
rect 1774 2281 1775 2285
rect 1779 2281 1780 2285
rect 1774 2280 1780 2281
rect 1934 2285 1940 2286
rect 1934 2281 1935 2285
rect 1939 2281 1940 2285
rect 1934 2280 1940 2281
rect 1776 2259 1778 2280
rect 1936 2259 1938 2280
rect 2008 2276 2010 2394
rect 2032 2389 2034 2417
rect 2072 2407 2074 2447
rect 2540 2444 2542 2562
rect 2616 2560 2618 2569
rect 2614 2559 2620 2560
rect 2614 2555 2615 2559
rect 2619 2555 2620 2559
rect 2614 2554 2620 2555
rect 2684 2552 2686 2582
rect 2752 2575 2754 2592
rect 2896 2575 2898 2592
rect 3024 2576 3026 2602
rect 3038 2597 3044 2598
rect 3128 2597 3130 2710
rect 3992 2705 3994 2733
rect 3990 2704 3996 2705
rect 3990 2700 3991 2704
rect 3995 2700 3996 2704
rect 3990 2699 3996 2700
rect 3990 2687 3996 2688
rect 3990 2683 3991 2687
rect 3995 2683 3996 2687
rect 3142 2682 3148 2683
rect 3142 2678 3143 2682
rect 3147 2678 3148 2682
rect 3142 2677 3148 2678
rect 3302 2682 3308 2683
rect 3302 2678 3303 2682
rect 3307 2678 3308 2682
rect 3302 2677 3308 2678
rect 3462 2682 3468 2683
rect 3462 2678 3463 2682
rect 3467 2678 3468 2682
rect 3462 2677 3468 2678
rect 3622 2682 3628 2683
rect 3990 2682 3996 2683
rect 3622 2678 3623 2682
rect 3627 2678 3628 2682
rect 3622 2677 3628 2678
rect 3144 2655 3146 2677
rect 3304 2655 3306 2677
rect 3464 2655 3466 2677
rect 3624 2655 3626 2677
rect 3992 2655 3994 2682
rect 3143 2654 3147 2655
rect 3143 2649 3147 2650
rect 3175 2654 3179 2655
rect 3175 2649 3179 2650
rect 3303 2654 3307 2655
rect 3303 2649 3307 2650
rect 3311 2654 3315 2655
rect 3311 2649 3315 2650
rect 3455 2654 3459 2655
rect 3455 2649 3459 2650
rect 3463 2654 3467 2655
rect 3463 2649 3467 2650
rect 3623 2654 3627 2655
rect 3623 2649 3627 2650
rect 3991 2654 3995 2655
rect 3991 2649 3995 2650
rect 3176 2639 3178 2649
rect 3312 2639 3314 2649
rect 3456 2639 3458 2649
rect 3174 2638 3180 2639
rect 3174 2634 3175 2638
rect 3179 2634 3180 2638
rect 3174 2633 3180 2634
rect 3310 2638 3316 2639
rect 3310 2634 3311 2638
rect 3315 2634 3316 2638
rect 3310 2633 3316 2634
rect 3454 2638 3460 2639
rect 3454 2634 3455 2638
rect 3459 2634 3460 2638
rect 3992 2634 3994 2649
rect 3454 2633 3460 2634
rect 3990 2633 3996 2634
rect 3990 2629 3991 2633
rect 3995 2629 3996 2633
rect 3990 2628 3996 2629
rect 3990 2616 3996 2617
rect 3990 2612 3991 2616
rect 3995 2612 3996 2616
rect 3990 2611 3996 2612
rect 3174 2597 3180 2598
rect 3038 2593 3039 2597
rect 3043 2593 3044 2597
rect 3038 2592 3044 2593
rect 3127 2596 3131 2597
rect 3174 2593 3175 2597
rect 3179 2593 3180 2597
rect 3174 2592 3180 2593
rect 3310 2597 3316 2598
rect 3310 2593 3311 2597
rect 3315 2593 3316 2597
rect 3310 2592 3316 2593
rect 3454 2597 3460 2598
rect 3454 2593 3455 2597
rect 3459 2593 3460 2597
rect 3454 2592 3460 2593
rect 3527 2596 3531 2597
rect 3022 2575 3028 2576
rect 3040 2575 3042 2592
rect 3127 2591 3131 2592
rect 3176 2575 3178 2592
rect 3312 2575 3314 2592
rect 3456 2575 3458 2592
rect 3527 2591 3531 2592
rect 3528 2588 3530 2591
rect 3526 2587 3532 2588
rect 3526 2583 3527 2587
rect 3531 2583 3532 2587
rect 3526 2582 3532 2583
rect 3992 2575 3994 2611
rect 2751 2574 2755 2575
rect 2751 2569 2755 2570
rect 2767 2574 2771 2575
rect 2767 2569 2771 2570
rect 2895 2574 2899 2575
rect 2895 2569 2899 2570
rect 2911 2574 2915 2575
rect 3022 2571 3023 2575
rect 3027 2571 3028 2575
rect 3022 2570 3028 2571
rect 3039 2574 3043 2575
rect 2911 2569 2915 2570
rect 3039 2569 3043 2570
rect 3047 2574 3051 2575
rect 3047 2569 3051 2570
rect 3175 2574 3179 2575
rect 3175 2569 3179 2570
rect 3183 2574 3187 2575
rect 3183 2569 3187 2570
rect 3311 2574 3315 2575
rect 3311 2569 3315 2570
rect 3319 2574 3323 2575
rect 3319 2569 3323 2570
rect 3455 2574 3459 2575
rect 3455 2569 3459 2570
rect 3991 2574 3995 2575
rect 3991 2569 3995 2570
rect 2768 2560 2770 2569
rect 2912 2560 2914 2569
rect 3048 2560 3050 2569
rect 3184 2560 3186 2569
rect 3320 2560 3322 2569
rect 2766 2559 2772 2560
rect 2766 2555 2767 2559
rect 2771 2555 2772 2559
rect 2766 2554 2772 2555
rect 2910 2559 2916 2560
rect 2910 2555 2911 2559
rect 2915 2555 2916 2559
rect 2910 2554 2916 2555
rect 3046 2559 3052 2560
rect 3046 2555 3047 2559
rect 3051 2555 3052 2559
rect 3046 2554 3052 2555
rect 3182 2559 3188 2560
rect 3182 2555 3183 2559
rect 3187 2555 3188 2559
rect 3182 2554 3188 2555
rect 3318 2559 3324 2560
rect 3318 2555 3319 2559
rect 3323 2555 3324 2559
rect 3318 2554 3324 2555
rect 2682 2551 2688 2552
rect 2682 2547 2683 2551
rect 2687 2547 2688 2551
rect 2682 2546 2688 2547
rect 2894 2551 2900 2552
rect 2894 2547 2895 2551
rect 2899 2547 2900 2551
rect 2894 2546 2900 2547
rect 2614 2518 2620 2519
rect 2614 2514 2615 2518
rect 2619 2514 2620 2518
rect 2614 2513 2620 2514
rect 2766 2518 2772 2519
rect 2766 2514 2767 2518
rect 2771 2514 2772 2518
rect 2766 2513 2772 2514
rect 2616 2491 2618 2513
rect 2768 2491 2770 2513
rect 2615 2490 2619 2491
rect 2615 2485 2619 2486
rect 2623 2490 2627 2491
rect 2623 2485 2627 2486
rect 2743 2490 2747 2491
rect 2743 2485 2747 2486
rect 2767 2490 2771 2491
rect 2767 2485 2771 2486
rect 2871 2490 2875 2491
rect 2871 2485 2875 2486
rect 2624 2475 2626 2485
rect 2744 2475 2746 2485
rect 2872 2475 2874 2485
rect 2622 2474 2628 2475
rect 2622 2470 2623 2474
rect 2627 2470 2628 2474
rect 2622 2469 2628 2470
rect 2742 2474 2748 2475
rect 2742 2470 2743 2474
rect 2747 2470 2748 2474
rect 2742 2469 2748 2470
rect 2870 2474 2876 2475
rect 2870 2470 2871 2474
rect 2875 2470 2876 2474
rect 2870 2469 2876 2470
rect 2538 2443 2544 2444
rect 2538 2439 2539 2443
rect 2543 2439 2544 2443
rect 2538 2438 2544 2439
rect 2622 2433 2628 2434
rect 2622 2429 2623 2433
rect 2627 2429 2628 2433
rect 2622 2428 2628 2429
rect 2742 2433 2748 2434
rect 2742 2429 2743 2433
rect 2747 2429 2748 2433
rect 2742 2428 2748 2429
rect 2870 2433 2876 2434
rect 2870 2429 2871 2433
rect 2875 2429 2876 2433
rect 2870 2428 2876 2429
rect 2582 2407 2588 2408
rect 2624 2407 2626 2428
rect 2744 2407 2746 2428
rect 2790 2423 2796 2424
rect 2790 2419 2791 2423
rect 2795 2419 2796 2423
rect 2790 2418 2796 2419
rect 2071 2406 2075 2407
rect 2071 2401 2075 2402
rect 2487 2406 2491 2407
rect 2582 2403 2583 2407
rect 2587 2403 2588 2407
rect 2582 2402 2588 2403
rect 2599 2406 2603 2407
rect 2487 2401 2491 2402
rect 2030 2388 2036 2389
rect 2030 2384 2031 2388
rect 2035 2384 2036 2388
rect 2030 2383 2036 2384
rect 2072 2373 2074 2401
rect 2488 2392 2490 2401
rect 2486 2391 2492 2392
rect 2486 2387 2487 2391
rect 2491 2387 2492 2391
rect 2486 2386 2492 2387
rect 2584 2384 2586 2402
rect 2599 2401 2603 2402
rect 2623 2406 2627 2407
rect 2623 2401 2627 2402
rect 2727 2406 2731 2407
rect 2727 2401 2731 2402
rect 2743 2406 2747 2407
rect 2743 2401 2747 2402
rect 2600 2392 2602 2401
rect 2662 2399 2668 2400
rect 2662 2395 2663 2399
rect 2667 2395 2668 2399
rect 2662 2394 2668 2395
rect 2598 2391 2604 2392
rect 2598 2387 2599 2391
rect 2603 2387 2604 2391
rect 2598 2386 2604 2387
rect 2582 2383 2588 2384
rect 2582 2379 2583 2383
rect 2587 2379 2588 2383
rect 2582 2378 2588 2379
rect 2070 2372 2076 2373
rect 2030 2371 2036 2372
rect 2030 2367 2031 2371
rect 2035 2367 2036 2371
rect 2070 2368 2071 2372
rect 2075 2368 2076 2372
rect 2070 2367 2076 2368
rect 2030 2366 2036 2367
rect 2032 2343 2034 2366
rect 2070 2355 2076 2356
rect 2070 2351 2071 2355
rect 2075 2351 2076 2355
rect 2070 2350 2076 2351
rect 2486 2350 2492 2351
rect 2031 2342 2035 2343
rect 2031 2337 2035 2338
rect 2032 2322 2034 2337
rect 2072 2323 2074 2350
rect 2486 2346 2487 2350
rect 2491 2346 2492 2350
rect 2486 2345 2492 2346
rect 2598 2350 2604 2351
rect 2598 2346 2599 2350
rect 2603 2346 2604 2350
rect 2598 2345 2604 2346
rect 2488 2323 2490 2345
rect 2600 2323 2602 2345
rect 2071 2322 2075 2323
rect 2030 2321 2036 2322
rect 2030 2317 2031 2321
rect 2035 2317 2036 2321
rect 2071 2317 2075 2318
rect 2111 2322 2115 2323
rect 2111 2317 2115 2318
rect 2223 2322 2227 2323
rect 2223 2317 2227 2318
rect 2359 2322 2363 2323
rect 2359 2317 2363 2318
rect 2487 2322 2491 2323
rect 2487 2317 2491 2318
rect 2511 2322 2515 2323
rect 2511 2317 2515 2318
rect 2599 2322 2603 2323
rect 2599 2317 2603 2318
rect 2030 2316 2036 2317
rect 2030 2304 2036 2305
rect 2030 2300 2031 2304
rect 2035 2300 2036 2304
rect 2072 2302 2074 2317
rect 2112 2307 2114 2317
rect 2224 2307 2226 2317
rect 2360 2307 2362 2317
rect 2512 2307 2514 2317
rect 2110 2306 2116 2307
rect 2110 2302 2111 2306
rect 2115 2302 2116 2306
rect 2030 2299 2036 2300
rect 2070 2301 2076 2302
rect 2110 2301 2116 2302
rect 2222 2306 2228 2307
rect 2222 2302 2223 2306
rect 2227 2302 2228 2306
rect 2222 2301 2228 2302
rect 2358 2306 2364 2307
rect 2358 2302 2359 2306
rect 2363 2302 2364 2306
rect 2358 2301 2364 2302
rect 2510 2306 2516 2307
rect 2510 2302 2511 2306
rect 2515 2302 2516 2306
rect 2510 2301 2516 2302
rect 2006 2275 2012 2276
rect 2006 2271 2007 2275
rect 2011 2271 2012 2275
rect 2006 2270 2012 2271
rect 2032 2259 2034 2299
rect 2070 2297 2071 2301
rect 2075 2297 2076 2301
rect 2070 2296 2076 2297
rect 2182 2295 2188 2296
rect 2182 2291 2183 2295
rect 2187 2291 2188 2295
rect 2182 2290 2188 2291
rect 2070 2284 2076 2285
rect 2070 2280 2071 2284
rect 2075 2280 2076 2284
rect 2070 2279 2076 2280
rect 1775 2258 1779 2259
rect 1775 2253 1779 2254
rect 1935 2258 1939 2259
rect 1935 2253 1939 2254
rect 2031 2258 2035 2259
rect 2031 2253 2035 2254
rect 1766 2251 1772 2252
rect 1766 2247 1767 2251
rect 1771 2247 1772 2251
rect 1766 2246 1772 2247
rect 1526 2243 1532 2244
rect 1526 2239 1527 2243
rect 1531 2239 1532 2243
rect 1526 2238 1532 2239
rect 1694 2243 1700 2244
rect 1694 2239 1695 2243
rect 1699 2239 1700 2243
rect 1694 2238 1700 2239
rect 1534 2231 1540 2232
rect 1534 2227 1535 2231
rect 1539 2227 1540 2231
rect 1534 2226 1540 2227
rect 1526 2202 1532 2203
rect 1526 2198 1527 2202
rect 1531 2198 1532 2202
rect 1526 2197 1532 2198
rect 1528 2175 1530 2197
rect 1463 2174 1467 2175
rect 1463 2169 1467 2170
rect 1527 2174 1531 2175
rect 1527 2169 1531 2170
rect 1464 2159 1466 2169
rect 1462 2158 1468 2159
rect 1462 2154 1463 2158
rect 1467 2154 1468 2158
rect 1462 2153 1468 2154
rect 238 2127 244 2128
rect 238 2123 239 2127
rect 243 2123 244 2127
rect 238 2122 244 2123
rect 450 2127 456 2128
rect 450 2123 451 2127
rect 455 2123 456 2127
rect 450 2122 456 2123
rect 534 2127 540 2128
rect 534 2123 535 2127
rect 539 2123 540 2127
rect 534 2122 540 2123
rect 878 2127 884 2128
rect 878 2123 879 2127
rect 883 2123 884 2127
rect 878 2122 884 2123
rect 918 2127 924 2128
rect 918 2123 919 2127
rect 923 2123 924 2127
rect 918 2122 924 2123
rect 1406 2127 1412 2128
rect 1406 2123 1407 2127
rect 1411 2123 1412 2127
rect 1406 2122 1412 2123
rect 240 2108 242 2122
rect 318 2117 324 2118
rect 318 2113 319 2117
rect 323 2113 324 2117
rect 318 2112 324 2113
rect 222 2107 228 2108
rect 222 2103 223 2107
rect 227 2103 228 2107
rect 222 2102 228 2103
rect 238 2107 244 2108
rect 238 2103 239 2107
rect 243 2103 244 2107
rect 238 2102 244 2103
rect 320 2095 322 2112
rect 452 2108 454 2122
rect 510 2117 516 2118
rect 510 2113 511 2117
rect 515 2113 516 2117
rect 510 2112 516 2113
rect 450 2107 456 2108
rect 450 2103 451 2107
rect 455 2103 456 2107
rect 450 2102 456 2103
rect 512 2095 514 2112
rect 111 2094 115 2095
rect 111 2089 115 2090
rect 151 2094 155 2095
rect 151 2089 155 2090
rect 303 2094 307 2095
rect 303 2089 307 2090
rect 319 2094 323 2095
rect 319 2089 323 2090
rect 479 2094 483 2095
rect 479 2089 483 2090
rect 511 2094 515 2095
rect 511 2089 515 2090
rect 112 2061 114 2089
rect 152 2080 154 2089
rect 304 2080 306 2089
rect 480 2080 482 2089
rect 536 2088 538 2122
rect 702 2117 708 2118
rect 702 2113 703 2117
rect 707 2113 708 2117
rect 702 2112 708 2113
rect 704 2095 706 2112
rect 880 2108 882 2122
rect 894 2117 900 2118
rect 894 2113 895 2117
rect 899 2113 900 2117
rect 894 2112 900 2113
rect 1086 2117 1092 2118
rect 1086 2113 1087 2117
rect 1091 2113 1092 2117
rect 1086 2112 1092 2113
rect 1278 2117 1284 2118
rect 1278 2113 1279 2117
rect 1283 2113 1284 2117
rect 1278 2112 1284 2113
rect 1462 2117 1468 2118
rect 1462 2113 1463 2117
rect 1467 2113 1468 2117
rect 1462 2112 1468 2113
rect 726 2107 732 2108
rect 726 2103 727 2107
rect 731 2103 732 2107
rect 726 2102 732 2103
rect 878 2107 884 2108
rect 878 2103 879 2107
rect 883 2103 884 2107
rect 878 2102 884 2103
rect 663 2094 667 2095
rect 663 2089 667 2090
rect 703 2094 707 2095
rect 703 2089 707 2090
rect 534 2087 540 2088
rect 534 2083 535 2087
rect 539 2083 540 2087
rect 534 2082 540 2083
rect 664 2080 666 2089
rect 150 2079 156 2080
rect 150 2075 151 2079
rect 155 2075 156 2079
rect 150 2074 156 2075
rect 302 2079 308 2080
rect 302 2075 303 2079
rect 307 2075 308 2079
rect 302 2074 308 2075
rect 478 2079 484 2080
rect 478 2075 479 2079
rect 483 2075 484 2079
rect 478 2074 484 2075
rect 662 2079 668 2080
rect 662 2075 663 2079
rect 667 2075 668 2079
rect 662 2074 668 2075
rect 728 2072 730 2102
rect 896 2095 898 2112
rect 1088 2095 1090 2112
rect 1114 2107 1120 2108
rect 1114 2103 1115 2107
rect 1119 2103 1120 2107
rect 1114 2102 1120 2103
rect 847 2094 851 2095
rect 847 2089 851 2090
rect 895 2094 899 2095
rect 895 2089 899 2090
rect 1039 2094 1043 2095
rect 1039 2089 1043 2090
rect 1087 2094 1091 2095
rect 1087 2089 1091 2090
rect 848 2080 850 2089
rect 918 2087 924 2088
rect 918 2083 919 2087
rect 923 2083 924 2087
rect 918 2082 924 2083
rect 846 2079 852 2080
rect 846 2075 847 2079
rect 851 2075 852 2079
rect 846 2074 852 2075
rect 222 2071 228 2072
rect 222 2067 223 2071
rect 227 2067 228 2071
rect 222 2066 228 2067
rect 726 2071 732 2072
rect 726 2067 727 2071
rect 731 2067 732 2071
rect 726 2066 732 2067
rect 110 2060 116 2061
rect 110 2056 111 2060
rect 115 2056 116 2060
rect 110 2055 116 2056
rect 110 2043 116 2044
rect 110 2039 111 2043
rect 115 2039 116 2043
rect 110 2038 116 2039
rect 150 2038 156 2039
rect 112 2015 114 2038
rect 150 2034 151 2038
rect 155 2034 156 2038
rect 150 2033 156 2034
rect 152 2015 154 2033
rect 111 2014 115 2015
rect 111 2009 115 2010
rect 151 2014 155 2015
rect 151 2009 155 2010
rect 112 1994 114 2009
rect 152 1999 154 2009
rect 150 1998 156 1999
rect 150 1994 151 1998
rect 155 1994 156 1998
rect 110 1993 116 1994
rect 150 1993 156 1994
rect 110 1989 111 1993
rect 115 1989 116 1993
rect 110 1988 116 1989
rect 110 1976 116 1977
rect 110 1972 111 1976
rect 115 1972 116 1976
rect 110 1971 116 1972
rect 112 1931 114 1971
rect 150 1957 156 1958
rect 150 1953 151 1957
rect 155 1953 156 1957
rect 150 1952 156 1953
rect 152 1931 154 1952
rect 224 1948 226 2066
rect 302 2038 308 2039
rect 302 2034 303 2038
rect 307 2034 308 2038
rect 302 2033 308 2034
rect 478 2038 484 2039
rect 478 2034 479 2038
rect 483 2034 484 2038
rect 478 2033 484 2034
rect 662 2038 668 2039
rect 662 2034 663 2038
rect 667 2034 668 2038
rect 662 2033 668 2034
rect 846 2038 852 2039
rect 846 2034 847 2038
rect 851 2034 852 2038
rect 846 2033 852 2034
rect 304 2015 306 2033
rect 480 2015 482 2033
rect 664 2015 666 2033
rect 848 2015 850 2033
rect 303 2014 307 2015
rect 303 2009 307 2010
rect 479 2014 483 2015
rect 479 2009 483 2010
rect 487 2014 491 2015
rect 487 2009 491 2010
rect 663 2014 667 2015
rect 663 2009 667 2010
rect 687 2014 691 2015
rect 687 2009 691 2010
rect 847 2014 851 2015
rect 847 2009 851 2010
rect 895 2014 899 2015
rect 895 2009 899 2010
rect 304 1999 306 2009
rect 488 1999 490 2009
rect 688 1999 690 2009
rect 896 1999 898 2009
rect 302 1998 308 1999
rect 302 1994 303 1998
rect 307 1994 308 1998
rect 302 1993 308 1994
rect 486 1998 492 1999
rect 486 1994 487 1998
rect 491 1994 492 1998
rect 486 1993 492 1994
rect 686 1998 692 1999
rect 686 1994 687 1998
rect 691 1994 692 1998
rect 686 1993 692 1994
rect 894 1998 900 1999
rect 894 1994 895 1998
rect 899 1994 900 1998
rect 894 1993 900 1994
rect 920 1968 922 2082
rect 1040 2080 1042 2089
rect 1038 2079 1044 2080
rect 1038 2075 1039 2079
rect 1043 2075 1044 2079
rect 1038 2074 1044 2075
rect 1116 2072 1118 2102
rect 1280 2095 1282 2112
rect 1464 2095 1466 2112
rect 1536 2108 1538 2226
rect 2032 2225 2034 2253
rect 2072 2243 2074 2279
rect 2110 2265 2116 2266
rect 2110 2261 2111 2265
rect 2115 2261 2116 2265
rect 2110 2260 2116 2261
rect 2112 2243 2114 2260
rect 2184 2256 2186 2290
rect 2664 2276 2666 2394
rect 2728 2392 2730 2401
rect 2726 2391 2732 2392
rect 2726 2387 2727 2391
rect 2731 2387 2732 2391
rect 2726 2386 2732 2387
rect 2792 2384 2794 2418
rect 2872 2407 2874 2428
rect 2896 2416 2898 2546
rect 3992 2541 3994 2569
rect 3990 2540 3996 2541
rect 3990 2536 3991 2540
rect 3995 2536 3996 2540
rect 3990 2535 3996 2536
rect 3990 2523 3996 2524
rect 3990 2519 3991 2523
rect 3995 2519 3996 2523
rect 2910 2518 2916 2519
rect 2910 2514 2911 2518
rect 2915 2514 2916 2518
rect 2910 2513 2916 2514
rect 3046 2518 3052 2519
rect 3046 2514 3047 2518
rect 3051 2514 3052 2518
rect 3046 2513 3052 2514
rect 3182 2518 3188 2519
rect 3182 2514 3183 2518
rect 3187 2514 3188 2518
rect 3182 2513 3188 2514
rect 3318 2518 3324 2519
rect 3990 2518 3996 2519
rect 3318 2514 3319 2518
rect 3323 2514 3324 2518
rect 3318 2513 3324 2514
rect 2912 2491 2914 2513
rect 3048 2491 3050 2513
rect 3184 2491 3186 2513
rect 3320 2491 3322 2513
rect 3992 2491 3994 2518
rect 2911 2490 2915 2491
rect 2911 2485 2915 2486
rect 3015 2490 3019 2491
rect 3015 2485 3019 2486
rect 3047 2490 3051 2491
rect 3047 2485 3051 2486
rect 3159 2490 3163 2491
rect 3159 2485 3163 2486
rect 3183 2490 3187 2491
rect 3183 2485 3187 2486
rect 3311 2490 3315 2491
rect 3311 2485 3315 2486
rect 3319 2490 3323 2491
rect 3319 2485 3323 2486
rect 3463 2490 3467 2491
rect 3463 2485 3467 2486
rect 3615 2490 3619 2491
rect 3615 2485 3619 2486
rect 3767 2490 3771 2491
rect 3767 2485 3771 2486
rect 3895 2490 3899 2491
rect 3895 2485 3899 2486
rect 3991 2490 3995 2491
rect 3991 2485 3995 2486
rect 3016 2475 3018 2485
rect 3160 2475 3162 2485
rect 3312 2475 3314 2485
rect 3464 2475 3466 2485
rect 3616 2475 3618 2485
rect 3768 2475 3770 2485
rect 3896 2475 3898 2485
rect 3014 2474 3020 2475
rect 3014 2470 3015 2474
rect 3019 2470 3020 2474
rect 3014 2469 3020 2470
rect 3158 2474 3164 2475
rect 3158 2470 3159 2474
rect 3163 2470 3164 2474
rect 3158 2469 3164 2470
rect 3310 2474 3316 2475
rect 3310 2470 3311 2474
rect 3315 2470 3316 2474
rect 3310 2469 3316 2470
rect 3462 2474 3468 2475
rect 3462 2470 3463 2474
rect 3467 2470 3468 2474
rect 3462 2469 3468 2470
rect 3614 2474 3620 2475
rect 3614 2470 3615 2474
rect 3619 2470 3620 2474
rect 3614 2469 3620 2470
rect 3766 2474 3772 2475
rect 3766 2470 3767 2474
rect 3771 2470 3772 2474
rect 3766 2469 3772 2470
rect 3894 2474 3900 2475
rect 3894 2470 3895 2474
rect 3899 2470 3900 2474
rect 3992 2470 3994 2485
rect 3894 2469 3900 2470
rect 3990 2469 3996 2470
rect 3990 2465 3991 2469
rect 3995 2465 3996 2469
rect 3990 2464 3996 2465
rect 3990 2452 3996 2453
rect 3990 2448 3991 2452
rect 3995 2448 3996 2452
rect 3990 2447 3996 2448
rect 2942 2443 2948 2444
rect 2942 2439 2943 2443
rect 2947 2439 2948 2443
rect 2942 2438 2948 2439
rect 3566 2443 3572 2444
rect 3566 2439 3567 2443
rect 3571 2439 3572 2443
rect 3566 2438 3572 2439
rect 3878 2443 3884 2444
rect 3878 2439 3879 2443
rect 3883 2439 3884 2443
rect 3878 2438 3884 2439
rect 3966 2443 3972 2444
rect 3966 2439 3967 2443
rect 3971 2439 3972 2443
rect 3966 2438 3972 2439
rect 2894 2415 2900 2416
rect 2894 2411 2895 2415
rect 2899 2411 2900 2415
rect 2894 2410 2900 2411
rect 2871 2406 2875 2407
rect 2871 2401 2875 2402
rect 2879 2406 2883 2407
rect 2879 2401 2883 2402
rect 2880 2392 2882 2401
rect 2944 2400 2946 2438
rect 3014 2433 3020 2434
rect 3014 2429 3015 2433
rect 3019 2429 3020 2433
rect 3014 2428 3020 2429
rect 3158 2433 3164 2434
rect 3158 2429 3159 2433
rect 3163 2429 3164 2433
rect 3158 2428 3164 2429
rect 3310 2433 3316 2434
rect 3310 2429 3311 2433
rect 3315 2429 3316 2433
rect 3310 2428 3316 2429
rect 3462 2433 3468 2434
rect 3462 2429 3463 2433
rect 3467 2429 3468 2433
rect 3462 2428 3468 2429
rect 3016 2407 3018 2428
rect 3038 2407 3044 2408
rect 3160 2407 3162 2428
rect 3312 2407 3314 2428
rect 3464 2407 3466 2428
rect 3568 2416 3570 2438
rect 3614 2433 3620 2434
rect 3614 2429 3615 2433
rect 3619 2429 3620 2433
rect 3614 2428 3620 2429
rect 3766 2433 3772 2434
rect 3766 2429 3767 2433
rect 3771 2429 3772 2433
rect 3766 2428 3772 2429
rect 3566 2415 3572 2416
rect 3566 2411 3567 2415
rect 3571 2411 3572 2415
rect 3566 2410 3572 2411
rect 3616 2407 3618 2428
rect 3686 2423 3692 2424
rect 3686 2419 3687 2423
rect 3691 2419 3692 2423
rect 3686 2418 3692 2419
rect 3015 2406 3019 2407
rect 3038 2403 3039 2407
rect 3043 2403 3044 2407
rect 3038 2402 3044 2403
rect 3055 2406 3059 2407
rect 3015 2401 3019 2402
rect 2942 2399 2948 2400
rect 2942 2395 2943 2399
rect 2947 2395 2948 2399
rect 2942 2394 2948 2395
rect 2878 2391 2884 2392
rect 2878 2387 2879 2391
rect 2883 2387 2884 2391
rect 2878 2386 2884 2387
rect 3040 2384 3042 2402
rect 3055 2401 3059 2402
rect 3159 2406 3163 2407
rect 3159 2401 3163 2402
rect 3247 2406 3251 2407
rect 3247 2401 3251 2402
rect 3311 2406 3315 2407
rect 3311 2401 3315 2402
rect 3455 2406 3459 2407
rect 3455 2401 3459 2402
rect 3463 2406 3467 2407
rect 3463 2401 3467 2402
rect 3615 2406 3619 2407
rect 3615 2401 3619 2402
rect 3679 2406 3683 2407
rect 3679 2401 3683 2402
rect 3056 2392 3058 2401
rect 3248 2392 3250 2401
rect 3456 2392 3458 2401
rect 3680 2392 3682 2401
rect 3054 2391 3060 2392
rect 3054 2387 3055 2391
rect 3059 2387 3060 2391
rect 3054 2386 3060 2387
rect 3246 2391 3252 2392
rect 3246 2387 3247 2391
rect 3251 2387 3252 2391
rect 3246 2386 3252 2387
rect 3454 2391 3460 2392
rect 3454 2387 3455 2391
rect 3459 2387 3460 2391
rect 3454 2386 3460 2387
rect 3678 2391 3684 2392
rect 3678 2387 3679 2391
rect 3683 2387 3684 2391
rect 3678 2386 3684 2387
rect 2790 2383 2796 2384
rect 2790 2379 2791 2383
rect 2795 2379 2796 2383
rect 2790 2378 2796 2379
rect 3038 2383 3044 2384
rect 3038 2379 3039 2383
rect 3043 2379 3044 2383
rect 3038 2378 3044 2379
rect 3118 2383 3124 2384
rect 3118 2379 3119 2383
rect 3123 2379 3124 2383
rect 3688 2380 3690 2418
rect 3768 2407 3770 2428
rect 3880 2424 3882 2438
rect 3894 2433 3900 2434
rect 3894 2429 3895 2433
rect 3899 2429 3900 2433
rect 3894 2428 3900 2429
rect 3878 2423 3884 2424
rect 3878 2419 3879 2423
rect 3883 2419 3884 2423
rect 3878 2418 3884 2419
rect 3896 2407 3898 2428
rect 3767 2406 3771 2407
rect 3767 2401 3771 2402
rect 3895 2406 3899 2407
rect 3895 2401 3899 2402
rect 3896 2392 3898 2401
rect 3968 2400 3970 2438
rect 3992 2407 3994 2447
rect 3991 2406 3995 2407
rect 3991 2401 3995 2402
rect 3966 2399 3972 2400
rect 3966 2395 3967 2399
rect 3971 2395 3972 2399
rect 3966 2394 3972 2395
rect 3894 2391 3900 2392
rect 3894 2387 3895 2391
rect 3899 2387 3900 2391
rect 3894 2386 3900 2387
rect 3958 2383 3964 2384
rect 3118 2378 3124 2379
rect 3686 2379 3692 2380
rect 2726 2350 2732 2351
rect 2726 2346 2727 2350
rect 2731 2346 2732 2350
rect 2726 2345 2732 2346
rect 2878 2350 2884 2351
rect 2878 2346 2879 2350
rect 2883 2346 2884 2350
rect 2878 2345 2884 2346
rect 3054 2350 3060 2351
rect 3054 2346 3055 2350
rect 3059 2346 3060 2350
rect 3054 2345 3060 2346
rect 2728 2323 2730 2345
rect 2880 2323 2882 2345
rect 3056 2323 3058 2345
rect 2671 2322 2675 2323
rect 2671 2317 2675 2318
rect 2727 2322 2731 2323
rect 2727 2317 2731 2318
rect 2847 2322 2851 2323
rect 2847 2317 2851 2318
rect 2879 2322 2883 2323
rect 2879 2317 2883 2318
rect 3039 2322 3043 2323
rect 3039 2317 3043 2318
rect 3055 2322 3059 2323
rect 3055 2317 3059 2318
rect 2672 2307 2674 2317
rect 2848 2307 2850 2317
rect 3040 2307 3042 2317
rect 2670 2306 2676 2307
rect 2670 2302 2671 2306
rect 2675 2302 2676 2306
rect 2670 2301 2676 2302
rect 2846 2306 2852 2307
rect 2846 2302 2847 2306
rect 2851 2302 2852 2306
rect 2846 2301 2852 2302
rect 3038 2306 3044 2307
rect 3038 2302 3039 2306
rect 3043 2302 3044 2306
rect 3038 2301 3044 2302
rect 2494 2275 2500 2276
rect 2494 2271 2495 2275
rect 2499 2271 2500 2275
rect 2494 2270 2500 2271
rect 2654 2275 2660 2276
rect 2654 2271 2655 2275
rect 2659 2271 2660 2275
rect 2654 2270 2660 2271
rect 2662 2275 2668 2276
rect 2662 2271 2663 2275
rect 2667 2271 2668 2275
rect 2662 2270 2668 2271
rect 3022 2275 3028 2276
rect 3022 2271 3023 2275
rect 3027 2271 3028 2275
rect 3022 2270 3028 2271
rect 2222 2265 2228 2266
rect 2222 2261 2223 2265
rect 2227 2261 2228 2265
rect 2222 2260 2228 2261
rect 2358 2265 2364 2266
rect 2358 2261 2359 2265
rect 2363 2261 2364 2265
rect 2358 2260 2364 2261
rect 2182 2255 2188 2256
rect 2182 2251 2183 2255
rect 2187 2251 2188 2255
rect 2182 2250 2188 2251
rect 2224 2243 2226 2260
rect 2360 2243 2362 2260
rect 2496 2256 2498 2270
rect 2510 2265 2516 2266
rect 2510 2261 2511 2265
rect 2515 2261 2516 2265
rect 2510 2260 2516 2261
rect 2434 2255 2440 2256
rect 2434 2251 2435 2255
rect 2439 2251 2440 2255
rect 2434 2250 2440 2251
rect 2494 2255 2500 2256
rect 2494 2251 2495 2255
rect 2499 2251 2500 2255
rect 2494 2250 2500 2251
rect 2071 2242 2075 2243
rect 2071 2237 2075 2238
rect 2111 2242 2115 2243
rect 2111 2237 2115 2238
rect 2223 2242 2227 2243
rect 2223 2237 2227 2238
rect 2279 2242 2283 2243
rect 2279 2237 2283 2238
rect 2359 2242 2363 2243
rect 2359 2237 2363 2238
rect 2030 2224 2036 2225
rect 2030 2220 2031 2224
rect 2035 2220 2036 2224
rect 2030 2219 2036 2220
rect 2072 2209 2074 2237
rect 2112 2228 2114 2237
rect 2280 2228 2282 2237
rect 2436 2236 2438 2250
rect 2512 2243 2514 2260
rect 2656 2256 2658 2270
rect 2670 2265 2676 2266
rect 2670 2261 2671 2265
rect 2675 2261 2676 2265
rect 2670 2260 2676 2261
rect 2846 2265 2852 2266
rect 2846 2261 2847 2265
rect 2851 2261 2852 2265
rect 2846 2260 2852 2261
rect 2654 2255 2660 2256
rect 2654 2251 2655 2255
rect 2659 2251 2660 2255
rect 2654 2250 2660 2251
rect 2672 2243 2674 2260
rect 2848 2243 2850 2260
rect 3024 2248 3026 2270
rect 3038 2265 3044 2266
rect 3038 2261 3039 2265
rect 3043 2261 3044 2265
rect 3038 2260 3044 2261
rect 3022 2247 3028 2248
rect 3022 2243 3023 2247
rect 3027 2243 3028 2247
rect 3040 2243 3042 2260
rect 3111 2255 3117 2256
rect 3111 2251 3112 2255
rect 3116 2254 3117 2255
rect 3120 2254 3122 2378
rect 3686 2375 3687 2379
rect 3691 2375 3692 2379
rect 3958 2379 3959 2383
rect 3963 2379 3964 2383
rect 3958 2378 3964 2379
rect 3686 2374 3692 2375
rect 3246 2350 3252 2351
rect 3246 2346 3247 2350
rect 3251 2346 3252 2350
rect 3246 2345 3252 2346
rect 3454 2350 3460 2351
rect 3454 2346 3455 2350
rect 3459 2346 3460 2350
rect 3454 2345 3460 2346
rect 3678 2350 3684 2351
rect 3678 2346 3679 2350
rect 3683 2346 3684 2350
rect 3678 2345 3684 2346
rect 3894 2350 3900 2351
rect 3894 2346 3895 2350
rect 3899 2346 3900 2350
rect 3894 2345 3900 2346
rect 3248 2323 3250 2345
rect 3456 2323 3458 2345
rect 3680 2323 3682 2345
rect 3896 2323 3898 2345
rect 3247 2322 3251 2323
rect 3247 2317 3251 2318
rect 3455 2322 3459 2323
rect 3455 2317 3459 2318
rect 3463 2322 3467 2323
rect 3463 2317 3467 2318
rect 3679 2322 3683 2323
rect 3679 2317 3683 2318
rect 3687 2322 3691 2323
rect 3687 2317 3691 2318
rect 3895 2322 3899 2323
rect 3895 2317 3899 2318
rect 3248 2307 3250 2317
rect 3464 2307 3466 2317
rect 3688 2307 3690 2317
rect 3896 2307 3898 2317
rect 3246 2306 3252 2307
rect 3246 2302 3247 2306
rect 3251 2302 3252 2306
rect 3246 2301 3252 2302
rect 3462 2306 3468 2307
rect 3462 2302 3463 2306
rect 3467 2302 3468 2306
rect 3462 2301 3468 2302
rect 3686 2306 3692 2307
rect 3686 2302 3687 2306
rect 3691 2302 3692 2306
rect 3686 2301 3692 2302
rect 3894 2306 3900 2307
rect 3894 2302 3895 2306
rect 3899 2302 3900 2306
rect 3894 2301 3900 2302
rect 3246 2265 3252 2266
rect 3246 2261 3247 2265
rect 3251 2261 3252 2265
rect 3246 2260 3252 2261
rect 3462 2265 3468 2266
rect 3462 2261 3463 2265
rect 3467 2261 3468 2265
rect 3462 2260 3468 2261
rect 3686 2265 3692 2266
rect 3686 2261 3687 2265
rect 3691 2261 3692 2265
rect 3686 2260 3692 2261
rect 3894 2265 3900 2266
rect 3894 2261 3895 2265
rect 3899 2261 3900 2265
rect 3894 2260 3900 2261
rect 3116 2252 3122 2254
rect 3154 2255 3160 2256
rect 3116 2251 3117 2252
rect 3111 2250 3117 2251
rect 3154 2251 3155 2255
rect 3159 2251 3160 2255
rect 3154 2250 3160 2251
rect 2479 2242 2483 2243
rect 2479 2237 2483 2238
rect 2511 2242 2515 2243
rect 2511 2237 2515 2238
rect 2671 2242 2675 2243
rect 2671 2237 2675 2238
rect 2679 2242 2683 2243
rect 2679 2237 2683 2238
rect 2847 2242 2851 2243
rect 2847 2237 2851 2238
rect 2879 2242 2883 2243
rect 3022 2242 3028 2243
rect 3039 2242 3043 2243
rect 2879 2237 2883 2238
rect 3039 2237 3043 2238
rect 3079 2242 3083 2243
rect 3079 2237 3083 2238
rect 2434 2235 2440 2236
rect 2434 2231 2435 2235
rect 2439 2231 2440 2235
rect 2434 2230 2440 2231
rect 2480 2228 2482 2237
rect 2680 2228 2682 2237
rect 2686 2235 2692 2236
rect 2686 2231 2687 2235
rect 2691 2231 2692 2235
rect 2686 2230 2692 2231
rect 2110 2227 2116 2228
rect 2110 2223 2111 2227
rect 2115 2223 2116 2227
rect 2110 2222 2116 2223
rect 2278 2227 2284 2228
rect 2278 2223 2279 2227
rect 2283 2223 2284 2227
rect 2278 2222 2284 2223
rect 2478 2227 2484 2228
rect 2478 2223 2479 2227
rect 2483 2223 2484 2227
rect 2478 2222 2484 2223
rect 2678 2227 2684 2228
rect 2678 2223 2679 2227
rect 2683 2223 2684 2227
rect 2678 2222 2684 2223
rect 2390 2219 2396 2220
rect 2390 2215 2391 2219
rect 2395 2215 2396 2219
rect 2390 2214 2396 2215
rect 2070 2208 2076 2209
rect 2030 2207 2036 2208
rect 2030 2203 2031 2207
rect 2035 2203 2036 2207
rect 2070 2204 2071 2208
rect 2075 2204 2076 2208
rect 2070 2203 2076 2204
rect 1694 2202 1700 2203
rect 2030 2202 2036 2203
rect 1694 2198 1695 2202
rect 1699 2198 1700 2202
rect 1694 2197 1700 2198
rect 1696 2175 1698 2197
rect 2032 2175 2034 2202
rect 2070 2191 2076 2192
rect 2070 2187 2071 2191
rect 2075 2187 2076 2191
rect 2070 2186 2076 2187
rect 2110 2186 2116 2187
rect 1655 2174 1659 2175
rect 1655 2169 1659 2170
rect 1695 2174 1699 2175
rect 1695 2169 1699 2170
rect 1847 2174 1851 2175
rect 1847 2169 1851 2170
rect 2031 2174 2035 2175
rect 2031 2169 2035 2170
rect 1656 2159 1658 2169
rect 1848 2159 1850 2169
rect 1654 2158 1660 2159
rect 1654 2154 1655 2158
rect 1659 2154 1660 2158
rect 1654 2153 1660 2154
rect 1846 2158 1852 2159
rect 1846 2154 1847 2158
rect 1851 2154 1852 2158
rect 2032 2154 2034 2169
rect 2072 2163 2074 2186
rect 2110 2182 2111 2186
rect 2115 2182 2116 2186
rect 2110 2181 2116 2182
rect 2278 2186 2284 2187
rect 2278 2182 2279 2186
rect 2283 2182 2284 2186
rect 2278 2181 2284 2182
rect 2112 2163 2114 2181
rect 2280 2163 2282 2181
rect 2071 2162 2075 2163
rect 2071 2157 2075 2158
rect 2111 2162 2115 2163
rect 2111 2157 2115 2158
rect 2143 2162 2147 2163
rect 2143 2157 2147 2158
rect 2279 2162 2283 2163
rect 2279 2157 2283 2158
rect 2319 2162 2323 2163
rect 2319 2157 2323 2158
rect 1846 2153 1852 2154
rect 2030 2153 2036 2154
rect 2030 2149 2031 2153
rect 2035 2149 2036 2153
rect 2030 2148 2036 2149
rect 2072 2142 2074 2157
rect 2144 2147 2146 2157
rect 2320 2147 2322 2157
rect 2142 2146 2148 2147
rect 2142 2142 2143 2146
rect 2147 2142 2148 2146
rect 2070 2141 2076 2142
rect 2142 2141 2148 2142
rect 2318 2146 2324 2147
rect 2318 2142 2319 2146
rect 2323 2142 2324 2146
rect 2318 2141 2324 2142
rect 2070 2137 2071 2141
rect 2075 2137 2076 2141
rect 2030 2136 2036 2137
rect 2070 2136 2076 2137
rect 2030 2132 2031 2136
rect 2035 2132 2036 2136
rect 2030 2131 2036 2132
rect 1638 2127 1644 2128
rect 1638 2123 1639 2127
rect 1643 2123 1644 2127
rect 1638 2122 1644 2123
rect 1640 2108 1642 2122
rect 1654 2117 1660 2118
rect 1654 2113 1655 2117
rect 1659 2113 1660 2117
rect 1654 2112 1660 2113
rect 1846 2117 1852 2118
rect 1846 2113 1847 2117
rect 1851 2113 1852 2117
rect 1846 2112 1852 2113
rect 1534 2107 1540 2108
rect 1534 2103 1535 2107
rect 1539 2103 1540 2107
rect 1534 2102 1540 2103
rect 1638 2107 1644 2108
rect 1638 2103 1639 2107
rect 1643 2103 1644 2107
rect 1638 2102 1644 2103
rect 1656 2095 1658 2112
rect 1738 2107 1744 2108
rect 1738 2103 1739 2107
rect 1743 2103 1744 2107
rect 1738 2102 1744 2103
rect 1239 2094 1243 2095
rect 1239 2089 1243 2090
rect 1279 2094 1283 2095
rect 1279 2089 1283 2090
rect 1447 2094 1451 2095
rect 1447 2089 1451 2090
rect 1463 2094 1467 2095
rect 1463 2089 1467 2090
rect 1655 2094 1659 2095
rect 1655 2089 1659 2090
rect 1663 2094 1667 2095
rect 1663 2089 1667 2090
rect 1240 2080 1242 2089
rect 1448 2080 1450 2089
rect 1454 2087 1460 2088
rect 1454 2083 1455 2087
rect 1459 2083 1460 2087
rect 1454 2082 1460 2083
rect 1238 2079 1244 2080
rect 1238 2075 1239 2079
rect 1243 2075 1244 2079
rect 1238 2074 1244 2075
rect 1446 2079 1452 2080
rect 1446 2075 1447 2079
rect 1451 2075 1452 2079
rect 1446 2074 1452 2075
rect 1114 2071 1120 2072
rect 1114 2067 1115 2071
rect 1119 2067 1120 2071
rect 1114 2066 1120 2067
rect 1038 2038 1044 2039
rect 1038 2034 1039 2038
rect 1043 2034 1044 2038
rect 1038 2033 1044 2034
rect 1238 2038 1244 2039
rect 1238 2034 1239 2038
rect 1243 2034 1244 2038
rect 1238 2033 1244 2034
rect 1446 2038 1452 2039
rect 1446 2034 1447 2038
rect 1451 2034 1452 2038
rect 1446 2033 1452 2034
rect 1040 2015 1042 2033
rect 1240 2015 1242 2033
rect 1448 2015 1450 2033
rect 1039 2014 1043 2015
rect 1039 2009 1043 2010
rect 1103 2014 1107 2015
rect 1103 2009 1107 2010
rect 1239 2014 1243 2015
rect 1239 2009 1243 2010
rect 1311 2014 1315 2015
rect 1311 2009 1315 2010
rect 1447 2014 1451 2015
rect 1447 2009 1451 2010
rect 1104 1999 1106 2009
rect 1312 1999 1314 2009
rect 1102 1998 1108 1999
rect 1102 1994 1103 1998
rect 1107 1994 1108 1998
rect 1102 1993 1108 1994
rect 1310 1998 1316 1999
rect 1310 1994 1311 1998
rect 1315 1994 1316 1998
rect 1310 1993 1316 1994
rect 1456 1968 1458 2082
rect 1664 2080 1666 2089
rect 1740 2088 1742 2102
rect 1848 2095 1850 2112
rect 2032 2095 2034 2131
rect 2070 2124 2076 2125
rect 2070 2120 2071 2124
rect 2075 2120 2076 2124
rect 2070 2119 2076 2120
rect 1847 2094 1851 2095
rect 1847 2089 1851 2090
rect 1879 2094 1883 2095
rect 1879 2089 1883 2090
rect 2031 2094 2035 2095
rect 2031 2089 2035 2090
rect 1738 2087 1744 2088
rect 1738 2083 1739 2087
rect 1743 2083 1744 2087
rect 1738 2082 1744 2083
rect 1880 2080 1882 2089
rect 1662 2079 1668 2080
rect 1662 2075 1663 2079
rect 1667 2075 1668 2079
rect 1662 2074 1668 2075
rect 1878 2079 1884 2080
rect 1878 2075 1879 2079
rect 1883 2075 1884 2079
rect 1878 2074 1884 2075
rect 2006 2071 2012 2072
rect 2006 2067 2007 2071
rect 2011 2067 2012 2071
rect 2006 2066 2012 2067
rect 1662 2038 1668 2039
rect 1662 2034 1663 2038
rect 1667 2034 1668 2038
rect 1662 2033 1668 2034
rect 1878 2038 1884 2039
rect 1878 2034 1879 2038
rect 1883 2034 1884 2038
rect 1878 2033 1884 2034
rect 1664 2015 1666 2033
rect 1880 2015 1882 2033
rect 1527 2014 1531 2015
rect 1527 2009 1531 2010
rect 1663 2014 1667 2015
rect 1663 2009 1667 2010
rect 1743 2014 1747 2015
rect 1743 2009 1747 2010
rect 1879 2014 1883 2015
rect 1879 2009 1883 2010
rect 1935 2014 1939 2015
rect 1935 2009 1939 2010
rect 1528 1999 1530 2009
rect 1744 1999 1746 2009
rect 1936 1999 1938 2009
rect 1526 1998 1532 1999
rect 1526 1994 1527 1998
rect 1531 1994 1532 1998
rect 1526 1993 1532 1994
rect 1742 1998 1748 1999
rect 1742 1994 1743 1998
rect 1747 1994 1748 1998
rect 1742 1993 1748 1994
rect 1934 1998 1940 1999
rect 1934 1994 1935 1998
rect 1939 1994 1940 1998
rect 1934 1993 1940 1994
rect 438 1967 444 1968
rect 438 1963 439 1967
rect 443 1963 444 1967
rect 438 1962 444 1963
rect 478 1967 484 1968
rect 478 1963 479 1967
rect 483 1963 484 1967
rect 478 1962 484 1963
rect 878 1967 884 1968
rect 878 1963 879 1967
rect 883 1963 884 1967
rect 878 1962 884 1963
rect 918 1967 924 1968
rect 918 1963 919 1967
rect 923 1963 924 1967
rect 918 1962 924 1963
rect 1294 1967 1300 1968
rect 1294 1963 1295 1967
rect 1299 1963 1300 1967
rect 1294 1962 1300 1963
rect 1454 1967 1460 1968
rect 1454 1963 1455 1967
rect 1459 1963 1460 1967
rect 1454 1962 1460 1963
rect 1670 1967 1676 1968
rect 1670 1963 1671 1967
rect 1675 1963 1676 1967
rect 1670 1962 1676 1963
rect 302 1957 308 1958
rect 302 1953 303 1957
rect 307 1953 308 1957
rect 302 1952 308 1953
rect 222 1947 228 1948
rect 222 1943 223 1947
rect 227 1943 228 1947
rect 222 1942 228 1943
rect 304 1931 306 1952
rect 440 1948 442 1962
rect 438 1947 444 1948
rect 438 1943 439 1947
rect 443 1943 444 1947
rect 438 1942 444 1943
rect 111 1930 115 1931
rect 111 1925 115 1926
rect 151 1930 155 1931
rect 151 1925 155 1926
rect 271 1930 275 1931
rect 271 1925 275 1926
rect 303 1930 307 1931
rect 303 1925 307 1926
rect 407 1930 411 1931
rect 407 1925 411 1926
rect 112 1897 114 1925
rect 152 1916 154 1925
rect 272 1916 274 1925
rect 408 1916 410 1925
rect 480 1924 482 1962
rect 486 1957 492 1958
rect 486 1953 487 1957
rect 491 1953 492 1957
rect 486 1952 492 1953
rect 686 1957 692 1958
rect 686 1953 687 1957
rect 691 1953 692 1957
rect 686 1952 692 1953
rect 488 1931 490 1952
rect 688 1931 690 1952
rect 880 1948 882 1962
rect 894 1957 900 1958
rect 894 1953 895 1957
rect 899 1953 900 1957
rect 894 1952 900 1953
rect 1102 1957 1108 1958
rect 1102 1953 1103 1957
rect 1107 1953 1108 1957
rect 1102 1952 1108 1953
rect 742 1947 748 1948
rect 742 1943 743 1947
rect 747 1943 748 1947
rect 742 1942 748 1943
rect 878 1947 884 1948
rect 878 1943 879 1947
rect 883 1943 884 1947
rect 878 1942 884 1943
rect 487 1930 491 1931
rect 487 1925 491 1926
rect 543 1930 547 1931
rect 543 1925 547 1926
rect 679 1930 683 1931
rect 679 1925 683 1926
rect 687 1930 691 1931
rect 687 1925 691 1926
rect 478 1923 484 1924
rect 478 1919 479 1923
rect 483 1919 484 1923
rect 478 1918 484 1919
rect 544 1916 546 1925
rect 614 1923 620 1924
rect 614 1919 615 1923
rect 619 1919 620 1923
rect 614 1918 620 1919
rect 150 1915 156 1916
rect 150 1911 151 1915
rect 155 1911 156 1915
rect 150 1910 156 1911
rect 270 1915 276 1916
rect 270 1911 271 1915
rect 275 1911 276 1915
rect 270 1910 276 1911
rect 406 1915 412 1916
rect 406 1911 407 1915
rect 411 1911 412 1915
rect 406 1910 412 1911
rect 542 1915 548 1916
rect 542 1911 543 1915
rect 547 1911 548 1915
rect 542 1910 548 1911
rect 222 1907 228 1908
rect 222 1903 223 1907
rect 227 1903 228 1907
rect 222 1902 228 1903
rect 110 1896 116 1897
rect 110 1892 111 1896
rect 115 1892 116 1896
rect 110 1891 116 1892
rect 110 1879 116 1880
rect 110 1875 111 1879
rect 115 1875 116 1879
rect 110 1874 116 1875
rect 150 1874 156 1875
rect 112 1851 114 1874
rect 150 1870 151 1874
rect 155 1870 156 1874
rect 150 1869 156 1870
rect 152 1851 154 1869
rect 111 1850 115 1851
rect 111 1845 115 1846
rect 151 1850 155 1851
rect 151 1845 155 1846
rect 112 1830 114 1845
rect 152 1835 154 1845
rect 150 1834 156 1835
rect 150 1830 151 1834
rect 155 1830 156 1834
rect 110 1829 116 1830
rect 150 1829 156 1830
rect 110 1825 111 1829
rect 115 1825 116 1829
rect 110 1824 116 1825
rect 110 1812 116 1813
rect 110 1808 111 1812
rect 115 1808 116 1812
rect 110 1807 116 1808
rect 112 1771 114 1807
rect 150 1793 156 1794
rect 150 1789 151 1793
rect 155 1789 156 1793
rect 150 1788 156 1789
rect 152 1771 154 1788
rect 224 1784 226 1902
rect 270 1874 276 1875
rect 270 1870 271 1874
rect 275 1870 276 1874
rect 270 1869 276 1870
rect 406 1874 412 1875
rect 406 1870 407 1874
rect 411 1870 412 1874
rect 406 1869 412 1870
rect 542 1874 548 1875
rect 542 1870 543 1874
rect 547 1870 548 1874
rect 542 1869 548 1870
rect 272 1851 274 1869
rect 408 1851 410 1869
rect 544 1851 546 1869
rect 271 1850 275 1851
rect 271 1845 275 1846
rect 287 1850 291 1851
rect 287 1845 291 1846
rect 407 1850 411 1851
rect 407 1845 411 1846
rect 447 1850 451 1851
rect 447 1845 451 1846
rect 543 1850 547 1851
rect 543 1845 547 1846
rect 599 1850 603 1851
rect 599 1845 603 1846
rect 288 1835 290 1845
rect 448 1835 450 1845
rect 600 1835 602 1845
rect 286 1834 292 1835
rect 286 1830 287 1834
rect 291 1830 292 1834
rect 286 1829 292 1830
rect 446 1834 452 1835
rect 446 1830 447 1834
rect 451 1830 452 1834
rect 446 1829 452 1830
rect 598 1834 604 1835
rect 598 1830 599 1834
rect 603 1830 604 1834
rect 598 1829 604 1830
rect 616 1804 618 1918
rect 680 1916 682 1925
rect 678 1915 684 1916
rect 678 1911 679 1915
rect 683 1911 684 1915
rect 678 1910 684 1911
rect 744 1908 746 1942
rect 896 1931 898 1952
rect 966 1939 972 1940
rect 966 1935 967 1939
rect 971 1935 972 1939
rect 966 1934 972 1935
rect 823 1930 827 1931
rect 823 1925 827 1926
rect 895 1930 899 1931
rect 895 1925 899 1926
rect 824 1916 826 1925
rect 822 1915 828 1916
rect 822 1911 823 1915
rect 827 1911 828 1915
rect 822 1910 828 1911
rect 968 1908 970 1934
rect 1104 1931 1106 1952
rect 1296 1948 1298 1962
rect 1310 1957 1316 1958
rect 1310 1953 1311 1957
rect 1315 1953 1316 1957
rect 1310 1952 1316 1953
rect 1526 1957 1532 1958
rect 1526 1953 1527 1957
rect 1531 1953 1532 1957
rect 1526 1952 1532 1953
rect 1294 1947 1300 1948
rect 1294 1943 1295 1947
rect 1299 1943 1300 1947
rect 1294 1942 1300 1943
rect 1312 1931 1314 1952
rect 1528 1931 1530 1952
rect 983 1930 987 1931
rect 983 1925 987 1926
rect 1103 1930 1107 1931
rect 1103 1925 1107 1926
rect 1159 1930 1163 1931
rect 1159 1925 1163 1926
rect 1311 1930 1315 1931
rect 1311 1925 1315 1926
rect 1343 1930 1347 1931
rect 1343 1925 1347 1926
rect 1527 1930 1531 1931
rect 1527 1925 1531 1926
rect 1543 1930 1547 1931
rect 1543 1925 1547 1926
rect 984 1916 986 1925
rect 1160 1916 1162 1925
rect 1344 1916 1346 1925
rect 1544 1916 1546 1925
rect 1672 1924 1674 1962
rect 1742 1957 1748 1958
rect 1742 1953 1743 1957
rect 1747 1953 1748 1957
rect 1742 1952 1748 1953
rect 1934 1957 1940 1958
rect 1934 1953 1935 1957
rect 1939 1953 1940 1957
rect 1934 1952 1940 1953
rect 1744 1931 1746 1952
rect 1936 1931 1938 1952
rect 2008 1948 2010 2066
rect 2032 2061 2034 2089
rect 2072 2079 2074 2119
rect 2214 2115 2220 2116
rect 2214 2111 2215 2115
rect 2219 2111 2220 2115
rect 2214 2110 2220 2111
rect 2142 2105 2148 2106
rect 2142 2101 2143 2105
rect 2147 2101 2148 2105
rect 2142 2100 2148 2101
rect 2144 2079 2146 2100
rect 2071 2078 2075 2079
rect 2071 2073 2075 2074
rect 2143 2078 2147 2079
rect 2143 2073 2147 2074
rect 2207 2078 2211 2079
rect 2207 2073 2211 2074
rect 2030 2060 2036 2061
rect 2030 2056 2031 2060
rect 2035 2056 2036 2060
rect 2030 2055 2036 2056
rect 2072 2045 2074 2073
rect 2208 2064 2210 2073
rect 2216 2072 2218 2110
rect 2318 2105 2324 2106
rect 2318 2101 2319 2105
rect 2323 2101 2324 2105
rect 2318 2100 2324 2101
rect 2320 2079 2322 2100
rect 2392 2096 2394 2214
rect 2478 2186 2484 2187
rect 2478 2182 2479 2186
rect 2483 2182 2484 2186
rect 2478 2181 2484 2182
rect 2678 2186 2684 2187
rect 2678 2182 2679 2186
rect 2683 2182 2684 2186
rect 2678 2181 2684 2182
rect 2480 2163 2482 2181
rect 2680 2163 2682 2181
rect 2479 2162 2483 2163
rect 2479 2157 2483 2158
rect 2495 2162 2499 2163
rect 2495 2157 2499 2158
rect 2679 2162 2683 2163
rect 2679 2157 2683 2158
rect 2496 2147 2498 2157
rect 2680 2147 2682 2157
rect 2494 2146 2500 2147
rect 2494 2142 2495 2146
rect 2499 2142 2500 2146
rect 2494 2141 2500 2142
rect 2678 2146 2684 2147
rect 2678 2142 2679 2146
rect 2683 2142 2684 2146
rect 2678 2141 2684 2142
rect 2688 2124 2690 2230
rect 2880 2228 2882 2237
rect 3063 2228 3067 2229
rect 3080 2228 3082 2237
rect 3156 2236 3158 2250
rect 3248 2243 3250 2260
rect 3464 2243 3466 2260
rect 3688 2243 3690 2260
rect 3770 2255 3776 2256
rect 3770 2251 3771 2255
rect 3775 2251 3776 2255
rect 3770 2250 3776 2251
rect 3247 2242 3251 2243
rect 3247 2237 3251 2238
rect 3279 2242 3283 2243
rect 3279 2237 3283 2238
rect 3463 2242 3467 2243
rect 3463 2237 3467 2238
rect 3487 2242 3491 2243
rect 3487 2237 3491 2238
rect 3687 2242 3691 2243
rect 3687 2237 3691 2238
rect 3703 2242 3707 2243
rect 3703 2237 3707 2238
rect 3154 2235 3160 2236
rect 3154 2231 3155 2235
rect 3159 2231 3160 2235
rect 3154 2230 3160 2231
rect 3258 2231 3264 2232
rect 2878 2227 2884 2228
rect 2878 2223 2879 2227
rect 2883 2223 2884 2227
rect 3063 2223 3067 2224
rect 3078 2227 3084 2228
rect 3078 2223 3079 2227
rect 3083 2223 3084 2227
rect 3258 2226 3259 2231
rect 3263 2226 3264 2231
rect 3280 2228 3282 2237
rect 3488 2228 3490 2237
rect 3704 2228 3706 2237
rect 3718 2235 3724 2236
rect 3718 2231 3719 2235
rect 3723 2231 3724 2235
rect 3718 2230 3724 2231
rect 3278 2227 3284 2228
rect 3259 2223 3263 2224
rect 3278 2223 3279 2227
rect 3283 2223 3284 2227
rect 2878 2222 2884 2223
rect 3064 2220 3066 2223
rect 3078 2222 3084 2223
rect 3278 2222 3284 2223
rect 3486 2227 3492 2228
rect 3486 2223 3487 2227
rect 3491 2223 3492 2227
rect 3486 2222 3492 2223
rect 3702 2227 3708 2228
rect 3702 2223 3703 2227
rect 3707 2223 3708 2227
rect 3702 2222 3708 2223
rect 3062 2219 3068 2220
rect 3062 2215 3063 2219
rect 3067 2215 3068 2219
rect 3062 2214 3068 2215
rect 3478 2215 3484 2216
rect 3478 2211 3479 2215
rect 3483 2211 3484 2215
rect 3478 2210 3484 2211
rect 2878 2186 2884 2187
rect 2878 2182 2879 2186
rect 2883 2182 2884 2186
rect 2878 2181 2884 2182
rect 3078 2186 3084 2187
rect 3078 2182 3079 2186
rect 3083 2182 3084 2186
rect 3078 2181 3084 2182
rect 3278 2186 3284 2187
rect 3278 2182 3279 2186
rect 3283 2182 3284 2186
rect 3278 2181 3284 2182
rect 2880 2163 2882 2181
rect 3080 2163 3082 2181
rect 3280 2163 3282 2181
rect 2863 2162 2867 2163
rect 2863 2157 2867 2158
rect 2879 2162 2883 2163
rect 2879 2157 2883 2158
rect 3039 2162 3043 2163
rect 3039 2157 3043 2158
rect 3079 2162 3083 2163
rect 3079 2157 3083 2158
rect 3215 2162 3219 2163
rect 3215 2157 3219 2158
rect 3279 2162 3283 2163
rect 3279 2157 3283 2158
rect 3391 2162 3395 2163
rect 3391 2157 3395 2158
rect 2864 2147 2866 2157
rect 3040 2147 3042 2157
rect 3216 2147 3218 2157
rect 3392 2147 3394 2157
rect 2862 2146 2868 2147
rect 2862 2142 2863 2146
rect 2867 2142 2868 2146
rect 2862 2141 2868 2142
rect 3038 2146 3044 2147
rect 3038 2142 3039 2146
rect 3043 2142 3044 2146
rect 3038 2141 3044 2142
rect 3214 2146 3220 2147
rect 3214 2142 3215 2146
rect 3219 2142 3220 2146
rect 3214 2141 3220 2142
rect 3390 2146 3396 2147
rect 3390 2142 3391 2146
rect 3395 2142 3396 2146
rect 3390 2141 3396 2142
rect 2686 2123 2692 2124
rect 2686 2119 2687 2123
rect 2691 2119 2692 2123
rect 2686 2118 2692 2119
rect 3110 2115 3116 2116
rect 3110 2111 3111 2115
rect 3115 2111 3116 2115
rect 3110 2110 3116 2111
rect 2494 2105 2500 2106
rect 2494 2101 2495 2105
rect 2499 2101 2500 2105
rect 2494 2100 2500 2101
rect 2678 2105 2684 2106
rect 2678 2101 2679 2105
rect 2683 2101 2684 2105
rect 2678 2100 2684 2101
rect 2862 2105 2868 2106
rect 2862 2101 2863 2105
rect 2867 2101 2868 2105
rect 2862 2100 2868 2101
rect 3038 2105 3044 2106
rect 3038 2101 3039 2105
rect 3043 2101 3044 2105
rect 3038 2100 3044 2101
rect 2390 2095 2396 2096
rect 2390 2091 2391 2095
rect 2395 2091 2396 2095
rect 2390 2090 2396 2091
rect 2496 2079 2498 2100
rect 2680 2079 2682 2100
rect 2864 2079 2866 2100
rect 2926 2095 2932 2096
rect 2926 2091 2927 2095
rect 2931 2091 2932 2095
rect 2926 2090 2932 2091
rect 2319 2078 2323 2079
rect 2319 2073 2323 2074
rect 2391 2078 2395 2079
rect 2391 2073 2395 2074
rect 2495 2078 2499 2079
rect 2495 2073 2499 2074
rect 2575 2078 2579 2079
rect 2575 2073 2579 2074
rect 2679 2078 2683 2079
rect 2679 2073 2683 2074
rect 2759 2078 2763 2079
rect 2759 2073 2763 2074
rect 2863 2078 2867 2079
rect 2863 2073 2867 2074
rect 2214 2071 2220 2072
rect 2214 2067 2215 2071
rect 2219 2067 2220 2071
rect 2214 2066 2220 2067
rect 2392 2064 2394 2073
rect 2576 2064 2578 2073
rect 2646 2071 2652 2072
rect 2646 2067 2647 2071
rect 2651 2067 2652 2071
rect 2646 2066 2652 2067
rect 2206 2063 2212 2064
rect 2206 2059 2207 2063
rect 2211 2059 2212 2063
rect 2206 2058 2212 2059
rect 2390 2063 2396 2064
rect 2390 2059 2391 2063
rect 2395 2059 2396 2063
rect 2390 2058 2396 2059
rect 2574 2063 2580 2064
rect 2574 2059 2575 2063
rect 2579 2059 2580 2063
rect 2574 2058 2580 2059
rect 2382 2051 2388 2052
rect 2382 2047 2383 2051
rect 2387 2047 2388 2051
rect 2382 2046 2388 2047
rect 2070 2044 2076 2045
rect 2030 2043 2036 2044
rect 2030 2039 2031 2043
rect 2035 2039 2036 2043
rect 2070 2040 2071 2044
rect 2075 2040 2076 2044
rect 2070 2039 2076 2040
rect 2030 2038 2036 2039
rect 2032 2015 2034 2038
rect 2070 2027 2076 2028
rect 2070 2023 2071 2027
rect 2075 2023 2076 2027
rect 2070 2022 2076 2023
rect 2206 2022 2212 2023
rect 2031 2014 2035 2015
rect 2031 2009 2035 2010
rect 2032 1994 2034 2009
rect 2072 1995 2074 2022
rect 2206 2018 2207 2022
rect 2211 2018 2212 2022
rect 2206 2017 2212 2018
rect 2208 1995 2210 2017
rect 2071 1994 2075 1995
rect 2030 1993 2036 1994
rect 2030 1989 2031 1993
rect 2035 1989 2036 1993
rect 2071 1989 2075 1990
rect 2207 1994 2211 1995
rect 2207 1989 2211 1990
rect 2279 1994 2283 1995
rect 2279 1989 2283 1990
rect 2030 1988 2036 1989
rect 2030 1976 2036 1977
rect 2030 1972 2031 1976
rect 2035 1972 2036 1976
rect 2072 1974 2074 1989
rect 2280 1979 2282 1989
rect 2278 1978 2284 1979
rect 2278 1974 2279 1978
rect 2283 1974 2284 1978
rect 2030 1971 2036 1972
rect 2070 1973 2076 1974
rect 2278 1973 2284 1974
rect 2006 1947 2012 1948
rect 2006 1943 2007 1947
rect 2011 1943 2012 1947
rect 2006 1942 2012 1943
rect 2032 1931 2034 1971
rect 2070 1969 2071 1973
rect 2075 1969 2076 1973
rect 2070 1968 2076 1969
rect 2070 1956 2076 1957
rect 2070 1952 2071 1956
rect 2075 1952 2076 1956
rect 2070 1951 2076 1952
rect 1743 1930 1747 1931
rect 1743 1925 1747 1926
rect 1751 1930 1755 1931
rect 1751 1925 1755 1926
rect 1935 1930 1939 1931
rect 1935 1925 1939 1926
rect 2031 1930 2035 1931
rect 2031 1925 2035 1926
rect 1550 1923 1556 1924
rect 1550 1919 1551 1923
rect 1555 1919 1556 1923
rect 1550 1918 1556 1919
rect 1670 1923 1676 1924
rect 1670 1919 1671 1923
rect 1675 1919 1676 1923
rect 1670 1918 1676 1919
rect 982 1915 988 1916
rect 982 1911 983 1915
rect 987 1911 988 1915
rect 982 1910 988 1911
rect 1158 1915 1164 1916
rect 1158 1911 1159 1915
rect 1163 1911 1164 1915
rect 1158 1910 1164 1911
rect 1342 1915 1348 1916
rect 1342 1911 1343 1915
rect 1347 1911 1348 1915
rect 1342 1910 1348 1911
rect 1542 1915 1548 1916
rect 1542 1911 1543 1915
rect 1547 1911 1548 1915
rect 1542 1910 1548 1911
rect 742 1907 748 1908
rect 742 1903 743 1907
rect 747 1903 748 1907
rect 742 1902 748 1903
rect 966 1907 972 1908
rect 966 1903 967 1907
rect 971 1903 972 1907
rect 966 1902 972 1903
rect 678 1874 684 1875
rect 678 1870 679 1874
rect 683 1870 684 1874
rect 678 1869 684 1870
rect 822 1874 828 1875
rect 822 1870 823 1874
rect 827 1870 828 1874
rect 822 1869 828 1870
rect 982 1874 988 1875
rect 982 1870 983 1874
rect 987 1870 988 1874
rect 982 1869 988 1870
rect 1158 1874 1164 1875
rect 1158 1870 1159 1874
rect 1163 1870 1164 1874
rect 1158 1869 1164 1870
rect 1342 1874 1348 1875
rect 1342 1870 1343 1874
rect 1347 1870 1348 1874
rect 1342 1869 1348 1870
rect 1542 1874 1548 1875
rect 1542 1870 1543 1874
rect 1547 1870 1548 1874
rect 1542 1869 1548 1870
rect 680 1851 682 1869
rect 824 1851 826 1869
rect 984 1851 986 1869
rect 1042 1855 1048 1856
rect 1042 1851 1043 1855
rect 1047 1851 1048 1855
rect 1160 1851 1162 1869
rect 1344 1851 1346 1869
rect 1544 1851 1546 1869
rect 1552 1856 1554 1918
rect 1752 1916 1754 1925
rect 1936 1916 1938 1925
rect 1750 1915 1756 1916
rect 1750 1911 1751 1915
rect 1755 1911 1756 1915
rect 1750 1910 1756 1911
rect 1934 1915 1940 1916
rect 1934 1911 1935 1915
rect 1939 1911 1940 1915
rect 1934 1910 1940 1911
rect 2006 1907 2012 1908
rect 2006 1903 2007 1907
rect 2011 1903 2012 1907
rect 2006 1902 2012 1903
rect 1750 1874 1756 1875
rect 1750 1870 1751 1874
rect 1755 1870 1756 1874
rect 1750 1869 1756 1870
rect 1934 1874 1940 1875
rect 1934 1870 1935 1874
rect 1939 1870 1940 1874
rect 1934 1869 1940 1870
rect 1550 1855 1556 1856
rect 1550 1851 1551 1855
rect 1555 1851 1556 1855
rect 1752 1851 1754 1869
rect 1936 1851 1938 1869
rect 679 1850 683 1851
rect 679 1845 683 1846
rect 751 1850 755 1851
rect 751 1845 755 1846
rect 823 1850 827 1851
rect 823 1845 827 1846
rect 919 1850 923 1851
rect 919 1845 923 1846
rect 983 1850 987 1851
rect 1042 1850 1048 1851
rect 1103 1850 1107 1851
rect 983 1845 987 1846
rect 752 1835 754 1845
rect 920 1835 922 1845
rect 750 1834 756 1835
rect 750 1830 751 1834
rect 755 1830 756 1834
rect 750 1829 756 1830
rect 918 1834 924 1835
rect 918 1830 919 1834
rect 923 1830 924 1834
rect 918 1829 924 1830
rect 1044 1804 1046 1850
rect 1103 1845 1107 1846
rect 1159 1850 1163 1851
rect 1159 1845 1163 1846
rect 1303 1850 1307 1851
rect 1303 1845 1307 1846
rect 1343 1850 1347 1851
rect 1343 1845 1347 1846
rect 1511 1850 1515 1851
rect 1511 1845 1515 1846
rect 1543 1850 1547 1851
rect 1550 1850 1556 1851
rect 1735 1850 1739 1851
rect 1543 1845 1547 1846
rect 1735 1845 1739 1846
rect 1751 1850 1755 1851
rect 1751 1845 1755 1846
rect 1935 1850 1939 1851
rect 1935 1845 1939 1846
rect 1104 1835 1106 1845
rect 1304 1835 1306 1845
rect 1512 1835 1514 1845
rect 1736 1835 1738 1845
rect 1936 1835 1938 1845
rect 1102 1834 1108 1835
rect 1102 1830 1103 1834
rect 1107 1830 1108 1834
rect 1102 1829 1108 1830
rect 1302 1834 1308 1835
rect 1302 1830 1303 1834
rect 1307 1830 1308 1834
rect 1302 1829 1308 1830
rect 1510 1834 1516 1835
rect 1510 1830 1511 1834
rect 1515 1830 1516 1834
rect 1510 1829 1516 1830
rect 1734 1834 1740 1835
rect 1734 1830 1735 1834
rect 1739 1830 1740 1834
rect 1734 1829 1740 1830
rect 1934 1834 1940 1835
rect 1934 1830 1935 1834
rect 1939 1830 1940 1834
rect 1934 1829 1940 1830
rect 426 1803 432 1804
rect 426 1799 427 1803
rect 431 1799 432 1803
rect 426 1798 432 1799
rect 614 1803 620 1804
rect 614 1799 615 1803
rect 619 1799 620 1803
rect 614 1798 620 1799
rect 1042 1803 1048 1804
rect 1042 1799 1043 1803
rect 1047 1799 1048 1803
rect 1042 1798 1048 1799
rect 286 1793 292 1794
rect 286 1789 287 1793
rect 291 1789 292 1793
rect 286 1788 292 1789
rect 222 1783 228 1784
rect 222 1779 223 1783
rect 227 1779 228 1783
rect 222 1778 228 1779
rect 288 1771 290 1788
rect 428 1784 430 1798
rect 446 1793 452 1794
rect 446 1789 447 1793
rect 451 1789 452 1793
rect 446 1788 452 1789
rect 598 1793 604 1794
rect 598 1789 599 1793
rect 603 1789 604 1793
rect 598 1788 604 1789
rect 750 1793 756 1794
rect 750 1789 751 1793
rect 755 1789 756 1793
rect 750 1788 756 1789
rect 918 1793 924 1794
rect 918 1789 919 1793
rect 923 1789 924 1793
rect 918 1788 924 1789
rect 1102 1793 1108 1794
rect 1102 1789 1103 1793
rect 1107 1789 1108 1793
rect 1102 1788 1108 1789
rect 1302 1793 1308 1794
rect 1302 1789 1303 1793
rect 1307 1789 1308 1793
rect 1302 1788 1308 1789
rect 1510 1793 1516 1794
rect 1510 1789 1511 1793
rect 1515 1789 1516 1793
rect 1510 1788 1516 1789
rect 1734 1793 1740 1794
rect 1734 1789 1735 1793
rect 1739 1789 1740 1793
rect 1734 1788 1740 1789
rect 1934 1793 1940 1794
rect 1934 1789 1935 1793
rect 1939 1789 1940 1793
rect 1934 1788 1940 1789
rect 426 1783 432 1784
rect 426 1779 427 1783
rect 431 1779 432 1783
rect 426 1778 432 1779
rect 448 1771 450 1788
rect 600 1771 602 1788
rect 752 1771 754 1788
rect 814 1783 820 1784
rect 814 1779 815 1783
rect 819 1779 820 1783
rect 814 1778 820 1779
rect 111 1770 115 1771
rect 111 1765 115 1766
rect 151 1770 155 1771
rect 151 1765 155 1766
rect 207 1770 211 1771
rect 207 1765 211 1766
rect 287 1770 291 1771
rect 287 1765 291 1766
rect 383 1770 387 1771
rect 383 1765 387 1766
rect 447 1770 451 1771
rect 447 1765 451 1766
rect 567 1770 571 1771
rect 567 1765 571 1766
rect 599 1770 603 1771
rect 599 1765 603 1766
rect 751 1770 755 1771
rect 751 1765 755 1766
rect 112 1737 114 1765
rect 208 1756 210 1765
rect 384 1756 386 1765
rect 568 1756 570 1765
rect 752 1756 754 1765
rect 206 1755 212 1756
rect 206 1751 207 1755
rect 211 1751 212 1755
rect 206 1750 212 1751
rect 382 1755 388 1756
rect 382 1751 383 1755
rect 387 1751 388 1755
rect 382 1750 388 1751
rect 566 1755 572 1756
rect 566 1751 567 1755
rect 571 1751 572 1755
rect 566 1750 572 1751
rect 750 1755 756 1756
rect 750 1751 751 1755
rect 755 1751 756 1755
rect 750 1750 756 1751
rect 816 1748 818 1778
rect 920 1771 922 1788
rect 1104 1771 1106 1788
rect 1304 1771 1306 1788
rect 1512 1771 1514 1788
rect 1736 1771 1738 1788
rect 1742 1783 1748 1784
rect 1742 1779 1743 1783
rect 1747 1779 1748 1783
rect 1742 1778 1748 1779
rect 919 1770 923 1771
rect 919 1765 923 1766
rect 935 1770 939 1771
rect 935 1765 939 1766
rect 1103 1770 1107 1771
rect 1103 1765 1107 1766
rect 1111 1770 1115 1771
rect 1111 1765 1115 1766
rect 1279 1770 1283 1771
rect 1279 1765 1283 1766
rect 1303 1770 1307 1771
rect 1303 1765 1307 1766
rect 1455 1770 1459 1771
rect 1455 1765 1459 1766
rect 1511 1770 1515 1771
rect 1511 1765 1515 1766
rect 1631 1770 1635 1771
rect 1631 1765 1635 1766
rect 1735 1770 1739 1771
rect 1735 1765 1739 1766
rect 936 1756 938 1765
rect 1006 1763 1012 1764
rect 1006 1759 1007 1763
rect 1011 1759 1012 1763
rect 1006 1758 1012 1759
rect 934 1755 940 1756
rect 934 1751 935 1755
rect 939 1751 940 1755
rect 934 1750 940 1751
rect 366 1747 372 1748
rect 366 1743 367 1747
rect 371 1743 372 1747
rect 366 1742 372 1743
rect 814 1747 820 1748
rect 814 1743 815 1747
rect 819 1743 820 1747
rect 814 1742 820 1743
rect 110 1736 116 1737
rect 110 1732 111 1736
rect 115 1732 116 1736
rect 110 1731 116 1732
rect 110 1719 116 1720
rect 110 1715 111 1719
rect 115 1715 116 1719
rect 110 1714 116 1715
rect 206 1714 212 1715
rect 112 1699 114 1714
rect 206 1710 207 1714
rect 211 1710 212 1714
rect 206 1709 212 1710
rect 208 1699 210 1709
rect 111 1698 115 1699
rect 111 1693 115 1694
rect 207 1698 211 1699
rect 207 1693 211 1694
rect 303 1698 307 1699
rect 303 1693 307 1694
rect 112 1678 114 1693
rect 304 1683 306 1693
rect 302 1682 308 1683
rect 302 1678 303 1682
rect 307 1678 308 1682
rect 110 1677 116 1678
rect 302 1677 308 1678
rect 110 1673 111 1677
rect 115 1673 116 1677
rect 110 1672 116 1673
rect 110 1660 116 1661
rect 110 1656 111 1660
rect 115 1656 116 1660
rect 110 1655 116 1656
rect 112 1623 114 1655
rect 302 1641 308 1642
rect 302 1637 303 1641
rect 307 1637 308 1641
rect 302 1636 308 1637
rect 304 1623 306 1636
rect 368 1632 370 1742
rect 382 1714 388 1715
rect 382 1710 383 1714
rect 387 1710 388 1714
rect 382 1709 388 1710
rect 566 1714 572 1715
rect 566 1710 567 1714
rect 571 1710 572 1714
rect 566 1709 572 1710
rect 750 1714 756 1715
rect 750 1710 751 1714
rect 755 1710 756 1714
rect 750 1709 756 1710
rect 934 1714 940 1715
rect 934 1710 935 1714
rect 939 1710 940 1714
rect 934 1709 940 1710
rect 384 1699 386 1709
rect 568 1699 570 1709
rect 752 1699 754 1709
rect 936 1699 938 1709
rect 383 1698 387 1699
rect 383 1693 387 1694
rect 535 1698 539 1699
rect 535 1693 539 1694
rect 567 1698 571 1699
rect 567 1693 571 1694
rect 751 1698 755 1699
rect 751 1693 755 1694
rect 767 1698 771 1699
rect 767 1693 771 1694
rect 935 1698 939 1699
rect 935 1693 939 1694
rect 983 1698 987 1699
rect 983 1693 987 1694
rect 536 1683 538 1693
rect 768 1683 770 1693
rect 984 1683 986 1693
rect 534 1682 540 1683
rect 534 1678 535 1682
rect 539 1678 540 1682
rect 534 1677 540 1678
rect 766 1682 772 1683
rect 766 1678 767 1682
rect 771 1678 772 1682
rect 766 1677 772 1678
rect 982 1682 988 1683
rect 982 1678 983 1682
rect 987 1678 988 1682
rect 982 1677 988 1678
rect 1008 1652 1010 1758
rect 1112 1756 1114 1765
rect 1280 1756 1282 1765
rect 1456 1756 1458 1765
rect 1632 1756 1634 1765
rect 1702 1763 1708 1764
rect 1702 1759 1703 1763
rect 1707 1759 1708 1763
rect 1702 1758 1708 1759
rect 1110 1755 1116 1756
rect 1110 1751 1111 1755
rect 1115 1751 1116 1755
rect 1110 1750 1116 1751
rect 1278 1755 1284 1756
rect 1278 1751 1279 1755
rect 1283 1751 1284 1755
rect 1278 1750 1284 1751
rect 1454 1755 1460 1756
rect 1454 1751 1455 1755
rect 1459 1751 1460 1755
rect 1454 1750 1460 1751
rect 1630 1755 1636 1756
rect 1630 1751 1631 1755
rect 1635 1751 1636 1755
rect 1630 1750 1636 1751
rect 1263 1748 1267 1749
rect 1262 1743 1263 1748
rect 1267 1743 1268 1748
rect 1262 1742 1268 1743
rect 1110 1714 1116 1715
rect 1110 1710 1111 1714
rect 1115 1710 1116 1714
rect 1110 1709 1116 1710
rect 1278 1714 1284 1715
rect 1278 1710 1279 1714
rect 1283 1710 1284 1714
rect 1278 1709 1284 1710
rect 1454 1714 1460 1715
rect 1454 1710 1455 1714
rect 1459 1710 1460 1714
rect 1454 1709 1460 1710
rect 1630 1714 1636 1715
rect 1630 1710 1631 1714
rect 1635 1710 1636 1714
rect 1630 1709 1636 1710
rect 1112 1699 1114 1709
rect 1280 1699 1282 1709
rect 1456 1699 1458 1709
rect 1632 1699 1634 1709
rect 1111 1698 1115 1699
rect 1111 1693 1115 1694
rect 1191 1698 1195 1699
rect 1191 1693 1195 1694
rect 1279 1698 1283 1699
rect 1279 1693 1283 1694
rect 1383 1698 1387 1699
rect 1383 1693 1387 1694
rect 1455 1698 1459 1699
rect 1455 1693 1459 1694
rect 1567 1698 1571 1699
rect 1567 1693 1571 1694
rect 1631 1698 1635 1699
rect 1631 1693 1635 1694
rect 1192 1683 1194 1693
rect 1384 1683 1386 1693
rect 1568 1683 1570 1693
rect 1190 1682 1196 1683
rect 1190 1678 1191 1682
rect 1195 1678 1196 1682
rect 1190 1677 1196 1678
rect 1382 1682 1388 1683
rect 1382 1678 1383 1682
rect 1387 1678 1388 1682
rect 1382 1677 1388 1678
rect 1566 1682 1572 1683
rect 1566 1678 1567 1682
rect 1571 1678 1572 1682
rect 1566 1677 1572 1678
rect 1704 1672 1706 1758
rect 1744 1749 1746 1778
rect 1936 1771 1938 1788
rect 2008 1784 2010 1902
rect 2032 1897 2034 1925
rect 2072 1915 2074 1951
rect 2278 1937 2284 1938
rect 2278 1933 2279 1937
rect 2283 1933 2284 1937
rect 2278 1932 2284 1933
rect 2280 1915 2282 1932
rect 2384 1928 2386 2046
rect 2390 2022 2396 2023
rect 2390 2018 2391 2022
rect 2395 2018 2396 2022
rect 2390 2017 2396 2018
rect 2574 2022 2580 2023
rect 2574 2018 2575 2022
rect 2579 2018 2580 2022
rect 2574 2017 2580 2018
rect 2392 1995 2394 2017
rect 2576 1995 2578 2017
rect 2391 1994 2395 1995
rect 2391 1989 2395 1990
rect 2463 1994 2467 1995
rect 2463 1989 2467 1990
rect 2575 1994 2579 1995
rect 2575 1989 2579 1990
rect 2639 1994 2643 1995
rect 2639 1989 2643 1990
rect 2464 1979 2466 1989
rect 2640 1979 2642 1989
rect 2462 1978 2468 1979
rect 2462 1974 2463 1978
rect 2467 1974 2468 1978
rect 2462 1973 2468 1974
rect 2638 1978 2644 1979
rect 2638 1974 2639 1978
rect 2643 1974 2644 1978
rect 2638 1973 2644 1974
rect 2648 1948 2650 2066
rect 2760 2064 2762 2073
rect 2758 2063 2764 2064
rect 2758 2059 2759 2063
rect 2763 2059 2764 2063
rect 2758 2058 2764 2059
rect 2928 2056 2930 2090
rect 3040 2079 3042 2100
rect 2935 2078 2939 2079
rect 2935 2073 2939 2074
rect 3039 2078 3043 2079
rect 3039 2073 3043 2074
rect 3103 2078 3107 2079
rect 3103 2073 3107 2074
rect 2936 2064 2938 2073
rect 3104 2064 3106 2073
rect 3112 2072 3114 2110
rect 3214 2105 3220 2106
rect 3214 2101 3215 2105
rect 3219 2101 3220 2105
rect 3214 2100 3220 2101
rect 3390 2105 3396 2106
rect 3390 2101 3391 2105
rect 3395 2101 3396 2105
rect 3390 2100 3396 2101
rect 3216 2079 3218 2100
rect 3246 2079 3252 2080
rect 3392 2079 3394 2100
rect 3480 2096 3482 2210
rect 3486 2186 3492 2187
rect 3486 2182 3487 2186
rect 3491 2182 3492 2186
rect 3486 2181 3492 2182
rect 3702 2186 3708 2187
rect 3702 2182 3703 2186
rect 3707 2182 3708 2186
rect 3702 2181 3708 2182
rect 3488 2163 3490 2181
rect 3704 2163 3706 2181
rect 3487 2162 3491 2163
rect 3487 2157 3491 2158
rect 3567 2162 3571 2163
rect 3567 2157 3571 2158
rect 3703 2162 3707 2163
rect 3703 2157 3707 2158
rect 3568 2147 3570 2157
rect 3566 2146 3572 2147
rect 3566 2142 3567 2146
rect 3571 2142 3572 2146
rect 3566 2141 3572 2142
rect 3720 2116 3722 2230
rect 3772 2220 3774 2250
rect 3896 2243 3898 2260
rect 3960 2256 3962 2378
rect 3992 2373 3994 2401
rect 3990 2372 3996 2373
rect 3990 2368 3991 2372
rect 3995 2368 3996 2372
rect 3990 2367 3996 2368
rect 3990 2355 3996 2356
rect 3990 2351 3991 2355
rect 3995 2351 3996 2355
rect 3990 2350 3996 2351
rect 3992 2323 3994 2350
rect 3991 2322 3995 2323
rect 3991 2317 3995 2318
rect 3992 2302 3994 2317
rect 3990 2301 3996 2302
rect 3990 2297 3991 2301
rect 3995 2297 3996 2301
rect 3990 2296 3996 2297
rect 3990 2284 3996 2285
rect 3990 2280 3991 2284
rect 3995 2280 3996 2284
rect 3990 2279 3996 2280
rect 3966 2275 3972 2276
rect 3966 2271 3967 2275
rect 3971 2271 3972 2275
rect 3966 2270 3972 2271
rect 3958 2255 3964 2256
rect 3958 2251 3959 2255
rect 3963 2251 3964 2255
rect 3958 2250 3964 2251
rect 3895 2242 3899 2243
rect 3895 2237 3899 2238
rect 3896 2228 3898 2237
rect 3968 2236 3970 2270
rect 3992 2243 3994 2279
rect 3991 2242 3995 2243
rect 3991 2237 3995 2238
rect 3966 2235 3972 2236
rect 3966 2231 3967 2235
rect 3971 2231 3972 2235
rect 3966 2230 3972 2231
rect 3894 2227 3900 2228
rect 3894 2223 3895 2227
rect 3899 2223 3900 2227
rect 3894 2222 3900 2223
rect 3770 2219 3776 2220
rect 3770 2215 3771 2219
rect 3775 2215 3776 2219
rect 3770 2214 3776 2215
rect 3958 2219 3964 2220
rect 3958 2215 3959 2219
rect 3963 2215 3964 2219
rect 3958 2214 3964 2215
rect 3894 2186 3900 2187
rect 3894 2182 3895 2186
rect 3899 2182 3900 2186
rect 3894 2181 3900 2182
rect 3896 2163 3898 2181
rect 3743 2162 3747 2163
rect 3743 2157 3747 2158
rect 3895 2162 3899 2163
rect 3895 2157 3899 2158
rect 3744 2147 3746 2157
rect 3896 2147 3898 2157
rect 3742 2146 3748 2147
rect 3742 2142 3743 2146
rect 3747 2142 3748 2146
rect 3742 2141 3748 2142
rect 3894 2146 3900 2147
rect 3894 2142 3895 2146
rect 3899 2142 3900 2146
rect 3894 2141 3900 2142
rect 3718 2115 3724 2116
rect 3718 2111 3719 2115
rect 3723 2111 3724 2115
rect 3718 2110 3724 2111
rect 3566 2105 3572 2106
rect 3566 2101 3567 2105
rect 3571 2101 3572 2105
rect 3566 2100 3572 2101
rect 3742 2105 3748 2106
rect 3742 2101 3743 2105
rect 3747 2101 3748 2105
rect 3742 2100 3748 2101
rect 3894 2105 3900 2106
rect 3894 2101 3895 2105
rect 3899 2101 3900 2105
rect 3894 2100 3900 2101
rect 3478 2095 3484 2096
rect 3478 2091 3479 2095
rect 3483 2091 3484 2095
rect 3478 2090 3484 2091
rect 3568 2079 3570 2100
rect 3744 2079 3746 2100
rect 3814 2095 3820 2096
rect 3814 2091 3815 2095
rect 3819 2091 3820 2095
rect 3814 2090 3820 2091
rect 3215 2078 3219 2079
rect 3246 2075 3247 2079
rect 3251 2075 3252 2079
rect 3246 2074 3252 2075
rect 3263 2078 3267 2079
rect 3215 2073 3219 2074
rect 3110 2071 3116 2072
rect 3110 2067 3111 2071
rect 3115 2067 3116 2071
rect 3110 2066 3116 2067
rect 2934 2063 2940 2064
rect 2934 2059 2935 2063
rect 2939 2059 2940 2063
rect 2934 2058 2940 2059
rect 3102 2063 3108 2064
rect 3102 2059 3103 2063
rect 3107 2059 3108 2063
rect 3102 2058 3108 2059
rect 3248 2056 3250 2074
rect 3263 2073 3267 2074
rect 3391 2078 3395 2079
rect 3391 2073 3395 2074
rect 3423 2078 3427 2079
rect 3423 2073 3427 2074
rect 3567 2078 3571 2079
rect 3567 2073 3571 2074
rect 3583 2078 3587 2079
rect 3583 2073 3587 2074
rect 3743 2078 3747 2079
rect 3743 2073 3747 2074
rect 3751 2078 3755 2079
rect 3751 2073 3755 2074
rect 3264 2064 3266 2073
rect 3424 2064 3426 2073
rect 3584 2064 3586 2073
rect 3638 2071 3644 2072
rect 3638 2067 3639 2071
rect 3643 2067 3644 2071
rect 3638 2066 3644 2067
rect 3262 2063 3268 2064
rect 3262 2059 3263 2063
rect 3267 2059 3268 2063
rect 3262 2058 3268 2059
rect 3422 2063 3428 2064
rect 3422 2059 3423 2063
rect 3427 2059 3428 2063
rect 3422 2058 3428 2059
rect 3582 2063 3588 2064
rect 3582 2059 3583 2063
rect 3587 2059 3588 2063
rect 3582 2058 3588 2059
rect 2926 2055 2932 2056
rect 2926 2051 2927 2055
rect 2931 2051 2932 2055
rect 2926 2050 2932 2051
rect 3246 2055 3252 2056
rect 3246 2051 3247 2055
rect 3251 2051 3252 2055
rect 3246 2050 3252 2051
rect 3254 2051 3260 2052
rect 3254 2047 3255 2051
rect 3259 2047 3260 2051
rect 3254 2046 3260 2047
rect 2758 2022 2764 2023
rect 2758 2018 2759 2022
rect 2763 2018 2764 2022
rect 2758 2017 2764 2018
rect 2934 2022 2940 2023
rect 2934 2018 2935 2022
rect 2939 2018 2940 2022
rect 2934 2017 2940 2018
rect 3102 2022 3108 2023
rect 3102 2018 3103 2022
rect 3107 2018 3108 2022
rect 3102 2017 3108 2018
rect 2760 1995 2762 2017
rect 2936 1995 2938 2017
rect 3104 1995 3106 2017
rect 2759 1994 2763 1995
rect 2759 1989 2763 1990
rect 2815 1994 2819 1995
rect 2815 1989 2819 1990
rect 2935 1994 2939 1995
rect 2935 1989 2939 1990
rect 2983 1994 2987 1995
rect 2983 1989 2987 1990
rect 3103 1994 3107 1995
rect 3103 1989 3107 1990
rect 3151 1994 3155 1995
rect 3151 1989 3155 1990
rect 2816 1979 2818 1989
rect 2984 1979 2986 1989
rect 3152 1979 3154 1989
rect 2814 1978 2820 1979
rect 2814 1974 2815 1978
rect 2819 1974 2820 1978
rect 2814 1973 2820 1974
rect 2982 1978 2988 1979
rect 2982 1974 2983 1978
rect 2987 1974 2988 1978
rect 2982 1973 2988 1974
rect 3150 1978 3156 1979
rect 3150 1974 3151 1978
rect 3155 1974 3156 1978
rect 3150 1973 3156 1974
rect 2446 1947 2452 1948
rect 2446 1943 2447 1947
rect 2451 1943 2452 1947
rect 2446 1942 2452 1943
rect 2590 1947 2596 1948
rect 2590 1943 2591 1947
rect 2595 1943 2596 1947
rect 2590 1942 2596 1943
rect 2646 1947 2652 1948
rect 2646 1943 2647 1947
rect 2651 1943 2652 1947
rect 2646 1942 2652 1943
rect 2448 1928 2450 1942
rect 2462 1937 2468 1938
rect 2462 1933 2463 1937
rect 2467 1933 2468 1937
rect 2462 1932 2468 1933
rect 2382 1927 2388 1928
rect 2382 1923 2383 1927
rect 2387 1923 2388 1927
rect 2382 1922 2388 1923
rect 2446 1927 2452 1928
rect 2446 1923 2447 1927
rect 2451 1923 2452 1927
rect 2446 1922 2452 1923
rect 2464 1915 2466 1932
rect 2592 1916 2594 1942
rect 2638 1937 2644 1938
rect 2638 1933 2639 1937
rect 2643 1933 2644 1937
rect 2638 1932 2644 1933
rect 2814 1937 2820 1938
rect 2814 1933 2815 1937
rect 2819 1933 2820 1937
rect 2814 1932 2820 1933
rect 2982 1937 2988 1938
rect 2982 1933 2983 1937
rect 2987 1933 2988 1937
rect 2982 1932 2988 1933
rect 3150 1937 3156 1938
rect 3150 1933 3151 1937
rect 3155 1933 3156 1937
rect 3150 1932 3156 1933
rect 2590 1915 2596 1916
rect 2640 1915 2642 1932
rect 2816 1915 2818 1932
rect 2984 1915 2986 1932
rect 3152 1915 3154 1932
rect 3256 1928 3258 2046
rect 3262 2022 3268 2023
rect 3262 2018 3263 2022
rect 3267 2018 3268 2022
rect 3262 2017 3268 2018
rect 3422 2022 3428 2023
rect 3422 2018 3423 2022
rect 3427 2018 3428 2022
rect 3422 2017 3428 2018
rect 3582 2022 3588 2023
rect 3582 2018 3583 2022
rect 3587 2018 3588 2022
rect 3582 2017 3588 2018
rect 3264 1995 3266 2017
rect 3424 1995 3426 2017
rect 3584 1995 3586 2017
rect 3263 1994 3267 1995
rect 3263 1989 3267 1990
rect 3311 1994 3315 1995
rect 3311 1989 3315 1990
rect 3423 1994 3427 1995
rect 3423 1989 3427 1990
rect 3463 1994 3467 1995
rect 3463 1989 3467 1990
rect 3583 1994 3587 1995
rect 3583 1989 3587 1990
rect 3615 1994 3619 1995
rect 3615 1989 3619 1990
rect 3312 1979 3314 1989
rect 3464 1979 3466 1989
rect 3616 1979 3618 1989
rect 3310 1978 3316 1979
rect 3310 1974 3311 1978
rect 3315 1974 3316 1978
rect 3310 1973 3316 1974
rect 3462 1978 3468 1979
rect 3462 1974 3463 1978
rect 3467 1974 3468 1978
rect 3462 1973 3468 1974
rect 3614 1978 3620 1979
rect 3614 1974 3615 1978
rect 3619 1974 3620 1978
rect 3614 1973 3620 1974
rect 3640 1948 3642 2066
rect 3752 2064 3754 2073
rect 3750 2063 3756 2064
rect 3750 2059 3751 2063
rect 3755 2059 3756 2063
rect 3750 2058 3756 2059
rect 3816 2056 3818 2090
rect 3896 2079 3898 2100
rect 3960 2096 3962 2214
rect 3992 2209 3994 2237
rect 3990 2208 3996 2209
rect 3990 2204 3991 2208
rect 3995 2204 3996 2208
rect 3990 2203 3996 2204
rect 3990 2191 3996 2192
rect 3990 2187 3991 2191
rect 3995 2187 3996 2191
rect 3990 2186 3996 2187
rect 3992 2163 3994 2186
rect 3991 2162 3995 2163
rect 3991 2157 3995 2158
rect 3992 2142 3994 2157
rect 3990 2141 3996 2142
rect 3990 2137 3991 2141
rect 3995 2137 3996 2141
rect 3990 2136 3996 2137
rect 3990 2124 3996 2125
rect 3990 2120 3991 2124
rect 3995 2120 3996 2124
rect 3990 2119 3996 2120
rect 3966 2115 3972 2116
rect 3966 2111 3967 2115
rect 3971 2111 3972 2115
rect 3966 2110 3972 2111
rect 3958 2095 3964 2096
rect 3958 2091 3959 2095
rect 3963 2091 3964 2095
rect 3958 2090 3964 2091
rect 3895 2078 3899 2079
rect 3895 2073 3899 2074
rect 3896 2064 3898 2073
rect 3968 2072 3970 2110
rect 3992 2079 3994 2119
rect 3991 2078 3995 2079
rect 3991 2073 3995 2074
rect 3966 2071 3972 2072
rect 3966 2067 3967 2071
rect 3971 2067 3972 2071
rect 3966 2066 3972 2067
rect 3894 2063 3900 2064
rect 3894 2059 3895 2063
rect 3899 2059 3900 2063
rect 3894 2058 3900 2059
rect 3814 2055 3820 2056
rect 3814 2051 3815 2055
rect 3819 2051 3820 2055
rect 3814 2050 3820 2051
rect 3958 2055 3964 2056
rect 3958 2051 3959 2055
rect 3963 2051 3964 2055
rect 3958 2050 3964 2051
rect 3750 2022 3756 2023
rect 3750 2018 3751 2022
rect 3755 2018 3756 2022
rect 3750 2017 3756 2018
rect 3894 2022 3900 2023
rect 3894 2018 3895 2022
rect 3899 2018 3900 2022
rect 3894 2017 3900 2018
rect 3752 1995 3754 2017
rect 3896 1995 3898 2017
rect 3751 1994 3755 1995
rect 3751 1989 3755 1990
rect 3767 1994 3771 1995
rect 3767 1989 3771 1990
rect 3895 1994 3899 1995
rect 3895 1989 3899 1990
rect 3768 1979 3770 1989
rect 3896 1979 3898 1989
rect 3766 1978 3772 1979
rect 3766 1974 3767 1978
rect 3771 1974 3772 1978
rect 3766 1973 3772 1974
rect 3894 1978 3900 1979
rect 3894 1974 3895 1978
rect 3899 1974 3900 1978
rect 3894 1973 3900 1974
rect 3294 1947 3300 1948
rect 3294 1943 3295 1947
rect 3299 1943 3300 1947
rect 3294 1942 3300 1943
rect 3446 1947 3452 1948
rect 3446 1943 3447 1947
rect 3451 1943 3452 1947
rect 3446 1942 3452 1943
rect 3638 1947 3644 1948
rect 3638 1943 3639 1947
rect 3643 1943 3644 1947
rect 3638 1942 3644 1943
rect 3296 1928 3298 1942
rect 3310 1937 3316 1938
rect 3310 1933 3311 1937
rect 3315 1933 3316 1937
rect 3310 1932 3316 1933
rect 3254 1927 3260 1928
rect 3254 1923 3255 1927
rect 3259 1923 3260 1927
rect 3254 1922 3260 1923
rect 3294 1927 3300 1928
rect 3294 1923 3295 1927
rect 3299 1923 3300 1927
rect 3294 1922 3300 1923
rect 3312 1915 3314 1932
rect 3448 1920 3450 1942
rect 3462 1937 3468 1938
rect 3462 1933 3463 1937
rect 3467 1933 3468 1937
rect 3462 1932 3468 1933
rect 3614 1937 3620 1938
rect 3614 1933 3615 1937
rect 3619 1933 3620 1937
rect 3614 1932 3620 1933
rect 3766 1937 3772 1938
rect 3766 1933 3767 1937
rect 3771 1933 3772 1937
rect 3766 1932 3772 1933
rect 3894 1937 3900 1938
rect 3894 1933 3895 1937
rect 3899 1933 3900 1937
rect 3894 1932 3900 1933
rect 3446 1919 3452 1920
rect 3446 1915 3447 1919
rect 3451 1915 3452 1919
rect 3464 1915 3466 1932
rect 3616 1915 3618 1932
rect 3768 1915 3770 1932
rect 3774 1927 3780 1928
rect 3774 1923 3775 1927
rect 3779 1923 3780 1927
rect 3774 1922 3780 1923
rect 2071 1914 2075 1915
rect 2071 1909 2075 1910
rect 2279 1914 2283 1915
rect 2279 1909 2283 1910
rect 2407 1914 2411 1915
rect 2407 1909 2411 1910
rect 2463 1914 2467 1915
rect 2590 1911 2591 1915
rect 2595 1911 2596 1915
rect 2590 1910 2596 1911
rect 2639 1914 2643 1915
rect 2463 1909 2467 1910
rect 2639 1909 2643 1910
rect 2655 1914 2659 1915
rect 2655 1909 2659 1910
rect 2815 1914 2819 1915
rect 2815 1909 2819 1910
rect 2887 1914 2891 1915
rect 2887 1909 2891 1910
rect 2983 1914 2987 1915
rect 2983 1909 2987 1910
rect 3103 1914 3107 1915
rect 3103 1909 3107 1910
rect 3151 1914 3155 1915
rect 3151 1909 3155 1910
rect 3311 1914 3315 1915
rect 3446 1914 3452 1915
rect 3463 1914 3467 1915
rect 3311 1909 3315 1910
rect 3463 1909 3467 1910
rect 3511 1914 3515 1915
rect 3511 1909 3515 1910
rect 3615 1914 3619 1915
rect 3615 1909 3619 1910
rect 3711 1914 3715 1915
rect 3711 1909 3715 1910
rect 3767 1914 3771 1915
rect 3767 1909 3771 1910
rect 2030 1896 2036 1897
rect 2030 1892 2031 1896
rect 2035 1892 2036 1896
rect 2030 1891 2036 1892
rect 2072 1881 2074 1909
rect 2408 1900 2410 1909
rect 2656 1900 2658 1909
rect 2862 1907 2868 1908
rect 2862 1903 2863 1907
rect 2867 1903 2868 1907
rect 2862 1902 2868 1903
rect 2406 1899 2412 1900
rect 2406 1895 2407 1899
rect 2411 1895 2412 1899
rect 2406 1894 2412 1895
rect 2654 1899 2660 1900
rect 2654 1895 2655 1899
rect 2659 1895 2660 1899
rect 2654 1894 2660 1895
rect 2430 1887 2436 1888
rect 2430 1883 2431 1887
rect 2435 1883 2436 1887
rect 2430 1882 2436 1883
rect 2070 1880 2076 1881
rect 2030 1879 2036 1880
rect 2030 1875 2031 1879
rect 2035 1875 2036 1879
rect 2070 1876 2071 1880
rect 2075 1876 2076 1880
rect 2070 1875 2076 1876
rect 2030 1874 2036 1875
rect 2032 1851 2034 1874
rect 2070 1863 2076 1864
rect 2070 1859 2071 1863
rect 2075 1859 2076 1863
rect 2070 1858 2076 1859
rect 2406 1858 2412 1859
rect 2031 1850 2035 1851
rect 2031 1845 2035 1846
rect 2032 1830 2034 1845
rect 2072 1843 2074 1858
rect 2406 1854 2407 1858
rect 2411 1854 2412 1858
rect 2406 1853 2412 1854
rect 2408 1843 2410 1853
rect 2071 1842 2075 1843
rect 2071 1837 2075 1838
rect 2111 1842 2115 1843
rect 2111 1837 2115 1838
rect 2383 1842 2387 1843
rect 2383 1837 2387 1838
rect 2407 1842 2411 1843
rect 2407 1837 2411 1838
rect 2030 1829 2036 1830
rect 2030 1825 2031 1829
rect 2035 1825 2036 1829
rect 2030 1824 2036 1825
rect 2072 1822 2074 1837
rect 2112 1827 2114 1837
rect 2384 1827 2386 1837
rect 2110 1826 2116 1827
rect 2110 1822 2111 1826
rect 2115 1822 2116 1826
rect 2070 1821 2076 1822
rect 2110 1821 2116 1822
rect 2382 1826 2388 1827
rect 2382 1822 2383 1826
rect 2387 1822 2388 1826
rect 2382 1821 2388 1822
rect 2070 1817 2071 1821
rect 2075 1817 2076 1821
rect 2070 1816 2076 1817
rect 2030 1812 2036 1813
rect 2030 1808 2031 1812
rect 2035 1808 2036 1812
rect 2030 1807 2036 1808
rect 2006 1783 2012 1784
rect 2006 1779 2007 1783
rect 2011 1779 2012 1783
rect 2006 1778 2012 1779
rect 2032 1771 2034 1807
rect 2070 1804 2076 1805
rect 2062 1803 2068 1804
rect 2062 1799 2063 1803
rect 2067 1799 2068 1803
rect 2070 1800 2071 1804
rect 2075 1800 2076 1804
rect 2070 1799 2076 1800
rect 2062 1798 2068 1799
rect 2064 1776 2066 1798
rect 2062 1775 2068 1776
rect 2062 1771 2063 1775
rect 2067 1771 2068 1775
rect 2072 1771 2074 1799
rect 2182 1795 2188 1796
rect 2182 1791 2183 1795
rect 2187 1791 2188 1795
rect 2182 1790 2188 1791
rect 2110 1785 2116 1786
rect 2110 1781 2111 1785
rect 2115 1781 2116 1785
rect 2110 1780 2116 1781
rect 2112 1771 2114 1780
rect 1935 1770 1939 1771
rect 1935 1765 1939 1766
rect 2031 1770 2035 1771
rect 2062 1770 2068 1771
rect 2071 1770 2075 1771
rect 2031 1765 2035 1766
rect 2071 1765 2075 1766
rect 2111 1770 2115 1771
rect 2111 1765 2115 1766
rect 1743 1748 1747 1749
rect 1743 1743 1747 1744
rect 2032 1737 2034 1765
rect 2072 1737 2074 1765
rect 2112 1756 2114 1765
rect 2184 1764 2186 1790
rect 2382 1785 2388 1786
rect 2382 1781 2383 1785
rect 2387 1781 2388 1785
rect 2382 1780 2388 1781
rect 2384 1771 2386 1780
rect 2432 1776 2434 1882
rect 2654 1858 2660 1859
rect 2654 1854 2655 1858
rect 2659 1854 2660 1858
rect 2654 1853 2660 1854
rect 2656 1843 2658 1853
rect 2647 1842 2651 1843
rect 2647 1837 2651 1838
rect 2655 1842 2659 1843
rect 2655 1837 2659 1838
rect 2648 1827 2650 1837
rect 2646 1826 2652 1827
rect 2646 1822 2647 1826
rect 2651 1822 2652 1826
rect 2646 1821 2652 1822
rect 2864 1796 2866 1902
rect 2888 1900 2890 1909
rect 3104 1900 3106 1909
rect 3312 1900 3314 1909
rect 3512 1900 3514 1909
rect 3606 1907 3612 1908
rect 3606 1903 3607 1907
rect 3611 1903 3612 1907
rect 3606 1902 3612 1903
rect 2886 1899 2892 1900
rect 2886 1895 2887 1899
rect 2891 1895 2892 1899
rect 2886 1894 2892 1895
rect 3102 1899 3108 1900
rect 3102 1895 3103 1899
rect 3107 1895 3108 1899
rect 3102 1894 3108 1895
rect 3310 1899 3316 1900
rect 3310 1895 3311 1899
rect 3315 1895 3316 1899
rect 3310 1894 3316 1895
rect 3510 1899 3516 1900
rect 3510 1895 3511 1899
rect 3515 1895 3516 1899
rect 3510 1894 3516 1895
rect 3166 1891 3172 1892
rect 3166 1887 3167 1891
rect 3171 1887 3172 1891
rect 3166 1886 3172 1887
rect 2886 1858 2892 1859
rect 2886 1854 2887 1858
rect 2891 1854 2892 1858
rect 2886 1853 2892 1854
rect 3102 1858 3108 1859
rect 3102 1854 3103 1858
rect 3107 1854 3108 1858
rect 3102 1853 3108 1854
rect 2888 1843 2890 1853
rect 3104 1843 3106 1853
rect 2887 1842 2891 1843
rect 2887 1837 2891 1838
rect 3095 1842 3099 1843
rect 3095 1837 3099 1838
rect 3103 1842 3107 1843
rect 3103 1837 3107 1838
rect 2888 1827 2890 1837
rect 3096 1827 3098 1837
rect 2886 1826 2892 1827
rect 2886 1822 2887 1826
rect 2891 1822 2892 1826
rect 2886 1821 2892 1822
rect 3094 1826 3100 1827
rect 3094 1822 3095 1826
rect 3099 1822 3100 1826
rect 3094 1821 3100 1822
rect 2578 1795 2584 1796
rect 2578 1791 2579 1795
rect 2583 1791 2584 1795
rect 2578 1790 2584 1791
rect 2862 1795 2868 1796
rect 2862 1791 2863 1795
rect 2867 1791 2868 1795
rect 2862 1790 2868 1791
rect 3078 1795 3084 1796
rect 3078 1791 3079 1795
rect 3083 1791 3084 1795
rect 3078 1790 3084 1791
rect 2430 1775 2436 1776
rect 2430 1771 2431 1775
rect 2435 1771 2436 1775
rect 2287 1770 2291 1771
rect 2287 1765 2291 1766
rect 2383 1770 2387 1771
rect 2430 1770 2436 1771
rect 2495 1770 2499 1771
rect 2383 1765 2387 1766
rect 2495 1765 2499 1766
rect 2182 1763 2188 1764
rect 2182 1759 2183 1763
rect 2187 1759 2188 1763
rect 2182 1758 2188 1759
rect 2288 1756 2290 1765
rect 2496 1756 2498 1765
rect 2580 1764 2582 1790
rect 2646 1785 2652 1786
rect 2646 1781 2647 1785
rect 2651 1781 2652 1785
rect 2646 1780 2652 1781
rect 2886 1785 2892 1786
rect 2886 1781 2887 1785
rect 2891 1781 2892 1785
rect 2886 1780 2892 1781
rect 2648 1771 2650 1780
rect 2888 1771 2890 1780
rect 2647 1770 2651 1771
rect 2647 1765 2651 1766
rect 2711 1770 2715 1771
rect 2711 1765 2715 1766
rect 2887 1770 2891 1771
rect 2887 1765 2891 1766
rect 2919 1770 2923 1771
rect 3080 1768 3082 1790
rect 3094 1785 3100 1786
rect 3094 1781 3095 1785
rect 3099 1781 3100 1785
rect 3094 1780 3100 1781
rect 3096 1771 3098 1780
rect 3168 1776 3170 1886
rect 3310 1858 3316 1859
rect 3310 1854 3311 1858
rect 3315 1854 3316 1858
rect 3310 1853 3316 1854
rect 3510 1858 3516 1859
rect 3510 1854 3511 1858
rect 3515 1854 3516 1858
rect 3510 1853 3516 1854
rect 3312 1843 3314 1853
rect 3512 1843 3514 1853
rect 3287 1842 3291 1843
rect 3287 1837 3291 1838
rect 3311 1842 3315 1843
rect 3311 1837 3315 1838
rect 3455 1842 3459 1843
rect 3455 1837 3459 1838
rect 3511 1842 3515 1843
rect 3511 1837 3515 1838
rect 3288 1827 3290 1837
rect 3456 1827 3458 1837
rect 3286 1826 3292 1827
rect 3286 1822 3287 1826
rect 3291 1822 3292 1826
rect 3286 1821 3292 1822
rect 3454 1826 3460 1827
rect 3454 1822 3455 1826
rect 3459 1822 3460 1826
rect 3454 1821 3460 1822
rect 3608 1796 3610 1902
rect 3712 1900 3714 1909
rect 3710 1899 3716 1900
rect 3710 1895 3711 1899
rect 3715 1895 3716 1899
rect 3710 1894 3716 1895
rect 3776 1892 3778 1922
rect 3896 1915 3898 1932
rect 3960 1928 3962 2050
rect 3992 2045 3994 2073
rect 3990 2044 3996 2045
rect 3990 2040 3991 2044
rect 3995 2040 3996 2044
rect 3990 2039 3996 2040
rect 3990 2027 3996 2028
rect 3990 2023 3991 2027
rect 3995 2023 3996 2027
rect 3990 2022 3996 2023
rect 3992 1995 3994 2022
rect 3991 1994 3995 1995
rect 3991 1989 3995 1990
rect 3992 1974 3994 1989
rect 3990 1973 3996 1974
rect 3990 1969 3991 1973
rect 3995 1969 3996 1973
rect 3990 1968 3996 1969
rect 3990 1956 3996 1957
rect 3990 1952 3991 1956
rect 3995 1952 3996 1956
rect 3990 1951 3996 1952
rect 3966 1947 3972 1948
rect 3966 1943 3967 1947
rect 3971 1943 3972 1947
rect 3966 1942 3972 1943
rect 3958 1927 3964 1928
rect 3958 1923 3959 1927
rect 3963 1923 3964 1927
rect 3958 1922 3964 1923
rect 3895 1914 3899 1915
rect 3895 1909 3899 1910
rect 3896 1900 3898 1909
rect 3968 1908 3970 1942
rect 3992 1915 3994 1951
rect 3991 1914 3995 1915
rect 3991 1909 3995 1910
rect 3966 1907 3972 1908
rect 3966 1903 3967 1907
rect 3971 1903 3972 1907
rect 3966 1902 3972 1903
rect 3894 1899 3900 1900
rect 3894 1895 3895 1899
rect 3899 1895 3900 1899
rect 3894 1894 3900 1895
rect 3774 1891 3780 1892
rect 3774 1887 3775 1891
rect 3779 1887 3780 1891
rect 3774 1886 3780 1887
rect 3886 1887 3892 1888
rect 3886 1883 3887 1887
rect 3891 1883 3892 1887
rect 3886 1882 3892 1883
rect 3710 1858 3716 1859
rect 3710 1854 3711 1858
rect 3715 1854 3716 1858
rect 3710 1853 3716 1854
rect 3712 1843 3714 1853
rect 3615 1842 3619 1843
rect 3615 1837 3619 1838
rect 3711 1842 3715 1843
rect 3711 1837 3715 1838
rect 3767 1842 3771 1843
rect 3767 1837 3771 1838
rect 3616 1827 3618 1837
rect 3768 1827 3770 1837
rect 3614 1826 3620 1827
rect 3614 1822 3615 1826
rect 3619 1822 3620 1826
rect 3614 1821 3620 1822
rect 3766 1826 3772 1827
rect 3766 1822 3767 1826
rect 3771 1822 3772 1826
rect 3766 1821 3772 1822
rect 3358 1795 3364 1796
rect 3358 1791 3359 1795
rect 3363 1791 3364 1795
rect 3358 1790 3364 1791
rect 3562 1795 3568 1796
rect 3562 1791 3563 1795
rect 3567 1791 3568 1795
rect 3562 1790 3568 1791
rect 3606 1795 3612 1796
rect 3606 1791 3607 1795
rect 3611 1791 3612 1795
rect 3606 1790 3612 1791
rect 3286 1785 3292 1786
rect 3286 1781 3287 1785
rect 3291 1781 3292 1785
rect 3286 1780 3292 1781
rect 3166 1775 3172 1776
rect 3166 1771 3167 1775
rect 3171 1771 3172 1775
rect 3288 1771 3290 1780
rect 3095 1770 3099 1771
rect 2919 1765 2923 1766
rect 3078 1767 3084 1768
rect 2578 1763 2584 1764
rect 2578 1759 2579 1763
rect 2583 1759 2584 1763
rect 2578 1758 2584 1759
rect 2712 1756 2714 1765
rect 2920 1756 2922 1765
rect 2990 1763 2996 1764
rect 2990 1759 2991 1763
rect 2995 1759 2996 1763
rect 3078 1763 3079 1767
rect 3083 1763 3084 1767
rect 3095 1765 3099 1766
rect 3119 1770 3123 1771
rect 3166 1770 3172 1771
rect 3287 1770 3291 1771
rect 3119 1765 3123 1766
rect 3287 1765 3291 1766
rect 3319 1770 3323 1771
rect 3319 1765 3323 1766
rect 3078 1762 3084 1763
rect 2990 1758 2996 1759
rect 2110 1755 2116 1756
rect 2110 1751 2111 1755
rect 2115 1751 2116 1755
rect 2110 1750 2116 1751
rect 2286 1755 2292 1756
rect 2286 1751 2287 1755
rect 2291 1751 2292 1755
rect 2286 1750 2292 1751
rect 2494 1755 2500 1756
rect 2494 1751 2495 1755
rect 2499 1751 2500 1755
rect 2494 1750 2500 1751
rect 2710 1755 2716 1756
rect 2710 1751 2711 1755
rect 2715 1751 2716 1755
rect 2710 1750 2716 1751
rect 2918 1755 2924 1756
rect 2918 1751 2919 1755
rect 2923 1751 2924 1755
rect 2918 1750 2924 1751
rect 2486 1743 2492 1744
rect 2486 1739 2487 1743
rect 2491 1739 2492 1743
rect 2486 1738 2492 1739
rect 2726 1743 2732 1744
rect 2726 1739 2727 1743
rect 2731 1739 2732 1743
rect 2726 1738 2732 1739
rect 2030 1736 2036 1737
rect 2030 1732 2031 1736
rect 2035 1732 2036 1736
rect 2030 1731 2036 1732
rect 2070 1736 2076 1737
rect 2070 1732 2071 1736
rect 2075 1732 2076 1736
rect 2070 1731 2076 1732
rect 2030 1719 2036 1720
rect 2030 1715 2031 1719
rect 2035 1715 2036 1719
rect 2030 1714 2036 1715
rect 2070 1719 2076 1720
rect 2070 1715 2071 1719
rect 2075 1715 2076 1719
rect 2070 1714 2076 1715
rect 2110 1714 2116 1715
rect 2032 1699 2034 1714
rect 1743 1698 1747 1699
rect 1743 1693 1747 1694
rect 1927 1698 1931 1699
rect 1927 1693 1931 1694
rect 2031 1698 2035 1699
rect 2031 1693 2035 1694
rect 1744 1683 1746 1693
rect 1928 1683 1930 1693
rect 1742 1682 1748 1683
rect 1742 1678 1743 1682
rect 1747 1678 1748 1682
rect 1742 1677 1748 1678
rect 1926 1682 1932 1683
rect 1926 1678 1927 1682
rect 1931 1678 1932 1682
rect 2032 1678 2034 1693
rect 2072 1691 2074 1714
rect 2110 1710 2111 1714
rect 2115 1710 2116 1714
rect 2110 1709 2116 1710
rect 2286 1714 2292 1715
rect 2286 1710 2287 1714
rect 2291 1710 2292 1714
rect 2286 1709 2292 1710
rect 2112 1691 2114 1709
rect 2288 1691 2290 1709
rect 2071 1690 2075 1691
rect 2071 1685 2075 1686
rect 2111 1690 2115 1691
rect 2111 1685 2115 1686
rect 2239 1690 2243 1691
rect 2239 1685 2243 1686
rect 2287 1690 2291 1691
rect 2287 1685 2291 1686
rect 2383 1690 2387 1691
rect 2383 1685 2387 1686
rect 1926 1677 1932 1678
rect 2030 1677 2036 1678
rect 2030 1673 2031 1677
rect 2035 1673 2036 1677
rect 2030 1672 2036 1673
rect 1702 1671 1708 1672
rect 1702 1667 1703 1671
rect 1707 1667 1708 1671
rect 2072 1670 2074 1685
rect 2112 1675 2114 1685
rect 2240 1675 2242 1685
rect 2384 1675 2386 1685
rect 2110 1674 2116 1675
rect 2110 1670 2111 1674
rect 2115 1670 2116 1674
rect 1702 1666 1708 1667
rect 2070 1669 2076 1670
rect 2110 1669 2116 1670
rect 2238 1674 2244 1675
rect 2238 1670 2239 1674
rect 2243 1670 2244 1674
rect 2238 1669 2244 1670
rect 2382 1674 2388 1675
rect 2382 1670 2383 1674
rect 2387 1670 2388 1674
rect 2382 1669 2388 1670
rect 2070 1665 2071 1669
rect 2075 1665 2076 1669
rect 2070 1664 2076 1665
rect 2030 1660 2036 1661
rect 2030 1656 2031 1660
rect 2035 1656 2036 1660
rect 2030 1655 2036 1656
rect 386 1651 392 1652
rect 386 1647 387 1651
rect 391 1647 392 1651
rect 386 1646 392 1647
rect 750 1651 756 1652
rect 750 1647 751 1651
rect 755 1647 756 1651
rect 750 1646 756 1647
rect 790 1651 796 1652
rect 790 1647 791 1651
rect 795 1647 796 1651
rect 790 1646 796 1647
rect 1006 1651 1012 1652
rect 1006 1647 1007 1651
rect 1011 1647 1012 1651
rect 1006 1646 1012 1647
rect 388 1632 390 1646
rect 534 1641 540 1642
rect 534 1637 535 1641
rect 539 1637 540 1641
rect 534 1636 540 1637
rect 366 1631 372 1632
rect 366 1627 367 1631
rect 371 1627 372 1631
rect 366 1626 372 1627
rect 386 1631 392 1632
rect 386 1627 387 1631
rect 391 1627 392 1631
rect 386 1626 392 1627
rect 536 1623 538 1636
rect 752 1632 754 1646
rect 766 1641 772 1642
rect 766 1637 767 1641
rect 771 1637 772 1641
rect 766 1636 772 1637
rect 750 1631 756 1632
rect 750 1627 751 1631
rect 755 1627 756 1631
rect 750 1626 756 1627
rect 768 1623 770 1636
rect 111 1622 115 1623
rect 111 1617 115 1618
rect 303 1622 307 1623
rect 303 1617 307 1618
rect 399 1622 403 1623
rect 399 1617 403 1618
rect 535 1622 539 1623
rect 535 1617 539 1618
rect 575 1622 579 1623
rect 575 1617 579 1618
rect 751 1622 755 1623
rect 751 1617 755 1618
rect 767 1622 771 1623
rect 767 1617 771 1618
rect 112 1589 114 1617
rect 400 1608 402 1617
rect 576 1608 578 1617
rect 752 1608 754 1617
rect 792 1616 794 1646
rect 982 1641 988 1642
rect 982 1637 983 1641
rect 987 1637 988 1641
rect 982 1636 988 1637
rect 1190 1641 1196 1642
rect 1190 1637 1191 1641
rect 1195 1637 1196 1641
rect 1190 1636 1196 1637
rect 1382 1641 1388 1642
rect 1382 1637 1383 1641
rect 1387 1637 1388 1641
rect 1382 1636 1388 1637
rect 1566 1641 1572 1642
rect 1566 1637 1567 1641
rect 1571 1637 1572 1641
rect 1566 1636 1572 1637
rect 1742 1641 1748 1642
rect 1742 1637 1743 1641
rect 1747 1637 1748 1641
rect 1742 1636 1748 1637
rect 1926 1641 1932 1642
rect 1926 1637 1927 1641
rect 1931 1637 1932 1641
rect 1926 1636 1932 1637
rect 984 1623 986 1636
rect 1192 1623 1194 1636
rect 1384 1623 1386 1636
rect 1430 1623 1436 1624
rect 1568 1623 1570 1636
rect 1744 1623 1746 1636
rect 1928 1623 1930 1636
rect 1998 1631 2004 1632
rect 1998 1627 1999 1631
rect 2003 1627 2004 1631
rect 1998 1626 2004 1627
rect 935 1622 939 1623
rect 935 1617 939 1618
rect 983 1622 987 1623
rect 983 1617 987 1618
rect 1111 1622 1115 1623
rect 1111 1617 1115 1618
rect 1191 1622 1195 1623
rect 1191 1617 1195 1618
rect 1279 1622 1283 1623
rect 1279 1617 1283 1618
rect 1383 1622 1387 1623
rect 1430 1619 1431 1623
rect 1435 1619 1436 1623
rect 1430 1618 1436 1619
rect 1447 1622 1451 1623
rect 1383 1617 1387 1618
rect 790 1615 796 1616
rect 790 1611 791 1615
rect 795 1611 796 1615
rect 790 1610 796 1611
rect 936 1608 938 1617
rect 990 1615 996 1616
rect 990 1611 991 1615
rect 995 1611 996 1615
rect 990 1610 996 1611
rect 398 1607 404 1608
rect 398 1603 399 1607
rect 403 1603 404 1607
rect 398 1602 404 1603
rect 574 1607 580 1608
rect 574 1603 575 1607
rect 579 1603 580 1607
rect 574 1602 580 1603
rect 750 1607 756 1608
rect 750 1603 751 1607
rect 755 1603 756 1607
rect 750 1602 756 1603
rect 934 1607 940 1608
rect 934 1603 935 1607
rect 939 1603 940 1607
rect 934 1602 940 1603
rect 558 1599 564 1600
rect 558 1595 559 1599
rect 563 1595 564 1599
rect 558 1594 564 1595
rect 110 1588 116 1589
rect 110 1584 111 1588
rect 115 1584 116 1588
rect 110 1583 116 1584
rect 110 1571 116 1572
rect 110 1567 111 1571
rect 115 1567 116 1571
rect 110 1566 116 1567
rect 398 1566 404 1567
rect 112 1543 114 1566
rect 398 1562 399 1566
rect 403 1562 404 1566
rect 398 1561 404 1562
rect 400 1543 402 1561
rect 111 1542 115 1543
rect 111 1537 115 1538
rect 399 1542 403 1543
rect 399 1537 403 1538
rect 503 1542 507 1543
rect 503 1537 507 1538
rect 112 1522 114 1537
rect 504 1527 506 1537
rect 502 1526 508 1527
rect 502 1522 503 1526
rect 507 1522 508 1526
rect 110 1521 116 1522
rect 502 1521 508 1522
rect 110 1517 111 1521
rect 115 1517 116 1521
rect 110 1516 116 1517
rect 110 1504 116 1505
rect 110 1500 111 1504
rect 115 1500 116 1504
rect 110 1499 116 1500
rect 112 1459 114 1499
rect 502 1485 508 1486
rect 502 1481 503 1485
rect 507 1481 508 1485
rect 502 1480 508 1481
rect 504 1459 506 1480
rect 560 1476 562 1594
rect 574 1566 580 1567
rect 574 1562 575 1566
rect 579 1562 580 1566
rect 574 1561 580 1562
rect 750 1566 756 1567
rect 750 1562 751 1566
rect 755 1562 756 1566
rect 750 1561 756 1562
rect 934 1566 940 1567
rect 934 1562 935 1566
rect 939 1562 940 1566
rect 934 1561 940 1562
rect 576 1543 578 1561
rect 752 1543 754 1561
rect 936 1543 938 1561
rect 575 1542 579 1543
rect 575 1537 579 1538
rect 615 1542 619 1543
rect 615 1537 619 1538
rect 735 1542 739 1543
rect 735 1537 739 1538
rect 751 1542 755 1543
rect 751 1537 755 1538
rect 855 1542 859 1543
rect 855 1537 859 1538
rect 935 1542 939 1543
rect 935 1537 939 1538
rect 967 1542 971 1543
rect 967 1537 971 1538
rect 616 1527 618 1537
rect 736 1527 738 1537
rect 856 1527 858 1537
rect 968 1527 970 1537
rect 614 1526 620 1527
rect 614 1522 615 1526
rect 619 1522 620 1526
rect 614 1521 620 1522
rect 734 1526 740 1527
rect 734 1522 735 1526
rect 739 1522 740 1526
rect 734 1521 740 1522
rect 854 1526 860 1527
rect 854 1522 855 1526
rect 859 1522 860 1526
rect 854 1521 860 1522
rect 966 1526 972 1527
rect 966 1522 967 1526
rect 971 1522 972 1526
rect 966 1521 972 1522
rect 992 1496 994 1610
rect 1112 1608 1114 1617
rect 1280 1608 1282 1617
rect 1110 1607 1116 1608
rect 1110 1603 1111 1607
rect 1115 1603 1116 1607
rect 1110 1602 1116 1603
rect 1278 1607 1284 1608
rect 1278 1603 1279 1607
rect 1283 1603 1284 1607
rect 1278 1602 1284 1603
rect 1432 1600 1434 1618
rect 1447 1617 1451 1618
rect 1567 1622 1571 1623
rect 1567 1617 1571 1618
rect 1607 1622 1611 1623
rect 1607 1617 1611 1618
rect 1743 1622 1747 1623
rect 1743 1617 1747 1618
rect 1767 1622 1771 1623
rect 1767 1617 1771 1618
rect 1927 1622 1931 1623
rect 1927 1617 1931 1618
rect 1935 1622 1939 1623
rect 1935 1617 1939 1618
rect 1448 1608 1450 1617
rect 1550 1615 1556 1616
rect 1550 1611 1551 1615
rect 1555 1611 1556 1615
rect 1550 1610 1556 1611
rect 1446 1607 1452 1608
rect 1446 1603 1447 1607
rect 1451 1603 1452 1607
rect 1446 1602 1452 1603
rect 1430 1599 1436 1600
rect 1430 1595 1431 1599
rect 1435 1595 1436 1599
rect 1430 1594 1436 1595
rect 1110 1566 1116 1567
rect 1110 1562 1111 1566
rect 1115 1562 1116 1566
rect 1110 1561 1116 1562
rect 1278 1566 1284 1567
rect 1278 1562 1279 1566
rect 1283 1562 1284 1566
rect 1278 1561 1284 1562
rect 1446 1566 1452 1567
rect 1446 1562 1447 1566
rect 1451 1562 1452 1566
rect 1446 1561 1452 1562
rect 1112 1543 1114 1561
rect 1280 1543 1282 1561
rect 1448 1543 1450 1561
rect 1079 1542 1083 1543
rect 1079 1537 1083 1538
rect 1111 1542 1115 1543
rect 1111 1537 1115 1538
rect 1199 1542 1203 1543
rect 1199 1537 1203 1538
rect 1279 1542 1283 1543
rect 1279 1537 1283 1538
rect 1319 1542 1323 1543
rect 1319 1537 1323 1538
rect 1439 1542 1443 1543
rect 1439 1537 1443 1538
rect 1447 1542 1451 1543
rect 1447 1537 1451 1538
rect 1080 1527 1082 1537
rect 1200 1527 1202 1537
rect 1320 1527 1322 1537
rect 1440 1527 1442 1537
rect 1078 1526 1084 1527
rect 1078 1522 1079 1526
rect 1083 1522 1084 1526
rect 1078 1521 1084 1522
rect 1198 1526 1204 1527
rect 1198 1522 1199 1526
rect 1203 1522 1204 1526
rect 1198 1521 1204 1522
rect 1318 1526 1324 1527
rect 1318 1522 1319 1526
rect 1323 1522 1324 1526
rect 1318 1521 1324 1522
rect 1438 1526 1444 1527
rect 1438 1522 1439 1526
rect 1443 1522 1444 1526
rect 1438 1521 1444 1522
rect 1552 1496 1554 1610
rect 1608 1608 1610 1617
rect 1768 1608 1770 1617
rect 1936 1608 1938 1617
rect 1606 1607 1612 1608
rect 1606 1603 1607 1607
rect 1611 1603 1612 1607
rect 1606 1602 1612 1603
rect 1766 1607 1772 1608
rect 1766 1603 1767 1607
rect 1771 1603 1772 1607
rect 1766 1602 1772 1603
rect 1934 1607 1940 1608
rect 1934 1603 1935 1607
rect 1939 1603 1940 1607
rect 1934 1602 1940 1603
rect 2000 1600 2002 1626
rect 2032 1623 2034 1655
rect 2070 1652 2076 1653
rect 2070 1648 2071 1652
rect 2075 1648 2076 1652
rect 2070 1647 2076 1648
rect 2031 1622 2035 1623
rect 2031 1617 2035 1618
rect 1998 1599 2004 1600
rect 1998 1595 1999 1599
rect 2003 1595 2004 1599
rect 1998 1594 2004 1595
rect 2032 1589 2034 1617
rect 2072 1607 2074 1647
rect 2182 1643 2188 1644
rect 2182 1639 2183 1643
rect 2187 1639 2188 1643
rect 2182 1638 2188 1639
rect 2110 1633 2116 1634
rect 2110 1629 2111 1633
rect 2115 1629 2116 1633
rect 2110 1628 2116 1629
rect 2112 1607 2114 1628
rect 2071 1606 2075 1607
rect 2071 1601 2075 1602
rect 2111 1606 2115 1607
rect 2111 1601 2115 1602
rect 2167 1606 2171 1607
rect 2167 1601 2171 1602
rect 2030 1588 2036 1589
rect 2030 1584 2031 1588
rect 2035 1584 2036 1588
rect 2030 1583 2036 1584
rect 2072 1573 2074 1601
rect 2168 1592 2170 1601
rect 2184 1600 2186 1638
rect 2238 1633 2244 1634
rect 2238 1629 2239 1633
rect 2243 1629 2244 1633
rect 2238 1628 2244 1629
rect 2382 1633 2388 1634
rect 2382 1629 2383 1633
rect 2387 1629 2388 1633
rect 2382 1628 2388 1629
rect 2240 1607 2242 1628
rect 2384 1607 2386 1628
rect 2488 1624 2490 1738
rect 2494 1714 2500 1715
rect 2494 1710 2495 1714
rect 2499 1710 2500 1714
rect 2494 1709 2500 1710
rect 2710 1714 2716 1715
rect 2710 1710 2711 1714
rect 2715 1710 2716 1714
rect 2710 1709 2716 1710
rect 2496 1691 2498 1709
rect 2712 1691 2714 1709
rect 2495 1690 2499 1691
rect 2495 1685 2499 1686
rect 2519 1690 2523 1691
rect 2519 1685 2523 1686
rect 2655 1690 2659 1691
rect 2655 1685 2659 1686
rect 2711 1690 2715 1691
rect 2711 1685 2715 1686
rect 2520 1675 2522 1685
rect 2656 1675 2658 1685
rect 2518 1674 2524 1675
rect 2518 1670 2519 1674
rect 2523 1670 2524 1674
rect 2518 1669 2524 1670
rect 2654 1674 2660 1675
rect 2654 1670 2655 1674
rect 2659 1670 2660 1674
rect 2654 1669 2660 1670
rect 2614 1643 2620 1644
rect 2614 1639 2615 1643
rect 2619 1639 2620 1643
rect 2614 1638 2620 1639
rect 2518 1633 2524 1634
rect 2518 1629 2519 1633
rect 2523 1629 2524 1633
rect 2518 1628 2524 1629
rect 2486 1623 2492 1624
rect 2486 1619 2487 1623
rect 2491 1619 2492 1623
rect 2486 1618 2492 1619
rect 2520 1607 2522 1628
rect 2239 1606 2243 1607
rect 2239 1601 2243 1602
rect 2287 1606 2291 1607
rect 2287 1601 2291 1602
rect 2383 1606 2387 1607
rect 2383 1601 2387 1602
rect 2407 1606 2411 1607
rect 2407 1601 2411 1602
rect 2519 1606 2523 1607
rect 2519 1601 2523 1602
rect 2527 1606 2531 1607
rect 2527 1601 2531 1602
rect 2182 1599 2188 1600
rect 2182 1595 2183 1599
rect 2187 1595 2188 1599
rect 2182 1594 2188 1595
rect 2288 1592 2290 1601
rect 2408 1592 2410 1601
rect 2528 1592 2530 1601
rect 2616 1600 2618 1638
rect 2654 1633 2660 1634
rect 2654 1629 2655 1633
rect 2659 1629 2660 1633
rect 2654 1628 2660 1629
rect 2656 1607 2658 1628
rect 2728 1624 2730 1738
rect 2918 1714 2924 1715
rect 2918 1710 2919 1714
rect 2923 1710 2924 1714
rect 2918 1709 2924 1710
rect 2920 1691 2922 1709
rect 2791 1690 2795 1691
rect 2791 1685 2795 1686
rect 2919 1690 2923 1691
rect 2919 1685 2923 1686
rect 2927 1690 2931 1691
rect 2927 1685 2931 1686
rect 2792 1675 2794 1685
rect 2928 1675 2930 1685
rect 2790 1674 2796 1675
rect 2790 1670 2791 1674
rect 2795 1670 2796 1674
rect 2790 1669 2796 1670
rect 2926 1674 2932 1675
rect 2926 1670 2927 1674
rect 2931 1670 2932 1674
rect 2926 1669 2932 1670
rect 2910 1643 2916 1644
rect 2910 1639 2911 1643
rect 2915 1639 2916 1643
rect 2992 1640 2994 1758
rect 3120 1756 3122 1765
rect 3320 1756 3322 1765
rect 3360 1764 3362 1790
rect 3454 1785 3460 1786
rect 3454 1781 3455 1785
rect 3459 1781 3460 1785
rect 3454 1780 3460 1781
rect 3456 1771 3458 1780
rect 3564 1776 3566 1790
rect 3614 1785 3620 1786
rect 3614 1781 3615 1785
rect 3619 1781 3620 1785
rect 3614 1780 3620 1781
rect 3766 1785 3772 1786
rect 3766 1781 3767 1785
rect 3771 1781 3772 1785
rect 3766 1780 3772 1781
rect 3526 1775 3532 1776
rect 3526 1771 3527 1775
rect 3531 1771 3532 1775
rect 3455 1770 3459 1771
rect 3455 1765 3459 1766
rect 3511 1770 3515 1771
rect 3526 1770 3532 1771
rect 3562 1775 3568 1776
rect 3562 1771 3563 1775
rect 3567 1771 3568 1775
rect 3616 1771 3618 1780
rect 3768 1771 3770 1780
rect 3888 1776 3890 1882
rect 3992 1881 3994 1909
rect 3990 1880 3996 1881
rect 3990 1876 3991 1880
rect 3995 1876 3996 1880
rect 3990 1875 3996 1876
rect 3990 1863 3996 1864
rect 3990 1859 3991 1863
rect 3995 1859 3996 1863
rect 3894 1858 3900 1859
rect 3990 1858 3996 1859
rect 3894 1854 3895 1858
rect 3899 1854 3900 1858
rect 3894 1853 3900 1854
rect 3896 1843 3898 1853
rect 3992 1843 3994 1858
rect 3895 1842 3899 1843
rect 3895 1837 3899 1838
rect 3991 1842 3995 1843
rect 3991 1837 3995 1838
rect 3896 1827 3898 1837
rect 3894 1826 3900 1827
rect 3894 1822 3895 1826
rect 3899 1822 3900 1826
rect 3992 1822 3994 1837
rect 3894 1821 3900 1822
rect 3990 1821 3996 1822
rect 3990 1817 3991 1821
rect 3995 1817 3996 1821
rect 3990 1816 3996 1817
rect 3990 1804 3996 1805
rect 3902 1803 3908 1804
rect 3902 1799 3903 1803
rect 3907 1799 3908 1803
rect 3990 1800 3991 1804
rect 3995 1800 3996 1804
rect 3990 1799 3996 1800
rect 3902 1798 3908 1799
rect 3894 1785 3900 1786
rect 3894 1781 3895 1785
rect 3899 1781 3900 1785
rect 3894 1780 3900 1781
rect 3886 1775 3892 1776
rect 3886 1771 3887 1775
rect 3891 1771 3892 1775
rect 3896 1771 3898 1780
rect 3904 1776 3906 1798
rect 3966 1795 3972 1796
rect 3966 1791 3967 1795
rect 3971 1791 3972 1795
rect 3966 1790 3972 1791
rect 3902 1775 3908 1776
rect 3902 1771 3903 1775
rect 3907 1771 3908 1775
rect 3562 1770 3568 1771
rect 3615 1770 3619 1771
rect 3511 1765 3515 1766
rect 3358 1763 3364 1764
rect 3358 1759 3359 1763
rect 3363 1759 3364 1763
rect 3358 1758 3364 1759
rect 3512 1756 3514 1765
rect 3118 1755 3124 1756
rect 3118 1751 3119 1755
rect 3123 1751 3124 1755
rect 3118 1750 3124 1751
rect 3318 1755 3324 1756
rect 3318 1751 3319 1755
rect 3323 1751 3324 1755
rect 3318 1750 3324 1751
rect 3510 1755 3516 1756
rect 3510 1751 3511 1755
rect 3515 1751 3516 1755
rect 3510 1750 3516 1751
rect 3528 1744 3530 1770
rect 3615 1765 3619 1766
rect 3703 1770 3707 1771
rect 3703 1765 3707 1766
rect 3767 1770 3771 1771
rect 3886 1770 3892 1771
rect 3895 1770 3899 1771
rect 3902 1770 3908 1771
rect 3767 1765 3771 1766
rect 3895 1765 3899 1766
rect 3704 1756 3706 1765
rect 3896 1756 3898 1765
rect 3968 1764 3970 1790
rect 3992 1771 3994 1799
rect 3991 1770 3995 1771
rect 3991 1765 3995 1766
rect 3966 1763 3972 1764
rect 3966 1759 3967 1763
rect 3971 1759 3972 1763
rect 3966 1758 3972 1759
rect 3702 1755 3708 1756
rect 3702 1751 3703 1755
rect 3707 1751 3708 1755
rect 3702 1750 3708 1751
rect 3894 1755 3900 1756
rect 3894 1751 3895 1755
rect 3899 1751 3900 1755
rect 3894 1750 3900 1751
rect 3134 1743 3140 1744
rect 3134 1739 3135 1743
rect 3139 1739 3140 1743
rect 3134 1738 3140 1739
rect 3526 1743 3532 1744
rect 3526 1739 3527 1743
rect 3531 1739 3532 1743
rect 3526 1738 3532 1739
rect 3118 1714 3124 1715
rect 3118 1710 3119 1714
rect 3123 1710 3124 1714
rect 3118 1709 3124 1710
rect 3120 1691 3122 1709
rect 3063 1690 3067 1691
rect 3063 1685 3067 1686
rect 3119 1690 3123 1691
rect 3119 1685 3123 1686
rect 3064 1675 3066 1685
rect 3062 1674 3068 1675
rect 3062 1670 3063 1674
rect 3067 1670 3068 1674
rect 3062 1669 3068 1670
rect 2910 1638 2916 1639
rect 2990 1639 2996 1640
rect 2790 1633 2796 1634
rect 2790 1629 2791 1633
rect 2795 1629 2796 1633
rect 2790 1628 2796 1629
rect 2726 1623 2732 1624
rect 2726 1619 2727 1623
rect 2731 1619 2732 1623
rect 2726 1618 2732 1619
rect 2792 1607 2794 1628
rect 2912 1624 2914 1638
rect 2990 1635 2991 1639
rect 2995 1635 2996 1639
rect 2990 1634 2996 1635
rect 2926 1633 2932 1634
rect 2926 1629 2927 1633
rect 2931 1629 2932 1633
rect 2926 1628 2932 1629
rect 3062 1633 3068 1634
rect 3062 1629 3063 1633
rect 3067 1629 3068 1633
rect 3062 1628 3068 1629
rect 2830 1623 2836 1624
rect 2830 1619 2831 1623
rect 2835 1619 2836 1623
rect 2830 1618 2836 1619
rect 2910 1623 2916 1624
rect 2910 1619 2911 1623
rect 2915 1619 2916 1623
rect 2910 1618 2916 1619
rect 2647 1606 2651 1607
rect 2647 1601 2651 1602
rect 2655 1606 2659 1607
rect 2655 1601 2659 1602
rect 2767 1606 2771 1607
rect 2767 1601 2771 1602
rect 2791 1606 2795 1607
rect 2791 1601 2795 1602
rect 2614 1599 2620 1600
rect 2614 1595 2615 1599
rect 2619 1595 2620 1599
rect 2614 1594 2620 1595
rect 2648 1592 2650 1601
rect 2768 1592 2770 1601
rect 2166 1591 2172 1592
rect 2166 1587 2167 1591
rect 2171 1587 2172 1591
rect 2166 1586 2172 1587
rect 2286 1591 2292 1592
rect 2286 1587 2287 1591
rect 2291 1587 2292 1591
rect 2286 1586 2292 1587
rect 2406 1591 2412 1592
rect 2406 1587 2407 1591
rect 2411 1587 2412 1591
rect 2406 1586 2412 1587
rect 2526 1591 2532 1592
rect 2526 1587 2527 1591
rect 2531 1587 2532 1591
rect 2526 1586 2532 1587
rect 2646 1591 2652 1592
rect 2646 1587 2647 1591
rect 2651 1587 2652 1591
rect 2646 1586 2652 1587
rect 2766 1591 2772 1592
rect 2766 1587 2767 1591
rect 2771 1587 2772 1591
rect 2766 1586 2772 1587
rect 2832 1584 2834 1618
rect 2928 1607 2930 1628
rect 3064 1607 3066 1628
rect 3136 1624 3138 1738
rect 3992 1737 3994 1765
rect 3990 1736 3996 1737
rect 3990 1732 3991 1736
rect 3995 1732 3996 1736
rect 3990 1731 3996 1732
rect 3990 1719 3996 1720
rect 3990 1715 3991 1719
rect 3995 1715 3996 1719
rect 3318 1714 3324 1715
rect 3318 1710 3319 1714
rect 3323 1710 3324 1714
rect 3318 1709 3324 1710
rect 3510 1714 3516 1715
rect 3510 1710 3511 1714
rect 3515 1710 3516 1714
rect 3510 1709 3516 1710
rect 3702 1714 3708 1715
rect 3702 1710 3703 1714
rect 3707 1710 3708 1714
rect 3702 1709 3708 1710
rect 3894 1714 3900 1715
rect 3990 1714 3996 1715
rect 3894 1710 3895 1714
rect 3899 1710 3900 1714
rect 3894 1709 3900 1710
rect 3320 1691 3322 1709
rect 3512 1691 3514 1709
rect 3704 1691 3706 1709
rect 3896 1691 3898 1709
rect 3992 1691 3994 1714
rect 3207 1690 3211 1691
rect 3207 1685 3211 1686
rect 3319 1690 3323 1691
rect 3319 1685 3323 1686
rect 3351 1690 3355 1691
rect 3351 1685 3355 1686
rect 3511 1690 3515 1691
rect 3511 1685 3515 1686
rect 3703 1690 3707 1691
rect 3703 1685 3707 1686
rect 3895 1690 3899 1691
rect 3895 1685 3899 1686
rect 3991 1690 3995 1691
rect 3991 1685 3995 1686
rect 3208 1675 3210 1685
rect 3352 1675 3354 1685
rect 3206 1674 3212 1675
rect 3206 1670 3207 1674
rect 3211 1670 3212 1674
rect 3206 1669 3212 1670
rect 3350 1674 3356 1675
rect 3350 1670 3351 1674
rect 3355 1670 3356 1674
rect 3992 1670 3994 1685
rect 3350 1669 3356 1670
rect 3990 1669 3996 1670
rect 3990 1665 3991 1669
rect 3995 1665 3996 1669
rect 3990 1664 3996 1665
rect 3990 1652 3996 1653
rect 3990 1648 3991 1652
rect 3995 1648 3996 1652
rect 3990 1647 3996 1648
rect 3190 1643 3196 1644
rect 3190 1639 3191 1643
rect 3195 1639 3196 1643
rect 3190 1638 3196 1639
rect 3192 1624 3194 1638
rect 3206 1633 3212 1634
rect 3206 1629 3207 1633
rect 3211 1629 3212 1633
rect 3206 1628 3212 1629
rect 3350 1633 3356 1634
rect 3350 1629 3351 1633
rect 3355 1629 3356 1633
rect 3350 1628 3356 1629
rect 3134 1623 3140 1624
rect 3134 1619 3135 1623
rect 3139 1619 3140 1623
rect 3134 1618 3140 1619
rect 3190 1623 3196 1624
rect 3190 1619 3191 1623
rect 3195 1619 3196 1623
rect 3190 1618 3196 1619
rect 3208 1607 3210 1628
rect 3330 1623 3336 1624
rect 3330 1619 3331 1623
rect 3335 1619 3336 1623
rect 3330 1618 3336 1619
rect 2887 1606 2891 1607
rect 2887 1601 2891 1602
rect 2927 1606 2931 1607
rect 2927 1601 2931 1602
rect 3007 1606 3011 1607
rect 3007 1601 3011 1602
rect 3063 1606 3067 1607
rect 3063 1601 3067 1602
rect 3127 1606 3131 1607
rect 3127 1601 3131 1602
rect 3207 1606 3211 1607
rect 3207 1601 3211 1602
rect 3255 1606 3259 1607
rect 3255 1601 3259 1602
rect 2888 1592 2890 1601
rect 2918 1599 2924 1600
rect 2918 1595 2919 1599
rect 2923 1595 2924 1599
rect 2918 1594 2924 1595
rect 2886 1591 2892 1592
rect 2886 1587 2887 1591
rect 2891 1587 2892 1591
rect 2886 1586 2892 1587
rect 2746 1583 2752 1584
rect 2534 1579 2540 1580
rect 2534 1575 2535 1579
rect 2539 1575 2540 1579
rect 2746 1579 2747 1583
rect 2751 1579 2752 1583
rect 2746 1578 2752 1579
rect 2830 1583 2836 1584
rect 2830 1579 2831 1583
rect 2835 1579 2836 1583
rect 2830 1578 2836 1579
rect 2534 1574 2540 1575
rect 2070 1572 2076 1573
rect 2030 1571 2036 1572
rect 2030 1567 2031 1571
rect 2035 1567 2036 1571
rect 2070 1568 2071 1572
rect 2075 1568 2076 1572
rect 2070 1567 2076 1568
rect 1606 1566 1612 1567
rect 1606 1562 1607 1566
rect 1611 1562 1612 1566
rect 1606 1561 1612 1562
rect 1766 1566 1772 1567
rect 1766 1562 1767 1566
rect 1771 1562 1772 1566
rect 1766 1561 1772 1562
rect 1934 1566 1940 1567
rect 2030 1566 2036 1567
rect 1934 1562 1935 1566
rect 1939 1562 1940 1566
rect 1934 1561 1940 1562
rect 1608 1543 1610 1561
rect 1768 1543 1770 1561
rect 1936 1543 1938 1561
rect 2032 1543 2034 1566
rect 2070 1555 2076 1556
rect 2070 1551 2071 1555
rect 2075 1551 2076 1555
rect 2070 1550 2076 1551
rect 2166 1550 2172 1551
rect 1559 1542 1563 1543
rect 1559 1537 1563 1538
rect 1607 1542 1611 1543
rect 1607 1537 1611 1538
rect 1767 1542 1771 1543
rect 1767 1537 1771 1538
rect 1935 1542 1939 1543
rect 1935 1537 1939 1538
rect 2031 1542 2035 1543
rect 2031 1537 2035 1538
rect 1560 1527 1562 1537
rect 1558 1526 1564 1527
rect 1558 1522 1559 1526
rect 1563 1522 1564 1526
rect 2032 1522 2034 1537
rect 2072 1527 2074 1550
rect 2166 1546 2167 1550
rect 2171 1546 2172 1550
rect 2166 1545 2172 1546
rect 2286 1550 2292 1551
rect 2286 1546 2287 1550
rect 2291 1546 2292 1550
rect 2286 1545 2292 1546
rect 2406 1550 2412 1551
rect 2406 1546 2407 1550
rect 2411 1546 2412 1550
rect 2406 1545 2412 1546
rect 2526 1550 2532 1551
rect 2526 1546 2527 1550
rect 2531 1546 2532 1550
rect 2526 1545 2532 1546
rect 2168 1527 2170 1545
rect 2288 1527 2290 1545
rect 2408 1527 2410 1545
rect 2528 1527 2530 1545
rect 2071 1526 2075 1527
rect 1558 1521 1564 1522
rect 2030 1521 2036 1522
rect 2071 1521 2075 1522
rect 2167 1526 2171 1527
rect 2167 1521 2171 1522
rect 2287 1526 2291 1527
rect 2287 1521 2291 1522
rect 2351 1526 2355 1527
rect 2351 1521 2355 1522
rect 2407 1526 2411 1527
rect 2407 1521 2411 1522
rect 2463 1526 2467 1527
rect 2463 1521 2467 1522
rect 2527 1526 2531 1527
rect 2527 1521 2531 1522
rect 2030 1517 2031 1521
rect 2035 1517 2036 1521
rect 2030 1516 2036 1517
rect 2072 1506 2074 1521
rect 2352 1511 2354 1521
rect 2464 1511 2466 1521
rect 2350 1510 2356 1511
rect 2350 1506 2351 1510
rect 2355 1506 2356 1510
rect 2070 1505 2076 1506
rect 2350 1505 2356 1506
rect 2462 1510 2468 1511
rect 2462 1506 2463 1510
rect 2467 1506 2468 1510
rect 2462 1505 2468 1506
rect 2030 1504 2036 1505
rect 2030 1500 2031 1504
rect 2035 1500 2036 1504
rect 2070 1501 2071 1505
rect 2075 1501 2076 1505
rect 2070 1500 2076 1501
rect 2030 1499 2036 1500
rect 598 1495 604 1496
rect 598 1491 599 1495
rect 603 1491 604 1495
rect 598 1490 604 1491
rect 718 1495 724 1496
rect 718 1491 719 1495
rect 723 1491 724 1495
rect 718 1490 724 1491
rect 758 1495 764 1496
rect 758 1491 759 1495
rect 763 1491 764 1495
rect 758 1490 764 1491
rect 950 1495 956 1496
rect 950 1491 951 1495
rect 955 1491 956 1495
rect 950 1490 956 1491
rect 990 1495 996 1496
rect 990 1491 991 1495
rect 995 1491 996 1495
rect 990 1490 996 1491
rect 1182 1495 1188 1496
rect 1182 1491 1183 1495
rect 1187 1491 1188 1495
rect 1182 1490 1188 1491
rect 1422 1495 1428 1496
rect 1422 1491 1423 1495
rect 1427 1491 1428 1495
rect 1422 1490 1428 1491
rect 1542 1495 1548 1496
rect 1542 1491 1543 1495
rect 1547 1491 1548 1495
rect 1542 1490 1548 1491
rect 1550 1495 1556 1496
rect 1550 1491 1551 1495
rect 1555 1491 1556 1495
rect 1550 1490 1556 1491
rect 600 1476 602 1490
rect 614 1485 620 1486
rect 614 1481 615 1485
rect 619 1481 620 1485
rect 614 1480 620 1481
rect 558 1475 564 1476
rect 558 1471 559 1475
rect 563 1471 564 1475
rect 558 1470 564 1471
rect 598 1475 604 1476
rect 598 1471 599 1475
rect 603 1471 604 1475
rect 598 1470 604 1471
rect 616 1459 618 1480
rect 720 1476 722 1490
rect 734 1485 740 1486
rect 734 1481 735 1485
rect 739 1481 740 1485
rect 734 1480 740 1481
rect 718 1475 724 1476
rect 718 1471 719 1475
rect 723 1471 724 1475
rect 718 1470 724 1471
rect 670 1459 676 1460
rect 736 1459 738 1480
rect 111 1458 115 1459
rect 111 1453 115 1454
rect 503 1458 507 1459
rect 503 1453 507 1454
rect 583 1458 587 1459
rect 583 1453 587 1454
rect 615 1458 619 1459
rect 670 1455 671 1459
rect 675 1455 676 1459
rect 670 1454 676 1455
rect 687 1458 691 1459
rect 615 1453 619 1454
rect 112 1425 114 1453
rect 584 1444 586 1453
rect 582 1443 588 1444
rect 582 1439 583 1443
rect 587 1439 588 1443
rect 582 1438 588 1439
rect 672 1436 674 1454
rect 687 1453 691 1454
rect 735 1458 739 1459
rect 735 1453 739 1454
rect 688 1444 690 1453
rect 760 1452 762 1490
rect 854 1485 860 1486
rect 854 1481 855 1485
rect 859 1481 860 1485
rect 854 1480 860 1481
rect 856 1459 858 1480
rect 952 1476 954 1490
rect 966 1485 972 1486
rect 966 1481 967 1485
rect 971 1481 972 1485
rect 966 1480 972 1481
rect 1078 1485 1084 1486
rect 1078 1481 1079 1485
rect 1083 1481 1084 1485
rect 1078 1480 1084 1481
rect 918 1475 924 1476
rect 918 1471 919 1475
rect 923 1471 924 1475
rect 918 1470 924 1471
rect 950 1475 956 1476
rect 950 1471 951 1475
rect 955 1471 956 1475
rect 950 1470 956 1471
rect 791 1458 795 1459
rect 791 1453 795 1454
rect 855 1458 859 1459
rect 855 1453 859 1454
rect 895 1458 899 1459
rect 895 1453 899 1454
rect 758 1451 764 1452
rect 758 1447 759 1451
rect 763 1447 764 1451
rect 758 1446 764 1447
rect 792 1444 794 1453
rect 896 1444 898 1453
rect 686 1443 692 1444
rect 686 1439 687 1443
rect 691 1439 692 1443
rect 686 1438 692 1439
rect 790 1443 796 1444
rect 790 1439 791 1443
rect 795 1439 796 1443
rect 790 1438 796 1439
rect 894 1443 900 1444
rect 894 1439 895 1443
rect 899 1439 900 1443
rect 894 1438 900 1439
rect 670 1435 676 1436
rect 670 1431 671 1435
rect 675 1431 676 1435
rect 670 1430 676 1431
rect 854 1435 860 1436
rect 854 1431 855 1435
rect 859 1431 860 1435
rect 920 1432 922 1470
rect 968 1459 970 1480
rect 1080 1459 1082 1480
rect 1184 1468 1186 1490
rect 1198 1485 1204 1486
rect 1198 1481 1199 1485
rect 1203 1481 1204 1485
rect 1198 1480 1204 1481
rect 1318 1485 1324 1486
rect 1318 1481 1319 1485
rect 1323 1481 1324 1485
rect 1318 1480 1324 1481
rect 1182 1467 1188 1468
rect 1182 1463 1183 1467
rect 1187 1463 1188 1467
rect 1182 1462 1188 1463
rect 1200 1459 1202 1480
rect 1270 1475 1276 1476
rect 1270 1471 1271 1475
rect 1275 1471 1276 1475
rect 1270 1470 1276 1471
rect 967 1458 971 1459
rect 967 1453 971 1454
rect 999 1458 1003 1459
rect 999 1453 1003 1454
rect 1079 1458 1083 1459
rect 1079 1453 1083 1454
rect 1103 1458 1107 1459
rect 1103 1453 1107 1454
rect 1199 1458 1203 1459
rect 1199 1453 1203 1454
rect 1207 1458 1211 1459
rect 1207 1453 1211 1454
rect 1000 1444 1002 1453
rect 1104 1444 1106 1453
rect 1166 1451 1172 1452
rect 1166 1447 1167 1451
rect 1171 1447 1172 1451
rect 1166 1446 1172 1447
rect 998 1443 1004 1444
rect 998 1439 999 1443
rect 1003 1439 1004 1443
rect 998 1438 1004 1439
rect 1102 1443 1108 1444
rect 1102 1439 1103 1443
rect 1107 1439 1108 1443
rect 1102 1438 1108 1439
rect 854 1430 860 1431
rect 918 1431 924 1432
rect 110 1424 116 1425
rect 110 1420 111 1424
rect 115 1420 116 1424
rect 110 1419 116 1420
rect 110 1407 116 1408
rect 110 1403 111 1407
rect 115 1403 116 1407
rect 110 1402 116 1403
rect 582 1402 588 1403
rect 112 1379 114 1402
rect 582 1398 583 1402
rect 587 1398 588 1402
rect 582 1397 588 1398
rect 686 1402 692 1403
rect 686 1398 687 1402
rect 691 1398 692 1402
rect 686 1397 692 1398
rect 790 1402 796 1403
rect 790 1398 791 1402
rect 795 1398 796 1402
rect 790 1397 796 1398
rect 584 1379 586 1397
rect 688 1379 690 1397
rect 792 1379 794 1397
rect 111 1378 115 1379
rect 111 1373 115 1374
rect 551 1378 555 1379
rect 551 1373 555 1374
rect 583 1378 587 1379
rect 583 1373 587 1374
rect 655 1378 659 1379
rect 655 1373 659 1374
rect 687 1378 691 1379
rect 687 1373 691 1374
rect 759 1378 763 1379
rect 759 1373 763 1374
rect 791 1378 795 1379
rect 791 1373 795 1374
rect 112 1358 114 1373
rect 552 1363 554 1373
rect 656 1363 658 1373
rect 760 1363 762 1373
rect 550 1362 556 1363
rect 550 1358 551 1362
rect 555 1358 556 1362
rect 110 1357 116 1358
rect 550 1357 556 1358
rect 654 1362 660 1363
rect 654 1358 655 1362
rect 659 1358 660 1362
rect 654 1357 660 1358
rect 758 1362 764 1363
rect 758 1358 759 1362
rect 763 1358 764 1362
rect 758 1357 764 1358
rect 110 1353 111 1357
rect 115 1353 116 1357
rect 110 1352 116 1353
rect 110 1340 116 1341
rect 110 1336 111 1340
rect 115 1336 116 1340
rect 110 1335 116 1336
rect 112 1303 114 1335
rect 638 1331 644 1332
rect 638 1327 639 1331
rect 643 1327 644 1331
rect 638 1326 644 1327
rect 550 1321 556 1322
rect 550 1317 551 1321
rect 555 1317 556 1321
rect 550 1316 556 1317
rect 552 1303 554 1316
rect 640 1304 642 1326
rect 654 1321 660 1322
rect 654 1317 655 1321
rect 659 1317 660 1321
rect 654 1316 660 1317
rect 758 1321 764 1322
rect 758 1317 759 1321
rect 763 1317 764 1321
rect 758 1316 764 1317
rect 638 1303 644 1304
rect 656 1303 658 1316
rect 760 1303 762 1316
rect 856 1304 858 1430
rect 918 1427 919 1431
rect 923 1427 924 1431
rect 918 1426 924 1427
rect 894 1402 900 1403
rect 894 1398 895 1402
rect 899 1398 900 1402
rect 894 1397 900 1398
rect 998 1402 1004 1403
rect 998 1398 999 1402
rect 1003 1398 1004 1402
rect 998 1397 1004 1398
rect 1102 1402 1108 1403
rect 1102 1398 1103 1402
rect 1107 1398 1108 1402
rect 1102 1397 1108 1398
rect 896 1379 898 1397
rect 1000 1379 1002 1397
rect 1104 1379 1106 1397
rect 863 1378 867 1379
rect 863 1373 867 1374
rect 895 1378 899 1379
rect 895 1373 899 1374
rect 975 1378 979 1379
rect 975 1373 979 1374
rect 999 1378 1003 1379
rect 999 1373 1003 1374
rect 1087 1378 1091 1379
rect 1087 1373 1091 1374
rect 1103 1378 1107 1379
rect 1103 1373 1107 1374
rect 864 1363 866 1373
rect 976 1363 978 1373
rect 1088 1363 1090 1373
rect 862 1362 868 1363
rect 862 1358 863 1362
rect 867 1358 868 1362
rect 862 1357 868 1358
rect 974 1362 980 1363
rect 974 1358 975 1362
rect 979 1358 980 1362
rect 974 1357 980 1358
rect 1086 1362 1092 1363
rect 1086 1358 1087 1362
rect 1091 1358 1092 1362
rect 1086 1357 1092 1358
rect 1168 1332 1170 1446
rect 1208 1444 1210 1453
rect 1206 1443 1212 1444
rect 1206 1439 1207 1443
rect 1211 1439 1212 1443
rect 1206 1438 1212 1439
rect 1272 1436 1274 1470
rect 1320 1459 1322 1480
rect 1424 1476 1426 1490
rect 1438 1485 1444 1486
rect 1438 1481 1439 1485
rect 1443 1481 1444 1485
rect 1438 1480 1444 1481
rect 1422 1475 1428 1476
rect 1422 1471 1423 1475
rect 1427 1471 1428 1475
rect 1422 1470 1428 1471
rect 1406 1459 1412 1460
rect 1440 1459 1442 1480
rect 1544 1476 1546 1490
rect 1558 1485 1564 1486
rect 1558 1481 1559 1485
rect 1563 1481 1564 1485
rect 1558 1480 1564 1481
rect 1542 1475 1548 1476
rect 1542 1471 1543 1475
rect 1547 1471 1548 1475
rect 1542 1470 1548 1471
rect 1560 1459 1562 1480
rect 2032 1459 2034 1499
rect 2070 1488 2076 1489
rect 2070 1484 2071 1488
rect 2075 1484 2076 1488
rect 2070 1483 2076 1484
rect 1311 1458 1315 1459
rect 1311 1453 1315 1454
rect 1319 1458 1323 1459
rect 1406 1455 1407 1459
rect 1411 1455 1412 1459
rect 1406 1454 1412 1455
rect 1415 1458 1419 1459
rect 1319 1453 1323 1454
rect 1312 1444 1314 1453
rect 1310 1443 1316 1444
rect 1310 1439 1311 1443
rect 1315 1439 1316 1443
rect 1310 1438 1316 1439
rect 1270 1435 1276 1436
rect 1270 1431 1271 1435
rect 1275 1431 1276 1435
rect 1270 1430 1276 1431
rect 1206 1402 1212 1403
rect 1206 1398 1207 1402
rect 1211 1398 1212 1402
rect 1206 1397 1212 1398
rect 1310 1402 1316 1403
rect 1310 1398 1311 1402
rect 1315 1398 1316 1402
rect 1310 1397 1316 1398
rect 1208 1379 1210 1397
rect 1312 1379 1314 1397
rect 1199 1378 1203 1379
rect 1199 1373 1203 1374
rect 1207 1378 1211 1379
rect 1207 1373 1211 1374
rect 1311 1378 1315 1379
rect 1311 1373 1315 1374
rect 1200 1363 1202 1373
rect 1312 1363 1314 1373
rect 1198 1362 1204 1363
rect 1198 1358 1199 1362
rect 1203 1358 1204 1362
rect 1198 1357 1204 1358
rect 1310 1362 1316 1363
rect 1310 1358 1311 1362
rect 1315 1358 1316 1362
rect 1310 1357 1316 1358
rect 1408 1332 1410 1454
rect 1415 1453 1419 1454
rect 1439 1458 1443 1459
rect 1439 1453 1443 1454
rect 1519 1458 1523 1459
rect 1519 1453 1523 1454
rect 1559 1458 1563 1459
rect 1559 1453 1563 1454
rect 2031 1458 2035 1459
rect 2031 1453 2035 1454
rect 1416 1444 1418 1453
rect 1520 1444 1522 1453
rect 1414 1443 1420 1444
rect 1414 1439 1415 1443
rect 1419 1439 1420 1443
rect 1414 1438 1420 1439
rect 1518 1443 1524 1444
rect 1518 1439 1519 1443
rect 1523 1439 1524 1443
rect 1518 1438 1524 1439
rect 2032 1425 2034 1453
rect 2072 1443 2074 1483
rect 2446 1479 2452 1480
rect 2446 1475 2447 1479
rect 2451 1475 2452 1479
rect 2446 1474 2452 1475
rect 2350 1469 2356 1470
rect 2448 1469 2450 1474
rect 2462 1469 2468 1470
rect 2350 1465 2351 1469
rect 2355 1465 2356 1469
rect 2350 1464 2356 1465
rect 2447 1468 2451 1469
rect 2462 1465 2463 1469
rect 2467 1465 2468 1469
rect 2462 1464 2468 1465
rect 2352 1443 2354 1464
rect 2447 1463 2451 1464
rect 2464 1443 2466 1464
rect 2536 1460 2538 1574
rect 2646 1550 2652 1551
rect 2646 1546 2647 1550
rect 2651 1546 2652 1550
rect 2646 1545 2652 1546
rect 2648 1527 2650 1545
rect 2575 1526 2579 1527
rect 2575 1521 2579 1522
rect 2647 1526 2651 1527
rect 2647 1521 2651 1522
rect 2695 1526 2699 1527
rect 2695 1521 2699 1522
rect 2576 1511 2578 1521
rect 2696 1511 2698 1521
rect 2574 1510 2580 1511
rect 2574 1506 2575 1510
rect 2579 1506 2580 1510
rect 2574 1505 2580 1506
rect 2694 1510 2700 1511
rect 2694 1506 2695 1510
rect 2699 1506 2700 1510
rect 2694 1505 2700 1506
rect 2638 1475 2644 1476
rect 2638 1471 2639 1475
rect 2643 1471 2644 1475
rect 2638 1470 2644 1471
rect 2574 1469 2580 1470
rect 2574 1465 2575 1469
rect 2579 1465 2580 1469
rect 2574 1464 2580 1465
rect 2534 1459 2540 1460
rect 2534 1455 2535 1459
rect 2539 1455 2540 1459
rect 2534 1454 2540 1455
rect 2576 1443 2578 1464
rect 2071 1442 2075 1443
rect 2071 1437 2075 1438
rect 2343 1442 2347 1443
rect 2343 1437 2347 1438
rect 2351 1442 2355 1443
rect 2351 1437 2355 1438
rect 2447 1442 2451 1443
rect 2447 1437 2451 1438
rect 2463 1442 2467 1443
rect 2463 1437 2467 1438
rect 2567 1442 2571 1443
rect 2567 1437 2571 1438
rect 2575 1442 2579 1443
rect 2575 1437 2579 1438
rect 2030 1424 2036 1425
rect 2030 1420 2031 1424
rect 2035 1420 2036 1424
rect 2030 1419 2036 1420
rect 2072 1409 2074 1437
rect 2344 1428 2346 1437
rect 2448 1428 2450 1437
rect 2568 1428 2570 1437
rect 2640 1436 2642 1470
rect 2694 1469 2700 1470
rect 2694 1465 2695 1469
rect 2699 1465 2700 1469
rect 2694 1464 2700 1465
rect 2748 1464 2750 1578
rect 2766 1550 2772 1551
rect 2766 1546 2767 1550
rect 2771 1546 2772 1550
rect 2766 1545 2772 1546
rect 2886 1550 2892 1551
rect 2886 1546 2887 1550
rect 2891 1546 2892 1550
rect 2886 1545 2892 1546
rect 2768 1527 2770 1545
rect 2888 1527 2890 1545
rect 2767 1526 2771 1527
rect 2767 1521 2771 1522
rect 2815 1526 2819 1527
rect 2815 1521 2819 1522
rect 2887 1526 2891 1527
rect 2887 1521 2891 1522
rect 2816 1511 2818 1521
rect 2814 1510 2820 1511
rect 2814 1506 2815 1510
rect 2819 1506 2820 1510
rect 2814 1505 2820 1506
rect 2920 1480 2922 1594
rect 3008 1592 3010 1601
rect 3128 1592 3130 1601
rect 3256 1592 3258 1601
rect 3332 1600 3334 1618
rect 3352 1607 3354 1628
rect 3992 1607 3994 1647
rect 3351 1606 3355 1607
rect 3351 1601 3355 1602
rect 3991 1606 3995 1607
rect 3991 1601 3995 1602
rect 3330 1599 3336 1600
rect 3330 1595 3331 1599
rect 3335 1595 3336 1599
rect 3330 1594 3336 1595
rect 3006 1591 3012 1592
rect 3006 1587 3007 1591
rect 3011 1587 3012 1591
rect 3006 1586 3012 1587
rect 3126 1591 3132 1592
rect 3126 1587 3127 1591
rect 3131 1587 3132 1591
rect 3126 1586 3132 1587
rect 3254 1591 3260 1592
rect 3254 1587 3255 1591
rect 3259 1587 3260 1591
rect 3254 1586 3260 1587
rect 2990 1583 2996 1584
rect 2990 1579 2991 1583
rect 2995 1579 2996 1583
rect 2990 1578 2996 1579
rect 2927 1526 2931 1527
rect 2927 1521 2931 1522
rect 2928 1511 2930 1521
rect 2926 1510 2932 1511
rect 2926 1506 2927 1510
rect 2931 1506 2932 1510
rect 2926 1505 2932 1506
rect 2886 1479 2892 1480
rect 2886 1475 2887 1479
rect 2891 1475 2892 1479
rect 2886 1474 2892 1475
rect 2918 1479 2924 1480
rect 2918 1475 2919 1479
rect 2923 1475 2924 1479
rect 2918 1474 2924 1475
rect 2814 1469 2820 1470
rect 2767 1468 2771 1469
rect 2814 1465 2815 1469
rect 2819 1465 2820 1469
rect 2814 1464 2820 1465
rect 2696 1443 2698 1464
rect 2746 1463 2752 1464
rect 2767 1463 2771 1464
rect 2746 1459 2747 1463
rect 2751 1459 2752 1463
rect 2768 1460 2770 1463
rect 2746 1458 2752 1459
rect 2766 1459 2772 1460
rect 2766 1455 2767 1459
rect 2771 1455 2772 1459
rect 2766 1454 2772 1455
rect 2816 1443 2818 1464
rect 2695 1442 2699 1443
rect 2695 1437 2699 1438
rect 2815 1442 2819 1443
rect 2815 1437 2819 1438
rect 2839 1442 2843 1443
rect 2839 1437 2843 1438
rect 2638 1435 2644 1436
rect 2638 1431 2639 1435
rect 2643 1431 2644 1435
rect 2638 1430 2644 1431
rect 2696 1428 2698 1437
rect 2840 1428 2842 1437
rect 2888 1436 2890 1474
rect 2926 1469 2932 1470
rect 2926 1465 2927 1469
rect 2931 1465 2932 1469
rect 2992 1468 2994 1578
rect 3992 1573 3994 1601
rect 3990 1572 3996 1573
rect 3990 1568 3991 1572
rect 3995 1568 3996 1572
rect 3990 1567 3996 1568
rect 3990 1555 3996 1556
rect 3990 1551 3991 1555
rect 3995 1551 3996 1555
rect 3006 1550 3012 1551
rect 3006 1546 3007 1550
rect 3011 1546 3012 1550
rect 3006 1545 3012 1546
rect 3126 1550 3132 1551
rect 3126 1546 3127 1550
rect 3131 1546 3132 1550
rect 3126 1545 3132 1546
rect 3254 1550 3260 1551
rect 3990 1550 3996 1551
rect 3254 1546 3255 1550
rect 3259 1546 3260 1550
rect 3254 1545 3260 1546
rect 3008 1527 3010 1545
rect 3128 1527 3130 1545
rect 3256 1527 3258 1545
rect 3992 1527 3994 1550
rect 3007 1526 3011 1527
rect 3007 1521 3011 1522
rect 3047 1526 3051 1527
rect 3047 1521 3051 1522
rect 3127 1526 3131 1527
rect 3127 1521 3131 1522
rect 3167 1526 3171 1527
rect 3167 1521 3171 1522
rect 3255 1526 3259 1527
rect 3255 1521 3259 1522
rect 3287 1526 3291 1527
rect 3287 1521 3291 1522
rect 3407 1526 3411 1527
rect 3407 1521 3411 1522
rect 3991 1526 3995 1527
rect 3991 1521 3995 1522
rect 3048 1511 3050 1521
rect 3168 1511 3170 1521
rect 3288 1511 3290 1521
rect 3408 1511 3410 1521
rect 3046 1510 3052 1511
rect 3046 1506 3047 1510
rect 3051 1506 3052 1510
rect 3046 1505 3052 1506
rect 3166 1510 3172 1511
rect 3166 1506 3167 1510
rect 3171 1506 3172 1510
rect 3166 1505 3172 1506
rect 3286 1510 3292 1511
rect 3286 1506 3287 1510
rect 3291 1506 3292 1510
rect 3286 1505 3292 1506
rect 3406 1510 3412 1511
rect 3406 1506 3407 1510
rect 3411 1506 3412 1510
rect 3992 1506 3994 1521
rect 3406 1505 3412 1506
rect 3990 1505 3996 1506
rect 3990 1501 3991 1505
rect 3995 1501 3996 1505
rect 3990 1500 3996 1501
rect 3990 1488 3996 1489
rect 3990 1484 3991 1488
rect 3995 1484 3996 1488
rect 3990 1483 3996 1484
rect 3150 1479 3156 1480
rect 3150 1475 3151 1479
rect 3155 1475 3156 1479
rect 3150 1474 3156 1475
rect 3270 1479 3276 1480
rect 3270 1475 3271 1479
rect 3275 1475 3276 1479
rect 3270 1474 3276 1475
rect 3046 1469 3052 1470
rect 2926 1464 2932 1465
rect 2990 1467 2996 1468
rect 2928 1443 2930 1464
rect 2990 1463 2991 1467
rect 2995 1463 2996 1467
rect 3046 1465 3047 1469
rect 3051 1465 3052 1469
rect 3046 1464 3052 1465
rect 2990 1462 2996 1463
rect 2998 1459 3004 1460
rect 2998 1455 2999 1459
rect 3003 1455 3004 1459
rect 2998 1454 3004 1455
rect 2927 1442 2931 1443
rect 2927 1437 2931 1438
rect 2991 1442 2995 1443
rect 2991 1437 2995 1438
rect 2886 1435 2892 1436
rect 2886 1431 2887 1435
rect 2891 1431 2892 1435
rect 2886 1430 2892 1431
rect 2992 1428 2994 1437
rect 2342 1427 2348 1428
rect 2342 1423 2343 1427
rect 2347 1423 2348 1427
rect 2342 1422 2348 1423
rect 2446 1427 2452 1428
rect 2446 1423 2447 1427
rect 2451 1423 2452 1427
rect 2446 1422 2452 1423
rect 2566 1427 2572 1428
rect 2566 1423 2567 1427
rect 2571 1423 2572 1427
rect 2566 1422 2572 1423
rect 2694 1427 2700 1428
rect 2694 1423 2695 1427
rect 2699 1423 2700 1427
rect 2694 1422 2700 1423
rect 2838 1427 2844 1428
rect 2838 1423 2839 1427
rect 2843 1423 2844 1427
rect 2838 1422 2844 1423
rect 2990 1427 2996 1428
rect 2990 1423 2991 1427
rect 2995 1423 2996 1427
rect 2990 1422 2996 1423
rect 2766 1419 2772 1420
rect 2358 1415 2364 1416
rect 2358 1411 2359 1415
rect 2363 1411 2364 1415
rect 2766 1415 2767 1419
rect 2771 1415 2772 1419
rect 3000 1416 3002 1454
rect 3048 1443 3050 1464
rect 3152 1460 3154 1474
rect 3166 1469 3172 1470
rect 3166 1465 3167 1469
rect 3171 1465 3172 1469
rect 3166 1464 3172 1465
rect 3150 1459 3156 1460
rect 3150 1455 3151 1459
rect 3155 1455 3156 1459
rect 3150 1454 3156 1455
rect 3168 1443 3170 1464
rect 3272 1460 3274 1474
rect 3286 1469 3292 1470
rect 3286 1465 3287 1469
rect 3291 1465 3292 1469
rect 3286 1464 3292 1465
rect 3406 1469 3412 1470
rect 3406 1465 3407 1469
rect 3411 1465 3412 1469
rect 3406 1464 3412 1465
rect 3270 1459 3276 1460
rect 3270 1455 3271 1459
rect 3275 1455 3276 1459
rect 3270 1454 3276 1455
rect 3288 1443 3290 1464
rect 3378 1459 3384 1460
rect 3378 1455 3379 1459
rect 3383 1455 3384 1459
rect 3378 1454 3384 1455
rect 3047 1442 3051 1443
rect 3047 1437 3051 1438
rect 3143 1442 3147 1443
rect 3143 1437 3147 1438
rect 3167 1442 3171 1443
rect 3167 1437 3171 1438
rect 3287 1442 3291 1443
rect 3287 1437 3291 1438
rect 3303 1442 3307 1443
rect 3303 1437 3307 1438
rect 3144 1428 3146 1437
rect 3206 1435 3212 1436
rect 3206 1431 3207 1435
rect 3211 1431 3212 1435
rect 3206 1430 3212 1431
rect 3142 1427 3148 1428
rect 3142 1423 3143 1427
rect 3147 1423 3148 1427
rect 3142 1422 3148 1423
rect 2766 1414 2772 1415
rect 2998 1415 3004 1416
rect 2358 1410 2364 1411
rect 2070 1408 2076 1409
rect 2030 1407 2036 1408
rect 2030 1403 2031 1407
rect 2035 1403 2036 1407
rect 2070 1404 2071 1408
rect 2075 1404 2076 1408
rect 2070 1403 2076 1404
rect 1414 1402 1420 1403
rect 1414 1398 1415 1402
rect 1419 1398 1420 1402
rect 1414 1397 1420 1398
rect 1518 1402 1524 1403
rect 2030 1402 2036 1403
rect 1518 1398 1519 1402
rect 1523 1398 1524 1402
rect 1518 1397 1524 1398
rect 1416 1379 1418 1397
rect 1520 1379 1522 1397
rect 2032 1379 2034 1402
rect 2070 1391 2076 1392
rect 2070 1387 2071 1391
rect 2075 1387 2076 1391
rect 2070 1386 2076 1387
rect 2342 1386 2348 1387
rect 1415 1378 1419 1379
rect 1415 1373 1419 1374
rect 1431 1378 1435 1379
rect 1431 1373 1435 1374
rect 1519 1378 1523 1379
rect 1519 1373 1523 1374
rect 1551 1378 1555 1379
rect 1551 1373 1555 1374
rect 2031 1378 2035 1379
rect 2031 1373 2035 1374
rect 1432 1363 1434 1373
rect 1552 1363 1554 1373
rect 1430 1362 1436 1363
rect 1430 1358 1431 1362
rect 1435 1358 1436 1362
rect 1430 1357 1436 1358
rect 1550 1362 1556 1363
rect 1550 1358 1551 1362
rect 1555 1358 1556 1362
rect 2032 1358 2034 1373
rect 2072 1363 2074 1386
rect 2342 1382 2343 1386
rect 2347 1382 2348 1386
rect 2342 1381 2348 1382
rect 2344 1363 2346 1381
rect 2071 1362 2075 1363
rect 1550 1357 1556 1358
rect 2030 1357 2036 1358
rect 2071 1357 2075 1358
rect 2287 1362 2291 1363
rect 2287 1357 2291 1358
rect 2343 1362 2347 1363
rect 2343 1357 2347 1358
rect 2030 1353 2031 1357
rect 2035 1353 2036 1357
rect 2030 1352 2036 1353
rect 2072 1342 2074 1357
rect 2288 1347 2290 1357
rect 2286 1346 2292 1347
rect 2286 1342 2287 1346
rect 2291 1342 2292 1346
rect 2070 1341 2076 1342
rect 2286 1341 2292 1342
rect 2030 1340 2036 1341
rect 2030 1336 2031 1340
rect 2035 1336 2036 1340
rect 2070 1337 2071 1341
rect 2075 1337 2076 1341
rect 2070 1336 2076 1337
rect 2030 1335 2036 1336
rect 1166 1331 1172 1332
rect 1166 1327 1167 1331
rect 1171 1327 1172 1331
rect 1166 1326 1172 1327
rect 1406 1331 1412 1332
rect 1406 1327 1407 1331
rect 1411 1327 1412 1331
rect 1406 1326 1412 1327
rect 862 1321 868 1322
rect 862 1317 863 1321
rect 867 1317 868 1321
rect 862 1316 868 1317
rect 974 1321 980 1322
rect 974 1317 975 1321
rect 979 1317 980 1321
rect 974 1316 980 1317
rect 1086 1321 1092 1322
rect 1086 1317 1087 1321
rect 1091 1317 1092 1321
rect 1086 1316 1092 1317
rect 1198 1321 1204 1322
rect 1198 1317 1199 1321
rect 1203 1317 1204 1321
rect 1198 1316 1204 1317
rect 1310 1321 1316 1322
rect 1310 1317 1311 1321
rect 1315 1317 1316 1321
rect 1310 1316 1316 1317
rect 1430 1321 1436 1322
rect 1430 1317 1431 1321
rect 1435 1317 1436 1321
rect 1430 1316 1436 1317
rect 1550 1321 1556 1322
rect 1550 1317 1551 1321
rect 1555 1317 1556 1321
rect 1550 1316 1556 1317
rect 854 1303 860 1304
rect 864 1303 866 1316
rect 976 1303 978 1316
rect 1088 1303 1090 1316
rect 1200 1303 1202 1316
rect 1254 1311 1260 1312
rect 1254 1307 1255 1311
rect 1259 1307 1260 1311
rect 1254 1306 1260 1307
rect 111 1302 115 1303
rect 111 1297 115 1298
rect 343 1302 347 1303
rect 343 1297 347 1298
rect 463 1302 467 1303
rect 463 1297 467 1298
rect 551 1302 555 1303
rect 551 1297 555 1298
rect 599 1302 603 1303
rect 638 1299 639 1303
rect 643 1299 644 1303
rect 638 1298 644 1299
rect 655 1302 659 1303
rect 599 1297 603 1298
rect 655 1297 659 1298
rect 743 1302 747 1303
rect 743 1297 747 1298
rect 759 1302 763 1303
rect 854 1299 855 1303
rect 859 1299 860 1303
rect 854 1298 860 1299
rect 863 1302 867 1303
rect 759 1297 763 1298
rect 863 1297 867 1298
rect 903 1302 907 1303
rect 903 1297 907 1298
rect 975 1302 979 1303
rect 975 1297 979 1298
rect 1063 1302 1067 1303
rect 1063 1297 1067 1298
rect 1087 1302 1091 1303
rect 1087 1297 1091 1298
rect 1199 1302 1203 1303
rect 1199 1297 1203 1298
rect 1231 1302 1235 1303
rect 1231 1297 1235 1298
rect 112 1269 114 1297
rect 344 1288 346 1297
rect 464 1288 466 1297
rect 600 1288 602 1297
rect 744 1288 746 1297
rect 904 1288 906 1297
rect 1064 1288 1066 1297
rect 1126 1295 1132 1296
rect 1126 1291 1127 1295
rect 1131 1291 1132 1295
rect 1126 1290 1132 1291
rect 342 1287 348 1288
rect 342 1283 343 1287
rect 347 1283 348 1287
rect 342 1282 348 1283
rect 462 1287 468 1288
rect 462 1283 463 1287
rect 467 1283 468 1287
rect 462 1282 468 1283
rect 598 1287 604 1288
rect 598 1283 599 1287
rect 603 1283 604 1287
rect 598 1282 604 1283
rect 742 1287 748 1288
rect 742 1283 743 1287
rect 747 1283 748 1287
rect 742 1282 748 1283
rect 902 1287 908 1288
rect 902 1283 903 1287
rect 907 1283 908 1287
rect 902 1282 908 1283
rect 1062 1287 1068 1288
rect 1062 1283 1063 1287
rect 1067 1283 1068 1287
rect 1062 1282 1068 1283
rect 446 1279 452 1280
rect 446 1275 447 1279
rect 451 1275 452 1279
rect 446 1274 452 1275
rect 110 1268 116 1269
rect 110 1264 111 1268
rect 115 1264 116 1268
rect 110 1263 116 1264
rect 110 1251 116 1252
rect 110 1247 111 1251
rect 115 1247 116 1251
rect 110 1246 116 1247
rect 342 1246 348 1247
rect 112 1231 114 1246
rect 342 1242 343 1246
rect 347 1242 348 1246
rect 342 1241 348 1242
rect 344 1231 346 1241
rect 448 1232 450 1274
rect 462 1246 468 1247
rect 462 1242 463 1246
rect 467 1242 468 1246
rect 462 1241 468 1242
rect 598 1246 604 1247
rect 598 1242 599 1246
rect 603 1242 604 1246
rect 598 1241 604 1242
rect 742 1246 748 1247
rect 742 1242 743 1246
rect 747 1242 748 1246
rect 742 1241 748 1242
rect 902 1246 908 1247
rect 902 1242 903 1246
rect 907 1242 908 1246
rect 902 1241 908 1242
rect 1062 1246 1068 1247
rect 1062 1242 1063 1246
rect 1067 1242 1068 1246
rect 1062 1241 1068 1242
rect 446 1231 452 1232
rect 464 1231 466 1241
rect 600 1231 602 1241
rect 744 1231 746 1241
rect 904 1231 906 1241
rect 990 1231 996 1232
rect 1064 1231 1066 1241
rect 111 1230 115 1231
rect 111 1225 115 1226
rect 183 1230 187 1231
rect 183 1225 187 1226
rect 343 1230 347 1231
rect 343 1225 347 1226
rect 351 1230 355 1231
rect 446 1227 447 1231
rect 451 1227 452 1231
rect 446 1226 452 1227
rect 463 1230 467 1231
rect 351 1225 355 1226
rect 463 1225 467 1226
rect 535 1230 539 1231
rect 535 1225 539 1226
rect 599 1230 603 1231
rect 599 1225 603 1226
rect 727 1230 731 1231
rect 727 1225 731 1226
rect 743 1230 747 1231
rect 743 1225 747 1226
rect 903 1230 907 1231
rect 903 1225 907 1226
rect 919 1230 923 1231
rect 990 1227 991 1231
rect 995 1227 996 1231
rect 990 1226 996 1227
rect 1063 1230 1067 1231
rect 919 1225 923 1226
rect 112 1210 114 1225
rect 184 1215 186 1225
rect 352 1215 354 1225
rect 536 1215 538 1225
rect 728 1215 730 1225
rect 920 1215 922 1225
rect 182 1214 188 1215
rect 182 1210 183 1214
rect 187 1210 188 1214
rect 110 1209 116 1210
rect 182 1209 188 1210
rect 350 1214 356 1215
rect 350 1210 351 1214
rect 355 1210 356 1214
rect 350 1209 356 1210
rect 534 1214 540 1215
rect 534 1210 535 1214
rect 539 1210 540 1214
rect 534 1209 540 1210
rect 726 1214 732 1215
rect 726 1210 727 1214
rect 731 1210 732 1214
rect 726 1209 732 1210
rect 918 1214 924 1215
rect 918 1210 919 1214
rect 923 1210 924 1214
rect 918 1209 924 1210
rect 110 1205 111 1209
rect 115 1205 116 1209
rect 110 1204 116 1205
rect 110 1192 116 1193
rect 110 1188 111 1192
rect 115 1188 116 1192
rect 110 1187 116 1188
rect 112 1151 114 1187
rect 334 1183 340 1184
rect 334 1179 335 1183
rect 339 1179 340 1183
rect 334 1178 340 1179
rect 182 1173 188 1174
rect 182 1169 183 1173
rect 187 1169 188 1173
rect 182 1168 188 1169
rect 184 1151 186 1168
rect 336 1152 338 1178
rect 350 1173 356 1174
rect 350 1169 351 1173
rect 355 1169 356 1173
rect 350 1168 356 1169
rect 534 1173 540 1174
rect 534 1169 535 1173
rect 539 1169 540 1173
rect 534 1168 540 1169
rect 726 1173 732 1174
rect 726 1169 727 1173
rect 731 1169 732 1173
rect 726 1168 732 1169
rect 918 1173 924 1174
rect 918 1169 919 1173
rect 923 1169 924 1173
rect 918 1168 924 1169
rect 334 1151 340 1152
rect 352 1151 354 1168
rect 536 1151 538 1168
rect 728 1151 730 1168
rect 920 1151 922 1168
rect 992 1164 994 1226
rect 1063 1225 1067 1226
rect 1103 1230 1107 1231
rect 1103 1225 1107 1226
rect 1104 1215 1106 1225
rect 1102 1214 1108 1215
rect 1102 1210 1103 1214
rect 1107 1210 1108 1214
rect 1102 1209 1108 1210
rect 1128 1184 1130 1290
rect 1232 1288 1234 1297
rect 1230 1287 1236 1288
rect 1230 1283 1231 1287
rect 1235 1283 1236 1287
rect 1230 1282 1236 1283
rect 1256 1276 1258 1306
rect 1312 1303 1314 1316
rect 1432 1303 1434 1316
rect 1552 1303 1554 1316
rect 1606 1311 1612 1312
rect 1606 1307 1607 1311
rect 1611 1307 1612 1311
rect 1606 1306 1612 1307
rect 1311 1302 1315 1303
rect 1311 1297 1315 1298
rect 1407 1302 1411 1303
rect 1407 1297 1411 1298
rect 1431 1302 1435 1303
rect 1431 1297 1435 1298
rect 1551 1302 1555 1303
rect 1551 1297 1555 1298
rect 1583 1302 1587 1303
rect 1583 1297 1587 1298
rect 1408 1288 1410 1297
rect 1414 1295 1420 1296
rect 1414 1291 1415 1295
rect 1419 1291 1420 1295
rect 1414 1290 1420 1291
rect 1406 1287 1412 1288
rect 1406 1283 1407 1287
rect 1411 1283 1412 1287
rect 1406 1282 1412 1283
rect 1254 1275 1260 1276
rect 1254 1271 1255 1275
rect 1259 1271 1260 1275
rect 1254 1270 1260 1271
rect 1230 1246 1236 1247
rect 1230 1242 1231 1246
rect 1235 1242 1236 1246
rect 1230 1241 1236 1242
rect 1406 1246 1412 1247
rect 1406 1242 1407 1246
rect 1411 1242 1412 1246
rect 1406 1241 1412 1242
rect 1232 1231 1234 1241
rect 1408 1231 1410 1241
rect 1231 1230 1235 1231
rect 1231 1225 1235 1226
rect 1287 1230 1291 1231
rect 1287 1225 1291 1226
rect 1407 1230 1411 1231
rect 1407 1225 1411 1226
rect 1288 1215 1290 1225
rect 1286 1214 1292 1215
rect 1286 1210 1287 1214
rect 1291 1210 1292 1214
rect 1286 1209 1292 1210
rect 1416 1184 1418 1290
rect 1584 1288 1586 1297
rect 1582 1287 1588 1288
rect 1582 1283 1583 1287
rect 1587 1283 1588 1287
rect 1582 1282 1588 1283
rect 1608 1276 1610 1306
rect 2032 1303 2034 1335
rect 2070 1324 2076 1325
rect 2070 1320 2071 1324
rect 2075 1320 2076 1324
rect 2070 1319 2076 1320
rect 2031 1302 2035 1303
rect 2031 1297 2035 1298
rect 1606 1275 1612 1276
rect 1606 1271 1607 1275
rect 1611 1271 1612 1275
rect 1606 1270 1612 1271
rect 2032 1269 2034 1297
rect 2072 1283 2074 1319
rect 2286 1305 2292 1306
rect 2286 1301 2287 1305
rect 2291 1301 2292 1305
rect 2286 1300 2292 1301
rect 2288 1283 2290 1300
rect 2360 1296 2362 1410
rect 2446 1386 2452 1387
rect 2446 1382 2447 1386
rect 2451 1382 2452 1386
rect 2446 1381 2452 1382
rect 2566 1386 2572 1387
rect 2566 1382 2567 1386
rect 2571 1382 2572 1386
rect 2566 1381 2572 1382
rect 2694 1386 2700 1387
rect 2694 1382 2695 1386
rect 2699 1382 2700 1386
rect 2694 1381 2700 1382
rect 2448 1363 2450 1381
rect 2568 1363 2570 1381
rect 2696 1363 2698 1381
rect 2407 1362 2411 1363
rect 2407 1357 2411 1358
rect 2447 1362 2451 1363
rect 2447 1357 2451 1358
rect 2543 1362 2547 1363
rect 2543 1357 2547 1358
rect 2567 1362 2571 1363
rect 2567 1357 2571 1358
rect 2695 1362 2699 1363
rect 2695 1357 2699 1358
rect 2408 1347 2410 1357
rect 2544 1347 2546 1357
rect 2696 1347 2698 1357
rect 2406 1346 2412 1347
rect 2406 1342 2407 1346
rect 2411 1342 2412 1346
rect 2406 1341 2412 1342
rect 2542 1346 2548 1347
rect 2542 1342 2543 1346
rect 2547 1342 2548 1346
rect 2542 1341 2548 1342
rect 2694 1346 2700 1347
rect 2694 1342 2695 1346
rect 2699 1342 2700 1346
rect 2694 1341 2700 1342
rect 2390 1315 2396 1316
rect 2390 1311 2391 1315
rect 2395 1311 2396 1315
rect 2390 1310 2396 1311
rect 2526 1315 2532 1316
rect 2526 1311 2527 1315
rect 2531 1311 2532 1315
rect 2526 1310 2532 1311
rect 2392 1296 2394 1310
rect 2406 1305 2412 1306
rect 2406 1301 2407 1305
rect 2411 1301 2412 1305
rect 2406 1300 2412 1301
rect 2358 1295 2364 1296
rect 2358 1291 2359 1295
rect 2363 1291 2364 1295
rect 2358 1290 2364 1291
rect 2390 1295 2396 1296
rect 2390 1291 2391 1295
rect 2395 1291 2396 1295
rect 2390 1290 2396 1291
rect 2408 1283 2410 1300
rect 2528 1296 2530 1310
rect 2542 1305 2548 1306
rect 2542 1301 2543 1305
rect 2547 1301 2548 1305
rect 2542 1300 2548 1301
rect 2694 1305 2700 1306
rect 2694 1301 2695 1305
rect 2699 1301 2700 1305
rect 2694 1300 2700 1301
rect 2526 1295 2532 1296
rect 2526 1291 2527 1295
rect 2531 1291 2532 1295
rect 2526 1290 2532 1291
rect 2544 1283 2546 1300
rect 2696 1283 2698 1300
rect 2768 1296 2770 1414
rect 2998 1411 2999 1415
rect 3003 1411 3004 1415
rect 2998 1410 3004 1411
rect 2838 1386 2844 1387
rect 2838 1382 2839 1386
rect 2843 1382 2844 1386
rect 2838 1381 2844 1382
rect 2990 1386 2996 1387
rect 2990 1382 2991 1386
rect 2995 1382 2996 1386
rect 2990 1381 2996 1382
rect 3142 1386 3148 1387
rect 3142 1382 3143 1386
rect 3147 1382 3148 1386
rect 3142 1381 3148 1382
rect 2840 1363 2842 1381
rect 2992 1363 2994 1381
rect 3144 1363 3146 1381
rect 2839 1362 2843 1363
rect 2839 1357 2843 1358
rect 2855 1362 2859 1363
rect 2855 1357 2859 1358
rect 2991 1362 2995 1363
rect 2991 1357 2995 1358
rect 3015 1362 3019 1363
rect 3015 1357 3019 1358
rect 3143 1362 3147 1363
rect 3143 1357 3147 1358
rect 3183 1362 3187 1363
rect 3183 1357 3187 1358
rect 2856 1347 2858 1357
rect 3016 1347 3018 1357
rect 3184 1347 3186 1357
rect 2854 1346 2860 1347
rect 2854 1342 2855 1346
rect 2859 1342 2860 1346
rect 2854 1341 2860 1342
rect 3014 1346 3020 1347
rect 3014 1342 3015 1346
rect 3019 1342 3020 1346
rect 3014 1341 3020 1342
rect 3182 1346 3188 1347
rect 3182 1342 3183 1346
rect 3187 1342 3188 1346
rect 3182 1341 3188 1342
rect 3208 1316 3210 1430
rect 3304 1428 3306 1437
rect 3380 1436 3382 1454
rect 3408 1443 3410 1464
rect 3992 1443 3994 1483
rect 3407 1442 3411 1443
rect 3407 1437 3411 1438
rect 3471 1442 3475 1443
rect 3471 1437 3475 1438
rect 3647 1442 3651 1443
rect 3647 1437 3651 1438
rect 3823 1442 3827 1443
rect 3823 1437 3827 1438
rect 3991 1442 3995 1443
rect 3991 1437 3995 1438
rect 3378 1435 3384 1436
rect 3378 1431 3379 1435
rect 3383 1431 3384 1435
rect 3378 1430 3384 1431
rect 3472 1428 3474 1437
rect 3648 1428 3650 1437
rect 3814 1435 3820 1436
rect 3814 1431 3815 1435
rect 3819 1431 3820 1435
rect 3814 1430 3820 1431
rect 3302 1427 3308 1428
rect 3302 1423 3303 1427
rect 3307 1423 3308 1427
rect 3302 1422 3308 1423
rect 3470 1427 3476 1428
rect 3470 1423 3471 1427
rect 3475 1423 3476 1427
rect 3470 1422 3476 1423
rect 3646 1427 3652 1428
rect 3646 1423 3647 1427
rect 3651 1423 3652 1427
rect 3646 1422 3652 1423
rect 3730 1419 3736 1420
rect 3730 1415 3731 1419
rect 3735 1415 3736 1419
rect 3730 1414 3736 1415
rect 3302 1386 3308 1387
rect 3302 1382 3303 1386
rect 3307 1382 3308 1386
rect 3302 1381 3308 1382
rect 3470 1386 3476 1387
rect 3470 1382 3471 1386
rect 3475 1382 3476 1386
rect 3470 1381 3476 1382
rect 3646 1386 3652 1387
rect 3646 1382 3647 1386
rect 3651 1382 3652 1386
rect 3646 1381 3652 1382
rect 3304 1363 3306 1381
rect 3472 1363 3474 1381
rect 3648 1363 3650 1381
rect 3303 1362 3307 1363
rect 3303 1357 3307 1358
rect 3351 1362 3355 1363
rect 3351 1357 3355 1358
rect 3471 1362 3475 1363
rect 3471 1357 3475 1358
rect 3519 1362 3523 1363
rect 3519 1357 3523 1358
rect 3647 1362 3651 1363
rect 3647 1357 3651 1358
rect 3687 1362 3691 1363
rect 3687 1357 3691 1358
rect 3352 1347 3354 1357
rect 3520 1347 3522 1357
rect 3688 1347 3690 1357
rect 3350 1346 3356 1347
rect 3350 1342 3351 1346
rect 3355 1342 3356 1346
rect 3350 1341 3356 1342
rect 3518 1346 3524 1347
rect 3518 1342 3519 1346
rect 3523 1342 3524 1346
rect 3518 1341 3524 1342
rect 3686 1346 3692 1347
rect 3686 1342 3687 1346
rect 3691 1342 3692 1346
rect 3686 1341 3692 1342
rect 2838 1315 2844 1316
rect 2838 1311 2839 1315
rect 2843 1311 2844 1315
rect 2838 1310 2844 1311
rect 2926 1315 2932 1316
rect 2926 1311 2927 1315
rect 2931 1311 2932 1315
rect 2926 1310 2932 1311
rect 3166 1315 3172 1316
rect 3166 1311 3167 1315
rect 3171 1311 3172 1315
rect 3166 1310 3172 1311
rect 3206 1315 3212 1316
rect 3206 1311 3207 1315
rect 3211 1311 3212 1315
rect 3206 1310 3212 1311
rect 2840 1296 2842 1310
rect 2854 1305 2860 1306
rect 2854 1301 2855 1305
rect 2859 1301 2860 1305
rect 2854 1300 2860 1301
rect 2766 1295 2772 1296
rect 2766 1291 2767 1295
rect 2771 1291 2772 1295
rect 2766 1290 2772 1291
rect 2838 1295 2844 1296
rect 2838 1291 2839 1295
rect 2843 1291 2844 1295
rect 2838 1290 2844 1291
rect 2856 1283 2858 1300
rect 2071 1282 2075 1283
rect 2071 1277 2075 1278
rect 2127 1282 2131 1283
rect 2127 1277 2131 1278
rect 2287 1282 2291 1283
rect 2287 1277 2291 1278
rect 2295 1282 2299 1283
rect 2295 1277 2299 1278
rect 2407 1282 2411 1283
rect 2407 1277 2411 1278
rect 2479 1282 2483 1283
rect 2479 1277 2483 1278
rect 2543 1282 2547 1283
rect 2543 1277 2547 1278
rect 2679 1282 2683 1283
rect 2679 1277 2683 1278
rect 2695 1282 2699 1283
rect 2695 1277 2699 1278
rect 2855 1282 2859 1283
rect 2855 1277 2859 1278
rect 2879 1282 2883 1283
rect 2879 1277 2883 1278
rect 2030 1268 2036 1269
rect 2030 1264 2031 1268
rect 2035 1264 2036 1268
rect 2030 1263 2036 1264
rect 2030 1251 2036 1252
rect 2030 1247 2031 1251
rect 2035 1247 2036 1251
rect 2072 1249 2074 1277
rect 2128 1268 2130 1277
rect 2296 1268 2298 1277
rect 2480 1268 2482 1277
rect 2680 1268 2682 1277
rect 2880 1268 2882 1277
rect 2928 1276 2930 1310
rect 3014 1305 3020 1306
rect 3014 1301 3015 1305
rect 3019 1301 3020 1305
rect 3014 1300 3020 1301
rect 3016 1283 3018 1300
rect 3168 1296 3170 1310
rect 3182 1305 3188 1306
rect 3182 1301 3183 1305
rect 3187 1301 3188 1305
rect 3182 1300 3188 1301
rect 3350 1305 3356 1306
rect 3350 1301 3351 1305
rect 3355 1301 3356 1305
rect 3350 1300 3356 1301
rect 3518 1305 3524 1306
rect 3518 1301 3519 1305
rect 3523 1301 3524 1305
rect 3518 1300 3524 1301
rect 3686 1305 3692 1306
rect 3686 1301 3687 1305
rect 3691 1301 3692 1305
rect 3686 1300 3692 1301
rect 3086 1295 3092 1296
rect 3086 1291 3087 1295
rect 3091 1291 3092 1295
rect 3086 1290 3092 1291
rect 3166 1295 3172 1296
rect 3166 1291 3167 1295
rect 3171 1291 3172 1295
rect 3166 1290 3172 1291
rect 3015 1282 3019 1283
rect 3015 1277 3019 1278
rect 3071 1282 3075 1283
rect 3071 1277 3075 1278
rect 2926 1275 2932 1276
rect 2926 1271 2927 1275
rect 2931 1271 2932 1275
rect 2926 1270 2932 1271
rect 3006 1275 3012 1276
rect 3006 1271 3007 1275
rect 3011 1271 3012 1275
rect 3006 1270 3012 1271
rect 2126 1267 2132 1268
rect 2126 1263 2127 1267
rect 2131 1263 2132 1267
rect 2126 1262 2132 1263
rect 2294 1267 2300 1268
rect 2294 1263 2295 1267
rect 2299 1263 2300 1267
rect 2294 1262 2300 1263
rect 2478 1267 2484 1268
rect 2478 1263 2479 1267
rect 2483 1263 2484 1267
rect 2478 1262 2484 1263
rect 2678 1267 2684 1268
rect 2678 1263 2679 1267
rect 2683 1263 2684 1267
rect 2678 1262 2684 1263
rect 2878 1267 2884 1268
rect 2878 1263 2879 1267
rect 2883 1263 2884 1267
rect 2878 1262 2884 1263
rect 2150 1255 2156 1256
rect 2150 1251 2151 1255
rect 2155 1251 2156 1255
rect 2150 1250 2156 1251
rect 2870 1255 2876 1256
rect 2870 1251 2871 1255
rect 2875 1251 2876 1255
rect 2870 1250 2876 1251
rect 1582 1246 1588 1247
rect 2030 1246 2036 1247
rect 2070 1248 2076 1249
rect 1582 1242 1583 1246
rect 1587 1242 1588 1246
rect 1582 1241 1588 1242
rect 1584 1231 1586 1241
rect 2032 1231 2034 1246
rect 2070 1244 2071 1248
rect 2075 1244 2076 1248
rect 2070 1243 2076 1244
rect 2070 1231 2076 1232
rect 1471 1230 1475 1231
rect 1471 1225 1475 1226
rect 1583 1230 1587 1231
rect 1583 1225 1587 1226
rect 1655 1230 1659 1231
rect 1655 1225 1659 1226
rect 1839 1230 1843 1231
rect 1839 1225 1843 1226
rect 2031 1230 2035 1231
rect 2070 1227 2071 1231
rect 2075 1227 2076 1231
rect 2070 1226 2076 1227
rect 2126 1226 2132 1227
rect 2031 1225 2035 1226
rect 1472 1215 1474 1225
rect 1656 1215 1658 1225
rect 1840 1215 1842 1225
rect 1470 1214 1476 1215
rect 1470 1210 1471 1214
rect 1475 1210 1476 1214
rect 1470 1209 1476 1210
rect 1654 1214 1660 1215
rect 1654 1210 1655 1214
rect 1659 1210 1660 1214
rect 1654 1209 1660 1210
rect 1838 1214 1844 1215
rect 1838 1210 1839 1214
rect 1843 1210 1844 1214
rect 2032 1210 2034 1225
rect 1838 1209 1844 1210
rect 2030 1209 2036 1210
rect 2030 1205 2031 1209
rect 2035 1205 2036 1209
rect 2030 1204 2036 1205
rect 2072 1199 2074 1226
rect 2126 1222 2127 1226
rect 2131 1222 2132 1226
rect 2126 1221 2132 1222
rect 2128 1199 2130 1221
rect 2071 1198 2075 1199
rect 2071 1193 2075 1194
rect 2111 1198 2115 1199
rect 2111 1193 2115 1194
rect 2127 1198 2131 1199
rect 2127 1193 2131 1194
rect 2030 1192 2036 1193
rect 2030 1188 2031 1192
rect 2035 1188 2036 1192
rect 2030 1187 2036 1188
rect 1126 1183 1132 1184
rect 1126 1179 1127 1183
rect 1131 1179 1132 1183
rect 1126 1178 1132 1179
rect 1414 1183 1420 1184
rect 1414 1179 1415 1183
rect 1419 1179 1420 1183
rect 1414 1178 1420 1179
rect 1102 1173 1108 1174
rect 1102 1169 1103 1173
rect 1107 1169 1108 1173
rect 1102 1168 1108 1169
rect 1286 1173 1292 1174
rect 1286 1169 1287 1173
rect 1291 1169 1292 1173
rect 1286 1168 1292 1169
rect 1470 1173 1476 1174
rect 1470 1169 1471 1173
rect 1475 1169 1476 1173
rect 1470 1168 1476 1169
rect 1654 1173 1660 1174
rect 1654 1169 1655 1173
rect 1659 1169 1660 1173
rect 1654 1168 1660 1169
rect 1838 1173 1844 1174
rect 1838 1169 1839 1173
rect 1843 1169 1844 1173
rect 1838 1168 1844 1169
rect 990 1163 996 1164
rect 990 1159 991 1163
rect 995 1159 996 1163
rect 990 1158 996 1159
rect 1104 1151 1106 1168
rect 1186 1163 1192 1164
rect 1186 1159 1187 1163
rect 1191 1159 1192 1163
rect 1186 1158 1192 1159
rect 111 1150 115 1151
rect 111 1145 115 1146
rect 151 1150 155 1151
rect 151 1145 155 1146
rect 183 1150 187 1151
rect 183 1145 187 1146
rect 303 1150 307 1151
rect 334 1147 335 1151
rect 339 1147 340 1151
rect 334 1146 340 1147
rect 351 1150 355 1151
rect 303 1145 307 1146
rect 351 1145 355 1146
rect 495 1150 499 1151
rect 495 1145 499 1146
rect 535 1150 539 1151
rect 535 1145 539 1146
rect 703 1150 707 1151
rect 703 1145 707 1146
rect 727 1150 731 1151
rect 727 1145 731 1146
rect 911 1150 915 1151
rect 911 1145 915 1146
rect 919 1150 923 1151
rect 919 1145 923 1146
rect 1103 1150 1107 1151
rect 1103 1145 1107 1146
rect 1119 1150 1123 1151
rect 1119 1145 1123 1146
rect 112 1117 114 1145
rect 152 1136 154 1145
rect 304 1136 306 1145
rect 496 1136 498 1145
rect 704 1136 706 1145
rect 912 1136 914 1145
rect 1082 1143 1088 1144
rect 1082 1139 1083 1143
rect 1087 1139 1088 1143
rect 1082 1138 1088 1139
rect 150 1135 156 1136
rect 150 1131 151 1135
rect 155 1131 156 1135
rect 150 1130 156 1131
rect 302 1135 308 1136
rect 302 1131 303 1135
rect 307 1131 308 1135
rect 302 1130 308 1131
rect 494 1135 500 1136
rect 494 1131 495 1135
rect 499 1131 500 1135
rect 494 1130 500 1131
rect 702 1135 708 1136
rect 702 1131 703 1135
rect 707 1131 708 1135
rect 702 1130 708 1131
rect 910 1135 916 1136
rect 910 1131 911 1135
rect 915 1131 916 1135
rect 910 1130 916 1131
rect 110 1116 116 1117
rect 110 1112 111 1116
rect 115 1112 116 1116
rect 110 1111 116 1112
rect 110 1099 116 1100
rect 110 1095 111 1099
rect 115 1095 116 1099
rect 110 1094 116 1095
rect 150 1094 156 1095
rect 112 1071 114 1094
rect 150 1090 151 1094
rect 155 1090 156 1094
rect 150 1089 156 1090
rect 302 1094 308 1095
rect 302 1090 303 1094
rect 307 1090 308 1094
rect 302 1089 308 1090
rect 494 1094 500 1095
rect 494 1090 495 1094
rect 499 1090 500 1094
rect 494 1089 500 1090
rect 702 1094 708 1095
rect 702 1090 703 1094
rect 707 1090 708 1094
rect 702 1089 708 1090
rect 910 1094 916 1095
rect 910 1090 911 1094
rect 915 1090 916 1094
rect 910 1089 916 1090
rect 152 1071 154 1089
rect 304 1071 306 1089
rect 496 1071 498 1089
rect 704 1071 706 1089
rect 912 1071 914 1089
rect 111 1070 115 1071
rect 111 1065 115 1066
rect 151 1070 155 1071
rect 151 1065 155 1066
rect 279 1070 283 1071
rect 279 1065 283 1066
rect 303 1070 307 1071
rect 303 1065 307 1066
rect 447 1070 451 1071
rect 447 1065 451 1066
rect 495 1070 499 1071
rect 495 1065 499 1066
rect 623 1070 627 1071
rect 623 1065 627 1066
rect 703 1070 707 1071
rect 703 1065 707 1066
rect 799 1070 803 1071
rect 799 1065 803 1066
rect 911 1070 915 1071
rect 911 1065 915 1066
rect 967 1070 971 1071
rect 967 1065 971 1066
rect 112 1050 114 1065
rect 152 1055 154 1065
rect 280 1055 282 1065
rect 448 1055 450 1065
rect 624 1055 626 1065
rect 800 1055 802 1065
rect 968 1055 970 1065
rect 150 1054 156 1055
rect 150 1050 151 1054
rect 155 1050 156 1054
rect 110 1049 116 1050
rect 150 1049 156 1050
rect 278 1054 284 1055
rect 278 1050 279 1054
rect 283 1050 284 1054
rect 278 1049 284 1050
rect 446 1054 452 1055
rect 446 1050 447 1054
rect 451 1050 452 1054
rect 446 1049 452 1050
rect 622 1054 628 1055
rect 622 1050 623 1054
rect 627 1050 628 1054
rect 622 1049 628 1050
rect 798 1054 804 1055
rect 798 1050 799 1054
rect 803 1050 804 1054
rect 798 1049 804 1050
rect 966 1054 972 1055
rect 966 1050 967 1054
rect 971 1050 972 1054
rect 966 1049 972 1050
rect 110 1045 111 1049
rect 115 1045 116 1049
rect 110 1044 116 1045
rect 110 1032 116 1033
rect 110 1028 111 1032
rect 115 1028 116 1032
rect 110 1027 116 1028
rect 112 987 114 1027
rect 1084 1024 1086 1138
rect 1120 1136 1122 1145
rect 1118 1135 1124 1136
rect 1118 1131 1119 1135
rect 1123 1131 1124 1135
rect 1118 1130 1124 1131
rect 1188 1128 1190 1158
rect 1288 1151 1290 1168
rect 1472 1151 1474 1168
rect 1656 1151 1658 1168
rect 1840 1151 1842 1168
rect 1910 1163 1916 1164
rect 1910 1159 1911 1163
rect 1915 1159 1916 1163
rect 1910 1158 1916 1159
rect 1287 1150 1291 1151
rect 1287 1145 1291 1146
rect 1319 1150 1323 1151
rect 1319 1145 1323 1146
rect 1471 1150 1475 1151
rect 1471 1145 1475 1146
rect 1519 1150 1523 1151
rect 1519 1145 1523 1146
rect 1655 1150 1659 1151
rect 1655 1145 1659 1146
rect 1719 1150 1723 1151
rect 1719 1145 1723 1146
rect 1839 1150 1843 1151
rect 1839 1145 1843 1146
rect 1210 1143 1216 1144
rect 1210 1139 1211 1143
rect 1215 1139 1216 1143
rect 1210 1138 1216 1139
rect 1186 1127 1192 1128
rect 1186 1123 1187 1127
rect 1191 1123 1192 1127
rect 1186 1122 1192 1123
rect 1118 1094 1124 1095
rect 1118 1090 1119 1094
rect 1123 1090 1124 1094
rect 1118 1089 1124 1090
rect 1120 1071 1122 1089
rect 1119 1070 1123 1071
rect 1119 1065 1123 1066
rect 1127 1070 1131 1071
rect 1127 1065 1131 1066
rect 1128 1055 1130 1065
rect 1126 1054 1132 1055
rect 1126 1050 1127 1054
rect 1131 1050 1132 1054
rect 1126 1049 1132 1050
rect 1212 1024 1214 1138
rect 1320 1136 1322 1145
rect 1520 1136 1522 1145
rect 1720 1136 1722 1145
rect 1318 1135 1324 1136
rect 1318 1131 1319 1135
rect 1323 1131 1324 1135
rect 1318 1130 1324 1131
rect 1518 1135 1524 1136
rect 1518 1131 1519 1135
rect 1523 1131 1524 1135
rect 1518 1130 1524 1131
rect 1718 1135 1724 1136
rect 1718 1131 1719 1135
rect 1723 1131 1724 1135
rect 1718 1130 1724 1131
rect 1912 1128 1914 1158
rect 2032 1151 2034 1187
rect 2072 1178 2074 1193
rect 2112 1183 2114 1193
rect 2110 1182 2116 1183
rect 2110 1178 2111 1182
rect 2115 1178 2116 1182
rect 2070 1177 2076 1178
rect 2110 1177 2116 1178
rect 2070 1173 2071 1177
rect 2075 1173 2076 1177
rect 2070 1172 2076 1173
rect 2070 1160 2076 1161
rect 2070 1156 2071 1160
rect 2075 1156 2076 1160
rect 2070 1155 2076 1156
rect 1919 1150 1923 1151
rect 1919 1145 1923 1146
rect 2031 1150 2035 1151
rect 2031 1145 2035 1146
rect 1920 1136 1922 1145
rect 1918 1135 1924 1136
rect 1918 1131 1919 1135
rect 1923 1131 1924 1135
rect 1918 1130 1924 1131
rect 1910 1127 1916 1128
rect 1910 1123 1911 1127
rect 1915 1123 1916 1127
rect 1910 1122 1916 1123
rect 2032 1117 2034 1145
rect 2072 1123 2074 1155
rect 2110 1141 2116 1142
rect 2110 1137 2111 1141
rect 2115 1137 2116 1141
rect 2110 1136 2116 1137
rect 2152 1136 2154 1250
rect 2294 1226 2300 1227
rect 2294 1222 2295 1226
rect 2299 1222 2300 1226
rect 2294 1221 2300 1222
rect 2478 1226 2484 1227
rect 2478 1222 2479 1226
rect 2483 1222 2484 1226
rect 2478 1221 2484 1222
rect 2678 1226 2684 1227
rect 2678 1222 2679 1226
rect 2683 1222 2684 1226
rect 2678 1221 2684 1222
rect 2296 1199 2298 1221
rect 2480 1199 2482 1221
rect 2680 1199 2682 1221
rect 2247 1198 2251 1199
rect 2247 1193 2251 1194
rect 2295 1198 2299 1199
rect 2295 1193 2299 1194
rect 2407 1198 2411 1199
rect 2407 1193 2411 1194
rect 2479 1198 2483 1199
rect 2479 1193 2483 1194
rect 2559 1198 2563 1199
rect 2559 1193 2563 1194
rect 2679 1198 2683 1199
rect 2679 1193 2683 1194
rect 2703 1198 2707 1199
rect 2703 1193 2707 1194
rect 2863 1198 2867 1199
rect 2863 1193 2867 1194
rect 2248 1183 2250 1193
rect 2408 1183 2410 1193
rect 2560 1183 2562 1193
rect 2704 1183 2706 1193
rect 2864 1183 2866 1193
rect 2246 1182 2252 1183
rect 2246 1178 2247 1182
rect 2251 1178 2252 1182
rect 2246 1177 2252 1178
rect 2406 1182 2412 1183
rect 2406 1178 2407 1182
rect 2411 1178 2412 1182
rect 2406 1177 2412 1178
rect 2558 1182 2564 1183
rect 2558 1178 2559 1182
rect 2563 1178 2564 1182
rect 2558 1177 2564 1178
rect 2702 1182 2708 1183
rect 2702 1178 2703 1182
rect 2707 1178 2708 1182
rect 2702 1177 2708 1178
rect 2862 1182 2868 1183
rect 2862 1178 2863 1182
rect 2867 1178 2868 1182
rect 2862 1177 2868 1178
rect 2230 1151 2236 1152
rect 2230 1147 2231 1151
rect 2235 1147 2236 1151
rect 2230 1146 2236 1147
rect 2390 1151 2396 1152
rect 2390 1147 2391 1151
rect 2395 1147 2396 1151
rect 2390 1146 2396 1147
rect 2662 1151 2668 1152
rect 2662 1147 2663 1151
rect 2667 1147 2668 1151
rect 2662 1146 2668 1147
rect 2112 1123 2114 1136
rect 2150 1135 2156 1136
rect 2150 1131 2151 1135
rect 2155 1131 2156 1135
rect 2232 1132 2234 1146
rect 2246 1141 2252 1142
rect 2246 1137 2247 1141
rect 2251 1137 2252 1141
rect 2246 1136 2252 1137
rect 2150 1130 2156 1131
rect 2230 1131 2236 1132
rect 2230 1127 2231 1131
rect 2235 1127 2236 1131
rect 2230 1126 2236 1127
rect 2248 1123 2250 1136
rect 2392 1132 2394 1146
rect 2406 1141 2412 1142
rect 2406 1137 2407 1141
rect 2411 1137 2412 1141
rect 2406 1136 2412 1137
rect 2558 1141 2564 1142
rect 2558 1137 2559 1141
rect 2563 1137 2564 1141
rect 2558 1136 2564 1137
rect 2390 1131 2396 1132
rect 2390 1127 2391 1131
rect 2395 1127 2396 1131
rect 2390 1126 2396 1127
rect 2408 1123 2410 1136
rect 2560 1123 2562 1136
rect 2071 1122 2075 1123
rect 2071 1117 2075 1118
rect 2111 1122 2115 1123
rect 2111 1117 2115 1118
rect 2247 1122 2251 1123
rect 2247 1117 2251 1118
rect 2303 1122 2307 1123
rect 2303 1117 2307 1118
rect 2407 1122 2411 1123
rect 2407 1117 2411 1118
rect 2511 1122 2515 1123
rect 2511 1117 2515 1118
rect 2559 1122 2563 1123
rect 2559 1117 2563 1118
rect 2030 1116 2036 1117
rect 2030 1112 2031 1116
rect 2035 1112 2036 1116
rect 2030 1111 2036 1112
rect 2030 1099 2036 1100
rect 2030 1095 2031 1099
rect 2035 1095 2036 1099
rect 1318 1094 1324 1095
rect 1318 1090 1319 1094
rect 1323 1090 1324 1094
rect 1318 1089 1324 1090
rect 1518 1094 1524 1095
rect 1518 1090 1519 1094
rect 1523 1090 1524 1094
rect 1518 1089 1524 1090
rect 1718 1094 1724 1095
rect 1718 1090 1719 1094
rect 1723 1090 1724 1094
rect 1718 1089 1724 1090
rect 1918 1094 1924 1095
rect 2030 1094 2036 1095
rect 1918 1090 1919 1094
rect 1923 1090 1924 1094
rect 1918 1089 1924 1090
rect 1320 1071 1322 1089
rect 1520 1071 1522 1089
rect 1720 1071 1722 1089
rect 1920 1071 1922 1089
rect 2032 1071 2034 1094
rect 2072 1089 2074 1117
rect 2112 1108 2114 1117
rect 2304 1108 2306 1117
rect 2512 1108 2514 1117
rect 2664 1116 2666 1146
rect 2702 1141 2708 1142
rect 2702 1137 2703 1141
rect 2707 1137 2708 1141
rect 2702 1136 2708 1137
rect 2862 1141 2868 1142
rect 2862 1137 2863 1141
rect 2867 1137 2868 1141
rect 2862 1136 2868 1137
rect 2704 1123 2706 1136
rect 2864 1123 2866 1136
rect 2872 1132 2874 1250
rect 2878 1226 2884 1227
rect 2878 1222 2879 1226
rect 2883 1222 2884 1226
rect 2878 1221 2884 1222
rect 2880 1199 2882 1221
rect 2879 1198 2883 1199
rect 2879 1193 2883 1194
rect 3008 1152 3010 1270
rect 3072 1268 3074 1277
rect 3070 1267 3076 1268
rect 3070 1263 3071 1267
rect 3075 1263 3076 1267
rect 3070 1262 3076 1263
rect 3088 1256 3090 1290
rect 3184 1283 3186 1300
rect 3322 1295 3328 1296
rect 3322 1291 3323 1295
rect 3327 1291 3328 1295
rect 3322 1290 3328 1291
rect 3183 1282 3187 1283
rect 3183 1277 3187 1278
rect 3247 1282 3251 1283
rect 3247 1277 3251 1278
rect 3248 1268 3250 1277
rect 3324 1276 3326 1290
rect 3352 1283 3354 1300
rect 3520 1283 3522 1300
rect 3688 1283 3690 1300
rect 3732 1296 3734 1414
rect 3730 1295 3736 1296
rect 3730 1291 3731 1295
rect 3735 1291 3736 1295
rect 3730 1290 3736 1291
rect 3351 1282 3355 1283
rect 3351 1277 3355 1278
rect 3415 1282 3419 1283
rect 3415 1277 3419 1278
rect 3519 1282 3523 1283
rect 3519 1277 3523 1278
rect 3583 1282 3587 1283
rect 3583 1277 3587 1278
rect 3687 1282 3691 1283
rect 3687 1277 3691 1278
rect 3751 1282 3755 1283
rect 3751 1277 3755 1278
rect 3322 1275 3328 1276
rect 3322 1271 3323 1275
rect 3327 1271 3328 1275
rect 3322 1270 3328 1271
rect 3416 1268 3418 1277
rect 3584 1268 3586 1277
rect 3752 1268 3754 1277
rect 3246 1267 3252 1268
rect 3246 1263 3247 1267
rect 3251 1263 3252 1267
rect 3246 1262 3252 1263
rect 3414 1267 3420 1268
rect 3414 1263 3415 1267
rect 3419 1263 3420 1267
rect 3414 1262 3420 1263
rect 3582 1267 3588 1268
rect 3582 1263 3583 1267
rect 3587 1263 3588 1267
rect 3582 1262 3588 1263
rect 3750 1267 3756 1268
rect 3750 1263 3751 1267
rect 3755 1263 3756 1267
rect 3750 1262 3756 1263
rect 3816 1260 3818 1430
rect 3824 1428 3826 1437
rect 3822 1427 3828 1428
rect 3822 1423 3823 1427
rect 3827 1423 3828 1427
rect 3822 1422 3828 1423
rect 3918 1419 3924 1420
rect 3918 1415 3919 1419
rect 3923 1415 3924 1419
rect 3918 1414 3924 1415
rect 3822 1386 3828 1387
rect 3822 1382 3823 1386
rect 3827 1382 3828 1386
rect 3822 1381 3828 1382
rect 3824 1363 3826 1381
rect 3823 1362 3827 1363
rect 3823 1357 3827 1358
rect 3855 1362 3859 1363
rect 3855 1357 3859 1358
rect 3856 1347 3858 1357
rect 3854 1346 3860 1347
rect 3854 1342 3855 1346
rect 3859 1342 3860 1346
rect 3854 1341 3860 1342
rect 3854 1305 3860 1306
rect 3854 1301 3855 1305
rect 3859 1301 3860 1305
rect 3854 1300 3860 1301
rect 3856 1283 3858 1300
rect 3920 1296 3922 1414
rect 3992 1409 3994 1437
rect 3990 1408 3996 1409
rect 3990 1404 3991 1408
rect 3995 1404 3996 1408
rect 3990 1403 3996 1404
rect 3990 1391 3996 1392
rect 3990 1387 3991 1391
rect 3995 1387 3996 1391
rect 3990 1386 3996 1387
rect 3992 1363 3994 1386
rect 3991 1362 3995 1363
rect 3991 1357 3995 1358
rect 3992 1342 3994 1357
rect 3990 1341 3996 1342
rect 3990 1337 3991 1341
rect 3995 1337 3996 1341
rect 3990 1336 3996 1337
rect 3990 1324 3996 1325
rect 3990 1320 3991 1324
rect 3995 1320 3996 1324
rect 3990 1319 3996 1320
rect 3926 1315 3932 1316
rect 3926 1311 3927 1315
rect 3931 1311 3932 1315
rect 3926 1310 3932 1311
rect 3918 1295 3924 1296
rect 3918 1291 3919 1295
rect 3923 1291 3924 1295
rect 3918 1290 3924 1291
rect 3855 1282 3859 1283
rect 3855 1277 3859 1278
rect 3895 1282 3899 1283
rect 3895 1277 3899 1278
rect 3896 1268 3898 1277
rect 3928 1276 3930 1310
rect 3992 1283 3994 1319
rect 3991 1282 3995 1283
rect 3991 1277 3995 1278
rect 3926 1275 3932 1276
rect 3926 1271 3927 1275
rect 3931 1271 3932 1275
rect 3926 1270 3932 1271
rect 3894 1267 3900 1268
rect 3894 1263 3895 1267
rect 3899 1263 3900 1267
rect 3894 1262 3900 1263
rect 3814 1259 3820 1260
rect 3086 1255 3092 1256
rect 3086 1251 3087 1255
rect 3091 1251 3092 1255
rect 3814 1255 3815 1259
rect 3819 1255 3820 1259
rect 3814 1254 3820 1255
rect 3958 1259 3964 1260
rect 3958 1255 3959 1259
rect 3963 1255 3964 1259
rect 3958 1254 3964 1255
rect 3086 1250 3092 1251
rect 3070 1226 3076 1227
rect 3070 1222 3071 1226
rect 3075 1222 3076 1226
rect 3070 1221 3076 1222
rect 3246 1226 3252 1227
rect 3246 1222 3247 1226
rect 3251 1222 3252 1226
rect 3246 1221 3252 1222
rect 3414 1226 3420 1227
rect 3414 1222 3415 1226
rect 3419 1222 3420 1226
rect 3414 1221 3420 1222
rect 3582 1226 3588 1227
rect 3582 1222 3583 1226
rect 3587 1222 3588 1226
rect 3582 1221 3588 1222
rect 3750 1226 3756 1227
rect 3750 1222 3751 1226
rect 3755 1222 3756 1226
rect 3750 1221 3756 1222
rect 3894 1226 3900 1227
rect 3894 1222 3895 1226
rect 3899 1222 3900 1226
rect 3894 1221 3900 1222
rect 3072 1199 3074 1221
rect 3248 1199 3250 1221
rect 3416 1199 3418 1221
rect 3584 1199 3586 1221
rect 3752 1199 3754 1221
rect 3896 1199 3898 1221
rect 3039 1198 3043 1199
rect 3039 1193 3043 1194
rect 3071 1198 3075 1199
rect 3071 1193 3075 1194
rect 3239 1198 3243 1199
rect 3239 1193 3243 1194
rect 3247 1198 3251 1199
rect 3247 1193 3251 1194
rect 3415 1198 3419 1199
rect 3415 1193 3419 1194
rect 3455 1198 3459 1199
rect 3455 1193 3459 1194
rect 3583 1198 3587 1199
rect 3583 1193 3587 1194
rect 3687 1198 3691 1199
rect 3687 1193 3691 1194
rect 3751 1198 3755 1199
rect 3751 1193 3755 1194
rect 3895 1198 3899 1199
rect 3895 1193 3899 1194
rect 3040 1183 3042 1193
rect 3240 1183 3242 1193
rect 3456 1183 3458 1193
rect 3688 1183 3690 1193
rect 3896 1183 3898 1193
rect 3038 1182 3044 1183
rect 3038 1178 3039 1182
rect 3043 1178 3044 1182
rect 3038 1177 3044 1178
rect 3238 1182 3244 1183
rect 3238 1178 3239 1182
rect 3243 1178 3244 1182
rect 3238 1177 3244 1178
rect 3454 1182 3460 1183
rect 3454 1178 3455 1182
rect 3459 1178 3460 1182
rect 3454 1177 3460 1178
rect 3686 1182 3692 1183
rect 3686 1178 3687 1182
rect 3691 1178 3692 1182
rect 3686 1177 3692 1178
rect 3894 1182 3900 1183
rect 3894 1178 3895 1182
rect 3899 1178 3900 1182
rect 3894 1177 3900 1178
rect 3006 1151 3012 1152
rect 3006 1147 3007 1151
rect 3011 1147 3012 1151
rect 3006 1146 3012 1147
rect 3038 1141 3044 1142
rect 3038 1137 3039 1141
rect 3043 1137 3044 1141
rect 3038 1136 3044 1137
rect 3238 1141 3244 1142
rect 3238 1137 3239 1141
rect 3243 1137 3244 1141
rect 3238 1136 3244 1137
rect 3454 1141 3460 1142
rect 3454 1137 3455 1141
rect 3459 1137 3460 1141
rect 3454 1136 3460 1137
rect 3686 1141 3692 1142
rect 3686 1137 3687 1141
rect 3691 1137 3692 1141
rect 3686 1136 3692 1137
rect 3894 1141 3900 1142
rect 3894 1137 3895 1141
rect 3899 1137 3900 1141
rect 3894 1136 3900 1137
rect 2870 1131 2876 1132
rect 2870 1127 2871 1131
rect 2875 1127 2876 1131
rect 2870 1126 2876 1127
rect 3040 1123 3042 1136
rect 3070 1123 3076 1124
rect 3240 1123 3242 1136
rect 3456 1123 3458 1136
rect 3688 1123 3690 1136
rect 3896 1123 3898 1136
rect 3960 1132 3962 1254
rect 3992 1249 3994 1277
rect 3990 1248 3996 1249
rect 3990 1244 3991 1248
rect 3995 1244 3996 1248
rect 3990 1243 3996 1244
rect 3990 1231 3996 1232
rect 3990 1227 3991 1231
rect 3995 1227 3996 1231
rect 3990 1226 3996 1227
rect 3992 1199 3994 1226
rect 3991 1198 3995 1199
rect 3991 1193 3995 1194
rect 3992 1178 3994 1193
rect 3990 1177 3996 1178
rect 3990 1173 3991 1177
rect 3995 1173 3996 1177
rect 3990 1172 3996 1173
rect 3990 1160 3996 1161
rect 3990 1156 3991 1160
rect 3995 1156 3996 1160
rect 3990 1155 3996 1156
rect 3966 1151 3972 1152
rect 3966 1147 3967 1151
rect 3971 1147 3972 1151
rect 3966 1146 3972 1147
rect 3958 1131 3964 1132
rect 3958 1127 3959 1131
rect 3963 1127 3964 1131
rect 3958 1126 3964 1127
rect 2703 1122 2707 1123
rect 2703 1117 2707 1118
rect 2863 1122 2867 1123
rect 2863 1117 2867 1118
rect 2895 1122 2899 1123
rect 2895 1117 2899 1118
rect 3039 1122 3043 1123
rect 3070 1119 3071 1123
rect 3075 1119 3076 1123
rect 3070 1118 3076 1119
rect 3087 1122 3091 1123
rect 3039 1117 3043 1118
rect 2662 1115 2668 1116
rect 2662 1111 2663 1115
rect 2667 1111 2668 1115
rect 2662 1110 2668 1111
rect 2704 1108 2706 1117
rect 2896 1108 2898 1117
rect 2110 1107 2116 1108
rect 2110 1103 2111 1107
rect 2115 1103 2116 1107
rect 2110 1102 2116 1103
rect 2302 1107 2308 1108
rect 2302 1103 2303 1107
rect 2307 1103 2308 1107
rect 2302 1102 2308 1103
rect 2510 1107 2516 1108
rect 2510 1103 2511 1107
rect 2515 1103 2516 1107
rect 2510 1102 2516 1103
rect 2702 1107 2708 1108
rect 2702 1103 2703 1107
rect 2707 1103 2708 1107
rect 2702 1102 2708 1103
rect 2894 1107 2900 1108
rect 2894 1103 2895 1107
rect 2899 1103 2900 1107
rect 2894 1102 2900 1103
rect 3072 1100 3074 1118
rect 3087 1117 3091 1118
rect 3239 1122 3243 1123
rect 3239 1117 3243 1118
rect 3287 1122 3291 1123
rect 3287 1117 3291 1118
rect 3455 1122 3459 1123
rect 3455 1117 3459 1118
rect 3495 1122 3499 1123
rect 3495 1117 3499 1118
rect 3687 1122 3691 1123
rect 3687 1117 3691 1118
rect 3703 1122 3707 1123
rect 3703 1117 3707 1118
rect 3895 1122 3899 1123
rect 3895 1117 3899 1118
rect 3088 1108 3090 1117
rect 3288 1108 3290 1117
rect 3496 1108 3498 1117
rect 3704 1108 3706 1117
rect 3758 1115 3764 1116
rect 3758 1111 3759 1115
rect 3763 1111 3764 1115
rect 3758 1110 3764 1111
rect 3086 1107 3092 1108
rect 3086 1103 3087 1107
rect 3091 1103 3092 1107
rect 3086 1102 3092 1103
rect 3286 1107 3292 1108
rect 3286 1103 3287 1107
rect 3291 1103 3292 1107
rect 3286 1102 3292 1103
rect 3494 1107 3500 1108
rect 3494 1103 3495 1107
rect 3499 1103 3500 1107
rect 3494 1102 3500 1103
rect 3702 1107 3708 1108
rect 3702 1103 3703 1107
rect 3707 1103 3708 1107
rect 3702 1102 3708 1103
rect 2878 1099 2884 1100
rect 2102 1095 2108 1096
rect 2102 1091 2103 1095
rect 2107 1091 2108 1095
rect 2878 1095 2879 1099
rect 2883 1095 2884 1099
rect 2878 1094 2884 1095
rect 3070 1099 3076 1100
rect 3070 1095 3071 1099
rect 3075 1095 3076 1099
rect 3070 1094 3076 1095
rect 2102 1090 2108 1091
rect 2070 1088 2076 1089
rect 2070 1084 2071 1088
rect 2075 1084 2076 1088
rect 2070 1083 2076 1084
rect 2070 1071 2076 1072
rect 1279 1070 1283 1071
rect 1279 1065 1283 1066
rect 1319 1070 1323 1071
rect 1319 1065 1323 1066
rect 1423 1070 1427 1071
rect 1423 1065 1427 1066
rect 1519 1070 1523 1071
rect 1519 1065 1523 1066
rect 1559 1070 1563 1071
rect 1559 1065 1563 1066
rect 1695 1070 1699 1071
rect 1695 1065 1699 1066
rect 1719 1070 1723 1071
rect 1719 1065 1723 1066
rect 1823 1070 1827 1071
rect 1823 1065 1827 1066
rect 1919 1070 1923 1071
rect 1919 1065 1923 1066
rect 1935 1070 1939 1071
rect 1935 1065 1939 1066
rect 2031 1070 2035 1071
rect 2070 1067 2071 1071
rect 2075 1067 2076 1071
rect 2070 1066 2076 1067
rect 2031 1065 2035 1066
rect 1280 1055 1282 1065
rect 1424 1055 1426 1065
rect 1560 1055 1562 1065
rect 1696 1055 1698 1065
rect 1824 1055 1826 1065
rect 1936 1055 1938 1065
rect 1278 1054 1284 1055
rect 1278 1050 1279 1054
rect 1283 1050 1284 1054
rect 1278 1049 1284 1050
rect 1422 1054 1428 1055
rect 1422 1050 1423 1054
rect 1427 1050 1428 1054
rect 1422 1049 1428 1050
rect 1558 1054 1564 1055
rect 1558 1050 1559 1054
rect 1563 1050 1564 1054
rect 1558 1049 1564 1050
rect 1694 1054 1700 1055
rect 1694 1050 1695 1054
rect 1699 1050 1700 1054
rect 1694 1049 1700 1050
rect 1822 1054 1828 1055
rect 1822 1050 1823 1054
rect 1827 1050 1828 1054
rect 1822 1049 1828 1050
rect 1934 1054 1940 1055
rect 1934 1050 1935 1054
rect 1939 1050 1940 1054
rect 2032 1050 2034 1065
rect 1934 1049 1940 1050
rect 2030 1049 2036 1050
rect 2030 1045 2031 1049
rect 2035 1045 2036 1049
rect 2030 1044 2036 1045
rect 2072 1035 2074 1066
rect 2071 1034 2075 1035
rect 2030 1032 2036 1033
rect 2030 1028 2031 1032
rect 2035 1028 2036 1032
rect 2071 1029 2075 1030
rect 2030 1027 2036 1028
rect 222 1023 228 1024
rect 222 1019 223 1023
rect 227 1019 228 1023
rect 222 1018 228 1019
rect 1082 1023 1088 1024
rect 1082 1019 1083 1023
rect 1087 1019 1088 1023
rect 1082 1018 1088 1019
rect 1210 1023 1216 1024
rect 1210 1019 1211 1023
rect 1215 1019 1216 1023
rect 1210 1018 1216 1019
rect 1406 1023 1412 1024
rect 1406 1019 1407 1023
rect 1411 1019 1412 1023
rect 1406 1018 1412 1019
rect 150 1013 156 1014
rect 150 1009 151 1013
rect 155 1009 156 1013
rect 150 1008 156 1009
rect 152 987 154 1008
rect 111 986 115 987
rect 111 981 115 982
rect 151 986 155 987
rect 151 981 155 982
rect 112 953 114 981
rect 152 972 154 981
rect 224 980 226 1018
rect 278 1013 284 1014
rect 278 1009 279 1013
rect 283 1009 284 1013
rect 278 1008 284 1009
rect 446 1013 452 1014
rect 446 1009 447 1013
rect 451 1009 452 1013
rect 446 1008 452 1009
rect 622 1013 628 1014
rect 622 1009 623 1013
rect 627 1009 628 1013
rect 622 1008 628 1009
rect 798 1013 804 1014
rect 798 1009 799 1013
rect 803 1009 804 1013
rect 798 1008 804 1009
rect 966 1013 972 1014
rect 966 1009 967 1013
rect 971 1009 972 1013
rect 966 1008 972 1009
rect 1126 1013 1132 1014
rect 1126 1009 1127 1013
rect 1131 1009 1132 1013
rect 1126 1008 1132 1009
rect 1278 1013 1284 1014
rect 1278 1009 1279 1013
rect 1283 1009 1284 1013
rect 1278 1008 1284 1009
rect 280 987 282 1008
rect 448 987 450 1008
rect 624 987 626 1008
rect 800 987 802 1008
rect 968 987 970 1008
rect 1042 1003 1048 1004
rect 1042 999 1043 1003
rect 1047 999 1048 1003
rect 1042 998 1048 999
rect 279 986 283 987
rect 279 981 283 982
rect 287 986 291 987
rect 287 981 291 982
rect 447 986 451 987
rect 447 981 451 982
rect 471 986 475 987
rect 471 981 475 982
rect 623 986 627 987
rect 623 981 627 982
rect 671 986 675 987
rect 671 981 675 982
rect 799 986 803 987
rect 799 981 803 982
rect 871 986 875 987
rect 871 981 875 982
rect 967 986 971 987
rect 967 981 971 982
rect 222 979 228 980
rect 222 975 223 979
rect 227 975 228 979
rect 222 974 228 975
rect 288 972 290 981
rect 472 972 474 981
rect 655 972 659 973
rect 672 972 674 981
rect 872 972 874 981
rect 1044 980 1046 998
rect 1128 987 1130 1008
rect 1202 1003 1208 1004
rect 1202 999 1203 1003
rect 1207 999 1208 1003
rect 1202 998 1208 999
rect 1079 986 1083 987
rect 1079 981 1083 982
rect 1127 986 1131 987
rect 1127 981 1131 982
rect 1042 979 1048 980
rect 934 975 940 976
rect 150 971 156 972
rect 150 967 151 971
rect 155 967 156 971
rect 150 966 156 967
rect 286 971 292 972
rect 286 967 287 971
rect 291 967 292 971
rect 286 966 292 967
rect 470 971 476 972
rect 470 967 471 971
rect 475 967 476 971
rect 655 967 659 968
rect 670 971 676 972
rect 670 967 671 971
rect 675 967 676 971
rect 470 966 476 967
rect 656 964 658 967
rect 670 966 676 967
rect 870 971 876 972
rect 870 967 871 971
rect 875 967 876 971
rect 934 970 935 975
rect 939 970 940 975
rect 1042 975 1043 979
rect 1047 975 1048 979
rect 1042 974 1048 975
rect 1080 972 1082 981
rect 1204 980 1206 998
rect 1280 987 1282 1008
rect 1408 988 1410 1018
rect 1422 1013 1428 1014
rect 1422 1009 1423 1013
rect 1427 1009 1428 1013
rect 1422 1008 1428 1009
rect 1558 1013 1564 1014
rect 1558 1009 1559 1013
rect 1563 1009 1564 1013
rect 1558 1008 1564 1009
rect 1694 1013 1700 1014
rect 1694 1009 1695 1013
rect 1699 1009 1700 1013
rect 1694 1008 1700 1009
rect 1822 1013 1828 1014
rect 1822 1009 1823 1013
rect 1827 1009 1828 1013
rect 1822 1008 1828 1009
rect 1934 1013 1940 1014
rect 1934 1009 1935 1013
rect 1939 1009 1940 1013
rect 1934 1008 1940 1009
rect 1406 987 1412 988
rect 1424 987 1426 1008
rect 1560 987 1562 1008
rect 1696 987 1698 1008
rect 1824 987 1826 1008
rect 1936 987 1938 1008
rect 2032 987 2034 1027
rect 2072 1014 2074 1029
rect 2070 1013 2076 1014
rect 2070 1009 2071 1013
rect 2075 1009 2076 1013
rect 2070 1008 2076 1009
rect 2104 1004 2106 1090
rect 2110 1066 2116 1067
rect 2110 1062 2111 1066
rect 2115 1062 2116 1066
rect 2110 1061 2116 1062
rect 2302 1066 2308 1067
rect 2302 1062 2303 1066
rect 2307 1062 2308 1066
rect 2302 1061 2308 1062
rect 2510 1066 2516 1067
rect 2510 1062 2511 1066
rect 2515 1062 2516 1066
rect 2510 1061 2516 1062
rect 2702 1066 2708 1067
rect 2702 1062 2703 1066
rect 2707 1062 2708 1066
rect 2702 1061 2708 1062
rect 2112 1035 2114 1061
rect 2304 1035 2306 1061
rect 2512 1035 2514 1061
rect 2704 1035 2706 1061
rect 2111 1034 2115 1035
rect 2111 1029 2115 1030
rect 2303 1034 2307 1035
rect 2303 1029 2307 1030
rect 2319 1034 2323 1035
rect 2319 1029 2323 1030
rect 2487 1034 2491 1035
rect 2487 1029 2491 1030
rect 2511 1034 2515 1035
rect 2511 1029 2515 1030
rect 2663 1034 2667 1035
rect 2663 1029 2667 1030
rect 2703 1034 2707 1035
rect 2703 1029 2707 1030
rect 2847 1034 2851 1035
rect 2847 1029 2851 1030
rect 2320 1019 2322 1029
rect 2488 1019 2490 1029
rect 2664 1019 2666 1029
rect 2848 1019 2850 1029
rect 2318 1018 2324 1019
rect 2318 1014 2319 1018
rect 2323 1014 2324 1018
rect 2318 1013 2324 1014
rect 2486 1018 2492 1019
rect 2486 1014 2487 1018
rect 2491 1014 2492 1018
rect 2486 1013 2492 1014
rect 2662 1018 2668 1019
rect 2662 1014 2663 1018
rect 2667 1014 2668 1018
rect 2662 1013 2668 1014
rect 2846 1018 2852 1019
rect 2846 1014 2847 1018
rect 2851 1014 2852 1018
rect 2846 1013 2852 1014
rect 2102 1003 2108 1004
rect 2102 999 2103 1003
rect 2107 999 2108 1003
rect 2102 998 2108 999
rect 2070 996 2076 997
rect 2070 992 2071 996
rect 2075 992 2076 996
rect 2070 991 2076 992
rect 1279 986 1283 987
rect 1279 981 1283 982
rect 1287 986 1291 987
rect 1406 983 1407 987
rect 1411 983 1412 987
rect 1406 982 1412 983
rect 1423 986 1427 987
rect 1287 981 1291 982
rect 1423 981 1427 982
rect 1495 986 1499 987
rect 1495 981 1499 982
rect 1559 986 1563 987
rect 1559 981 1563 982
rect 1695 986 1699 987
rect 1695 981 1699 982
rect 1703 986 1707 987
rect 1703 981 1707 982
rect 1823 986 1827 987
rect 1823 981 1827 982
rect 1911 986 1915 987
rect 1911 981 1915 982
rect 1935 986 1939 987
rect 1935 981 1939 982
rect 2031 986 2035 987
rect 2031 981 2035 982
rect 1202 979 1208 980
rect 1202 975 1203 979
rect 1207 975 1208 979
rect 1202 974 1208 975
rect 1288 972 1290 981
rect 1496 972 1498 981
rect 1502 979 1508 980
rect 1502 975 1503 979
rect 1507 975 1508 979
rect 1502 974 1508 975
rect 998 971 1004 972
rect 935 967 939 968
rect 998 967 999 971
rect 1003 967 1004 971
rect 870 966 876 967
rect 998 966 1004 967
rect 1078 971 1084 972
rect 1078 967 1079 971
rect 1083 967 1084 971
rect 1078 966 1084 967
rect 1286 971 1292 972
rect 1286 967 1287 971
rect 1291 967 1292 971
rect 1286 966 1292 967
rect 1494 971 1500 972
rect 1494 967 1495 971
rect 1499 967 1500 971
rect 1494 966 1500 967
rect 654 963 660 964
rect 654 959 655 963
rect 659 959 660 963
rect 654 958 660 959
rect 662 959 668 960
rect 662 955 663 959
rect 667 955 668 959
rect 662 954 668 955
rect 110 952 116 953
rect 110 948 111 952
rect 115 948 116 952
rect 110 947 116 948
rect 110 935 116 936
rect 110 931 111 935
rect 115 931 116 935
rect 110 930 116 931
rect 150 930 156 931
rect 112 907 114 930
rect 150 926 151 930
rect 155 926 156 930
rect 150 925 156 926
rect 286 930 292 931
rect 286 926 287 930
rect 291 926 292 930
rect 286 925 292 926
rect 470 930 476 931
rect 470 926 471 930
rect 475 926 476 930
rect 470 925 476 926
rect 152 907 154 925
rect 288 907 290 925
rect 472 907 474 925
rect 111 906 115 907
rect 111 901 115 902
rect 151 906 155 907
rect 151 901 155 902
rect 287 906 291 907
rect 287 901 291 902
rect 319 906 323 907
rect 319 901 323 902
rect 471 906 475 907
rect 471 901 475 902
rect 519 906 523 907
rect 519 901 523 902
rect 112 886 114 901
rect 152 891 154 901
rect 320 891 322 901
rect 520 891 522 901
rect 150 890 156 891
rect 150 886 151 890
rect 155 886 156 890
rect 110 885 116 886
rect 150 885 156 886
rect 318 890 324 891
rect 318 886 319 890
rect 323 886 324 890
rect 318 885 324 886
rect 518 890 524 891
rect 518 886 519 890
rect 523 886 524 890
rect 518 885 524 886
rect 110 881 111 885
rect 115 881 116 885
rect 110 880 116 881
rect 110 868 116 869
rect 110 864 111 868
rect 115 864 116 868
rect 110 863 116 864
rect 112 823 114 863
rect 230 859 236 860
rect 230 855 231 859
rect 235 855 236 859
rect 230 854 236 855
rect 150 849 156 850
rect 150 845 151 849
rect 155 845 156 849
rect 150 844 156 845
rect 152 823 154 844
rect 232 832 234 854
rect 318 849 324 850
rect 318 845 319 849
rect 323 845 324 849
rect 318 844 324 845
rect 518 849 524 850
rect 518 845 519 849
rect 523 845 524 849
rect 518 844 524 845
rect 230 831 236 832
rect 230 827 231 831
rect 235 827 236 831
rect 230 826 236 827
rect 320 823 322 844
rect 520 823 522 844
rect 664 840 666 954
rect 670 930 676 931
rect 670 926 671 930
rect 675 926 676 930
rect 670 925 676 926
rect 870 930 876 931
rect 870 926 871 930
rect 875 926 876 930
rect 870 925 876 926
rect 672 907 674 925
rect 872 907 874 925
rect 671 906 675 907
rect 671 901 675 902
rect 727 906 731 907
rect 727 901 731 902
rect 871 906 875 907
rect 871 901 875 902
rect 935 906 939 907
rect 935 901 939 902
rect 728 891 730 901
rect 936 891 938 901
rect 726 890 732 891
rect 726 886 727 890
rect 731 886 732 890
rect 726 885 732 886
rect 934 890 940 891
rect 934 886 935 890
rect 939 886 940 890
rect 934 885 940 886
rect 750 859 756 860
rect 750 855 751 859
rect 755 855 756 859
rect 750 854 756 855
rect 726 849 732 850
rect 726 845 727 849
rect 731 845 732 849
rect 726 844 732 845
rect 662 839 668 840
rect 662 835 663 839
rect 667 835 668 839
rect 662 834 668 835
rect 728 823 730 844
rect 111 822 115 823
rect 111 817 115 818
rect 151 822 155 823
rect 151 817 155 818
rect 263 822 267 823
rect 263 817 267 818
rect 319 822 323 823
rect 319 817 323 818
rect 367 822 371 823
rect 367 817 371 818
rect 479 822 483 823
rect 479 817 483 818
rect 519 822 523 823
rect 519 817 523 818
rect 591 822 595 823
rect 591 817 595 818
rect 711 822 715 823
rect 711 817 715 818
rect 727 822 731 823
rect 727 817 731 818
rect 112 789 114 817
rect 264 808 266 817
rect 368 808 370 817
rect 480 808 482 817
rect 592 808 594 817
rect 712 808 714 817
rect 752 816 754 854
rect 934 849 940 850
rect 934 845 935 849
rect 939 845 940 849
rect 934 844 940 845
rect 936 823 938 844
rect 855 822 859 823
rect 855 817 859 818
rect 935 822 939 823
rect 935 817 939 818
rect 750 815 756 816
rect 750 811 751 815
rect 755 811 756 815
rect 750 810 756 811
rect 856 808 858 817
rect 262 807 268 808
rect 262 803 263 807
rect 267 803 268 807
rect 262 802 268 803
rect 366 807 372 808
rect 366 803 367 807
rect 371 803 372 807
rect 366 802 372 803
rect 478 807 484 808
rect 478 803 479 807
rect 483 803 484 807
rect 478 802 484 803
rect 590 807 596 808
rect 590 803 591 807
rect 595 803 596 807
rect 590 802 596 803
rect 710 807 716 808
rect 710 803 711 807
rect 715 803 716 807
rect 710 802 716 803
rect 854 807 860 808
rect 854 803 855 807
rect 859 803 860 807
rect 854 802 860 803
rect 1000 800 1002 966
rect 1078 930 1084 931
rect 1078 926 1079 930
rect 1083 926 1084 930
rect 1078 925 1084 926
rect 1286 930 1292 931
rect 1286 926 1287 930
rect 1291 926 1292 930
rect 1286 925 1292 926
rect 1494 930 1500 931
rect 1494 926 1495 930
rect 1499 926 1500 930
rect 1494 925 1500 926
rect 1080 907 1082 925
rect 1288 907 1290 925
rect 1496 907 1498 925
rect 1504 912 1506 974
rect 1704 972 1706 981
rect 1912 972 1914 981
rect 1702 971 1708 972
rect 1702 967 1703 971
rect 1707 967 1708 971
rect 1702 966 1708 967
rect 1910 971 1916 972
rect 1910 967 1911 971
rect 1915 967 1916 971
rect 1910 966 1916 967
rect 1982 963 1988 964
rect 1982 959 1983 963
rect 1987 959 1988 963
rect 1982 958 1988 959
rect 1702 930 1708 931
rect 1702 926 1703 930
rect 1707 926 1708 930
rect 1702 925 1708 926
rect 1910 930 1916 931
rect 1910 926 1911 930
rect 1915 926 1916 930
rect 1910 925 1916 926
rect 1502 911 1508 912
rect 1502 907 1503 911
rect 1507 907 1508 911
rect 1704 907 1706 925
rect 1912 907 1914 925
rect 1079 906 1083 907
rect 1079 901 1083 902
rect 1143 906 1147 907
rect 1143 901 1147 902
rect 1287 906 1291 907
rect 1287 901 1291 902
rect 1335 906 1339 907
rect 1335 901 1339 902
rect 1495 906 1499 907
rect 1502 906 1508 907
rect 1527 906 1531 907
rect 1495 901 1499 902
rect 1527 901 1531 902
rect 1703 906 1707 907
rect 1703 901 1707 902
rect 1719 906 1723 907
rect 1719 901 1723 902
rect 1911 906 1915 907
rect 1911 901 1915 902
rect 1144 891 1146 901
rect 1336 891 1338 901
rect 1528 891 1530 901
rect 1720 891 1722 901
rect 1912 891 1914 901
rect 1142 890 1148 891
rect 1142 886 1143 890
rect 1147 886 1148 890
rect 1142 885 1148 886
rect 1334 890 1340 891
rect 1334 886 1335 890
rect 1339 886 1340 890
rect 1334 885 1340 886
rect 1526 890 1532 891
rect 1526 886 1527 890
rect 1531 886 1532 890
rect 1526 885 1532 886
rect 1718 890 1724 891
rect 1718 886 1719 890
rect 1723 886 1724 890
rect 1718 885 1724 886
rect 1910 890 1916 891
rect 1910 886 1911 890
rect 1915 886 1916 890
rect 1910 885 1916 886
rect 1142 849 1148 850
rect 1142 845 1143 849
rect 1147 845 1148 849
rect 1142 844 1148 845
rect 1334 849 1340 850
rect 1334 845 1335 849
rect 1339 845 1340 849
rect 1334 844 1340 845
rect 1526 849 1532 850
rect 1526 845 1527 849
rect 1531 845 1532 849
rect 1526 844 1532 845
rect 1718 849 1724 850
rect 1718 845 1719 849
rect 1723 845 1724 849
rect 1718 844 1724 845
rect 1910 849 1916 850
rect 1910 845 1911 849
rect 1915 845 1916 849
rect 1910 844 1916 845
rect 1144 823 1146 844
rect 1336 823 1338 844
rect 1528 823 1530 844
rect 1720 823 1722 844
rect 1912 823 1914 844
rect 1984 840 1986 958
rect 2032 953 2034 981
rect 2072 959 2074 991
rect 2318 977 2324 978
rect 2318 973 2319 977
rect 2323 973 2324 977
rect 2318 972 2324 973
rect 2486 977 2492 978
rect 2486 973 2487 977
rect 2491 973 2492 977
rect 2486 972 2492 973
rect 2662 977 2668 978
rect 2662 973 2663 977
rect 2667 973 2668 977
rect 2662 972 2668 973
rect 2846 977 2852 978
rect 2846 973 2847 977
rect 2851 973 2852 977
rect 2846 972 2852 973
rect 2320 959 2322 972
rect 2488 959 2490 972
rect 2664 959 2666 972
rect 2670 967 2676 968
rect 2670 963 2671 967
rect 2675 963 2676 967
rect 2670 962 2676 963
rect 2071 958 2075 959
rect 2071 953 2075 954
rect 2151 958 2155 959
rect 2151 953 2155 954
rect 2287 958 2291 959
rect 2287 953 2291 954
rect 2319 958 2323 959
rect 2319 953 2323 954
rect 2431 958 2435 959
rect 2431 953 2435 954
rect 2487 958 2491 959
rect 2487 953 2491 954
rect 2591 958 2595 959
rect 2591 953 2595 954
rect 2663 958 2667 959
rect 2663 953 2667 954
rect 2030 952 2036 953
rect 2030 948 2031 952
rect 2035 948 2036 952
rect 2030 947 2036 948
rect 2030 935 2036 936
rect 2030 931 2031 935
rect 2035 931 2036 935
rect 2030 930 2036 931
rect 2032 907 2034 930
rect 2072 925 2074 953
rect 2152 944 2154 953
rect 2288 944 2290 953
rect 2432 944 2434 953
rect 2592 944 2594 953
rect 2150 943 2156 944
rect 2150 939 2151 943
rect 2155 939 2156 943
rect 2150 938 2156 939
rect 2286 943 2292 944
rect 2286 939 2287 943
rect 2291 939 2292 943
rect 2286 938 2292 939
rect 2430 943 2436 944
rect 2430 939 2431 943
rect 2435 939 2436 943
rect 2430 938 2436 939
rect 2590 943 2596 944
rect 2590 939 2591 943
rect 2595 939 2596 943
rect 2590 938 2596 939
rect 2672 936 2674 962
rect 2848 959 2850 972
rect 2880 968 2882 1094
rect 2894 1066 2900 1067
rect 2894 1062 2895 1066
rect 2899 1062 2900 1066
rect 2894 1061 2900 1062
rect 3086 1066 3092 1067
rect 3086 1062 3087 1066
rect 3091 1062 3092 1066
rect 3086 1061 3092 1062
rect 3286 1066 3292 1067
rect 3286 1062 3287 1066
rect 3291 1062 3292 1066
rect 3286 1061 3292 1062
rect 3494 1066 3500 1067
rect 3494 1062 3495 1066
rect 3499 1062 3500 1066
rect 3494 1061 3500 1062
rect 3702 1066 3708 1067
rect 3702 1062 3703 1066
rect 3707 1062 3708 1066
rect 3702 1061 3708 1062
rect 2896 1035 2898 1061
rect 3088 1035 3090 1061
rect 3288 1035 3290 1061
rect 3496 1035 3498 1061
rect 3704 1035 3706 1061
rect 2895 1034 2899 1035
rect 2895 1029 2899 1030
rect 3039 1034 3043 1035
rect 3039 1029 3043 1030
rect 3087 1034 3091 1035
rect 3087 1029 3091 1030
rect 3247 1034 3251 1035
rect 3247 1029 3251 1030
rect 3287 1034 3291 1035
rect 3287 1029 3291 1030
rect 3463 1034 3467 1035
rect 3463 1029 3467 1030
rect 3495 1034 3499 1035
rect 3495 1029 3499 1030
rect 3687 1034 3691 1035
rect 3687 1029 3691 1030
rect 3703 1034 3707 1035
rect 3703 1029 3707 1030
rect 3040 1019 3042 1029
rect 3248 1019 3250 1029
rect 3464 1019 3466 1029
rect 3688 1019 3690 1029
rect 3038 1018 3044 1019
rect 3038 1014 3039 1018
rect 3043 1014 3044 1018
rect 3038 1013 3044 1014
rect 3246 1018 3252 1019
rect 3246 1014 3247 1018
rect 3251 1014 3252 1018
rect 3246 1013 3252 1014
rect 3462 1018 3468 1019
rect 3462 1014 3463 1018
rect 3467 1014 3468 1018
rect 3462 1013 3468 1014
rect 3686 1018 3692 1019
rect 3686 1014 3687 1018
rect 3691 1014 3692 1018
rect 3686 1013 3692 1014
rect 3760 988 3762 1110
rect 3896 1108 3898 1117
rect 3968 1116 3970 1146
rect 3992 1123 3994 1155
rect 3991 1122 3995 1123
rect 3991 1117 3995 1118
rect 3966 1115 3972 1116
rect 3966 1111 3967 1115
rect 3971 1111 3972 1115
rect 3966 1110 3972 1111
rect 3894 1107 3900 1108
rect 3894 1103 3895 1107
rect 3899 1103 3900 1107
rect 3894 1102 3900 1103
rect 3958 1099 3964 1100
rect 3958 1095 3959 1099
rect 3963 1095 3964 1099
rect 3958 1094 3964 1095
rect 3894 1066 3900 1067
rect 3894 1062 3895 1066
rect 3899 1062 3900 1066
rect 3894 1061 3900 1062
rect 3896 1035 3898 1061
rect 3895 1034 3899 1035
rect 3895 1029 3899 1030
rect 3896 1019 3898 1029
rect 3894 1018 3900 1019
rect 3894 1014 3895 1018
rect 3899 1014 3900 1018
rect 3894 1013 3900 1014
rect 3446 987 3452 988
rect 3446 983 3447 987
rect 3451 983 3452 987
rect 3446 982 3452 983
rect 3758 987 3764 988
rect 3758 983 3759 987
rect 3763 983 3764 987
rect 3758 982 3764 983
rect 3038 977 3044 978
rect 3038 973 3039 977
rect 3043 973 3044 977
rect 3038 972 3044 973
rect 3246 977 3252 978
rect 3246 973 3247 977
rect 3251 973 3252 977
rect 3246 972 3252 973
rect 2878 967 2884 968
rect 2878 963 2879 967
rect 2883 963 2884 967
rect 2878 962 2884 963
rect 3040 959 3042 972
rect 3214 967 3220 968
rect 3214 963 3215 967
rect 3219 963 3220 967
rect 3214 962 3220 963
rect 2759 958 2763 959
rect 2759 953 2763 954
rect 2847 958 2851 959
rect 2847 953 2851 954
rect 2935 958 2939 959
rect 2935 953 2939 954
rect 3039 958 3043 959
rect 3039 953 3043 954
rect 3119 958 3123 959
rect 3119 953 3123 954
rect 2760 944 2762 953
rect 2830 951 2836 952
rect 2830 947 2831 951
rect 2835 947 2836 951
rect 2830 946 2836 947
rect 2758 943 2764 944
rect 2758 939 2759 943
rect 2763 939 2764 943
rect 2758 938 2764 939
rect 2270 935 2276 936
rect 2270 931 2271 935
rect 2275 931 2276 935
rect 2270 930 2276 931
rect 2670 935 2676 936
rect 2670 931 2671 935
rect 2675 931 2676 935
rect 2670 930 2676 931
rect 2070 924 2076 925
rect 2070 920 2071 924
rect 2075 920 2076 924
rect 2070 919 2076 920
rect 2070 907 2076 908
rect 2031 906 2035 907
rect 2070 903 2071 907
rect 2075 903 2076 907
rect 2070 902 2076 903
rect 2150 902 2156 903
rect 2031 901 2035 902
rect 2032 886 2034 901
rect 2030 885 2036 886
rect 2030 881 2031 885
rect 2035 881 2036 885
rect 2030 880 2036 881
rect 2072 875 2074 902
rect 2150 898 2151 902
rect 2155 898 2156 902
rect 2150 897 2156 898
rect 2152 875 2154 897
rect 2071 874 2075 875
rect 2071 869 2075 870
rect 2111 874 2115 875
rect 2111 869 2115 870
rect 2151 874 2155 875
rect 2151 869 2155 870
rect 2239 874 2243 875
rect 2239 869 2243 870
rect 2030 868 2036 869
rect 2030 864 2031 868
rect 2035 864 2036 868
rect 2030 863 2036 864
rect 1982 839 1988 840
rect 1982 835 1983 839
rect 1987 835 1988 839
rect 1982 834 1988 835
rect 2032 823 2034 863
rect 2072 854 2074 869
rect 2112 859 2114 869
rect 2240 859 2242 869
rect 2110 858 2116 859
rect 2110 854 2111 858
rect 2115 854 2116 858
rect 2070 853 2076 854
rect 2110 853 2116 854
rect 2238 858 2244 859
rect 2238 854 2239 858
rect 2243 854 2244 858
rect 2238 853 2244 854
rect 2070 849 2071 853
rect 2075 849 2076 853
rect 2070 848 2076 849
rect 2070 836 2076 837
rect 2070 832 2071 836
rect 2075 832 2076 836
rect 2070 831 2076 832
rect 1031 822 1035 823
rect 1031 817 1035 818
rect 1143 822 1147 823
rect 1143 817 1147 818
rect 1239 822 1243 823
rect 1239 817 1243 818
rect 1335 822 1339 823
rect 1335 817 1339 818
rect 1471 822 1475 823
rect 1471 817 1475 818
rect 1527 822 1531 823
rect 1527 817 1531 818
rect 1711 822 1715 823
rect 1711 817 1715 818
rect 1719 822 1723 823
rect 1719 817 1723 818
rect 1911 822 1915 823
rect 1911 817 1915 818
rect 1935 822 1939 823
rect 1935 817 1939 818
rect 2031 822 2035 823
rect 2031 817 2035 818
rect 1032 808 1034 817
rect 1240 808 1242 817
rect 1472 808 1474 817
rect 1712 808 1714 817
rect 1726 815 1732 816
rect 1726 811 1727 815
rect 1731 811 1732 815
rect 1726 810 1732 811
rect 1030 807 1036 808
rect 1030 803 1031 807
rect 1035 803 1036 807
rect 1030 802 1036 803
rect 1238 807 1244 808
rect 1238 803 1239 807
rect 1243 803 1244 807
rect 1238 802 1244 803
rect 1470 807 1476 808
rect 1470 803 1471 807
rect 1475 803 1476 807
rect 1470 802 1476 803
rect 1710 807 1716 808
rect 1710 803 1711 807
rect 1715 803 1716 807
rect 1710 802 1716 803
rect 350 799 356 800
rect 350 795 351 799
rect 355 795 356 799
rect 350 794 356 795
rect 998 799 1004 800
rect 998 795 999 799
rect 1003 795 1004 799
rect 998 794 1004 795
rect 110 788 116 789
rect 110 784 111 788
rect 115 784 116 788
rect 110 783 116 784
rect 110 771 116 772
rect 110 767 111 771
rect 115 767 116 771
rect 110 766 116 767
rect 262 766 268 767
rect 112 747 114 766
rect 262 762 263 766
rect 267 762 268 766
rect 262 761 268 762
rect 264 747 266 761
rect 111 746 115 747
rect 111 741 115 742
rect 263 746 267 747
rect 263 741 267 742
rect 112 726 114 741
rect 110 725 116 726
rect 110 721 111 725
rect 115 721 116 725
rect 110 720 116 721
rect 110 708 116 709
rect 110 704 111 708
rect 115 704 116 708
rect 110 703 116 704
rect 112 663 114 703
rect 352 680 354 794
rect 366 766 372 767
rect 366 762 367 766
rect 371 762 372 766
rect 366 761 372 762
rect 478 766 484 767
rect 478 762 479 766
rect 483 762 484 766
rect 478 761 484 762
rect 590 766 596 767
rect 590 762 591 766
rect 595 762 596 766
rect 590 761 596 762
rect 710 766 716 767
rect 710 762 711 766
rect 715 762 716 766
rect 710 761 716 762
rect 854 766 860 767
rect 854 762 855 766
rect 859 762 860 766
rect 854 761 860 762
rect 1030 766 1036 767
rect 1030 762 1031 766
rect 1035 762 1036 766
rect 1030 761 1036 762
rect 1238 766 1244 767
rect 1238 762 1239 766
rect 1243 762 1244 766
rect 1238 761 1244 762
rect 1470 766 1476 767
rect 1470 762 1471 766
rect 1475 762 1476 766
rect 1470 761 1476 762
rect 1710 766 1716 767
rect 1710 762 1711 766
rect 1715 762 1716 766
rect 1710 761 1716 762
rect 368 747 370 761
rect 480 747 482 761
rect 592 747 594 761
rect 712 747 714 761
rect 856 747 858 761
rect 1032 747 1034 761
rect 1078 747 1084 748
rect 1240 747 1242 761
rect 1472 747 1474 761
rect 1712 747 1714 761
rect 1728 748 1730 810
rect 1936 808 1938 817
rect 2010 815 2016 816
rect 2010 811 2011 815
rect 2015 811 2016 815
rect 2010 810 2016 811
rect 1934 807 1940 808
rect 1934 803 1935 807
rect 1939 803 1940 807
rect 1934 802 1940 803
rect 2012 796 2014 810
rect 1926 795 1932 796
rect 1926 791 1927 795
rect 1931 791 1932 795
rect 1926 790 1932 791
rect 2010 795 2016 796
rect 2010 791 2011 795
rect 2015 791 2016 795
rect 2010 790 2016 791
rect 1726 747 1732 748
rect 367 746 371 747
rect 367 741 371 742
rect 423 746 427 747
rect 423 741 427 742
rect 479 746 483 747
rect 479 741 483 742
rect 527 746 531 747
rect 527 741 531 742
rect 591 746 595 747
rect 591 741 595 742
rect 639 746 643 747
rect 639 741 643 742
rect 711 746 715 747
rect 711 741 715 742
rect 759 746 763 747
rect 759 741 763 742
rect 855 746 859 747
rect 855 741 859 742
rect 879 746 883 747
rect 879 741 883 742
rect 1007 746 1011 747
rect 1007 741 1011 742
rect 1031 746 1035 747
rect 1078 743 1079 747
rect 1083 743 1084 747
rect 1078 742 1084 743
rect 1143 746 1147 747
rect 1031 741 1035 742
rect 424 731 426 741
rect 528 731 530 741
rect 640 731 642 741
rect 760 731 762 741
rect 880 731 882 741
rect 1008 731 1010 741
rect 422 730 428 731
rect 422 726 423 730
rect 427 726 428 730
rect 422 725 428 726
rect 526 730 532 731
rect 526 726 527 730
rect 531 726 532 730
rect 526 725 532 726
rect 638 730 644 731
rect 638 726 639 730
rect 643 726 644 730
rect 638 725 644 726
rect 758 730 764 731
rect 758 726 759 730
rect 763 726 764 730
rect 758 725 764 726
rect 878 730 884 731
rect 878 726 879 730
rect 883 726 884 730
rect 878 725 884 726
rect 1006 730 1012 731
rect 1006 726 1007 730
rect 1011 726 1012 730
rect 1006 725 1012 726
rect 1080 700 1082 742
rect 1143 741 1147 742
rect 1239 746 1243 747
rect 1239 741 1243 742
rect 1287 746 1291 747
rect 1287 741 1291 742
rect 1447 746 1451 747
rect 1447 741 1451 742
rect 1471 746 1475 747
rect 1471 741 1475 742
rect 1615 746 1619 747
rect 1615 741 1619 742
rect 1711 746 1715 747
rect 1726 743 1727 747
rect 1731 743 1732 747
rect 1726 742 1732 743
rect 1783 746 1787 747
rect 1711 741 1715 742
rect 1783 741 1787 742
rect 1144 731 1146 741
rect 1288 731 1290 741
rect 1448 731 1450 741
rect 1616 731 1618 741
rect 1784 731 1786 741
rect 1142 730 1148 731
rect 1142 726 1143 730
rect 1147 726 1148 730
rect 1142 725 1148 726
rect 1286 730 1292 731
rect 1286 726 1287 730
rect 1291 726 1292 730
rect 1286 725 1292 726
rect 1446 730 1452 731
rect 1446 726 1447 730
rect 1451 726 1452 730
rect 1446 725 1452 726
rect 1614 730 1620 731
rect 1614 726 1615 730
rect 1619 726 1620 730
rect 1614 725 1620 726
rect 1782 730 1788 731
rect 1782 726 1783 730
rect 1787 726 1788 730
rect 1782 725 1788 726
rect 510 699 516 700
rect 510 695 511 699
rect 515 695 516 699
rect 510 694 516 695
rect 622 699 628 700
rect 622 695 623 699
rect 627 695 628 699
rect 622 694 628 695
rect 742 699 748 700
rect 742 695 743 699
rect 747 695 748 699
rect 742 694 748 695
rect 862 699 868 700
rect 862 695 863 699
rect 867 695 868 699
rect 862 694 868 695
rect 870 699 876 700
rect 870 695 871 699
rect 875 695 876 699
rect 870 694 876 695
rect 1078 699 1084 700
rect 1078 695 1079 699
rect 1083 695 1084 699
rect 1078 694 1084 695
rect 1890 699 1896 700
rect 1890 695 1891 699
rect 1895 695 1896 699
rect 1890 694 1896 695
rect 422 689 428 690
rect 422 685 423 689
rect 427 685 428 689
rect 422 684 428 685
rect 350 679 356 680
rect 350 675 351 679
rect 355 675 356 679
rect 350 674 356 675
rect 424 663 426 684
rect 512 680 514 694
rect 526 689 532 690
rect 526 685 527 689
rect 531 685 532 689
rect 526 684 532 685
rect 510 679 516 680
rect 510 675 511 679
rect 515 675 516 679
rect 510 674 516 675
rect 528 663 530 684
rect 624 680 626 694
rect 638 689 644 690
rect 638 685 639 689
rect 643 685 644 689
rect 638 684 644 685
rect 622 679 628 680
rect 622 675 623 679
rect 627 675 628 679
rect 622 674 628 675
rect 640 663 642 684
rect 744 680 746 694
rect 758 689 764 690
rect 758 685 759 689
rect 763 685 764 689
rect 758 684 764 685
rect 742 679 748 680
rect 742 675 743 679
rect 747 675 748 679
rect 742 674 748 675
rect 678 667 684 668
rect 678 663 679 667
rect 683 663 684 667
rect 760 663 762 684
rect 864 680 866 694
rect 862 679 868 680
rect 862 675 863 679
rect 867 675 868 679
rect 862 674 868 675
rect 111 662 115 663
rect 111 657 115 658
rect 423 662 427 663
rect 423 657 427 658
rect 527 662 531 663
rect 527 657 531 658
rect 591 662 595 663
rect 591 657 595 658
rect 639 662 643 663
rect 678 662 684 663
rect 695 662 699 663
rect 639 657 643 658
rect 112 629 114 657
rect 592 648 594 657
rect 590 647 596 648
rect 590 643 591 647
rect 595 643 596 647
rect 590 642 596 643
rect 680 640 682 662
rect 695 657 699 658
rect 759 662 763 663
rect 759 657 763 658
rect 807 662 811 663
rect 872 660 874 694
rect 878 689 884 690
rect 878 685 879 689
rect 883 685 884 689
rect 878 684 884 685
rect 1006 689 1012 690
rect 1006 685 1007 689
rect 1011 685 1012 689
rect 1006 684 1012 685
rect 1142 689 1148 690
rect 1142 685 1143 689
rect 1147 685 1148 689
rect 1142 684 1148 685
rect 1286 689 1292 690
rect 1286 685 1287 689
rect 1291 685 1292 689
rect 1286 684 1292 685
rect 1446 689 1452 690
rect 1446 685 1447 689
rect 1451 685 1452 689
rect 1446 684 1452 685
rect 1614 689 1620 690
rect 1614 685 1615 689
rect 1619 685 1620 689
rect 1614 684 1620 685
rect 1782 689 1788 690
rect 1782 685 1783 689
rect 1787 685 1788 689
rect 1782 684 1788 685
rect 880 663 882 684
rect 1008 663 1010 684
rect 1144 663 1146 684
rect 1246 671 1252 672
rect 1246 667 1247 671
rect 1251 667 1252 671
rect 1246 666 1252 667
rect 879 662 883 663
rect 807 657 811 658
rect 870 659 876 660
rect 696 648 698 657
rect 808 648 810 657
rect 870 655 871 659
rect 875 655 876 659
rect 879 657 883 658
rect 919 662 923 663
rect 919 657 923 658
rect 1007 662 1011 663
rect 1007 657 1011 658
rect 1031 662 1035 663
rect 1031 657 1035 658
rect 1143 662 1147 663
rect 1143 657 1147 658
rect 870 654 876 655
rect 920 648 922 657
rect 1032 648 1034 657
rect 1144 648 1146 657
rect 694 647 700 648
rect 694 643 695 647
rect 699 643 700 647
rect 694 642 700 643
rect 806 647 812 648
rect 806 643 807 647
rect 811 643 812 647
rect 806 642 812 643
rect 918 647 924 648
rect 918 643 919 647
rect 923 643 924 647
rect 918 642 924 643
rect 1030 647 1036 648
rect 1030 643 1031 647
rect 1035 643 1036 647
rect 1030 642 1036 643
rect 1142 647 1148 648
rect 1142 643 1143 647
rect 1147 643 1148 647
rect 1142 642 1148 643
rect 1248 640 1250 666
rect 1288 663 1290 684
rect 1448 663 1450 684
rect 1616 663 1618 684
rect 1784 663 1786 684
rect 1892 672 1894 694
rect 1928 680 1930 790
rect 2032 789 2034 817
rect 2072 803 2074 831
rect 2182 827 2188 828
rect 2182 823 2183 827
rect 2187 823 2188 827
rect 2182 822 2188 823
rect 2110 817 2116 818
rect 2110 813 2111 817
rect 2115 813 2116 817
rect 2110 812 2116 813
rect 2112 803 2114 812
rect 2071 802 2075 803
rect 2071 797 2075 798
rect 2111 802 2115 803
rect 2111 797 2115 798
rect 2030 788 2036 789
rect 2030 784 2031 788
rect 2035 784 2036 788
rect 2030 783 2036 784
rect 2030 771 2036 772
rect 2030 767 2031 771
rect 2035 767 2036 771
rect 2072 769 2074 797
rect 2112 788 2114 797
rect 2184 796 2186 822
rect 2238 817 2244 818
rect 2238 813 2239 817
rect 2243 813 2244 817
rect 2238 812 2244 813
rect 2240 803 2242 812
rect 2272 808 2274 930
rect 2286 902 2292 903
rect 2286 898 2287 902
rect 2291 898 2292 902
rect 2286 897 2292 898
rect 2430 902 2436 903
rect 2430 898 2431 902
rect 2435 898 2436 902
rect 2430 897 2436 898
rect 2590 902 2596 903
rect 2590 898 2591 902
rect 2595 898 2596 902
rect 2590 897 2596 898
rect 2758 902 2764 903
rect 2758 898 2759 902
rect 2763 898 2764 902
rect 2758 897 2764 898
rect 2288 875 2290 897
rect 2432 875 2434 897
rect 2592 875 2594 897
rect 2760 875 2762 897
rect 2287 874 2291 875
rect 2287 869 2291 870
rect 2407 874 2411 875
rect 2407 869 2411 870
rect 2431 874 2435 875
rect 2431 869 2435 870
rect 2575 874 2579 875
rect 2575 869 2579 870
rect 2591 874 2595 875
rect 2591 869 2595 870
rect 2751 874 2755 875
rect 2751 869 2755 870
rect 2759 874 2763 875
rect 2759 869 2763 870
rect 2408 859 2410 869
rect 2576 859 2578 869
rect 2752 859 2754 869
rect 2406 858 2412 859
rect 2406 854 2407 858
rect 2411 854 2412 858
rect 2406 853 2412 854
rect 2574 858 2580 859
rect 2574 854 2575 858
rect 2579 854 2580 858
rect 2574 853 2580 854
rect 2750 858 2756 859
rect 2750 854 2751 858
rect 2755 854 2756 858
rect 2750 853 2756 854
rect 2832 828 2834 946
rect 2936 944 2938 953
rect 3120 944 3122 953
rect 2934 943 2940 944
rect 2934 939 2935 943
rect 2939 939 2940 943
rect 2934 938 2940 939
rect 3118 943 3124 944
rect 3118 939 3119 943
rect 3123 939 3124 943
rect 3118 938 3124 939
rect 3216 936 3218 962
rect 3248 959 3250 972
rect 3448 968 3450 982
rect 3462 977 3468 978
rect 3462 973 3463 977
rect 3467 973 3468 977
rect 3462 972 3468 973
rect 3686 977 3692 978
rect 3686 973 3687 977
rect 3691 973 3692 977
rect 3686 972 3692 973
rect 3894 977 3900 978
rect 3894 973 3895 977
rect 3899 973 3900 977
rect 3894 972 3900 973
rect 3446 967 3452 968
rect 3446 963 3447 967
rect 3451 963 3452 967
rect 3446 962 3452 963
rect 3464 959 3466 972
rect 3688 959 3690 972
rect 3896 959 3898 972
rect 3960 968 3962 1094
rect 3992 1089 3994 1117
rect 3990 1088 3996 1089
rect 3990 1084 3991 1088
rect 3995 1084 3996 1088
rect 3990 1083 3996 1084
rect 3990 1071 3996 1072
rect 3990 1067 3991 1071
rect 3995 1067 3996 1071
rect 3990 1066 3996 1067
rect 3992 1035 3994 1066
rect 3991 1034 3995 1035
rect 3991 1029 3995 1030
rect 3992 1014 3994 1029
rect 3990 1013 3996 1014
rect 3990 1009 3991 1013
rect 3995 1009 3996 1013
rect 3990 1008 3996 1009
rect 3990 996 3996 997
rect 3990 992 3991 996
rect 3995 992 3996 996
rect 3990 991 3996 992
rect 3966 987 3972 988
rect 3966 983 3967 987
rect 3971 983 3972 987
rect 3966 982 3972 983
rect 3958 967 3964 968
rect 3958 963 3959 967
rect 3963 963 3964 967
rect 3958 962 3964 963
rect 3247 958 3251 959
rect 3247 953 3251 954
rect 3311 958 3315 959
rect 3311 953 3315 954
rect 3463 958 3467 959
rect 3463 953 3467 954
rect 3511 958 3515 959
rect 3511 953 3515 954
rect 3687 958 3691 959
rect 3687 953 3691 954
rect 3711 958 3715 959
rect 3711 953 3715 954
rect 3895 958 3899 959
rect 3895 953 3899 954
rect 3312 944 3314 953
rect 3512 944 3514 953
rect 3712 944 3714 953
rect 3782 951 3788 952
rect 3782 947 3783 951
rect 3787 947 3788 951
rect 3782 946 3788 947
rect 3310 943 3316 944
rect 3310 939 3311 943
rect 3315 939 3316 943
rect 3310 938 3316 939
rect 3510 943 3516 944
rect 3510 939 3511 943
rect 3515 939 3516 943
rect 3510 938 3516 939
rect 3710 943 3716 944
rect 3710 939 3711 943
rect 3715 939 3716 943
rect 3710 938 3716 939
rect 3214 935 3220 936
rect 3214 931 3215 935
rect 3219 931 3220 935
rect 3214 930 3220 931
rect 2934 902 2940 903
rect 2934 898 2935 902
rect 2939 898 2940 902
rect 2934 897 2940 898
rect 3118 902 3124 903
rect 3118 898 3119 902
rect 3123 898 3124 902
rect 3118 897 3124 898
rect 3310 902 3316 903
rect 3310 898 3311 902
rect 3315 898 3316 902
rect 3310 897 3316 898
rect 3510 902 3516 903
rect 3510 898 3511 902
rect 3515 898 3516 902
rect 3510 897 3516 898
rect 3710 902 3716 903
rect 3710 898 3711 902
rect 3715 898 3716 902
rect 3710 897 3716 898
rect 2936 875 2938 897
rect 3120 875 3122 897
rect 3312 875 3314 897
rect 3512 875 3514 897
rect 3712 875 3714 897
rect 2935 874 2939 875
rect 2935 869 2939 870
rect 3119 874 3123 875
rect 3119 869 3123 870
rect 3311 874 3315 875
rect 3311 869 3315 870
rect 3511 874 3515 875
rect 3511 869 3515 870
rect 3711 874 3715 875
rect 3711 869 3715 870
rect 2936 859 2938 869
rect 3120 859 3122 869
rect 3312 859 3314 869
rect 3512 859 3514 869
rect 3712 859 3714 869
rect 2934 858 2940 859
rect 2934 854 2935 858
rect 2939 854 2940 858
rect 2934 853 2940 854
rect 3118 858 3124 859
rect 3118 854 3119 858
rect 3123 854 3124 858
rect 3118 853 3124 854
rect 3310 858 3316 859
rect 3310 854 3311 858
rect 3315 854 3316 858
rect 3310 853 3316 854
rect 3510 858 3516 859
rect 3510 854 3511 858
rect 3515 854 3516 858
rect 3510 853 3516 854
rect 3710 858 3716 859
rect 3710 854 3711 858
rect 3715 854 3716 858
rect 3710 853 3716 854
rect 3784 828 3786 946
rect 3896 944 3898 953
rect 3968 952 3970 982
rect 3992 959 3994 991
rect 3991 958 3995 959
rect 3991 953 3995 954
rect 3966 951 3972 952
rect 3966 947 3967 951
rect 3971 947 3972 951
rect 3966 946 3972 947
rect 3894 943 3900 944
rect 3894 939 3895 943
rect 3899 939 3900 943
rect 3894 938 3900 939
rect 3958 935 3964 936
rect 3958 931 3959 935
rect 3963 931 3964 935
rect 3958 930 3964 931
rect 3894 902 3900 903
rect 3894 898 3895 902
rect 3899 898 3900 902
rect 3894 897 3900 898
rect 3896 875 3898 897
rect 3895 874 3899 875
rect 3895 869 3899 870
rect 3896 859 3898 869
rect 3894 858 3900 859
rect 3894 854 3895 858
rect 3899 854 3900 858
rect 3894 853 3900 854
rect 2558 827 2564 828
rect 2558 823 2559 827
rect 2563 823 2564 827
rect 2558 822 2564 823
rect 2734 827 2740 828
rect 2734 823 2735 827
rect 2739 823 2740 827
rect 2734 822 2740 823
rect 2830 827 2836 828
rect 2830 823 2831 827
rect 2835 823 2836 827
rect 2830 822 2836 823
rect 3494 827 3500 828
rect 3494 823 3495 827
rect 3499 823 3500 827
rect 3494 822 3500 823
rect 3694 827 3700 828
rect 3694 823 3695 827
rect 3699 823 3700 827
rect 3694 822 3700 823
rect 3782 827 3788 828
rect 3782 823 3783 827
rect 3787 823 3788 827
rect 3782 822 3788 823
rect 2406 817 2412 818
rect 2406 813 2407 817
rect 2411 813 2412 817
rect 2406 812 2412 813
rect 2270 807 2276 808
rect 2270 803 2271 807
rect 2275 803 2276 807
rect 2408 803 2410 812
rect 2560 808 2562 822
rect 2574 817 2580 818
rect 2574 813 2575 817
rect 2579 813 2580 817
rect 2574 812 2580 813
rect 2454 807 2460 808
rect 2454 803 2455 807
rect 2459 803 2460 807
rect 2239 802 2243 803
rect 2270 802 2276 803
rect 2391 802 2395 803
rect 2239 797 2243 798
rect 2391 797 2395 798
rect 2407 802 2411 803
rect 2454 802 2460 803
rect 2558 807 2564 808
rect 2558 803 2559 807
rect 2563 803 2564 807
rect 2576 803 2578 812
rect 2736 808 2738 822
rect 2750 817 2756 818
rect 2750 813 2751 817
rect 2755 813 2756 817
rect 2750 812 2756 813
rect 2934 817 2940 818
rect 2934 813 2935 817
rect 2939 813 2940 817
rect 2934 812 2940 813
rect 3118 817 3124 818
rect 3118 813 3119 817
rect 3123 813 3124 817
rect 3118 812 3124 813
rect 3310 817 3316 818
rect 3310 813 3311 817
rect 3315 813 3316 817
rect 3310 812 3316 813
rect 2734 807 2740 808
rect 2734 803 2735 807
rect 2739 803 2740 807
rect 2752 803 2754 812
rect 2936 803 2938 812
rect 3120 803 3122 812
rect 3270 807 3276 808
rect 3270 803 3271 807
rect 3275 803 3276 807
rect 3312 803 3314 812
rect 3496 808 3498 822
rect 3510 817 3516 818
rect 3510 813 3511 817
rect 3515 813 3516 817
rect 3510 812 3516 813
rect 3494 807 3500 808
rect 3494 803 3495 807
rect 3499 803 3500 807
rect 3512 803 3514 812
rect 3696 808 3698 822
rect 3710 817 3716 818
rect 3710 813 3711 817
rect 3715 813 3716 817
rect 3710 812 3716 813
rect 3894 817 3900 818
rect 3894 813 3895 817
rect 3899 813 3900 817
rect 3894 812 3900 813
rect 3694 807 3700 808
rect 3694 803 3695 807
rect 3699 803 3700 807
rect 3712 803 3714 812
rect 3896 803 3898 812
rect 3960 808 3962 930
rect 3992 925 3994 953
rect 3990 924 3996 925
rect 3990 920 3991 924
rect 3995 920 3996 924
rect 3990 919 3996 920
rect 3990 907 3996 908
rect 3990 903 3991 907
rect 3995 903 3996 907
rect 3990 902 3996 903
rect 3992 875 3994 902
rect 3991 874 3995 875
rect 3991 869 3995 870
rect 3992 854 3994 869
rect 3990 853 3996 854
rect 3990 849 3991 853
rect 3995 849 3996 853
rect 3990 848 3996 849
rect 3990 836 3996 837
rect 3990 832 3991 836
rect 3995 832 3996 836
rect 3990 831 3996 832
rect 3966 827 3972 828
rect 3966 823 3967 827
rect 3971 823 3972 827
rect 3966 822 3972 823
rect 3958 807 3964 808
rect 3958 803 3959 807
rect 3963 803 3964 807
rect 2558 802 2564 803
rect 2575 802 2579 803
rect 2407 797 2411 798
rect 2182 795 2188 796
rect 2182 791 2183 795
rect 2187 791 2188 795
rect 2182 790 2188 791
rect 2392 788 2394 797
rect 2110 787 2116 788
rect 2110 783 2111 787
rect 2115 783 2116 787
rect 2110 782 2116 783
rect 2390 787 2396 788
rect 2390 783 2391 787
rect 2395 783 2396 787
rect 2390 782 2396 783
rect 2456 780 2458 802
rect 2575 797 2579 798
rect 2679 802 2683 803
rect 2734 802 2740 803
rect 2751 802 2755 803
rect 2679 797 2683 798
rect 2751 797 2755 798
rect 2935 802 2939 803
rect 2935 797 2939 798
rect 2951 802 2955 803
rect 2951 797 2955 798
rect 3119 802 3123 803
rect 3119 797 3123 798
rect 3199 802 3203 803
rect 3270 802 3276 803
rect 3311 802 3315 803
rect 3199 797 3203 798
rect 2462 795 2468 796
rect 2462 791 2463 795
rect 2467 791 2468 795
rect 2462 790 2468 791
rect 2454 779 2460 780
rect 2454 775 2455 779
rect 2459 775 2460 779
rect 2454 774 2460 775
rect 1934 766 1940 767
rect 2030 766 2036 767
rect 2070 768 2076 769
rect 1934 762 1935 766
rect 1939 762 1940 766
rect 1934 761 1940 762
rect 1936 747 1938 761
rect 2032 747 2034 766
rect 2070 764 2071 768
rect 2075 764 2076 768
rect 2070 763 2076 764
rect 2070 751 2076 752
rect 2070 747 2071 751
rect 2075 747 2076 751
rect 1935 746 1939 747
rect 1935 741 1939 742
rect 2031 746 2035 747
rect 2070 746 2076 747
rect 2110 746 2116 747
rect 2031 741 2035 742
rect 1936 731 1938 741
rect 1934 730 1940 731
rect 1934 726 1935 730
rect 1939 726 1940 730
rect 2032 726 2034 741
rect 1934 725 1940 726
rect 2030 725 2036 726
rect 2030 721 2031 725
rect 2035 721 2036 725
rect 2072 723 2074 746
rect 2110 742 2111 746
rect 2115 742 2116 746
rect 2110 741 2116 742
rect 2390 746 2396 747
rect 2390 742 2391 746
rect 2395 742 2396 746
rect 2390 741 2396 742
rect 2112 723 2114 741
rect 2392 723 2394 741
rect 2030 720 2036 721
rect 2071 722 2075 723
rect 2071 717 2075 718
rect 2111 722 2115 723
rect 2111 717 2115 718
rect 2327 722 2331 723
rect 2327 717 2331 718
rect 2391 722 2395 723
rect 2391 717 2395 718
rect 2030 708 2036 709
rect 2030 704 2031 708
rect 2035 704 2036 708
rect 2030 703 2036 704
rect 1934 689 1940 690
rect 1934 685 1935 689
rect 1939 685 1940 689
rect 1934 684 1940 685
rect 1926 679 1932 680
rect 1926 675 1927 679
rect 1931 675 1932 679
rect 1926 674 1932 675
rect 1890 671 1896 672
rect 1890 667 1891 671
rect 1895 667 1896 671
rect 1890 666 1896 667
rect 1936 663 1938 684
rect 2032 663 2034 703
rect 2072 702 2074 717
rect 2112 707 2114 717
rect 2328 707 2330 717
rect 2110 706 2116 707
rect 2110 702 2111 706
rect 2115 702 2116 706
rect 2070 701 2076 702
rect 2110 701 2116 702
rect 2326 706 2332 707
rect 2326 702 2327 706
rect 2331 702 2332 706
rect 2326 701 2332 702
rect 2062 699 2068 700
rect 2062 695 2063 699
rect 2067 695 2068 699
rect 2070 697 2071 701
rect 2075 697 2076 701
rect 2070 696 2076 697
rect 2062 694 2068 695
rect 1263 662 1267 663
rect 1263 657 1267 658
rect 1287 662 1291 663
rect 1287 657 1291 658
rect 1383 662 1387 663
rect 1383 657 1387 658
rect 1447 662 1451 663
rect 1447 657 1451 658
rect 1503 662 1507 663
rect 1503 657 1507 658
rect 1615 662 1619 663
rect 1615 657 1619 658
rect 1623 662 1627 663
rect 1623 657 1627 658
rect 1783 662 1787 663
rect 1783 657 1787 658
rect 1935 662 1939 663
rect 1935 657 1939 658
rect 2031 662 2035 663
rect 2031 657 2035 658
rect 1264 648 1266 657
rect 1384 648 1386 657
rect 1504 648 1506 657
rect 1624 648 1626 657
rect 1262 647 1268 648
rect 1262 643 1263 647
rect 1267 643 1268 647
rect 1262 642 1268 643
rect 1382 647 1388 648
rect 1382 643 1383 647
rect 1387 643 1388 647
rect 1382 642 1388 643
rect 1502 647 1508 648
rect 1502 643 1503 647
rect 1507 643 1508 647
rect 1502 642 1508 643
rect 1566 647 1572 648
rect 1566 643 1567 647
rect 1571 643 1572 647
rect 1566 642 1572 643
rect 1622 647 1628 648
rect 1622 643 1623 647
rect 1627 643 1628 647
rect 1622 642 1628 643
rect 678 639 684 640
rect 678 635 679 639
rect 683 635 684 639
rect 1246 639 1252 640
rect 678 634 684 635
rect 942 635 948 636
rect 942 631 943 635
rect 947 631 948 635
rect 1246 635 1247 639
rect 1251 635 1252 639
rect 1246 634 1252 635
rect 942 630 948 631
rect 110 628 116 629
rect 110 624 111 628
rect 115 624 116 628
rect 110 623 116 624
rect 110 611 116 612
rect 110 607 111 611
rect 115 607 116 611
rect 110 606 116 607
rect 590 606 596 607
rect 112 583 114 606
rect 590 602 591 606
rect 595 602 596 606
rect 590 601 596 602
rect 694 606 700 607
rect 694 602 695 606
rect 699 602 700 606
rect 694 601 700 602
rect 806 606 812 607
rect 806 602 807 606
rect 811 602 812 606
rect 806 601 812 602
rect 918 606 924 607
rect 918 602 919 606
rect 923 602 924 606
rect 918 601 924 602
rect 592 583 594 601
rect 696 583 698 601
rect 808 583 810 601
rect 920 583 922 601
rect 111 582 115 583
rect 111 577 115 578
rect 591 582 595 583
rect 591 577 595 578
rect 663 582 667 583
rect 663 577 667 578
rect 695 582 699 583
rect 695 577 699 578
rect 775 582 779 583
rect 775 577 779 578
rect 807 582 811 583
rect 807 577 811 578
rect 895 582 899 583
rect 895 577 899 578
rect 919 582 923 583
rect 919 577 923 578
rect 112 562 114 577
rect 664 567 666 577
rect 776 567 778 577
rect 896 567 898 577
rect 662 566 668 567
rect 662 562 663 566
rect 667 562 668 566
rect 110 561 116 562
rect 662 561 668 562
rect 774 566 780 567
rect 774 562 775 566
rect 779 562 780 566
rect 774 561 780 562
rect 894 566 900 567
rect 894 562 895 566
rect 899 562 900 566
rect 894 561 900 562
rect 110 557 111 561
rect 115 557 116 561
rect 110 556 116 557
rect 110 544 116 545
rect 110 540 111 544
rect 115 540 116 544
rect 110 539 116 540
rect 112 495 114 539
rect 878 535 884 536
rect 878 531 879 535
rect 883 531 884 535
rect 878 530 884 531
rect 662 525 668 526
rect 662 521 663 525
rect 667 521 668 525
rect 662 520 668 521
rect 774 525 780 526
rect 774 521 775 525
rect 779 521 780 525
rect 774 520 780 521
rect 664 495 666 520
rect 776 495 778 520
rect 880 508 882 530
rect 894 525 900 526
rect 894 521 895 525
rect 899 521 900 525
rect 894 520 900 521
rect 878 507 884 508
rect 878 503 879 507
rect 883 503 884 507
rect 878 502 884 503
rect 896 495 898 520
rect 944 516 946 630
rect 1030 606 1036 607
rect 1030 602 1031 606
rect 1035 602 1036 606
rect 1030 601 1036 602
rect 1142 606 1148 607
rect 1142 602 1143 606
rect 1147 602 1148 606
rect 1142 601 1148 602
rect 1262 606 1268 607
rect 1262 602 1263 606
rect 1267 602 1268 606
rect 1262 601 1268 602
rect 1382 606 1388 607
rect 1382 602 1383 606
rect 1387 602 1388 606
rect 1382 601 1388 602
rect 1502 606 1508 607
rect 1502 602 1503 606
rect 1507 602 1508 606
rect 1502 601 1508 602
rect 1032 583 1034 601
rect 1144 583 1146 601
rect 1264 583 1266 601
rect 1384 583 1386 601
rect 1504 583 1506 601
rect 1023 582 1027 583
rect 1023 577 1027 578
rect 1031 582 1035 583
rect 1031 577 1035 578
rect 1143 582 1147 583
rect 1143 577 1147 578
rect 1159 582 1163 583
rect 1159 577 1163 578
rect 1263 582 1267 583
rect 1263 577 1267 578
rect 1303 582 1307 583
rect 1303 577 1307 578
rect 1383 582 1387 583
rect 1383 577 1387 578
rect 1447 582 1451 583
rect 1447 577 1451 578
rect 1503 582 1507 583
rect 1503 577 1507 578
rect 1024 567 1026 577
rect 1160 567 1162 577
rect 1304 567 1306 577
rect 1448 567 1450 577
rect 1022 566 1028 567
rect 1022 562 1023 566
rect 1027 562 1028 566
rect 1022 561 1028 562
rect 1158 566 1164 567
rect 1158 562 1159 566
rect 1163 562 1164 566
rect 1158 561 1164 562
rect 1302 566 1308 567
rect 1302 562 1303 566
rect 1307 562 1308 566
rect 1302 561 1308 562
rect 1446 566 1452 567
rect 1446 562 1447 566
rect 1451 562 1452 566
rect 1446 561 1452 562
rect 1568 536 1570 642
rect 2032 629 2034 657
rect 2064 656 2066 694
rect 2070 684 2076 685
rect 2070 680 2071 684
rect 2075 680 2076 684
rect 2070 679 2076 680
rect 2062 655 2068 656
rect 2062 651 2063 655
rect 2067 651 2068 655
rect 2062 650 2068 651
rect 2072 647 2074 679
rect 2464 676 2466 790
rect 2680 788 2682 797
rect 2952 788 2954 797
rect 3200 788 3202 797
rect 2678 787 2684 788
rect 2678 783 2679 787
rect 2683 783 2684 787
rect 2678 782 2684 783
rect 2950 787 2956 788
rect 2950 783 2951 787
rect 2955 783 2956 787
rect 2950 782 2956 783
rect 3198 787 3204 788
rect 3198 783 3199 787
rect 3203 783 3204 787
rect 3198 782 3204 783
rect 3272 780 3274 802
rect 3311 797 3315 798
rect 3439 802 3443 803
rect 3494 802 3500 803
rect 3511 802 3515 803
rect 3439 797 3443 798
rect 3511 797 3515 798
rect 3671 802 3675 803
rect 3694 802 3700 803
rect 3711 802 3715 803
rect 3671 797 3675 798
rect 3711 797 3715 798
rect 3895 802 3899 803
rect 3958 802 3964 803
rect 3895 797 3899 798
rect 3440 788 3442 797
rect 3672 788 3674 797
rect 3822 795 3828 796
rect 3822 791 3823 795
rect 3827 791 3828 795
rect 3822 790 3828 791
rect 3438 787 3444 788
rect 3438 783 3439 787
rect 3443 783 3444 787
rect 3438 782 3444 783
rect 3670 787 3676 788
rect 3670 783 3671 787
rect 3675 783 3676 787
rect 3670 782 3676 783
rect 3062 779 3068 780
rect 3062 775 3063 779
rect 3067 775 3068 779
rect 3062 774 3068 775
rect 3270 779 3276 780
rect 3270 775 3271 779
rect 3275 775 3276 779
rect 3270 774 3276 775
rect 2678 746 2684 747
rect 2678 742 2679 746
rect 2683 742 2684 746
rect 2678 741 2684 742
rect 2950 746 2956 747
rect 2950 742 2951 746
rect 2955 742 2956 746
rect 2950 741 2956 742
rect 2680 723 2682 741
rect 2952 723 2954 741
rect 2551 722 2555 723
rect 2551 717 2555 718
rect 2679 722 2683 723
rect 2679 717 2683 718
rect 2775 722 2779 723
rect 2775 717 2779 718
rect 2951 722 2955 723
rect 2951 717 2955 718
rect 2991 722 2995 723
rect 2991 717 2995 718
rect 2552 707 2554 717
rect 2776 707 2778 717
rect 2992 707 2994 717
rect 2550 706 2556 707
rect 2550 702 2551 706
rect 2555 702 2556 706
rect 2550 701 2556 702
rect 2774 706 2780 707
rect 2774 702 2775 706
rect 2779 702 2780 706
rect 2774 701 2780 702
rect 2990 706 2996 707
rect 2990 702 2991 706
rect 2995 702 2996 706
rect 2990 701 2996 702
rect 2182 675 2188 676
rect 2182 671 2183 675
rect 2187 671 2188 675
rect 2182 670 2188 671
rect 2462 675 2468 676
rect 2462 671 2463 675
rect 2467 671 2468 675
rect 2462 670 2468 671
rect 2110 665 2116 666
rect 2110 661 2111 665
rect 2115 661 2116 665
rect 2110 660 2116 661
rect 2112 647 2114 660
rect 2071 646 2075 647
rect 2071 641 2075 642
rect 2111 646 2115 647
rect 2111 641 2115 642
rect 2127 646 2131 647
rect 2127 641 2131 642
rect 2030 628 2036 629
rect 2030 624 2031 628
rect 2035 624 2036 628
rect 2030 623 2036 624
rect 2072 613 2074 641
rect 2128 632 2130 641
rect 2184 640 2186 670
rect 2326 665 2332 666
rect 2326 661 2327 665
rect 2331 661 2332 665
rect 2326 660 2332 661
rect 2550 665 2556 666
rect 2550 661 2551 665
rect 2555 661 2556 665
rect 2550 660 2556 661
rect 2774 665 2780 666
rect 2774 661 2775 665
rect 2779 661 2780 665
rect 2774 660 2780 661
rect 2990 665 2996 666
rect 2990 661 2991 665
rect 2995 661 2996 665
rect 2990 660 2996 661
rect 2328 647 2330 660
rect 2552 647 2554 660
rect 2722 647 2728 648
rect 2776 647 2778 660
rect 2992 647 2994 660
rect 3064 656 3066 774
rect 3198 746 3204 747
rect 3198 742 3199 746
rect 3203 742 3204 746
rect 3198 741 3204 742
rect 3438 746 3444 747
rect 3438 742 3439 746
rect 3443 742 3444 746
rect 3438 741 3444 742
rect 3670 746 3676 747
rect 3670 742 3671 746
rect 3675 742 3676 746
rect 3670 741 3676 742
rect 3200 723 3202 741
rect 3440 723 3442 741
rect 3672 723 3674 741
rect 3199 722 3203 723
rect 3199 717 3203 718
rect 3207 722 3211 723
rect 3207 717 3211 718
rect 3415 722 3419 723
rect 3415 717 3419 718
rect 3439 722 3443 723
rect 3439 717 3443 718
rect 3623 722 3627 723
rect 3623 717 3627 718
rect 3671 722 3675 723
rect 3671 717 3675 718
rect 3208 707 3210 717
rect 3416 707 3418 717
rect 3624 707 3626 717
rect 3206 706 3212 707
rect 3206 702 3207 706
rect 3211 702 3212 706
rect 3206 701 3212 702
rect 3414 706 3420 707
rect 3414 702 3415 706
rect 3419 702 3420 706
rect 3414 701 3420 702
rect 3622 706 3628 707
rect 3622 702 3623 706
rect 3627 702 3628 706
rect 3622 701 3628 702
rect 3824 676 3826 790
rect 3896 788 3898 797
rect 3968 796 3970 822
rect 3992 803 3994 831
rect 3991 802 3995 803
rect 3991 797 3995 798
rect 3966 795 3972 796
rect 3966 791 3967 795
rect 3971 791 3972 795
rect 3966 790 3972 791
rect 3894 787 3900 788
rect 3894 783 3895 787
rect 3899 783 3900 787
rect 3894 782 3900 783
rect 3918 775 3924 776
rect 3918 771 3919 775
rect 3923 771 3924 775
rect 3918 770 3924 771
rect 3894 746 3900 747
rect 3894 742 3895 746
rect 3899 742 3900 746
rect 3894 741 3900 742
rect 3896 723 3898 741
rect 3831 722 3835 723
rect 3831 717 3835 718
rect 3895 722 3899 723
rect 3895 717 3899 718
rect 3832 707 3834 717
rect 3830 706 3836 707
rect 3830 702 3831 706
rect 3835 702 3836 706
rect 3830 701 3836 702
rect 3190 675 3196 676
rect 3190 671 3191 675
rect 3195 671 3196 675
rect 3190 670 3196 671
rect 3198 675 3204 676
rect 3198 671 3199 675
rect 3203 671 3204 675
rect 3198 670 3204 671
rect 3546 675 3552 676
rect 3546 671 3547 675
rect 3551 671 3552 675
rect 3546 670 3552 671
rect 3822 675 3828 676
rect 3822 671 3823 675
rect 3827 671 3828 675
rect 3822 670 3828 671
rect 3192 656 3194 670
rect 3062 655 3068 656
rect 3062 651 3063 655
rect 3067 651 3068 655
rect 3062 650 3068 651
rect 3190 655 3196 656
rect 3190 651 3191 655
rect 3195 651 3196 655
rect 3190 650 3196 651
rect 3110 647 3116 648
rect 2295 646 2299 647
rect 2295 641 2299 642
rect 2327 646 2331 647
rect 2327 641 2331 642
rect 2455 646 2459 647
rect 2455 641 2459 642
rect 2551 646 2555 647
rect 2551 641 2555 642
rect 2615 646 2619 647
rect 2722 643 2723 647
rect 2727 643 2728 647
rect 2722 642 2728 643
rect 2775 646 2779 647
rect 2615 641 2619 642
rect 2182 639 2188 640
rect 2182 635 2183 639
rect 2187 635 2188 639
rect 2182 634 2188 635
rect 2296 632 2298 641
rect 2456 632 2458 641
rect 2616 632 2618 641
rect 2126 631 2132 632
rect 2126 627 2127 631
rect 2131 627 2132 631
rect 2126 626 2132 627
rect 2294 631 2300 632
rect 2294 627 2295 631
rect 2299 627 2300 631
rect 2294 626 2300 627
rect 2454 631 2460 632
rect 2454 627 2455 631
rect 2459 627 2460 631
rect 2454 626 2460 627
rect 2614 631 2620 632
rect 2614 627 2615 631
rect 2619 627 2620 631
rect 2614 626 2620 627
rect 2724 624 2726 642
rect 2775 641 2779 642
rect 2783 646 2787 647
rect 2783 641 2787 642
rect 2951 646 2955 647
rect 2951 641 2955 642
rect 2991 646 2995 647
rect 3110 643 3111 647
rect 3115 643 3116 647
rect 3110 642 3116 643
rect 3127 646 3131 647
rect 2991 641 2995 642
rect 2784 632 2786 641
rect 2870 639 2876 640
rect 2870 635 2871 639
rect 2875 635 2876 639
rect 2870 634 2876 635
rect 2782 631 2788 632
rect 2782 627 2783 631
rect 2787 627 2788 631
rect 2782 626 2788 627
rect 2518 623 2524 624
rect 2518 619 2519 623
rect 2523 619 2524 623
rect 2518 618 2524 619
rect 2722 623 2728 624
rect 2722 619 2723 623
rect 2727 619 2728 623
rect 2722 618 2728 619
rect 2070 612 2076 613
rect 2030 611 2036 612
rect 2030 607 2031 611
rect 2035 607 2036 611
rect 2070 608 2071 612
rect 2075 608 2076 612
rect 2070 607 2076 608
rect 1622 606 1628 607
rect 2030 606 2036 607
rect 1622 602 1623 606
rect 1627 602 1628 606
rect 1622 601 1628 602
rect 1624 583 1626 601
rect 2032 583 2034 606
rect 2070 595 2076 596
rect 2070 591 2071 595
rect 2075 591 2076 595
rect 2070 590 2076 591
rect 2126 590 2132 591
rect 1591 582 1595 583
rect 1591 577 1595 578
rect 1623 582 1627 583
rect 1623 577 1627 578
rect 1735 582 1739 583
rect 1735 577 1739 578
rect 1879 582 1883 583
rect 1879 577 1883 578
rect 2031 582 2035 583
rect 2031 577 2035 578
rect 1592 567 1594 577
rect 1736 567 1738 577
rect 1880 567 1882 577
rect 1590 566 1596 567
rect 1590 562 1591 566
rect 1595 562 1596 566
rect 1590 561 1596 562
rect 1734 566 1740 567
rect 1734 562 1735 566
rect 1739 562 1740 566
rect 1734 561 1740 562
rect 1878 566 1884 567
rect 1878 562 1879 566
rect 1883 562 1884 566
rect 2032 562 2034 577
rect 2072 567 2074 590
rect 2126 586 2127 590
rect 2131 586 2132 590
rect 2126 585 2132 586
rect 2294 590 2300 591
rect 2294 586 2295 590
rect 2299 586 2300 590
rect 2294 585 2300 586
rect 2454 590 2460 591
rect 2454 586 2455 590
rect 2459 586 2460 590
rect 2454 585 2460 586
rect 2128 567 2130 585
rect 2296 567 2298 585
rect 2456 567 2458 585
rect 2071 566 2075 567
rect 1878 561 1884 562
rect 2030 561 2036 562
rect 2071 561 2075 562
rect 2127 566 2131 567
rect 2127 561 2131 562
rect 2295 566 2299 567
rect 2295 561 2299 562
rect 2303 566 2307 567
rect 2303 561 2307 562
rect 2447 566 2451 567
rect 2447 561 2451 562
rect 2455 566 2459 567
rect 2455 561 2459 562
rect 2030 557 2031 561
rect 2035 557 2036 561
rect 2030 556 2036 557
rect 2072 546 2074 561
rect 2304 551 2306 561
rect 2448 551 2450 561
rect 2302 550 2308 551
rect 2302 546 2303 550
rect 2307 546 2308 550
rect 2070 545 2076 546
rect 2302 545 2308 546
rect 2446 550 2452 551
rect 2446 546 2447 550
rect 2451 546 2452 550
rect 2446 545 2452 546
rect 2030 544 2036 545
rect 2030 540 2031 544
rect 2035 540 2036 544
rect 2070 541 2071 545
rect 2075 541 2076 545
rect 2070 540 2076 541
rect 2030 539 2036 540
rect 1266 535 1272 536
rect 1266 531 1267 535
rect 1271 531 1272 535
rect 1266 530 1272 531
rect 1326 535 1332 536
rect 1326 531 1327 535
rect 1331 531 1332 535
rect 1326 530 1332 531
rect 1566 535 1572 536
rect 1566 531 1567 535
rect 1571 531 1572 535
rect 1566 530 1572 531
rect 1022 525 1028 526
rect 1022 521 1023 525
rect 1027 521 1028 525
rect 1022 520 1028 521
rect 1158 525 1164 526
rect 1158 521 1159 525
rect 1163 521 1164 525
rect 1158 520 1164 521
rect 942 515 948 516
rect 942 511 943 515
rect 947 511 948 515
rect 942 510 948 511
rect 1024 495 1026 520
rect 1160 495 1162 520
rect 1268 516 1270 530
rect 1302 525 1308 526
rect 1302 521 1303 525
rect 1307 521 1308 525
rect 1302 520 1308 521
rect 1266 515 1272 516
rect 1266 511 1267 515
rect 1271 511 1272 515
rect 1266 510 1272 511
rect 1304 495 1306 520
rect 111 494 115 495
rect 111 489 115 490
rect 535 494 539 495
rect 535 489 539 490
rect 639 494 643 495
rect 639 489 643 490
rect 663 494 667 495
rect 663 489 667 490
rect 743 494 747 495
rect 743 489 747 490
rect 775 494 779 495
rect 775 489 779 490
rect 847 494 851 495
rect 847 489 851 490
rect 895 494 899 495
rect 895 489 899 490
rect 967 494 971 495
rect 967 489 971 490
rect 1023 494 1027 495
rect 1023 489 1027 490
rect 1103 494 1107 495
rect 1103 489 1107 490
rect 1159 494 1163 495
rect 1159 489 1163 490
rect 1255 494 1259 495
rect 1255 489 1259 490
rect 1303 494 1307 495
rect 1303 489 1307 490
rect 112 461 114 489
rect 536 480 538 489
rect 640 480 642 489
rect 744 480 746 489
rect 848 480 850 489
rect 968 480 970 489
rect 1038 487 1044 488
rect 1038 483 1039 487
rect 1043 483 1044 487
rect 1038 482 1044 483
rect 534 479 540 480
rect 534 475 535 479
rect 539 475 540 479
rect 534 474 540 475
rect 638 479 644 480
rect 638 475 639 479
rect 643 475 644 479
rect 638 474 644 475
rect 742 479 748 480
rect 742 475 743 479
rect 747 475 748 479
rect 742 474 748 475
rect 846 479 852 480
rect 846 475 847 479
rect 851 475 852 479
rect 846 474 852 475
rect 966 479 972 480
rect 966 475 967 479
rect 971 475 972 479
rect 966 474 972 475
rect 558 467 564 468
rect 558 463 559 467
rect 563 463 564 467
rect 558 462 564 463
rect 110 460 116 461
rect 110 456 111 460
rect 115 456 116 460
rect 110 455 116 456
rect 110 443 116 444
rect 110 439 111 443
rect 115 439 116 443
rect 110 438 116 439
rect 534 438 540 439
rect 112 419 114 438
rect 534 434 535 438
rect 539 434 540 438
rect 534 433 540 434
rect 536 419 538 433
rect 111 418 115 419
rect 111 413 115 414
rect 495 418 499 419
rect 495 413 499 414
rect 535 418 539 419
rect 535 413 539 414
rect 112 398 114 413
rect 496 403 498 413
rect 494 402 500 403
rect 494 398 495 402
rect 499 398 500 402
rect 110 397 116 398
rect 494 397 500 398
rect 110 393 111 397
rect 115 393 116 397
rect 110 392 116 393
rect 110 380 116 381
rect 110 376 111 380
rect 115 376 116 380
rect 110 375 116 376
rect 112 335 114 375
rect 494 361 500 362
rect 494 357 495 361
rect 499 357 500 361
rect 494 356 500 357
rect 446 335 452 336
rect 496 335 498 356
rect 560 352 562 462
rect 638 438 644 439
rect 638 434 639 438
rect 643 434 644 438
rect 638 433 644 434
rect 742 438 748 439
rect 742 434 743 438
rect 747 434 748 438
rect 742 433 748 434
rect 846 438 852 439
rect 846 434 847 438
rect 851 434 852 438
rect 846 433 852 434
rect 966 438 972 439
rect 966 434 967 438
rect 971 434 972 438
rect 966 433 972 434
rect 640 419 642 433
rect 744 419 746 433
rect 848 419 850 433
rect 968 419 970 433
rect 631 418 635 419
rect 631 413 635 414
rect 639 418 643 419
rect 639 413 643 414
rect 743 418 747 419
rect 743 413 747 414
rect 767 418 771 419
rect 767 413 771 414
rect 847 418 851 419
rect 847 413 851 414
rect 911 418 915 419
rect 911 413 915 414
rect 967 418 971 419
rect 967 413 971 414
rect 632 403 634 413
rect 768 403 770 413
rect 912 403 914 413
rect 630 402 636 403
rect 630 398 631 402
rect 635 398 636 402
rect 630 397 636 398
rect 766 402 772 403
rect 766 398 767 402
rect 771 398 772 402
rect 766 397 772 398
rect 910 402 916 403
rect 910 398 911 402
rect 915 398 916 402
rect 910 397 916 398
rect 1040 372 1042 482
rect 1104 480 1106 489
rect 1256 480 1258 489
rect 1328 488 1330 530
rect 1446 525 1452 526
rect 1446 521 1447 525
rect 1451 521 1452 525
rect 1446 520 1452 521
rect 1590 525 1596 526
rect 1590 521 1591 525
rect 1595 521 1596 525
rect 1590 520 1596 521
rect 1734 525 1740 526
rect 1734 521 1735 525
rect 1739 521 1740 525
rect 1734 520 1740 521
rect 1878 525 1884 526
rect 1878 521 1879 525
rect 1883 521 1884 525
rect 1878 520 1884 521
rect 1448 495 1450 520
rect 1592 495 1594 520
rect 1736 495 1738 520
rect 1880 495 1882 520
rect 1950 515 1956 516
rect 1950 511 1951 515
rect 1955 511 1956 515
rect 1950 510 1956 511
rect 1415 494 1419 495
rect 1415 489 1419 490
rect 1447 494 1451 495
rect 1447 489 1451 490
rect 1591 494 1595 495
rect 1591 489 1595 490
rect 1735 494 1739 495
rect 1735 489 1739 490
rect 1775 494 1779 495
rect 1775 489 1779 490
rect 1879 494 1883 495
rect 1879 489 1883 490
rect 1935 494 1939 495
rect 1935 489 1939 490
rect 1326 487 1332 488
rect 1326 483 1327 487
rect 1331 483 1332 487
rect 1326 482 1332 483
rect 1416 480 1418 489
rect 1592 480 1594 489
rect 1598 487 1604 488
rect 1598 483 1599 487
rect 1603 483 1604 487
rect 1598 482 1604 483
rect 1102 479 1108 480
rect 1102 475 1103 479
rect 1107 475 1108 479
rect 1254 479 1260 480
rect 1102 474 1108 475
rect 1239 476 1243 477
rect 1254 475 1255 479
rect 1259 475 1260 479
rect 1254 474 1260 475
rect 1414 479 1420 480
rect 1414 475 1415 479
rect 1419 475 1420 479
rect 1414 474 1420 475
rect 1590 479 1596 480
rect 1590 475 1591 479
rect 1595 475 1596 479
rect 1600 477 1602 482
rect 1776 480 1778 489
rect 1846 487 1852 488
rect 1846 483 1847 487
rect 1851 483 1852 487
rect 1846 482 1852 483
rect 1774 479 1780 480
rect 1590 474 1596 475
rect 1599 476 1603 477
rect 1774 475 1775 479
rect 1779 475 1780 479
rect 1774 474 1780 475
rect 1238 471 1244 472
rect 1599 471 1603 472
rect 1238 467 1239 471
rect 1243 467 1244 471
rect 1238 466 1244 467
rect 1406 467 1412 468
rect 1406 463 1407 467
rect 1411 463 1412 467
rect 1406 462 1412 463
rect 1102 438 1108 439
rect 1102 434 1103 438
rect 1107 434 1108 438
rect 1102 433 1108 434
rect 1254 438 1260 439
rect 1254 434 1255 438
rect 1259 434 1260 438
rect 1254 433 1260 434
rect 1104 419 1106 433
rect 1256 419 1258 433
rect 1047 418 1051 419
rect 1047 413 1051 414
rect 1103 418 1107 419
rect 1103 413 1107 414
rect 1183 418 1187 419
rect 1183 413 1187 414
rect 1255 418 1259 419
rect 1255 413 1259 414
rect 1319 418 1323 419
rect 1319 413 1323 414
rect 1048 403 1050 413
rect 1184 403 1186 413
rect 1320 403 1322 413
rect 1046 402 1052 403
rect 1046 398 1047 402
rect 1051 398 1052 402
rect 1046 397 1052 398
rect 1182 402 1188 403
rect 1182 398 1183 402
rect 1187 398 1188 402
rect 1182 397 1188 398
rect 1318 402 1324 403
rect 1318 398 1319 402
rect 1323 398 1324 402
rect 1318 397 1324 398
rect 614 371 620 372
rect 614 367 615 371
rect 619 367 620 371
rect 614 366 620 367
rect 750 371 756 372
rect 750 367 751 371
rect 755 367 756 371
rect 750 366 756 367
rect 838 371 844 372
rect 838 367 839 371
rect 843 367 844 371
rect 838 366 844 367
rect 1030 371 1036 372
rect 1030 367 1031 371
rect 1035 367 1036 371
rect 1030 366 1036 367
rect 1038 371 1044 372
rect 1038 367 1039 371
rect 1043 367 1044 371
rect 1038 366 1044 367
rect 1302 371 1308 372
rect 1302 367 1303 371
rect 1307 367 1308 371
rect 1302 366 1308 367
rect 616 352 618 366
rect 630 361 636 362
rect 630 357 631 361
rect 635 357 636 361
rect 630 356 636 357
rect 558 351 564 352
rect 558 347 559 351
rect 563 347 564 351
rect 558 346 564 347
rect 614 351 620 352
rect 614 347 615 351
rect 619 347 620 351
rect 614 346 620 347
rect 632 335 634 356
rect 752 352 754 366
rect 766 361 772 362
rect 766 357 767 361
rect 771 357 772 361
rect 766 356 772 357
rect 750 351 756 352
rect 750 347 751 351
rect 755 347 756 351
rect 750 346 756 347
rect 768 335 770 356
rect 111 334 115 335
rect 111 329 115 330
rect 335 334 339 335
rect 446 331 447 335
rect 451 331 452 335
rect 446 330 452 331
rect 463 334 467 335
rect 335 329 339 330
rect 112 301 114 329
rect 336 320 338 329
rect 334 319 340 320
rect 334 315 335 319
rect 339 315 340 319
rect 334 314 340 315
rect 448 312 450 330
rect 463 329 467 330
rect 495 334 499 335
rect 495 329 499 330
rect 607 334 611 335
rect 607 329 611 330
rect 631 334 635 335
rect 631 329 635 330
rect 767 334 771 335
rect 767 329 771 330
rect 464 320 466 329
rect 608 320 610 329
rect 768 320 770 329
rect 840 328 842 366
rect 910 361 916 362
rect 910 357 911 361
rect 915 357 916 361
rect 910 356 916 357
rect 854 335 860 336
rect 912 335 914 356
rect 1032 352 1034 366
rect 1046 361 1052 362
rect 1046 357 1047 361
rect 1051 357 1052 361
rect 1046 356 1052 357
rect 1182 361 1188 362
rect 1182 357 1183 361
rect 1187 357 1188 361
rect 1182 356 1188 357
rect 966 351 972 352
rect 966 347 967 351
rect 971 347 972 351
rect 966 346 972 347
rect 1030 351 1036 352
rect 1030 347 1031 351
rect 1035 347 1036 351
rect 1030 346 1036 347
rect 854 331 855 335
rect 859 331 860 335
rect 854 330 860 331
rect 911 334 915 335
rect 838 327 844 328
rect 838 323 839 327
rect 843 323 844 327
rect 838 322 844 323
rect 462 319 468 320
rect 462 315 463 319
rect 467 315 468 319
rect 462 314 468 315
rect 606 319 612 320
rect 606 315 607 319
rect 611 315 612 319
rect 606 314 612 315
rect 766 319 772 320
rect 766 315 767 319
rect 771 315 772 319
rect 766 314 772 315
rect 446 311 452 312
rect 446 307 447 311
rect 451 307 452 311
rect 446 306 452 307
rect 110 300 116 301
rect 110 296 111 300
rect 115 296 116 300
rect 110 295 116 296
rect 110 283 116 284
rect 110 279 111 283
rect 115 279 116 283
rect 110 278 116 279
rect 334 278 340 279
rect 112 255 114 278
rect 334 274 335 278
rect 339 274 340 278
rect 334 273 340 274
rect 462 278 468 279
rect 462 274 463 278
rect 467 274 468 278
rect 462 273 468 274
rect 606 278 612 279
rect 606 274 607 278
rect 611 274 612 278
rect 606 273 612 274
rect 766 278 772 279
rect 766 274 767 278
rect 771 274 772 278
rect 766 273 772 274
rect 336 255 338 273
rect 464 255 466 273
rect 608 255 610 273
rect 768 255 770 273
rect 111 254 115 255
rect 111 249 115 250
rect 151 254 155 255
rect 151 249 155 250
rect 279 254 283 255
rect 279 249 283 250
rect 335 254 339 255
rect 335 249 339 250
rect 431 254 435 255
rect 431 249 435 250
rect 463 254 467 255
rect 463 249 467 250
rect 599 254 603 255
rect 599 249 603 250
rect 607 254 611 255
rect 607 249 611 250
rect 767 254 771 255
rect 767 249 771 250
rect 783 254 787 255
rect 783 249 787 250
rect 112 234 114 249
rect 152 239 154 249
rect 280 239 282 249
rect 432 239 434 249
rect 600 239 602 249
rect 784 239 786 249
rect 150 238 156 239
rect 150 234 151 238
rect 155 234 156 238
rect 110 233 116 234
rect 150 233 156 234
rect 278 238 284 239
rect 278 234 279 238
rect 283 234 284 238
rect 278 233 284 234
rect 430 238 436 239
rect 430 234 431 238
rect 435 234 436 238
rect 430 233 436 234
rect 598 238 604 239
rect 598 234 599 238
rect 603 234 604 238
rect 598 233 604 234
rect 782 238 788 239
rect 782 234 783 238
rect 787 234 788 238
rect 782 233 788 234
rect 110 229 111 233
rect 115 229 116 233
rect 110 228 116 229
rect 110 216 116 217
rect 110 212 111 216
rect 115 212 116 216
rect 110 211 116 212
rect 112 159 114 211
rect 230 207 236 208
rect 230 203 231 207
rect 235 203 236 207
rect 230 202 236 203
rect 150 197 156 198
rect 150 193 151 197
rect 155 193 156 197
rect 150 192 156 193
rect 152 159 154 192
rect 232 160 234 202
rect 278 197 284 198
rect 278 193 279 197
rect 283 193 284 197
rect 278 192 284 193
rect 430 197 436 198
rect 430 193 431 197
rect 435 193 436 197
rect 430 192 436 193
rect 598 197 604 198
rect 598 193 599 197
rect 603 193 604 197
rect 598 192 604 193
rect 782 197 788 198
rect 782 193 783 197
rect 787 193 788 197
rect 782 192 788 193
rect 230 159 236 160
rect 280 159 282 192
rect 432 159 434 192
rect 600 159 602 192
rect 784 159 786 192
rect 856 188 858 330
rect 911 329 915 330
rect 943 334 947 335
rect 943 329 947 330
rect 944 320 946 329
rect 942 319 948 320
rect 942 315 943 319
rect 947 315 948 319
rect 942 314 948 315
rect 968 308 970 346
rect 1048 335 1050 356
rect 1184 335 1186 356
rect 1304 344 1306 366
rect 1318 361 1324 362
rect 1318 357 1319 361
rect 1323 357 1324 361
rect 1318 356 1324 357
rect 1302 343 1308 344
rect 1302 339 1303 343
rect 1307 339 1308 343
rect 1302 338 1308 339
rect 1320 335 1322 356
rect 1408 352 1410 462
rect 1414 438 1420 439
rect 1414 434 1415 438
rect 1419 434 1420 438
rect 1414 433 1420 434
rect 1590 438 1596 439
rect 1590 434 1591 438
rect 1595 434 1596 438
rect 1590 433 1596 434
rect 1774 438 1780 439
rect 1774 434 1775 438
rect 1779 434 1780 438
rect 1774 433 1780 434
rect 1416 419 1418 433
rect 1592 419 1594 433
rect 1776 419 1778 433
rect 1415 418 1419 419
rect 1415 413 1419 414
rect 1447 418 1451 419
rect 1447 413 1451 414
rect 1575 418 1579 419
rect 1575 413 1579 414
rect 1591 418 1595 419
rect 1591 413 1595 414
rect 1703 418 1707 419
rect 1703 413 1707 414
rect 1775 418 1779 419
rect 1775 413 1779 414
rect 1831 418 1835 419
rect 1831 413 1835 414
rect 1448 403 1450 413
rect 1576 403 1578 413
rect 1704 403 1706 413
rect 1832 403 1834 413
rect 1446 402 1452 403
rect 1446 398 1447 402
rect 1451 398 1452 402
rect 1446 397 1452 398
rect 1574 402 1580 403
rect 1574 398 1575 402
rect 1579 398 1580 402
rect 1574 397 1580 398
rect 1702 402 1708 403
rect 1702 398 1703 402
rect 1707 398 1708 402
rect 1702 397 1708 398
rect 1830 402 1836 403
rect 1830 398 1831 402
rect 1835 398 1836 402
rect 1830 397 1836 398
rect 1848 372 1850 482
rect 1936 480 1938 489
rect 1934 479 1940 480
rect 1934 475 1935 479
rect 1939 475 1940 479
rect 1934 474 1940 475
rect 1952 468 1954 510
rect 2032 495 2034 539
rect 2070 528 2076 529
rect 2070 524 2071 528
rect 2075 524 2076 528
rect 2070 523 2076 524
rect 2031 494 2035 495
rect 2031 489 2035 490
rect 1950 467 1956 468
rect 1950 463 1951 467
rect 1955 463 1956 467
rect 1950 462 1956 463
rect 2032 461 2034 489
rect 2072 487 2074 523
rect 2430 519 2436 520
rect 2430 515 2431 519
rect 2435 515 2436 519
rect 2430 514 2436 515
rect 2302 509 2308 510
rect 2302 505 2303 509
rect 2307 505 2308 509
rect 2302 504 2308 505
rect 2304 487 2306 504
rect 2432 492 2434 514
rect 2446 509 2452 510
rect 2446 505 2447 509
rect 2451 505 2452 509
rect 2446 504 2452 505
rect 2430 491 2436 492
rect 2430 487 2431 491
rect 2435 487 2436 491
rect 2448 487 2450 504
rect 2520 500 2522 618
rect 2614 590 2620 591
rect 2614 586 2615 590
rect 2619 586 2620 590
rect 2614 585 2620 586
rect 2782 590 2788 591
rect 2782 586 2783 590
rect 2787 586 2788 590
rect 2782 585 2788 586
rect 2616 567 2618 585
rect 2784 567 2786 585
rect 2591 566 2595 567
rect 2591 561 2595 562
rect 2615 566 2619 567
rect 2615 561 2619 562
rect 2735 566 2739 567
rect 2735 561 2739 562
rect 2783 566 2787 567
rect 2783 561 2787 562
rect 2592 551 2594 561
rect 2736 551 2738 561
rect 2590 550 2596 551
rect 2590 546 2591 550
rect 2595 546 2596 550
rect 2590 545 2596 546
rect 2734 550 2740 551
rect 2734 546 2735 550
rect 2739 546 2740 550
rect 2734 545 2740 546
rect 2872 520 2874 634
rect 2952 632 2954 641
rect 2950 631 2956 632
rect 2950 627 2951 631
rect 2955 627 2956 631
rect 2950 626 2956 627
rect 3112 624 3114 642
rect 3127 641 3131 642
rect 3128 632 3130 641
rect 3200 640 3202 670
rect 3206 665 3212 666
rect 3206 661 3207 665
rect 3211 661 3212 665
rect 3206 660 3212 661
rect 3414 665 3420 666
rect 3414 661 3415 665
rect 3419 661 3420 665
rect 3414 660 3420 661
rect 3208 647 3210 660
rect 3416 647 3418 660
rect 3548 648 3550 670
rect 3622 665 3628 666
rect 3622 661 3623 665
rect 3627 661 3628 665
rect 3622 660 3628 661
rect 3830 665 3836 666
rect 3830 661 3831 665
rect 3835 661 3836 665
rect 3830 660 3836 661
rect 3546 647 3552 648
rect 3624 647 3626 660
rect 3694 655 3700 656
rect 3694 651 3695 655
rect 3699 651 3700 655
rect 3694 650 3700 651
rect 3207 646 3211 647
rect 3207 641 3211 642
rect 3303 646 3307 647
rect 3303 641 3307 642
rect 3415 646 3419 647
rect 3415 641 3419 642
rect 3487 646 3491 647
rect 3546 643 3547 647
rect 3551 643 3552 647
rect 3546 642 3552 643
rect 3623 646 3627 647
rect 3487 641 3491 642
rect 3623 641 3627 642
rect 3679 646 3683 647
rect 3679 641 3683 642
rect 3198 639 3204 640
rect 3198 635 3199 639
rect 3203 635 3204 639
rect 3198 634 3204 635
rect 3304 632 3306 641
rect 3488 632 3490 641
rect 3680 632 3682 641
rect 3126 631 3132 632
rect 3126 627 3127 631
rect 3131 627 3132 631
rect 3126 626 3132 627
rect 3302 631 3308 632
rect 3302 627 3303 631
rect 3307 627 3308 631
rect 3302 626 3308 627
rect 3486 631 3492 632
rect 3486 627 3487 631
rect 3491 627 3492 631
rect 3486 626 3492 627
rect 3678 631 3684 632
rect 3678 627 3679 631
rect 3683 627 3684 631
rect 3678 626 3684 627
rect 3110 623 3116 624
rect 3110 619 3111 623
rect 3115 619 3116 623
rect 3696 620 3698 650
rect 3832 647 3834 660
rect 3831 646 3835 647
rect 3831 641 3835 642
rect 3879 646 3883 647
rect 3920 644 3922 770
rect 3992 769 3994 797
rect 3990 768 3996 769
rect 3990 764 3991 768
rect 3995 764 3996 768
rect 3990 763 3996 764
rect 3990 751 3996 752
rect 3990 747 3991 751
rect 3995 747 3996 751
rect 3990 746 3996 747
rect 3992 723 3994 746
rect 3991 722 3995 723
rect 3991 717 3995 718
rect 3992 702 3994 717
rect 3990 701 3996 702
rect 3990 697 3991 701
rect 3995 697 3996 701
rect 3990 696 3996 697
rect 3990 684 3996 685
rect 3990 680 3991 684
rect 3995 680 3996 684
rect 3990 679 3996 680
rect 3992 647 3994 679
rect 3991 646 3995 647
rect 3879 641 3883 642
rect 3918 643 3924 644
rect 3814 639 3820 640
rect 3814 635 3815 639
rect 3819 635 3820 639
rect 3814 634 3820 635
rect 3110 618 3116 619
rect 3478 619 3484 620
rect 3478 615 3479 619
rect 3483 615 3484 619
rect 3478 614 3484 615
rect 3694 619 3700 620
rect 3694 615 3695 619
rect 3699 615 3700 619
rect 3694 614 3700 615
rect 2950 590 2956 591
rect 2950 586 2951 590
rect 2955 586 2956 590
rect 2950 585 2956 586
rect 3126 590 3132 591
rect 3126 586 3127 590
rect 3131 586 3132 590
rect 3126 585 3132 586
rect 3302 590 3308 591
rect 3302 586 3303 590
rect 3307 586 3308 590
rect 3302 585 3308 586
rect 2952 567 2954 585
rect 3128 567 3130 585
rect 3304 567 3306 585
rect 2879 566 2883 567
rect 2879 561 2883 562
rect 2951 566 2955 567
rect 2951 561 2955 562
rect 3031 566 3035 567
rect 3031 561 3035 562
rect 3127 566 3131 567
rect 3127 561 3131 562
rect 3183 566 3187 567
rect 3183 561 3187 562
rect 3303 566 3307 567
rect 3303 561 3307 562
rect 3335 566 3339 567
rect 3335 561 3339 562
rect 2880 551 2882 561
rect 3032 551 3034 561
rect 3184 551 3186 561
rect 3336 551 3338 561
rect 2878 550 2884 551
rect 2878 546 2879 550
rect 2883 546 2884 550
rect 2878 545 2884 546
rect 3030 550 3036 551
rect 3030 546 3031 550
rect 3035 546 3036 550
rect 3030 545 3036 546
rect 3182 550 3188 551
rect 3182 546 3183 550
rect 3187 546 3188 550
rect 3182 545 3188 546
rect 3334 550 3340 551
rect 3334 546 3335 550
rect 3339 546 3340 550
rect 3334 545 3340 546
rect 2718 519 2724 520
rect 2718 515 2719 519
rect 2723 515 2724 519
rect 2718 514 2724 515
rect 2806 519 2812 520
rect 2806 515 2807 519
rect 2811 515 2812 519
rect 2806 514 2812 515
rect 2870 519 2876 520
rect 2870 515 2871 519
rect 2875 515 2876 519
rect 2870 514 2876 515
rect 3166 519 3172 520
rect 3166 515 3167 519
rect 3171 515 3172 519
rect 3166 514 3172 515
rect 2590 509 2596 510
rect 2590 505 2591 509
rect 2595 505 2596 509
rect 2590 504 2596 505
rect 2518 499 2524 500
rect 2518 495 2519 499
rect 2523 495 2524 499
rect 2518 494 2524 495
rect 2592 487 2594 504
rect 2720 500 2722 514
rect 2734 509 2740 510
rect 2734 505 2735 509
rect 2739 505 2740 509
rect 2734 504 2740 505
rect 2718 499 2724 500
rect 2718 495 2719 499
rect 2723 495 2724 499
rect 2718 494 2724 495
rect 2598 487 2604 488
rect 2736 487 2738 504
rect 2071 486 2075 487
rect 2071 481 2075 482
rect 2303 486 2307 487
rect 2430 486 2436 487
rect 2447 486 2451 487
rect 2303 481 2307 482
rect 2447 481 2451 482
rect 2511 486 2515 487
rect 2511 481 2515 482
rect 2591 486 2595 487
rect 2598 483 2599 487
rect 2603 483 2604 487
rect 2598 482 2604 483
rect 2615 486 2619 487
rect 2591 481 2595 482
rect 2030 460 2036 461
rect 2030 456 2031 460
rect 2035 456 2036 460
rect 2030 455 2036 456
rect 2072 453 2074 481
rect 2512 472 2514 481
rect 2510 471 2516 472
rect 2510 467 2511 471
rect 2515 467 2516 471
rect 2510 466 2516 467
rect 2600 464 2602 482
rect 2615 481 2619 482
rect 2735 486 2739 487
rect 2735 481 2739 482
rect 2616 472 2618 481
rect 2736 472 2738 481
rect 2808 480 2810 514
rect 2878 509 2884 510
rect 2878 505 2879 509
rect 2883 505 2884 509
rect 2878 504 2884 505
rect 3030 509 3036 510
rect 3168 509 3170 514
rect 3182 509 3188 510
rect 3030 505 3031 509
rect 3035 505 3036 509
rect 3030 504 3036 505
rect 3167 508 3171 509
rect 3182 505 3183 509
rect 3187 505 3188 509
rect 3182 504 3188 505
rect 3334 509 3340 510
rect 3334 505 3335 509
rect 3339 505 3340 509
rect 3334 504 3340 505
rect 2880 487 2882 504
rect 2954 499 2960 500
rect 2954 495 2955 499
rect 2959 495 2960 499
rect 2954 494 2960 495
rect 2863 486 2867 487
rect 2863 481 2867 482
rect 2879 486 2883 487
rect 2879 481 2883 482
rect 2806 479 2812 480
rect 2806 475 2807 479
rect 2811 475 2812 479
rect 2806 474 2812 475
rect 2864 472 2866 481
rect 2956 480 2958 494
rect 3032 487 3034 504
rect 3167 503 3171 504
rect 3184 487 3186 504
rect 3336 487 3338 504
rect 3480 500 3482 614
rect 3486 590 3492 591
rect 3486 586 3487 590
rect 3491 586 3492 590
rect 3486 585 3492 586
rect 3678 590 3684 591
rect 3678 586 3679 590
rect 3683 586 3684 590
rect 3678 585 3684 586
rect 3488 567 3490 585
rect 3680 567 3682 585
rect 3487 566 3491 567
rect 3487 561 3491 562
rect 3495 566 3499 567
rect 3495 561 3499 562
rect 3655 566 3659 567
rect 3655 561 3659 562
rect 3679 566 3683 567
rect 3679 561 3683 562
rect 3496 551 3498 561
rect 3656 551 3658 561
rect 3494 550 3500 551
rect 3494 546 3495 550
rect 3499 546 3500 550
rect 3494 545 3500 546
rect 3654 550 3660 551
rect 3654 546 3655 550
rect 3659 546 3660 550
rect 3654 545 3660 546
rect 3816 520 3818 634
rect 3880 632 3882 641
rect 3918 639 3919 643
rect 3923 639 3924 643
rect 3991 641 3995 642
rect 3918 638 3924 639
rect 3878 631 3884 632
rect 3878 627 3879 631
rect 3883 627 3884 631
rect 3878 626 3884 627
rect 3894 619 3900 620
rect 3894 615 3895 619
rect 3899 615 3900 619
rect 3894 614 3900 615
rect 3878 590 3884 591
rect 3878 586 3879 590
rect 3883 586 3884 590
rect 3878 585 3884 586
rect 3880 567 3882 585
rect 3823 566 3827 567
rect 3823 561 3827 562
rect 3879 566 3883 567
rect 3879 561 3883 562
rect 3824 551 3826 561
rect 3822 550 3828 551
rect 3822 546 3823 550
rect 3827 546 3828 550
rect 3822 545 3828 546
rect 3814 519 3820 520
rect 3718 515 3724 516
rect 3718 511 3719 515
rect 3723 511 3724 515
rect 3814 515 3815 519
rect 3819 515 3820 519
rect 3814 514 3820 515
rect 3718 510 3724 511
rect 3494 509 3500 510
rect 3654 509 3660 510
rect 3494 505 3495 509
rect 3499 505 3500 509
rect 3494 504 3500 505
rect 3567 508 3571 509
rect 3654 505 3655 509
rect 3659 505 3660 509
rect 3654 504 3660 505
rect 3478 499 3484 500
rect 3478 495 3479 499
rect 3483 495 3484 499
rect 3478 494 3484 495
rect 3496 487 3498 504
rect 3567 503 3571 504
rect 3568 500 3570 503
rect 3566 499 3572 500
rect 3566 495 3567 499
rect 3571 495 3572 499
rect 3566 494 3572 495
rect 3656 487 3658 504
rect 3007 486 3011 487
rect 3007 481 3011 482
rect 3031 486 3035 487
rect 3031 481 3035 482
rect 3159 486 3163 487
rect 3159 481 3163 482
rect 3183 486 3187 487
rect 3183 481 3187 482
rect 3319 486 3323 487
rect 3319 481 3323 482
rect 3335 486 3339 487
rect 3335 481 3339 482
rect 3479 486 3483 487
rect 3479 481 3483 482
rect 3495 486 3499 487
rect 3495 481 3499 482
rect 3647 486 3651 487
rect 3647 481 3651 482
rect 3655 486 3659 487
rect 3655 481 3659 482
rect 2954 479 2960 480
rect 2954 475 2955 479
rect 2959 475 2960 479
rect 2954 474 2960 475
rect 3008 472 3010 481
rect 3160 472 3162 481
rect 3320 472 3322 481
rect 3390 479 3396 480
rect 3390 475 3391 479
rect 3395 475 3396 479
rect 3390 474 3396 475
rect 2614 471 2620 472
rect 2614 467 2615 471
rect 2619 467 2620 471
rect 2614 466 2620 467
rect 2734 471 2740 472
rect 2734 467 2735 471
rect 2739 467 2740 471
rect 2734 466 2740 467
rect 2862 471 2868 472
rect 2862 467 2863 471
rect 2867 467 2868 471
rect 2862 466 2868 467
rect 3006 471 3012 472
rect 3006 467 3007 471
rect 3011 467 3012 471
rect 3006 466 3012 467
rect 3158 471 3164 472
rect 3158 467 3159 471
rect 3163 467 3164 471
rect 3158 466 3164 467
rect 3318 471 3324 472
rect 3318 467 3319 471
rect 3323 467 3324 471
rect 3318 466 3324 467
rect 2598 463 2604 464
rect 2598 459 2599 463
rect 2603 459 2604 463
rect 2598 458 2604 459
rect 2886 459 2892 460
rect 2886 455 2887 459
rect 2891 455 2892 459
rect 2886 454 2892 455
rect 2070 452 2076 453
rect 2070 448 2071 452
rect 2075 448 2076 452
rect 2070 447 2076 448
rect 2030 443 2036 444
rect 2030 439 2031 443
rect 2035 439 2036 443
rect 1934 438 1940 439
rect 2030 438 2036 439
rect 1934 434 1935 438
rect 1939 434 1940 438
rect 1934 433 1940 434
rect 1936 419 1938 433
rect 2032 419 2034 438
rect 2070 435 2076 436
rect 2070 431 2071 435
rect 2075 431 2076 435
rect 2070 430 2076 431
rect 2510 430 2516 431
rect 1935 418 1939 419
rect 1935 413 1939 414
rect 2031 418 2035 419
rect 2031 413 2035 414
rect 1936 403 1938 413
rect 1934 402 1940 403
rect 1934 398 1935 402
rect 1939 398 1940 402
rect 2032 398 2034 413
rect 2072 403 2074 430
rect 2510 426 2511 430
rect 2515 426 2516 430
rect 2510 425 2516 426
rect 2614 430 2620 431
rect 2614 426 2615 430
rect 2619 426 2620 430
rect 2614 425 2620 426
rect 2734 430 2740 431
rect 2734 426 2735 430
rect 2739 426 2740 430
rect 2734 425 2740 426
rect 2862 430 2868 431
rect 2862 426 2863 430
rect 2867 426 2868 430
rect 2862 425 2868 426
rect 2512 403 2514 425
rect 2616 403 2618 425
rect 2736 403 2738 425
rect 2864 403 2866 425
rect 2071 402 2075 403
rect 1934 397 1940 398
rect 2030 397 2036 398
rect 2071 397 2075 398
rect 2511 402 2515 403
rect 2511 397 2515 398
rect 2591 402 2595 403
rect 2591 397 2595 398
rect 2615 402 2619 403
rect 2615 397 2619 398
rect 2695 402 2699 403
rect 2695 397 2699 398
rect 2735 402 2739 403
rect 2735 397 2739 398
rect 2815 402 2819 403
rect 2815 397 2819 398
rect 2863 402 2867 403
rect 2863 397 2867 398
rect 2030 393 2031 397
rect 2035 393 2036 397
rect 2030 392 2036 393
rect 2072 382 2074 397
rect 2592 387 2594 397
rect 2696 387 2698 397
rect 2816 387 2818 397
rect 2590 386 2596 387
rect 2590 382 2591 386
rect 2595 382 2596 386
rect 2070 381 2076 382
rect 2590 381 2596 382
rect 2694 386 2700 387
rect 2694 382 2695 386
rect 2699 382 2700 386
rect 2694 381 2700 382
rect 2814 386 2820 387
rect 2814 382 2815 386
rect 2819 382 2820 386
rect 2814 381 2820 382
rect 2030 380 2036 381
rect 2030 376 2031 380
rect 2035 376 2036 380
rect 2070 377 2071 381
rect 2075 377 2076 381
rect 2070 376 2076 377
rect 2030 375 2036 376
rect 1558 371 1564 372
rect 1558 367 1559 371
rect 1563 367 1564 371
rect 1558 366 1564 367
rect 1686 371 1692 372
rect 1686 367 1687 371
rect 1691 367 1692 371
rect 1686 366 1692 367
rect 1774 371 1780 372
rect 1774 367 1775 371
rect 1779 367 1780 371
rect 1774 366 1780 367
rect 1846 371 1852 372
rect 1846 367 1847 371
rect 1851 367 1852 371
rect 1846 366 1852 367
rect 1446 361 1452 362
rect 1446 357 1447 361
rect 1451 357 1452 361
rect 1446 356 1452 357
rect 1406 351 1412 352
rect 1406 347 1407 351
rect 1411 347 1412 351
rect 1406 346 1412 347
rect 1448 335 1450 356
rect 1560 352 1562 366
rect 1574 361 1580 362
rect 1574 357 1575 361
rect 1579 357 1580 361
rect 1574 356 1580 357
rect 1558 351 1564 352
rect 1558 347 1559 351
rect 1563 347 1564 351
rect 1558 346 1564 347
rect 1576 335 1578 356
rect 1688 352 1690 366
rect 1702 361 1708 362
rect 1702 357 1703 361
rect 1707 357 1708 361
rect 1702 356 1708 357
rect 1686 351 1692 352
rect 1686 347 1687 351
rect 1691 347 1692 351
rect 1686 346 1692 347
rect 1686 335 1692 336
rect 1704 335 1706 356
rect 1047 334 1051 335
rect 1047 329 1051 330
rect 1127 334 1131 335
rect 1127 329 1131 330
rect 1183 334 1187 335
rect 1183 329 1187 330
rect 1311 334 1315 335
rect 1311 329 1315 330
rect 1319 334 1323 335
rect 1319 329 1323 330
rect 1447 334 1451 335
rect 1447 329 1451 330
rect 1503 334 1507 335
rect 1503 329 1507 330
rect 1575 334 1579 335
rect 1686 331 1687 335
rect 1691 331 1692 335
rect 1686 330 1692 331
rect 1703 334 1707 335
rect 1575 329 1579 330
rect 1128 320 1130 329
rect 1312 320 1314 329
rect 1382 327 1388 328
rect 1382 323 1383 327
rect 1387 323 1388 327
rect 1382 322 1388 323
rect 1126 319 1132 320
rect 1126 315 1127 319
rect 1131 315 1132 319
rect 1126 314 1132 315
rect 1310 319 1316 320
rect 1310 315 1311 319
rect 1315 315 1316 319
rect 1310 314 1316 315
rect 966 307 972 308
rect 966 303 967 307
rect 971 303 972 307
rect 966 302 972 303
rect 942 278 948 279
rect 942 274 943 278
rect 947 274 948 278
rect 942 273 948 274
rect 1126 278 1132 279
rect 1126 274 1127 278
rect 1131 274 1132 278
rect 1126 273 1132 274
rect 1310 278 1316 279
rect 1310 274 1311 278
rect 1315 274 1316 278
rect 1310 273 1316 274
rect 944 255 946 273
rect 1128 255 1130 273
rect 1312 255 1314 273
rect 943 254 947 255
rect 943 249 947 250
rect 975 254 979 255
rect 975 249 979 250
rect 1127 254 1131 255
rect 1127 249 1131 250
rect 1175 254 1179 255
rect 1175 249 1179 250
rect 1311 254 1315 255
rect 1311 249 1315 250
rect 1375 254 1379 255
rect 1375 249 1379 250
rect 976 239 978 249
rect 1176 239 1178 249
rect 1376 239 1378 249
rect 974 238 980 239
rect 974 234 975 238
rect 979 234 980 238
rect 974 233 980 234
rect 1174 238 1180 239
rect 1174 234 1175 238
rect 1179 234 1180 238
rect 1174 233 1180 234
rect 1374 238 1380 239
rect 1374 234 1375 238
rect 1379 234 1380 238
rect 1374 233 1380 234
rect 1384 208 1386 322
rect 1504 320 1506 329
rect 1502 319 1508 320
rect 1502 315 1503 319
rect 1507 315 1508 319
rect 1502 314 1508 315
rect 1688 312 1690 330
rect 1703 329 1707 330
rect 1704 320 1706 329
rect 1776 328 1778 366
rect 1830 361 1836 362
rect 1830 357 1831 361
rect 1835 357 1836 361
rect 1830 356 1836 357
rect 1934 361 1940 362
rect 1934 357 1935 361
rect 1939 357 1940 361
rect 1934 356 1940 357
rect 1832 335 1834 356
rect 1936 335 1938 356
rect 2032 335 2034 375
rect 2070 364 2076 365
rect 2070 360 2071 364
rect 2075 360 2076 364
rect 2070 359 2076 360
rect 1831 334 1835 335
rect 1831 329 1835 330
rect 1903 334 1907 335
rect 1903 329 1907 330
rect 1935 334 1939 335
rect 1935 329 1939 330
rect 2031 334 2035 335
rect 2072 331 2074 359
rect 2094 351 2100 352
rect 2094 347 2095 351
rect 2099 347 2100 351
rect 2094 346 2100 347
rect 2031 329 2035 330
rect 2071 330 2075 331
rect 1774 327 1780 328
rect 1774 323 1775 327
rect 1779 323 1780 327
rect 1774 322 1780 323
rect 1904 320 1906 329
rect 1702 319 1708 320
rect 1702 315 1703 319
rect 1707 315 1708 319
rect 1702 314 1708 315
rect 1902 319 1908 320
rect 1902 315 1903 319
rect 1907 315 1908 319
rect 1902 314 1908 315
rect 1686 311 1692 312
rect 1686 307 1687 311
rect 1691 307 1692 311
rect 1686 306 1692 307
rect 1894 307 1900 308
rect 1894 303 1895 307
rect 1899 303 1900 307
rect 1894 302 1900 303
rect 1502 278 1508 279
rect 1502 274 1503 278
rect 1507 274 1508 278
rect 1502 273 1508 274
rect 1702 278 1708 279
rect 1702 274 1703 278
rect 1707 274 1708 278
rect 1702 273 1708 274
rect 1504 255 1506 273
rect 1704 255 1706 273
rect 1503 254 1507 255
rect 1503 249 1507 250
rect 1583 254 1587 255
rect 1583 249 1587 250
rect 1703 254 1707 255
rect 1703 249 1707 250
rect 1799 254 1803 255
rect 1799 249 1803 250
rect 1584 239 1586 249
rect 1800 239 1802 249
rect 1582 238 1588 239
rect 1582 234 1583 238
rect 1587 234 1588 238
rect 1582 233 1588 234
rect 1798 238 1804 239
rect 1798 234 1799 238
rect 1803 234 1804 238
rect 1798 233 1804 234
rect 1158 207 1164 208
rect 1158 203 1159 207
rect 1163 203 1164 207
rect 1158 202 1164 203
rect 1358 207 1364 208
rect 1358 203 1359 207
rect 1363 203 1364 207
rect 1358 202 1364 203
rect 1382 207 1388 208
rect 1382 203 1383 207
rect 1387 203 1388 207
rect 1382 202 1388 203
rect 974 197 980 198
rect 974 193 975 197
rect 979 193 980 197
rect 974 192 980 193
rect 854 187 860 188
rect 854 183 855 187
rect 859 183 860 187
rect 854 182 860 183
rect 976 159 978 192
rect 1160 188 1162 202
rect 1174 197 1180 198
rect 1174 193 1175 197
rect 1179 193 1180 197
rect 1174 192 1180 193
rect 1038 187 1044 188
rect 1038 183 1039 187
rect 1043 183 1044 187
rect 1038 182 1044 183
rect 1158 187 1164 188
rect 1158 183 1159 187
rect 1163 183 1164 187
rect 1158 182 1164 183
rect 111 158 115 159
rect 111 153 115 154
rect 151 158 155 159
rect 230 155 231 159
rect 235 155 236 159
rect 230 154 236 155
rect 255 158 259 159
rect 151 153 155 154
rect 255 153 259 154
rect 279 158 283 159
rect 279 153 283 154
rect 359 158 363 159
rect 359 153 363 154
rect 431 158 435 159
rect 431 153 435 154
rect 471 158 475 159
rect 471 153 475 154
rect 599 158 603 159
rect 599 153 603 154
rect 607 158 611 159
rect 607 153 611 154
rect 743 158 747 159
rect 743 153 747 154
rect 783 158 787 159
rect 783 153 787 154
rect 879 158 883 159
rect 879 153 883 154
rect 975 158 979 159
rect 975 153 979 154
rect 1015 158 1019 159
rect 1015 153 1019 154
rect 112 125 114 153
rect 152 144 154 153
rect 256 144 258 153
rect 360 144 362 153
rect 472 144 474 153
rect 608 144 610 153
rect 744 144 746 153
rect 880 144 882 153
rect 1016 144 1018 153
rect 150 143 156 144
rect 150 139 151 143
rect 155 139 156 143
rect 150 138 156 139
rect 254 143 260 144
rect 254 139 255 143
rect 259 139 260 143
rect 254 138 260 139
rect 358 143 364 144
rect 358 139 359 143
rect 363 139 364 143
rect 358 138 364 139
rect 470 143 476 144
rect 470 139 471 143
rect 475 139 476 143
rect 470 138 476 139
rect 606 143 612 144
rect 606 139 607 143
rect 611 139 612 143
rect 606 138 612 139
rect 742 143 748 144
rect 742 139 743 143
rect 747 139 748 143
rect 742 138 748 139
rect 878 143 884 144
rect 878 139 879 143
rect 883 139 884 143
rect 878 138 884 139
rect 1014 143 1020 144
rect 1014 139 1015 143
rect 1019 139 1020 143
rect 1014 138 1020 139
rect 1040 132 1042 182
rect 1176 159 1178 192
rect 1360 188 1362 202
rect 1374 197 1380 198
rect 1374 193 1375 197
rect 1379 193 1380 197
rect 1374 192 1380 193
rect 1582 197 1588 198
rect 1582 193 1583 197
rect 1587 193 1588 197
rect 1582 192 1588 193
rect 1798 197 1804 198
rect 1798 193 1799 197
rect 1803 193 1804 197
rect 1798 192 1804 193
rect 1358 187 1364 188
rect 1358 183 1359 187
rect 1363 183 1364 187
rect 1358 182 1364 183
rect 1376 159 1378 192
rect 1584 159 1586 192
rect 1800 159 1802 192
rect 1896 188 1898 302
rect 2032 301 2034 329
rect 2071 325 2075 326
rect 2030 300 2036 301
rect 2030 296 2031 300
rect 2035 296 2036 300
rect 2072 297 2074 325
rect 2096 324 2098 346
rect 2590 345 2596 346
rect 2590 341 2591 345
rect 2595 341 2596 345
rect 2590 340 2596 341
rect 2694 345 2700 346
rect 2694 341 2695 345
rect 2699 341 2700 345
rect 2694 340 2700 341
rect 2814 345 2820 346
rect 2814 341 2815 345
rect 2819 341 2820 345
rect 2814 340 2820 341
rect 2592 331 2594 340
rect 2696 331 2698 340
rect 2816 331 2818 340
rect 2888 336 2890 454
rect 3006 430 3012 431
rect 3006 426 3007 430
rect 3011 426 3012 430
rect 3006 425 3012 426
rect 3158 430 3164 431
rect 3158 426 3159 430
rect 3163 426 3164 430
rect 3158 425 3164 426
rect 3318 430 3324 431
rect 3318 426 3319 430
rect 3323 426 3324 430
rect 3318 425 3324 426
rect 3008 403 3010 425
rect 3160 403 3162 425
rect 3320 403 3322 425
rect 3392 416 3394 474
rect 3480 472 3482 481
rect 3648 472 3650 481
rect 3720 480 3722 510
rect 3822 509 3828 510
rect 3822 505 3823 509
rect 3827 505 3828 509
rect 3822 504 3828 505
rect 3824 487 3826 504
rect 3896 500 3898 614
rect 3992 613 3994 641
rect 3990 612 3996 613
rect 3990 608 3991 612
rect 3995 608 3996 612
rect 3990 607 3996 608
rect 3990 595 3996 596
rect 3990 591 3991 595
rect 3995 591 3996 595
rect 3990 590 3996 591
rect 3992 567 3994 590
rect 3991 566 3995 567
rect 3991 561 3995 562
rect 3992 546 3994 561
rect 3990 545 3996 546
rect 3990 541 3991 545
rect 3995 541 3996 545
rect 3990 540 3996 541
rect 3990 528 3996 529
rect 3990 524 3991 528
rect 3995 524 3996 528
rect 3990 523 3996 524
rect 3894 499 3900 500
rect 3894 495 3895 499
rect 3899 495 3900 499
rect 3894 494 3900 495
rect 3992 487 3994 523
rect 3823 486 3827 487
rect 3823 481 3827 482
rect 3991 486 3995 487
rect 3991 481 3995 482
rect 3718 479 3724 480
rect 3718 475 3719 479
rect 3723 475 3724 479
rect 3718 474 3724 475
rect 3824 472 3826 481
rect 3838 479 3844 480
rect 3838 475 3839 479
rect 3843 475 3844 479
rect 3838 474 3844 475
rect 3478 471 3484 472
rect 3478 467 3479 471
rect 3483 467 3484 471
rect 3478 466 3484 467
rect 3646 471 3652 472
rect 3646 467 3647 471
rect 3651 467 3652 471
rect 3646 466 3652 467
rect 3822 471 3828 472
rect 3822 467 3823 471
rect 3827 467 3828 471
rect 3822 466 3828 467
rect 3586 463 3592 464
rect 3586 459 3587 463
rect 3591 459 3592 463
rect 3586 458 3592 459
rect 3478 430 3484 431
rect 3478 426 3479 430
rect 3483 426 3484 430
rect 3478 425 3484 426
rect 3390 415 3396 416
rect 3390 411 3391 415
rect 3395 411 3396 415
rect 3390 410 3396 411
rect 3480 403 3482 425
rect 3588 404 3590 458
rect 3646 430 3652 431
rect 3646 426 3647 430
rect 3651 426 3652 430
rect 3646 425 3652 426
rect 3822 430 3828 431
rect 3822 426 3823 430
rect 3827 426 3828 430
rect 3822 425 3828 426
rect 3586 403 3592 404
rect 3648 403 3650 425
rect 3782 403 3788 404
rect 3824 403 3826 425
rect 2959 402 2963 403
rect 2959 397 2963 398
rect 3007 402 3011 403
rect 3007 397 3011 398
rect 3119 402 3123 403
rect 3119 397 3123 398
rect 3159 402 3163 403
rect 3159 397 3163 398
rect 3303 402 3307 403
rect 3303 397 3307 398
rect 3319 402 3323 403
rect 3319 397 3323 398
rect 3479 402 3483 403
rect 3479 397 3483 398
rect 3503 402 3507 403
rect 3586 399 3587 403
rect 3591 399 3592 403
rect 3586 398 3592 399
rect 3647 402 3651 403
rect 3503 397 3507 398
rect 3647 397 3651 398
rect 3711 402 3715 403
rect 3782 399 3783 403
rect 3787 399 3788 403
rect 3782 398 3788 399
rect 3823 402 3827 403
rect 3711 397 3715 398
rect 2960 387 2962 397
rect 3120 387 3122 397
rect 3304 387 3306 397
rect 3504 387 3506 397
rect 3712 387 3714 397
rect 2958 386 2964 387
rect 2958 382 2959 386
rect 2963 382 2964 386
rect 2958 381 2964 382
rect 3118 386 3124 387
rect 3118 382 3119 386
rect 3123 382 3124 386
rect 3118 381 3124 382
rect 3302 386 3308 387
rect 3302 382 3303 386
rect 3307 382 3308 386
rect 3302 381 3308 382
rect 3502 386 3508 387
rect 3502 382 3503 386
rect 3507 382 3508 386
rect 3502 381 3508 382
rect 3710 386 3716 387
rect 3710 382 3711 386
rect 3715 382 3716 386
rect 3710 381 3716 382
rect 2958 345 2964 346
rect 2958 341 2959 345
rect 2963 341 2964 345
rect 2958 340 2964 341
rect 3118 345 3124 346
rect 3118 341 3119 345
rect 3123 341 3124 345
rect 3118 340 3124 341
rect 3302 345 3308 346
rect 3302 341 3303 345
rect 3307 341 3308 345
rect 3302 340 3308 341
rect 3502 345 3508 346
rect 3502 341 3503 345
rect 3507 341 3508 345
rect 3502 340 3508 341
rect 3710 345 3716 346
rect 3710 341 3711 345
rect 3715 341 3716 345
rect 3710 340 3716 341
rect 2886 335 2892 336
rect 2886 331 2887 335
rect 2891 331 2892 335
rect 2960 331 2962 340
rect 3120 331 3122 340
rect 3304 331 3306 340
rect 3504 331 3506 340
rect 3510 335 3516 336
rect 3510 331 3511 335
rect 3515 331 3516 335
rect 3712 331 3714 340
rect 3784 336 3786 398
rect 3823 397 3827 398
rect 3840 356 3842 474
rect 3958 463 3964 464
rect 3958 459 3959 463
rect 3963 459 3964 463
rect 3958 458 3964 459
rect 3895 402 3899 403
rect 3895 397 3899 398
rect 3896 387 3898 397
rect 3894 386 3900 387
rect 3894 382 3895 386
rect 3899 382 3900 386
rect 3894 381 3900 382
rect 3838 355 3844 356
rect 3838 351 3839 355
rect 3843 351 3844 355
rect 3838 350 3844 351
rect 3894 345 3900 346
rect 3894 341 3895 345
rect 3899 341 3900 345
rect 3894 340 3900 341
rect 3782 335 3788 336
rect 3782 331 3783 335
rect 3787 331 3788 335
rect 3896 331 3898 340
rect 3960 336 3962 458
rect 3992 453 3994 481
rect 3990 452 3996 453
rect 3990 448 3991 452
rect 3995 448 3996 452
rect 3990 447 3996 448
rect 3990 435 3996 436
rect 3990 431 3991 435
rect 3995 431 3996 435
rect 3990 430 3996 431
rect 3992 403 3994 430
rect 3991 402 3995 403
rect 3991 397 3995 398
rect 3992 382 3994 397
rect 3990 381 3996 382
rect 3990 377 3991 381
rect 3995 377 3996 381
rect 3990 376 3996 377
rect 3990 364 3996 365
rect 3990 360 3991 364
rect 3995 360 3996 364
rect 3990 359 3996 360
rect 3966 355 3972 356
rect 3966 351 3967 355
rect 3971 351 3972 355
rect 3966 350 3972 351
rect 3958 335 3964 336
rect 3958 331 3959 335
rect 3963 331 3964 335
rect 2111 330 2115 331
rect 2111 325 2115 326
rect 2271 330 2275 331
rect 2271 325 2275 326
rect 2455 330 2459 331
rect 2455 325 2459 326
rect 2591 330 2595 331
rect 2591 325 2595 326
rect 2631 330 2635 331
rect 2631 325 2635 326
rect 2695 330 2699 331
rect 2695 325 2699 326
rect 2807 330 2811 331
rect 2807 325 2811 326
rect 2815 330 2819 331
rect 2886 330 2892 331
rect 2959 330 2963 331
rect 2815 325 2819 326
rect 2959 325 2963 326
rect 2999 330 3003 331
rect 2999 325 3003 326
rect 3119 330 3123 331
rect 3119 325 3123 326
rect 3215 330 3219 331
rect 3215 325 3219 326
rect 3303 330 3307 331
rect 3303 325 3307 326
rect 3439 330 3443 331
rect 3439 325 3443 326
rect 3503 330 3507 331
rect 3510 330 3516 331
rect 3679 330 3683 331
rect 3503 325 3507 326
rect 2094 323 2100 324
rect 2094 319 2095 323
rect 2099 319 2100 323
rect 2094 318 2100 319
rect 2112 316 2114 325
rect 2272 316 2274 325
rect 2456 316 2458 325
rect 2462 323 2468 324
rect 2462 319 2463 323
rect 2467 319 2468 323
rect 2462 318 2468 319
rect 2110 315 2116 316
rect 2110 311 2111 315
rect 2115 311 2116 315
rect 2110 310 2116 311
rect 2270 315 2276 316
rect 2270 311 2271 315
rect 2275 311 2276 315
rect 2270 310 2276 311
rect 2454 315 2460 316
rect 2454 311 2455 315
rect 2459 311 2460 315
rect 2454 310 2460 311
rect 2030 295 2036 296
rect 2070 296 2076 297
rect 2070 292 2071 296
rect 2075 292 2076 296
rect 2070 291 2076 292
rect 2030 283 2036 284
rect 2030 279 2031 283
rect 2035 279 2036 283
rect 1902 278 1908 279
rect 2030 278 2036 279
rect 2070 279 2076 280
rect 1902 274 1903 278
rect 1907 274 1908 278
rect 1902 273 1908 274
rect 1904 255 1906 273
rect 2032 255 2034 278
rect 2070 275 2071 279
rect 2075 275 2076 279
rect 2070 274 2076 275
rect 2110 274 2116 275
rect 2072 259 2074 274
rect 2110 270 2111 274
rect 2115 270 2116 274
rect 2110 269 2116 270
rect 2270 274 2276 275
rect 2270 270 2271 274
rect 2275 270 2276 274
rect 2270 269 2276 270
rect 2454 274 2460 275
rect 2454 270 2455 274
rect 2459 270 2460 274
rect 2454 269 2460 270
rect 2112 259 2114 269
rect 2272 259 2274 269
rect 2456 259 2458 269
rect 2071 258 2075 259
rect 1903 254 1907 255
rect 1903 249 1907 250
rect 2031 254 2035 255
rect 2071 253 2075 254
rect 2111 258 2115 259
rect 2111 253 2115 254
rect 2271 258 2275 259
rect 2271 253 2275 254
rect 2455 258 2459 259
rect 2455 253 2459 254
rect 2031 249 2035 250
rect 2032 234 2034 249
rect 2072 238 2074 253
rect 2112 243 2114 253
rect 2272 243 2274 253
rect 2110 242 2116 243
rect 2110 238 2111 242
rect 2115 238 2116 242
rect 2070 237 2076 238
rect 2110 237 2116 238
rect 2270 242 2276 243
rect 2270 238 2271 242
rect 2275 238 2276 242
rect 2270 237 2276 238
rect 2030 233 2036 234
rect 2030 229 2031 233
rect 2035 229 2036 233
rect 2070 233 2071 237
rect 2075 233 2076 237
rect 2070 232 2076 233
rect 2030 228 2036 229
rect 2070 220 2076 221
rect 2030 216 2036 217
rect 2030 212 2031 216
rect 2035 212 2036 216
rect 2070 216 2071 220
rect 2075 216 2076 220
rect 2070 215 2076 216
rect 2030 211 2036 212
rect 1894 187 1900 188
rect 1894 183 1895 187
rect 1899 183 1900 187
rect 1894 182 1900 183
rect 2032 159 2034 211
rect 2072 159 2074 215
rect 2464 212 2466 318
rect 2632 316 2634 325
rect 2808 316 2810 325
rect 2983 316 2987 317
rect 3000 316 3002 325
rect 3216 316 3218 325
rect 3440 316 3442 325
rect 3512 317 3514 330
rect 3679 325 3683 326
rect 3711 330 3715 331
rect 3782 330 3788 331
rect 3895 330 3899 331
rect 3958 330 3964 331
rect 3711 325 3715 326
rect 3895 325 3899 326
rect 3511 316 3515 317
rect 3680 316 3682 325
rect 3686 323 3692 324
rect 3686 319 3687 323
rect 3691 319 3692 323
rect 3686 318 3692 319
rect 2630 315 2636 316
rect 2630 311 2631 315
rect 2635 311 2636 315
rect 2630 310 2636 311
rect 2806 315 2812 316
rect 2806 311 2807 315
rect 2811 311 2812 315
rect 2983 311 2987 312
rect 2998 315 3004 316
rect 2998 311 2999 315
rect 3003 311 3004 315
rect 2806 310 2812 311
rect 2984 308 2986 311
rect 2998 310 3004 311
rect 3214 315 3220 316
rect 3214 311 3215 315
rect 3219 311 3220 315
rect 3214 310 3220 311
rect 3438 315 3444 316
rect 3438 311 3439 315
rect 3443 311 3444 315
rect 3511 311 3515 312
rect 3678 315 3684 316
rect 3678 311 3679 315
rect 3683 311 3684 315
rect 3438 310 3444 311
rect 3678 310 3684 311
rect 2758 307 2764 308
rect 2758 303 2759 307
rect 2763 303 2764 307
rect 2758 302 2764 303
rect 2982 307 2988 308
rect 2982 303 2983 307
rect 2987 303 2988 307
rect 2982 302 2988 303
rect 2630 274 2636 275
rect 2630 270 2631 274
rect 2635 270 2636 274
rect 2630 269 2636 270
rect 2632 259 2634 269
rect 2471 258 2475 259
rect 2471 253 2475 254
rect 2631 258 2635 259
rect 2631 253 2635 254
rect 2687 258 2691 259
rect 2687 253 2691 254
rect 2472 243 2474 253
rect 2688 243 2690 253
rect 2470 242 2476 243
rect 2470 238 2471 242
rect 2475 238 2476 242
rect 2470 237 2476 238
rect 2686 242 2692 243
rect 2686 238 2687 242
rect 2691 238 2692 242
rect 2686 237 2692 238
rect 2254 211 2260 212
rect 2254 207 2255 211
rect 2259 207 2260 211
rect 2254 206 2260 207
rect 2454 211 2460 212
rect 2454 207 2455 211
rect 2459 207 2460 211
rect 2454 206 2460 207
rect 2462 211 2468 212
rect 2462 207 2463 211
rect 2467 207 2468 211
rect 2462 206 2468 207
rect 2110 201 2116 202
rect 2110 197 2111 201
rect 2115 197 2116 201
rect 2110 196 2116 197
rect 2112 159 2114 196
rect 2256 192 2258 206
rect 2270 201 2276 202
rect 2270 197 2271 201
rect 2275 197 2276 201
rect 2270 196 2276 197
rect 2174 191 2180 192
rect 2174 187 2175 191
rect 2179 187 2180 191
rect 2174 186 2180 187
rect 2254 191 2260 192
rect 2254 187 2255 191
rect 2259 187 2260 191
rect 2254 186 2260 187
rect 1151 158 1155 159
rect 1151 153 1155 154
rect 1175 158 1179 159
rect 1175 153 1179 154
rect 1279 158 1283 159
rect 1279 153 1283 154
rect 1375 158 1379 159
rect 1375 153 1379 154
rect 1399 158 1403 159
rect 1399 153 1403 154
rect 1519 158 1523 159
rect 1519 153 1523 154
rect 1583 158 1587 159
rect 1583 153 1587 154
rect 1647 158 1651 159
rect 1647 153 1651 154
rect 1775 158 1779 159
rect 1775 153 1779 154
rect 1799 158 1803 159
rect 1799 153 1803 154
rect 2031 158 2035 159
rect 2031 153 2035 154
rect 2071 158 2075 159
rect 2071 153 2075 154
rect 2111 158 2115 159
rect 2111 153 2115 154
rect 1152 144 1154 153
rect 1280 144 1282 153
rect 1400 144 1402 153
rect 1520 144 1522 153
rect 1648 144 1650 153
rect 1776 144 1778 153
rect 1150 143 1156 144
rect 1150 139 1151 143
rect 1155 139 1156 143
rect 1150 138 1156 139
rect 1278 143 1284 144
rect 1278 139 1279 143
rect 1283 139 1284 143
rect 1278 138 1284 139
rect 1398 143 1404 144
rect 1398 139 1399 143
rect 1403 139 1404 143
rect 1398 138 1404 139
rect 1518 143 1524 144
rect 1518 139 1519 143
rect 1523 139 1524 143
rect 1518 138 1524 139
rect 1646 143 1652 144
rect 1646 139 1647 143
rect 1651 139 1652 143
rect 1646 138 1652 139
rect 1774 143 1780 144
rect 1774 139 1775 143
rect 1779 139 1780 143
rect 1774 138 1780 139
rect 1038 131 1044 132
rect 1038 127 1039 131
rect 1043 127 1044 131
rect 1038 126 1044 127
rect 2032 125 2034 153
rect 2072 125 2074 153
rect 2112 144 2114 153
rect 2110 143 2116 144
rect 2110 139 2111 143
rect 2115 139 2116 143
rect 2110 138 2116 139
rect 2176 136 2178 186
rect 2272 159 2274 196
rect 2456 192 2458 206
rect 2470 201 2476 202
rect 2470 197 2471 201
rect 2475 197 2476 201
rect 2470 196 2476 197
rect 2686 201 2692 202
rect 2686 197 2687 201
rect 2691 197 2692 201
rect 2686 196 2692 197
rect 2454 191 2460 192
rect 2454 187 2455 191
rect 2459 187 2460 191
rect 2454 186 2460 187
rect 2472 159 2474 196
rect 2688 159 2690 196
rect 2760 192 2762 302
rect 2806 274 2812 275
rect 2806 270 2807 274
rect 2811 270 2812 274
rect 2806 269 2812 270
rect 2998 274 3004 275
rect 2998 270 2999 274
rect 3003 270 3004 274
rect 2998 269 3004 270
rect 3214 274 3220 275
rect 3214 270 3215 274
rect 3219 270 3220 274
rect 3214 269 3220 270
rect 3438 274 3444 275
rect 3438 270 3439 274
rect 3443 270 3444 274
rect 3438 269 3444 270
rect 3678 274 3684 275
rect 3678 270 3679 274
rect 3683 270 3684 274
rect 3678 269 3684 270
rect 2808 259 2810 269
rect 3000 259 3002 269
rect 3216 259 3218 269
rect 3440 259 3442 269
rect 3680 259 3682 269
rect 2807 258 2811 259
rect 2807 253 2811 254
rect 2903 258 2907 259
rect 2903 253 2907 254
rect 2999 258 3003 259
rect 2999 253 3003 254
rect 3111 258 3115 259
rect 3111 253 3115 254
rect 3215 258 3219 259
rect 3215 253 3219 254
rect 3319 258 3323 259
rect 3319 253 3323 254
rect 3439 258 3443 259
rect 3439 253 3443 254
rect 3519 258 3523 259
rect 3519 253 3523 254
rect 3679 258 3683 259
rect 3679 253 3683 254
rect 2904 243 2906 253
rect 3112 243 3114 253
rect 3320 243 3322 253
rect 3520 243 3522 253
rect 2902 242 2908 243
rect 2902 238 2903 242
rect 2907 238 2908 242
rect 2902 237 2908 238
rect 3110 242 3116 243
rect 3110 238 3111 242
rect 3115 238 3116 242
rect 3110 237 3116 238
rect 3318 242 3324 243
rect 3318 238 3319 242
rect 3323 238 3324 242
rect 3318 237 3324 238
rect 3518 242 3524 243
rect 3518 238 3519 242
rect 3523 238 3524 242
rect 3518 237 3524 238
rect 3688 232 3690 318
rect 3896 316 3898 325
rect 3968 324 3970 350
rect 3992 331 3994 359
rect 3991 330 3995 331
rect 3991 325 3995 326
rect 3966 323 3972 324
rect 3966 319 3967 323
rect 3971 319 3972 323
rect 3966 318 3972 319
rect 3894 315 3900 316
rect 3894 311 3895 315
rect 3899 311 3900 315
rect 3894 310 3900 311
rect 3958 307 3964 308
rect 3958 303 3959 307
rect 3963 303 3964 307
rect 3958 302 3964 303
rect 3894 274 3900 275
rect 3894 270 3895 274
rect 3899 270 3900 274
rect 3894 269 3900 270
rect 3896 259 3898 269
rect 3719 258 3723 259
rect 3719 253 3723 254
rect 3895 258 3899 259
rect 3895 253 3899 254
rect 3720 243 3722 253
rect 3896 243 3898 253
rect 3718 242 3724 243
rect 3718 238 3719 242
rect 3723 238 3724 242
rect 3718 237 3724 238
rect 3894 242 3900 243
rect 3894 238 3895 242
rect 3899 238 3900 242
rect 3894 237 3900 238
rect 3302 231 3308 232
rect 3302 227 3303 231
rect 3307 227 3308 231
rect 3302 226 3308 227
rect 3686 231 3692 232
rect 3686 227 3687 231
rect 3691 227 3692 231
rect 3686 226 3692 227
rect 3304 212 3306 226
rect 3302 211 3308 212
rect 3302 207 3303 211
rect 3307 207 3308 211
rect 3302 206 3308 207
rect 2902 201 2908 202
rect 2902 197 2903 201
rect 2907 197 2908 201
rect 2902 196 2908 197
rect 3110 201 3116 202
rect 3110 197 3111 201
rect 3115 197 3116 201
rect 3110 196 3116 197
rect 3318 201 3324 202
rect 3318 197 3319 201
rect 3323 197 3324 201
rect 3318 196 3324 197
rect 3518 201 3524 202
rect 3518 197 3519 201
rect 3523 197 3524 201
rect 3518 196 3524 197
rect 3718 201 3724 202
rect 3718 197 3719 201
rect 3723 197 3724 201
rect 3718 196 3724 197
rect 3894 201 3900 202
rect 3894 197 3895 201
rect 3899 197 3900 201
rect 3894 196 3900 197
rect 2758 191 2764 192
rect 2758 187 2759 191
rect 2763 187 2764 191
rect 2758 186 2764 187
rect 2904 159 2906 196
rect 2998 191 3004 192
rect 2998 187 2999 191
rect 3003 187 3004 191
rect 2998 186 3004 187
rect 2215 158 2219 159
rect 2215 153 2219 154
rect 2271 158 2275 159
rect 2271 153 2275 154
rect 2319 158 2323 159
rect 2319 153 2323 154
rect 2423 158 2427 159
rect 2423 153 2427 154
rect 2471 158 2475 159
rect 2471 153 2475 154
rect 2527 158 2531 159
rect 2527 153 2531 154
rect 2655 158 2659 159
rect 2655 153 2659 154
rect 2687 158 2691 159
rect 2687 153 2691 154
rect 2775 158 2779 159
rect 2775 153 2779 154
rect 2895 158 2899 159
rect 2895 153 2899 154
rect 2903 158 2907 159
rect 2903 153 2907 154
rect 2216 144 2218 153
rect 2320 144 2322 153
rect 2424 144 2426 153
rect 2528 144 2530 153
rect 2656 144 2658 153
rect 2776 144 2778 153
rect 2896 144 2898 153
rect 2214 143 2220 144
rect 2214 139 2215 143
rect 2219 139 2220 143
rect 2214 138 2220 139
rect 2318 143 2324 144
rect 2318 139 2319 143
rect 2323 139 2324 143
rect 2318 138 2324 139
rect 2422 143 2428 144
rect 2422 139 2423 143
rect 2427 139 2428 143
rect 2422 138 2428 139
rect 2526 143 2532 144
rect 2526 139 2527 143
rect 2531 139 2532 143
rect 2526 138 2532 139
rect 2654 143 2660 144
rect 2654 139 2655 143
rect 2659 139 2660 143
rect 2654 138 2660 139
rect 2774 143 2780 144
rect 2774 139 2775 143
rect 2779 139 2780 143
rect 2774 138 2780 139
rect 2894 143 2900 144
rect 2894 139 2895 143
rect 2899 139 2900 143
rect 2894 138 2900 139
rect 3000 136 3002 186
rect 3112 159 3114 196
rect 3320 159 3322 196
rect 3520 159 3522 196
rect 3720 159 3722 196
rect 3782 191 3788 192
rect 3782 187 3783 191
rect 3787 187 3788 191
rect 3782 186 3788 187
rect 3015 158 3019 159
rect 3015 153 3019 154
rect 3111 158 3115 159
rect 3111 153 3115 154
rect 3135 158 3139 159
rect 3135 153 3139 154
rect 3247 158 3251 159
rect 3247 153 3251 154
rect 3319 158 3323 159
rect 3319 153 3323 154
rect 3359 158 3363 159
rect 3359 153 3363 154
rect 3471 158 3475 159
rect 3471 153 3475 154
rect 3519 158 3523 159
rect 3519 153 3523 154
rect 3583 158 3587 159
rect 3583 153 3587 154
rect 3687 158 3691 159
rect 3687 153 3691 154
rect 3719 158 3723 159
rect 3719 153 3723 154
rect 3016 144 3018 153
rect 3136 144 3138 153
rect 3248 144 3250 153
rect 3360 144 3362 153
rect 3472 144 3474 153
rect 3584 144 3586 153
rect 3688 144 3690 153
rect 3014 143 3020 144
rect 3014 139 3015 143
rect 3019 139 3020 143
rect 3014 138 3020 139
rect 3134 143 3140 144
rect 3134 139 3135 143
rect 3139 139 3140 143
rect 3134 138 3140 139
rect 3246 143 3252 144
rect 3246 139 3247 143
rect 3251 139 3252 143
rect 3246 138 3252 139
rect 3358 143 3364 144
rect 3358 139 3359 143
rect 3363 139 3364 143
rect 3358 138 3364 139
rect 3470 143 3476 144
rect 3470 139 3471 143
rect 3475 139 3476 143
rect 3470 138 3476 139
rect 3582 143 3588 144
rect 3582 139 3583 143
rect 3587 139 3588 143
rect 3582 138 3588 139
rect 3686 143 3692 144
rect 3686 139 3687 143
rect 3691 139 3692 143
rect 3686 138 3692 139
rect 3784 136 3786 186
rect 3896 159 3898 196
rect 3960 192 3962 302
rect 3992 297 3994 325
rect 3990 296 3996 297
rect 3990 292 3991 296
rect 3995 292 3996 296
rect 3990 291 3996 292
rect 3990 279 3996 280
rect 3990 275 3991 279
rect 3995 275 3996 279
rect 3990 274 3996 275
rect 3992 259 3994 274
rect 3991 258 3995 259
rect 3991 253 3995 254
rect 3992 238 3994 253
rect 3990 237 3996 238
rect 3990 233 3991 237
rect 3995 233 3996 237
rect 3990 232 3996 233
rect 3990 220 3996 221
rect 3990 216 3991 220
rect 3995 216 3996 220
rect 3990 215 3996 216
rect 3966 211 3972 212
rect 3966 207 3967 211
rect 3971 207 3972 211
rect 3966 206 3972 207
rect 3958 191 3964 192
rect 3958 187 3959 191
rect 3963 187 3964 191
rect 3958 186 3964 187
rect 3791 158 3795 159
rect 3791 153 3795 154
rect 3895 158 3899 159
rect 3895 153 3899 154
rect 3792 144 3794 153
rect 3896 144 3898 153
rect 3968 152 3970 206
rect 3992 159 3994 215
rect 3991 158 3995 159
rect 3991 153 3995 154
rect 3966 151 3972 152
rect 3966 147 3967 151
rect 3971 147 3972 151
rect 3966 146 3972 147
rect 3790 143 3796 144
rect 3790 139 3791 143
rect 3795 139 3796 143
rect 3790 138 3796 139
rect 3894 143 3900 144
rect 3894 139 3895 143
rect 3899 139 3900 143
rect 3894 138 3900 139
rect 2174 135 2180 136
rect 2174 131 2175 135
rect 2179 131 2180 135
rect 2174 130 2180 131
rect 2998 135 3004 136
rect 2998 131 2999 135
rect 3003 131 3004 135
rect 2998 130 3004 131
rect 3782 135 3788 136
rect 3782 131 3783 135
rect 3787 131 3788 135
rect 3782 130 3788 131
rect 3992 125 3994 153
rect 110 124 116 125
rect 110 120 111 124
rect 115 120 116 124
rect 110 119 116 120
rect 2030 124 2036 125
rect 2030 120 2031 124
rect 2035 120 2036 124
rect 2030 119 2036 120
rect 2070 124 2076 125
rect 2070 120 2071 124
rect 2075 120 2076 124
rect 2070 119 2076 120
rect 3990 124 3996 125
rect 3990 120 3991 124
rect 3995 120 3996 124
rect 3990 119 3996 120
rect 110 107 116 108
rect 110 103 111 107
rect 115 103 116 107
rect 2030 107 2036 108
rect 2030 103 2031 107
rect 2035 103 2036 107
rect 110 102 116 103
rect 150 102 156 103
rect 112 87 114 102
rect 150 98 151 102
rect 155 98 156 102
rect 150 97 156 98
rect 254 102 260 103
rect 254 98 255 102
rect 259 98 260 102
rect 254 97 260 98
rect 358 102 364 103
rect 358 98 359 102
rect 363 98 364 102
rect 358 97 364 98
rect 470 102 476 103
rect 470 98 471 102
rect 475 98 476 102
rect 470 97 476 98
rect 606 102 612 103
rect 606 98 607 102
rect 611 98 612 102
rect 606 97 612 98
rect 742 102 748 103
rect 742 98 743 102
rect 747 98 748 102
rect 742 97 748 98
rect 878 102 884 103
rect 878 98 879 102
rect 883 98 884 102
rect 878 97 884 98
rect 1014 102 1020 103
rect 1014 98 1015 102
rect 1019 98 1020 102
rect 1014 97 1020 98
rect 1150 102 1156 103
rect 1150 98 1151 102
rect 1155 98 1156 102
rect 1150 97 1156 98
rect 1278 102 1284 103
rect 1278 98 1279 102
rect 1283 98 1284 102
rect 1278 97 1284 98
rect 1398 102 1404 103
rect 1398 98 1399 102
rect 1403 98 1404 102
rect 1398 97 1404 98
rect 1518 102 1524 103
rect 1518 98 1519 102
rect 1523 98 1524 102
rect 1518 97 1524 98
rect 1646 102 1652 103
rect 1646 98 1647 102
rect 1651 98 1652 102
rect 1646 97 1652 98
rect 1774 102 1780 103
rect 2030 102 2036 103
rect 2070 107 2076 108
rect 2070 103 2071 107
rect 2075 103 2076 107
rect 3990 107 3996 108
rect 3990 103 3991 107
rect 3995 103 3996 107
rect 2070 102 2076 103
rect 2110 102 2116 103
rect 1774 98 1775 102
rect 1779 98 1780 102
rect 1774 97 1780 98
rect 152 87 154 97
rect 256 87 258 97
rect 360 87 362 97
rect 472 87 474 97
rect 608 87 610 97
rect 744 87 746 97
rect 880 87 882 97
rect 1016 87 1018 97
rect 1152 87 1154 97
rect 1280 87 1282 97
rect 1400 87 1402 97
rect 1520 87 1522 97
rect 1648 87 1650 97
rect 1776 87 1778 97
rect 2032 87 2034 102
rect 2072 87 2074 102
rect 2110 98 2111 102
rect 2115 98 2116 102
rect 2110 97 2116 98
rect 2214 102 2220 103
rect 2214 98 2215 102
rect 2219 98 2220 102
rect 2214 97 2220 98
rect 2318 102 2324 103
rect 2318 98 2319 102
rect 2323 98 2324 102
rect 2318 97 2324 98
rect 2422 102 2428 103
rect 2422 98 2423 102
rect 2427 98 2428 102
rect 2422 97 2428 98
rect 2526 102 2532 103
rect 2526 98 2527 102
rect 2531 98 2532 102
rect 2526 97 2532 98
rect 2654 102 2660 103
rect 2654 98 2655 102
rect 2659 98 2660 102
rect 2654 97 2660 98
rect 2774 102 2780 103
rect 2774 98 2775 102
rect 2779 98 2780 102
rect 2774 97 2780 98
rect 2894 102 2900 103
rect 2894 98 2895 102
rect 2899 98 2900 102
rect 2894 97 2900 98
rect 3014 102 3020 103
rect 3014 98 3015 102
rect 3019 98 3020 102
rect 3014 97 3020 98
rect 3134 102 3140 103
rect 3134 98 3135 102
rect 3139 98 3140 102
rect 3134 97 3140 98
rect 3246 102 3252 103
rect 3246 98 3247 102
rect 3251 98 3252 102
rect 3246 97 3252 98
rect 3358 102 3364 103
rect 3358 98 3359 102
rect 3363 98 3364 102
rect 3358 97 3364 98
rect 3470 102 3476 103
rect 3470 98 3471 102
rect 3475 98 3476 102
rect 3470 97 3476 98
rect 3582 102 3588 103
rect 3582 98 3583 102
rect 3587 98 3588 102
rect 3582 97 3588 98
rect 3686 102 3692 103
rect 3686 98 3687 102
rect 3691 98 3692 102
rect 3686 97 3692 98
rect 3790 102 3796 103
rect 3790 98 3791 102
rect 3795 98 3796 102
rect 3790 97 3796 98
rect 3894 102 3900 103
rect 3990 102 3996 103
rect 3894 98 3895 102
rect 3899 98 3900 102
rect 3894 97 3900 98
rect 2112 87 2114 97
rect 2216 87 2218 97
rect 2320 87 2322 97
rect 2424 87 2426 97
rect 2528 87 2530 97
rect 2656 87 2658 97
rect 2776 87 2778 97
rect 2896 87 2898 97
rect 3016 87 3018 97
rect 3136 87 3138 97
rect 3248 87 3250 97
rect 3360 87 3362 97
rect 3472 87 3474 97
rect 3584 87 3586 97
rect 3688 87 3690 97
rect 3792 87 3794 97
rect 3896 87 3898 97
rect 3992 87 3994 102
rect 111 86 115 87
rect 111 81 115 82
rect 151 86 155 87
rect 151 81 155 82
rect 255 86 259 87
rect 255 81 259 82
rect 359 86 363 87
rect 359 81 363 82
rect 471 86 475 87
rect 471 81 475 82
rect 607 86 611 87
rect 607 81 611 82
rect 743 86 747 87
rect 743 81 747 82
rect 879 86 883 87
rect 879 81 883 82
rect 1015 86 1019 87
rect 1015 81 1019 82
rect 1151 86 1155 87
rect 1151 81 1155 82
rect 1279 86 1283 87
rect 1279 81 1283 82
rect 1399 86 1403 87
rect 1399 81 1403 82
rect 1519 86 1523 87
rect 1519 81 1523 82
rect 1647 86 1651 87
rect 1647 81 1651 82
rect 1775 86 1779 87
rect 1775 81 1779 82
rect 2031 86 2035 87
rect 2031 81 2035 82
rect 2071 86 2075 87
rect 2071 81 2075 82
rect 2111 86 2115 87
rect 2111 81 2115 82
rect 2215 86 2219 87
rect 2215 81 2219 82
rect 2319 86 2323 87
rect 2319 81 2323 82
rect 2423 86 2427 87
rect 2423 81 2427 82
rect 2527 86 2531 87
rect 2527 81 2531 82
rect 2655 86 2659 87
rect 2655 81 2659 82
rect 2775 86 2779 87
rect 2775 81 2779 82
rect 2895 86 2899 87
rect 2895 81 2899 82
rect 3015 86 3019 87
rect 3015 81 3019 82
rect 3135 86 3139 87
rect 3135 81 3139 82
rect 3247 86 3251 87
rect 3247 81 3251 82
rect 3359 86 3363 87
rect 3359 81 3363 82
rect 3471 86 3475 87
rect 3471 81 3475 82
rect 3583 86 3587 87
rect 3583 81 3587 82
rect 3687 86 3691 87
rect 3687 81 3691 82
rect 3791 86 3795 87
rect 3791 81 3795 82
rect 3895 86 3899 87
rect 3895 81 3899 82
rect 3991 86 3995 87
rect 3991 81 3995 82
<< m4c >>
rect 111 4062 115 4066
rect 327 4062 331 4066
rect 431 4062 435 4066
rect 535 4062 539 4066
rect 639 4062 643 4066
rect 743 4062 747 4066
rect 847 4062 851 4066
rect 951 4062 955 4066
rect 1055 4062 1059 4066
rect 1159 4062 1163 4066
rect 1263 4062 1267 4066
rect 1367 4062 1371 4066
rect 1471 4062 1475 4066
rect 2031 4062 2035 4066
rect 2071 4062 2075 4066
rect 2263 4062 2267 4066
rect 2367 4062 2371 4066
rect 2471 4062 2475 4066
rect 2575 4062 2579 4066
rect 2679 4062 2683 4066
rect 3991 4062 3995 4066
rect 111 3986 115 3990
rect 175 3986 179 3990
rect 327 3986 331 3990
rect 383 3986 387 3990
rect 431 3986 435 3990
rect 535 3986 539 3990
rect 591 3986 595 3990
rect 639 3986 643 3990
rect 743 3986 747 3990
rect 791 3986 795 3990
rect 847 3986 851 3990
rect 951 3986 955 3990
rect 983 3986 987 3990
rect 1055 3986 1059 3990
rect 1159 3986 1163 3990
rect 1167 3986 1171 3990
rect 1263 3986 1267 3990
rect 1343 3986 1347 3990
rect 1367 3986 1371 3990
rect 1471 3986 1475 3990
rect 1519 3986 1523 3990
rect 1703 3986 1707 3990
rect 2031 3986 2035 3990
rect 2071 3990 2075 3994
rect 2231 3990 2235 3994
rect 2263 3990 2267 3994
rect 111 3914 115 3918
rect 175 3914 179 3918
rect 359 3914 363 3918
rect 383 3914 387 3918
rect 551 3914 555 3918
rect 591 3914 595 3918
rect 735 3914 739 3918
rect 791 3914 795 3918
rect 535 3904 539 3908
rect 1075 3976 1079 3980
rect 1287 3979 1291 3980
rect 1287 3976 1291 3979
rect 1503 3976 1507 3980
rect 1775 3979 1779 3980
rect 1775 3976 1779 3979
rect 919 3914 923 3918
rect 983 3914 987 3918
rect 1087 3914 1091 3918
rect 1167 3914 1171 3918
rect 1247 3914 1251 3918
rect 1343 3914 1347 3918
rect 1399 3914 1403 3918
rect 863 3904 867 3908
rect 111 3842 115 3846
rect 359 3842 363 3846
rect 551 3842 555 3846
rect 583 3842 587 3846
rect 2367 3990 2371 3994
rect 2391 3990 2395 3994
rect 1519 3914 1523 3918
rect 1543 3914 1547 3918
rect 1679 3914 1683 3918
rect 1703 3914 1707 3918
rect 1815 3914 1819 3918
rect 1935 3914 1939 3918
rect 2031 3914 2035 3918
rect 2071 3918 2075 3922
rect 2223 3918 2227 3922
rect 2231 3918 2235 3922
rect 735 3842 739 3846
rect 887 3842 891 3846
rect 919 3842 923 3846
rect 1031 3842 1035 3846
rect 1087 3842 1091 3846
rect 1175 3842 1179 3846
rect 1247 3842 1251 3846
rect 1311 3842 1315 3846
rect 1399 3842 1403 3846
rect 1447 3842 1451 3846
rect 1543 3842 1547 3846
rect 1575 3842 1579 3846
rect 1679 3842 1683 3846
rect 1703 3842 1707 3846
rect 1815 3842 1819 3846
rect 1831 3842 1835 3846
rect 1935 3842 1939 3846
rect 111 3758 115 3762
rect 583 3758 587 3762
rect 599 3758 603 3762
rect 719 3758 723 3762
rect 735 3758 739 3762
rect 847 3758 851 3762
rect 887 3758 891 3762
rect 983 3758 987 3762
rect 1031 3758 1035 3762
rect 2471 3990 2475 3994
rect 2551 3990 2555 3994
rect 2575 3990 2579 3994
rect 2679 3990 2683 3994
rect 2703 3990 2707 3994
rect 2847 3990 2851 3994
rect 2983 3990 2987 3994
rect 3119 3990 3123 3994
rect 3247 3990 3251 3994
rect 3367 3990 3371 3994
rect 3479 3990 3483 3994
rect 3599 3990 3603 3994
rect 3719 3990 3723 3994
rect 3839 3990 3843 3994
rect 3991 3990 3995 3994
rect 2391 3918 2395 3922
rect 2455 3918 2459 3922
rect 2551 3918 2555 3922
rect 2671 3918 2675 3922
rect 2703 3918 2707 3922
rect 2031 3842 2035 3846
rect 2071 3846 2075 3850
rect 2191 3846 2195 3850
rect 2223 3846 2227 3850
rect 2455 3846 2459 3850
rect 2487 3846 2491 3850
rect 2071 3774 2075 3778
rect 2111 3774 2115 3778
rect 2191 3774 2195 3778
rect 1111 3758 1115 3762
rect 1175 3758 1179 3762
rect 1239 3758 1243 3762
rect 1311 3758 1315 3762
rect 1367 3758 1371 3762
rect 1447 3758 1451 3762
rect 1495 3758 1499 3762
rect 1575 3758 1579 3762
rect 1631 3758 1635 3762
rect 1703 3758 1707 3762
rect 1767 3758 1771 3762
rect 1831 3758 1835 3762
rect 1935 3758 1939 3762
rect 111 3682 115 3686
rect 471 3682 475 3686
rect 599 3682 603 3686
rect 615 3682 619 3686
rect 719 3682 723 3686
rect 759 3682 763 3686
rect 599 3664 603 3668
rect 111 3610 115 3614
rect 247 3610 251 3614
rect 375 3610 379 3614
rect 471 3610 475 3614
rect 519 3610 523 3614
rect 615 3610 619 3614
rect 679 3610 683 3614
rect 2031 3758 2035 3762
rect 2847 3918 2851 3922
rect 2879 3918 2883 3922
rect 2983 3918 2987 3922
rect 3071 3918 3075 3922
rect 3119 3918 3123 3922
rect 3247 3918 3251 3922
rect 3367 3918 3371 3922
rect 3415 3918 3419 3922
rect 3479 3918 3483 3922
rect 3583 3918 3587 3922
rect 3599 3918 3603 3922
rect 3719 3918 3723 3922
rect 3751 3918 3755 3922
rect 3839 3918 3843 3922
rect 3991 3918 3995 3922
rect 3055 3856 3059 3860
rect 3487 3856 3491 3860
rect 2671 3846 2675 3850
rect 2759 3846 2763 3850
rect 2879 3846 2883 3850
rect 2999 3846 3003 3850
rect 3071 3846 3075 3850
rect 3215 3846 3219 3850
rect 3247 3846 3251 3850
rect 3407 3846 3411 3850
rect 3415 3846 3419 3850
rect 3583 3846 3587 3850
rect 3751 3846 3755 3850
rect 3895 3846 3899 3850
rect 3991 3846 3995 3850
rect 2335 3774 2339 3778
rect 2487 3774 2491 3778
rect 2559 3774 2563 3778
rect 2759 3774 2763 3778
rect 2775 3774 2779 3778
rect 2975 3774 2979 3778
rect 2999 3774 3003 3778
rect 3159 3774 3163 3778
rect 3215 3774 3219 3778
rect 3327 3774 3331 3778
rect 3407 3774 3411 3778
rect 3479 3774 3483 3778
rect 3583 3774 3587 3778
rect 2071 3690 2075 3694
rect 2111 3690 2115 3694
rect 2255 3690 2259 3694
rect 2335 3690 2339 3694
rect 2439 3690 2443 3694
rect 2559 3690 2563 3694
rect 2623 3690 2627 3694
rect 2775 3690 2779 3694
rect 2815 3690 2819 3694
rect 847 3682 851 3686
rect 903 3682 907 3686
rect 983 3682 987 3686
rect 1047 3682 1051 3686
rect 1111 3682 1115 3686
rect 1191 3682 1195 3686
rect 1239 3682 1243 3686
rect 1335 3682 1339 3686
rect 1367 3682 1371 3686
rect 1479 3682 1483 3686
rect 1495 3682 1499 3686
rect 1631 3682 1635 3686
rect 1767 3682 1771 3686
rect 2031 3682 2035 3686
rect 911 3664 915 3668
rect 759 3610 763 3614
rect 847 3610 851 3614
rect 903 3610 907 3614
rect 1023 3610 1027 3614
rect 1047 3610 1051 3614
rect 111 3526 115 3530
rect 151 3526 155 3530
rect 247 3526 251 3530
rect 263 3526 267 3530
rect 375 3526 379 3530
rect 399 3526 403 3530
rect 111 3454 115 3458
rect 151 3454 155 3458
rect 263 3454 267 3458
rect 399 3454 403 3458
rect 519 3526 523 3530
rect 543 3526 547 3530
rect 679 3526 683 3530
rect 687 3526 691 3530
rect 831 3526 835 3530
rect 847 3526 851 3530
rect 967 3526 971 3530
rect 1023 3526 1027 3530
rect 1191 3610 1195 3614
rect 1207 3610 1211 3614
rect 1335 3610 1339 3614
rect 1391 3610 1395 3614
rect 1479 3610 1483 3614
rect 1575 3610 1579 3614
rect 1767 3610 1771 3614
rect 1935 3610 1939 3614
rect 2031 3610 2035 3614
rect 1175 3552 1179 3556
rect 1463 3552 1467 3556
rect 1095 3526 1099 3530
rect 1207 3526 1211 3530
rect 1223 3526 1227 3530
rect 1343 3526 1347 3530
rect 1391 3526 1395 3530
rect 1463 3526 1467 3530
rect 1575 3526 1579 3530
rect 423 3454 427 3458
rect 543 3454 547 3458
rect 687 3454 691 3458
rect 743 3454 747 3458
rect 831 3454 835 3458
rect 967 3454 971 3458
rect 1071 3454 1075 3458
rect 1095 3454 1099 3458
rect 1223 3454 1227 3458
rect 1343 3454 1347 3458
rect 1399 3454 1403 3458
rect 111 3358 115 3362
rect 151 3358 155 3362
rect 1463 3454 1467 3458
rect 1583 3526 1587 3530
rect 3623 3774 3627 3778
rect 3751 3774 3755 3778
rect 3767 3774 3771 3778
rect 3895 3774 3899 3778
rect 3991 3774 3995 3778
rect 2975 3690 2979 3694
rect 3007 3690 3011 3694
rect 3159 3690 3163 3694
rect 3199 3690 3203 3694
rect 3327 3690 3331 3694
rect 3391 3690 3395 3694
rect 3479 3690 3483 3694
rect 3583 3690 3587 3694
rect 3623 3690 3627 3694
rect 3767 3690 3771 3694
rect 3895 3690 3899 3694
rect 3991 3690 3995 3694
rect 2071 3606 2075 3610
rect 2111 3606 2115 3610
rect 2255 3606 2259 3610
rect 2359 3606 2363 3610
rect 2439 3606 2443 3610
rect 2583 3606 2587 3610
rect 2623 3606 2627 3610
rect 2799 3606 2803 3610
rect 2815 3606 2819 3610
rect 3007 3606 3011 3610
rect 3199 3606 3203 3610
rect 3215 3606 3219 3610
rect 3391 3606 3395 3610
rect 3431 3606 3435 3610
rect 3583 3606 3587 3610
rect 3991 3606 3995 3610
rect 1711 3526 1715 3530
rect 1767 3526 1771 3530
rect 1935 3526 1939 3530
rect 2031 3526 2035 3530
rect 2071 3530 2075 3534
rect 2359 3530 2363 3534
rect 2439 3530 2443 3534
rect 2575 3530 2579 3534
rect 2583 3530 2587 3534
rect 2703 3530 2707 3534
rect 2799 3530 2803 3534
rect 2831 3530 2835 3534
rect 2951 3530 2955 3534
rect 3007 3530 3011 3534
rect 3071 3530 3075 3534
rect 3199 3530 3203 3534
rect 3215 3530 3219 3534
rect 3327 3530 3331 3534
rect 3431 3530 3435 3534
rect 3991 3530 3995 3534
rect 1583 3454 1587 3458
rect 1711 3454 1715 3458
rect 2031 3454 2035 3458
rect 2071 3458 2075 3462
rect 2359 3458 2363 3462
rect 2439 3458 2443 3462
rect 2463 3458 2467 3462
rect 2567 3458 2571 3462
rect 2575 3458 2579 3462
rect 2671 3458 2675 3462
rect 2703 3458 2707 3462
rect 2775 3458 2779 3462
rect 319 3358 323 3362
rect 423 3358 427 3362
rect 527 3358 531 3362
rect 743 3358 747 3362
rect 959 3358 963 3362
rect 1071 3358 1075 3362
rect 1167 3358 1171 3362
rect 1367 3358 1371 3362
rect 1399 3358 1403 3362
rect 1559 3358 1563 3362
rect 1751 3358 1755 3362
rect 1935 3358 1939 3362
rect 2031 3358 2035 3362
rect 2071 3358 2075 3362
rect 2359 3358 2363 3362
rect 2439 3358 2443 3362
rect 2463 3358 2467 3362
rect 111 3278 115 3282
rect 151 3278 155 3282
rect 311 3278 315 3282
rect 319 3278 323 3282
rect 479 3278 483 3282
rect 527 3278 531 3282
rect 655 3278 659 3282
rect 743 3278 747 3282
rect 847 3278 851 3282
rect 959 3278 963 3282
rect 1039 3278 1043 3282
rect 1167 3278 1171 3282
rect 1231 3278 1235 3282
rect 1367 3278 1371 3282
rect 1431 3278 1435 3282
rect 1559 3278 1563 3282
rect 1631 3278 1635 3282
rect 1751 3278 1755 3282
rect 1831 3278 1835 3282
rect 1935 3278 1939 3282
rect 2543 3358 2547 3362
rect 2567 3358 2571 3362
rect 2831 3458 2835 3462
rect 2879 3458 2883 3462
rect 2951 3458 2955 3462
rect 2983 3458 2987 3462
rect 3071 3458 3075 3462
rect 3087 3458 3091 3462
rect 3191 3458 3195 3462
rect 3199 3458 3203 3462
rect 3327 3458 3331 3462
rect 3991 3458 3995 3462
rect 2647 3358 2651 3362
rect 2671 3358 2675 3362
rect 2751 3358 2755 3362
rect 2775 3358 2779 3362
rect 2855 3358 2859 3362
rect 2879 3358 2883 3362
rect 2959 3358 2963 3362
rect 2983 3358 2987 3362
rect 3087 3358 3091 3362
rect 3191 3358 3195 3362
rect 3991 3358 3995 3362
rect 2071 3286 2075 3290
rect 2439 3286 2443 3290
rect 2527 3286 2531 3290
rect 2543 3286 2547 3290
rect 2031 3278 2035 3282
rect 111 3202 115 3206
rect 311 3202 315 3206
rect 479 3202 483 3206
rect 623 3202 627 3206
rect 655 3202 659 3206
rect 759 3202 763 3206
rect 847 3202 851 3206
rect 903 3202 907 3206
rect 1039 3202 1043 3206
rect 743 3192 747 3196
rect 1055 3202 1059 3206
rect 1207 3202 1211 3206
rect 1231 3202 1235 3206
rect 1047 3192 1051 3196
rect 111 3130 115 3134
rect 599 3130 603 3134
rect 623 3130 627 3134
rect 703 3130 707 3134
rect 759 3130 763 3134
rect 807 3130 811 3134
rect 903 3130 907 3134
rect 911 3130 915 3134
rect 1039 3130 1043 3134
rect 1055 3130 1059 3134
rect 1351 3202 1355 3206
rect 1431 3202 1435 3206
rect 1503 3202 1507 3206
rect 1631 3202 1635 3206
rect 1655 3202 1659 3206
rect 2631 3286 2635 3290
rect 2647 3286 2651 3290
rect 2735 3286 2739 3290
rect 2751 3286 2755 3290
rect 2839 3286 2843 3290
rect 2855 3286 2859 3290
rect 2071 3214 2075 3218
rect 2399 3214 2403 3218
rect 2527 3214 2531 3218
rect 2719 3224 2723 3228
rect 2943 3286 2947 3290
rect 2959 3286 2963 3290
rect 3047 3286 3051 3290
rect 3151 3286 3155 3290
rect 3255 3286 3259 3290
rect 3991 3286 3995 3290
rect 3015 3224 3019 3228
rect 2551 3214 2555 3218
rect 2631 3214 2635 3218
rect 2695 3214 2699 3218
rect 2735 3214 2739 3218
rect 2839 3214 2843 3218
rect 2943 3214 2947 3218
rect 2975 3214 2979 3218
rect 3047 3214 3051 3218
rect 3111 3214 3115 3218
rect 3151 3214 3155 3218
rect 1807 3202 1811 3206
rect 1831 3202 1835 3206
rect 1935 3202 1939 3206
rect 2031 3202 2035 3206
rect 1183 3130 1187 3134
rect 1207 3130 1211 3134
rect 1351 3130 1355 3134
rect 1359 3130 1363 3134
rect 1503 3130 1507 3134
rect 1551 3130 1555 3134
rect 111 3050 115 3054
rect 311 3050 315 3054
rect 415 3050 419 3054
rect 527 3050 531 3054
rect 599 3050 603 3054
rect 639 3050 643 3054
rect 111 2970 115 2974
rect 151 2970 155 2974
rect 271 2970 275 2974
rect 311 2970 315 2974
rect 415 2970 419 2974
rect 431 2970 435 2974
rect 527 2970 531 2974
rect 1655 3130 1659 3134
rect 1751 3130 1755 3134
rect 1807 3130 1811 3134
rect 1935 3130 1939 3134
rect 3247 3214 3251 3218
rect 3255 3214 3259 3218
rect 3391 3214 3395 3218
rect 3991 3214 3995 3218
rect 2959 3195 2963 3196
rect 2959 3192 2963 3195
rect 3399 3192 3403 3196
rect 2031 3130 2035 3134
rect 2071 3130 2075 3134
rect 2111 3130 2115 3134
rect 2343 3130 2347 3134
rect 2399 3130 2403 3134
rect 703 3050 707 3054
rect 751 3050 755 3054
rect 807 3050 811 3054
rect 863 3050 867 3054
rect 911 3050 915 3054
rect 975 3050 979 3054
rect 1039 3050 1043 3054
rect 1095 3050 1099 3054
rect 1183 3050 1187 3054
rect 1215 3050 1219 3054
rect 1335 3050 1339 3054
rect 1359 3050 1363 3054
rect 1551 3050 1555 3054
rect 1751 3050 1755 3054
rect 1935 3050 1939 3054
rect 2031 3050 2035 3054
rect 2071 3054 2075 3058
rect 2111 3054 2115 3058
rect 607 2970 611 2974
rect 639 2970 643 2974
rect 751 2970 755 2974
rect 783 2970 787 2974
rect 863 2970 867 2974
rect 959 2970 963 2974
rect 975 2970 979 2974
rect 1095 2970 1099 2974
rect 1135 2970 1139 2974
rect 111 2886 115 2890
rect 151 2886 155 2890
rect 271 2886 275 2890
rect 287 2886 291 2890
rect 431 2886 435 2890
rect 447 2886 451 2890
rect 111 2802 115 2806
rect 151 2802 155 2806
rect 599 2886 603 2890
rect 607 2886 611 2890
rect 759 2886 763 2890
rect 783 2886 787 2890
rect 927 2886 931 2890
rect 959 2886 963 2890
rect 2551 3130 2555 3134
rect 2583 3130 2587 3134
rect 2695 3130 2699 3134
rect 2799 3130 2803 3134
rect 2839 3130 2843 3134
rect 2975 3130 2979 3134
rect 2999 3130 3003 3134
rect 3111 3130 3115 3134
rect 3191 3130 3195 3134
rect 3247 3130 3251 3134
rect 2263 3054 2267 3058
rect 2343 3054 2347 3058
rect 2455 3054 2459 3058
rect 2583 3054 2587 3058
rect 2655 3054 2659 3058
rect 3375 3130 3379 3134
rect 3391 3130 3395 3134
rect 3567 3130 3571 3134
rect 3991 3130 3995 3134
rect 2799 3054 2803 3058
rect 2855 3054 2859 3058
rect 2999 3054 3003 3058
rect 3055 3054 3059 3058
rect 3191 3054 3195 3058
rect 3255 3054 3259 3058
rect 3375 3054 3379 3058
rect 3455 3054 3459 3058
rect 3567 3054 3571 3058
rect 3655 3054 3659 3058
rect 3991 3054 3995 3058
rect 2071 2982 2075 2986
rect 2111 2982 2115 2986
rect 2263 2982 2267 2986
rect 2359 2982 2363 2986
rect 1215 2970 1219 2974
rect 1303 2970 1307 2974
rect 1335 2970 1339 2974
rect 1471 2970 1475 2974
rect 1647 2970 1651 2974
rect 2031 2970 2035 2974
rect 1103 2886 1107 2890
rect 1135 2886 1139 2890
rect 1287 2886 1291 2890
rect 1303 2886 1307 2890
rect 1471 2886 1475 2890
rect 1479 2886 1483 2890
rect 1647 2886 1651 2890
rect 1671 2886 1675 2890
rect 287 2802 291 2806
rect 319 2802 323 2806
rect 447 2802 451 2806
rect 503 2802 507 2806
rect 111 2726 115 2730
rect 151 2726 155 2730
rect 183 2726 187 2730
rect 319 2726 323 2730
rect 383 2726 387 2730
rect 111 2646 115 2650
rect 183 2646 187 2650
rect 599 2802 603 2806
rect 687 2802 691 2806
rect 759 2802 763 2806
rect 871 2802 875 2806
rect 927 2802 931 2806
rect 1055 2802 1059 2806
rect 1103 2802 1107 2806
rect 1239 2802 1243 2806
rect 1287 2802 1291 2806
rect 1431 2802 1435 2806
rect 1479 2802 1483 2806
rect 2455 2982 2459 2986
rect 2607 2982 2611 2986
rect 2655 2982 2659 2986
rect 2847 2982 2851 2986
rect 2855 2982 2859 2986
rect 2071 2902 2075 2906
rect 2111 2902 2115 2906
rect 2279 2902 2283 2906
rect 2359 2902 2363 2906
rect 2031 2886 2035 2890
rect 1631 2802 1635 2806
rect 1671 2802 1675 2806
rect 503 2726 507 2730
rect 583 2726 587 2730
rect 687 2726 691 2730
rect 783 2726 787 2730
rect 871 2726 875 2730
rect 983 2726 987 2730
rect 3055 2982 3059 2986
rect 3079 2982 3083 2986
rect 3255 2982 3259 2986
rect 3303 2982 3307 2986
rect 3455 2982 3459 2986
rect 3535 2982 3539 2986
rect 3655 2982 3659 2986
rect 3767 2982 3771 2986
rect 3991 2982 3995 2986
rect 2487 2902 2491 2906
rect 2607 2902 2611 2906
rect 2695 2902 2699 2906
rect 2847 2902 2851 2906
rect 2903 2902 2907 2906
rect 3079 2902 3083 2906
rect 3111 2902 3115 2906
rect 3303 2902 3307 2906
rect 3495 2902 3499 2906
rect 3535 2902 3539 2906
rect 3687 2902 3691 2906
rect 3767 2902 3771 2906
rect 3879 2902 3883 2906
rect 3991 2902 3995 2906
rect 2071 2818 2075 2822
rect 2111 2818 2115 2822
rect 2143 2818 2147 2822
rect 1831 2802 1835 2806
rect 2031 2802 2035 2806
rect 1055 2726 1059 2730
rect 1199 2726 1203 2730
rect 1239 2726 1243 2730
rect 1415 2726 1419 2730
rect 1431 2726 1435 2730
rect 1631 2726 1635 2730
rect 1639 2726 1643 2730
rect 1831 2726 1835 2730
rect 1871 2726 1875 2730
rect 255 2646 259 2650
rect 383 2646 387 2650
rect 423 2646 427 2650
rect 583 2646 587 2650
rect 599 2646 603 2650
rect 775 2646 779 2650
rect 783 2646 787 2650
rect 959 2646 963 2650
rect 983 2646 987 2650
rect 1151 2646 1155 2650
rect 1199 2646 1203 2650
rect 1343 2646 1347 2650
rect 1415 2646 1419 2650
rect 1535 2646 1539 2650
rect 1639 2646 1643 2650
rect 2071 2734 2075 2738
rect 2111 2734 2115 2738
rect 2143 2734 2147 2738
rect 2031 2726 2035 2730
rect 1727 2646 1731 2650
rect 1871 2646 1875 2650
rect 1927 2646 1931 2650
rect 111 2570 115 2574
rect 255 2570 259 2574
rect 319 2570 323 2574
rect 423 2570 427 2574
rect 535 2570 539 2574
rect 599 2570 603 2574
rect 743 2570 747 2574
rect 775 2570 779 2574
rect 111 2498 115 2502
rect 279 2498 283 2502
rect 319 2498 323 2502
rect 951 2570 955 2574
rect 959 2570 963 2574
rect 1151 2570 1155 2574
rect 1159 2570 1163 2574
rect 1343 2570 1347 2574
rect 1359 2570 1363 2574
rect 1535 2570 1539 2574
rect 1559 2570 1563 2574
rect 439 2498 443 2502
rect 535 2498 539 2502
rect 607 2498 611 2502
rect 743 2498 747 2502
rect 783 2498 787 2502
rect 951 2498 955 2502
rect 959 2498 963 2502
rect 111 2418 115 2422
rect 279 2418 283 2422
rect 327 2418 331 2422
rect 439 2418 443 2422
rect 471 2418 475 2422
rect 607 2418 611 2422
rect 623 2418 627 2422
rect 1127 2498 1131 2502
rect 1159 2498 1163 2502
rect 1295 2498 1299 2502
rect 1359 2498 1363 2502
rect 1727 2570 1731 2574
rect 1759 2570 1763 2574
rect 2279 2818 2283 2822
rect 2319 2818 2323 2822
rect 2487 2818 2491 2822
rect 2503 2818 2507 2822
rect 2695 2818 2699 2822
rect 2887 2818 2891 2822
rect 2903 2818 2907 2822
rect 3079 2818 3083 2822
rect 3111 2818 3115 2822
rect 3263 2818 3267 2822
rect 3303 2818 3307 2822
rect 3439 2818 3443 2822
rect 3495 2818 3499 2822
rect 3615 2818 3619 2822
rect 3687 2818 3691 2822
rect 3791 2818 3795 2822
rect 3879 2818 3883 2822
rect 2279 2734 2283 2738
rect 2319 2734 2323 2738
rect 2455 2734 2459 2738
rect 2503 2734 2507 2738
rect 3991 2818 3995 2822
rect 2639 2734 2643 2738
rect 2695 2734 2699 2738
rect 2815 2734 2819 2738
rect 2887 2734 2891 2738
rect 2983 2734 2987 2738
rect 3079 2734 3083 2738
rect 3143 2734 3147 2738
rect 3263 2734 3267 2738
rect 3303 2734 3307 2738
rect 3439 2734 3443 2738
rect 3463 2734 3467 2738
rect 3615 2734 3619 2738
rect 3623 2734 3627 2738
rect 3791 2734 3795 2738
rect 3991 2734 3995 2738
rect 2031 2646 2035 2650
rect 2071 2650 2075 2654
rect 2111 2650 2115 2654
rect 2263 2650 2267 2654
rect 2279 2650 2283 2654
rect 1927 2570 1931 2574
rect 1935 2570 1939 2574
rect 2031 2570 2035 2574
rect 2071 2570 2075 2574
rect 2111 2570 2115 2574
rect 1463 2498 1467 2502
rect 1559 2498 1563 2502
rect 1623 2498 1627 2502
rect 1759 2498 1763 2502
rect 1791 2498 1795 2502
rect 783 2418 787 2422
rect 943 2418 947 2422
rect 959 2418 963 2422
rect 1095 2418 1099 2422
rect 1127 2418 1131 2422
rect 1247 2418 1251 2422
rect 1295 2418 1299 2422
rect 111 2338 115 2342
rect 327 2338 331 2342
rect 359 2338 363 2342
rect 471 2338 475 2342
rect 495 2338 499 2342
rect 623 2338 627 2342
rect 639 2338 643 2342
rect 783 2338 787 2342
rect 935 2338 939 2342
rect 943 2338 947 2342
rect 1391 2418 1395 2422
rect 1463 2418 1467 2422
rect 1535 2418 1539 2422
rect 1623 2418 1627 2422
rect 1671 2418 1675 2422
rect 1935 2498 1939 2502
rect 1791 2418 1795 2422
rect 1815 2418 1819 2422
rect 2431 2650 2435 2654
rect 2455 2650 2459 2654
rect 2599 2650 2603 2654
rect 2639 2650 2643 2654
rect 2751 2650 2755 2654
rect 2815 2650 2819 2654
rect 2895 2650 2899 2654
rect 2983 2650 2987 2654
rect 3039 2650 3043 2654
rect 2263 2570 2267 2574
rect 2271 2570 2275 2574
rect 2431 2570 2435 2574
rect 2447 2570 2451 2574
rect 2599 2570 2603 2574
rect 2615 2570 2619 2574
rect 2031 2498 2035 2502
rect 2071 2486 2075 2490
rect 2111 2486 2115 2490
rect 2271 2486 2275 2490
rect 2447 2486 2451 2490
rect 1935 2418 1939 2422
rect 2031 2418 2035 2422
rect 1087 2338 1091 2342
rect 1095 2338 1099 2342
rect 1247 2338 1251 2342
rect 1391 2338 1395 2342
rect 1415 2338 1419 2342
rect 111 2254 115 2258
rect 239 2254 243 2258
rect 359 2254 363 2258
rect 391 2254 395 2258
rect 495 2254 499 2258
rect 551 2254 555 2258
rect 639 2254 643 2258
rect 711 2254 715 2258
rect 783 2254 787 2258
rect 871 2254 875 2258
rect 935 2254 939 2258
rect 1031 2254 1035 2258
rect 1087 2254 1091 2258
rect 111 2170 115 2174
rect 151 2170 155 2174
rect 239 2170 243 2174
rect 319 2170 323 2174
rect 391 2170 395 2174
rect 511 2170 515 2174
rect 551 2170 555 2174
rect 703 2170 707 2174
rect 711 2170 715 2174
rect 871 2170 875 2174
rect 895 2170 899 2174
rect 1535 2338 1539 2342
rect 1591 2338 1595 2342
rect 1671 2338 1675 2342
rect 1775 2338 1779 2342
rect 1815 2338 1819 2342
rect 1935 2338 1939 2342
rect 1191 2254 1195 2258
rect 1247 2254 1251 2258
rect 1359 2254 1363 2258
rect 1415 2254 1419 2258
rect 1527 2254 1531 2258
rect 1591 2254 1595 2258
rect 1695 2254 1699 2258
rect 1031 2170 1035 2174
rect 1087 2170 1091 2174
rect 1191 2170 1195 2174
rect 1279 2170 1283 2174
rect 1359 2170 1363 2174
rect 3143 2650 3147 2654
rect 3175 2650 3179 2654
rect 3303 2650 3307 2654
rect 3311 2650 3315 2654
rect 3455 2650 3459 2654
rect 3463 2650 3467 2654
rect 3623 2650 3627 2654
rect 3991 2650 3995 2654
rect 3127 2592 3131 2596
rect 3527 2592 3531 2596
rect 2751 2570 2755 2574
rect 2767 2570 2771 2574
rect 2895 2570 2899 2574
rect 2911 2570 2915 2574
rect 3039 2570 3043 2574
rect 3047 2570 3051 2574
rect 3175 2570 3179 2574
rect 3183 2570 3187 2574
rect 3311 2570 3315 2574
rect 3319 2570 3323 2574
rect 3455 2570 3459 2574
rect 3991 2570 3995 2574
rect 2615 2486 2619 2490
rect 2623 2486 2627 2490
rect 2743 2486 2747 2490
rect 2767 2486 2771 2490
rect 2871 2486 2875 2490
rect 2071 2402 2075 2406
rect 2487 2402 2491 2406
rect 2599 2402 2603 2406
rect 2623 2402 2627 2406
rect 2727 2402 2731 2406
rect 2743 2402 2747 2406
rect 2031 2338 2035 2342
rect 2071 2318 2075 2322
rect 2111 2318 2115 2322
rect 2223 2318 2227 2322
rect 2359 2318 2363 2322
rect 2487 2318 2491 2322
rect 2511 2318 2515 2322
rect 2599 2318 2603 2322
rect 1775 2254 1779 2258
rect 1935 2254 1939 2258
rect 2031 2254 2035 2258
rect 1463 2170 1467 2174
rect 1527 2170 1531 2174
rect 111 2090 115 2094
rect 151 2090 155 2094
rect 303 2090 307 2094
rect 319 2090 323 2094
rect 479 2090 483 2094
rect 511 2090 515 2094
rect 663 2090 667 2094
rect 703 2090 707 2094
rect 847 2090 851 2094
rect 895 2090 899 2094
rect 1039 2090 1043 2094
rect 1087 2090 1091 2094
rect 111 2010 115 2014
rect 151 2010 155 2014
rect 303 2010 307 2014
rect 479 2010 483 2014
rect 487 2010 491 2014
rect 663 2010 667 2014
rect 687 2010 691 2014
rect 847 2010 851 2014
rect 895 2010 899 2014
rect 2911 2486 2915 2490
rect 3015 2486 3019 2490
rect 3047 2486 3051 2490
rect 3159 2486 3163 2490
rect 3183 2486 3187 2490
rect 3311 2486 3315 2490
rect 3319 2486 3323 2490
rect 3463 2486 3467 2490
rect 3615 2486 3619 2490
rect 3767 2486 3771 2490
rect 3895 2486 3899 2490
rect 3991 2486 3995 2490
rect 2871 2402 2875 2406
rect 2879 2402 2883 2406
rect 3015 2402 3019 2406
rect 3055 2402 3059 2406
rect 3159 2402 3163 2406
rect 3247 2402 3251 2406
rect 3311 2402 3315 2406
rect 3455 2402 3459 2406
rect 3463 2402 3467 2406
rect 3615 2402 3619 2406
rect 3679 2402 3683 2406
rect 3767 2402 3771 2406
rect 3895 2402 3899 2406
rect 3991 2402 3995 2406
rect 2671 2318 2675 2322
rect 2727 2318 2731 2322
rect 2847 2318 2851 2322
rect 2879 2318 2883 2322
rect 3039 2318 3043 2322
rect 3055 2318 3059 2322
rect 2071 2238 2075 2242
rect 2111 2238 2115 2242
rect 2223 2238 2227 2242
rect 2279 2238 2283 2242
rect 2359 2238 2363 2242
rect 3247 2318 3251 2322
rect 3455 2318 3459 2322
rect 3463 2318 3467 2322
rect 3679 2318 3683 2322
rect 3687 2318 3691 2322
rect 3895 2318 3899 2322
rect 2479 2238 2483 2242
rect 2511 2238 2515 2242
rect 2671 2238 2675 2242
rect 2679 2238 2683 2242
rect 2847 2238 2851 2242
rect 2879 2238 2883 2242
rect 3039 2238 3043 2242
rect 3079 2238 3083 2242
rect 1655 2170 1659 2174
rect 1695 2170 1699 2174
rect 1847 2170 1851 2174
rect 2031 2170 2035 2174
rect 2071 2158 2075 2162
rect 2111 2158 2115 2162
rect 2143 2158 2147 2162
rect 2279 2158 2283 2162
rect 2319 2158 2323 2162
rect 1239 2090 1243 2094
rect 1279 2090 1283 2094
rect 1447 2090 1451 2094
rect 1463 2090 1467 2094
rect 1655 2090 1659 2094
rect 1663 2090 1667 2094
rect 1039 2010 1043 2014
rect 1103 2010 1107 2014
rect 1239 2010 1243 2014
rect 1311 2010 1315 2014
rect 1447 2010 1451 2014
rect 1847 2090 1851 2094
rect 1879 2090 1883 2094
rect 2031 2090 2035 2094
rect 1527 2010 1531 2014
rect 1663 2010 1667 2014
rect 1743 2010 1747 2014
rect 1879 2010 1883 2014
rect 1935 2010 1939 2014
rect 111 1926 115 1930
rect 151 1926 155 1930
rect 271 1926 275 1930
rect 303 1926 307 1930
rect 407 1926 411 1930
rect 487 1926 491 1930
rect 543 1926 547 1930
rect 679 1926 683 1930
rect 687 1926 691 1930
rect 111 1846 115 1850
rect 151 1846 155 1850
rect 271 1846 275 1850
rect 287 1846 291 1850
rect 407 1846 411 1850
rect 447 1846 451 1850
rect 543 1846 547 1850
rect 599 1846 603 1850
rect 823 1926 827 1930
rect 895 1926 899 1930
rect 983 1926 987 1930
rect 1103 1926 1107 1930
rect 1159 1926 1163 1930
rect 1311 1926 1315 1930
rect 1343 1926 1347 1930
rect 1527 1926 1531 1930
rect 1543 1926 1547 1930
rect 2071 2074 2075 2078
rect 2143 2074 2147 2078
rect 2207 2074 2211 2078
rect 2479 2158 2483 2162
rect 2495 2158 2499 2162
rect 2679 2158 2683 2162
rect 3247 2238 3251 2242
rect 3279 2238 3283 2242
rect 3463 2238 3467 2242
rect 3487 2238 3491 2242
rect 3687 2238 3691 2242
rect 3703 2238 3707 2242
rect 3063 2224 3067 2228
rect 3259 2227 3263 2228
rect 3259 2224 3263 2227
rect 2863 2158 2867 2162
rect 2879 2158 2883 2162
rect 3039 2158 3043 2162
rect 3079 2158 3083 2162
rect 3215 2158 3219 2162
rect 3279 2158 3283 2162
rect 3391 2158 3395 2162
rect 2319 2074 2323 2078
rect 2391 2074 2395 2078
rect 2495 2074 2499 2078
rect 2575 2074 2579 2078
rect 2679 2074 2683 2078
rect 2759 2074 2763 2078
rect 2863 2074 2867 2078
rect 2031 2010 2035 2014
rect 2071 1990 2075 1994
rect 2207 1990 2211 1994
rect 2279 1990 2283 1994
rect 1743 1926 1747 1930
rect 1751 1926 1755 1930
rect 1935 1926 1939 1930
rect 2031 1926 2035 1930
rect 679 1846 683 1850
rect 751 1846 755 1850
rect 823 1846 827 1850
rect 919 1846 923 1850
rect 983 1846 987 1850
rect 1103 1846 1107 1850
rect 1159 1846 1163 1850
rect 1303 1846 1307 1850
rect 1343 1846 1347 1850
rect 1511 1846 1515 1850
rect 1543 1846 1547 1850
rect 1735 1846 1739 1850
rect 1751 1846 1755 1850
rect 1935 1846 1939 1850
rect 111 1766 115 1770
rect 151 1766 155 1770
rect 207 1766 211 1770
rect 287 1766 291 1770
rect 383 1766 387 1770
rect 447 1766 451 1770
rect 567 1766 571 1770
rect 599 1766 603 1770
rect 751 1766 755 1770
rect 919 1766 923 1770
rect 935 1766 939 1770
rect 1103 1766 1107 1770
rect 1111 1766 1115 1770
rect 1279 1766 1283 1770
rect 1303 1766 1307 1770
rect 1455 1766 1459 1770
rect 1511 1766 1515 1770
rect 1631 1766 1635 1770
rect 1735 1766 1739 1770
rect 111 1694 115 1698
rect 207 1694 211 1698
rect 303 1694 307 1698
rect 383 1694 387 1698
rect 535 1694 539 1698
rect 567 1694 571 1698
rect 751 1694 755 1698
rect 767 1694 771 1698
rect 935 1694 939 1698
rect 983 1694 987 1698
rect 1263 1747 1267 1748
rect 1263 1744 1267 1747
rect 1111 1694 1115 1698
rect 1191 1694 1195 1698
rect 1279 1694 1283 1698
rect 1383 1694 1387 1698
rect 1455 1694 1459 1698
rect 1567 1694 1571 1698
rect 1631 1694 1635 1698
rect 2391 1990 2395 1994
rect 2463 1990 2467 1994
rect 2575 1990 2579 1994
rect 2639 1990 2643 1994
rect 2935 2074 2939 2078
rect 3039 2074 3043 2078
rect 3103 2074 3107 2078
rect 3487 2158 3491 2162
rect 3567 2158 3571 2162
rect 3703 2158 3707 2162
rect 3991 2318 3995 2322
rect 3895 2238 3899 2242
rect 3991 2238 3995 2242
rect 3743 2158 3747 2162
rect 3895 2158 3899 2162
rect 3215 2074 3219 2078
rect 3263 2074 3267 2078
rect 3391 2074 3395 2078
rect 3423 2074 3427 2078
rect 3567 2074 3571 2078
rect 3583 2074 3587 2078
rect 3743 2074 3747 2078
rect 3751 2074 3755 2078
rect 2759 1990 2763 1994
rect 2815 1990 2819 1994
rect 2935 1990 2939 1994
rect 2983 1990 2987 1994
rect 3103 1990 3107 1994
rect 3151 1990 3155 1994
rect 3263 1990 3267 1994
rect 3311 1990 3315 1994
rect 3423 1990 3427 1994
rect 3463 1990 3467 1994
rect 3583 1990 3587 1994
rect 3615 1990 3619 1994
rect 3991 2158 3995 2162
rect 3895 2074 3899 2078
rect 3991 2074 3995 2078
rect 3751 1990 3755 1994
rect 3767 1990 3771 1994
rect 3895 1990 3899 1994
rect 2071 1910 2075 1914
rect 2279 1910 2283 1914
rect 2407 1910 2411 1914
rect 2463 1910 2467 1914
rect 2639 1910 2643 1914
rect 2655 1910 2659 1914
rect 2815 1910 2819 1914
rect 2887 1910 2891 1914
rect 2983 1910 2987 1914
rect 3103 1910 3107 1914
rect 3151 1910 3155 1914
rect 3311 1910 3315 1914
rect 3463 1910 3467 1914
rect 3511 1910 3515 1914
rect 3615 1910 3619 1914
rect 3711 1910 3715 1914
rect 3767 1910 3771 1914
rect 2031 1846 2035 1850
rect 2071 1838 2075 1842
rect 2111 1838 2115 1842
rect 2383 1838 2387 1842
rect 2407 1838 2411 1842
rect 1935 1766 1939 1770
rect 2031 1766 2035 1770
rect 2071 1766 2075 1770
rect 2111 1766 2115 1770
rect 1743 1744 1747 1748
rect 2647 1838 2651 1842
rect 2655 1838 2659 1842
rect 2887 1838 2891 1842
rect 3095 1838 3099 1842
rect 3103 1838 3107 1842
rect 2287 1766 2291 1770
rect 2383 1766 2387 1770
rect 2495 1766 2499 1770
rect 2647 1766 2651 1770
rect 2711 1766 2715 1770
rect 2887 1766 2891 1770
rect 2919 1766 2923 1770
rect 3287 1838 3291 1842
rect 3311 1838 3315 1842
rect 3455 1838 3459 1842
rect 3511 1838 3515 1842
rect 3991 1990 3995 1994
rect 3895 1910 3899 1914
rect 3991 1910 3995 1914
rect 3615 1838 3619 1842
rect 3711 1838 3715 1842
rect 3767 1838 3771 1842
rect 3095 1766 3099 1770
rect 3119 1766 3123 1770
rect 3287 1766 3291 1770
rect 3319 1766 3323 1770
rect 1743 1694 1747 1698
rect 1927 1694 1931 1698
rect 2031 1694 2035 1698
rect 2071 1686 2075 1690
rect 2111 1686 2115 1690
rect 2239 1686 2243 1690
rect 2287 1686 2291 1690
rect 2383 1686 2387 1690
rect 111 1618 115 1622
rect 303 1618 307 1622
rect 399 1618 403 1622
rect 535 1618 539 1622
rect 575 1618 579 1622
rect 751 1618 755 1622
rect 767 1618 771 1622
rect 935 1618 939 1622
rect 983 1618 987 1622
rect 1111 1618 1115 1622
rect 1191 1618 1195 1622
rect 1279 1618 1283 1622
rect 1383 1618 1387 1622
rect 1447 1618 1451 1622
rect 111 1538 115 1542
rect 399 1538 403 1542
rect 503 1538 507 1542
rect 575 1538 579 1542
rect 615 1538 619 1542
rect 735 1538 739 1542
rect 751 1538 755 1542
rect 855 1538 859 1542
rect 935 1538 939 1542
rect 967 1538 971 1542
rect 1567 1618 1571 1622
rect 1607 1618 1611 1622
rect 1743 1618 1747 1622
rect 1767 1618 1771 1622
rect 1927 1618 1931 1622
rect 1935 1618 1939 1622
rect 1079 1538 1083 1542
rect 1111 1538 1115 1542
rect 1199 1538 1203 1542
rect 1279 1538 1283 1542
rect 1319 1538 1323 1542
rect 1439 1538 1443 1542
rect 1447 1538 1451 1542
rect 2031 1618 2035 1622
rect 2071 1602 2075 1606
rect 2111 1602 2115 1606
rect 2167 1602 2171 1606
rect 2495 1686 2499 1690
rect 2519 1686 2523 1690
rect 2655 1686 2659 1690
rect 2711 1686 2715 1690
rect 2239 1602 2243 1606
rect 2287 1602 2291 1606
rect 2383 1602 2387 1606
rect 2407 1602 2411 1606
rect 2519 1602 2523 1606
rect 2527 1602 2531 1606
rect 2791 1686 2795 1690
rect 2919 1686 2923 1690
rect 2927 1686 2931 1690
rect 3455 1766 3459 1770
rect 3895 1838 3899 1842
rect 3991 1838 3995 1842
rect 3511 1766 3515 1770
rect 3615 1766 3619 1770
rect 3703 1766 3707 1770
rect 3767 1766 3771 1770
rect 3895 1766 3899 1770
rect 3991 1766 3995 1770
rect 3063 1686 3067 1690
rect 3119 1686 3123 1690
rect 2647 1602 2651 1606
rect 2655 1602 2659 1606
rect 2767 1602 2771 1606
rect 2791 1602 2795 1606
rect 3207 1686 3211 1690
rect 3319 1686 3323 1690
rect 3351 1686 3355 1690
rect 3511 1686 3515 1690
rect 3703 1686 3707 1690
rect 3895 1686 3899 1690
rect 3991 1686 3995 1690
rect 2887 1602 2891 1606
rect 2927 1602 2931 1606
rect 3007 1602 3011 1606
rect 3063 1602 3067 1606
rect 3127 1602 3131 1606
rect 3207 1602 3211 1606
rect 3255 1602 3259 1606
rect 1559 1538 1563 1542
rect 1607 1538 1611 1542
rect 1767 1538 1771 1542
rect 1935 1538 1939 1542
rect 2031 1538 2035 1542
rect 2071 1522 2075 1526
rect 2167 1522 2171 1526
rect 2287 1522 2291 1526
rect 2351 1522 2355 1526
rect 2407 1522 2411 1526
rect 2463 1522 2467 1526
rect 2527 1522 2531 1526
rect 111 1454 115 1458
rect 503 1454 507 1458
rect 583 1454 587 1458
rect 615 1454 619 1458
rect 687 1454 691 1458
rect 735 1454 739 1458
rect 791 1454 795 1458
rect 855 1454 859 1458
rect 895 1454 899 1458
rect 967 1454 971 1458
rect 999 1454 1003 1458
rect 1079 1454 1083 1458
rect 1103 1454 1107 1458
rect 1199 1454 1203 1458
rect 1207 1454 1211 1458
rect 111 1374 115 1378
rect 551 1374 555 1378
rect 583 1374 587 1378
rect 655 1374 659 1378
rect 687 1374 691 1378
rect 759 1374 763 1378
rect 791 1374 795 1378
rect 863 1374 867 1378
rect 895 1374 899 1378
rect 975 1374 979 1378
rect 999 1374 1003 1378
rect 1087 1374 1091 1378
rect 1103 1374 1107 1378
rect 1311 1454 1315 1458
rect 1319 1454 1323 1458
rect 1415 1454 1419 1458
rect 1199 1374 1203 1378
rect 1207 1374 1211 1378
rect 1311 1374 1315 1378
rect 1439 1454 1443 1458
rect 1519 1454 1523 1458
rect 1559 1454 1563 1458
rect 2031 1454 2035 1458
rect 2447 1464 2451 1468
rect 2575 1522 2579 1526
rect 2647 1522 2651 1526
rect 2695 1522 2699 1526
rect 2071 1438 2075 1442
rect 2343 1438 2347 1442
rect 2351 1438 2355 1442
rect 2447 1438 2451 1442
rect 2463 1438 2467 1442
rect 2567 1438 2571 1442
rect 2575 1438 2579 1442
rect 2767 1522 2771 1526
rect 2815 1522 2819 1526
rect 2887 1522 2891 1526
rect 3351 1602 3355 1606
rect 3991 1602 3995 1606
rect 2927 1522 2931 1526
rect 2767 1464 2771 1468
rect 2695 1438 2699 1442
rect 2815 1438 2819 1442
rect 2839 1438 2843 1442
rect 3007 1522 3011 1526
rect 3047 1522 3051 1526
rect 3127 1522 3131 1526
rect 3167 1522 3171 1526
rect 3255 1522 3259 1526
rect 3287 1522 3291 1526
rect 3407 1522 3411 1526
rect 3991 1522 3995 1526
rect 2927 1438 2931 1442
rect 2991 1438 2995 1442
rect 3047 1438 3051 1442
rect 3143 1438 3147 1442
rect 3167 1438 3171 1442
rect 3287 1438 3291 1442
rect 3303 1438 3307 1442
rect 1415 1374 1419 1378
rect 1431 1374 1435 1378
rect 1519 1374 1523 1378
rect 1551 1374 1555 1378
rect 2031 1374 2035 1378
rect 2071 1358 2075 1362
rect 2287 1358 2291 1362
rect 2343 1358 2347 1362
rect 111 1298 115 1302
rect 343 1298 347 1302
rect 463 1298 467 1302
rect 551 1298 555 1302
rect 599 1298 603 1302
rect 655 1298 659 1302
rect 743 1298 747 1302
rect 759 1298 763 1302
rect 863 1298 867 1302
rect 903 1298 907 1302
rect 975 1298 979 1302
rect 1063 1298 1067 1302
rect 1087 1298 1091 1302
rect 1199 1298 1203 1302
rect 1231 1298 1235 1302
rect 111 1226 115 1230
rect 183 1226 187 1230
rect 343 1226 347 1230
rect 351 1226 355 1230
rect 463 1226 467 1230
rect 535 1226 539 1230
rect 599 1226 603 1230
rect 727 1226 731 1230
rect 743 1226 747 1230
rect 903 1226 907 1230
rect 919 1226 923 1230
rect 1063 1226 1067 1230
rect 1103 1226 1107 1230
rect 1311 1298 1315 1302
rect 1407 1298 1411 1302
rect 1431 1298 1435 1302
rect 1551 1298 1555 1302
rect 1583 1298 1587 1302
rect 1231 1226 1235 1230
rect 1287 1226 1291 1230
rect 1407 1226 1411 1230
rect 2031 1298 2035 1302
rect 2407 1358 2411 1362
rect 2447 1358 2451 1362
rect 2543 1358 2547 1362
rect 2567 1358 2571 1362
rect 2695 1358 2699 1362
rect 2839 1358 2843 1362
rect 2855 1358 2859 1362
rect 2991 1358 2995 1362
rect 3015 1358 3019 1362
rect 3143 1358 3147 1362
rect 3183 1358 3187 1362
rect 3407 1438 3411 1442
rect 3471 1438 3475 1442
rect 3647 1438 3651 1442
rect 3823 1438 3827 1442
rect 3991 1438 3995 1442
rect 3303 1358 3307 1362
rect 3351 1358 3355 1362
rect 3471 1358 3475 1362
rect 3519 1358 3523 1362
rect 3647 1358 3651 1362
rect 3687 1358 3691 1362
rect 2071 1278 2075 1282
rect 2127 1278 2131 1282
rect 2287 1278 2291 1282
rect 2295 1278 2299 1282
rect 2407 1278 2411 1282
rect 2479 1278 2483 1282
rect 2543 1278 2547 1282
rect 2679 1278 2683 1282
rect 2695 1278 2699 1282
rect 2855 1278 2859 1282
rect 2879 1278 2883 1282
rect 3015 1278 3019 1282
rect 3071 1278 3075 1282
rect 1471 1226 1475 1230
rect 1583 1226 1587 1230
rect 1655 1226 1659 1230
rect 1839 1226 1843 1230
rect 2031 1226 2035 1230
rect 2071 1194 2075 1198
rect 2111 1194 2115 1198
rect 2127 1194 2131 1198
rect 111 1146 115 1150
rect 151 1146 155 1150
rect 183 1146 187 1150
rect 303 1146 307 1150
rect 351 1146 355 1150
rect 495 1146 499 1150
rect 535 1146 539 1150
rect 703 1146 707 1150
rect 727 1146 731 1150
rect 911 1146 915 1150
rect 919 1146 923 1150
rect 1103 1146 1107 1150
rect 1119 1146 1123 1150
rect 111 1066 115 1070
rect 151 1066 155 1070
rect 279 1066 283 1070
rect 303 1066 307 1070
rect 447 1066 451 1070
rect 495 1066 499 1070
rect 623 1066 627 1070
rect 703 1066 707 1070
rect 799 1066 803 1070
rect 911 1066 915 1070
rect 967 1066 971 1070
rect 1287 1146 1291 1150
rect 1319 1146 1323 1150
rect 1471 1146 1475 1150
rect 1519 1146 1523 1150
rect 1655 1146 1659 1150
rect 1719 1146 1723 1150
rect 1839 1146 1843 1150
rect 1119 1066 1123 1070
rect 1127 1066 1131 1070
rect 1919 1146 1923 1150
rect 2031 1146 2035 1150
rect 2247 1194 2251 1198
rect 2295 1194 2299 1198
rect 2407 1194 2411 1198
rect 2479 1194 2483 1198
rect 2559 1194 2563 1198
rect 2679 1194 2683 1198
rect 2703 1194 2707 1198
rect 2863 1194 2867 1198
rect 2071 1118 2075 1122
rect 2111 1118 2115 1122
rect 2247 1118 2251 1122
rect 2303 1118 2307 1122
rect 2407 1118 2411 1122
rect 2511 1118 2515 1122
rect 2559 1118 2563 1122
rect 2879 1194 2883 1198
rect 3183 1278 3187 1282
rect 3247 1278 3251 1282
rect 3351 1278 3355 1282
rect 3415 1278 3419 1282
rect 3519 1278 3523 1282
rect 3583 1278 3587 1282
rect 3687 1278 3691 1282
rect 3751 1278 3755 1282
rect 3823 1358 3827 1362
rect 3855 1358 3859 1362
rect 3991 1358 3995 1362
rect 3855 1278 3859 1282
rect 3895 1278 3899 1282
rect 3991 1278 3995 1282
rect 3039 1194 3043 1198
rect 3071 1194 3075 1198
rect 3239 1194 3243 1198
rect 3247 1194 3251 1198
rect 3415 1194 3419 1198
rect 3455 1194 3459 1198
rect 3583 1194 3587 1198
rect 3687 1194 3691 1198
rect 3751 1194 3755 1198
rect 3895 1194 3899 1198
rect 3991 1194 3995 1198
rect 2703 1118 2707 1122
rect 2863 1118 2867 1122
rect 2895 1118 2899 1122
rect 3039 1118 3043 1122
rect 3087 1118 3091 1122
rect 3239 1118 3243 1122
rect 3287 1118 3291 1122
rect 3455 1118 3459 1122
rect 3495 1118 3499 1122
rect 3687 1118 3691 1122
rect 3703 1118 3707 1122
rect 3895 1118 3899 1122
rect 1279 1066 1283 1070
rect 1319 1066 1323 1070
rect 1423 1066 1427 1070
rect 1519 1066 1523 1070
rect 1559 1066 1563 1070
rect 1695 1066 1699 1070
rect 1719 1066 1723 1070
rect 1823 1066 1827 1070
rect 1919 1066 1923 1070
rect 1935 1066 1939 1070
rect 2031 1066 2035 1070
rect 2071 1030 2075 1034
rect 111 982 115 986
rect 151 982 155 986
rect 279 982 283 986
rect 287 982 291 986
rect 447 982 451 986
rect 471 982 475 986
rect 623 982 627 986
rect 671 982 675 986
rect 799 982 803 986
rect 871 982 875 986
rect 967 982 971 986
rect 1079 982 1083 986
rect 1127 982 1131 986
rect 655 968 659 972
rect 935 971 939 972
rect 935 968 939 971
rect 2111 1030 2115 1034
rect 2303 1030 2307 1034
rect 2319 1030 2323 1034
rect 2487 1030 2491 1034
rect 2511 1030 2515 1034
rect 2663 1030 2667 1034
rect 2703 1030 2707 1034
rect 2847 1030 2851 1034
rect 1279 982 1283 986
rect 1287 982 1291 986
rect 1423 982 1427 986
rect 1495 982 1499 986
rect 1559 982 1563 986
rect 1695 982 1699 986
rect 1703 982 1707 986
rect 1823 982 1827 986
rect 1911 982 1915 986
rect 1935 982 1939 986
rect 2031 982 2035 986
rect 111 902 115 906
rect 151 902 155 906
rect 287 902 291 906
rect 319 902 323 906
rect 471 902 475 906
rect 519 902 523 906
rect 671 902 675 906
rect 727 902 731 906
rect 871 902 875 906
rect 935 902 939 906
rect 111 818 115 822
rect 151 818 155 822
rect 263 818 267 822
rect 319 818 323 822
rect 367 818 371 822
rect 479 818 483 822
rect 519 818 523 822
rect 591 818 595 822
rect 711 818 715 822
rect 727 818 731 822
rect 855 818 859 822
rect 935 818 939 822
rect 1079 902 1083 906
rect 1143 902 1147 906
rect 1287 902 1291 906
rect 1335 902 1339 906
rect 1495 902 1499 906
rect 1527 902 1531 906
rect 1703 902 1707 906
rect 1719 902 1723 906
rect 1911 902 1915 906
rect 2071 954 2075 958
rect 2151 954 2155 958
rect 2287 954 2291 958
rect 2319 954 2323 958
rect 2431 954 2435 958
rect 2487 954 2491 958
rect 2591 954 2595 958
rect 2663 954 2667 958
rect 2895 1030 2899 1034
rect 3039 1030 3043 1034
rect 3087 1030 3091 1034
rect 3247 1030 3251 1034
rect 3287 1030 3291 1034
rect 3463 1030 3467 1034
rect 3495 1030 3499 1034
rect 3687 1030 3691 1034
rect 3703 1030 3707 1034
rect 3991 1118 3995 1122
rect 3895 1030 3899 1034
rect 2759 954 2763 958
rect 2847 954 2851 958
rect 2935 954 2939 958
rect 3039 954 3043 958
rect 3119 954 3123 958
rect 2031 902 2035 906
rect 2071 870 2075 874
rect 2111 870 2115 874
rect 2151 870 2155 874
rect 2239 870 2243 874
rect 1031 818 1035 822
rect 1143 818 1147 822
rect 1239 818 1243 822
rect 1335 818 1339 822
rect 1471 818 1475 822
rect 1527 818 1531 822
rect 1711 818 1715 822
rect 1719 818 1723 822
rect 1911 818 1915 822
rect 1935 818 1939 822
rect 2031 818 2035 822
rect 111 742 115 746
rect 263 742 267 746
rect 367 742 371 746
rect 423 742 427 746
rect 479 742 483 746
rect 527 742 531 746
rect 591 742 595 746
rect 639 742 643 746
rect 711 742 715 746
rect 759 742 763 746
rect 855 742 859 746
rect 879 742 883 746
rect 1007 742 1011 746
rect 1031 742 1035 746
rect 1143 742 1147 746
rect 1239 742 1243 746
rect 1287 742 1291 746
rect 1447 742 1451 746
rect 1471 742 1475 746
rect 1615 742 1619 746
rect 1711 742 1715 746
rect 1783 742 1787 746
rect 111 658 115 662
rect 423 658 427 662
rect 527 658 531 662
rect 591 658 595 662
rect 639 658 643 662
rect 695 658 699 662
rect 759 658 763 662
rect 807 658 811 662
rect 879 658 883 662
rect 919 658 923 662
rect 1007 658 1011 662
rect 1031 658 1035 662
rect 1143 658 1147 662
rect 2071 798 2075 802
rect 2111 798 2115 802
rect 2287 870 2291 874
rect 2407 870 2411 874
rect 2431 870 2435 874
rect 2575 870 2579 874
rect 2591 870 2595 874
rect 2751 870 2755 874
rect 2759 870 2763 874
rect 3991 1030 3995 1034
rect 3247 954 3251 958
rect 3311 954 3315 958
rect 3463 954 3467 958
rect 3511 954 3515 958
rect 3687 954 3691 958
rect 3711 954 3715 958
rect 3895 954 3899 958
rect 2935 870 2939 874
rect 3119 870 3123 874
rect 3311 870 3315 874
rect 3511 870 3515 874
rect 3711 870 3715 874
rect 3991 954 3995 958
rect 3895 870 3899 874
rect 2239 798 2243 802
rect 2391 798 2395 802
rect 3991 870 3995 874
rect 2407 798 2411 802
rect 2575 798 2579 802
rect 2679 798 2683 802
rect 2751 798 2755 802
rect 2935 798 2939 802
rect 2951 798 2955 802
rect 3119 798 3123 802
rect 3199 798 3203 802
rect 1935 742 1939 746
rect 2031 742 2035 746
rect 2071 718 2075 722
rect 2111 718 2115 722
rect 2327 718 2331 722
rect 2391 718 2395 722
rect 1263 658 1267 662
rect 1287 658 1291 662
rect 1383 658 1387 662
rect 1447 658 1451 662
rect 1503 658 1507 662
rect 1615 658 1619 662
rect 1623 658 1627 662
rect 1783 658 1787 662
rect 1935 658 1939 662
rect 2031 658 2035 662
rect 111 578 115 582
rect 591 578 595 582
rect 663 578 667 582
rect 695 578 699 582
rect 775 578 779 582
rect 807 578 811 582
rect 895 578 899 582
rect 919 578 923 582
rect 1023 578 1027 582
rect 1031 578 1035 582
rect 1143 578 1147 582
rect 1159 578 1163 582
rect 1263 578 1267 582
rect 1303 578 1307 582
rect 1383 578 1387 582
rect 1447 578 1451 582
rect 1503 578 1507 582
rect 3311 798 3315 802
rect 3439 798 3443 802
rect 3511 798 3515 802
rect 3671 798 3675 802
rect 3711 798 3715 802
rect 3895 798 3899 802
rect 2551 718 2555 722
rect 2679 718 2683 722
rect 2775 718 2779 722
rect 2951 718 2955 722
rect 2991 718 2995 722
rect 2071 642 2075 646
rect 2111 642 2115 646
rect 2127 642 2131 646
rect 3199 718 3203 722
rect 3207 718 3211 722
rect 3415 718 3419 722
rect 3439 718 3443 722
rect 3623 718 3627 722
rect 3671 718 3675 722
rect 3991 798 3995 802
rect 3831 718 3835 722
rect 3895 718 3899 722
rect 2295 642 2299 646
rect 2327 642 2331 646
rect 2455 642 2459 646
rect 2551 642 2555 646
rect 2615 642 2619 646
rect 2775 642 2779 646
rect 2783 642 2787 646
rect 2951 642 2955 646
rect 2991 642 2995 646
rect 3127 642 3131 646
rect 1591 578 1595 582
rect 1623 578 1627 582
rect 1735 578 1739 582
rect 1879 578 1883 582
rect 2031 578 2035 582
rect 2071 562 2075 566
rect 2127 562 2131 566
rect 2295 562 2299 566
rect 2303 562 2307 566
rect 2447 562 2451 566
rect 2455 562 2459 566
rect 111 490 115 494
rect 535 490 539 494
rect 639 490 643 494
rect 663 490 667 494
rect 743 490 747 494
rect 775 490 779 494
rect 847 490 851 494
rect 895 490 899 494
rect 967 490 971 494
rect 1023 490 1027 494
rect 1103 490 1107 494
rect 1159 490 1163 494
rect 1255 490 1259 494
rect 1303 490 1307 494
rect 111 414 115 418
rect 495 414 499 418
rect 535 414 539 418
rect 631 414 635 418
rect 639 414 643 418
rect 743 414 747 418
rect 767 414 771 418
rect 847 414 851 418
rect 911 414 915 418
rect 967 414 971 418
rect 1415 490 1419 494
rect 1447 490 1451 494
rect 1591 490 1595 494
rect 1735 490 1739 494
rect 1775 490 1779 494
rect 1879 490 1883 494
rect 1935 490 1939 494
rect 1239 472 1243 476
rect 1599 472 1603 476
rect 1047 414 1051 418
rect 1103 414 1107 418
rect 1183 414 1187 418
rect 1255 414 1259 418
rect 1319 414 1323 418
rect 111 330 115 334
rect 335 330 339 334
rect 463 330 467 334
rect 495 330 499 334
rect 607 330 611 334
rect 631 330 635 334
rect 767 330 771 334
rect 911 330 915 334
rect 111 250 115 254
rect 151 250 155 254
rect 279 250 283 254
rect 335 250 339 254
rect 431 250 435 254
rect 463 250 467 254
rect 599 250 603 254
rect 607 250 611 254
rect 767 250 771 254
rect 783 250 787 254
rect 943 330 947 334
rect 1415 414 1419 418
rect 1447 414 1451 418
rect 1575 414 1579 418
rect 1591 414 1595 418
rect 1703 414 1707 418
rect 1775 414 1779 418
rect 1831 414 1835 418
rect 2031 490 2035 494
rect 2591 562 2595 566
rect 2615 562 2619 566
rect 2735 562 2739 566
rect 2783 562 2787 566
rect 3207 642 3211 646
rect 3303 642 3307 646
rect 3415 642 3419 646
rect 3487 642 3491 646
rect 3623 642 3627 646
rect 3679 642 3683 646
rect 3831 642 3835 646
rect 3879 642 3883 646
rect 3991 718 3995 722
rect 2879 562 2883 566
rect 2951 562 2955 566
rect 3031 562 3035 566
rect 3127 562 3131 566
rect 3183 562 3187 566
rect 3303 562 3307 566
rect 3335 562 3339 566
rect 2071 482 2075 486
rect 2303 482 2307 486
rect 2447 482 2451 486
rect 2511 482 2515 486
rect 2591 482 2595 486
rect 2615 482 2619 486
rect 2735 482 2739 486
rect 3167 504 3171 508
rect 2863 482 2867 486
rect 2879 482 2883 486
rect 3487 562 3491 566
rect 3495 562 3499 566
rect 3655 562 3659 566
rect 3679 562 3683 566
rect 3991 642 3995 646
rect 3823 562 3827 566
rect 3879 562 3883 566
rect 3567 504 3571 508
rect 3007 482 3011 486
rect 3031 482 3035 486
rect 3159 482 3163 486
rect 3183 482 3187 486
rect 3319 482 3323 486
rect 3335 482 3339 486
rect 3479 482 3483 486
rect 3495 482 3499 486
rect 3647 482 3651 486
rect 3655 482 3659 486
rect 1935 414 1939 418
rect 2031 414 2035 418
rect 2071 398 2075 402
rect 2511 398 2515 402
rect 2591 398 2595 402
rect 2615 398 2619 402
rect 2695 398 2699 402
rect 2735 398 2739 402
rect 2815 398 2819 402
rect 2863 398 2867 402
rect 1047 330 1051 334
rect 1127 330 1131 334
rect 1183 330 1187 334
rect 1311 330 1315 334
rect 1319 330 1323 334
rect 1447 330 1451 334
rect 1503 330 1507 334
rect 1575 330 1579 334
rect 1703 330 1707 334
rect 943 250 947 254
rect 975 250 979 254
rect 1127 250 1131 254
rect 1175 250 1179 254
rect 1311 250 1315 254
rect 1375 250 1379 254
rect 1831 330 1835 334
rect 1903 330 1907 334
rect 1935 330 1939 334
rect 2031 330 2035 334
rect 1503 250 1507 254
rect 1583 250 1587 254
rect 1703 250 1707 254
rect 1799 250 1803 254
rect 111 154 115 158
rect 151 154 155 158
rect 255 154 259 158
rect 279 154 283 158
rect 359 154 363 158
rect 431 154 435 158
rect 471 154 475 158
rect 599 154 603 158
rect 607 154 611 158
rect 743 154 747 158
rect 783 154 787 158
rect 879 154 883 158
rect 975 154 979 158
rect 1015 154 1019 158
rect 2071 326 2075 330
rect 3991 562 3995 566
rect 3823 482 3827 486
rect 3991 482 3995 486
rect 2959 398 2963 402
rect 3007 398 3011 402
rect 3119 398 3123 402
rect 3159 398 3163 402
rect 3303 398 3307 402
rect 3319 398 3323 402
rect 3479 398 3483 402
rect 3503 398 3507 402
rect 3647 398 3651 402
rect 3711 398 3715 402
rect 3823 398 3827 402
rect 3895 398 3899 402
rect 3991 398 3995 402
rect 2111 326 2115 330
rect 2271 326 2275 330
rect 2455 326 2459 330
rect 2591 326 2595 330
rect 2631 326 2635 330
rect 2695 326 2699 330
rect 2807 326 2811 330
rect 2815 326 2819 330
rect 2959 326 2963 330
rect 2999 326 3003 330
rect 3119 326 3123 330
rect 3215 326 3219 330
rect 3303 326 3307 330
rect 3439 326 3443 330
rect 3503 326 3507 330
rect 1903 250 1907 254
rect 2031 250 2035 254
rect 2071 254 2075 258
rect 2111 254 2115 258
rect 2271 254 2275 258
rect 2455 254 2459 258
rect 3679 326 3683 330
rect 3711 326 3715 330
rect 3895 326 3899 330
rect 2983 312 2987 316
rect 3511 312 3515 316
rect 2471 254 2475 258
rect 2631 254 2635 258
rect 2687 254 2691 258
rect 1151 154 1155 158
rect 1175 154 1179 158
rect 1279 154 1283 158
rect 1375 154 1379 158
rect 1399 154 1403 158
rect 1519 154 1523 158
rect 1583 154 1587 158
rect 1647 154 1651 158
rect 1775 154 1779 158
rect 1799 154 1803 158
rect 2031 154 2035 158
rect 2071 154 2075 158
rect 2111 154 2115 158
rect 2807 254 2811 258
rect 2903 254 2907 258
rect 2999 254 3003 258
rect 3111 254 3115 258
rect 3215 254 3219 258
rect 3319 254 3323 258
rect 3439 254 3443 258
rect 3519 254 3523 258
rect 3679 254 3683 258
rect 3991 326 3995 330
rect 3719 254 3723 258
rect 3895 254 3899 258
rect 2215 154 2219 158
rect 2271 154 2275 158
rect 2319 154 2323 158
rect 2423 154 2427 158
rect 2471 154 2475 158
rect 2527 154 2531 158
rect 2655 154 2659 158
rect 2687 154 2691 158
rect 2775 154 2779 158
rect 2895 154 2899 158
rect 2903 154 2907 158
rect 3015 154 3019 158
rect 3111 154 3115 158
rect 3135 154 3139 158
rect 3247 154 3251 158
rect 3319 154 3323 158
rect 3359 154 3363 158
rect 3471 154 3475 158
rect 3519 154 3523 158
rect 3583 154 3587 158
rect 3687 154 3691 158
rect 3719 154 3723 158
rect 3991 254 3995 258
rect 3791 154 3795 158
rect 3895 154 3899 158
rect 3991 154 3995 158
rect 111 82 115 86
rect 151 82 155 86
rect 255 82 259 86
rect 359 82 363 86
rect 471 82 475 86
rect 607 82 611 86
rect 743 82 747 86
rect 879 82 883 86
rect 1015 82 1019 86
rect 1151 82 1155 86
rect 1279 82 1283 86
rect 1399 82 1403 86
rect 1519 82 1523 86
rect 1647 82 1651 86
rect 1775 82 1779 86
rect 2031 82 2035 86
rect 2071 82 2075 86
rect 2111 82 2115 86
rect 2215 82 2219 86
rect 2319 82 2323 86
rect 2423 82 2427 86
rect 2527 82 2531 86
rect 2655 82 2659 86
rect 2775 82 2779 86
rect 2895 82 2899 86
rect 3015 82 3019 86
rect 3135 82 3139 86
rect 3247 82 3251 86
rect 3359 82 3363 86
rect 3471 82 3475 86
rect 3583 82 3587 86
rect 3687 82 3691 86
rect 3791 82 3795 86
rect 3895 82 3899 86
rect 3991 82 3995 86
<< m4 >>
rect 84 4061 85 4067
rect 91 4066 2043 4067
rect 91 4062 111 4066
rect 115 4062 327 4066
rect 331 4062 431 4066
rect 435 4062 535 4066
rect 539 4062 639 4066
rect 643 4062 743 4066
rect 747 4062 847 4066
rect 851 4062 951 4066
rect 955 4062 1055 4066
rect 1059 4062 1159 4066
rect 1163 4062 1263 4066
rect 1267 4062 1367 4066
rect 1371 4062 1471 4066
rect 1475 4062 2031 4066
rect 2035 4062 2043 4066
rect 91 4061 2043 4062
rect 2049 4066 4022 4067
rect 2049 4062 2071 4066
rect 2075 4062 2263 4066
rect 2267 4062 2367 4066
rect 2371 4062 2471 4066
rect 2475 4062 2575 4066
rect 2579 4062 2679 4066
rect 2683 4062 3991 4066
rect 3995 4062 4022 4066
rect 2049 4061 4022 4062
rect 2054 3994 4034 3995
rect 2054 3991 2071 3994
rect 96 3985 97 3991
rect 103 3990 2055 3991
rect 103 3986 111 3990
rect 115 3986 175 3990
rect 179 3986 327 3990
rect 331 3986 383 3990
rect 387 3986 431 3990
rect 435 3986 535 3990
rect 539 3986 591 3990
rect 595 3986 639 3990
rect 643 3986 743 3990
rect 747 3986 791 3990
rect 795 3986 847 3990
rect 851 3986 951 3990
rect 955 3986 983 3990
rect 987 3986 1055 3990
rect 1059 3986 1159 3990
rect 1163 3986 1167 3990
rect 1171 3986 1263 3990
rect 1267 3986 1343 3990
rect 1347 3986 1367 3990
rect 1371 3986 1471 3990
rect 1475 3986 1519 3990
rect 1523 3986 1703 3990
rect 1707 3986 2031 3990
rect 2035 3986 2055 3990
rect 103 3985 2055 3986
rect 2061 3990 2071 3991
rect 2075 3990 2231 3994
rect 2235 3990 2263 3994
rect 2267 3990 2367 3994
rect 2371 3990 2391 3994
rect 2395 3990 2471 3994
rect 2475 3990 2551 3994
rect 2555 3990 2575 3994
rect 2579 3990 2679 3994
rect 2683 3990 2703 3994
rect 2707 3990 2847 3994
rect 2851 3990 2983 3994
rect 2987 3990 3119 3994
rect 3123 3990 3247 3994
rect 3251 3990 3367 3994
rect 3371 3990 3479 3994
rect 3483 3990 3599 3994
rect 3603 3990 3719 3994
rect 3723 3990 3839 3994
rect 3843 3990 3991 3994
rect 3995 3990 4034 3994
rect 2061 3989 4034 3990
rect 2061 3985 2062 3989
rect 1074 3980 1080 3981
rect 1286 3980 1292 3981
rect 1074 3976 1075 3980
rect 1079 3976 1287 3980
rect 1291 3976 1292 3980
rect 1074 3975 1080 3976
rect 1286 3975 1292 3976
rect 1502 3980 1508 3981
rect 1774 3980 1780 3981
rect 1502 3976 1503 3980
rect 1507 3976 1775 3980
rect 1779 3976 1780 3980
rect 1502 3975 1508 3976
rect 1774 3975 1780 3976
rect 2042 3922 4022 3923
rect 2042 3919 2071 3922
rect 84 3913 85 3919
rect 91 3918 2043 3919
rect 91 3914 111 3918
rect 115 3914 175 3918
rect 179 3914 359 3918
rect 363 3914 383 3918
rect 387 3914 551 3918
rect 555 3914 591 3918
rect 595 3914 735 3918
rect 739 3914 791 3918
rect 795 3914 919 3918
rect 923 3914 983 3918
rect 987 3914 1087 3918
rect 1091 3914 1167 3918
rect 1171 3914 1247 3918
rect 1251 3914 1343 3918
rect 1347 3914 1399 3918
rect 1403 3914 1519 3918
rect 1523 3914 1543 3918
rect 1547 3914 1679 3918
rect 1683 3914 1703 3918
rect 1707 3914 1815 3918
rect 1819 3914 1935 3918
rect 1939 3914 2031 3918
rect 2035 3914 2043 3918
rect 91 3913 2043 3914
rect 2049 3918 2071 3919
rect 2075 3918 2223 3922
rect 2227 3918 2231 3922
rect 2235 3918 2391 3922
rect 2395 3918 2455 3922
rect 2459 3918 2551 3922
rect 2555 3918 2671 3922
rect 2675 3918 2703 3922
rect 2707 3918 2847 3922
rect 2851 3918 2879 3922
rect 2883 3918 2983 3922
rect 2987 3918 3071 3922
rect 3075 3918 3119 3922
rect 3123 3918 3247 3922
rect 3251 3918 3367 3922
rect 3371 3918 3415 3922
rect 3419 3918 3479 3922
rect 3483 3918 3583 3922
rect 3587 3918 3599 3922
rect 3603 3918 3719 3922
rect 3723 3918 3751 3922
rect 3755 3918 3839 3922
rect 3843 3918 3991 3922
rect 3995 3918 4022 3922
rect 2049 3917 4022 3918
rect 2049 3913 2050 3917
rect 534 3908 540 3909
rect 862 3908 868 3909
rect 534 3904 535 3908
rect 539 3904 863 3908
rect 867 3904 868 3908
rect 534 3903 540 3904
rect 862 3903 868 3904
rect 3054 3860 3060 3861
rect 3486 3860 3492 3861
rect 3054 3856 3055 3860
rect 3059 3856 3487 3860
rect 3491 3856 3492 3860
rect 3054 3855 3060 3856
rect 3486 3855 3492 3856
rect 2054 3850 4034 3851
rect 2054 3847 2071 3850
rect 96 3841 97 3847
rect 103 3846 2055 3847
rect 103 3842 111 3846
rect 115 3842 359 3846
rect 363 3842 551 3846
rect 555 3842 583 3846
rect 587 3842 735 3846
rect 739 3842 887 3846
rect 891 3842 919 3846
rect 923 3842 1031 3846
rect 1035 3842 1087 3846
rect 1091 3842 1175 3846
rect 1179 3842 1247 3846
rect 1251 3842 1311 3846
rect 1315 3842 1399 3846
rect 1403 3842 1447 3846
rect 1451 3842 1543 3846
rect 1547 3842 1575 3846
rect 1579 3842 1679 3846
rect 1683 3842 1703 3846
rect 1707 3842 1815 3846
rect 1819 3842 1831 3846
rect 1835 3842 1935 3846
rect 1939 3842 2031 3846
rect 2035 3842 2055 3846
rect 103 3841 2055 3842
rect 2061 3846 2071 3847
rect 2075 3846 2191 3850
rect 2195 3846 2223 3850
rect 2227 3846 2455 3850
rect 2459 3846 2487 3850
rect 2491 3846 2671 3850
rect 2675 3846 2759 3850
rect 2763 3846 2879 3850
rect 2883 3846 2999 3850
rect 3003 3846 3071 3850
rect 3075 3846 3215 3850
rect 3219 3846 3247 3850
rect 3251 3846 3407 3850
rect 3411 3846 3415 3850
rect 3419 3846 3583 3850
rect 3587 3846 3751 3850
rect 3755 3846 3895 3850
rect 3899 3846 3991 3850
rect 3995 3846 4034 3850
rect 2061 3845 4034 3846
rect 2061 3841 2062 3845
rect 2042 3773 2043 3779
rect 2049 3778 4015 3779
rect 2049 3774 2071 3778
rect 2075 3774 2111 3778
rect 2115 3774 2191 3778
rect 2195 3774 2335 3778
rect 2339 3774 2487 3778
rect 2491 3774 2559 3778
rect 2563 3774 2759 3778
rect 2763 3774 2775 3778
rect 2779 3774 2975 3778
rect 2979 3774 2999 3778
rect 3003 3774 3159 3778
rect 3163 3774 3215 3778
rect 3219 3774 3327 3778
rect 3331 3774 3407 3778
rect 3411 3774 3479 3778
rect 3483 3774 3583 3778
rect 3587 3774 3623 3778
rect 3627 3774 3751 3778
rect 3755 3774 3767 3778
rect 3771 3774 3895 3778
rect 3899 3774 3991 3778
rect 3995 3774 4015 3778
rect 2049 3773 4015 3774
rect 4021 3773 4022 3779
rect 84 3757 85 3763
rect 91 3762 2043 3763
rect 91 3758 111 3762
rect 115 3758 583 3762
rect 587 3758 599 3762
rect 603 3758 719 3762
rect 723 3758 735 3762
rect 739 3758 847 3762
rect 851 3758 887 3762
rect 891 3758 983 3762
rect 987 3758 1031 3762
rect 1035 3758 1111 3762
rect 1115 3758 1175 3762
rect 1179 3758 1239 3762
rect 1243 3758 1311 3762
rect 1315 3758 1367 3762
rect 1371 3758 1447 3762
rect 1451 3758 1495 3762
rect 1499 3758 1575 3762
rect 1579 3758 1631 3762
rect 1635 3758 1703 3762
rect 1707 3758 1767 3762
rect 1771 3758 1831 3762
rect 1835 3758 1935 3762
rect 1939 3758 2031 3762
rect 2035 3758 2043 3762
rect 91 3757 2043 3758
rect 2049 3757 2050 3763
rect 2054 3689 2055 3695
rect 2061 3694 4027 3695
rect 2061 3690 2071 3694
rect 2075 3690 2111 3694
rect 2115 3690 2255 3694
rect 2259 3690 2335 3694
rect 2339 3690 2439 3694
rect 2443 3690 2559 3694
rect 2563 3690 2623 3694
rect 2627 3690 2775 3694
rect 2779 3690 2815 3694
rect 2819 3690 2975 3694
rect 2979 3690 3007 3694
rect 3011 3690 3159 3694
rect 3163 3690 3199 3694
rect 3203 3690 3327 3694
rect 3331 3690 3391 3694
rect 3395 3690 3479 3694
rect 3483 3690 3583 3694
rect 3587 3690 3623 3694
rect 3627 3690 3767 3694
rect 3771 3690 3895 3694
rect 3899 3690 3991 3694
rect 3995 3690 4027 3694
rect 2061 3689 4027 3690
rect 4033 3689 4034 3695
rect 2054 3687 2062 3689
rect 96 3681 97 3687
rect 103 3686 2055 3687
rect 103 3682 111 3686
rect 115 3682 471 3686
rect 475 3682 599 3686
rect 603 3682 615 3686
rect 619 3682 719 3686
rect 723 3682 759 3686
rect 763 3682 847 3686
rect 851 3682 903 3686
rect 907 3682 983 3686
rect 987 3682 1047 3686
rect 1051 3682 1111 3686
rect 1115 3682 1191 3686
rect 1195 3682 1239 3686
rect 1243 3682 1335 3686
rect 1339 3682 1367 3686
rect 1371 3682 1479 3686
rect 1483 3682 1495 3686
rect 1499 3682 1631 3686
rect 1635 3682 1767 3686
rect 1771 3682 2031 3686
rect 2035 3682 2055 3686
rect 103 3681 2055 3682
rect 2061 3681 2062 3687
rect 598 3668 604 3669
rect 910 3668 916 3669
rect 598 3664 599 3668
rect 603 3664 911 3668
rect 915 3664 916 3668
rect 598 3663 604 3664
rect 910 3663 916 3664
rect 84 3609 85 3615
rect 91 3614 2043 3615
rect 91 3610 111 3614
rect 115 3610 247 3614
rect 251 3610 375 3614
rect 379 3610 471 3614
rect 475 3610 519 3614
rect 523 3610 615 3614
rect 619 3610 679 3614
rect 683 3610 759 3614
rect 763 3610 847 3614
rect 851 3610 903 3614
rect 907 3610 1023 3614
rect 1027 3610 1047 3614
rect 1051 3610 1191 3614
rect 1195 3610 1207 3614
rect 1211 3610 1335 3614
rect 1339 3610 1391 3614
rect 1395 3610 1479 3614
rect 1483 3610 1575 3614
rect 1579 3610 1767 3614
rect 1771 3610 1935 3614
rect 1939 3610 2031 3614
rect 2035 3610 2043 3614
rect 91 3609 2043 3610
rect 2049 3611 2050 3615
rect 2049 3610 4022 3611
rect 2049 3609 2071 3610
rect 2042 3606 2071 3609
rect 2075 3606 2111 3610
rect 2115 3606 2255 3610
rect 2259 3606 2359 3610
rect 2363 3606 2439 3610
rect 2443 3606 2583 3610
rect 2587 3606 2623 3610
rect 2627 3606 2799 3610
rect 2803 3606 2815 3610
rect 2819 3606 3007 3610
rect 3011 3606 3199 3610
rect 3203 3606 3215 3610
rect 3219 3606 3391 3610
rect 3395 3606 3431 3610
rect 3435 3606 3583 3610
rect 3587 3606 3991 3610
rect 3995 3606 4022 3610
rect 2042 3605 4022 3606
rect 1174 3556 1180 3557
rect 1462 3556 1468 3557
rect 1174 3552 1175 3556
rect 1179 3552 1463 3556
rect 1467 3552 1468 3556
rect 1174 3551 1180 3552
rect 1462 3551 1468 3552
rect 2054 3534 4034 3535
rect 2054 3531 2071 3534
rect 96 3525 97 3531
rect 103 3530 2055 3531
rect 103 3526 111 3530
rect 115 3526 151 3530
rect 155 3526 247 3530
rect 251 3526 263 3530
rect 267 3526 375 3530
rect 379 3526 399 3530
rect 403 3526 519 3530
rect 523 3526 543 3530
rect 547 3526 679 3530
rect 683 3526 687 3530
rect 691 3526 831 3530
rect 835 3526 847 3530
rect 851 3526 967 3530
rect 971 3526 1023 3530
rect 1027 3526 1095 3530
rect 1099 3526 1207 3530
rect 1211 3526 1223 3530
rect 1227 3526 1343 3530
rect 1347 3526 1391 3530
rect 1395 3526 1463 3530
rect 1467 3526 1575 3530
rect 1579 3526 1583 3530
rect 1587 3526 1711 3530
rect 1715 3526 1767 3530
rect 1771 3526 1935 3530
rect 1939 3526 2031 3530
rect 2035 3526 2055 3530
rect 103 3525 2055 3526
rect 2061 3530 2071 3531
rect 2075 3530 2359 3534
rect 2363 3530 2439 3534
rect 2443 3530 2575 3534
rect 2579 3530 2583 3534
rect 2587 3530 2703 3534
rect 2707 3530 2799 3534
rect 2803 3530 2831 3534
rect 2835 3530 2951 3534
rect 2955 3530 3007 3534
rect 3011 3530 3071 3534
rect 3075 3530 3199 3534
rect 3203 3530 3215 3534
rect 3219 3530 3327 3534
rect 3331 3530 3431 3534
rect 3435 3530 3991 3534
rect 3995 3530 4034 3534
rect 2061 3529 4034 3530
rect 2061 3525 2062 3529
rect 2042 3462 4022 3463
rect 2042 3459 2071 3462
rect 84 3453 85 3459
rect 91 3458 2043 3459
rect 91 3454 111 3458
rect 115 3454 151 3458
rect 155 3454 263 3458
rect 267 3454 399 3458
rect 403 3454 423 3458
rect 427 3454 543 3458
rect 547 3454 687 3458
rect 691 3454 743 3458
rect 747 3454 831 3458
rect 835 3454 967 3458
rect 971 3454 1071 3458
rect 1075 3454 1095 3458
rect 1099 3454 1223 3458
rect 1227 3454 1343 3458
rect 1347 3454 1399 3458
rect 1403 3454 1463 3458
rect 1467 3454 1583 3458
rect 1587 3454 1711 3458
rect 1715 3454 2031 3458
rect 2035 3454 2043 3458
rect 91 3453 2043 3454
rect 2049 3458 2071 3459
rect 2075 3458 2359 3462
rect 2363 3458 2439 3462
rect 2443 3458 2463 3462
rect 2467 3458 2567 3462
rect 2571 3458 2575 3462
rect 2579 3458 2671 3462
rect 2675 3458 2703 3462
rect 2707 3458 2775 3462
rect 2779 3458 2831 3462
rect 2835 3458 2879 3462
rect 2883 3458 2951 3462
rect 2955 3458 2983 3462
rect 2987 3458 3071 3462
rect 3075 3458 3087 3462
rect 3091 3458 3191 3462
rect 3195 3458 3199 3462
rect 3203 3458 3327 3462
rect 3331 3458 3991 3462
rect 3995 3458 4022 3462
rect 2049 3457 4022 3458
rect 2049 3453 2050 3457
rect 96 3357 97 3363
rect 103 3362 2055 3363
rect 103 3358 111 3362
rect 115 3358 151 3362
rect 155 3358 319 3362
rect 323 3358 423 3362
rect 427 3358 527 3362
rect 531 3358 743 3362
rect 747 3358 959 3362
rect 963 3358 1071 3362
rect 1075 3358 1167 3362
rect 1171 3358 1367 3362
rect 1371 3358 1399 3362
rect 1403 3358 1559 3362
rect 1563 3358 1751 3362
rect 1755 3358 1935 3362
rect 1939 3358 2031 3362
rect 2035 3358 2055 3362
rect 103 3357 2055 3358
rect 2061 3362 4034 3363
rect 2061 3358 2071 3362
rect 2075 3358 2359 3362
rect 2363 3358 2439 3362
rect 2443 3358 2463 3362
rect 2467 3358 2543 3362
rect 2547 3358 2567 3362
rect 2571 3358 2647 3362
rect 2651 3358 2671 3362
rect 2675 3358 2751 3362
rect 2755 3358 2775 3362
rect 2779 3358 2855 3362
rect 2859 3358 2879 3362
rect 2883 3358 2959 3362
rect 2963 3358 2983 3362
rect 2987 3358 3087 3362
rect 3091 3358 3191 3362
rect 3195 3358 3991 3362
rect 3995 3358 4034 3362
rect 2061 3357 4034 3358
rect 2042 3285 2043 3291
rect 2049 3290 4015 3291
rect 2049 3286 2071 3290
rect 2075 3286 2439 3290
rect 2443 3286 2527 3290
rect 2531 3286 2543 3290
rect 2547 3286 2631 3290
rect 2635 3286 2647 3290
rect 2651 3286 2735 3290
rect 2739 3286 2751 3290
rect 2755 3286 2839 3290
rect 2843 3286 2855 3290
rect 2859 3286 2943 3290
rect 2947 3286 2959 3290
rect 2963 3286 3047 3290
rect 3051 3286 3151 3290
rect 3155 3286 3255 3290
rect 3259 3286 3991 3290
rect 3995 3286 4015 3290
rect 2049 3285 4015 3286
rect 4021 3285 4022 3291
rect 2042 3283 2050 3285
rect 84 3277 85 3283
rect 91 3282 2043 3283
rect 91 3278 111 3282
rect 115 3278 151 3282
rect 155 3278 311 3282
rect 315 3278 319 3282
rect 323 3278 479 3282
rect 483 3278 527 3282
rect 531 3278 655 3282
rect 659 3278 743 3282
rect 747 3278 847 3282
rect 851 3278 959 3282
rect 963 3278 1039 3282
rect 1043 3278 1167 3282
rect 1171 3278 1231 3282
rect 1235 3278 1367 3282
rect 1371 3278 1431 3282
rect 1435 3278 1559 3282
rect 1563 3278 1631 3282
rect 1635 3278 1751 3282
rect 1755 3278 1831 3282
rect 1835 3278 1935 3282
rect 1939 3278 2031 3282
rect 2035 3278 2043 3282
rect 91 3277 2043 3278
rect 2049 3277 2050 3283
rect 2718 3228 2724 3229
rect 3014 3228 3020 3229
rect 2718 3224 2719 3228
rect 2723 3224 3015 3228
rect 3019 3224 3020 3228
rect 2718 3223 2724 3224
rect 3014 3223 3020 3224
rect 2054 3213 2055 3219
rect 2061 3218 4027 3219
rect 2061 3214 2071 3218
rect 2075 3214 2399 3218
rect 2403 3214 2527 3218
rect 2531 3214 2551 3218
rect 2555 3214 2631 3218
rect 2635 3214 2695 3218
rect 2699 3214 2735 3218
rect 2739 3214 2839 3218
rect 2843 3214 2943 3218
rect 2947 3214 2975 3218
rect 2979 3214 3047 3218
rect 3051 3214 3111 3218
rect 3115 3214 3151 3218
rect 3155 3214 3247 3218
rect 3251 3214 3255 3218
rect 3259 3214 3391 3218
rect 3395 3214 3991 3218
rect 3995 3214 4027 3218
rect 2061 3213 4027 3214
rect 4033 3213 4034 3219
rect 96 3201 97 3207
rect 103 3206 2055 3207
rect 103 3202 111 3206
rect 115 3202 311 3206
rect 315 3202 479 3206
rect 483 3202 623 3206
rect 627 3202 655 3206
rect 659 3202 759 3206
rect 763 3202 847 3206
rect 851 3202 903 3206
rect 907 3202 1039 3206
rect 1043 3202 1055 3206
rect 1059 3202 1207 3206
rect 1211 3202 1231 3206
rect 1235 3202 1351 3206
rect 1355 3202 1431 3206
rect 1435 3202 1503 3206
rect 1507 3202 1631 3206
rect 1635 3202 1655 3206
rect 1659 3202 1807 3206
rect 1811 3202 1831 3206
rect 1835 3202 1935 3206
rect 1939 3202 2031 3206
rect 2035 3202 2055 3206
rect 103 3201 2055 3202
rect 2061 3201 2062 3207
rect 742 3196 748 3197
rect 1046 3196 1052 3197
rect 742 3192 743 3196
rect 747 3192 1047 3196
rect 1051 3192 1052 3196
rect 742 3191 748 3192
rect 1046 3191 1052 3192
rect 2958 3196 2964 3197
rect 3398 3196 3404 3197
rect 2958 3192 2959 3196
rect 2963 3192 3399 3196
rect 3403 3192 3404 3196
rect 2958 3191 2964 3192
rect 3398 3191 3404 3192
rect 84 3129 85 3135
rect 91 3134 2043 3135
rect 91 3130 111 3134
rect 115 3130 599 3134
rect 603 3130 623 3134
rect 627 3130 703 3134
rect 707 3130 759 3134
rect 763 3130 807 3134
rect 811 3130 903 3134
rect 907 3130 911 3134
rect 915 3130 1039 3134
rect 1043 3130 1055 3134
rect 1059 3130 1183 3134
rect 1187 3130 1207 3134
rect 1211 3130 1351 3134
rect 1355 3130 1359 3134
rect 1363 3130 1503 3134
rect 1507 3130 1551 3134
rect 1555 3130 1655 3134
rect 1659 3130 1751 3134
rect 1755 3130 1807 3134
rect 1811 3130 1935 3134
rect 1939 3130 2031 3134
rect 2035 3130 2043 3134
rect 91 3129 2043 3130
rect 2049 3134 4022 3135
rect 2049 3130 2071 3134
rect 2075 3130 2111 3134
rect 2115 3130 2343 3134
rect 2347 3130 2399 3134
rect 2403 3130 2551 3134
rect 2555 3130 2583 3134
rect 2587 3130 2695 3134
rect 2699 3130 2799 3134
rect 2803 3130 2839 3134
rect 2843 3130 2975 3134
rect 2979 3130 2999 3134
rect 3003 3130 3111 3134
rect 3115 3130 3191 3134
rect 3195 3130 3247 3134
rect 3251 3130 3375 3134
rect 3379 3130 3391 3134
rect 3395 3130 3567 3134
rect 3571 3130 3991 3134
rect 3995 3130 4022 3134
rect 2049 3129 4022 3130
rect 2054 3058 4034 3059
rect 2054 3055 2071 3058
rect 96 3049 97 3055
rect 103 3054 2055 3055
rect 103 3050 111 3054
rect 115 3050 311 3054
rect 315 3050 415 3054
rect 419 3050 527 3054
rect 531 3050 599 3054
rect 603 3050 639 3054
rect 643 3050 703 3054
rect 707 3050 751 3054
rect 755 3050 807 3054
rect 811 3050 863 3054
rect 867 3050 911 3054
rect 915 3050 975 3054
rect 979 3050 1039 3054
rect 1043 3050 1095 3054
rect 1099 3050 1183 3054
rect 1187 3050 1215 3054
rect 1219 3050 1335 3054
rect 1339 3050 1359 3054
rect 1363 3050 1551 3054
rect 1555 3050 1751 3054
rect 1755 3050 1935 3054
rect 1939 3050 2031 3054
rect 2035 3050 2055 3054
rect 103 3049 2055 3050
rect 2061 3054 2071 3055
rect 2075 3054 2111 3058
rect 2115 3054 2263 3058
rect 2267 3054 2343 3058
rect 2347 3054 2455 3058
rect 2459 3054 2583 3058
rect 2587 3054 2655 3058
rect 2659 3054 2799 3058
rect 2803 3054 2855 3058
rect 2859 3054 2999 3058
rect 3003 3054 3055 3058
rect 3059 3054 3191 3058
rect 3195 3054 3255 3058
rect 3259 3054 3375 3058
rect 3379 3054 3455 3058
rect 3459 3054 3567 3058
rect 3571 3054 3655 3058
rect 3659 3054 3991 3058
rect 3995 3054 4034 3058
rect 2061 3053 4034 3054
rect 2061 3049 2062 3053
rect 2042 2981 2043 2987
rect 2049 2986 4015 2987
rect 2049 2982 2071 2986
rect 2075 2982 2111 2986
rect 2115 2982 2263 2986
rect 2267 2982 2359 2986
rect 2363 2982 2455 2986
rect 2459 2982 2607 2986
rect 2611 2982 2655 2986
rect 2659 2982 2847 2986
rect 2851 2982 2855 2986
rect 2859 2982 3055 2986
rect 3059 2982 3079 2986
rect 3083 2982 3255 2986
rect 3259 2982 3303 2986
rect 3307 2982 3455 2986
rect 3459 2982 3535 2986
rect 3539 2982 3655 2986
rect 3659 2982 3767 2986
rect 3771 2982 3991 2986
rect 3995 2982 4015 2986
rect 2049 2981 4015 2982
rect 4021 2981 4022 2987
rect 84 2969 85 2975
rect 91 2974 2043 2975
rect 91 2970 111 2974
rect 115 2970 151 2974
rect 155 2970 271 2974
rect 275 2970 311 2974
rect 315 2970 415 2974
rect 419 2970 431 2974
rect 435 2970 527 2974
rect 531 2970 607 2974
rect 611 2970 639 2974
rect 643 2970 751 2974
rect 755 2970 783 2974
rect 787 2970 863 2974
rect 867 2970 959 2974
rect 963 2970 975 2974
rect 979 2970 1095 2974
rect 1099 2970 1135 2974
rect 1139 2970 1215 2974
rect 1219 2970 1303 2974
rect 1307 2970 1335 2974
rect 1339 2970 1471 2974
rect 1475 2970 1647 2974
rect 1651 2970 2031 2974
rect 2035 2970 2043 2974
rect 91 2969 2043 2970
rect 2049 2969 2050 2975
rect 2054 2901 2055 2907
rect 2061 2906 4027 2907
rect 2061 2902 2071 2906
rect 2075 2902 2111 2906
rect 2115 2902 2279 2906
rect 2283 2902 2359 2906
rect 2363 2902 2487 2906
rect 2491 2902 2607 2906
rect 2611 2902 2695 2906
rect 2699 2902 2847 2906
rect 2851 2902 2903 2906
rect 2907 2902 3079 2906
rect 3083 2902 3111 2906
rect 3115 2902 3303 2906
rect 3307 2902 3495 2906
rect 3499 2902 3535 2906
rect 3539 2902 3687 2906
rect 3691 2902 3767 2906
rect 3771 2902 3879 2906
rect 3883 2902 3991 2906
rect 3995 2902 4027 2906
rect 2061 2901 4027 2902
rect 4033 2901 4034 2907
rect 96 2885 97 2891
rect 103 2890 2055 2891
rect 103 2886 111 2890
rect 115 2886 151 2890
rect 155 2886 271 2890
rect 275 2886 287 2890
rect 291 2886 431 2890
rect 435 2886 447 2890
rect 451 2886 599 2890
rect 603 2886 607 2890
rect 611 2886 759 2890
rect 763 2886 783 2890
rect 787 2886 927 2890
rect 931 2886 959 2890
rect 963 2886 1103 2890
rect 1107 2886 1135 2890
rect 1139 2886 1287 2890
rect 1291 2886 1303 2890
rect 1307 2886 1471 2890
rect 1475 2886 1479 2890
rect 1483 2886 1647 2890
rect 1651 2886 1671 2890
rect 1675 2886 2031 2890
rect 2035 2886 2055 2890
rect 103 2885 2055 2886
rect 2061 2885 2062 2891
rect 2042 2817 2043 2823
rect 2049 2822 4015 2823
rect 2049 2818 2071 2822
rect 2075 2818 2111 2822
rect 2115 2818 2143 2822
rect 2147 2818 2279 2822
rect 2283 2818 2319 2822
rect 2323 2818 2487 2822
rect 2491 2818 2503 2822
rect 2507 2818 2695 2822
rect 2699 2818 2887 2822
rect 2891 2818 2903 2822
rect 2907 2818 3079 2822
rect 3083 2818 3111 2822
rect 3115 2818 3263 2822
rect 3267 2818 3303 2822
rect 3307 2818 3439 2822
rect 3443 2818 3495 2822
rect 3499 2818 3615 2822
rect 3619 2818 3687 2822
rect 3691 2818 3791 2822
rect 3795 2818 3879 2822
rect 3883 2818 3991 2822
rect 3995 2818 4015 2822
rect 2049 2817 4015 2818
rect 4021 2817 4022 2823
rect 84 2801 85 2807
rect 91 2806 2043 2807
rect 91 2802 111 2806
rect 115 2802 151 2806
rect 155 2802 287 2806
rect 291 2802 319 2806
rect 323 2802 447 2806
rect 451 2802 503 2806
rect 507 2802 599 2806
rect 603 2802 687 2806
rect 691 2802 759 2806
rect 763 2802 871 2806
rect 875 2802 927 2806
rect 931 2802 1055 2806
rect 1059 2802 1103 2806
rect 1107 2802 1239 2806
rect 1243 2802 1287 2806
rect 1291 2802 1431 2806
rect 1435 2802 1479 2806
rect 1483 2802 1631 2806
rect 1635 2802 1671 2806
rect 1675 2802 1831 2806
rect 1835 2802 2031 2806
rect 2035 2802 2043 2806
rect 91 2801 2043 2802
rect 2049 2801 2050 2807
rect 2054 2733 2055 2739
rect 2061 2738 4027 2739
rect 2061 2734 2071 2738
rect 2075 2734 2111 2738
rect 2115 2734 2143 2738
rect 2147 2734 2279 2738
rect 2283 2734 2319 2738
rect 2323 2734 2455 2738
rect 2459 2734 2503 2738
rect 2507 2734 2639 2738
rect 2643 2734 2695 2738
rect 2699 2734 2815 2738
rect 2819 2734 2887 2738
rect 2891 2734 2983 2738
rect 2987 2734 3079 2738
rect 3083 2734 3143 2738
rect 3147 2734 3263 2738
rect 3267 2734 3303 2738
rect 3307 2734 3439 2738
rect 3443 2734 3463 2738
rect 3467 2734 3615 2738
rect 3619 2734 3623 2738
rect 3627 2734 3791 2738
rect 3795 2734 3991 2738
rect 3995 2734 4027 2738
rect 2061 2733 4027 2734
rect 4033 2733 4034 2739
rect 2054 2731 2062 2733
rect 96 2725 97 2731
rect 103 2730 2055 2731
rect 103 2726 111 2730
rect 115 2726 151 2730
rect 155 2726 183 2730
rect 187 2726 319 2730
rect 323 2726 383 2730
rect 387 2726 503 2730
rect 507 2726 583 2730
rect 587 2726 687 2730
rect 691 2726 783 2730
rect 787 2726 871 2730
rect 875 2726 983 2730
rect 987 2726 1055 2730
rect 1059 2726 1199 2730
rect 1203 2726 1239 2730
rect 1243 2726 1415 2730
rect 1419 2726 1431 2730
rect 1435 2726 1631 2730
rect 1635 2726 1639 2730
rect 1643 2726 1831 2730
rect 1835 2726 1871 2730
rect 1875 2726 2031 2730
rect 2035 2726 2055 2730
rect 103 2725 2055 2726
rect 2061 2725 2062 2731
rect 2042 2654 4022 2655
rect 2042 2651 2071 2654
rect 84 2645 85 2651
rect 91 2650 2043 2651
rect 91 2646 111 2650
rect 115 2646 183 2650
rect 187 2646 255 2650
rect 259 2646 383 2650
rect 387 2646 423 2650
rect 427 2646 583 2650
rect 587 2646 599 2650
rect 603 2646 775 2650
rect 779 2646 783 2650
rect 787 2646 959 2650
rect 963 2646 983 2650
rect 987 2646 1151 2650
rect 1155 2646 1199 2650
rect 1203 2646 1343 2650
rect 1347 2646 1415 2650
rect 1419 2646 1535 2650
rect 1539 2646 1639 2650
rect 1643 2646 1727 2650
rect 1731 2646 1871 2650
rect 1875 2646 1927 2650
rect 1931 2646 2031 2650
rect 2035 2646 2043 2650
rect 91 2645 2043 2646
rect 2049 2650 2071 2651
rect 2075 2650 2111 2654
rect 2115 2650 2263 2654
rect 2267 2650 2279 2654
rect 2283 2650 2431 2654
rect 2435 2650 2455 2654
rect 2459 2650 2599 2654
rect 2603 2650 2639 2654
rect 2643 2650 2751 2654
rect 2755 2650 2815 2654
rect 2819 2650 2895 2654
rect 2899 2650 2983 2654
rect 2987 2650 3039 2654
rect 3043 2650 3143 2654
rect 3147 2650 3175 2654
rect 3179 2650 3303 2654
rect 3307 2650 3311 2654
rect 3315 2650 3455 2654
rect 3459 2650 3463 2654
rect 3467 2650 3623 2654
rect 3627 2650 3991 2654
rect 3995 2650 4022 2654
rect 2049 2649 4022 2650
rect 2049 2645 2050 2649
rect 3126 2596 3132 2597
rect 3526 2596 3532 2597
rect 3126 2592 3127 2596
rect 3131 2592 3527 2596
rect 3531 2592 3532 2596
rect 3126 2591 3132 2592
rect 3526 2591 3532 2592
rect 96 2569 97 2575
rect 103 2574 2055 2575
rect 103 2570 111 2574
rect 115 2570 255 2574
rect 259 2570 319 2574
rect 323 2570 423 2574
rect 427 2570 535 2574
rect 539 2570 599 2574
rect 603 2570 743 2574
rect 747 2570 775 2574
rect 779 2570 951 2574
rect 955 2570 959 2574
rect 963 2570 1151 2574
rect 1155 2570 1159 2574
rect 1163 2570 1343 2574
rect 1347 2570 1359 2574
rect 1363 2570 1535 2574
rect 1539 2570 1559 2574
rect 1563 2570 1727 2574
rect 1731 2570 1759 2574
rect 1763 2570 1927 2574
rect 1931 2570 1935 2574
rect 1939 2570 2031 2574
rect 2035 2570 2055 2574
rect 103 2569 2055 2570
rect 2061 2574 4034 2575
rect 2061 2570 2071 2574
rect 2075 2570 2111 2574
rect 2115 2570 2263 2574
rect 2267 2570 2271 2574
rect 2275 2570 2431 2574
rect 2435 2570 2447 2574
rect 2451 2570 2599 2574
rect 2603 2570 2615 2574
rect 2619 2570 2751 2574
rect 2755 2570 2767 2574
rect 2771 2570 2895 2574
rect 2899 2570 2911 2574
rect 2915 2570 3039 2574
rect 3043 2570 3047 2574
rect 3051 2570 3175 2574
rect 3179 2570 3183 2574
rect 3187 2570 3311 2574
rect 3315 2570 3319 2574
rect 3323 2570 3455 2574
rect 3459 2570 3991 2574
rect 3995 2570 4034 2574
rect 2061 2569 4034 2570
rect 84 2497 85 2503
rect 91 2502 2043 2503
rect 91 2498 111 2502
rect 115 2498 279 2502
rect 283 2498 319 2502
rect 323 2498 439 2502
rect 443 2498 535 2502
rect 539 2498 607 2502
rect 611 2498 743 2502
rect 747 2498 783 2502
rect 787 2498 951 2502
rect 955 2498 959 2502
rect 963 2498 1127 2502
rect 1131 2498 1159 2502
rect 1163 2498 1295 2502
rect 1299 2498 1359 2502
rect 1363 2498 1463 2502
rect 1467 2498 1559 2502
rect 1563 2498 1623 2502
rect 1627 2498 1759 2502
rect 1763 2498 1791 2502
rect 1795 2498 1935 2502
rect 1939 2498 2031 2502
rect 2035 2498 2043 2502
rect 91 2497 2043 2498
rect 2049 2497 2050 2503
rect 2042 2485 2043 2491
rect 2049 2490 4015 2491
rect 2049 2486 2071 2490
rect 2075 2486 2111 2490
rect 2115 2486 2271 2490
rect 2275 2486 2447 2490
rect 2451 2486 2615 2490
rect 2619 2486 2623 2490
rect 2627 2486 2743 2490
rect 2747 2486 2767 2490
rect 2771 2486 2871 2490
rect 2875 2486 2911 2490
rect 2915 2486 3015 2490
rect 3019 2486 3047 2490
rect 3051 2486 3159 2490
rect 3163 2486 3183 2490
rect 3187 2486 3311 2490
rect 3315 2486 3319 2490
rect 3323 2486 3463 2490
rect 3467 2486 3615 2490
rect 3619 2486 3767 2490
rect 3771 2486 3895 2490
rect 3899 2486 3991 2490
rect 3995 2486 4015 2490
rect 2049 2485 4015 2486
rect 4021 2485 4022 2491
rect 96 2417 97 2423
rect 103 2422 2055 2423
rect 103 2418 111 2422
rect 115 2418 279 2422
rect 283 2418 327 2422
rect 331 2418 439 2422
rect 443 2418 471 2422
rect 475 2418 607 2422
rect 611 2418 623 2422
rect 627 2418 783 2422
rect 787 2418 943 2422
rect 947 2418 959 2422
rect 963 2418 1095 2422
rect 1099 2418 1127 2422
rect 1131 2418 1247 2422
rect 1251 2418 1295 2422
rect 1299 2418 1391 2422
rect 1395 2418 1463 2422
rect 1467 2418 1535 2422
rect 1539 2418 1623 2422
rect 1627 2418 1671 2422
rect 1675 2418 1791 2422
rect 1795 2418 1815 2422
rect 1819 2418 1935 2422
rect 1939 2418 2031 2422
rect 2035 2418 2055 2422
rect 103 2417 2055 2418
rect 2061 2417 2062 2423
rect 2054 2401 2055 2407
rect 2061 2406 4027 2407
rect 2061 2402 2071 2406
rect 2075 2402 2487 2406
rect 2491 2402 2599 2406
rect 2603 2402 2623 2406
rect 2627 2402 2727 2406
rect 2731 2402 2743 2406
rect 2747 2402 2871 2406
rect 2875 2402 2879 2406
rect 2883 2402 3015 2406
rect 3019 2402 3055 2406
rect 3059 2402 3159 2406
rect 3163 2402 3247 2406
rect 3251 2402 3311 2406
rect 3315 2402 3455 2406
rect 3459 2402 3463 2406
rect 3467 2402 3615 2406
rect 3619 2402 3679 2406
rect 3683 2402 3767 2406
rect 3771 2402 3895 2406
rect 3899 2402 3991 2406
rect 3995 2402 4027 2406
rect 2061 2401 4027 2402
rect 4033 2401 4034 2407
rect 84 2337 85 2343
rect 91 2342 2043 2343
rect 91 2338 111 2342
rect 115 2338 327 2342
rect 331 2338 359 2342
rect 363 2338 471 2342
rect 475 2338 495 2342
rect 499 2338 623 2342
rect 627 2338 639 2342
rect 643 2338 783 2342
rect 787 2338 935 2342
rect 939 2338 943 2342
rect 947 2338 1087 2342
rect 1091 2338 1095 2342
rect 1099 2338 1247 2342
rect 1251 2338 1391 2342
rect 1395 2338 1415 2342
rect 1419 2338 1535 2342
rect 1539 2338 1591 2342
rect 1595 2338 1671 2342
rect 1675 2338 1775 2342
rect 1779 2338 1815 2342
rect 1819 2338 1935 2342
rect 1939 2338 2031 2342
rect 2035 2338 2043 2342
rect 91 2337 2043 2338
rect 2049 2337 2050 2343
rect 2042 2317 2043 2323
rect 2049 2322 4015 2323
rect 2049 2318 2071 2322
rect 2075 2318 2111 2322
rect 2115 2318 2223 2322
rect 2227 2318 2359 2322
rect 2363 2318 2487 2322
rect 2491 2318 2511 2322
rect 2515 2318 2599 2322
rect 2603 2318 2671 2322
rect 2675 2318 2727 2322
rect 2731 2318 2847 2322
rect 2851 2318 2879 2322
rect 2883 2318 3039 2322
rect 3043 2318 3055 2322
rect 3059 2318 3247 2322
rect 3251 2318 3455 2322
rect 3459 2318 3463 2322
rect 3467 2318 3679 2322
rect 3683 2318 3687 2322
rect 3691 2318 3895 2322
rect 3899 2318 3991 2322
rect 3995 2318 4015 2322
rect 2049 2317 4015 2318
rect 4021 2317 4022 2323
rect 96 2253 97 2259
rect 103 2258 2055 2259
rect 103 2254 111 2258
rect 115 2254 239 2258
rect 243 2254 359 2258
rect 363 2254 391 2258
rect 395 2254 495 2258
rect 499 2254 551 2258
rect 555 2254 639 2258
rect 643 2254 711 2258
rect 715 2254 783 2258
rect 787 2254 871 2258
rect 875 2254 935 2258
rect 939 2254 1031 2258
rect 1035 2254 1087 2258
rect 1091 2254 1191 2258
rect 1195 2254 1247 2258
rect 1251 2254 1359 2258
rect 1363 2254 1415 2258
rect 1419 2254 1527 2258
rect 1531 2254 1591 2258
rect 1595 2254 1695 2258
rect 1699 2254 1775 2258
rect 1779 2254 1935 2258
rect 1939 2254 2031 2258
rect 2035 2254 2055 2258
rect 103 2253 2055 2254
rect 2061 2253 2062 2259
rect 2054 2237 2055 2243
rect 2061 2242 4027 2243
rect 2061 2238 2071 2242
rect 2075 2238 2111 2242
rect 2115 2238 2223 2242
rect 2227 2238 2279 2242
rect 2283 2238 2359 2242
rect 2363 2238 2479 2242
rect 2483 2238 2511 2242
rect 2515 2238 2671 2242
rect 2675 2238 2679 2242
rect 2683 2238 2847 2242
rect 2851 2238 2879 2242
rect 2883 2238 3039 2242
rect 3043 2238 3079 2242
rect 3083 2238 3247 2242
rect 3251 2238 3279 2242
rect 3283 2238 3463 2242
rect 3467 2238 3487 2242
rect 3491 2238 3687 2242
rect 3691 2238 3703 2242
rect 3707 2238 3895 2242
rect 3899 2238 3991 2242
rect 3995 2238 4027 2242
rect 2061 2237 4027 2238
rect 4033 2237 4034 2243
rect 3062 2228 3068 2229
rect 3258 2228 3264 2229
rect 3062 2224 3063 2228
rect 3067 2224 3259 2228
rect 3263 2224 3264 2228
rect 3062 2223 3068 2224
rect 3258 2223 3264 2224
rect 84 2169 85 2175
rect 91 2174 2043 2175
rect 91 2170 111 2174
rect 115 2170 151 2174
rect 155 2170 239 2174
rect 243 2170 319 2174
rect 323 2170 391 2174
rect 395 2170 511 2174
rect 515 2170 551 2174
rect 555 2170 703 2174
rect 707 2170 711 2174
rect 715 2170 871 2174
rect 875 2170 895 2174
rect 899 2170 1031 2174
rect 1035 2170 1087 2174
rect 1091 2170 1191 2174
rect 1195 2170 1279 2174
rect 1283 2170 1359 2174
rect 1363 2170 1463 2174
rect 1467 2170 1527 2174
rect 1531 2170 1655 2174
rect 1659 2170 1695 2174
rect 1699 2170 1847 2174
rect 1851 2170 2031 2174
rect 2035 2170 2043 2174
rect 91 2169 2043 2170
rect 2049 2169 2050 2175
rect 2042 2157 2043 2163
rect 2049 2162 4015 2163
rect 2049 2158 2071 2162
rect 2075 2158 2111 2162
rect 2115 2158 2143 2162
rect 2147 2158 2279 2162
rect 2283 2158 2319 2162
rect 2323 2158 2479 2162
rect 2483 2158 2495 2162
rect 2499 2158 2679 2162
rect 2683 2158 2863 2162
rect 2867 2158 2879 2162
rect 2883 2158 3039 2162
rect 3043 2158 3079 2162
rect 3083 2158 3215 2162
rect 3219 2158 3279 2162
rect 3283 2158 3391 2162
rect 3395 2158 3487 2162
rect 3491 2158 3567 2162
rect 3571 2158 3703 2162
rect 3707 2158 3743 2162
rect 3747 2158 3895 2162
rect 3899 2158 3991 2162
rect 3995 2158 4015 2162
rect 2049 2157 4015 2158
rect 4021 2157 4022 2163
rect 96 2089 97 2095
rect 103 2094 2055 2095
rect 103 2090 111 2094
rect 115 2090 151 2094
rect 155 2090 303 2094
rect 307 2090 319 2094
rect 323 2090 479 2094
rect 483 2090 511 2094
rect 515 2090 663 2094
rect 667 2090 703 2094
rect 707 2090 847 2094
rect 851 2090 895 2094
rect 899 2090 1039 2094
rect 1043 2090 1087 2094
rect 1091 2090 1239 2094
rect 1243 2090 1279 2094
rect 1283 2090 1447 2094
rect 1451 2090 1463 2094
rect 1467 2090 1655 2094
rect 1659 2090 1663 2094
rect 1667 2090 1847 2094
rect 1851 2090 1879 2094
rect 1883 2090 2031 2094
rect 2035 2090 2055 2094
rect 103 2089 2055 2090
rect 2061 2089 2062 2095
rect 2054 2073 2055 2079
rect 2061 2078 4027 2079
rect 2061 2074 2071 2078
rect 2075 2074 2143 2078
rect 2147 2074 2207 2078
rect 2211 2074 2319 2078
rect 2323 2074 2391 2078
rect 2395 2074 2495 2078
rect 2499 2074 2575 2078
rect 2579 2074 2679 2078
rect 2683 2074 2759 2078
rect 2763 2074 2863 2078
rect 2867 2074 2935 2078
rect 2939 2074 3039 2078
rect 3043 2074 3103 2078
rect 3107 2074 3215 2078
rect 3219 2074 3263 2078
rect 3267 2074 3391 2078
rect 3395 2074 3423 2078
rect 3427 2074 3567 2078
rect 3571 2074 3583 2078
rect 3587 2074 3743 2078
rect 3747 2074 3751 2078
rect 3755 2074 3895 2078
rect 3899 2074 3991 2078
rect 3995 2074 4027 2078
rect 2061 2073 4027 2074
rect 4033 2073 4034 2079
rect 84 2009 85 2015
rect 91 2014 2043 2015
rect 91 2010 111 2014
rect 115 2010 151 2014
rect 155 2010 303 2014
rect 307 2010 479 2014
rect 483 2010 487 2014
rect 491 2010 663 2014
rect 667 2010 687 2014
rect 691 2010 847 2014
rect 851 2010 895 2014
rect 899 2010 1039 2014
rect 1043 2010 1103 2014
rect 1107 2010 1239 2014
rect 1243 2010 1311 2014
rect 1315 2010 1447 2014
rect 1451 2010 1527 2014
rect 1531 2010 1663 2014
rect 1667 2010 1743 2014
rect 1747 2010 1879 2014
rect 1883 2010 1935 2014
rect 1939 2010 2031 2014
rect 2035 2010 2043 2014
rect 91 2009 2043 2010
rect 2049 2009 2050 2015
rect 2042 1989 2043 1995
rect 2049 1994 4015 1995
rect 2049 1990 2071 1994
rect 2075 1990 2207 1994
rect 2211 1990 2279 1994
rect 2283 1990 2391 1994
rect 2395 1990 2463 1994
rect 2467 1990 2575 1994
rect 2579 1990 2639 1994
rect 2643 1990 2759 1994
rect 2763 1990 2815 1994
rect 2819 1990 2935 1994
rect 2939 1990 2983 1994
rect 2987 1990 3103 1994
rect 3107 1990 3151 1994
rect 3155 1990 3263 1994
rect 3267 1990 3311 1994
rect 3315 1990 3423 1994
rect 3427 1990 3463 1994
rect 3467 1990 3583 1994
rect 3587 1990 3615 1994
rect 3619 1990 3751 1994
rect 3755 1990 3767 1994
rect 3771 1990 3895 1994
rect 3899 1990 3991 1994
rect 3995 1990 4015 1994
rect 2049 1989 4015 1990
rect 4021 1989 4022 1995
rect 96 1925 97 1931
rect 103 1930 2055 1931
rect 103 1926 111 1930
rect 115 1926 151 1930
rect 155 1926 271 1930
rect 275 1926 303 1930
rect 307 1926 407 1930
rect 411 1926 487 1930
rect 491 1926 543 1930
rect 547 1926 679 1930
rect 683 1926 687 1930
rect 691 1926 823 1930
rect 827 1926 895 1930
rect 899 1926 983 1930
rect 987 1926 1103 1930
rect 1107 1926 1159 1930
rect 1163 1926 1311 1930
rect 1315 1926 1343 1930
rect 1347 1926 1527 1930
rect 1531 1926 1543 1930
rect 1547 1926 1743 1930
rect 1747 1926 1751 1930
rect 1755 1926 1935 1930
rect 1939 1926 2031 1930
rect 2035 1926 2055 1930
rect 103 1925 2055 1926
rect 2061 1925 2062 1931
rect 2054 1909 2055 1915
rect 2061 1914 4027 1915
rect 2061 1910 2071 1914
rect 2075 1910 2279 1914
rect 2283 1910 2407 1914
rect 2411 1910 2463 1914
rect 2467 1910 2639 1914
rect 2643 1910 2655 1914
rect 2659 1910 2815 1914
rect 2819 1910 2887 1914
rect 2891 1910 2983 1914
rect 2987 1910 3103 1914
rect 3107 1910 3151 1914
rect 3155 1910 3311 1914
rect 3315 1910 3463 1914
rect 3467 1910 3511 1914
rect 3515 1910 3615 1914
rect 3619 1910 3711 1914
rect 3715 1910 3767 1914
rect 3771 1910 3895 1914
rect 3899 1910 3991 1914
rect 3995 1910 4027 1914
rect 2061 1909 4027 1910
rect 4033 1909 4034 1915
rect 84 1845 85 1851
rect 91 1850 2043 1851
rect 91 1846 111 1850
rect 115 1846 151 1850
rect 155 1846 271 1850
rect 275 1846 287 1850
rect 291 1846 407 1850
rect 411 1846 447 1850
rect 451 1846 543 1850
rect 547 1846 599 1850
rect 603 1846 679 1850
rect 683 1846 751 1850
rect 755 1846 823 1850
rect 827 1846 919 1850
rect 923 1846 983 1850
rect 987 1846 1103 1850
rect 1107 1846 1159 1850
rect 1163 1846 1303 1850
rect 1307 1846 1343 1850
rect 1347 1846 1511 1850
rect 1515 1846 1543 1850
rect 1547 1846 1735 1850
rect 1739 1846 1751 1850
rect 1755 1846 1935 1850
rect 1939 1846 2031 1850
rect 2035 1846 2043 1850
rect 91 1845 2043 1846
rect 2049 1845 2050 1851
rect 2042 1843 2050 1845
rect 2042 1837 2043 1843
rect 2049 1842 4015 1843
rect 2049 1838 2071 1842
rect 2075 1838 2111 1842
rect 2115 1838 2383 1842
rect 2387 1838 2407 1842
rect 2411 1838 2647 1842
rect 2651 1838 2655 1842
rect 2659 1838 2887 1842
rect 2891 1838 3095 1842
rect 3099 1838 3103 1842
rect 3107 1838 3287 1842
rect 3291 1838 3311 1842
rect 3315 1838 3455 1842
rect 3459 1838 3511 1842
rect 3515 1838 3615 1842
rect 3619 1838 3711 1842
rect 3715 1838 3767 1842
rect 3771 1838 3895 1842
rect 3899 1838 3991 1842
rect 3995 1838 4015 1842
rect 2049 1837 4015 1838
rect 4021 1837 4022 1843
rect 96 1765 97 1771
rect 103 1770 2055 1771
rect 103 1766 111 1770
rect 115 1766 151 1770
rect 155 1766 207 1770
rect 211 1766 287 1770
rect 291 1766 383 1770
rect 387 1766 447 1770
rect 451 1766 567 1770
rect 571 1766 599 1770
rect 603 1766 751 1770
rect 755 1766 919 1770
rect 923 1766 935 1770
rect 939 1766 1103 1770
rect 1107 1766 1111 1770
rect 1115 1766 1279 1770
rect 1283 1766 1303 1770
rect 1307 1766 1455 1770
rect 1459 1766 1511 1770
rect 1515 1766 1631 1770
rect 1635 1766 1735 1770
rect 1739 1766 1935 1770
rect 1939 1766 2031 1770
rect 2035 1766 2055 1770
rect 103 1765 2055 1766
rect 2061 1770 4034 1771
rect 2061 1766 2071 1770
rect 2075 1766 2111 1770
rect 2115 1766 2287 1770
rect 2291 1766 2383 1770
rect 2387 1766 2495 1770
rect 2499 1766 2647 1770
rect 2651 1766 2711 1770
rect 2715 1766 2887 1770
rect 2891 1766 2919 1770
rect 2923 1766 3095 1770
rect 3099 1766 3119 1770
rect 3123 1766 3287 1770
rect 3291 1766 3319 1770
rect 3323 1766 3455 1770
rect 3459 1766 3511 1770
rect 3515 1766 3615 1770
rect 3619 1766 3703 1770
rect 3707 1766 3767 1770
rect 3771 1766 3895 1770
rect 3899 1766 3991 1770
rect 3995 1766 4034 1770
rect 2061 1765 4034 1766
rect 1262 1748 1268 1749
rect 1742 1748 1748 1749
rect 1262 1744 1263 1748
rect 1267 1744 1743 1748
rect 1747 1744 1748 1748
rect 1262 1743 1268 1744
rect 1742 1743 1748 1744
rect 84 1693 85 1699
rect 91 1698 2043 1699
rect 91 1694 111 1698
rect 115 1694 207 1698
rect 211 1694 303 1698
rect 307 1694 383 1698
rect 387 1694 535 1698
rect 539 1694 567 1698
rect 571 1694 751 1698
rect 755 1694 767 1698
rect 771 1694 935 1698
rect 939 1694 983 1698
rect 987 1694 1111 1698
rect 1115 1694 1191 1698
rect 1195 1694 1279 1698
rect 1283 1694 1383 1698
rect 1387 1694 1455 1698
rect 1459 1694 1567 1698
rect 1571 1694 1631 1698
rect 1635 1694 1743 1698
rect 1747 1694 1927 1698
rect 1931 1694 2031 1698
rect 2035 1694 2043 1698
rect 91 1693 2043 1694
rect 2049 1693 2050 1699
rect 2042 1691 2050 1693
rect 2042 1685 2043 1691
rect 2049 1690 4015 1691
rect 2049 1686 2071 1690
rect 2075 1686 2111 1690
rect 2115 1686 2239 1690
rect 2243 1686 2287 1690
rect 2291 1686 2383 1690
rect 2387 1686 2495 1690
rect 2499 1686 2519 1690
rect 2523 1686 2655 1690
rect 2659 1686 2711 1690
rect 2715 1686 2791 1690
rect 2795 1686 2919 1690
rect 2923 1686 2927 1690
rect 2931 1686 3063 1690
rect 3067 1686 3119 1690
rect 3123 1686 3207 1690
rect 3211 1686 3319 1690
rect 3323 1686 3351 1690
rect 3355 1686 3511 1690
rect 3515 1686 3703 1690
rect 3707 1686 3895 1690
rect 3899 1686 3991 1690
rect 3995 1686 4015 1690
rect 2049 1685 4015 1686
rect 4021 1685 4022 1691
rect 96 1617 97 1623
rect 103 1622 2055 1623
rect 103 1618 111 1622
rect 115 1618 303 1622
rect 307 1618 399 1622
rect 403 1618 535 1622
rect 539 1618 575 1622
rect 579 1618 751 1622
rect 755 1618 767 1622
rect 771 1618 935 1622
rect 939 1618 983 1622
rect 987 1618 1111 1622
rect 1115 1618 1191 1622
rect 1195 1618 1279 1622
rect 1283 1618 1383 1622
rect 1387 1618 1447 1622
rect 1451 1618 1567 1622
rect 1571 1618 1607 1622
rect 1611 1618 1743 1622
rect 1747 1618 1767 1622
rect 1771 1618 1927 1622
rect 1931 1618 1935 1622
rect 1939 1618 2031 1622
rect 2035 1618 2055 1622
rect 103 1617 2055 1618
rect 2061 1617 2062 1623
rect 2054 1601 2055 1607
rect 2061 1606 4027 1607
rect 2061 1602 2071 1606
rect 2075 1602 2111 1606
rect 2115 1602 2167 1606
rect 2171 1602 2239 1606
rect 2243 1602 2287 1606
rect 2291 1602 2383 1606
rect 2387 1602 2407 1606
rect 2411 1602 2519 1606
rect 2523 1602 2527 1606
rect 2531 1602 2647 1606
rect 2651 1602 2655 1606
rect 2659 1602 2767 1606
rect 2771 1602 2791 1606
rect 2795 1602 2887 1606
rect 2891 1602 2927 1606
rect 2931 1602 3007 1606
rect 3011 1602 3063 1606
rect 3067 1602 3127 1606
rect 3131 1602 3207 1606
rect 3211 1602 3255 1606
rect 3259 1602 3351 1606
rect 3355 1602 3991 1606
rect 3995 1602 4027 1606
rect 2061 1601 4027 1602
rect 4033 1601 4034 1607
rect 84 1537 85 1543
rect 91 1542 2043 1543
rect 91 1538 111 1542
rect 115 1538 399 1542
rect 403 1538 503 1542
rect 507 1538 575 1542
rect 579 1538 615 1542
rect 619 1538 735 1542
rect 739 1538 751 1542
rect 755 1538 855 1542
rect 859 1538 935 1542
rect 939 1538 967 1542
rect 971 1538 1079 1542
rect 1083 1538 1111 1542
rect 1115 1538 1199 1542
rect 1203 1538 1279 1542
rect 1283 1538 1319 1542
rect 1323 1538 1439 1542
rect 1443 1538 1447 1542
rect 1451 1538 1559 1542
rect 1563 1538 1607 1542
rect 1611 1538 1767 1542
rect 1771 1538 1935 1542
rect 1939 1538 2031 1542
rect 2035 1538 2043 1542
rect 91 1537 2043 1538
rect 2049 1537 2050 1543
rect 2042 1521 2043 1527
rect 2049 1526 4015 1527
rect 2049 1522 2071 1526
rect 2075 1522 2167 1526
rect 2171 1522 2287 1526
rect 2291 1522 2351 1526
rect 2355 1522 2407 1526
rect 2411 1522 2463 1526
rect 2467 1522 2527 1526
rect 2531 1522 2575 1526
rect 2579 1522 2647 1526
rect 2651 1522 2695 1526
rect 2699 1522 2767 1526
rect 2771 1522 2815 1526
rect 2819 1522 2887 1526
rect 2891 1522 2927 1526
rect 2931 1522 3007 1526
rect 3011 1522 3047 1526
rect 3051 1522 3127 1526
rect 3131 1522 3167 1526
rect 3171 1522 3255 1526
rect 3259 1522 3287 1526
rect 3291 1522 3407 1526
rect 3411 1522 3991 1526
rect 3995 1522 4015 1526
rect 2049 1521 4015 1522
rect 4021 1521 4022 1527
rect 2446 1468 2452 1469
rect 2766 1468 2772 1469
rect 2446 1464 2447 1468
rect 2451 1464 2767 1468
rect 2771 1464 2772 1468
rect 2446 1463 2452 1464
rect 2766 1463 2772 1464
rect 96 1453 97 1459
rect 103 1458 2055 1459
rect 103 1454 111 1458
rect 115 1454 503 1458
rect 507 1454 583 1458
rect 587 1454 615 1458
rect 619 1454 687 1458
rect 691 1454 735 1458
rect 739 1454 791 1458
rect 795 1454 855 1458
rect 859 1454 895 1458
rect 899 1454 967 1458
rect 971 1454 999 1458
rect 1003 1454 1079 1458
rect 1083 1454 1103 1458
rect 1107 1454 1199 1458
rect 1203 1454 1207 1458
rect 1211 1454 1311 1458
rect 1315 1454 1319 1458
rect 1323 1454 1415 1458
rect 1419 1454 1439 1458
rect 1443 1454 1519 1458
rect 1523 1454 1559 1458
rect 1563 1454 2031 1458
rect 2035 1454 2055 1458
rect 103 1453 2055 1454
rect 2061 1453 2062 1459
rect 2054 1437 2055 1443
rect 2061 1442 4027 1443
rect 2061 1438 2071 1442
rect 2075 1438 2343 1442
rect 2347 1438 2351 1442
rect 2355 1438 2447 1442
rect 2451 1438 2463 1442
rect 2467 1438 2567 1442
rect 2571 1438 2575 1442
rect 2579 1438 2695 1442
rect 2699 1438 2815 1442
rect 2819 1438 2839 1442
rect 2843 1438 2927 1442
rect 2931 1438 2991 1442
rect 2995 1438 3047 1442
rect 3051 1438 3143 1442
rect 3147 1438 3167 1442
rect 3171 1438 3287 1442
rect 3291 1438 3303 1442
rect 3307 1438 3407 1442
rect 3411 1438 3471 1442
rect 3475 1438 3647 1442
rect 3651 1438 3823 1442
rect 3827 1438 3991 1442
rect 3995 1438 4027 1442
rect 2061 1437 4027 1438
rect 4033 1437 4034 1443
rect 84 1373 85 1379
rect 91 1378 2043 1379
rect 91 1374 111 1378
rect 115 1374 551 1378
rect 555 1374 583 1378
rect 587 1374 655 1378
rect 659 1374 687 1378
rect 691 1374 759 1378
rect 763 1374 791 1378
rect 795 1374 863 1378
rect 867 1374 895 1378
rect 899 1374 975 1378
rect 979 1374 999 1378
rect 1003 1374 1087 1378
rect 1091 1374 1103 1378
rect 1107 1374 1199 1378
rect 1203 1374 1207 1378
rect 1211 1374 1311 1378
rect 1315 1374 1415 1378
rect 1419 1374 1431 1378
rect 1435 1374 1519 1378
rect 1523 1374 1551 1378
rect 1555 1374 2031 1378
rect 2035 1374 2043 1378
rect 91 1373 2043 1374
rect 2049 1373 2050 1379
rect 2042 1357 2043 1363
rect 2049 1362 4015 1363
rect 2049 1358 2071 1362
rect 2075 1358 2287 1362
rect 2291 1358 2343 1362
rect 2347 1358 2407 1362
rect 2411 1358 2447 1362
rect 2451 1358 2543 1362
rect 2547 1358 2567 1362
rect 2571 1358 2695 1362
rect 2699 1358 2839 1362
rect 2843 1358 2855 1362
rect 2859 1358 2991 1362
rect 2995 1358 3015 1362
rect 3019 1358 3143 1362
rect 3147 1358 3183 1362
rect 3187 1358 3303 1362
rect 3307 1358 3351 1362
rect 3355 1358 3471 1362
rect 3475 1358 3519 1362
rect 3523 1358 3647 1362
rect 3651 1358 3687 1362
rect 3691 1358 3823 1362
rect 3827 1358 3855 1362
rect 3859 1358 3991 1362
rect 3995 1358 4015 1362
rect 2049 1357 4015 1358
rect 4021 1357 4022 1363
rect 96 1297 97 1303
rect 103 1302 2055 1303
rect 103 1298 111 1302
rect 115 1298 343 1302
rect 347 1298 463 1302
rect 467 1298 551 1302
rect 555 1298 599 1302
rect 603 1298 655 1302
rect 659 1298 743 1302
rect 747 1298 759 1302
rect 763 1298 863 1302
rect 867 1298 903 1302
rect 907 1298 975 1302
rect 979 1298 1063 1302
rect 1067 1298 1087 1302
rect 1091 1298 1199 1302
rect 1203 1298 1231 1302
rect 1235 1298 1311 1302
rect 1315 1298 1407 1302
rect 1411 1298 1431 1302
rect 1435 1298 1551 1302
rect 1555 1298 1583 1302
rect 1587 1298 2031 1302
rect 2035 1298 2055 1302
rect 103 1297 2055 1298
rect 2061 1297 2062 1303
rect 2054 1277 2055 1283
rect 2061 1282 4027 1283
rect 2061 1278 2071 1282
rect 2075 1278 2127 1282
rect 2131 1278 2287 1282
rect 2291 1278 2295 1282
rect 2299 1278 2407 1282
rect 2411 1278 2479 1282
rect 2483 1278 2543 1282
rect 2547 1278 2679 1282
rect 2683 1278 2695 1282
rect 2699 1278 2855 1282
rect 2859 1278 2879 1282
rect 2883 1278 3015 1282
rect 3019 1278 3071 1282
rect 3075 1278 3183 1282
rect 3187 1278 3247 1282
rect 3251 1278 3351 1282
rect 3355 1278 3415 1282
rect 3419 1278 3519 1282
rect 3523 1278 3583 1282
rect 3587 1278 3687 1282
rect 3691 1278 3751 1282
rect 3755 1278 3855 1282
rect 3859 1278 3895 1282
rect 3899 1278 3991 1282
rect 3995 1278 4027 1282
rect 2061 1277 4027 1278
rect 4033 1277 4034 1283
rect 84 1225 85 1231
rect 91 1230 2043 1231
rect 91 1226 111 1230
rect 115 1226 183 1230
rect 187 1226 343 1230
rect 347 1226 351 1230
rect 355 1226 463 1230
rect 467 1226 535 1230
rect 539 1226 599 1230
rect 603 1226 727 1230
rect 731 1226 743 1230
rect 747 1226 903 1230
rect 907 1226 919 1230
rect 923 1226 1063 1230
rect 1067 1226 1103 1230
rect 1107 1226 1231 1230
rect 1235 1226 1287 1230
rect 1291 1226 1407 1230
rect 1411 1226 1471 1230
rect 1475 1226 1583 1230
rect 1587 1226 1655 1230
rect 1659 1226 1839 1230
rect 1843 1226 2031 1230
rect 2035 1226 2043 1230
rect 91 1225 2043 1226
rect 2049 1225 2050 1231
rect 2042 1193 2043 1199
rect 2049 1198 4015 1199
rect 2049 1194 2071 1198
rect 2075 1194 2111 1198
rect 2115 1194 2127 1198
rect 2131 1194 2247 1198
rect 2251 1194 2295 1198
rect 2299 1194 2407 1198
rect 2411 1194 2479 1198
rect 2483 1194 2559 1198
rect 2563 1194 2679 1198
rect 2683 1194 2703 1198
rect 2707 1194 2863 1198
rect 2867 1194 2879 1198
rect 2883 1194 3039 1198
rect 3043 1194 3071 1198
rect 3075 1194 3239 1198
rect 3243 1194 3247 1198
rect 3251 1194 3415 1198
rect 3419 1194 3455 1198
rect 3459 1194 3583 1198
rect 3587 1194 3687 1198
rect 3691 1194 3751 1198
rect 3755 1194 3895 1198
rect 3899 1194 3991 1198
rect 3995 1194 4015 1198
rect 2049 1193 4015 1194
rect 4021 1193 4022 1199
rect 96 1145 97 1151
rect 103 1150 2055 1151
rect 103 1146 111 1150
rect 115 1146 151 1150
rect 155 1146 183 1150
rect 187 1146 303 1150
rect 307 1146 351 1150
rect 355 1146 495 1150
rect 499 1146 535 1150
rect 539 1146 703 1150
rect 707 1146 727 1150
rect 731 1146 911 1150
rect 915 1146 919 1150
rect 923 1146 1103 1150
rect 1107 1146 1119 1150
rect 1123 1146 1287 1150
rect 1291 1146 1319 1150
rect 1323 1146 1471 1150
rect 1475 1146 1519 1150
rect 1523 1146 1655 1150
rect 1659 1146 1719 1150
rect 1723 1146 1839 1150
rect 1843 1146 1919 1150
rect 1923 1146 2031 1150
rect 2035 1146 2055 1150
rect 103 1145 2055 1146
rect 2061 1145 2062 1151
rect 2054 1117 2055 1123
rect 2061 1122 4027 1123
rect 2061 1118 2071 1122
rect 2075 1118 2111 1122
rect 2115 1118 2247 1122
rect 2251 1118 2303 1122
rect 2307 1118 2407 1122
rect 2411 1118 2511 1122
rect 2515 1118 2559 1122
rect 2563 1118 2703 1122
rect 2707 1118 2863 1122
rect 2867 1118 2895 1122
rect 2899 1118 3039 1122
rect 3043 1118 3087 1122
rect 3091 1118 3239 1122
rect 3243 1118 3287 1122
rect 3291 1118 3455 1122
rect 3459 1118 3495 1122
rect 3499 1118 3687 1122
rect 3691 1118 3703 1122
rect 3707 1118 3895 1122
rect 3899 1118 3991 1122
rect 3995 1118 4027 1122
rect 2061 1117 4027 1118
rect 4033 1117 4034 1123
rect 84 1065 85 1071
rect 91 1070 2043 1071
rect 91 1066 111 1070
rect 115 1066 151 1070
rect 155 1066 279 1070
rect 283 1066 303 1070
rect 307 1066 447 1070
rect 451 1066 495 1070
rect 499 1066 623 1070
rect 627 1066 703 1070
rect 707 1066 799 1070
rect 803 1066 911 1070
rect 915 1066 967 1070
rect 971 1066 1119 1070
rect 1123 1066 1127 1070
rect 1131 1066 1279 1070
rect 1283 1066 1319 1070
rect 1323 1066 1423 1070
rect 1427 1066 1519 1070
rect 1523 1066 1559 1070
rect 1563 1066 1695 1070
rect 1699 1066 1719 1070
rect 1723 1066 1823 1070
rect 1827 1066 1919 1070
rect 1923 1066 1935 1070
rect 1939 1066 2031 1070
rect 2035 1066 2043 1070
rect 91 1065 2043 1066
rect 2049 1065 2050 1071
rect 2042 1029 2043 1035
rect 2049 1034 4015 1035
rect 2049 1030 2071 1034
rect 2075 1030 2111 1034
rect 2115 1030 2303 1034
rect 2307 1030 2319 1034
rect 2323 1030 2487 1034
rect 2491 1030 2511 1034
rect 2515 1030 2663 1034
rect 2667 1030 2703 1034
rect 2707 1030 2847 1034
rect 2851 1030 2895 1034
rect 2899 1030 3039 1034
rect 3043 1030 3087 1034
rect 3091 1030 3247 1034
rect 3251 1030 3287 1034
rect 3291 1030 3463 1034
rect 3467 1030 3495 1034
rect 3499 1030 3687 1034
rect 3691 1030 3703 1034
rect 3707 1030 3895 1034
rect 3899 1030 3991 1034
rect 3995 1030 4015 1034
rect 2049 1029 4015 1030
rect 4021 1029 4022 1035
rect 96 981 97 987
rect 103 986 2055 987
rect 103 982 111 986
rect 115 982 151 986
rect 155 982 279 986
rect 283 982 287 986
rect 291 982 447 986
rect 451 982 471 986
rect 475 982 623 986
rect 627 982 671 986
rect 675 982 799 986
rect 803 982 871 986
rect 875 982 967 986
rect 971 982 1079 986
rect 1083 982 1127 986
rect 1131 982 1279 986
rect 1283 982 1287 986
rect 1291 982 1423 986
rect 1427 982 1495 986
rect 1499 982 1559 986
rect 1563 982 1695 986
rect 1699 982 1703 986
rect 1707 982 1823 986
rect 1827 982 1911 986
rect 1915 982 1935 986
rect 1939 982 2031 986
rect 2035 982 2055 986
rect 103 981 2055 982
rect 2061 981 2062 987
rect 654 972 660 973
rect 934 972 940 973
rect 654 968 655 972
rect 659 968 935 972
rect 939 968 940 972
rect 654 967 660 968
rect 934 967 940 968
rect 2054 953 2055 959
rect 2061 958 4027 959
rect 2061 954 2071 958
rect 2075 954 2151 958
rect 2155 954 2287 958
rect 2291 954 2319 958
rect 2323 954 2431 958
rect 2435 954 2487 958
rect 2491 954 2591 958
rect 2595 954 2663 958
rect 2667 954 2759 958
rect 2763 954 2847 958
rect 2851 954 2935 958
rect 2939 954 3039 958
rect 3043 954 3119 958
rect 3123 954 3247 958
rect 3251 954 3311 958
rect 3315 954 3463 958
rect 3467 954 3511 958
rect 3515 954 3687 958
rect 3691 954 3711 958
rect 3715 954 3895 958
rect 3899 954 3991 958
rect 3995 954 4027 958
rect 2061 953 4027 954
rect 4033 953 4034 959
rect 84 901 85 907
rect 91 906 2043 907
rect 91 902 111 906
rect 115 902 151 906
rect 155 902 287 906
rect 291 902 319 906
rect 323 902 471 906
rect 475 902 519 906
rect 523 902 671 906
rect 675 902 727 906
rect 731 902 871 906
rect 875 902 935 906
rect 939 902 1079 906
rect 1083 902 1143 906
rect 1147 902 1287 906
rect 1291 902 1335 906
rect 1339 902 1495 906
rect 1499 902 1527 906
rect 1531 902 1703 906
rect 1707 902 1719 906
rect 1723 902 1911 906
rect 1915 902 2031 906
rect 2035 902 2043 906
rect 91 901 2043 902
rect 2049 901 2050 907
rect 2042 869 2043 875
rect 2049 874 4015 875
rect 2049 870 2071 874
rect 2075 870 2111 874
rect 2115 870 2151 874
rect 2155 870 2239 874
rect 2243 870 2287 874
rect 2291 870 2407 874
rect 2411 870 2431 874
rect 2435 870 2575 874
rect 2579 870 2591 874
rect 2595 870 2751 874
rect 2755 870 2759 874
rect 2763 870 2935 874
rect 2939 870 3119 874
rect 3123 870 3311 874
rect 3315 870 3511 874
rect 3515 870 3711 874
rect 3715 870 3895 874
rect 3899 870 3991 874
rect 3995 870 4015 874
rect 2049 869 4015 870
rect 4021 869 4022 875
rect 96 817 97 823
rect 103 822 2055 823
rect 103 818 111 822
rect 115 818 151 822
rect 155 818 263 822
rect 267 818 319 822
rect 323 818 367 822
rect 371 818 479 822
rect 483 818 519 822
rect 523 818 591 822
rect 595 818 711 822
rect 715 818 727 822
rect 731 818 855 822
rect 859 818 935 822
rect 939 818 1031 822
rect 1035 818 1143 822
rect 1147 818 1239 822
rect 1243 818 1335 822
rect 1339 818 1471 822
rect 1475 818 1527 822
rect 1531 818 1711 822
rect 1715 818 1719 822
rect 1723 818 1911 822
rect 1915 818 1935 822
rect 1939 818 2031 822
rect 2035 818 2055 822
rect 103 817 2055 818
rect 2061 817 2062 823
rect 2054 797 2055 803
rect 2061 802 4027 803
rect 2061 798 2071 802
rect 2075 798 2111 802
rect 2115 798 2239 802
rect 2243 798 2391 802
rect 2395 798 2407 802
rect 2411 798 2575 802
rect 2579 798 2679 802
rect 2683 798 2751 802
rect 2755 798 2935 802
rect 2939 798 2951 802
rect 2955 798 3119 802
rect 3123 798 3199 802
rect 3203 798 3311 802
rect 3315 798 3439 802
rect 3443 798 3511 802
rect 3515 798 3671 802
rect 3675 798 3711 802
rect 3715 798 3895 802
rect 3899 798 3991 802
rect 3995 798 4027 802
rect 2061 797 4027 798
rect 4033 797 4034 803
rect 84 741 85 747
rect 91 746 2043 747
rect 91 742 111 746
rect 115 742 263 746
rect 267 742 367 746
rect 371 742 423 746
rect 427 742 479 746
rect 483 742 527 746
rect 531 742 591 746
rect 595 742 639 746
rect 643 742 711 746
rect 715 742 759 746
rect 763 742 855 746
rect 859 742 879 746
rect 883 742 1007 746
rect 1011 742 1031 746
rect 1035 742 1143 746
rect 1147 742 1239 746
rect 1243 742 1287 746
rect 1291 742 1447 746
rect 1451 742 1471 746
rect 1475 742 1615 746
rect 1619 742 1711 746
rect 1715 742 1783 746
rect 1787 742 1935 746
rect 1939 742 2031 746
rect 2035 742 2043 746
rect 91 741 2043 742
rect 2049 741 2050 747
rect 2042 717 2043 723
rect 2049 722 4015 723
rect 2049 718 2071 722
rect 2075 718 2111 722
rect 2115 718 2327 722
rect 2331 718 2391 722
rect 2395 718 2551 722
rect 2555 718 2679 722
rect 2683 718 2775 722
rect 2779 718 2951 722
rect 2955 718 2991 722
rect 2995 718 3199 722
rect 3203 718 3207 722
rect 3211 718 3415 722
rect 3419 718 3439 722
rect 3443 718 3623 722
rect 3627 718 3671 722
rect 3675 718 3831 722
rect 3835 718 3895 722
rect 3899 718 3991 722
rect 3995 718 4015 722
rect 2049 717 4015 718
rect 4021 717 4022 723
rect 96 657 97 663
rect 103 662 2055 663
rect 103 658 111 662
rect 115 658 423 662
rect 427 658 527 662
rect 531 658 591 662
rect 595 658 639 662
rect 643 658 695 662
rect 699 658 759 662
rect 763 658 807 662
rect 811 658 879 662
rect 883 658 919 662
rect 923 658 1007 662
rect 1011 658 1031 662
rect 1035 658 1143 662
rect 1147 658 1263 662
rect 1267 658 1287 662
rect 1291 658 1383 662
rect 1387 658 1447 662
rect 1451 658 1503 662
rect 1507 658 1615 662
rect 1619 658 1623 662
rect 1627 658 1783 662
rect 1787 658 1935 662
rect 1939 658 2031 662
rect 2035 658 2055 662
rect 103 657 2055 658
rect 2061 657 2062 663
rect 2054 641 2055 647
rect 2061 646 4027 647
rect 2061 642 2071 646
rect 2075 642 2111 646
rect 2115 642 2127 646
rect 2131 642 2295 646
rect 2299 642 2327 646
rect 2331 642 2455 646
rect 2459 642 2551 646
rect 2555 642 2615 646
rect 2619 642 2775 646
rect 2779 642 2783 646
rect 2787 642 2951 646
rect 2955 642 2991 646
rect 2995 642 3127 646
rect 3131 642 3207 646
rect 3211 642 3303 646
rect 3307 642 3415 646
rect 3419 642 3487 646
rect 3491 642 3623 646
rect 3627 642 3679 646
rect 3683 642 3831 646
rect 3835 642 3879 646
rect 3883 642 3991 646
rect 3995 642 4027 646
rect 2061 641 4027 642
rect 4033 641 4034 647
rect 84 577 85 583
rect 91 582 2043 583
rect 91 578 111 582
rect 115 578 591 582
rect 595 578 663 582
rect 667 578 695 582
rect 699 578 775 582
rect 779 578 807 582
rect 811 578 895 582
rect 899 578 919 582
rect 923 578 1023 582
rect 1027 578 1031 582
rect 1035 578 1143 582
rect 1147 578 1159 582
rect 1163 578 1263 582
rect 1267 578 1303 582
rect 1307 578 1383 582
rect 1387 578 1447 582
rect 1451 578 1503 582
rect 1507 578 1591 582
rect 1595 578 1623 582
rect 1627 578 1735 582
rect 1739 578 1879 582
rect 1883 578 2031 582
rect 2035 578 2043 582
rect 91 577 2043 578
rect 2049 577 2050 583
rect 2042 561 2043 567
rect 2049 566 4015 567
rect 2049 562 2071 566
rect 2075 562 2127 566
rect 2131 562 2295 566
rect 2299 562 2303 566
rect 2307 562 2447 566
rect 2451 562 2455 566
rect 2459 562 2591 566
rect 2595 562 2615 566
rect 2619 562 2735 566
rect 2739 562 2783 566
rect 2787 562 2879 566
rect 2883 562 2951 566
rect 2955 562 3031 566
rect 3035 562 3127 566
rect 3131 562 3183 566
rect 3187 562 3303 566
rect 3307 562 3335 566
rect 3339 562 3487 566
rect 3491 562 3495 566
rect 3499 562 3655 566
rect 3659 562 3679 566
rect 3683 562 3823 566
rect 3827 562 3879 566
rect 3883 562 3991 566
rect 3995 562 4015 566
rect 2049 561 4015 562
rect 4021 561 4022 567
rect 3166 508 3172 509
rect 3566 508 3572 509
rect 3166 504 3167 508
rect 3171 504 3567 508
rect 3571 504 3572 508
rect 3166 503 3172 504
rect 3566 503 3572 504
rect 96 489 97 495
rect 103 494 2055 495
rect 103 490 111 494
rect 115 490 535 494
rect 539 490 639 494
rect 643 490 663 494
rect 667 490 743 494
rect 747 490 775 494
rect 779 490 847 494
rect 851 490 895 494
rect 899 490 967 494
rect 971 490 1023 494
rect 1027 490 1103 494
rect 1107 490 1159 494
rect 1163 490 1255 494
rect 1259 490 1303 494
rect 1307 490 1415 494
rect 1419 490 1447 494
rect 1451 490 1591 494
rect 1595 490 1735 494
rect 1739 490 1775 494
rect 1779 490 1879 494
rect 1883 490 1935 494
rect 1939 490 2031 494
rect 2035 490 2055 494
rect 103 489 2055 490
rect 2061 489 2062 495
rect 2054 487 2062 489
rect 2054 481 2055 487
rect 2061 486 4027 487
rect 2061 482 2071 486
rect 2075 482 2303 486
rect 2307 482 2447 486
rect 2451 482 2511 486
rect 2515 482 2591 486
rect 2595 482 2615 486
rect 2619 482 2735 486
rect 2739 482 2863 486
rect 2867 482 2879 486
rect 2883 482 3007 486
rect 3011 482 3031 486
rect 3035 482 3159 486
rect 3163 482 3183 486
rect 3187 482 3319 486
rect 3323 482 3335 486
rect 3339 482 3479 486
rect 3483 482 3495 486
rect 3499 482 3647 486
rect 3651 482 3655 486
rect 3659 482 3823 486
rect 3827 482 3991 486
rect 3995 482 4027 486
rect 2061 481 4027 482
rect 4033 481 4034 487
rect 1238 476 1244 477
rect 1598 476 1604 477
rect 1238 472 1239 476
rect 1243 472 1599 476
rect 1603 472 1604 476
rect 1238 471 1244 472
rect 1598 471 1604 472
rect 84 413 85 419
rect 91 418 2043 419
rect 91 414 111 418
rect 115 414 495 418
rect 499 414 535 418
rect 539 414 631 418
rect 635 414 639 418
rect 643 414 743 418
rect 747 414 767 418
rect 771 414 847 418
rect 851 414 911 418
rect 915 414 967 418
rect 971 414 1047 418
rect 1051 414 1103 418
rect 1107 414 1183 418
rect 1187 414 1255 418
rect 1259 414 1319 418
rect 1323 414 1415 418
rect 1419 414 1447 418
rect 1451 414 1575 418
rect 1579 414 1591 418
rect 1595 414 1703 418
rect 1707 414 1775 418
rect 1779 414 1831 418
rect 1835 414 1935 418
rect 1939 414 2031 418
rect 2035 414 2043 418
rect 91 413 2043 414
rect 2049 413 2050 419
rect 2042 397 2043 403
rect 2049 402 4015 403
rect 2049 398 2071 402
rect 2075 398 2511 402
rect 2515 398 2591 402
rect 2595 398 2615 402
rect 2619 398 2695 402
rect 2699 398 2735 402
rect 2739 398 2815 402
rect 2819 398 2863 402
rect 2867 398 2959 402
rect 2963 398 3007 402
rect 3011 398 3119 402
rect 3123 398 3159 402
rect 3163 398 3303 402
rect 3307 398 3319 402
rect 3323 398 3479 402
rect 3483 398 3503 402
rect 3507 398 3647 402
rect 3651 398 3711 402
rect 3715 398 3823 402
rect 3827 398 3895 402
rect 3899 398 3991 402
rect 3995 398 4015 402
rect 2049 397 4015 398
rect 4021 397 4022 403
rect 96 329 97 335
rect 103 334 2055 335
rect 103 330 111 334
rect 115 330 335 334
rect 339 330 463 334
rect 467 330 495 334
rect 499 330 607 334
rect 611 330 631 334
rect 635 330 767 334
rect 771 330 911 334
rect 915 330 943 334
rect 947 330 1047 334
rect 1051 330 1127 334
rect 1131 330 1183 334
rect 1187 330 1311 334
rect 1315 330 1319 334
rect 1323 330 1447 334
rect 1451 330 1503 334
rect 1507 330 1575 334
rect 1579 330 1703 334
rect 1707 330 1831 334
rect 1835 330 1903 334
rect 1907 330 1935 334
rect 1939 330 2031 334
rect 2035 330 2055 334
rect 103 329 2055 330
rect 2061 331 2062 335
rect 2061 330 4034 331
rect 2061 329 2071 330
rect 2054 326 2071 329
rect 2075 326 2111 330
rect 2115 326 2271 330
rect 2275 326 2455 330
rect 2459 326 2591 330
rect 2595 326 2631 330
rect 2635 326 2695 330
rect 2699 326 2807 330
rect 2811 326 2815 330
rect 2819 326 2959 330
rect 2963 326 2999 330
rect 3003 326 3119 330
rect 3123 326 3215 330
rect 3219 326 3303 330
rect 3307 326 3439 330
rect 3443 326 3503 330
rect 3507 326 3679 330
rect 3683 326 3711 330
rect 3715 326 3895 330
rect 3899 326 3991 330
rect 3995 326 4034 330
rect 2054 325 4034 326
rect 2982 316 2988 317
rect 3510 316 3516 317
rect 2982 312 2983 316
rect 2987 312 3511 316
rect 3515 312 3516 316
rect 2982 311 2988 312
rect 3510 311 3516 312
rect 2042 258 4022 259
rect 2042 255 2071 258
rect 84 249 85 255
rect 91 254 2043 255
rect 91 250 111 254
rect 115 250 151 254
rect 155 250 279 254
rect 283 250 335 254
rect 339 250 431 254
rect 435 250 463 254
rect 467 250 599 254
rect 603 250 607 254
rect 611 250 767 254
rect 771 250 783 254
rect 787 250 943 254
rect 947 250 975 254
rect 979 250 1127 254
rect 1131 250 1175 254
rect 1179 250 1311 254
rect 1315 250 1375 254
rect 1379 250 1503 254
rect 1507 250 1583 254
rect 1587 250 1703 254
rect 1707 250 1799 254
rect 1803 250 1903 254
rect 1907 250 2031 254
rect 2035 250 2043 254
rect 91 249 2043 250
rect 2049 254 2071 255
rect 2075 254 2111 258
rect 2115 254 2271 258
rect 2275 254 2455 258
rect 2459 254 2471 258
rect 2475 254 2631 258
rect 2635 254 2687 258
rect 2691 254 2807 258
rect 2811 254 2903 258
rect 2907 254 2999 258
rect 3003 254 3111 258
rect 3115 254 3215 258
rect 3219 254 3319 258
rect 3323 254 3439 258
rect 3443 254 3519 258
rect 3523 254 3679 258
rect 3683 254 3719 258
rect 3723 254 3895 258
rect 3899 254 3991 258
rect 3995 254 4022 258
rect 2049 253 4022 254
rect 2049 249 2050 253
rect 96 153 97 159
rect 103 158 2055 159
rect 103 154 111 158
rect 115 154 151 158
rect 155 154 255 158
rect 259 154 279 158
rect 283 154 359 158
rect 363 154 431 158
rect 435 154 471 158
rect 475 154 599 158
rect 603 154 607 158
rect 611 154 743 158
rect 747 154 783 158
rect 787 154 879 158
rect 883 154 975 158
rect 979 154 1015 158
rect 1019 154 1151 158
rect 1155 154 1175 158
rect 1179 154 1279 158
rect 1283 154 1375 158
rect 1379 154 1399 158
rect 1403 154 1519 158
rect 1523 154 1583 158
rect 1587 154 1647 158
rect 1651 154 1775 158
rect 1779 154 1799 158
rect 1803 154 2031 158
rect 2035 154 2055 158
rect 103 153 2055 154
rect 2061 158 4034 159
rect 2061 154 2071 158
rect 2075 154 2111 158
rect 2115 154 2215 158
rect 2219 154 2271 158
rect 2275 154 2319 158
rect 2323 154 2423 158
rect 2427 154 2471 158
rect 2475 154 2527 158
rect 2531 154 2655 158
rect 2659 154 2687 158
rect 2691 154 2775 158
rect 2779 154 2895 158
rect 2899 154 2903 158
rect 2907 154 3015 158
rect 3019 154 3111 158
rect 3115 154 3135 158
rect 3139 154 3247 158
rect 3251 154 3319 158
rect 3323 154 3359 158
rect 3363 154 3471 158
rect 3475 154 3519 158
rect 3523 154 3583 158
rect 3587 154 3687 158
rect 3691 154 3719 158
rect 3723 154 3791 158
rect 3795 154 3895 158
rect 3899 154 3991 158
rect 3995 154 4034 158
rect 2061 153 4034 154
rect 84 81 85 87
rect 91 86 2043 87
rect 91 82 111 86
rect 115 82 151 86
rect 155 82 255 86
rect 259 82 359 86
rect 363 82 471 86
rect 475 82 607 86
rect 611 82 743 86
rect 747 82 879 86
rect 883 82 1015 86
rect 1019 82 1151 86
rect 1155 82 1279 86
rect 1283 82 1399 86
rect 1403 82 1519 86
rect 1523 82 1647 86
rect 1651 82 1775 86
rect 1779 82 2031 86
rect 2035 82 2043 86
rect 91 81 2043 82
rect 2049 86 4022 87
rect 2049 82 2071 86
rect 2075 82 2111 86
rect 2115 82 2215 86
rect 2219 82 2319 86
rect 2323 82 2423 86
rect 2427 82 2527 86
rect 2531 82 2655 86
rect 2659 82 2775 86
rect 2779 82 2895 86
rect 2899 82 3015 86
rect 3019 82 3135 86
rect 3139 82 3247 86
rect 3251 82 3359 86
rect 3363 82 3471 86
rect 3475 82 3583 86
rect 3587 82 3687 86
rect 3691 82 3791 86
rect 3795 82 3895 86
rect 3899 82 3991 86
rect 3995 82 4022 86
rect 2049 81 4022 82
<< m5c >>
rect 85 4061 91 4067
rect 2043 4061 2049 4067
rect 97 3985 103 3991
rect 2055 3985 2061 3991
rect 85 3913 91 3919
rect 2043 3913 2049 3919
rect 97 3841 103 3847
rect 2055 3841 2061 3847
rect 2043 3773 2049 3779
rect 4015 3773 4021 3779
rect 85 3757 91 3763
rect 2043 3757 2049 3763
rect 2055 3689 2061 3695
rect 4027 3689 4033 3695
rect 97 3681 103 3687
rect 2055 3681 2061 3687
rect 85 3609 91 3615
rect 2043 3609 2049 3615
rect 97 3525 103 3531
rect 2055 3525 2061 3531
rect 85 3453 91 3459
rect 2043 3453 2049 3459
rect 97 3357 103 3363
rect 2055 3357 2061 3363
rect 2043 3285 2049 3291
rect 4015 3285 4021 3291
rect 85 3277 91 3283
rect 2043 3277 2049 3283
rect 2055 3213 2061 3219
rect 4027 3213 4033 3219
rect 97 3201 103 3207
rect 2055 3201 2061 3207
rect 85 3129 91 3135
rect 2043 3129 2049 3135
rect 97 3049 103 3055
rect 2055 3049 2061 3055
rect 2043 2981 2049 2987
rect 4015 2981 4021 2987
rect 85 2969 91 2975
rect 2043 2969 2049 2975
rect 2055 2901 2061 2907
rect 4027 2901 4033 2907
rect 97 2885 103 2891
rect 2055 2885 2061 2891
rect 2043 2817 2049 2823
rect 4015 2817 4021 2823
rect 85 2801 91 2807
rect 2043 2801 2049 2807
rect 2055 2733 2061 2739
rect 4027 2733 4033 2739
rect 97 2725 103 2731
rect 2055 2725 2061 2731
rect 85 2645 91 2651
rect 2043 2645 2049 2651
rect 97 2569 103 2575
rect 2055 2569 2061 2575
rect 85 2497 91 2503
rect 2043 2497 2049 2503
rect 2043 2485 2049 2491
rect 4015 2485 4021 2491
rect 97 2417 103 2423
rect 2055 2417 2061 2423
rect 2055 2401 2061 2407
rect 4027 2401 4033 2407
rect 85 2337 91 2343
rect 2043 2337 2049 2343
rect 2043 2317 2049 2323
rect 4015 2317 4021 2323
rect 97 2253 103 2259
rect 2055 2253 2061 2259
rect 2055 2237 2061 2243
rect 4027 2237 4033 2243
rect 85 2169 91 2175
rect 2043 2169 2049 2175
rect 2043 2157 2049 2163
rect 4015 2157 4021 2163
rect 97 2089 103 2095
rect 2055 2089 2061 2095
rect 2055 2073 2061 2079
rect 4027 2073 4033 2079
rect 85 2009 91 2015
rect 2043 2009 2049 2015
rect 2043 1989 2049 1995
rect 4015 1989 4021 1995
rect 97 1925 103 1931
rect 2055 1925 2061 1931
rect 2055 1909 2061 1915
rect 4027 1909 4033 1915
rect 85 1845 91 1851
rect 2043 1845 2049 1851
rect 2043 1837 2049 1843
rect 4015 1837 4021 1843
rect 97 1765 103 1771
rect 2055 1765 2061 1771
rect 85 1693 91 1699
rect 2043 1693 2049 1699
rect 2043 1685 2049 1691
rect 4015 1685 4021 1691
rect 97 1617 103 1623
rect 2055 1617 2061 1623
rect 2055 1601 2061 1607
rect 4027 1601 4033 1607
rect 85 1537 91 1543
rect 2043 1537 2049 1543
rect 2043 1521 2049 1527
rect 4015 1521 4021 1527
rect 97 1453 103 1459
rect 2055 1453 2061 1459
rect 2055 1437 2061 1443
rect 4027 1437 4033 1443
rect 85 1373 91 1379
rect 2043 1373 2049 1379
rect 2043 1357 2049 1363
rect 4015 1357 4021 1363
rect 97 1297 103 1303
rect 2055 1297 2061 1303
rect 2055 1277 2061 1283
rect 4027 1277 4033 1283
rect 85 1225 91 1231
rect 2043 1225 2049 1231
rect 2043 1193 2049 1199
rect 4015 1193 4021 1199
rect 97 1145 103 1151
rect 2055 1145 2061 1151
rect 2055 1117 2061 1123
rect 4027 1117 4033 1123
rect 85 1065 91 1071
rect 2043 1065 2049 1071
rect 2043 1029 2049 1035
rect 4015 1029 4021 1035
rect 97 981 103 987
rect 2055 981 2061 987
rect 2055 953 2061 959
rect 4027 953 4033 959
rect 85 901 91 907
rect 2043 901 2049 907
rect 2043 869 2049 875
rect 4015 869 4021 875
rect 97 817 103 823
rect 2055 817 2061 823
rect 2055 797 2061 803
rect 4027 797 4033 803
rect 85 741 91 747
rect 2043 741 2049 747
rect 2043 717 2049 723
rect 4015 717 4021 723
rect 97 657 103 663
rect 2055 657 2061 663
rect 2055 641 2061 647
rect 4027 641 4033 647
rect 85 577 91 583
rect 2043 577 2049 583
rect 2043 561 2049 567
rect 4015 561 4021 567
rect 97 489 103 495
rect 2055 489 2061 495
rect 2055 481 2061 487
rect 4027 481 4033 487
rect 85 413 91 419
rect 2043 413 2049 419
rect 2043 397 2049 403
rect 4015 397 4021 403
rect 97 329 103 335
rect 2055 329 2061 335
rect 85 249 91 255
rect 2043 249 2049 255
rect 97 153 103 159
rect 2055 153 2061 159
rect 85 81 91 87
rect 2043 81 2049 87
<< m5 >>
rect 84 4067 92 4104
rect 84 4061 85 4067
rect 91 4061 92 4067
rect 84 3919 92 4061
rect 84 3913 85 3919
rect 91 3913 92 3919
rect 84 3763 92 3913
rect 84 3757 85 3763
rect 91 3757 92 3763
rect 84 3615 92 3757
rect 84 3609 85 3615
rect 91 3609 92 3615
rect 84 3459 92 3609
rect 84 3453 85 3459
rect 91 3453 92 3459
rect 84 3283 92 3453
rect 84 3277 85 3283
rect 91 3277 92 3283
rect 84 3135 92 3277
rect 84 3129 85 3135
rect 91 3129 92 3135
rect 84 2975 92 3129
rect 84 2969 85 2975
rect 91 2969 92 2975
rect 84 2807 92 2969
rect 84 2801 85 2807
rect 91 2801 92 2807
rect 84 2651 92 2801
rect 84 2645 85 2651
rect 91 2645 92 2651
rect 84 2503 92 2645
rect 84 2497 85 2503
rect 91 2497 92 2503
rect 84 2343 92 2497
rect 84 2337 85 2343
rect 91 2337 92 2343
rect 84 2175 92 2337
rect 84 2169 85 2175
rect 91 2169 92 2175
rect 84 2015 92 2169
rect 84 2009 85 2015
rect 91 2009 92 2015
rect 84 1851 92 2009
rect 84 1845 85 1851
rect 91 1845 92 1851
rect 84 1699 92 1845
rect 84 1693 85 1699
rect 91 1693 92 1699
rect 84 1543 92 1693
rect 84 1537 85 1543
rect 91 1537 92 1543
rect 84 1379 92 1537
rect 84 1373 85 1379
rect 91 1373 92 1379
rect 84 1231 92 1373
rect 84 1225 85 1231
rect 91 1225 92 1231
rect 84 1071 92 1225
rect 84 1065 85 1071
rect 91 1065 92 1071
rect 84 907 92 1065
rect 84 901 85 907
rect 91 901 92 907
rect 84 747 92 901
rect 84 741 85 747
rect 91 741 92 747
rect 84 583 92 741
rect 84 577 85 583
rect 91 577 92 583
rect 84 419 92 577
rect 84 413 85 419
rect 91 413 92 419
rect 84 255 92 413
rect 84 249 85 255
rect 91 249 92 255
rect 84 87 92 249
rect 84 81 85 87
rect 91 81 92 87
rect 84 72 92 81
rect 96 3991 104 4104
rect 96 3985 97 3991
rect 103 3985 104 3991
rect 96 3847 104 3985
rect 96 3841 97 3847
rect 103 3841 104 3847
rect 96 3687 104 3841
rect 96 3681 97 3687
rect 103 3681 104 3687
rect 96 3531 104 3681
rect 96 3525 97 3531
rect 103 3525 104 3531
rect 96 3363 104 3525
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3207 104 3357
rect 96 3201 97 3207
rect 103 3201 104 3207
rect 96 3055 104 3201
rect 96 3049 97 3055
rect 103 3049 104 3055
rect 96 2891 104 3049
rect 96 2885 97 2891
rect 103 2885 104 2891
rect 96 2731 104 2885
rect 96 2725 97 2731
rect 103 2725 104 2731
rect 96 2575 104 2725
rect 96 2569 97 2575
rect 103 2569 104 2575
rect 96 2423 104 2569
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2259 104 2417
rect 96 2253 97 2259
rect 103 2253 104 2259
rect 96 2095 104 2253
rect 96 2089 97 2095
rect 103 2089 104 2095
rect 96 1931 104 2089
rect 96 1925 97 1931
rect 103 1925 104 1931
rect 96 1771 104 1925
rect 96 1765 97 1771
rect 103 1765 104 1771
rect 96 1623 104 1765
rect 96 1617 97 1623
rect 103 1617 104 1623
rect 96 1459 104 1617
rect 96 1453 97 1459
rect 103 1453 104 1459
rect 96 1303 104 1453
rect 96 1297 97 1303
rect 103 1297 104 1303
rect 96 1151 104 1297
rect 96 1145 97 1151
rect 103 1145 104 1151
rect 96 987 104 1145
rect 96 981 97 987
rect 103 981 104 987
rect 96 823 104 981
rect 96 817 97 823
rect 103 817 104 823
rect 96 663 104 817
rect 96 657 97 663
rect 103 657 104 663
rect 96 495 104 657
rect 96 489 97 495
rect 103 489 104 495
rect 96 335 104 489
rect 96 329 97 335
rect 103 329 104 335
rect 96 159 104 329
rect 96 153 97 159
rect 103 153 104 159
rect 96 72 104 153
rect 2042 4067 2050 4104
rect 2042 4061 2043 4067
rect 2049 4061 2050 4067
rect 2042 3919 2050 4061
rect 2042 3913 2043 3919
rect 2049 3913 2050 3919
rect 2042 3779 2050 3913
rect 2042 3773 2043 3779
rect 2049 3773 2050 3779
rect 2042 3763 2050 3773
rect 2042 3757 2043 3763
rect 2049 3757 2050 3763
rect 2042 3615 2050 3757
rect 2042 3609 2043 3615
rect 2049 3609 2050 3615
rect 2042 3459 2050 3609
rect 2042 3453 2043 3459
rect 2049 3453 2050 3459
rect 2042 3291 2050 3453
rect 2042 3285 2043 3291
rect 2049 3285 2050 3291
rect 2042 3283 2050 3285
rect 2042 3277 2043 3283
rect 2049 3277 2050 3283
rect 2042 3135 2050 3277
rect 2042 3129 2043 3135
rect 2049 3129 2050 3135
rect 2042 2987 2050 3129
rect 2042 2981 2043 2987
rect 2049 2981 2050 2987
rect 2042 2975 2050 2981
rect 2042 2969 2043 2975
rect 2049 2969 2050 2975
rect 2042 2823 2050 2969
rect 2042 2817 2043 2823
rect 2049 2817 2050 2823
rect 2042 2807 2050 2817
rect 2042 2801 2043 2807
rect 2049 2801 2050 2807
rect 2042 2651 2050 2801
rect 2042 2645 2043 2651
rect 2049 2645 2050 2651
rect 2042 2503 2050 2645
rect 2042 2497 2043 2503
rect 2049 2497 2050 2503
rect 2042 2491 2050 2497
rect 2042 2485 2043 2491
rect 2049 2485 2050 2491
rect 2042 2343 2050 2485
rect 2042 2337 2043 2343
rect 2049 2337 2050 2343
rect 2042 2323 2050 2337
rect 2042 2317 2043 2323
rect 2049 2317 2050 2323
rect 2042 2175 2050 2317
rect 2042 2169 2043 2175
rect 2049 2169 2050 2175
rect 2042 2163 2050 2169
rect 2042 2157 2043 2163
rect 2049 2157 2050 2163
rect 2042 2015 2050 2157
rect 2042 2009 2043 2015
rect 2049 2009 2050 2015
rect 2042 1995 2050 2009
rect 2042 1989 2043 1995
rect 2049 1989 2050 1995
rect 2042 1851 2050 1989
rect 2042 1845 2043 1851
rect 2049 1845 2050 1851
rect 2042 1843 2050 1845
rect 2042 1837 2043 1843
rect 2049 1837 2050 1843
rect 2042 1699 2050 1837
rect 2042 1693 2043 1699
rect 2049 1693 2050 1699
rect 2042 1691 2050 1693
rect 2042 1685 2043 1691
rect 2049 1685 2050 1691
rect 2042 1543 2050 1685
rect 2042 1537 2043 1543
rect 2049 1537 2050 1543
rect 2042 1527 2050 1537
rect 2042 1521 2043 1527
rect 2049 1521 2050 1527
rect 2042 1379 2050 1521
rect 2042 1373 2043 1379
rect 2049 1373 2050 1379
rect 2042 1363 2050 1373
rect 2042 1357 2043 1363
rect 2049 1357 2050 1363
rect 2042 1231 2050 1357
rect 2042 1225 2043 1231
rect 2049 1225 2050 1231
rect 2042 1199 2050 1225
rect 2042 1193 2043 1199
rect 2049 1193 2050 1199
rect 2042 1071 2050 1193
rect 2042 1065 2043 1071
rect 2049 1065 2050 1071
rect 2042 1035 2050 1065
rect 2042 1029 2043 1035
rect 2049 1029 2050 1035
rect 2042 907 2050 1029
rect 2042 901 2043 907
rect 2049 901 2050 907
rect 2042 875 2050 901
rect 2042 869 2043 875
rect 2049 869 2050 875
rect 2042 747 2050 869
rect 2042 741 2043 747
rect 2049 741 2050 747
rect 2042 723 2050 741
rect 2042 717 2043 723
rect 2049 717 2050 723
rect 2042 583 2050 717
rect 2042 577 2043 583
rect 2049 577 2050 583
rect 2042 567 2050 577
rect 2042 561 2043 567
rect 2049 561 2050 567
rect 2042 419 2050 561
rect 2042 413 2043 419
rect 2049 413 2050 419
rect 2042 403 2050 413
rect 2042 397 2043 403
rect 2049 397 2050 403
rect 2042 255 2050 397
rect 2042 249 2043 255
rect 2049 249 2050 255
rect 2042 87 2050 249
rect 2042 81 2043 87
rect 2049 81 2050 87
rect 2042 72 2050 81
rect 2054 3991 2062 4104
rect 2054 3985 2055 3991
rect 2061 3985 2062 3991
rect 2054 3847 2062 3985
rect 2054 3841 2055 3847
rect 2061 3841 2062 3847
rect 2054 3695 2062 3841
rect 2054 3689 2055 3695
rect 2061 3689 2062 3695
rect 2054 3687 2062 3689
rect 2054 3681 2055 3687
rect 2061 3681 2062 3687
rect 2054 3531 2062 3681
rect 2054 3525 2055 3531
rect 2061 3525 2062 3531
rect 2054 3363 2062 3525
rect 2054 3357 2055 3363
rect 2061 3357 2062 3363
rect 2054 3219 2062 3357
rect 2054 3213 2055 3219
rect 2061 3213 2062 3219
rect 2054 3207 2062 3213
rect 2054 3201 2055 3207
rect 2061 3201 2062 3207
rect 2054 3055 2062 3201
rect 2054 3049 2055 3055
rect 2061 3049 2062 3055
rect 2054 2907 2062 3049
rect 2054 2901 2055 2907
rect 2061 2901 2062 2907
rect 2054 2891 2062 2901
rect 2054 2885 2055 2891
rect 2061 2885 2062 2891
rect 2054 2739 2062 2885
rect 2054 2733 2055 2739
rect 2061 2733 2062 2739
rect 2054 2731 2062 2733
rect 2054 2725 2055 2731
rect 2061 2725 2062 2731
rect 2054 2575 2062 2725
rect 2054 2569 2055 2575
rect 2061 2569 2062 2575
rect 2054 2423 2062 2569
rect 2054 2417 2055 2423
rect 2061 2417 2062 2423
rect 2054 2407 2062 2417
rect 2054 2401 2055 2407
rect 2061 2401 2062 2407
rect 2054 2259 2062 2401
rect 2054 2253 2055 2259
rect 2061 2253 2062 2259
rect 2054 2243 2062 2253
rect 2054 2237 2055 2243
rect 2061 2237 2062 2243
rect 2054 2095 2062 2237
rect 2054 2089 2055 2095
rect 2061 2089 2062 2095
rect 2054 2079 2062 2089
rect 2054 2073 2055 2079
rect 2061 2073 2062 2079
rect 2054 1931 2062 2073
rect 2054 1925 2055 1931
rect 2061 1925 2062 1931
rect 2054 1915 2062 1925
rect 2054 1909 2055 1915
rect 2061 1909 2062 1915
rect 2054 1771 2062 1909
rect 2054 1765 2055 1771
rect 2061 1765 2062 1771
rect 2054 1623 2062 1765
rect 2054 1617 2055 1623
rect 2061 1617 2062 1623
rect 2054 1607 2062 1617
rect 2054 1601 2055 1607
rect 2061 1601 2062 1607
rect 2054 1459 2062 1601
rect 2054 1453 2055 1459
rect 2061 1453 2062 1459
rect 2054 1443 2062 1453
rect 2054 1437 2055 1443
rect 2061 1437 2062 1443
rect 2054 1303 2062 1437
rect 2054 1297 2055 1303
rect 2061 1297 2062 1303
rect 2054 1283 2062 1297
rect 2054 1277 2055 1283
rect 2061 1277 2062 1283
rect 2054 1151 2062 1277
rect 2054 1145 2055 1151
rect 2061 1145 2062 1151
rect 2054 1123 2062 1145
rect 2054 1117 2055 1123
rect 2061 1117 2062 1123
rect 2054 987 2062 1117
rect 2054 981 2055 987
rect 2061 981 2062 987
rect 2054 959 2062 981
rect 2054 953 2055 959
rect 2061 953 2062 959
rect 2054 823 2062 953
rect 2054 817 2055 823
rect 2061 817 2062 823
rect 2054 803 2062 817
rect 2054 797 2055 803
rect 2061 797 2062 803
rect 2054 663 2062 797
rect 2054 657 2055 663
rect 2061 657 2062 663
rect 2054 647 2062 657
rect 2054 641 2055 647
rect 2061 641 2062 647
rect 2054 495 2062 641
rect 2054 489 2055 495
rect 2061 489 2062 495
rect 2054 487 2062 489
rect 2054 481 2055 487
rect 2061 481 2062 487
rect 2054 335 2062 481
rect 2054 329 2055 335
rect 2061 329 2062 335
rect 2054 159 2062 329
rect 2054 153 2055 159
rect 2061 153 2062 159
rect 2054 72 2062 153
rect 4014 3779 4022 4104
rect 4014 3773 4015 3779
rect 4021 3773 4022 3779
rect 4014 3291 4022 3773
rect 4014 3285 4015 3291
rect 4021 3285 4022 3291
rect 4014 2987 4022 3285
rect 4014 2981 4015 2987
rect 4021 2981 4022 2987
rect 4014 2823 4022 2981
rect 4014 2817 4015 2823
rect 4021 2817 4022 2823
rect 4014 2491 4022 2817
rect 4014 2485 4015 2491
rect 4021 2485 4022 2491
rect 4014 2323 4022 2485
rect 4014 2317 4015 2323
rect 4021 2317 4022 2323
rect 4014 2163 4022 2317
rect 4014 2157 4015 2163
rect 4021 2157 4022 2163
rect 4014 1995 4022 2157
rect 4014 1989 4015 1995
rect 4021 1989 4022 1995
rect 4014 1843 4022 1989
rect 4014 1837 4015 1843
rect 4021 1837 4022 1843
rect 4014 1691 4022 1837
rect 4014 1685 4015 1691
rect 4021 1685 4022 1691
rect 4014 1527 4022 1685
rect 4014 1521 4015 1527
rect 4021 1521 4022 1527
rect 4014 1363 4022 1521
rect 4014 1357 4015 1363
rect 4021 1357 4022 1363
rect 4014 1199 4022 1357
rect 4014 1193 4015 1199
rect 4021 1193 4022 1199
rect 4014 1035 4022 1193
rect 4014 1029 4015 1035
rect 4021 1029 4022 1035
rect 4014 875 4022 1029
rect 4014 869 4015 875
rect 4021 869 4022 875
rect 4014 723 4022 869
rect 4014 717 4015 723
rect 4021 717 4022 723
rect 4014 567 4022 717
rect 4014 561 4015 567
rect 4021 561 4022 567
rect 4014 403 4022 561
rect 4014 397 4015 403
rect 4021 397 4022 403
rect 4014 72 4022 397
rect 4026 3695 4034 4104
rect 4026 3689 4027 3695
rect 4033 3689 4034 3695
rect 4026 3219 4034 3689
rect 4026 3213 4027 3219
rect 4033 3213 4034 3219
rect 4026 2907 4034 3213
rect 4026 2901 4027 2907
rect 4033 2901 4034 2907
rect 4026 2739 4034 2901
rect 4026 2733 4027 2739
rect 4033 2733 4034 2739
rect 4026 2407 4034 2733
rect 4026 2401 4027 2407
rect 4033 2401 4034 2407
rect 4026 2243 4034 2401
rect 4026 2237 4027 2243
rect 4033 2237 4034 2243
rect 4026 2079 4034 2237
rect 4026 2073 4027 2079
rect 4033 2073 4034 2079
rect 4026 1915 4034 2073
rect 4026 1909 4027 1915
rect 4033 1909 4034 1915
rect 4026 1607 4034 1909
rect 4026 1601 4027 1607
rect 4033 1601 4034 1607
rect 4026 1443 4034 1601
rect 4026 1437 4027 1443
rect 4033 1437 4034 1443
rect 4026 1283 4034 1437
rect 4026 1277 4027 1283
rect 4033 1277 4034 1283
rect 4026 1123 4034 1277
rect 4026 1117 4027 1123
rect 4033 1117 4034 1123
rect 4026 959 4034 1117
rect 4026 953 4027 959
rect 4033 953 4034 959
rect 4026 803 4034 953
rect 4026 797 4027 803
rect 4033 797 4034 803
rect 4026 647 4034 797
rect 4026 641 4027 647
rect 4033 641 4034 647
rect 4026 487 4034 641
rect 4026 481 4027 487
rect 4033 481 4034 487
rect 4026 72 4034 481
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__199
timestamp 1731220555
transform 1 0 3984 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220555
transform 1 0 2064 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220555
transform 1 0 3984 0 1 3936
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220555
transform 1 0 2064 0 1 3936
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220555
transform 1 0 3984 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220555
transform 1 0 2064 0 -1 3904
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220555
transform 1 0 3984 0 1 3792
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220555
transform 1 0 2064 0 1 3792
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220555
transform 1 0 3984 0 -1 3760
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220555
transform 1 0 2064 0 -1 3760
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220555
transform 1 0 3984 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220555
transform 1 0 2064 0 1 3636
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220555
transform 1 0 3984 0 -1 3592
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220555
transform 1 0 2064 0 -1 3592
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220555
transform 1 0 3984 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220555
transform 1 0 2064 0 1 3476
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220555
transform 1 0 3984 0 -1 3444
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220555
transform 1 0 2064 0 -1 3444
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220555
transform 1 0 3984 0 1 3304
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220555
transform 1 0 2064 0 1 3304
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220555
transform 1 0 3984 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220555
transform 1 0 2064 0 -1 3272
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220555
transform 1 0 3984 0 1 3160
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220555
transform 1 0 2064 0 1 3160
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220555
transform 1 0 3984 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220555
transform 1 0 2064 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220555
transform 1 0 3984 0 1 3000
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220555
transform 1 0 2064 0 1 3000
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220555
transform 1 0 3984 0 -1 2968
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220555
transform 1 0 2064 0 -1 2968
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220555
transform 1 0 3984 0 1 2848
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220555
transform 1 0 2064 0 1 2848
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220555
transform 1 0 3984 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220555
transform 1 0 2064 0 -1 2804
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220555
transform 1 0 3984 0 1 2680
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220555
transform 1 0 2064 0 1 2680
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220555
transform 1 0 3984 0 -1 2636
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220555
transform 1 0 2064 0 -1 2636
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220555
transform 1 0 3984 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220555
transform 1 0 2064 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220555
transform 1 0 3984 0 -1 2472
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220555
transform 1 0 2064 0 -1 2472
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220555
transform 1 0 3984 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220555
transform 1 0 2064 0 1 2348
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220555
transform 1 0 3984 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220555
transform 1 0 2064 0 -1 2304
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220555
transform 1 0 3984 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220555
transform 1 0 2064 0 1 2184
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220555
transform 1 0 3984 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220555
transform 1 0 2064 0 -1 2144
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220555
transform 1 0 3984 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220555
transform 1 0 2064 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220555
transform 1 0 3984 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220555
transform 1 0 2064 0 -1 1976
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220555
transform 1 0 3984 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220555
transform 1 0 2064 0 1 1856
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220555
transform 1 0 3984 0 -1 1824
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220555
transform 1 0 2064 0 -1 1824
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220555
transform 1 0 3984 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220555
transform 1 0 2064 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220555
transform 1 0 3984 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220555
transform 1 0 2064 0 -1 1672
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220555
transform 1 0 3984 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220555
transform 1 0 2064 0 1 1548
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220555
transform 1 0 3984 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220555
transform 1 0 2064 0 -1 1508
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220555
transform 1 0 3984 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220555
transform 1 0 2064 0 1 1384
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220555
transform 1 0 3984 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220555
transform 1 0 2064 0 -1 1344
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220555
transform 1 0 3984 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220555
transform 1 0 2064 0 1 1224
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220555
transform 1 0 3984 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220555
transform 1 0 2064 0 -1 1180
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220555
transform 1 0 3984 0 1 1064
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220555
transform 1 0 2064 0 1 1064
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220555
transform 1 0 3984 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220555
transform 1 0 2064 0 -1 1016
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220555
transform 1 0 3984 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220555
transform 1 0 2064 0 1 900
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220555
transform 1 0 3984 0 -1 856
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220555
transform 1 0 2064 0 -1 856
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220555
transform 1 0 3984 0 1 744
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220555
transform 1 0 2064 0 1 744
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220555
transform 1 0 3984 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220555
transform 1 0 2064 0 -1 704
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220555
transform 1 0 3984 0 1 588
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220555
transform 1 0 2064 0 1 588
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220555
transform 1 0 3984 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220555
transform 1 0 2064 0 -1 548
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220555
transform 1 0 3984 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220555
transform 1 0 2064 0 1 428
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220555
transform 1 0 3984 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220555
transform 1 0 2064 0 -1 384
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220555
transform 1 0 3984 0 1 272
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220555
transform 1 0 2064 0 1 272
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220555
transform 1 0 3984 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220555
transform 1 0 2064 0 -1 240
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220555
transform 1 0 3984 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220555
transform 1 0 2064 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220555
transform 1 0 2024 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220555
transform 1 0 104 0 -1 4048
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220555
transform 1 0 2024 0 1 3932
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220555
transform 1 0 104 0 1 3932
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220555
transform 1 0 2024 0 -1 3900
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220555
transform 1 0 104 0 -1 3900
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220555
transform 1 0 2024 0 1 3788
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220555
transform 1 0 104 0 1 3788
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220555
transform 1 0 2024 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220555
transform 1 0 104 0 -1 3744
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220555
transform 1 0 2024 0 1 3628
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220555
transform 1 0 104 0 1 3628
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220555
transform 1 0 2024 0 -1 3596
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220555
transform 1 0 104 0 -1 3596
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220555
transform 1 0 2024 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220555
transform 1 0 104 0 1 3472
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220555
transform 1 0 2024 0 -1 3440
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220555
transform 1 0 104 0 -1 3440
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220555
transform 1 0 2024 0 1 3304
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220555
transform 1 0 104 0 1 3304
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220555
transform 1 0 2024 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220555
transform 1 0 104 0 -1 3264
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220555
transform 1 0 2024 0 1 3148
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220555
transform 1 0 104 0 1 3148
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220555
transform 1 0 2024 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220555
transform 1 0 104 0 -1 3116
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220555
transform 1 0 2024 0 1 2996
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220555
transform 1 0 104 0 1 2996
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220555
transform 1 0 2024 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220555
transform 1 0 104 0 -1 2956
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220555
transform 1 0 2024 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220555
transform 1 0 104 0 1 2832
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220555
transform 1 0 2024 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220555
transform 1 0 104 0 -1 2788
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220555
transform 1 0 2024 0 1 2672
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220555
transform 1 0 104 0 1 2672
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220555
transform 1 0 2024 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220555
transform 1 0 104 0 -1 2632
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220555
transform 1 0 2024 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220555
transform 1 0 104 0 1 2516
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220555
transform 1 0 2024 0 -1 2484
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220555
transform 1 0 104 0 -1 2484
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220555
transform 1 0 2024 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220555
transform 1 0 104 0 1 2364
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220555
transform 1 0 2024 0 -1 2324
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220555
transform 1 0 104 0 -1 2324
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220555
transform 1 0 2024 0 1 2200
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220555
transform 1 0 104 0 1 2200
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220555
transform 1 0 2024 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220555
transform 1 0 104 0 -1 2156
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220555
transform 1 0 2024 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220555
transform 1 0 104 0 1 2036
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220555
transform 1 0 2024 0 -1 1996
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220555
transform 1 0 104 0 -1 1996
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220555
transform 1 0 2024 0 1 1872
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220555
transform 1 0 104 0 1 1872
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220555
transform 1 0 2024 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220555
transform 1 0 104 0 -1 1832
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220555
transform 1 0 2024 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220555
transform 1 0 104 0 1 1712
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220555
transform 1 0 2024 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220555
transform 1 0 104 0 -1 1680
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220555
transform 1 0 2024 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220555
transform 1 0 104 0 1 1564
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220555
transform 1 0 2024 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220555
transform 1 0 104 0 -1 1524
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220555
transform 1 0 2024 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220555
transform 1 0 104 0 1 1400
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220555
transform 1 0 2024 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220555
transform 1 0 104 0 -1 1360
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220555
transform 1 0 2024 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220555
transform 1 0 104 0 1 1244
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220555
transform 1 0 2024 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220555
transform 1 0 104 0 -1 1212
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220555
transform 1 0 2024 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220555
transform 1 0 104 0 1 1092
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220555
transform 1 0 2024 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220555
transform 1 0 104 0 -1 1052
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220555
transform 1 0 2024 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220555
transform 1 0 104 0 1 928
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220555
transform 1 0 2024 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220555
transform 1 0 104 0 -1 888
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220555
transform 1 0 2024 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220555
transform 1 0 104 0 1 764
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220555
transform 1 0 2024 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220555
transform 1 0 104 0 -1 728
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220555
transform 1 0 2024 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220555
transform 1 0 104 0 1 604
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220555
transform 1 0 2024 0 -1 564
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220555
transform 1 0 104 0 -1 564
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220555
transform 1 0 2024 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220555
transform 1 0 104 0 1 436
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220555
transform 1 0 2024 0 -1 400
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220555
transform 1 0 104 0 -1 400
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220555
transform 1 0 2024 0 1 276
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220555
transform 1 0 104 0 1 276
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220555
transform 1 0 2024 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220555
transform 1 0 104 0 -1 236
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220555
transform 1 0 2024 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220555
transform 1 0 104 0 1 100
box 7 3 12 24
use _0_0std_0_0cells_0_0LATCH  tst_5999_6
timestamp 1731220555
transform 1 0 128 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5998_6
timestamp 1731220555
transform 1 0 232 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5997_6
timestamp 1731220555
transform 1 0 336 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5996_6
timestamp 1731220555
transform 1 0 448 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5995_6
timestamp 1731220555
transform 1 0 584 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5994_6
timestamp 1731220555
transform 1 0 720 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5993_6
timestamp 1731220555
transform 1 0 856 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5992_6
timestamp 1731220555
transform 1 0 128 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5991_6
timestamp 1731220555
transform 1 0 256 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5990_6
timestamp 1731220555
transform 1 0 408 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5989_6
timestamp 1731220555
transform 1 0 576 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5988_6
timestamp 1731220555
transform 1 0 760 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5987_6
timestamp 1731220555
transform 1 0 312 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5986_6
timestamp 1731220555
transform 1 0 440 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5985_6
timestamp 1731220555
transform 1 0 584 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5984_6
timestamp 1731220555
transform 1 0 744 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5983_6
timestamp 1731220555
transform 1 0 744 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5982_6
timestamp 1731220555
transform 1 0 608 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5981_6
timestamp 1731220555
transform 1 0 472 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5980_6
timestamp 1731220555
transform 1 0 512 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5979_6
timestamp 1731220555
transform 1 0 616 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5978_6
timestamp 1731220555
transform 1 0 720 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5977_6
timestamp 1731220555
transform 1 0 640 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5976_6
timestamp 1731220555
transform 1 0 824 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5975_6
timestamp 1731220555
transform 1 0 944 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5974_6
timestamp 1731220555
transform 1 0 1024 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5973_6
timestamp 1731220555
transform 1 0 888 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5972_6
timestamp 1731220555
transform 1 0 920 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5971_6
timestamp 1731220555
transform 1 0 1104 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5970_6
timestamp 1731220555
transform 1 0 1288 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5969_6
timestamp 1731220555
transform 1 0 1352 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5968_6
timestamp 1731220555
transform 1 0 1152 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5967_6
timestamp 1731220555
transform 1 0 952 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5966_6
timestamp 1731220555
transform 1 0 992 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5965_6
timestamp 1731220555
transform 1 0 1128 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5964_6
timestamp 1731220555
transform 1 0 1256 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5963_6
timestamp 1731220555
transform 1 0 1376 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5962_6
timestamp 1731220555
transform 1 0 1496 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5961_6
timestamp 1731220555
transform 1 0 1624 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5960_6
timestamp 1731220555
transform 1 0 1752 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5959_6
timestamp 1731220555
transform 1 0 1560 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5958_6
timestamp 1731220555
transform 1 0 1776 0 -1 252
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5957_6
timestamp 1731220555
transform 1 0 1880 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5956_6
timestamp 1731220555
transform 1 0 1480 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5955_6
timestamp 1731220555
transform 1 0 1680 0 1 260
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5954_6
timestamp 1731220555
transform 1 0 1680 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5953_6
timestamp 1731220555
transform 1 0 1552 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5952_6
timestamp 1731220555
transform 1 0 1424 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5951_6
timestamp 1731220555
transform 1 0 1160 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5950_6
timestamp 1731220555
transform 1 0 1296 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5949_6
timestamp 1731220555
transform 1 0 1392 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5948_6
timestamp 1731220555
transform 1 0 1568 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5947_6
timestamp 1731220555
transform 1 0 1080 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5946_6
timestamp 1731220555
transform 1 0 1232 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5945_6
timestamp 1731220555
transform 1 0 1280 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5944_6
timestamp 1731220555
transform 1 0 1136 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5943_6
timestamp 1731220555
transform 1 0 1000 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5942_6
timestamp 1731220555
transform 1 0 752 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5941_6
timestamp 1731220555
transform 1 0 872 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5940_6
timestamp 1731220555
transform 1 0 896 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5939_6
timestamp 1731220555
transform 1 0 1008 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5938_6
timestamp 1731220555
transform 1 0 568 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5937_6
timestamp 1731220555
transform 1 0 672 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5936_6
timestamp 1731220555
transform 1 0 784 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5935_6
timestamp 1731220555
transform 1 0 856 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5934_6
timestamp 1731220555
transform 1 0 736 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5933_6
timestamp 1731220555
transform 1 0 616 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5932_6
timestamp 1731220555
transform 1 0 504 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5931_6
timestamp 1731220555
transform 1 0 400 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5930_6
timestamp 1731220555
transform 1 0 240 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5929_6
timestamp 1731220555
transform 1 0 344 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5928_6
timestamp 1731220555
transform 1 0 456 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5927_6
timestamp 1731220555
transform 1 0 568 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5926_6
timestamp 1731220555
transform 1 0 688 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5925_6
timestamp 1731220555
transform 1 0 704 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5924_6
timestamp 1731220555
transform 1 0 912 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5923_6
timestamp 1731220555
transform 1 0 128 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5922_6
timestamp 1731220555
transform 1 0 296 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5921_6
timestamp 1731220555
transform 1 0 496 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5920_6
timestamp 1731220555
transform 1 0 648 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5919_6
timestamp 1731220555
transform 1 0 848 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5918_6
timestamp 1731220555
transform 1 0 448 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5917_6
timestamp 1731220555
transform 1 0 264 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5916_6
timestamp 1731220555
transform 1 0 128 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5915_6
timestamp 1731220555
transform 1 0 128 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5914_6
timestamp 1731220555
transform 1 0 256 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5913_6
timestamp 1731220555
transform 1 0 424 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5912_6
timestamp 1731220555
transform 1 0 600 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5911_6
timestamp 1731220555
transform 1 0 776 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5910_6
timestamp 1731220555
transform 1 0 128 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5909_6
timestamp 1731220555
transform 1 0 280 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5908_6
timestamp 1731220555
transform 1 0 472 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5907_6
timestamp 1731220555
transform 1 0 680 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5906_6
timestamp 1731220555
transform 1 0 888 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5905_6
timestamp 1731220555
transform 1 0 160 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5904_6
timestamp 1731220555
transform 1 0 328 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5903_6
timestamp 1731220555
transform 1 0 512 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5902_6
timestamp 1731220555
transform 1 0 704 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5901_6
timestamp 1731220555
transform 1 0 896 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5900_6
timestamp 1731220555
transform 1 0 320 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5899_6
timestamp 1731220555
transform 1 0 440 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5898_6
timestamp 1731220555
transform 1 0 576 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5897_6
timestamp 1731220555
transform 1 0 720 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5896_6
timestamp 1731220555
transform 1 0 880 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5895_6
timestamp 1731220555
transform 1 0 528 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5894_6
timestamp 1731220555
transform 1 0 632 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5893_6
timestamp 1731220555
transform 1 0 736 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5892_6
timestamp 1731220555
transform 1 0 840 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5891_6
timestamp 1731220555
transform 1 0 952 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5890_6
timestamp 1731220555
transform 1 0 768 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5889_6
timestamp 1731220555
transform 1 0 560 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5888_6
timestamp 1731220555
transform 1 0 664 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5887_6
timestamp 1731220555
transform 1 0 712 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5886_6
timestamp 1731220555
transform 1 0 592 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5885_6
timestamp 1731220555
transform 1 0 480 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5884_6
timestamp 1731220555
transform 1 0 376 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5883_6
timestamp 1731220555
transform 1 0 552 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5882_6
timestamp 1731220555
transform 1 0 728 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5881_6
timestamp 1731220555
transform 1 0 744 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5880_6
timestamp 1731220555
transform 1 0 512 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5879_6
timestamp 1731220555
transform 1 0 280 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5878_6
timestamp 1731220555
transform 1 0 184 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5877_6
timestamp 1731220555
transform 1 0 360 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5876_6
timestamp 1731220555
transform 1 0 544 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5875_6
timestamp 1731220555
transform 1 0 424 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5874_6
timestamp 1731220555
transform 1 0 264 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5873_6
timestamp 1731220555
transform 1 0 128 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5872_6
timestamp 1731220555
transform 1 0 128 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5871_6
timestamp 1731220555
transform 1 0 248 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5870_6
timestamp 1731220555
transform 1 0 384 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5869_6
timestamp 1731220555
transform 1 0 464 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5868_6
timestamp 1731220555
transform 1 0 280 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5867_6
timestamp 1731220555
transform 1 0 128 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5866_6
timestamp 1731220555
transform 1 0 128 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5865_6
timestamp 1731220555
transform 1 0 280 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5864_6
timestamp 1731220555
transform 1 0 456 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5863_6
timestamp 1731220555
transform 1 0 488 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5862_6
timestamp 1731220555
transform 1 0 296 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5861_6
timestamp 1731220555
transform 1 0 128 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5860_6
timestamp 1731220555
transform 1 0 216 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5859_6
timestamp 1731220555
transform 1 0 368 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5858_6
timestamp 1731220555
transform 1 0 528 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5857_6
timestamp 1731220555
transform 1 0 336 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5856_6
timestamp 1731220555
transform 1 0 472 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5855_6
timestamp 1731220555
transform 1 0 760 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5854_6
timestamp 1731220555
transform 1 0 920 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5853_6
timestamp 1731220555
transform 1 0 912 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5852_6
timestamp 1731220555
transform 1 0 760 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5851_6
timestamp 1731220555
transform 1 0 616 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5850_6
timestamp 1731220555
transform 1 0 688 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5849_6
timestamp 1731220555
transform 1 0 848 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5848_6
timestamp 1731220555
transform 1 0 872 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5847_6
timestamp 1731220555
transform 1 0 680 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5846_6
timestamp 1731220555
transform 1 0 640 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5845_6
timestamp 1731220555
transform 1 0 824 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5844_6
timestamp 1731220555
transform 1 0 872 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5843_6
timestamp 1731220555
transform 1 0 664 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5842_6
timestamp 1731220555
transform 1 0 656 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5841_6
timestamp 1731220555
transform 1 0 520 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5840_6
timestamp 1731220555
transform 1 0 576 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5839_6
timestamp 1731220555
transform 1 0 728 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5838_6
timestamp 1731220555
transform 1 0 728 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5837_6
timestamp 1731220555
transform 1 0 912 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5836_6
timestamp 1731220555
transform 1 0 960 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5835_6
timestamp 1731220555
transform 1 0 1088 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5834_6
timestamp 1731220555
transform 1 0 912 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5833_6
timestamp 1731220555
transform 1 0 944 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5832_6
timestamp 1731220555
transform 1 0 832 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5831_6
timestamp 1731220555
transform 1 0 872 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5830_6
timestamp 1731220555
transform 1 0 976 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5829_6
timestamp 1731220555
transform 1 0 1080 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5828_6
timestamp 1731220555
transform 1 0 1064 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5827_6
timestamp 1731220555
transform 1 0 1176 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5826_6
timestamp 1731220555
transform 1 0 1208 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5825_6
timestamp 1731220555
transform 1 0 1040 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5824_6
timestamp 1731220555
transform 1 0 1080 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5823_6
timestamp 1731220555
transform 1 0 1096 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5822_6
timestamp 1731220555
transform 1 0 944 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5821_6
timestamp 1731220555
transform 1 0 1056 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5820_6
timestamp 1731220555
transform 1 0 832 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5819_6
timestamp 1731220555
transform 1 0 1008 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5818_6
timestamp 1731220555
transform 1 0 1216 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5817_6
timestamp 1731220555
transform 1 0 1448 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5816_6
timestamp 1731220555
transform 1 0 1688 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5815_6
timestamp 1731220555
transform 1 0 984 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5814_6
timestamp 1731220555
transform 1 0 1120 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5813_6
timestamp 1731220555
transform 1 0 1264 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5812_6
timestamp 1731220555
transform 1 0 1424 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5811_6
timestamp 1731220555
transform 1 0 1592 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5810_6
timestamp 1731220555
transform 1 0 1120 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5809_6
timestamp 1731220555
transform 1 0 1240 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5808_6
timestamp 1731220555
transform 1 0 1360 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5807_6
timestamp 1731220555
transform 1 0 1480 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5806_6
timestamp 1731220555
transform 1 0 1600 0 1 588
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5805_6
timestamp 1731220555
transform 1 0 1424 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5804_6
timestamp 1731220555
transform 1 0 1568 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5803_6
timestamp 1731220555
transform 1 0 1712 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5802_6
timestamp 1731220555
transform 1 0 1856 0 -1 580
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5801_6
timestamp 1731220555
transform 1 0 1912 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5800_6
timestamp 1731220555
transform 1 0 1752 0 1 420
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5799_6
timestamp 1731220555
transform 1 0 1808 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5798_6
timestamp 1731220555
transform 1 0 1912 0 -1 416
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5797_6
timestamp 1731220555
transform 1 0 2088 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5796_6
timestamp 1731220555
transform 1 0 2248 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5795_6
timestamp 1731220555
transform 1 0 2448 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5794_6
timestamp 1731220555
transform 1 0 2248 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5793_6
timestamp 1731220555
transform 1 0 2088 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5792_6
timestamp 1731220555
transform 1 0 2088 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5791_6
timestamp 1731220555
transform 1 0 2192 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5790_6
timestamp 1731220555
transform 1 0 2296 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5789_6
timestamp 1731220555
transform 1 0 2400 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5788_6
timestamp 1731220555
transform 1 0 2504 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5787_6
timestamp 1731220555
transform 1 0 2632 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5786_6
timestamp 1731220555
transform 1 0 2752 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5785_6
timestamp 1731220555
transform 1 0 2880 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5784_6
timestamp 1731220555
transform 1 0 2664 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5783_6
timestamp 1731220555
transform 1 0 2608 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5782_6
timestamp 1731220555
transform 1 0 2432 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5781_6
timestamp 1731220555
transform 1 0 2568 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5780_6
timestamp 1731220555
transform 1 0 2672 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5779_6
timestamp 1731220555
transform 1 0 2792 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5778_6
timestamp 1731220555
transform 1 0 2840 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5777_6
timestamp 1731220555
transform 1 0 2488 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5776_6
timestamp 1731220555
transform 1 0 2592 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5775_6
timestamp 1731220555
transform 1 0 2712 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5774_6
timestamp 1731220555
transform 1 0 2712 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5773_6
timestamp 1731220555
transform 1 0 2568 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5772_6
timestamp 1731220555
transform 1 0 2280 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5771_6
timestamp 1731220555
transform 1 0 2424 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5770_6
timestamp 1731220555
transform 1 0 2432 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5769_6
timestamp 1731220555
transform 1 0 2272 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5768_6
timestamp 1731220555
transform 1 0 2104 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5767_6
timestamp 1731220555
transform 1 0 2088 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5766_6
timestamp 1731220555
transform 1 0 1912 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5765_6
timestamp 1731220555
transform 1 0 1760 0 -1 744
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5764_6
timestamp 1731220555
transform 1 0 1912 0 1 748
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5763_6
timestamp 1731220555
transform 1 0 2088 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5762_6
timestamp 1731220555
transform 1 0 2088 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5761_6
timestamp 1731220555
transform 1 0 2216 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5760_6
timestamp 1731220555
transform 1 0 2128 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5759_6
timestamp 1731220555
transform 1 0 2264 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5758_6
timestamp 1731220555
transform 1 0 2408 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5757_6
timestamp 1731220555
transform 1 0 2296 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5756_6
timestamp 1731220555
transform 1 0 2464 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5755_6
timestamp 1731220555
transform 1 0 2640 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5754_6
timestamp 1731220555
transform 1 0 2568 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5753_6
timestamp 1731220555
transform 1 0 2736 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5752_6
timestamp 1731220555
transform 1 0 2728 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5751_6
timestamp 1731220555
transform 1 0 2552 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5750_6
timestamp 1731220555
transform 1 0 2384 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5749_6
timestamp 1731220555
transform 1 0 2368 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5748_6
timestamp 1731220555
transform 1 0 2304 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5747_6
timestamp 1731220555
transform 1 0 2528 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5746_6
timestamp 1731220555
transform 1 0 2752 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5745_6
timestamp 1731220555
transform 1 0 2592 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5744_6
timestamp 1731220555
transform 1 0 2760 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5743_6
timestamp 1731220555
transform 1 0 2856 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5742_6
timestamp 1731220555
transform 1 0 2984 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5741_6
timestamp 1731220555
transform 1 0 3136 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5740_6
timestamp 1731220555
transform 1 0 3296 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5739_6
timestamp 1731220555
transform 1 0 2936 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5738_6
timestamp 1731220555
transform 1 0 3096 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5737_6
timestamp 1731220555
transform 1 0 3280 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5736_6
timestamp 1731220555
transform 1 0 3480 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5735_6
timestamp 1731220555
transform 1 0 2784 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5734_6
timestamp 1731220555
transform 1 0 2976 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5733_6
timestamp 1731220555
transform 1 0 3192 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5732_6
timestamp 1731220555
transform 1 0 3416 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5731_6
timestamp 1731220555
transform 1 0 3656 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5730_6
timestamp 1731220555
transform 1 0 3088 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5729_6
timestamp 1731220555
transform 1 0 2872 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5728_6
timestamp 1731220555
transform 1 0 2992 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5727_6
timestamp 1731220555
transform 1 0 3112 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5726_6
timestamp 1731220555
transform 1 0 3224 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5725_6
timestamp 1731220555
transform 1 0 3336 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5724_6
timestamp 1731220555
transform 1 0 3448 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5723_6
timestamp 1731220555
transform 1 0 3560 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5722_6
timestamp 1731220555
transform 1 0 3664 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5721_6
timestamp 1731220555
transform 1 0 3296 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5720_6
timestamp 1731220555
transform 1 0 3496 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5719_6
timestamp 1731220555
transform 1 0 3696 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5718_6
timestamp 1731220555
transform 1 0 3768 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5717_6
timestamp 1731220555
transform 1 0 3872 0 1 84
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5716_6
timestamp 1731220555
transform 1 0 3872 0 -1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5715_6
timestamp 1731220555
transform 1 0 3872 0 1 256
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5714_6
timestamp 1731220555
transform 1 0 3872 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5713_6
timestamp 1731220555
transform 1 0 3800 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5712_6
timestamp 1731220555
transform 1 0 3688 0 -1 400
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5711_6
timestamp 1731220555
transform 1 0 3456 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5710_6
timestamp 1731220555
transform 1 0 3624 0 1 412
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5709_6
timestamp 1731220555
transform 1 0 3632 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5708_6
timestamp 1731220555
transform 1 0 3472 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5707_6
timestamp 1731220555
transform 1 0 3008 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5706_6
timestamp 1731220555
transform 1 0 3160 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5705_6
timestamp 1731220555
transform 1 0 3312 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5704_6
timestamp 1731220555
transform 1 0 3464 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5703_6
timestamp 1731220555
transform 1 0 3280 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5702_6
timestamp 1731220555
transform 1 0 2928 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5701_6
timestamp 1731220555
transform 1 0 3104 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5700_6
timestamp 1731220555
transform 1 0 3184 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5699_6
timestamp 1731220555
transform 1 0 2968 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5698_6
timestamp 1731220555
transform 1 0 2928 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5697_6
timestamp 1731220555
transform 1 0 2656 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5696_6
timestamp 1731220555
transform 1 0 2912 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5695_6
timestamp 1731220555
transform 1 0 3096 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5694_6
timestamp 1731220555
transform 1 0 2912 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5693_6
timestamp 1731220555
transform 1 0 3016 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5692_6
timestamp 1731220555
transform 1 0 2824 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5691_6
timestamp 1731220555
transform 1 0 2680 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5690_6
timestamp 1731220555
transform 1 0 2536 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5689_6
timestamp 1731220555
transform 1 0 2680 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5688_6
timestamp 1731220555
transform 1 0 2856 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5687_6
timestamp 1731220555
transform 1 0 2832 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5686_6
timestamp 1731220555
transform 1 0 2672 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5685_6
timestamp 1731220555
transform 1 0 2672 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5684_6
timestamp 1731220555
transform 1 0 2816 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5683_6
timestamp 1731220555
transform 1 0 2792 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5682_6
timestamp 1731220555
transform 1 0 2624 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5681_6
timestamp 1731220555
transform 1 0 2496 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5680_6
timestamp 1731220555
transform 1 0 2632 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5679_6
timestamp 1731220555
transform 1 0 2688 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5678_6
timestamp 1731220555
transform 1 0 2360 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5677_6
timestamp 1731220555
transform 1 0 2384 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5676_6
timestamp 1731220555
transform 1 0 2632 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5675_6
timestamp 1731220555
transform 1 0 2440 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5674_6
timestamp 1731220555
transform 1 0 2256 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5673_6
timestamp 1731220555
transform 1 0 2368 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5672_6
timestamp 1731220555
transform 1 0 2184 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5671_6
timestamp 1731220555
transform 1 0 2120 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5670_6
timestamp 1731220555
transform 1 0 2296 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5669_6
timestamp 1731220555
transform 1 0 2256 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5668_6
timestamp 1731220555
transform 1 0 2088 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5667_6
timestamp 1731220555
transform 1 0 2200 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5666_6
timestamp 1731220555
transform 1 0 2088 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5665_6
timestamp 1731220555
transform 1 0 1912 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5664_6
timestamp 1731220555
transform 1 0 1912 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5663_6
timestamp 1731220555
transform 1 0 1792 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5662_6
timestamp 1731220555
transform 1 0 1912 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5661_6
timestamp 1731220555
transform 1 0 1912 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5660_6
timestamp 1731220555
transform 1 0 2088 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5659_6
timestamp 1731220555
transform 1 0 2088 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5658_6
timestamp 1731220555
transform 1 0 2240 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5657_6
timestamp 1731220555
transform 1 0 2256 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5656_6
timestamp 1731220555
transform 1 0 2088 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5655_6
timestamp 1731220555
transform 1 0 2120 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5654_6
timestamp 1731220555
transform 1 0 2296 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5653_6
timestamp 1731220555
transform 1 0 2088 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5652_6
timestamp 1731220555
transform 1 0 2256 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5651_6
timestamp 1731220555
transform 1 0 2584 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5650_6
timestamp 1731220555
transform 1 0 2824 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5649_6
timestamp 1731220555
transform 1 0 2832 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5648_6
timestamp 1731220555
transform 1 0 2632 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5647_6
timestamp 1731220555
transform 1 0 2560 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5646_6
timestamp 1731220555
transform 1 0 2320 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5645_6
timestamp 1731220555
transform 1 0 2376 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5644_6
timestamp 1731220555
transform 1 0 2528 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5643_6
timestamp 1731220555
transform 1 0 2672 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5642_6
timestamp 1731220555
transform 1 0 2504 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5641_6
timestamp 1731220555
transform 1 0 2520 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5640_6
timestamp 1731220555
transform 1 0 2416 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5639_6
timestamp 1731220555
transform 1 0 2440 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5638_6
timestamp 1731220555
transform 1 0 2336 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5637_6
timestamp 1731220555
transform 1 0 2416 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5636_6
timestamp 1731220555
transform 1 0 2552 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5635_6
timestamp 1731220555
transform 1 0 2560 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5634_6
timestamp 1731220555
transform 1 0 2336 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5633_6
timestamp 1731220555
transform 1 0 2416 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5632_6
timestamp 1731220555
transform 1 0 2600 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5631_6
timestamp 1731220555
transform 1 0 2792 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5630_6
timestamp 1731220555
transform 1 0 2752 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5629_6
timestamp 1731220555
transform 1 0 2536 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5628_6
timestamp 1731220555
transform 1 0 2464 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5627_6
timestamp 1731220555
transform 1 0 2432 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5626_6
timestamp 1731220555
transform 1 0 2648 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5625_6
timestamp 1731220555
transform 1 0 2680 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5624_6
timestamp 1731220555
transform 1 0 2528 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5623_6
timestamp 1731220555
transform 1 0 2552 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5622_6
timestamp 1731220555
transform 1 0 2656 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5621_6
timestamp 1731220555
transform 1 0 2448 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5620_6
timestamp 1731220555
transform 1 0 2240 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5619_6
timestamp 1731220555
transform 1 0 2344 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5618_6
timestamp 1731220555
transform 1 0 2368 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5617_6
timestamp 1731220555
transform 1 0 2208 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5616_6
timestamp 1731220555
transform 1 0 2200 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5615_6
timestamp 1731220555
transform 1 0 2168 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5614_6
timestamp 1731220555
transform 1 0 2088 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5613_6
timestamp 1731220555
transform 1 0 2312 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5612_6
timestamp 1731220555
transform 1 0 2232 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5611_6
timestamp 1731220555
transform 1 0 2088 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5610_6
timestamp 1731220555
transform 1 0 1912 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5609_6
timestamp 1731220555
transform 1 0 1744 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5608_6
timestamp 1731220555
transform 1 0 1552 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5607_6
timestamp 1731220555
transform 1 0 1560 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5606_6
timestamp 1731220555
transform 1 0 1688 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5605_6
timestamp 1731220555
transform 1 0 1440 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5604_6
timestamp 1731220555
transform 1 0 1376 0 -1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5603_6
timestamp 1731220555
transform 1 0 1320 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5602_6
timestamp 1731220555
transform 1 0 1200 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5601_6
timestamp 1731220555
transform 1 0 1072 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5600_6
timestamp 1731220555
transform 1 0 808 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5599_6
timestamp 1731220555
transform 1 0 944 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5598_6
timestamp 1731220555
transform 1 0 1000 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5597_6
timestamp 1731220555
transform 1 0 1184 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5596_6
timestamp 1731220555
transform 1 0 1368 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5595_6
timestamp 1731220555
transform 1 0 1024 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5594_6
timestamp 1731220555
transform 1 0 1168 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5593_6
timestamp 1731220555
transform 1 0 1312 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5592_6
timestamp 1731220555
transform 1 0 1456 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5591_6
timestamp 1731220555
transform 1 0 1216 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5590_6
timestamp 1731220555
transform 1 0 1344 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5589_6
timestamp 1731220555
transform 1 0 1472 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5588_6
timestamp 1731220555
transform 1 0 1608 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5587_6
timestamp 1731220555
transform 1 0 1744 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5586_6
timestamp 1731220555
transform 1 0 1152 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5585_6
timestamp 1731220555
transform 1 0 1288 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5584_6
timestamp 1731220555
transform 1 0 1424 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5583_6
timestamp 1731220555
transform 1 0 1552 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5582_6
timestamp 1731220555
transform 1 0 1680 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5581_6
timestamp 1731220555
transform 1 0 1808 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5580_6
timestamp 1731220555
transform 1 0 1912 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5579_6
timestamp 1731220555
transform 1 0 1912 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5578_6
timestamp 1731220555
transform 1 0 1792 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5577_6
timestamp 1731220555
transform 1 0 1656 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5576_6
timestamp 1731220555
transform 1 0 1520 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5575_6
timestamp 1731220555
transform 1 0 1064 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5574_6
timestamp 1731220555
transform 1 0 1224 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5573_6
timestamp 1731220555
transform 1 0 1376 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5572_6
timestamp 1731220555
transform 1 0 1496 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5571_6
timestamp 1731220555
transform 1 0 1680 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5570_6
timestamp 1731220555
transform 1 0 1320 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5569_6
timestamp 1731220555
transform 1 0 960 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5568_6
timestamp 1731220555
transform 1 0 1144 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5567_6
timestamp 1731220555
transform 1 0 1240 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5566_6
timestamp 1731220555
transform 1 0 1344 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5565_6
timestamp 1731220555
transform 1 0 1448 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5564_6
timestamp 1731220555
transform 1 0 1136 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5563_6
timestamp 1731220555
transform 1 0 1032 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5562_6
timestamp 1731220555
transform 1 0 928 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5561_6
timestamp 1731220555
transform 1 0 824 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5560_6
timestamp 1731220555
transform 1 0 720 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5559_6
timestamp 1731220555
transform 1 0 616 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5558_6
timestamp 1731220555
transform 1 0 512 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5557_6
timestamp 1731220555
transform 1 0 408 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5556_6
timestamp 1731220555
transform 1 0 304 0 -1 4064
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5555_6
timestamp 1731220555
transform 1 0 152 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5554_6
timestamp 1731220555
transform 1 0 360 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5553_6
timestamp 1731220555
transform 1 0 568 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5552_6
timestamp 1731220555
transform 1 0 768 0 1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5551_6
timestamp 1731220555
transform 1 0 336 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5550_6
timestamp 1731220555
transform 1 0 528 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5549_6
timestamp 1731220555
transform 1 0 712 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5548_6
timestamp 1731220555
transform 1 0 896 0 -1 3916
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5547_6
timestamp 1731220555
transform 1 0 560 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5546_6
timestamp 1731220555
transform 1 0 712 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5545_6
timestamp 1731220555
transform 1 0 864 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5544_6
timestamp 1731220555
transform 1 0 1008 0 1 3772
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5543_6
timestamp 1731220555
transform 1 0 1088 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5542_6
timestamp 1731220555
transform 1 0 960 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5541_6
timestamp 1731220555
transform 1 0 824 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5540_6
timestamp 1731220555
transform 1 0 576 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5539_6
timestamp 1731220555
transform 1 0 696 0 -1 3760
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5538_6
timestamp 1731220555
transform 1 0 736 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5537_6
timestamp 1731220555
transform 1 0 880 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5536_6
timestamp 1731220555
transform 1 0 448 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5535_6
timestamp 1731220555
transform 1 0 592 0 1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5534_6
timestamp 1731220555
transform 1 0 656 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5533_6
timestamp 1731220555
transform 1 0 824 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5532_6
timestamp 1731220555
transform 1 0 496 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5531_6
timestamp 1731220555
transform 1 0 224 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5530_6
timestamp 1731220555
transform 1 0 352 0 -1 3612
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5529_6
timestamp 1731220555
transform 1 0 376 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5528_6
timestamp 1731220555
transform 1 0 520 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5527_6
timestamp 1731220555
transform 1 0 664 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5526_6
timestamp 1731220555
transform 1 0 128 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5525_6
timestamp 1731220555
transform 1 0 240 0 1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5524_6
timestamp 1731220555
transform 1 0 400 0 -1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5523_6
timestamp 1731220555
transform 1 0 720 0 -1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5522_6
timestamp 1731220555
transform 1 0 1048 0 -1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5521_6
timestamp 1731220555
transform 1 0 128 0 -1 3456
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5520_6
timestamp 1731220555
transform 1 0 128 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5519_6
timestamp 1731220555
transform 1 0 296 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5518_6
timestamp 1731220555
transform 1 0 504 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5517_6
timestamp 1731220555
transform 1 0 720 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5516_6
timestamp 1731220555
transform 1 0 936 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5515_6
timestamp 1731220555
transform 1 0 288 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5514_6
timestamp 1731220555
transform 1 0 456 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5513_6
timestamp 1731220555
transform 1 0 632 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5512_6
timestamp 1731220555
transform 1 0 824 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5511_6
timestamp 1731220555
transform 1 0 1016 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5510_6
timestamp 1731220555
transform 1 0 600 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5509_6
timestamp 1731220555
transform 1 0 736 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5508_6
timestamp 1731220555
transform 1 0 880 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5507_6
timestamp 1731220555
transform 1 0 1032 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5506_6
timestamp 1731220555
transform 1 0 1016 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5505_6
timestamp 1731220555
transform 1 0 888 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5504_6
timestamp 1731220555
transform 1 0 784 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5503_6
timestamp 1731220555
transform 1 0 680 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5502_6
timestamp 1731220555
transform 1 0 576 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5501_6
timestamp 1731220555
transform 1 0 616 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5500_6
timestamp 1731220555
transform 1 0 728 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5499_6
timestamp 1731220555
transform 1 0 288 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5498_6
timestamp 1731220555
transform 1 0 392 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5497_6
timestamp 1731220555
transform 1 0 504 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5496_6
timestamp 1731220555
transform 1 0 584 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5495_6
timestamp 1731220555
transform 1 0 760 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5494_6
timestamp 1731220555
transform 1 0 128 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5493_6
timestamp 1731220555
transform 1 0 248 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5492_6
timestamp 1731220555
transform 1 0 408 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5491_6
timestamp 1731220555
transform 1 0 424 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5490_6
timestamp 1731220555
transform 1 0 264 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5489_6
timestamp 1731220555
transform 1 0 128 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5488_6
timestamp 1731220555
transform 1 0 128 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5487_6
timestamp 1731220555
transform 1 0 296 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5486_6
timestamp 1731220555
transform 1 0 360 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5485_6
timestamp 1731220555
transform 1 0 160 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5484_6
timestamp 1731220555
transform 1 0 232 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5483_6
timestamp 1731220555
transform 1 0 400 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5482_6
timestamp 1731220555
transform 1 0 512 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5481_6
timestamp 1731220555
transform 1 0 296 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5480_6
timestamp 1731220555
transform 1 0 416 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5479_6
timestamp 1731220555
transform 1 0 256 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5478_6
timestamp 1731220555
transform 1 0 304 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5477_6
timestamp 1731220555
transform 1 0 448 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5476_6
timestamp 1731220555
transform 1 0 600 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5475_6
timestamp 1731220555
transform 1 0 584 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5474_6
timestamp 1731220555
transform 1 0 760 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5473_6
timestamp 1731220555
transform 1 0 936 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5472_6
timestamp 1731220555
transform 1 0 928 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5471_6
timestamp 1731220555
transform 1 0 720 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5470_6
timestamp 1731220555
transform 1 0 752 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5469_6
timestamp 1731220555
transform 1 0 936 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5468_6
timestamp 1731220555
transform 1 0 576 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5467_6
timestamp 1731220555
transform 1 0 560 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5466_6
timestamp 1731220555
transform 1 0 760 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5465_6
timestamp 1731220555
transform 1 0 848 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5464_6
timestamp 1731220555
transform 1 0 664 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5463_6
timestamp 1731220555
transform 1 0 480 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5462_6
timestamp 1731220555
transform 1 0 576 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5461_6
timestamp 1731220555
transform 1 0 736 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5460_6
timestamp 1731220555
transform 1 0 904 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5459_6
timestamp 1731220555
transform 1 0 936 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5458_6
timestamp 1731220555
transform 1 0 1080 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5457_6
timestamp 1731220555
transform 1 0 1264 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5456_6
timestamp 1731220555
transform 1 0 1456 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5455_6
timestamp 1731220555
transform 1 0 1408 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5454_6
timestamp 1731220555
transform 1 0 1216 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5453_6
timestamp 1731220555
transform 1 0 1032 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5452_6
timestamp 1731220555
transform 1 0 960 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5451_6
timestamp 1731220555
transform 1 0 1176 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5450_6
timestamp 1731220555
transform 1 0 1392 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5449_6
timestamp 1731220555
transform 1 0 1616 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5448_6
timestamp 1731220555
transform 1 0 1128 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5447_6
timestamp 1731220555
transform 1 0 1320 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5446_6
timestamp 1731220555
transform 1 0 1512 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5445_6
timestamp 1731220555
transform 1 0 1536 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5444_6
timestamp 1731220555
transform 1 0 1136 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5443_6
timestamp 1731220555
transform 1 0 1336 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5442_6
timestamp 1731220555
transform 1 0 1440 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5441_6
timestamp 1731220555
transform 1 0 1104 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5440_6
timestamp 1731220555
transform 1 0 1272 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5439_6
timestamp 1731220555
transform 1 0 1368 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5438_6
timestamp 1731220555
transform 1 0 1224 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5437_6
timestamp 1731220555
transform 1 0 1072 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5436_6
timestamp 1731220555
transform 1 0 1224 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5435_6
timestamp 1731220555
transform 1 0 1064 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5434_6
timestamp 1731220555
transform 1 0 1008 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5433_6
timestamp 1731220555
transform 1 0 1168 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5432_6
timestamp 1731220555
transform 1 0 1336 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5431_6
timestamp 1731220555
transform 1 0 1256 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5430_6
timestamp 1731220555
transform 1 0 1064 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5429_6
timestamp 1731220555
transform 1 0 1016 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5428_6
timestamp 1731220555
transform 1 0 1216 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5427_6
timestamp 1731220555
transform 1 0 1424 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5426_6
timestamp 1731220555
transform 1 0 1288 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5425_6
timestamp 1731220555
transform 1 0 1080 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5424_6
timestamp 1731220555
transform 1 0 800 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5423_6
timestamp 1731220555
transform 1 0 960 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5422_6
timestamp 1731220555
transform 1 0 1136 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5421_6
timestamp 1731220555
transform 1 0 1320 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5420_6
timestamp 1731220555
transform 1 0 1520 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5419_6
timestamp 1731220555
transform 1 0 896 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5418_6
timestamp 1731220555
transform 1 0 1080 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5417_6
timestamp 1731220555
transform 1 0 1280 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5416_6
timestamp 1731220555
transform 1 0 1488 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5415_6
timestamp 1731220555
transform 1 0 1712 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5414_6
timestamp 1731220555
transform 1 0 1088 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5413_6
timestamp 1731220555
transform 1 0 1256 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5412_6
timestamp 1731220555
transform 1 0 1432 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5411_6
timestamp 1731220555
transform 1 0 1608 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5410_6
timestamp 1731220555
transform 1 0 1168 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5409_6
timestamp 1731220555
transform 1 0 1360 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5408_6
timestamp 1731220555
transform 1 0 1544 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5407_6
timestamp 1731220555
transform 1 0 1720 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5406_6
timestamp 1731220555
transform 1 0 1904 0 -1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5405_6
timestamp 1731220555
transform 1 0 1912 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5404_6
timestamp 1731220555
transform 1 0 1744 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5403_6
timestamp 1731220555
transform 1 0 1584 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5402_6
timestamp 1731220555
transform 1 0 1256 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5401_6
timestamp 1731220555
transform 1 0 1424 0 1 1548
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5400_6
timestamp 1731220555
transform 1 0 1536 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5399_6
timestamp 1731220555
transform 1 0 1416 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5398_6
timestamp 1731220555
transform 1 0 1296 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5397_6
timestamp 1731220555
transform 1 0 1056 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5396_6
timestamp 1731220555
transform 1 0 1176 0 -1 1540
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5395_6
timestamp 1731220555
transform 1 0 1184 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5394_6
timestamp 1731220555
transform 1 0 1288 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5393_6
timestamp 1731220555
transform 1 0 1392 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5392_6
timestamp 1731220555
transform 1 0 1496 0 1 1384
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5391_6
timestamp 1731220555
transform 1 0 1288 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5390_6
timestamp 1731220555
transform 1 0 1408 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5389_6
timestamp 1731220555
transform 1 0 1528 0 -1 1376
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5388_6
timestamp 1731220555
transform 1 0 1560 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5387_6
timestamp 1731220555
transform 1 0 1384 0 1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5386_6
timestamp 1731220555
transform 1 0 1264 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5385_6
timestamp 1731220555
transform 1 0 1448 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5384_6
timestamp 1731220555
transform 1 0 1632 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5383_6
timestamp 1731220555
transform 1 0 1816 0 -1 1228
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5382_6
timestamp 1731220555
transform 1 0 1896 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5381_6
timestamp 1731220555
transform 1 0 1696 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5380_6
timestamp 1731220555
transform 1 0 1496 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5379_6
timestamp 1731220555
transform 1 0 1296 0 1 1076
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5378_6
timestamp 1731220555
transform 1 0 1104 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5377_6
timestamp 1731220555
transform 1 0 1264 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5376_6
timestamp 1731220555
transform 1 0 1472 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5375_6
timestamp 1731220555
transform 1 0 1120 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5374_6
timestamp 1731220555
transform 1 0 1312 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5373_6
timestamp 1731220555
transform 1 0 1504 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5372_6
timestamp 1731220555
transform 1 0 1696 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5371_6
timestamp 1731220555
transform 1 0 1888 0 -1 904
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5370_6
timestamp 1731220555
transform 1 0 1888 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5369_6
timestamp 1731220555
transform 1 0 1680 0 1 912
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5368_6
timestamp 1731220555
transform 1 0 1256 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5367_6
timestamp 1731220555
transform 1 0 1400 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5366_6
timestamp 1731220555
transform 1 0 1536 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5365_6
timestamp 1731220555
transform 1 0 1672 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5364_6
timestamp 1731220555
transform 1 0 1800 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5363_6
timestamp 1731220555
transform 1 0 1912 0 -1 1068
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5362_6
timestamp 1731220555
transform 1 0 2088 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5361_6
timestamp 1731220555
transform 1 0 2280 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5360_6
timestamp 1731220555
transform 1 0 2488 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5359_6
timestamp 1731220555
transform 1 0 2384 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5358_6
timestamp 1731220555
transform 1 0 2224 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5357_6
timestamp 1731220555
transform 1 0 2088 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5356_6
timestamp 1731220555
transform 1 0 2104 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5355_6
timestamp 1731220555
transform 1 0 2272 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5354_6
timestamp 1731220555
transform 1 0 2456 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5353_6
timestamp 1731220555
transform 1 0 2656 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5352_6
timestamp 1731220555
transform 1 0 2520 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5351_6
timestamp 1731220555
transform 1 0 2384 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5350_6
timestamp 1731220555
transform 1 0 2264 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5349_6
timestamp 1731220555
transform 1 0 2320 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5348_6
timestamp 1731220555
transform 1 0 2424 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5347_6
timestamp 1731220555
transform 1 0 2544 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5346_6
timestamp 1731220555
transform 1 0 2552 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5345_6
timestamp 1731220555
transform 1 0 2672 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5344_6
timestamp 1731220555
transform 1 0 2328 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5343_6
timestamp 1731220555
transform 1 0 2440 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5342_6
timestamp 1731220555
transform 1 0 2504 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5341_6
timestamp 1731220555
transform 1 0 2384 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5340_6
timestamp 1731220555
transform 1 0 2264 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5339_6
timestamp 1731220555
transform 1 0 2144 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5338_6
timestamp 1731220555
transform 1 0 2088 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5337_6
timestamp 1731220555
transform 1 0 2216 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5336_6
timestamp 1731220555
transform 1 0 2360 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5335_6
timestamp 1731220555
transform 1 0 2472 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5334_6
timestamp 1731220555
transform 1 0 2264 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5333_6
timestamp 1731220555
transform 1 0 2088 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5332_6
timestamp 1731220555
transform 1 0 2088 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5331_6
timestamp 1731220555
transform 1 0 1912 0 -1 1848
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5330_6
timestamp 1731220555
transform 1 0 1912 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5329_6
timestamp 1731220555
transform 1 0 1728 0 1 1856
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5328_6
timestamp 1731220555
transform 1 0 1504 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5327_6
timestamp 1731220555
transform 1 0 1720 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5326_6
timestamp 1731220555
transform 1 0 1912 0 -1 2012
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5325_6
timestamp 1731220555
transform 1 0 1856 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5324_6
timestamp 1731220555
transform 1 0 1640 0 1 2020
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5323_6
timestamp 1731220555
transform 1 0 1824 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5322_6
timestamp 1731220555
transform 1 0 1632 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5321_6
timestamp 1731220555
transform 1 0 1440 0 -1 2172
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5320_6
timestamp 1731220555
transform 1 0 1504 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5319_6
timestamp 1731220555
transform 1 0 1672 0 1 2184
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5318_6
timestamp 1731220555
transform 1 0 1752 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5317_6
timestamp 1731220555
transform 1 0 1568 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5316_6
timestamp 1731220555
transform 1 0 1392 0 -1 2340
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5315_6
timestamp 1731220555
transform 1 0 1512 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5314_6
timestamp 1731220555
transform 1 0 1648 0 1 2348
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5313_6
timestamp 1731220555
transform 1 0 1600 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5312_6
timestamp 1731220555
transform 1 0 1768 0 -1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5311_6
timestamp 1731220555
transform 1 0 1736 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5310_6
timestamp 1731220555
transform 1 0 1704 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5309_6
timestamp 1731220555
transform 1 0 1904 0 -1 2648
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5308_6
timestamp 1731220555
transform 1 0 1848 0 1 2656
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5307_6
timestamp 1731220555
transform 1 0 1808 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5306_6
timestamp 1731220555
transform 1 0 1608 0 -1 2804
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5305_6
timestamp 1731220555
transform 1 0 1648 0 1 2816
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5304_6
timestamp 1731220555
transform 1 0 1624 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5303_6
timestamp 1731220555
transform 1 0 1448 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5302_6
timestamp 1731220555
transform 1 0 1280 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5301_6
timestamp 1731220555
transform 1 0 1112 0 -1 2972
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5300_6
timestamp 1731220555
transform 1 0 1192 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5299_6
timestamp 1731220555
transform 1 0 1312 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5298_6
timestamp 1731220555
transform 1 0 840 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5297_6
timestamp 1731220555
transform 1 0 952 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5296_6
timestamp 1731220555
transform 1 0 1072 0 1 2980
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5295_6
timestamp 1731220555
transform 1 0 1160 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5294_6
timestamp 1731220555
transform 1 0 1336 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5293_6
timestamp 1731220555
transform 1 0 1528 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5292_6
timestamp 1731220555
transform 1 0 1728 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5291_6
timestamp 1731220555
transform 1 0 1480 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5290_6
timestamp 1731220555
transform 1 0 1328 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5289_6
timestamp 1731220555
transform 1 0 1184 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5288_6
timestamp 1731220555
transform 1 0 1208 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5287_6
timestamp 1731220555
transform 1 0 1408 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5286_6
timestamp 1731220555
transform 1 0 1608 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5285_6
timestamp 1731220555
transform 1 0 1144 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5284_6
timestamp 1731220555
transform 1 0 1344 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5283_6
timestamp 1731220555
transform 1 0 1536 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5282_6
timestamp 1731220555
transform 1 0 1728 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5281_6
timestamp 1731220555
transform 1 0 1912 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5280_6
timestamp 1731220555
transform 1 0 1808 0 -1 3280
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5279_6
timestamp 1731220555
transform 1 0 1632 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5278_6
timestamp 1731220555
transform 1 0 1784 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5277_6
timestamp 1731220555
transform 1 0 1912 0 1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5276_6
timestamp 1731220555
transform 1 0 1912 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5275_6
timestamp 1731220555
transform 1 0 2088 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5274_6
timestamp 1731220555
transform 1 0 2088 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5273_6
timestamp 1731220555
transform 1 0 2240 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5272_6
timestamp 1731220555
transform 1 0 2432 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5271_6
timestamp 1731220555
transform 1 0 2088 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5270_6
timestamp 1731220555
transform 1 0 2336 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5269_6
timestamp 1731220555
transform 1 0 2464 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5268_6
timestamp 1731220555
transform 1 0 2672 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5267_6
timestamp 1731220555
transform 1 0 2880 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5266_6
timestamp 1731220555
transform 1 0 2864 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5265_6
timestamp 1731220555
transform 1 0 2672 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5264_6
timestamp 1731220555
transform 1 0 2480 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5263_6
timestamp 1731220555
transform 1 0 2432 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5262_6
timestamp 1731220555
transform 1 0 2616 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5261_6
timestamp 1731220555
transform 1 0 2792 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5260_6
timestamp 1731220555
transform 1 0 2728 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5259_6
timestamp 1731220555
transform 1 0 2408 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5258_6
timestamp 1731220555
transform 1 0 2576 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5257_6
timestamp 1731220555
transform 1 0 2592 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5256_6
timestamp 1731220555
transform 1 0 2248 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5255_6
timestamp 1731220555
transform 1 0 2424 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5254_6
timestamp 1731220555
transform 1 0 2600 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5253_6
timestamp 1731220555
transform 1 0 2720 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5252_6
timestamp 1731220555
transform 1 0 2704 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5251_6
timestamp 1731220555
transform 1 0 2464 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5250_6
timestamp 1731220555
transform 1 0 2576 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5249_6
timestamp 1731220555
transform 1 0 2648 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5248_6
timestamp 1731220555
transform 1 0 2488 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5247_6
timestamp 1731220555
transform 1 0 2336 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5246_6
timestamp 1731220555
transform 1 0 2456 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5245_6
timestamp 1731220555
transform 1 0 2656 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5244_6
timestamp 1731220555
transform 1 0 2472 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5243_6
timestamp 1731220555
transform 1 0 2656 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5242_6
timestamp 1731220555
transform 1 0 2840 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5241_6
timestamp 1731220555
transform 1 0 2912 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5240_6
timestamp 1731220555
transform 1 0 2736 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5239_6
timestamp 1731220555
transform 1 0 2552 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5238_6
timestamp 1731220555
transform 1 0 2616 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5237_6
timestamp 1731220555
transform 1 0 2792 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5236_6
timestamp 1731220555
transform 1 0 2960 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5235_6
timestamp 1731220555
transform 1 0 2864 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5234_6
timestamp 1731220555
transform 1 0 2624 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5233_6
timestamp 1731220555
transform 1 0 2896 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5232_6
timestamp 1731220555
transform 1 0 2904 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5231_6
timestamp 1731220555
transform 1 0 2768 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5230_6
timestamp 1731220555
transform 1 0 2744 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5229_6
timestamp 1731220555
transform 1 0 2904 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5228_6
timestamp 1731220555
transform 1 0 2968 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5227_6
timestamp 1731220555
transform 1 0 3120 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5226_6
timestamp 1731220555
transform 1 0 3160 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5225_6
timestamp 1731220555
transform 1 0 2992 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5224_6
timestamp 1731220555
transform 1 0 3048 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5223_6
timestamp 1731220555
transform 1 0 2840 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5222_6
timestamp 1731220555
transform 1 0 3016 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5221_6
timestamp 1731220555
transform 1 0 3216 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5220_6
timestamp 1731220555
transform 1 0 3432 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5219_6
timestamp 1731220555
transform 1 0 3664 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5218_6
timestamp 1731220555
transform 1 0 2872 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5217_6
timestamp 1731220555
transform 1 0 3064 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5216_6
timestamp 1731220555
transform 1 0 3264 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5215_6
timestamp 1731220555
transform 1 0 3472 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5214_6
timestamp 1731220555
transform 1 0 3680 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5213_6
timestamp 1731220555
transform 1 0 3664 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5212_6
timestamp 1731220555
transform 1 0 3440 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5211_6
timestamp 1731220555
transform 1 0 3224 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5210_6
timestamp 1731220555
transform 1 0 3096 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5209_6
timestamp 1731220555
transform 1 0 3288 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5208_6
timestamp 1731220555
transform 1 0 3488 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5207_6
timestamp 1731220555
transform 1 0 3688 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5206_6
timestamp 1731220555
transform 1 0 3688 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5205_6
timestamp 1731220555
transform 1 0 3488 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5204_6
timestamp 1731220555
transform 1 0 3288 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5203_6
timestamp 1731220555
transform 1 0 3176 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5202_6
timestamp 1731220555
transform 1 0 3416 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5201_6
timestamp 1731220555
transform 1 0 3648 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5200_6
timestamp 1731220555
transform 1 0 3808 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5199_6
timestamp 1731220555
transform 1 0 3392 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5198_6
timestamp 1731220555
transform 1 0 3600 0 -1 720
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5197_6
timestamp 1731220555
transform 1 0 3656 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5196_6
timestamp 1731220555
transform 1 0 3800 0 -1 564
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5195_6
timestamp 1731220555
transform 1 0 3856 0 1 572
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5194_6
timestamp 1731220555
transform 1 0 3872 0 1 728
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5193_6
timestamp 1731220555
transform 1 0 3872 0 -1 872
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5192_6
timestamp 1731220555
transform 1 0 3872 0 1 884
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5191_6
timestamp 1731220555
transform 1 0 3872 0 -1 1032
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5190_6
timestamp 1731220555
transform 1 0 3872 0 1 1048
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5189_6
timestamp 1731220555
transform 1 0 3872 0 -1 1196
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5188_6
timestamp 1731220555
transform 1 0 3872 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5187_6
timestamp 1731220555
transform 1 0 3832 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5186_6
timestamp 1731220555
transform 1 0 3800 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5185_6
timestamp 1731220555
transform 1 0 3728 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5184_6
timestamp 1731220555
transform 1 0 3560 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5183_6
timestamp 1731220555
transform 1 0 3392 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5182_6
timestamp 1731220555
transform 1 0 3224 0 1 1208
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5181_6
timestamp 1731220555
transform 1 0 3328 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5180_6
timestamp 1731220555
transform 1 0 3496 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5179_6
timestamp 1731220555
transform 1 0 3664 0 -1 1360
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5178_6
timestamp 1731220555
transform 1 0 3624 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5177_6
timestamp 1731220555
transform 1 0 3448 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5176_6
timestamp 1731220555
transform 1 0 3280 0 1 1368
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5175_6
timestamp 1731220555
transform 1 0 3384 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5174_6
timestamp 1731220555
transform 1 0 3264 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5173_6
timestamp 1731220555
transform 1 0 3144 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5172_6
timestamp 1731220555
transform 1 0 3024 0 -1 1524
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5171_6
timestamp 1731220555
transform 1 0 2864 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5170_6
timestamp 1731220555
transform 1 0 2984 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5169_6
timestamp 1731220555
transform 1 0 3104 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5168_6
timestamp 1731220555
transform 1 0 3232 0 1 1532
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5167_6
timestamp 1731220555
transform 1 0 3328 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5166_6
timestamp 1731220555
transform 1 0 3184 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5165_6
timestamp 1731220555
transform 1 0 3040 0 -1 1688
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5164_6
timestamp 1731220555
transform 1 0 3096 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5163_6
timestamp 1731220555
transform 1 0 3296 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5162_6
timestamp 1731220555
transform 1 0 3264 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5161_6
timestamp 1731220555
transform 1 0 2864 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5160_6
timestamp 1731220555
transform 1 0 3072 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5159_6
timestamp 1731220555
transform 1 0 3080 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5158_6
timestamp 1731220555
transform 1 0 3288 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5157_6
timestamp 1731220555
transform 1 0 3440 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5156_6
timestamp 1731220555
transform 1 0 3744 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5155_6
timestamp 1731220555
transform 1 0 3688 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5154_6
timestamp 1731220555
transform 1 0 3488 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5153_6
timestamp 1731220555
transform 1 0 3592 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5152_6
timestamp 1731220555
transform 1 0 3432 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5151_6
timestamp 1731220555
transform 1 0 3488 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5150_6
timestamp 1731220555
transform 1 0 3680 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5149_6
timestamp 1731220555
transform 1 0 3872 0 1 1696
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5148_6
timestamp 1731220555
transform 1 0 3872 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5147_6
timestamp 1731220555
transform 1 0 3744 0 -1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5146_6
timestamp 1731220555
transform 1 0 3872 0 1 1840
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5145_6
timestamp 1731220555
transform 1 0 3872 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5144_6
timestamp 1731220555
transform 1 0 3872 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5143_6
timestamp 1731220555
transform 1 0 3872 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5142_6
timestamp 1731220555
transform 1 0 3872 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5141_6
timestamp 1731220555
transform 1 0 3872 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5140_6
timestamp 1731220555
transform 1 0 3872 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5139_6
timestamp 1731220555
transform 1 0 3872 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5138_6
timestamp 1731220555
transform 1 0 3744 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5137_6
timestamp 1731220555
transform 1 0 3440 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5136_6
timestamp 1731220555
transform 1 0 3592 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5135_6
timestamp 1731220555
transform 1 0 3656 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5134_6
timestamp 1731220555
transform 1 0 3664 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5133_6
timestamp 1731220555
transform 1 0 3680 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5132_6
timestamp 1731220555
transform 1 0 3544 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5131_6
timestamp 1731220555
transform 1 0 3720 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5130_6
timestamp 1731220555
transform 1 0 3728 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5129_6
timestamp 1731220555
transform 1 0 3560 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5128_6
timestamp 1731220555
transform 1 0 3592 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5127_6
timestamp 1731220555
transform 1 0 3288 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5126_6
timestamp 1731220555
transform 1 0 3128 0 -1 1992
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5125_6
timestamp 1731220555
transform 1 0 3240 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5124_6
timestamp 1731220555
transform 1 0 3400 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5123_6
timestamp 1731220555
transform 1 0 3080 0 1 2004
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5122_6
timestamp 1731220555
transform 1 0 3016 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5121_6
timestamp 1731220555
transform 1 0 3192 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5120_6
timestamp 1731220555
transform 1 0 3368 0 -1 2160
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5119_6
timestamp 1731220555
transform 1 0 3464 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5118_6
timestamp 1731220555
transform 1 0 3256 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5117_6
timestamp 1731220555
transform 1 0 2856 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5116_6
timestamp 1731220555
transform 1 0 3056 0 1 2168
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5115_6
timestamp 1731220555
transform 1 0 3224 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5114_6
timestamp 1731220555
transform 1 0 3440 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5113_6
timestamp 1731220555
transform 1 0 2824 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5112_6
timestamp 1731220555
transform 1 0 3016 0 -1 2320
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5111_6
timestamp 1731220555
transform 1 0 3032 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5110_6
timestamp 1731220555
transform 1 0 3224 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5109_6
timestamp 1731220555
transform 1 0 3432 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5108_6
timestamp 1731220555
transform 1 0 2856 0 1 2332
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5107_6
timestamp 1731220555
transform 1 0 2848 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5106_6
timestamp 1731220555
transform 1 0 2992 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5105_6
timestamp 1731220555
transform 1 0 3136 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5104_6
timestamp 1731220555
transform 1 0 3288 0 -1 2488
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5103_6
timestamp 1731220555
transform 1 0 2744 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5102_6
timestamp 1731220555
transform 1 0 2888 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5101_6
timestamp 1731220555
transform 1 0 3024 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_5100_6
timestamp 1731220555
transform 1 0 3160 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_599_6
timestamp 1731220555
transform 1 0 3296 0 1 2500
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_598_6
timestamp 1731220555
transform 1 0 2872 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_597_6
timestamp 1731220555
transform 1 0 3016 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_596_6
timestamp 1731220555
transform 1 0 3152 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_595_6
timestamp 1731220555
transform 1 0 3288 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_594_6
timestamp 1731220555
transform 1 0 3432 0 -1 2652
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_593_6
timestamp 1731220555
transform 1 0 2960 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_592_6
timestamp 1731220555
transform 1 0 3120 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_591_6
timestamp 1731220555
transform 1 0 3280 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_590_6
timestamp 1731220555
transform 1 0 3440 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_589_6
timestamp 1731220555
transform 1 0 3600 0 1 2664
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_588_6
timestamp 1731220555
transform 1 0 3056 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_587_6
timestamp 1731220555
transform 1 0 3240 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_586_6
timestamp 1731220555
transform 1 0 3416 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_585_6
timestamp 1731220555
transform 1 0 3592 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_584_6
timestamp 1731220555
transform 1 0 3768 0 -1 2820
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_583_6
timestamp 1731220555
transform 1 0 3088 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_582_6
timestamp 1731220555
transform 1 0 3280 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_581_6
timestamp 1731220555
transform 1 0 3472 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_580_6
timestamp 1731220555
transform 1 0 3664 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_579_6
timestamp 1731220555
transform 1 0 3856 0 1 2832
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_578_6
timestamp 1731220555
transform 1 0 3744 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_577_6
timestamp 1731220555
transform 1 0 3512 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_576_6
timestamp 1731220555
transform 1 0 3280 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_575_6
timestamp 1731220555
transform 1 0 3056 0 -1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_574_6
timestamp 1731220555
transform 1 0 3032 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_573_6
timestamp 1731220555
transform 1 0 3232 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_572_6
timestamp 1731220555
transform 1 0 3432 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_571_6
timestamp 1731220555
transform 1 0 3632 0 1 2984
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_570_6
timestamp 1731220555
transform 1 0 3544 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_569_6
timestamp 1731220555
transform 1 0 3352 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_568_6
timestamp 1731220555
transform 1 0 2776 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_567_6
timestamp 1731220555
transform 1 0 2976 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_566_6
timestamp 1731220555
transform 1 0 3168 0 -1 3132
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_565_6
timestamp 1731220555
transform 1 0 3224 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_564_6
timestamp 1731220555
transform 1 0 3368 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_563_6
timestamp 1731220555
transform 1 0 2816 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_562_6
timestamp 1731220555
transform 1 0 2952 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_561_6
timestamp 1731220555
transform 1 0 3088 0 1 3144
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_560_6
timestamp 1731220555
transform 1 0 3128 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_559_6
timestamp 1731220555
transform 1 0 3232 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_558_6
timestamp 1731220555
transform 1 0 3024 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_557_6
timestamp 1731220555
transform 1 0 2920 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_556_6
timestamp 1731220555
transform 1 0 2608 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_555_6
timestamp 1731220555
transform 1 0 2712 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_554_6
timestamp 1731220555
transform 1 0 2816 0 -1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_553_6
timestamp 1731220555
transform 1 0 2832 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_552_6
timestamp 1731220555
transform 1 0 2936 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_551_6
timestamp 1731220555
transform 1 0 2728 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_550_6
timestamp 1731220555
transform 1 0 2624 0 1 3288
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_549_6
timestamp 1731220555
transform 1 0 2544 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_548_6
timestamp 1731220555
transform 1 0 2648 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_547_6
timestamp 1731220555
transform 1 0 2752 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_546_6
timestamp 1731220555
transform 1 0 2856 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_545_6
timestamp 1731220555
transform 1 0 2960 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_544_6
timestamp 1731220555
transform 1 0 3064 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_543_6
timestamp 1731220555
transform 1 0 3168 0 -1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_542_6
timestamp 1731220555
transform 1 0 2680 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_541_6
timestamp 1731220555
transform 1 0 2808 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_540_6
timestamp 1731220555
transform 1 0 2928 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_539_6
timestamp 1731220555
transform 1 0 3048 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_538_6
timestamp 1731220555
transform 1 0 3176 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_537_6
timestamp 1731220555
transform 1 0 3304 0 1 3460
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_536_6
timestamp 1731220555
transform 1 0 2776 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_535_6
timestamp 1731220555
transform 1 0 2984 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_534_6
timestamp 1731220555
transform 1 0 3192 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_533_6
timestamp 1731220555
transform 1 0 3408 0 -1 3608
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_532_6
timestamp 1731220555
transform 1 0 2984 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_531_6
timestamp 1731220555
transform 1 0 3176 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_530_6
timestamp 1731220555
transform 1 0 3368 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_529_6
timestamp 1731220555
transform 1 0 3560 0 1 3620
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_528_6
timestamp 1731220555
transform 1 0 2952 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_527_6
timestamp 1731220555
transform 1 0 3136 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_526_6
timestamp 1731220555
transform 1 0 3304 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_525_6
timestamp 1731220555
transform 1 0 3456 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_524_6
timestamp 1731220555
transform 1 0 3192 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_523_6
timestamp 1731220555
transform 1 0 2736 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_522_6
timestamp 1731220555
transform 1 0 2976 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_521_6
timestamp 1731220555
transform 1 0 3048 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_520_6
timestamp 1731220555
transform 1 0 3224 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_519_6
timestamp 1731220555
transform 1 0 3392 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_518_6
timestamp 1731220555
transform 1 0 2856 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_517_6
timestamp 1731220555
transform 1 0 2824 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_516_6
timestamp 1731220555
transform 1 0 2960 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_515_6
timestamp 1731220555
transform 1 0 3096 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_514_6
timestamp 1731220555
transform 1 0 3224 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_513_6
timestamp 1731220555
transform 1 0 3344 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_512_6
timestamp 1731220555
transform 1 0 3456 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_511_6
timestamp 1731220555
transform 1 0 3576 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_510_6
timestamp 1731220555
transform 1 0 3696 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_59_6
timestamp 1731220555
transform 1 0 3816 0 1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_58_6
timestamp 1731220555
transform 1 0 3728 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_57_6
timestamp 1731220555
transform 1 0 3560 0 -1 3920
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_56_6
timestamp 1731220555
transform 1 0 3384 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_55_6
timestamp 1731220555
transform 1 0 3560 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_54_6
timestamp 1731220555
transform 1 0 3600 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_53_6
timestamp 1731220555
transform 1 0 3744 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_52_6
timestamp 1731220555
transform 1 0 3872 0 -1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_51_6
timestamp 1731220555
transform 1 0 3872 0 1 3776
box 8 5 100 68
use _0_0std_0_0cells_0_0LATCH  tst_50_6
timestamp 1731220555
transform 1 0 3728 0 1 3776
box 8 5 100 68
<< end >>
