magic
tech sky130l
timestamp 1731220412
<< m2 >>
rect 110 5729 116 5730
rect 1934 5729 1940 5730
rect 110 5725 111 5729
rect 115 5725 116 5729
rect 110 5724 116 5725
rect 158 5728 164 5729
rect 158 5724 159 5728
rect 163 5724 164 5728
rect 158 5723 164 5724
rect 294 5728 300 5729
rect 294 5724 295 5728
rect 299 5724 300 5728
rect 1934 5725 1935 5729
rect 1939 5725 1940 5729
rect 1934 5724 1940 5725
rect 294 5723 300 5724
rect 130 5713 136 5714
rect 110 5712 116 5713
rect 110 5708 111 5712
rect 115 5708 116 5712
rect 130 5709 131 5713
rect 135 5709 136 5713
rect 130 5708 136 5709
rect 266 5713 272 5714
rect 266 5709 267 5713
rect 271 5709 272 5713
rect 266 5708 272 5709
rect 1934 5712 1940 5713
rect 1934 5708 1935 5712
rect 1939 5708 1940 5712
rect 110 5707 116 5708
rect 1934 5707 1940 5708
rect 1974 5629 1980 5630
rect 3798 5629 3804 5630
rect 1974 5625 1975 5629
rect 1979 5625 1980 5629
rect 1974 5624 1980 5625
rect 2022 5628 2028 5629
rect 2022 5624 2023 5628
rect 2027 5624 2028 5628
rect 2022 5623 2028 5624
rect 2182 5628 2188 5629
rect 2182 5624 2183 5628
rect 2187 5624 2188 5628
rect 2182 5623 2188 5624
rect 2366 5628 2372 5629
rect 2366 5624 2367 5628
rect 2371 5624 2372 5628
rect 2366 5623 2372 5624
rect 2550 5628 2556 5629
rect 2550 5624 2551 5628
rect 2555 5624 2556 5628
rect 2550 5623 2556 5624
rect 2726 5628 2732 5629
rect 2726 5624 2727 5628
rect 2731 5624 2732 5628
rect 2726 5623 2732 5624
rect 2894 5628 2900 5629
rect 2894 5624 2895 5628
rect 2899 5624 2900 5628
rect 2894 5623 2900 5624
rect 3062 5628 3068 5629
rect 3062 5624 3063 5628
rect 3067 5624 3068 5628
rect 3062 5623 3068 5624
rect 3222 5628 3228 5629
rect 3222 5624 3223 5628
rect 3227 5624 3228 5628
rect 3222 5623 3228 5624
rect 3382 5628 3388 5629
rect 3382 5624 3383 5628
rect 3387 5624 3388 5628
rect 3382 5623 3388 5624
rect 3542 5628 3548 5629
rect 3542 5624 3543 5628
rect 3547 5624 3548 5628
rect 3542 5623 3548 5624
rect 3678 5628 3684 5629
rect 3678 5624 3679 5628
rect 3683 5624 3684 5628
rect 3798 5625 3799 5629
rect 3803 5625 3804 5629
rect 3798 5624 3804 5625
rect 3838 5625 3844 5626
rect 5662 5625 5668 5626
rect 3678 5623 3684 5624
rect 3838 5621 3839 5625
rect 3843 5621 3844 5625
rect 3838 5620 3844 5621
rect 4334 5624 4340 5625
rect 4334 5620 4335 5624
rect 4339 5620 4340 5624
rect 4334 5619 4340 5620
rect 4470 5624 4476 5625
rect 4470 5620 4471 5624
rect 4475 5620 4476 5624
rect 4470 5619 4476 5620
rect 4606 5624 4612 5625
rect 4606 5620 4607 5624
rect 4611 5620 4612 5624
rect 4606 5619 4612 5620
rect 4742 5624 4748 5625
rect 4742 5620 4743 5624
rect 4747 5620 4748 5624
rect 4742 5619 4748 5620
rect 4878 5624 4884 5625
rect 4878 5620 4879 5624
rect 4883 5620 4884 5624
rect 4878 5619 4884 5620
rect 5014 5624 5020 5625
rect 5014 5620 5015 5624
rect 5019 5620 5020 5624
rect 5662 5621 5663 5625
rect 5667 5621 5668 5625
rect 5662 5620 5668 5621
rect 5014 5619 5020 5620
rect 1994 5613 2000 5614
rect 1974 5612 1980 5613
rect 1974 5608 1975 5612
rect 1979 5608 1980 5612
rect 1994 5609 1995 5613
rect 1999 5609 2000 5613
rect 1994 5608 2000 5609
rect 2154 5613 2160 5614
rect 2154 5609 2155 5613
rect 2159 5609 2160 5613
rect 2154 5608 2160 5609
rect 2338 5613 2344 5614
rect 2338 5609 2339 5613
rect 2343 5609 2344 5613
rect 2338 5608 2344 5609
rect 2522 5613 2528 5614
rect 2522 5609 2523 5613
rect 2527 5609 2528 5613
rect 2522 5608 2528 5609
rect 2698 5613 2704 5614
rect 2698 5609 2699 5613
rect 2703 5609 2704 5613
rect 2698 5608 2704 5609
rect 2866 5613 2872 5614
rect 2866 5609 2867 5613
rect 2871 5609 2872 5613
rect 2866 5608 2872 5609
rect 3034 5613 3040 5614
rect 3034 5609 3035 5613
rect 3039 5609 3040 5613
rect 3034 5608 3040 5609
rect 3194 5613 3200 5614
rect 3194 5609 3195 5613
rect 3199 5609 3200 5613
rect 3194 5608 3200 5609
rect 3354 5613 3360 5614
rect 3354 5609 3355 5613
rect 3359 5609 3360 5613
rect 3354 5608 3360 5609
rect 3514 5613 3520 5614
rect 3514 5609 3515 5613
rect 3519 5609 3520 5613
rect 3514 5608 3520 5609
rect 3650 5613 3656 5614
rect 3650 5609 3651 5613
rect 3655 5609 3656 5613
rect 3650 5608 3656 5609
rect 3798 5612 3804 5613
rect 3798 5608 3799 5612
rect 3803 5608 3804 5612
rect 4306 5609 4312 5610
rect 1974 5607 1980 5608
rect 3798 5607 3804 5608
rect 3838 5608 3844 5609
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 4306 5605 4307 5609
rect 4311 5605 4312 5609
rect 4306 5604 4312 5605
rect 4442 5609 4448 5610
rect 4442 5605 4443 5609
rect 4447 5605 4448 5609
rect 4442 5604 4448 5605
rect 4578 5609 4584 5610
rect 4578 5605 4579 5609
rect 4583 5605 4584 5609
rect 4578 5604 4584 5605
rect 4714 5609 4720 5610
rect 4714 5605 4715 5609
rect 4719 5605 4720 5609
rect 4714 5604 4720 5605
rect 4850 5609 4856 5610
rect 4850 5605 4851 5609
rect 4855 5605 4856 5609
rect 4850 5604 4856 5605
rect 4986 5609 4992 5610
rect 4986 5605 4987 5609
rect 4991 5605 4992 5609
rect 4986 5604 4992 5605
rect 5662 5608 5668 5609
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 3838 5603 3844 5604
rect 5662 5603 5668 5604
rect 110 5580 116 5581
rect 1934 5580 1940 5581
rect 110 5576 111 5580
rect 115 5576 116 5580
rect 110 5575 116 5576
rect 130 5579 136 5580
rect 130 5575 131 5579
rect 135 5575 136 5579
rect 130 5574 136 5575
rect 274 5579 280 5580
rect 274 5575 275 5579
rect 279 5575 280 5579
rect 274 5574 280 5575
rect 474 5579 480 5580
rect 474 5575 475 5579
rect 479 5575 480 5579
rect 474 5574 480 5575
rect 698 5579 704 5580
rect 698 5575 699 5579
rect 703 5575 704 5579
rect 698 5574 704 5575
rect 954 5579 960 5580
rect 954 5575 955 5579
rect 959 5575 960 5579
rect 954 5574 960 5575
rect 1226 5579 1232 5580
rect 1226 5575 1227 5579
rect 1231 5575 1232 5579
rect 1226 5574 1232 5575
rect 1514 5579 1520 5580
rect 1514 5575 1515 5579
rect 1519 5575 1520 5579
rect 1514 5574 1520 5575
rect 1786 5579 1792 5580
rect 1786 5575 1787 5579
rect 1791 5575 1792 5579
rect 1934 5576 1935 5580
rect 1939 5576 1940 5580
rect 1934 5575 1940 5576
rect 1786 5574 1792 5575
rect 158 5564 164 5565
rect 110 5563 116 5564
rect 110 5559 111 5563
rect 115 5559 116 5563
rect 158 5560 159 5564
rect 163 5560 164 5564
rect 158 5559 164 5560
rect 302 5564 308 5565
rect 302 5560 303 5564
rect 307 5560 308 5564
rect 302 5559 308 5560
rect 502 5564 508 5565
rect 502 5560 503 5564
rect 507 5560 508 5564
rect 502 5559 508 5560
rect 726 5564 732 5565
rect 726 5560 727 5564
rect 731 5560 732 5564
rect 726 5559 732 5560
rect 982 5564 988 5565
rect 982 5560 983 5564
rect 987 5560 988 5564
rect 982 5559 988 5560
rect 1254 5564 1260 5565
rect 1254 5560 1255 5564
rect 1259 5560 1260 5564
rect 1254 5559 1260 5560
rect 1542 5564 1548 5565
rect 1542 5560 1543 5564
rect 1547 5560 1548 5564
rect 1542 5559 1548 5560
rect 1814 5564 1820 5565
rect 1814 5560 1815 5564
rect 1819 5560 1820 5564
rect 1814 5559 1820 5560
rect 1934 5563 1940 5564
rect 1934 5559 1935 5563
rect 1939 5559 1940 5563
rect 110 5558 116 5559
rect 1934 5558 1940 5559
rect 110 5505 116 5506
rect 1934 5505 1940 5506
rect 110 5501 111 5505
rect 115 5501 116 5505
rect 110 5500 116 5501
rect 278 5504 284 5505
rect 278 5500 279 5504
rect 283 5500 284 5504
rect 278 5499 284 5500
rect 518 5504 524 5505
rect 518 5500 519 5504
rect 523 5500 524 5504
rect 518 5499 524 5500
rect 766 5504 772 5505
rect 766 5500 767 5504
rect 771 5500 772 5504
rect 766 5499 772 5500
rect 1014 5504 1020 5505
rect 1014 5500 1015 5504
rect 1019 5500 1020 5504
rect 1014 5499 1020 5500
rect 1262 5504 1268 5505
rect 1262 5500 1263 5504
rect 1267 5500 1268 5504
rect 1262 5499 1268 5500
rect 1510 5504 1516 5505
rect 1510 5500 1511 5504
rect 1515 5500 1516 5504
rect 1510 5499 1516 5500
rect 1766 5504 1772 5505
rect 1766 5500 1767 5504
rect 1771 5500 1772 5504
rect 1934 5501 1935 5505
rect 1939 5501 1940 5505
rect 1934 5500 1940 5501
rect 1766 5499 1772 5500
rect 250 5489 256 5490
rect 110 5488 116 5489
rect 110 5484 111 5488
rect 115 5484 116 5488
rect 250 5485 251 5489
rect 255 5485 256 5489
rect 250 5484 256 5485
rect 490 5489 496 5490
rect 490 5485 491 5489
rect 495 5485 496 5489
rect 490 5484 496 5485
rect 738 5489 744 5490
rect 738 5485 739 5489
rect 743 5485 744 5489
rect 738 5484 744 5485
rect 986 5489 992 5490
rect 986 5485 987 5489
rect 991 5485 992 5489
rect 986 5484 992 5485
rect 1234 5489 1240 5490
rect 1234 5485 1235 5489
rect 1239 5485 1240 5489
rect 1234 5484 1240 5485
rect 1482 5489 1488 5490
rect 1482 5485 1483 5489
rect 1487 5485 1488 5489
rect 1482 5484 1488 5485
rect 1738 5489 1744 5490
rect 1738 5485 1739 5489
rect 1743 5485 1744 5489
rect 1738 5484 1744 5485
rect 1934 5488 1940 5489
rect 1934 5484 1935 5488
rect 1939 5484 1940 5488
rect 110 5483 116 5484
rect 1934 5483 1940 5484
rect 1974 5480 1980 5481
rect 3798 5480 3804 5481
rect 1974 5476 1975 5480
rect 1979 5476 1980 5480
rect 1974 5475 1980 5476
rect 2138 5479 2144 5480
rect 2138 5475 2139 5479
rect 2143 5475 2144 5479
rect 2138 5474 2144 5475
rect 2354 5479 2360 5480
rect 2354 5475 2355 5479
rect 2359 5475 2360 5479
rect 2354 5474 2360 5475
rect 2562 5479 2568 5480
rect 2562 5475 2563 5479
rect 2567 5475 2568 5479
rect 2562 5474 2568 5475
rect 2754 5479 2760 5480
rect 2754 5475 2755 5479
rect 2759 5475 2760 5479
rect 2754 5474 2760 5475
rect 2938 5479 2944 5480
rect 2938 5475 2939 5479
rect 2943 5475 2944 5479
rect 2938 5474 2944 5475
rect 3114 5479 3120 5480
rect 3114 5475 3115 5479
rect 3119 5475 3120 5479
rect 3114 5474 3120 5475
rect 3290 5479 3296 5480
rect 3290 5475 3291 5479
rect 3295 5475 3296 5479
rect 3290 5474 3296 5475
rect 3466 5479 3472 5480
rect 3466 5475 3467 5479
rect 3471 5475 3472 5479
rect 3466 5474 3472 5475
rect 3642 5479 3648 5480
rect 3642 5475 3643 5479
rect 3647 5475 3648 5479
rect 3798 5476 3799 5480
rect 3803 5476 3804 5480
rect 3798 5475 3804 5476
rect 3838 5476 3844 5477
rect 5662 5476 5668 5477
rect 3642 5474 3648 5475
rect 3838 5472 3839 5476
rect 3843 5472 3844 5476
rect 3838 5471 3844 5472
rect 4250 5475 4256 5476
rect 4250 5471 4251 5475
rect 4255 5471 4256 5475
rect 4250 5470 4256 5471
rect 4402 5475 4408 5476
rect 4402 5471 4403 5475
rect 4407 5471 4408 5475
rect 4402 5470 4408 5471
rect 4554 5475 4560 5476
rect 4554 5471 4555 5475
rect 4559 5471 4560 5475
rect 4554 5470 4560 5471
rect 4706 5475 4712 5476
rect 4706 5471 4707 5475
rect 4711 5471 4712 5475
rect 4706 5470 4712 5471
rect 4858 5475 4864 5476
rect 4858 5471 4859 5475
rect 4863 5471 4864 5475
rect 4858 5470 4864 5471
rect 5018 5475 5024 5476
rect 5018 5471 5019 5475
rect 5023 5471 5024 5475
rect 5662 5472 5663 5476
rect 5667 5472 5668 5476
rect 5662 5471 5668 5472
rect 5018 5470 5024 5471
rect 2166 5464 2172 5465
rect 1974 5463 1980 5464
rect 1974 5459 1975 5463
rect 1979 5459 1980 5463
rect 2166 5460 2167 5464
rect 2171 5460 2172 5464
rect 2166 5459 2172 5460
rect 2382 5464 2388 5465
rect 2382 5460 2383 5464
rect 2387 5460 2388 5464
rect 2382 5459 2388 5460
rect 2590 5464 2596 5465
rect 2590 5460 2591 5464
rect 2595 5460 2596 5464
rect 2590 5459 2596 5460
rect 2782 5464 2788 5465
rect 2782 5460 2783 5464
rect 2787 5460 2788 5464
rect 2782 5459 2788 5460
rect 2966 5464 2972 5465
rect 2966 5460 2967 5464
rect 2971 5460 2972 5464
rect 2966 5459 2972 5460
rect 3142 5464 3148 5465
rect 3142 5460 3143 5464
rect 3147 5460 3148 5464
rect 3142 5459 3148 5460
rect 3318 5464 3324 5465
rect 3318 5460 3319 5464
rect 3323 5460 3324 5464
rect 3318 5459 3324 5460
rect 3494 5464 3500 5465
rect 3494 5460 3495 5464
rect 3499 5460 3500 5464
rect 3494 5459 3500 5460
rect 3670 5464 3676 5465
rect 3670 5460 3671 5464
rect 3675 5460 3676 5464
rect 3670 5459 3676 5460
rect 3798 5463 3804 5464
rect 3798 5459 3799 5463
rect 3803 5459 3804 5463
rect 4278 5460 4284 5461
rect 1974 5458 1980 5459
rect 3798 5458 3804 5459
rect 3838 5459 3844 5460
rect 3838 5455 3839 5459
rect 3843 5455 3844 5459
rect 4278 5456 4279 5460
rect 4283 5456 4284 5460
rect 4278 5455 4284 5456
rect 4430 5460 4436 5461
rect 4430 5456 4431 5460
rect 4435 5456 4436 5460
rect 4430 5455 4436 5456
rect 4582 5460 4588 5461
rect 4582 5456 4583 5460
rect 4587 5456 4588 5460
rect 4582 5455 4588 5456
rect 4734 5460 4740 5461
rect 4734 5456 4735 5460
rect 4739 5456 4740 5460
rect 4734 5455 4740 5456
rect 4886 5460 4892 5461
rect 4886 5456 4887 5460
rect 4891 5456 4892 5460
rect 4886 5455 4892 5456
rect 5046 5460 5052 5461
rect 5046 5456 5047 5460
rect 5051 5456 5052 5460
rect 5046 5455 5052 5456
rect 5662 5459 5668 5460
rect 5662 5455 5663 5459
rect 5667 5455 5668 5459
rect 3838 5454 3844 5455
rect 5662 5454 5668 5455
rect 1974 5397 1980 5398
rect 3798 5397 3804 5398
rect 1974 5393 1975 5397
rect 1979 5393 1980 5397
rect 1974 5392 1980 5393
rect 2310 5396 2316 5397
rect 2310 5392 2311 5396
rect 2315 5392 2316 5396
rect 2310 5391 2316 5392
rect 2510 5396 2516 5397
rect 2510 5392 2511 5396
rect 2515 5392 2516 5396
rect 2510 5391 2516 5392
rect 2702 5396 2708 5397
rect 2702 5392 2703 5396
rect 2707 5392 2708 5396
rect 2702 5391 2708 5392
rect 2886 5396 2892 5397
rect 2886 5392 2887 5396
rect 2891 5392 2892 5396
rect 2886 5391 2892 5392
rect 3070 5396 3076 5397
rect 3070 5392 3071 5396
rect 3075 5392 3076 5396
rect 3070 5391 3076 5392
rect 3246 5396 3252 5397
rect 3246 5392 3247 5396
rect 3251 5392 3252 5396
rect 3246 5391 3252 5392
rect 3422 5396 3428 5397
rect 3422 5392 3423 5396
rect 3427 5392 3428 5396
rect 3422 5391 3428 5392
rect 3606 5396 3612 5397
rect 3606 5392 3607 5396
rect 3611 5392 3612 5396
rect 3798 5393 3799 5397
rect 3803 5393 3804 5397
rect 3798 5392 3804 5393
rect 3606 5391 3612 5392
rect 2282 5381 2288 5382
rect 1974 5380 1980 5381
rect 1974 5376 1975 5380
rect 1979 5376 1980 5380
rect 2282 5377 2283 5381
rect 2287 5377 2288 5381
rect 2282 5376 2288 5377
rect 2482 5381 2488 5382
rect 2482 5377 2483 5381
rect 2487 5377 2488 5381
rect 2482 5376 2488 5377
rect 2674 5381 2680 5382
rect 2674 5377 2675 5381
rect 2679 5377 2680 5381
rect 2674 5376 2680 5377
rect 2858 5381 2864 5382
rect 2858 5377 2859 5381
rect 2863 5377 2864 5381
rect 2858 5376 2864 5377
rect 3042 5381 3048 5382
rect 3042 5377 3043 5381
rect 3047 5377 3048 5381
rect 3042 5376 3048 5377
rect 3218 5381 3224 5382
rect 3218 5377 3219 5381
rect 3223 5377 3224 5381
rect 3218 5376 3224 5377
rect 3394 5381 3400 5382
rect 3394 5377 3395 5381
rect 3399 5377 3400 5381
rect 3394 5376 3400 5377
rect 3578 5381 3584 5382
rect 3838 5381 3844 5382
rect 5662 5381 5668 5382
rect 3578 5377 3579 5381
rect 3583 5377 3584 5381
rect 3578 5376 3584 5377
rect 3798 5380 3804 5381
rect 3798 5376 3799 5380
rect 3803 5376 3804 5380
rect 3838 5377 3839 5381
rect 3843 5377 3844 5381
rect 3838 5376 3844 5377
rect 4278 5380 4284 5381
rect 4278 5376 4279 5380
rect 4283 5376 4284 5380
rect 1974 5375 1980 5376
rect 3798 5375 3804 5376
rect 4278 5375 4284 5376
rect 4486 5380 4492 5381
rect 4486 5376 4487 5380
rect 4491 5376 4492 5380
rect 4486 5375 4492 5376
rect 4694 5380 4700 5381
rect 4694 5376 4695 5380
rect 4699 5376 4700 5380
rect 4694 5375 4700 5376
rect 4910 5380 4916 5381
rect 4910 5376 4911 5380
rect 4915 5376 4916 5380
rect 4910 5375 4916 5376
rect 5126 5380 5132 5381
rect 5126 5376 5127 5380
rect 5131 5376 5132 5380
rect 5662 5377 5663 5381
rect 5667 5377 5668 5381
rect 5662 5376 5668 5377
rect 5126 5375 5132 5376
rect 4250 5365 4256 5366
rect 3838 5364 3844 5365
rect 3838 5360 3839 5364
rect 3843 5360 3844 5364
rect 4250 5361 4251 5365
rect 4255 5361 4256 5365
rect 4250 5360 4256 5361
rect 4458 5365 4464 5366
rect 4458 5361 4459 5365
rect 4463 5361 4464 5365
rect 4458 5360 4464 5361
rect 4666 5365 4672 5366
rect 4666 5361 4667 5365
rect 4671 5361 4672 5365
rect 4666 5360 4672 5361
rect 4882 5365 4888 5366
rect 4882 5361 4883 5365
rect 4887 5361 4888 5365
rect 4882 5360 4888 5361
rect 5098 5365 5104 5366
rect 5098 5361 5099 5365
rect 5103 5361 5104 5365
rect 5098 5360 5104 5361
rect 5662 5364 5668 5365
rect 5662 5360 5663 5364
rect 5667 5360 5668 5364
rect 3838 5359 3844 5360
rect 5662 5359 5668 5360
rect 110 5356 116 5357
rect 1934 5356 1940 5357
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 110 5351 116 5352
rect 410 5355 416 5356
rect 410 5351 411 5355
rect 415 5351 416 5355
rect 410 5350 416 5351
rect 610 5355 616 5356
rect 610 5351 611 5355
rect 615 5351 616 5355
rect 610 5350 616 5351
rect 818 5355 824 5356
rect 818 5351 819 5355
rect 823 5351 824 5355
rect 818 5350 824 5351
rect 1034 5355 1040 5356
rect 1034 5351 1035 5355
rect 1039 5351 1040 5355
rect 1034 5350 1040 5351
rect 1258 5355 1264 5356
rect 1258 5351 1259 5355
rect 1263 5351 1264 5355
rect 1258 5350 1264 5351
rect 1490 5355 1496 5356
rect 1490 5351 1491 5355
rect 1495 5351 1496 5355
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 1934 5351 1940 5352
rect 1490 5350 1496 5351
rect 438 5340 444 5341
rect 110 5339 116 5340
rect 110 5335 111 5339
rect 115 5335 116 5339
rect 438 5336 439 5340
rect 443 5336 444 5340
rect 438 5335 444 5336
rect 638 5340 644 5341
rect 638 5336 639 5340
rect 643 5336 644 5340
rect 638 5335 644 5336
rect 846 5340 852 5341
rect 846 5336 847 5340
rect 851 5336 852 5340
rect 846 5335 852 5336
rect 1062 5340 1068 5341
rect 1062 5336 1063 5340
rect 1067 5336 1068 5340
rect 1062 5335 1068 5336
rect 1286 5340 1292 5341
rect 1286 5336 1287 5340
rect 1291 5336 1292 5340
rect 1286 5335 1292 5336
rect 1518 5340 1524 5341
rect 1518 5336 1519 5340
rect 1523 5336 1524 5340
rect 1518 5335 1524 5336
rect 1934 5339 1940 5340
rect 1934 5335 1935 5339
rect 1939 5335 1940 5339
rect 110 5334 116 5335
rect 1934 5334 1940 5335
rect 110 5281 116 5282
rect 1934 5281 1940 5282
rect 110 5277 111 5281
rect 115 5277 116 5281
rect 110 5276 116 5277
rect 590 5280 596 5281
rect 590 5276 591 5280
rect 595 5276 596 5280
rect 590 5275 596 5276
rect 726 5280 732 5281
rect 726 5276 727 5280
rect 731 5276 732 5280
rect 726 5275 732 5276
rect 862 5280 868 5281
rect 862 5276 863 5280
rect 867 5276 868 5280
rect 862 5275 868 5276
rect 998 5280 1004 5281
rect 998 5276 999 5280
rect 1003 5276 1004 5280
rect 998 5275 1004 5276
rect 1134 5280 1140 5281
rect 1134 5276 1135 5280
rect 1139 5276 1140 5280
rect 1134 5275 1140 5276
rect 1270 5280 1276 5281
rect 1270 5276 1271 5280
rect 1275 5276 1276 5280
rect 1270 5275 1276 5276
rect 1406 5280 1412 5281
rect 1406 5276 1407 5280
rect 1411 5276 1412 5280
rect 1406 5275 1412 5276
rect 1542 5280 1548 5281
rect 1542 5276 1543 5280
rect 1547 5276 1548 5280
rect 1934 5277 1935 5281
rect 1939 5277 1940 5281
rect 1934 5276 1940 5277
rect 1542 5275 1548 5276
rect 562 5265 568 5266
rect 110 5264 116 5265
rect 110 5260 111 5264
rect 115 5260 116 5264
rect 562 5261 563 5265
rect 567 5261 568 5265
rect 562 5260 568 5261
rect 698 5265 704 5266
rect 698 5261 699 5265
rect 703 5261 704 5265
rect 698 5260 704 5261
rect 834 5265 840 5266
rect 834 5261 835 5265
rect 839 5261 840 5265
rect 834 5260 840 5261
rect 970 5265 976 5266
rect 970 5261 971 5265
rect 975 5261 976 5265
rect 970 5260 976 5261
rect 1106 5265 1112 5266
rect 1106 5261 1107 5265
rect 1111 5261 1112 5265
rect 1106 5260 1112 5261
rect 1242 5265 1248 5266
rect 1242 5261 1243 5265
rect 1247 5261 1248 5265
rect 1242 5260 1248 5261
rect 1378 5265 1384 5266
rect 1378 5261 1379 5265
rect 1383 5261 1384 5265
rect 1378 5260 1384 5261
rect 1514 5265 1520 5266
rect 1514 5261 1515 5265
rect 1519 5261 1520 5265
rect 1514 5260 1520 5261
rect 1934 5264 1940 5265
rect 1934 5260 1935 5264
rect 1939 5260 1940 5264
rect 110 5259 116 5260
rect 1934 5259 1940 5260
rect 1974 5248 1980 5249
rect 3798 5248 3804 5249
rect 1974 5244 1975 5248
rect 1979 5244 1980 5248
rect 1974 5243 1980 5244
rect 2194 5247 2200 5248
rect 2194 5243 2195 5247
rect 2199 5243 2200 5247
rect 2194 5242 2200 5243
rect 2338 5247 2344 5248
rect 2338 5243 2339 5247
rect 2343 5243 2344 5247
rect 2338 5242 2344 5243
rect 2490 5247 2496 5248
rect 2490 5243 2491 5247
rect 2495 5243 2496 5247
rect 2490 5242 2496 5243
rect 2650 5247 2656 5248
rect 2650 5243 2651 5247
rect 2655 5243 2656 5247
rect 2650 5242 2656 5243
rect 2818 5247 2824 5248
rect 2818 5243 2819 5247
rect 2823 5243 2824 5247
rect 2818 5242 2824 5243
rect 3002 5247 3008 5248
rect 3002 5243 3003 5247
rect 3007 5243 3008 5247
rect 3002 5242 3008 5243
rect 3186 5247 3192 5248
rect 3186 5243 3187 5247
rect 3191 5243 3192 5247
rect 3186 5242 3192 5243
rect 3378 5247 3384 5248
rect 3378 5243 3379 5247
rect 3383 5243 3384 5247
rect 3378 5242 3384 5243
rect 3578 5247 3584 5248
rect 3578 5243 3579 5247
rect 3583 5243 3584 5247
rect 3798 5244 3799 5248
rect 3803 5244 3804 5248
rect 3798 5243 3804 5244
rect 3578 5242 3584 5243
rect 2222 5232 2228 5233
rect 1974 5231 1980 5232
rect 1974 5227 1975 5231
rect 1979 5227 1980 5231
rect 2222 5228 2223 5232
rect 2227 5228 2228 5232
rect 2222 5227 2228 5228
rect 2366 5232 2372 5233
rect 2366 5228 2367 5232
rect 2371 5228 2372 5232
rect 2366 5227 2372 5228
rect 2518 5232 2524 5233
rect 2518 5228 2519 5232
rect 2523 5228 2524 5232
rect 2518 5227 2524 5228
rect 2678 5232 2684 5233
rect 2678 5228 2679 5232
rect 2683 5228 2684 5232
rect 2678 5227 2684 5228
rect 2846 5232 2852 5233
rect 2846 5228 2847 5232
rect 2851 5228 2852 5232
rect 2846 5227 2852 5228
rect 3030 5232 3036 5233
rect 3030 5228 3031 5232
rect 3035 5228 3036 5232
rect 3030 5227 3036 5228
rect 3214 5232 3220 5233
rect 3214 5228 3215 5232
rect 3219 5228 3220 5232
rect 3214 5227 3220 5228
rect 3406 5232 3412 5233
rect 3406 5228 3407 5232
rect 3411 5228 3412 5232
rect 3406 5227 3412 5228
rect 3606 5232 3612 5233
rect 3606 5228 3607 5232
rect 3611 5228 3612 5232
rect 3606 5227 3612 5228
rect 3798 5231 3804 5232
rect 3798 5227 3799 5231
rect 3803 5227 3804 5231
rect 1974 5226 1980 5227
rect 3798 5226 3804 5227
rect 3838 5216 3844 5217
rect 5662 5216 5668 5217
rect 3838 5212 3839 5216
rect 3843 5212 3844 5216
rect 3838 5211 3844 5212
rect 4250 5215 4256 5216
rect 4250 5211 4251 5215
rect 4255 5211 4256 5215
rect 4250 5210 4256 5211
rect 4482 5215 4488 5216
rect 4482 5211 4483 5215
rect 4487 5211 4488 5215
rect 4482 5210 4488 5211
rect 4714 5215 4720 5216
rect 4714 5211 4715 5215
rect 4719 5211 4720 5215
rect 4714 5210 4720 5211
rect 4946 5215 4952 5216
rect 4946 5211 4947 5215
rect 4951 5211 4952 5215
rect 4946 5210 4952 5211
rect 5186 5215 5192 5216
rect 5186 5211 5187 5215
rect 5191 5211 5192 5215
rect 5662 5212 5663 5216
rect 5667 5212 5668 5216
rect 5662 5211 5668 5212
rect 5186 5210 5192 5211
rect 4278 5200 4284 5201
rect 3838 5199 3844 5200
rect 3838 5195 3839 5199
rect 3843 5195 3844 5199
rect 4278 5196 4279 5200
rect 4283 5196 4284 5200
rect 4278 5195 4284 5196
rect 4510 5200 4516 5201
rect 4510 5196 4511 5200
rect 4515 5196 4516 5200
rect 4510 5195 4516 5196
rect 4742 5200 4748 5201
rect 4742 5196 4743 5200
rect 4747 5196 4748 5200
rect 4742 5195 4748 5196
rect 4974 5200 4980 5201
rect 4974 5196 4975 5200
rect 4979 5196 4980 5200
rect 4974 5195 4980 5196
rect 5214 5200 5220 5201
rect 5214 5196 5215 5200
rect 5219 5196 5220 5200
rect 5214 5195 5220 5196
rect 5662 5199 5668 5200
rect 5662 5195 5663 5199
rect 5667 5195 5668 5199
rect 3838 5194 3844 5195
rect 5662 5194 5668 5195
rect 1974 5173 1980 5174
rect 3798 5173 3804 5174
rect 1974 5169 1975 5173
rect 1979 5169 1980 5173
rect 1974 5168 1980 5169
rect 2022 5172 2028 5173
rect 2022 5168 2023 5172
rect 2027 5168 2028 5172
rect 2022 5167 2028 5168
rect 2158 5172 2164 5173
rect 2158 5168 2159 5172
rect 2163 5168 2164 5172
rect 2158 5167 2164 5168
rect 2326 5172 2332 5173
rect 2326 5168 2327 5172
rect 2331 5168 2332 5172
rect 2326 5167 2332 5168
rect 2510 5172 2516 5173
rect 2510 5168 2511 5172
rect 2515 5168 2516 5172
rect 2510 5167 2516 5168
rect 2694 5172 2700 5173
rect 2694 5168 2695 5172
rect 2699 5168 2700 5172
rect 2694 5167 2700 5168
rect 2886 5172 2892 5173
rect 2886 5168 2887 5172
rect 2891 5168 2892 5172
rect 2886 5167 2892 5168
rect 3086 5172 3092 5173
rect 3086 5168 3087 5172
rect 3091 5168 3092 5172
rect 3086 5167 3092 5168
rect 3286 5172 3292 5173
rect 3286 5168 3287 5172
rect 3291 5168 3292 5172
rect 3286 5167 3292 5168
rect 3494 5172 3500 5173
rect 3494 5168 3495 5172
rect 3499 5168 3500 5172
rect 3494 5167 3500 5168
rect 3678 5172 3684 5173
rect 3678 5168 3679 5172
rect 3683 5168 3684 5172
rect 3798 5169 3799 5173
rect 3803 5169 3804 5173
rect 3798 5168 3804 5169
rect 3678 5167 3684 5168
rect 1994 5157 2000 5158
rect 1974 5156 1980 5157
rect 1974 5152 1975 5156
rect 1979 5152 1980 5156
rect 1994 5153 1995 5157
rect 1999 5153 2000 5157
rect 1994 5152 2000 5153
rect 2130 5157 2136 5158
rect 2130 5153 2131 5157
rect 2135 5153 2136 5157
rect 2130 5152 2136 5153
rect 2298 5157 2304 5158
rect 2298 5153 2299 5157
rect 2303 5153 2304 5157
rect 2298 5152 2304 5153
rect 2482 5157 2488 5158
rect 2482 5153 2483 5157
rect 2487 5153 2488 5157
rect 2482 5152 2488 5153
rect 2666 5157 2672 5158
rect 2666 5153 2667 5157
rect 2671 5153 2672 5157
rect 2666 5152 2672 5153
rect 2858 5157 2864 5158
rect 2858 5153 2859 5157
rect 2863 5153 2864 5157
rect 2858 5152 2864 5153
rect 3058 5157 3064 5158
rect 3058 5153 3059 5157
rect 3063 5153 3064 5157
rect 3058 5152 3064 5153
rect 3258 5157 3264 5158
rect 3258 5153 3259 5157
rect 3263 5153 3264 5157
rect 3258 5152 3264 5153
rect 3466 5157 3472 5158
rect 3466 5153 3467 5157
rect 3471 5153 3472 5157
rect 3466 5152 3472 5153
rect 3650 5157 3656 5158
rect 3650 5153 3651 5157
rect 3655 5153 3656 5157
rect 3650 5152 3656 5153
rect 3798 5156 3804 5157
rect 3798 5152 3799 5156
rect 3803 5152 3804 5156
rect 1974 5151 1980 5152
rect 3798 5151 3804 5152
rect 3838 5113 3844 5114
rect 5662 5113 5668 5114
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 3886 5107 3892 5108
rect 4134 5112 4140 5113
rect 4134 5108 4135 5112
rect 4139 5108 4140 5112
rect 4134 5107 4140 5108
rect 4406 5112 4412 5113
rect 4406 5108 4407 5112
rect 4411 5108 4412 5112
rect 4406 5107 4412 5108
rect 4678 5112 4684 5113
rect 4678 5108 4679 5112
rect 4683 5108 4684 5112
rect 4678 5107 4684 5108
rect 4958 5112 4964 5113
rect 4958 5108 4959 5112
rect 4963 5108 4964 5112
rect 4958 5107 4964 5108
rect 5238 5112 5244 5113
rect 5238 5108 5239 5112
rect 5243 5108 5244 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5238 5107 5244 5108
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4106 5097 4112 5098
rect 4106 5093 4107 5097
rect 4111 5093 4112 5097
rect 4106 5092 4112 5093
rect 4378 5097 4384 5098
rect 4378 5093 4379 5097
rect 4383 5093 4384 5097
rect 4378 5092 4384 5093
rect 4650 5097 4656 5098
rect 4650 5093 4651 5097
rect 4655 5093 4656 5097
rect 4650 5092 4656 5093
rect 4930 5097 4936 5098
rect 4930 5093 4931 5097
rect 4935 5093 4936 5097
rect 4930 5092 4936 5093
rect 5210 5097 5216 5098
rect 5210 5093 5211 5097
rect 5215 5093 5216 5097
rect 5210 5092 5216 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 3838 5091 3844 5092
rect 5662 5091 5668 5092
rect 110 5028 116 5029
rect 1934 5028 1940 5029
rect 110 5024 111 5028
rect 115 5024 116 5028
rect 110 5023 116 5024
rect 346 5027 352 5028
rect 346 5023 347 5027
rect 351 5023 352 5027
rect 346 5022 352 5023
rect 482 5027 488 5028
rect 482 5023 483 5027
rect 487 5023 488 5027
rect 482 5022 488 5023
rect 618 5027 624 5028
rect 618 5023 619 5027
rect 623 5023 624 5027
rect 618 5022 624 5023
rect 754 5027 760 5028
rect 754 5023 755 5027
rect 759 5023 760 5027
rect 754 5022 760 5023
rect 890 5027 896 5028
rect 890 5023 891 5027
rect 895 5023 896 5027
rect 890 5022 896 5023
rect 1034 5027 1040 5028
rect 1034 5023 1035 5027
rect 1039 5023 1040 5027
rect 1034 5022 1040 5023
rect 1186 5027 1192 5028
rect 1186 5023 1187 5027
rect 1191 5023 1192 5027
rect 1186 5022 1192 5023
rect 1338 5027 1344 5028
rect 1338 5023 1339 5027
rect 1343 5023 1344 5027
rect 1338 5022 1344 5023
rect 1490 5027 1496 5028
rect 1490 5023 1491 5027
rect 1495 5023 1496 5027
rect 1490 5022 1496 5023
rect 1650 5027 1656 5028
rect 1650 5023 1651 5027
rect 1655 5023 1656 5027
rect 1650 5022 1656 5023
rect 1786 5027 1792 5028
rect 1786 5023 1787 5027
rect 1791 5023 1792 5027
rect 1934 5024 1935 5028
rect 1939 5024 1940 5028
rect 1934 5023 1940 5024
rect 1974 5024 1980 5025
rect 3798 5024 3804 5025
rect 1786 5022 1792 5023
rect 1974 5020 1975 5024
rect 1979 5020 1980 5024
rect 1974 5019 1980 5020
rect 1994 5023 2000 5024
rect 1994 5019 1995 5023
rect 1999 5019 2000 5023
rect 1994 5018 2000 5019
rect 2530 5023 2536 5024
rect 2530 5019 2531 5023
rect 2535 5019 2536 5023
rect 2530 5018 2536 5019
rect 3098 5023 3104 5024
rect 3098 5019 3099 5023
rect 3103 5019 3104 5023
rect 3098 5018 3104 5019
rect 3650 5023 3656 5024
rect 3650 5019 3651 5023
rect 3655 5019 3656 5023
rect 3798 5020 3799 5024
rect 3803 5020 3804 5024
rect 3798 5019 3804 5020
rect 3650 5018 3656 5019
rect 374 5012 380 5013
rect 110 5011 116 5012
rect 110 5007 111 5011
rect 115 5007 116 5011
rect 374 5008 375 5012
rect 379 5008 380 5012
rect 374 5007 380 5008
rect 510 5012 516 5013
rect 510 5008 511 5012
rect 515 5008 516 5012
rect 510 5007 516 5008
rect 646 5012 652 5013
rect 646 5008 647 5012
rect 651 5008 652 5012
rect 646 5007 652 5008
rect 782 5012 788 5013
rect 782 5008 783 5012
rect 787 5008 788 5012
rect 782 5007 788 5008
rect 918 5012 924 5013
rect 918 5008 919 5012
rect 923 5008 924 5012
rect 918 5007 924 5008
rect 1062 5012 1068 5013
rect 1062 5008 1063 5012
rect 1067 5008 1068 5012
rect 1062 5007 1068 5008
rect 1214 5012 1220 5013
rect 1214 5008 1215 5012
rect 1219 5008 1220 5012
rect 1214 5007 1220 5008
rect 1366 5012 1372 5013
rect 1366 5008 1367 5012
rect 1371 5008 1372 5012
rect 1366 5007 1372 5008
rect 1518 5012 1524 5013
rect 1518 5008 1519 5012
rect 1523 5008 1524 5012
rect 1518 5007 1524 5008
rect 1678 5012 1684 5013
rect 1678 5008 1679 5012
rect 1683 5008 1684 5012
rect 1678 5007 1684 5008
rect 1814 5012 1820 5013
rect 1814 5008 1815 5012
rect 1819 5008 1820 5012
rect 1814 5007 1820 5008
rect 1934 5011 1940 5012
rect 1934 5007 1935 5011
rect 1939 5007 1940 5011
rect 2022 5008 2028 5009
rect 110 5006 116 5007
rect 1934 5006 1940 5007
rect 1974 5007 1980 5008
rect 1974 5003 1975 5007
rect 1979 5003 1980 5007
rect 2022 5004 2023 5008
rect 2027 5004 2028 5008
rect 2022 5003 2028 5004
rect 2558 5008 2564 5009
rect 2558 5004 2559 5008
rect 2563 5004 2564 5008
rect 2558 5003 2564 5004
rect 3126 5008 3132 5009
rect 3126 5004 3127 5008
rect 3131 5004 3132 5008
rect 3126 5003 3132 5004
rect 3678 5008 3684 5009
rect 3678 5004 3679 5008
rect 3683 5004 3684 5008
rect 3678 5003 3684 5004
rect 3798 5007 3804 5008
rect 3798 5003 3799 5007
rect 3803 5003 3804 5007
rect 1974 5002 1980 5003
rect 3798 5002 3804 5003
rect 110 4953 116 4954
rect 1934 4953 1940 4954
rect 110 4949 111 4953
rect 115 4949 116 4953
rect 110 4948 116 4949
rect 158 4952 164 4953
rect 158 4948 159 4952
rect 163 4948 164 4952
rect 158 4947 164 4948
rect 342 4952 348 4953
rect 342 4948 343 4952
rect 347 4948 348 4952
rect 342 4947 348 4948
rect 550 4952 556 4953
rect 550 4948 551 4952
rect 555 4948 556 4952
rect 550 4947 556 4948
rect 750 4952 756 4953
rect 750 4948 751 4952
rect 755 4948 756 4952
rect 750 4947 756 4948
rect 942 4952 948 4953
rect 942 4948 943 4952
rect 947 4948 948 4952
rect 942 4947 948 4948
rect 1126 4952 1132 4953
rect 1126 4948 1127 4952
rect 1131 4948 1132 4952
rect 1126 4947 1132 4948
rect 1310 4952 1316 4953
rect 1310 4948 1311 4952
rect 1315 4948 1316 4952
rect 1310 4947 1316 4948
rect 1486 4952 1492 4953
rect 1486 4948 1487 4952
rect 1491 4948 1492 4952
rect 1486 4947 1492 4948
rect 1662 4952 1668 4953
rect 1662 4948 1663 4952
rect 1667 4948 1668 4952
rect 1662 4947 1668 4948
rect 1814 4952 1820 4953
rect 1814 4948 1815 4952
rect 1819 4948 1820 4952
rect 1934 4949 1935 4953
rect 1939 4949 1940 4953
rect 1934 4948 1940 4949
rect 3838 4952 3844 4953
rect 5662 4952 5668 4953
rect 3838 4948 3839 4952
rect 3843 4948 3844 4952
rect 1814 4947 1820 4948
rect 3838 4947 3844 4948
rect 3858 4951 3864 4952
rect 3858 4947 3859 4951
rect 3863 4947 3864 4951
rect 3858 4946 3864 4947
rect 4018 4951 4024 4952
rect 4018 4947 4019 4951
rect 4023 4947 4024 4951
rect 4018 4946 4024 4947
rect 4210 4951 4216 4952
rect 4210 4947 4211 4951
rect 4215 4947 4216 4951
rect 4210 4946 4216 4947
rect 4410 4951 4416 4952
rect 4410 4947 4411 4951
rect 4415 4947 4416 4951
rect 4410 4946 4416 4947
rect 4626 4951 4632 4952
rect 4626 4947 4627 4951
rect 4631 4947 4632 4951
rect 4626 4946 4632 4947
rect 4842 4951 4848 4952
rect 4842 4947 4843 4951
rect 4847 4947 4848 4951
rect 4842 4946 4848 4947
rect 5066 4951 5072 4952
rect 5066 4947 5067 4951
rect 5071 4947 5072 4951
rect 5066 4946 5072 4947
rect 5298 4951 5304 4952
rect 5298 4947 5299 4951
rect 5303 4947 5304 4951
rect 5662 4948 5663 4952
rect 5667 4948 5668 4952
rect 5662 4947 5668 4948
rect 5298 4946 5304 4947
rect 130 4937 136 4938
rect 110 4936 116 4937
rect 110 4932 111 4936
rect 115 4932 116 4936
rect 130 4933 131 4937
rect 135 4933 136 4937
rect 130 4932 136 4933
rect 314 4937 320 4938
rect 314 4933 315 4937
rect 319 4933 320 4937
rect 314 4932 320 4933
rect 522 4937 528 4938
rect 522 4933 523 4937
rect 527 4933 528 4937
rect 522 4932 528 4933
rect 722 4937 728 4938
rect 722 4933 723 4937
rect 727 4933 728 4937
rect 722 4932 728 4933
rect 914 4937 920 4938
rect 914 4933 915 4937
rect 919 4933 920 4937
rect 914 4932 920 4933
rect 1098 4937 1104 4938
rect 1098 4933 1099 4937
rect 1103 4933 1104 4937
rect 1098 4932 1104 4933
rect 1282 4937 1288 4938
rect 1282 4933 1283 4937
rect 1287 4933 1288 4937
rect 1282 4932 1288 4933
rect 1458 4937 1464 4938
rect 1458 4933 1459 4937
rect 1463 4933 1464 4937
rect 1458 4932 1464 4933
rect 1634 4937 1640 4938
rect 1634 4933 1635 4937
rect 1639 4933 1640 4937
rect 1634 4932 1640 4933
rect 1786 4937 1792 4938
rect 1786 4933 1787 4937
rect 1791 4933 1792 4937
rect 1786 4932 1792 4933
rect 1934 4936 1940 4937
rect 3886 4936 3892 4937
rect 1934 4932 1935 4936
rect 1939 4932 1940 4936
rect 110 4931 116 4932
rect 1934 4931 1940 4932
rect 3838 4935 3844 4936
rect 3838 4931 3839 4935
rect 3843 4931 3844 4935
rect 3886 4932 3887 4936
rect 3891 4932 3892 4936
rect 3886 4931 3892 4932
rect 4046 4936 4052 4937
rect 4046 4932 4047 4936
rect 4051 4932 4052 4936
rect 4046 4931 4052 4932
rect 4238 4936 4244 4937
rect 4238 4932 4239 4936
rect 4243 4932 4244 4936
rect 4238 4931 4244 4932
rect 4438 4936 4444 4937
rect 4438 4932 4439 4936
rect 4443 4932 4444 4936
rect 4438 4931 4444 4932
rect 4654 4936 4660 4937
rect 4654 4932 4655 4936
rect 4659 4932 4660 4936
rect 4654 4931 4660 4932
rect 4870 4936 4876 4937
rect 4870 4932 4871 4936
rect 4875 4932 4876 4936
rect 4870 4931 4876 4932
rect 5094 4936 5100 4937
rect 5094 4932 5095 4936
rect 5099 4932 5100 4936
rect 5094 4931 5100 4932
rect 5326 4936 5332 4937
rect 5326 4932 5327 4936
rect 5331 4932 5332 4936
rect 5326 4931 5332 4932
rect 5662 4935 5668 4936
rect 5662 4931 5663 4935
rect 5667 4931 5668 4935
rect 3838 4930 3844 4931
rect 5662 4930 5668 4931
rect 1974 4917 1980 4918
rect 3798 4917 3804 4918
rect 1974 4913 1975 4917
rect 1979 4913 1980 4917
rect 1974 4912 1980 4913
rect 2870 4916 2876 4917
rect 2870 4912 2871 4916
rect 2875 4912 2876 4916
rect 2870 4911 2876 4912
rect 3006 4916 3012 4917
rect 3006 4912 3007 4916
rect 3011 4912 3012 4916
rect 3798 4913 3799 4917
rect 3803 4913 3804 4917
rect 3798 4912 3804 4913
rect 3006 4911 3012 4912
rect 2842 4901 2848 4902
rect 1974 4900 1980 4901
rect 1974 4896 1975 4900
rect 1979 4896 1980 4900
rect 2842 4897 2843 4901
rect 2847 4897 2848 4901
rect 2842 4896 2848 4897
rect 2978 4901 2984 4902
rect 2978 4897 2979 4901
rect 2983 4897 2984 4901
rect 2978 4896 2984 4897
rect 3798 4900 3804 4901
rect 3798 4896 3799 4900
rect 3803 4896 3804 4900
rect 1974 4895 1980 4896
rect 3798 4895 3804 4896
rect 3838 4857 3844 4858
rect 5662 4857 5668 4858
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3886 4856 3892 4857
rect 3886 4852 3887 4856
rect 3891 4852 3892 4856
rect 3886 4851 3892 4852
rect 4070 4856 4076 4857
rect 4070 4852 4071 4856
rect 4075 4852 4076 4856
rect 4070 4851 4076 4852
rect 4286 4856 4292 4857
rect 4286 4852 4287 4856
rect 4291 4852 4292 4856
rect 4286 4851 4292 4852
rect 4510 4856 4516 4857
rect 4510 4852 4511 4856
rect 4515 4852 4516 4856
rect 4510 4851 4516 4852
rect 4734 4856 4740 4857
rect 4734 4852 4735 4856
rect 4739 4852 4740 4856
rect 4734 4851 4740 4852
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5182 4856 5188 4857
rect 5182 4852 5183 4856
rect 5187 4852 5188 4856
rect 5182 4851 5188 4852
rect 5406 4856 5412 4857
rect 5406 4852 5407 4856
rect 5411 4852 5412 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5406 4851 5412 4852
rect 3858 4841 3864 4842
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3858 4837 3859 4841
rect 3863 4837 3864 4841
rect 3858 4836 3864 4837
rect 4042 4841 4048 4842
rect 4042 4837 4043 4841
rect 4047 4837 4048 4841
rect 4042 4836 4048 4837
rect 4258 4841 4264 4842
rect 4258 4837 4259 4841
rect 4263 4837 4264 4841
rect 4258 4836 4264 4837
rect 4482 4841 4488 4842
rect 4482 4837 4483 4841
rect 4487 4837 4488 4841
rect 4482 4836 4488 4837
rect 4706 4841 4712 4842
rect 4706 4837 4707 4841
rect 4711 4837 4712 4841
rect 4706 4836 4712 4837
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5154 4841 5160 4842
rect 5154 4837 5155 4841
rect 5159 4837 5160 4841
rect 5154 4836 5160 4837
rect 5378 4841 5384 4842
rect 5378 4837 5379 4841
rect 5383 4837 5384 4841
rect 5378 4836 5384 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 3838 4835 3844 4836
rect 5662 4835 5668 4836
rect 110 4796 116 4797
rect 1934 4796 1940 4797
rect 110 4792 111 4796
rect 115 4792 116 4796
rect 110 4791 116 4792
rect 130 4795 136 4796
rect 130 4791 131 4795
rect 135 4791 136 4795
rect 130 4790 136 4791
rect 266 4795 272 4796
rect 266 4791 267 4795
rect 271 4791 272 4795
rect 266 4790 272 4791
rect 402 4795 408 4796
rect 402 4791 403 4795
rect 407 4791 408 4795
rect 402 4790 408 4791
rect 538 4795 544 4796
rect 538 4791 539 4795
rect 543 4791 544 4795
rect 538 4790 544 4791
rect 674 4795 680 4796
rect 674 4791 675 4795
rect 679 4791 680 4795
rect 1934 4792 1935 4796
rect 1939 4792 1940 4796
rect 1934 4791 1940 4792
rect 674 4790 680 4791
rect 158 4780 164 4781
rect 110 4779 116 4780
rect 110 4775 111 4779
rect 115 4775 116 4779
rect 158 4776 159 4780
rect 163 4776 164 4780
rect 158 4775 164 4776
rect 294 4780 300 4781
rect 294 4776 295 4780
rect 299 4776 300 4780
rect 294 4775 300 4776
rect 430 4780 436 4781
rect 430 4776 431 4780
rect 435 4776 436 4780
rect 430 4775 436 4776
rect 566 4780 572 4781
rect 566 4776 567 4780
rect 571 4776 572 4780
rect 566 4775 572 4776
rect 702 4780 708 4781
rect 702 4776 703 4780
rect 707 4776 708 4780
rect 702 4775 708 4776
rect 1934 4779 1940 4780
rect 1934 4775 1935 4779
rect 1939 4775 1940 4779
rect 110 4774 116 4775
rect 1934 4774 1940 4775
rect 1974 4744 1980 4745
rect 3798 4744 3804 4745
rect 1974 4740 1975 4744
rect 1979 4740 1980 4744
rect 1974 4739 1980 4740
rect 1994 4743 2000 4744
rect 1994 4739 1995 4743
rect 1999 4739 2000 4743
rect 1994 4738 2000 4739
rect 2154 4743 2160 4744
rect 2154 4739 2155 4743
rect 2159 4739 2160 4743
rect 2154 4738 2160 4739
rect 2346 4743 2352 4744
rect 2346 4739 2347 4743
rect 2351 4739 2352 4743
rect 2346 4738 2352 4739
rect 2538 4743 2544 4744
rect 2538 4739 2539 4743
rect 2543 4739 2544 4743
rect 2538 4738 2544 4739
rect 2730 4743 2736 4744
rect 2730 4739 2731 4743
rect 2735 4739 2736 4743
rect 2730 4738 2736 4739
rect 2930 4743 2936 4744
rect 2930 4739 2931 4743
rect 2935 4739 2936 4743
rect 2930 4738 2936 4739
rect 3130 4743 3136 4744
rect 3130 4739 3131 4743
rect 3135 4739 3136 4743
rect 3798 4740 3799 4744
rect 3803 4740 3804 4744
rect 3798 4739 3804 4740
rect 3130 4738 3136 4739
rect 2022 4728 2028 4729
rect 1974 4727 1980 4728
rect 1974 4723 1975 4727
rect 1979 4723 1980 4727
rect 2022 4724 2023 4728
rect 2027 4724 2028 4728
rect 2022 4723 2028 4724
rect 2182 4728 2188 4729
rect 2182 4724 2183 4728
rect 2187 4724 2188 4728
rect 2182 4723 2188 4724
rect 2374 4728 2380 4729
rect 2374 4724 2375 4728
rect 2379 4724 2380 4728
rect 2374 4723 2380 4724
rect 2566 4728 2572 4729
rect 2566 4724 2567 4728
rect 2571 4724 2572 4728
rect 2566 4723 2572 4724
rect 2758 4728 2764 4729
rect 2758 4724 2759 4728
rect 2763 4724 2764 4728
rect 2758 4723 2764 4724
rect 2958 4728 2964 4729
rect 2958 4724 2959 4728
rect 2963 4724 2964 4728
rect 2958 4723 2964 4724
rect 3158 4728 3164 4729
rect 3158 4724 3159 4728
rect 3163 4724 3164 4728
rect 3158 4723 3164 4724
rect 3798 4727 3804 4728
rect 3798 4723 3799 4727
rect 3803 4723 3804 4727
rect 1974 4722 1980 4723
rect 3798 4722 3804 4723
rect 110 4713 116 4714
rect 1934 4713 1940 4714
rect 110 4709 111 4713
rect 115 4709 116 4713
rect 110 4708 116 4709
rect 158 4712 164 4713
rect 158 4708 159 4712
rect 163 4708 164 4712
rect 158 4707 164 4708
rect 342 4712 348 4713
rect 342 4708 343 4712
rect 347 4708 348 4712
rect 342 4707 348 4708
rect 566 4712 572 4713
rect 566 4708 567 4712
rect 571 4708 572 4712
rect 566 4707 572 4708
rect 806 4712 812 4713
rect 806 4708 807 4712
rect 811 4708 812 4712
rect 806 4707 812 4708
rect 1054 4712 1060 4713
rect 1054 4708 1055 4712
rect 1059 4708 1060 4712
rect 1054 4707 1060 4708
rect 1310 4712 1316 4713
rect 1310 4708 1311 4712
rect 1315 4708 1316 4712
rect 1310 4707 1316 4708
rect 1574 4712 1580 4713
rect 1574 4708 1575 4712
rect 1579 4708 1580 4712
rect 1574 4707 1580 4708
rect 1814 4712 1820 4713
rect 1814 4708 1815 4712
rect 1819 4708 1820 4712
rect 1934 4709 1935 4713
rect 1939 4709 1940 4713
rect 1934 4708 1940 4709
rect 1814 4707 1820 4708
rect 3838 4704 3844 4705
rect 5662 4704 5668 4705
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 3838 4699 3844 4700
rect 3914 4703 3920 4704
rect 3914 4699 3915 4703
rect 3919 4699 3920 4703
rect 3914 4698 3920 4699
rect 4186 4703 4192 4704
rect 4186 4699 4187 4703
rect 4191 4699 4192 4703
rect 4186 4698 4192 4699
rect 4466 4703 4472 4704
rect 4466 4699 4467 4703
rect 4471 4699 4472 4703
rect 4466 4698 4472 4699
rect 4762 4703 4768 4704
rect 4762 4699 4763 4703
rect 4767 4699 4768 4703
rect 4762 4698 4768 4699
rect 5066 4703 5072 4704
rect 5066 4699 5067 4703
rect 5071 4699 5072 4703
rect 5066 4698 5072 4699
rect 5370 4703 5376 4704
rect 5370 4699 5371 4703
rect 5375 4699 5376 4703
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 5662 4699 5668 4700
rect 5370 4698 5376 4699
rect 130 4697 136 4698
rect 110 4696 116 4697
rect 110 4692 111 4696
rect 115 4692 116 4696
rect 130 4693 131 4697
rect 135 4693 136 4697
rect 130 4692 136 4693
rect 314 4697 320 4698
rect 314 4693 315 4697
rect 319 4693 320 4697
rect 314 4692 320 4693
rect 538 4697 544 4698
rect 538 4693 539 4697
rect 543 4693 544 4697
rect 538 4692 544 4693
rect 778 4697 784 4698
rect 778 4693 779 4697
rect 783 4693 784 4697
rect 778 4692 784 4693
rect 1026 4697 1032 4698
rect 1026 4693 1027 4697
rect 1031 4693 1032 4697
rect 1026 4692 1032 4693
rect 1282 4697 1288 4698
rect 1282 4693 1283 4697
rect 1287 4693 1288 4697
rect 1282 4692 1288 4693
rect 1546 4697 1552 4698
rect 1546 4693 1547 4697
rect 1551 4693 1552 4697
rect 1546 4692 1552 4693
rect 1786 4697 1792 4698
rect 1786 4693 1787 4697
rect 1791 4693 1792 4697
rect 1786 4692 1792 4693
rect 1934 4696 1940 4697
rect 1934 4692 1935 4696
rect 1939 4692 1940 4696
rect 110 4691 116 4692
rect 1934 4691 1940 4692
rect 3942 4688 3948 4689
rect 3838 4687 3844 4688
rect 3838 4683 3839 4687
rect 3843 4683 3844 4687
rect 3942 4684 3943 4688
rect 3947 4684 3948 4688
rect 3942 4683 3948 4684
rect 4214 4688 4220 4689
rect 4214 4684 4215 4688
rect 4219 4684 4220 4688
rect 4214 4683 4220 4684
rect 4494 4688 4500 4689
rect 4494 4684 4495 4688
rect 4499 4684 4500 4688
rect 4494 4683 4500 4684
rect 4790 4688 4796 4689
rect 4790 4684 4791 4688
rect 4795 4684 4796 4688
rect 4790 4683 4796 4684
rect 5094 4688 5100 4689
rect 5094 4684 5095 4688
rect 5099 4684 5100 4688
rect 5094 4683 5100 4684
rect 5398 4688 5404 4689
rect 5398 4684 5399 4688
rect 5403 4684 5404 4688
rect 5398 4683 5404 4684
rect 5662 4687 5668 4688
rect 5662 4683 5663 4687
rect 5667 4683 5668 4687
rect 3838 4682 3844 4683
rect 5662 4682 5668 4683
rect 1974 4665 1980 4666
rect 3798 4665 3804 4666
rect 1974 4661 1975 4665
rect 1979 4661 1980 4665
rect 1974 4660 1980 4661
rect 2022 4664 2028 4665
rect 2022 4660 2023 4664
rect 2027 4660 2028 4664
rect 2022 4659 2028 4660
rect 2238 4664 2244 4665
rect 2238 4660 2239 4664
rect 2243 4660 2244 4664
rect 2238 4659 2244 4660
rect 2470 4664 2476 4665
rect 2470 4660 2471 4664
rect 2475 4660 2476 4664
rect 2470 4659 2476 4660
rect 2694 4664 2700 4665
rect 2694 4660 2695 4664
rect 2699 4660 2700 4664
rect 2694 4659 2700 4660
rect 2918 4664 2924 4665
rect 2918 4660 2919 4664
rect 2923 4660 2924 4664
rect 2918 4659 2924 4660
rect 3142 4664 3148 4665
rect 3142 4660 3143 4664
rect 3147 4660 3148 4664
rect 3142 4659 3148 4660
rect 3366 4664 3372 4665
rect 3366 4660 3367 4664
rect 3371 4660 3372 4664
rect 3798 4661 3799 4665
rect 3803 4661 3804 4665
rect 3798 4660 3804 4661
rect 3366 4659 3372 4660
rect 1994 4649 2000 4650
rect 1974 4648 1980 4649
rect 1974 4644 1975 4648
rect 1979 4644 1980 4648
rect 1994 4645 1995 4649
rect 1999 4645 2000 4649
rect 1994 4644 2000 4645
rect 2210 4649 2216 4650
rect 2210 4645 2211 4649
rect 2215 4645 2216 4649
rect 2210 4644 2216 4645
rect 2442 4649 2448 4650
rect 2442 4645 2443 4649
rect 2447 4645 2448 4649
rect 2442 4644 2448 4645
rect 2666 4649 2672 4650
rect 2666 4645 2667 4649
rect 2671 4645 2672 4649
rect 2666 4644 2672 4645
rect 2890 4649 2896 4650
rect 2890 4645 2891 4649
rect 2895 4645 2896 4649
rect 2890 4644 2896 4645
rect 3114 4649 3120 4650
rect 3114 4645 3115 4649
rect 3119 4645 3120 4649
rect 3114 4644 3120 4645
rect 3338 4649 3344 4650
rect 3338 4645 3339 4649
rect 3343 4645 3344 4649
rect 3338 4644 3344 4645
rect 3798 4648 3804 4649
rect 3798 4644 3799 4648
rect 3803 4644 3804 4648
rect 1974 4643 1980 4644
rect 3798 4643 3804 4644
rect 3838 4629 3844 4630
rect 5662 4629 5668 4630
rect 3838 4625 3839 4629
rect 3843 4625 3844 4629
rect 3838 4624 3844 4625
rect 4062 4628 4068 4629
rect 4062 4624 4063 4628
rect 4067 4624 4068 4628
rect 4062 4623 4068 4624
rect 4326 4628 4332 4629
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4326 4623 4332 4624
rect 4598 4628 4604 4629
rect 4598 4624 4599 4628
rect 4603 4624 4604 4628
rect 4598 4623 4604 4624
rect 4870 4628 4876 4629
rect 4870 4624 4871 4628
rect 4875 4624 4876 4628
rect 4870 4623 4876 4624
rect 5150 4628 5156 4629
rect 5150 4624 5151 4628
rect 5155 4624 5156 4628
rect 5150 4623 5156 4624
rect 5438 4628 5444 4629
rect 5438 4624 5439 4628
rect 5443 4624 5444 4628
rect 5662 4625 5663 4629
rect 5667 4625 5668 4629
rect 5662 4624 5668 4625
rect 5438 4623 5444 4624
rect 4034 4613 4040 4614
rect 3838 4612 3844 4613
rect 3838 4608 3839 4612
rect 3843 4608 3844 4612
rect 4034 4609 4035 4613
rect 4039 4609 4040 4613
rect 4034 4608 4040 4609
rect 4298 4613 4304 4614
rect 4298 4609 4299 4613
rect 4303 4609 4304 4613
rect 4298 4608 4304 4609
rect 4570 4613 4576 4614
rect 4570 4609 4571 4613
rect 4575 4609 4576 4613
rect 4570 4608 4576 4609
rect 4842 4613 4848 4614
rect 4842 4609 4843 4613
rect 4847 4609 4848 4613
rect 4842 4608 4848 4609
rect 5122 4613 5128 4614
rect 5122 4609 5123 4613
rect 5127 4609 5128 4613
rect 5122 4608 5128 4609
rect 5410 4613 5416 4614
rect 5410 4609 5411 4613
rect 5415 4609 5416 4613
rect 5410 4608 5416 4609
rect 5662 4612 5668 4613
rect 5662 4608 5663 4612
rect 5667 4608 5668 4612
rect 3838 4607 3844 4608
rect 5662 4607 5668 4608
rect 110 4548 116 4549
rect 1934 4548 1940 4549
rect 110 4544 111 4548
rect 115 4544 116 4548
rect 110 4543 116 4544
rect 170 4547 176 4548
rect 170 4543 171 4547
rect 175 4543 176 4547
rect 170 4542 176 4543
rect 394 4547 400 4548
rect 394 4543 395 4547
rect 399 4543 400 4547
rect 394 4542 400 4543
rect 642 4547 648 4548
rect 642 4543 643 4547
rect 647 4543 648 4547
rect 642 4542 648 4543
rect 906 4547 912 4548
rect 906 4543 907 4547
rect 911 4543 912 4547
rect 906 4542 912 4543
rect 1194 4547 1200 4548
rect 1194 4543 1195 4547
rect 1199 4543 1200 4547
rect 1194 4542 1200 4543
rect 1490 4547 1496 4548
rect 1490 4543 1491 4547
rect 1495 4543 1496 4547
rect 1490 4542 1496 4543
rect 1786 4547 1792 4548
rect 1786 4543 1787 4547
rect 1791 4543 1792 4547
rect 1934 4544 1935 4548
rect 1939 4544 1940 4548
rect 1934 4543 1940 4544
rect 1786 4542 1792 4543
rect 198 4532 204 4533
rect 110 4531 116 4532
rect 110 4527 111 4531
rect 115 4527 116 4531
rect 198 4528 199 4532
rect 203 4528 204 4532
rect 198 4527 204 4528
rect 422 4532 428 4533
rect 422 4528 423 4532
rect 427 4528 428 4532
rect 422 4527 428 4528
rect 670 4532 676 4533
rect 670 4528 671 4532
rect 675 4528 676 4532
rect 670 4527 676 4528
rect 934 4532 940 4533
rect 934 4528 935 4532
rect 939 4528 940 4532
rect 934 4527 940 4528
rect 1222 4532 1228 4533
rect 1222 4528 1223 4532
rect 1227 4528 1228 4532
rect 1222 4527 1228 4528
rect 1518 4532 1524 4533
rect 1518 4528 1519 4532
rect 1523 4528 1524 4532
rect 1518 4527 1524 4528
rect 1814 4532 1820 4533
rect 1814 4528 1815 4532
rect 1819 4528 1820 4532
rect 1814 4527 1820 4528
rect 1934 4531 1940 4532
rect 1934 4527 1935 4531
rect 1939 4527 1940 4531
rect 110 4526 116 4527
rect 1934 4526 1940 4527
rect 1974 4512 1980 4513
rect 3798 4512 3804 4513
rect 1974 4508 1975 4512
rect 1979 4508 1980 4512
rect 1974 4507 1980 4508
rect 2098 4511 2104 4512
rect 2098 4507 2099 4511
rect 2103 4507 2104 4511
rect 2098 4506 2104 4507
rect 2346 4511 2352 4512
rect 2346 4507 2347 4511
rect 2351 4507 2352 4511
rect 2346 4506 2352 4507
rect 2578 4511 2584 4512
rect 2578 4507 2579 4511
rect 2583 4507 2584 4511
rect 2578 4506 2584 4507
rect 2794 4511 2800 4512
rect 2794 4507 2795 4511
rect 2799 4507 2800 4511
rect 2794 4506 2800 4507
rect 3002 4511 3008 4512
rect 3002 4507 3003 4511
rect 3007 4507 3008 4511
rect 3002 4506 3008 4507
rect 3202 4511 3208 4512
rect 3202 4507 3203 4511
rect 3207 4507 3208 4511
rect 3202 4506 3208 4507
rect 3402 4511 3408 4512
rect 3402 4507 3403 4511
rect 3407 4507 3408 4511
rect 3402 4506 3408 4507
rect 3610 4511 3616 4512
rect 3610 4507 3611 4511
rect 3615 4507 3616 4511
rect 3798 4508 3799 4512
rect 3803 4508 3804 4512
rect 3798 4507 3804 4508
rect 3610 4506 3616 4507
rect 2126 4496 2132 4497
rect 1974 4495 1980 4496
rect 1974 4491 1975 4495
rect 1979 4491 1980 4495
rect 2126 4492 2127 4496
rect 2131 4492 2132 4496
rect 2126 4491 2132 4492
rect 2374 4496 2380 4497
rect 2374 4492 2375 4496
rect 2379 4492 2380 4496
rect 2374 4491 2380 4492
rect 2606 4496 2612 4497
rect 2606 4492 2607 4496
rect 2611 4492 2612 4496
rect 2606 4491 2612 4492
rect 2822 4496 2828 4497
rect 2822 4492 2823 4496
rect 2827 4492 2828 4496
rect 2822 4491 2828 4492
rect 3030 4496 3036 4497
rect 3030 4492 3031 4496
rect 3035 4492 3036 4496
rect 3030 4491 3036 4492
rect 3230 4496 3236 4497
rect 3230 4492 3231 4496
rect 3235 4492 3236 4496
rect 3230 4491 3236 4492
rect 3430 4496 3436 4497
rect 3430 4492 3431 4496
rect 3435 4492 3436 4496
rect 3430 4491 3436 4492
rect 3638 4496 3644 4497
rect 3638 4492 3639 4496
rect 3643 4492 3644 4496
rect 3638 4491 3644 4492
rect 3798 4495 3804 4496
rect 3798 4491 3799 4495
rect 3803 4491 3804 4495
rect 1974 4490 1980 4491
rect 3798 4490 3804 4491
rect 3838 4480 3844 4481
rect 5662 4480 5668 4481
rect 3838 4476 3839 4480
rect 3843 4476 3844 4480
rect 3838 4475 3844 4476
rect 4178 4479 4184 4480
rect 4178 4475 4179 4479
rect 4183 4475 4184 4479
rect 4178 4474 4184 4475
rect 4410 4479 4416 4480
rect 4410 4475 4411 4479
rect 4415 4475 4416 4479
rect 4410 4474 4416 4475
rect 4658 4479 4664 4480
rect 4658 4475 4659 4479
rect 4663 4475 4664 4479
rect 4658 4474 4664 4475
rect 4914 4479 4920 4480
rect 4914 4475 4915 4479
rect 4919 4475 4920 4479
rect 4914 4474 4920 4475
rect 5178 4479 5184 4480
rect 5178 4475 5179 4479
rect 5183 4475 5184 4479
rect 5178 4474 5184 4475
rect 5442 4479 5448 4480
rect 5442 4475 5443 4479
rect 5447 4475 5448 4479
rect 5662 4476 5663 4480
rect 5667 4476 5668 4480
rect 5662 4475 5668 4476
rect 5442 4474 5448 4475
rect 110 4469 116 4470
rect 1934 4469 1940 4470
rect 110 4465 111 4469
rect 115 4465 116 4469
rect 110 4464 116 4465
rect 446 4468 452 4469
rect 446 4464 447 4468
rect 451 4464 452 4468
rect 446 4463 452 4464
rect 654 4468 660 4469
rect 654 4464 655 4468
rect 659 4464 660 4468
rect 654 4463 660 4464
rect 886 4468 892 4469
rect 886 4464 887 4468
rect 891 4464 892 4468
rect 886 4463 892 4464
rect 1142 4468 1148 4469
rect 1142 4464 1143 4468
rect 1147 4464 1148 4468
rect 1142 4463 1148 4464
rect 1406 4468 1412 4469
rect 1406 4464 1407 4468
rect 1411 4464 1412 4468
rect 1406 4463 1412 4464
rect 1678 4468 1684 4469
rect 1678 4464 1679 4468
rect 1683 4464 1684 4468
rect 1934 4465 1935 4469
rect 1939 4465 1940 4469
rect 1934 4464 1940 4465
rect 4206 4464 4212 4465
rect 1678 4463 1684 4464
rect 3838 4463 3844 4464
rect 3838 4459 3839 4463
rect 3843 4459 3844 4463
rect 4206 4460 4207 4464
rect 4211 4460 4212 4464
rect 4206 4459 4212 4460
rect 4438 4464 4444 4465
rect 4438 4460 4439 4464
rect 4443 4460 4444 4464
rect 4438 4459 4444 4460
rect 4686 4464 4692 4465
rect 4686 4460 4687 4464
rect 4691 4460 4692 4464
rect 4686 4459 4692 4460
rect 4942 4464 4948 4465
rect 4942 4460 4943 4464
rect 4947 4460 4948 4464
rect 4942 4459 4948 4460
rect 5206 4464 5212 4465
rect 5206 4460 5207 4464
rect 5211 4460 5212 4464
rect 5206 4459 5212 4460
rect 5470 4464 5476 4465
rect 5470 4460 5471 4464
rect 5475 4460 5476 4464
rect 5470 4459 5476 4460
rect 5662 4463 5668 4464
rect 5662 4459 5663 4463
rect 5667 4459 5668 4463
rect 3838 4458 3844 4459
rect 5662 4458 5668 4459
rect 418 4453 424 4454
rect 110 4452 116 4453
rect 110 4448 111 4452
rect 115 4448 116 4452
rect 418 4449 419 4453
rect 423 4449 424 4453
rect 418 4448 424 4449
rect 626 4453 632 4454
rect 626 4449 627 4453
rect 631 4449 632 4453
rect 626 4448 632 4449
rect 858 4453 864 4454
rect 858 4449 859 4453
rect 863 4449 864 4453
rect 858 4448 864 4449
rect 1114 4453 1120 4454
rect 1114 4449 1115 4453
rect 1119 4449 1120 4453
rect 1114 4448 1120 4449
rect 1378 4453 1384 4454
rect 1378 4449 1379 4453
rect 1383 4449 1384 4453
rect 1378 4448 1384 4449
rect 1650 4453 1656 4454
rect 1650 4449 1651 4453
rect 1655 4449 1656 4453
rect 1650 4448 1656 4449
rect 1934 4452 1940 4453
rect 1934 4448 1935 4452
rect 1939 4448 1940 4452
rect 110 4447 116 4448
rect 1934 4447 1940 4448
rect 1974 4429 1980 4430
rect 3798 4429 3804 4430
rect 1974 4425 1975 4429
rect 1979 4425 1980 4429
rect 1974 4424 1980 4425
rect 2230 4428 2236 4429
rect 2230 4424 2231 4428
rect 2235 4424 2236 4428
rect 2230 4423 2236 4424
rect 2446 4428 2452 4429
rect 2446 4424 2447 4428
rect 2451 4424 2452 4428
rect 2446 4423 2452 4424
rect 2662 4428 2668 4429
rect 2662 4424 2663 4428
rect 2667 4424 2668 4428
rect 2662 4423 2668 4424
rect 2870 4428 2876 4429
rect 2870 4424 2871 4428
rect 2875 4424 2876 4428
rect 2870 4423 2876 4424
rect 3078 4428 3084 4429
rect 3078 4424 3079 4428
rect 3083 4424 3084 4428
rect 3078 4423 3084 4424
rect 3286 4428 3292 4429
rect 3286 4424 3287 4428
rect 3291 4424 3292 4428
rect 3286 4423 3292 4424
rect 3494 4428 3500 4429
rect 3494 4424 3495 4428
rect 3499 4424 3500 4428
rect 3494 4423 3500 4424
rect 3678 4428 3684 4429
rect 3678 4424 3679 4428
rect 3683 4424 3684 4428
rect 3798 4425 3799 4429
rect 3803 4425 3804 4429
rect 3798 4424 3804 4425
rect 3678 4423 3684 4424
rect 2202 4413 2208 4414
rect 1974 4412 1980 4413
rect 1974 4408 1975 4412
rect 1979 4408 1980 4412
rect 2202 4409 2203 4413
rect 2207 4409 2208 4413
rect 2202 4408 2208 4409
rect 2418 4413 2424 4414
rect 2418 4409 2419 4413
rect 2423 4409 2424 4413
rect 2418 4408 2424 4409
rect 2634 4413 2640 4414
rect 2634 4409 2635 4413
rect 2639 4409 2640 4413
rect 2634 4408 2640 4409
rect 2842 4413 2848 4414
rect 2842 4409 2843 4413
rect 2847 4409 2848 4413
rect 2842 4408 2848 4409
rect 3050 4413 3056 4414
rect 3050 4409 3051 4413
rect 3055 4409 3056 4413
rect 3050 4408 3056 4409
rect 3258 4413 3264 4414
rect 3258 4409 3259 4413
rect 3263 4409 3264 4413
rect 3258 4408 3264 4409
rect 3466 4413 3472 4414
rect 3466 4409 3467 4413
rect 3471 4409 3472 4413
rect 3466 4408 3472 4409
rect 3650 4413 3656 4414
rect 3650 4409 3651 4413
rect 3655 4409 3656 4413
rect 3650 4408 3656 4409
rect 3798 4412 3804 4413
rect 3798 4408 3799 4412
rect 3803 4408 3804 4412
rect 1974 4407 1980 4408
rect 3798 4407 3804 4408
rect 3838 4397 3844 4398
rect 5662 4397 5668 4398
rect 3838 4393 3839 4397
rect 3843 4393 3844 4397
rect 3838 4392 3844 4393
rect 4358 4396 4364 4397
rect 4358 4392 4359 4396
rect 4363 4392 4364 4396
rect 4358 4391 4364 4392
rect 4518 4396 4524 4397
rect 4518 4392 4519 4396
rect 4523 4392 4524 4396
rect 4518 4391 4524 4392
rect 4686 4396 4692 4397
rect 4686 4392 4687 4396
rect 4691 4392 4692 4396
rect 4686 4391 4692 4392
rect 4878 4396 4884 4397
rect 4878 4392 4879 4396
rect 4883 4392 4884 4396
rect 4878 4391 4884 4392
rect 5078 4396 5084 4397
rect 5078 4392 5079 4396
rect 5083 4392 5084 4396
rect 5078 4391 5084 4392
rect 5286 4396 5292 4397
rect 5286 4392 5287 4396
rect 5291 4392 5292 4396
rect 5286 4391 5292 4392
rect 5502 4396 5508 4397
rect 5502 4392 5503 4396
rect 5507 4392 5508 4396
rect 5662 4393 5663 4397
rect 5667 4393 5668 4397
rect 5662 4392 5668 4393
rect 5502 4391 5508 4392
rect 4330 4381 4336 4382
rect 3838 4380 3844 4381
rect 3838 4376 3839 4380
rect 3843 4376 3844 4380
rect 4330 4377 4331 4381
rect 4335 4377 4336 4381
rect 4330 4376 4336 4377
rect 4490 4381 4496 4382
rect 4490 4377 4491 4381
rect 4495 4377 4496 4381
rect 4490 4376 4496 4377
rect 4658 4381 4664 4382
rect 4658 4377 4659 4381
rect 4663 4377 4664 4381
rect 4658 4376 4664 4377
rect 4850 4381 4856 4382
rect 4850 4377 4851 4381
rect 4855 4377 4856 4381
rect 4850 4376 4856 4377
rect 5050 4381 5056 4382
rect 5050 4377 5051 4381
rect 5055 4377 5056 4381
rect 5050 4376 5056 4377
rect 5258 4381 5264 4382
rect 5258 4377 5259 4381
rect 5263 4377 5264 4381
rect 5258 4376 5264 4377
rect 5474 4381 5480 4382
rect 5474 4377 5475 4381
rect 5479 4377 5480 4381
rect 5474 4376 5480 4377
rect 5662 4380 5668 4381
rect 5662 4376 5663 4380
rect 5667 4376 5668 4380
rect 3838 4375 3844 4376
rect 5662 4375 5668 4376
rect 110 4316 116 4317
rect 1934 4316 1940 4317
rect 110 4312 111 4316
rect 115 4312 116 4316
rect 110 4311 116 4312
rect 666 4315 672 4316
rect 666 4311 667 4315
rect 671 4311 672 4315
rect 666 4310 672 4311
rect 810 4315 816 4316
rect 810 4311 811 4315
rect 815 4311 816 4315
rect 810 4310 816 4311
rect 962 4315 968 4316
rect 962 4311 963 4315
rect 967 4311 968 4315
rect 962 4310 968 4311
rect 1122 4315 1128 4316
rect 1122 4311 1123 4315
rect 1127 4311 1128 4315
rect 1122 4310 1128 4311
rect 1290 4315 1296 4316
rect 1290 4311 1291 4315
rect 1295 4311 1296 4315
rect 1290 4310 1296 4311
rect 1466 4315 1472 4316
rect 1466 4311 1467 4315
rect 1471 4311 1472 4315
rect 1466 4310 1472 4311
rect 1650 4315 1656 4316
rect 1650 4311 1651 4315
rect 1655 4311 1656 4315
rect 1934 4312 1935 4316
rect 1939 4312 1940 4316
rect 1934 4311 1940 4312
rect 1650 4310 1656 4311
rect 694 4300 700 4301
rect 110 4299 116 4300
rect 110 4295 111 4299
rect 115 4295 116 4299
rect 694 4296 695 4300
rect 699 4296 700 4300
rect 694 4295 700 4296
rect 838 4300 844 4301
rect 838 4296 839 4300
rect 843 4296 844 4300
rect 838 4295 844 4296
rect 990 4300 996 4301
rect 990 4296 991 4300
rect 995 4296 996 4300
rect 990 4295 996 4296
rect 1150 4300 1156 4301
rect 1150 4296 1151 4300
rect 1155 4296 1156 4300
rect 1150 4295 1156 4296
rect 1318 4300 1324 4301
rect 1318 4296 1319 4300
rect 1323 4296 1324 4300
rect 1318 4295 1324 4296
rect 1494 4300 1500 4301
rect 1494 4296 1495 4300
rect 1499 4296 1500 4300
rect 1494 4295 1500 4296
rect 1678 4300 1684 4301
rect 1678 4296 1679 4300
rect 1683 4296 1684 4300
rect 1678 4295 1684 4296
rect 1934 4299 1940 4300
rect 1934 4295 1935 4299
rect 1939 4295 1940 4299
rect 110 4294 116 4295
rect 1934 4294 1940 4295
rect 1974 4272 1980 4273
rect 3798 4272 3804 4273
rect 1974 4268 1975 4272
rect 1979 4268 1980 4272
rect 1974 4267 1980 4268
rect 2306 4271 2312 4272
rect 2306 4267 2307 4271
rect 2311 4267 2312 4271
rect 2306 4266 2312 4267
rect 2458 4271 2464 4272
rect 2458 4267 2459 4271
rect 2463 4267 2464 4271
rect 2458 4266 2464 4267
rect 2626 4271 2632 4272
rect 2626 4267 2627 4271
rect 2631 4267 2632 4271
rect 2626 4266 2632 4267
rect 2810 4271 2816 4272
rect 2810 4267 2811 4271
rect 2815 4267 2816 4271
rect 2810 4266 2816 4267
rect 3010 4271 3016 4272
rect 3010 4267 3011 4271
rect 3015 4267 3016 4271
rect 3010 4266 3016 4267
rect 3226 4271 3232 4272
rect 3226 4267 3227 4271
rect 3231 4267 3232 4271
rect 3226 4266 3232 4267
rect 3450 4271 3456 4272
rect 3450 4267 3451 4271
rect 3455 4267 3456 4271
rect 3450 4266 3456 4267
rect 3650 4271 3656 4272
rect 3650 4267 3651 4271
rect 3655 4267 3656 4271
rect 3798 4268 3799 4272
rect 3803 4268 3804 4272
rect 3798 4267 3804 4268
rect 3650 4266 3656 4267
rect 2334 4256 2340 4257
rect 1974 4255 1980 4256
rect 1974 4251 1975 4255
rect 1979 4251 1980 4255
rect 2334 4252 2335 4256
rect 2339 4252 2340 4256
rect 2334 4251 2340 4252
rect 2486 4256 2492 4257
rect 2486 4252 2487 4256
rect 2491 4252 2492 4256
rect 2486 4251 2492 4252
rect 2654 4256 2660 4257
rect 2654 4252 2655 4256
rect 2659 4252 2660 4256
rect 2654 4251 2660 4252
rect 2838 4256 2844 4257
rect 2838 4252 2839 4256
rect 2843 4252 2844 4256
rect 2838 4251 2844 4252
rect 3038 4256 3044 4257
rect 3038 4252 3039 4256
rect 3043 4252 3044 4256
rect 3038 4251 3044 4252
rect 3254 4256 3260 4257
rect 3254 4252 3255 4256
rect 3259 4252 3260 4256
rect 3254 4251 3260 4252
rect 3478 4256 3484 4257
rect 3478 4252 3479 4256
rect 3483 4252 3484 4256
rect 3478 4251 3484 4252
rect 3678 4256 3684 4257
rect 3678 4252 3679 4256
rect 3683 4252 3684 4256
rect 3678 4251 3684 4252
rect 3798 4255 3804 4256
rect 3798 4251 3799 4255
rect 3803 4251 3804 4255
rect 1974 4250 1980 4251
rect 3798 4250 3804 4251
rect 3838 4248 3844 4249
rect 5662 4248 5668 4249
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 3838 4243 3844 4244
rect 3858 4247 3864 4248
rect 3858 4243 3859 4247
rect 3863 4243 3864 4247
rect 3858 4242 3864 4243
rect 4042 4247 4048 4248
rect 4042 4243 4043 4247
rect 4047 4243 4048 4247
rect 4042 4242 4048 4243
rect 4250 4247 4256 4248
rect 4250 4243 4251 4247
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4474 4247 4480 4248
rect 4474 4243 4475 4247
rect 4479 4243 4480 4247
rect 4474 4242 4480 4243
rect 4714 4247 4720 4248
rect 4714 4243 4715 4247
rect 4719 4243 4720 4247
rect 4714 4242 4720 4243
rect 4970 4247 4976 4248
rect 4970 4243 4971 4247
rect 4975 4243 4976 4247
rect 4970 4242 4976 4243
rect 5234 4247 5240 4248
rect 5234 4243 5235 4247
rect 5239 4243 5240 4247
rect 5234 4242 5240 4243
rect 5498 4247 5504 4248
rect 5498 4243 5499 4247
rect 5503 4243 5504 4247
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 5662 4243 5668 4244
rect 5498 4242 5504 4243
rect 3886 4232 3892 4233
rect 3838 4231 3844 4232
rect 3838 4227 3839 4231
rect 3843 4227 3844 4231
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 3886 4227 3892 4228
rect 4070 4232 4076 4233
rect 4070 4228 4071 4232
rect 4075 4228 4076 4232
rect 4070 4227 4076 4228
rect 4278 4232 4284 4233
rect 4278 4228 4279 4232
rect 4283 4228 4284 4232
rect 4278 4227 4284 4228
rect 4502 4232 4508 4233
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4742 4232 4748 4233
rect 4742 4228 4743 4232
rect 4747 4228 4748 4232
rect 4742 4227 4748 4228
rect 4998 4232 5004 4233
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5262 4232 5268 4233
rect 5262 4228 5263 4232
rect 5267 4228 5268 4232
rect 5262 4227 5268 4228
rect 5526 4232 5532 4233
rect 5526 4228 5527 4232
rect 5531 4228 5532 4232
rect 5526 4227 5532 4228
rect 5662 4231 5668 4232
rect 5662 4227 5663 4231
rect 5667 4227 5668 4231
rect 3838 4226 3844 4227
rect 5662 4226 5668 4227
rect 110 4225 116 4226
rect 1934 4225 1940 4226
rect 110 4221 111 4225
rect 115 4221 116 4225
rect 110 4220 116 4221
rect 814 4224 820 4225
rect 814 4220 815 4224
rect 819 4220 820 4224
rect 814 4219 820 4220
rect 950 4224 956 4225
rect 950 4220 951 4224
rect 955 4220 956 4224
rect 950 4219 956 4220
rect 1086 4224 1092 4225
rect 1086 4220 1087 4224
rect 1091 4220 1092 4224
rect 1086 4219 1092 4220
rect 1222 4224 1228 4225
rect 1222 4220 1223 4224
rect 1227 4220 1228 4224
rect 1222 4219 1228 4220
rect 1358 4224 1364 4225
rect 1358 4220 1359 4224
rect 1363 4220 1364 4224
rect 1358 4219 1364 4220
rect 1494 4224 1500 4225
rect 1494 4220 1495 4224
rect 1499 4220 1500 4224
rect 1494 4219 1500 4220
rect 1630 4224 1636 4225
rect 1630 4220 1631 4224
rect 1635 4220 1636 4224
rect 1630 4219 1636 4220
rect 1766 4224 1772 4225
rect 1766 4220 1767 4224
rect 1771 4220 1772 4224
rect 1934 4221 1935 4225
rect 1939 4221 1940 4225
rect 1934 4220 1940 4221
rect 1766 4219 1772 4220
rect 786 4209 792 4210
rect 110 4208 116 4209
rect 110 4204 111 4208
rect 115 4204 116 4208
rect 786 4205 787 4209
rect 791 4205 792 4209
rect 786 4204 792 4205
rect 922 4209 928 4210
rect 922 4205 923 4209
rect 927 4205 928 4209
rect 922 4204 928 4205
rect 1058 4209 1064 4210
rect 1058 4205 1059 4209
rect 1063 4205 1064 4209
rect 1058 4204 1064 4205
rect 1194 4209 1200 4210
rect 1194 4205 1195 4209
rect 1199 4205 1200 4209
rect 1194 4204 1200 4205
rect 1330 4209 1336 4210
rect 1330 4205 1331 4209
rect 1335 4205 1336 4209
rect 1330 4204 1336 4205
rect 1466 4209 1472 4210
rect 1466 4205 1467 4209
rect 1471 4205 1472 4209
rect 1466 4204 1472 4205
rect 1602 4209 1608 4210
rect 1602 4205 1603 4209
rect 1607 4205 1608 4209
rect 1602 4204 1608 4205
rect 1738 4209 1744 4210
rect 1738 4205 1739 4209
rect 1743 4205 1744 4209
rect 1738 4204 1744 4205
rect 1934 4208 1940 4209
rect 1934 4204 1935 4208
rect 1939 4204 1940 4208
rect 110 4203 116 4204
rect 1934 4203 1940 4204
rect 1974 4189 1980 4190
rect 3798 4189 3804 4190
rect 1974 4185 1975 4189
rect 1979 4185 1980 4189
rect 1974 4184 1980 4185
rect 2566 4188 2572 4189
rect 2566 4184 2567 4188
rect 2571 4184 2572 4188
rect 2566 4183 2572 4184
rect 2702 4188 2708 4189
rect 2702 4184 2703 4188
rect 2707 4184 2708 4188
rect 2702 4183 2708 4184
rect 2838 4188 2844 4189
rect 2838 4184 2839 4188
rect 2843 4184 2844 4188
rect 2838 4183 2844 4184
rect 2974 4188 2980 4189
rect 2974 4184 2975 4188
rect 2979 4184 2980 4188
rect 3798 4185 3799 4189
rect 3803 4185 3804 4189
rect 3798 4184 3804 4185
rect 2974 4183 2980 4184
rect 2538 4173 2544 4174
rect 1974 4172 1980 4173
rect 1974 4168 1975 4172
rect 1979 4168 1980 4172
rect 2538 4169 2539 4173
rect 2543 4169 2544 4173
rect 2538 4168 2544 4169
rect 2674 4173 2680 4174
rect 2674 4169 2675 4173
rect 2679 4169 2680 4173
rect 2674 4168 2680 4169
rect 2810 4173 2816 4174
rect 2810 4169 2811 4173
rect 2815 4169 2816 4173
rect 2810 4168 2816 4169
rect 2946 4173 2952 4174
rect 2946 4169 2947 4173
rect 2951 4169 2952 4173
rect 2946 4168 2952 4169
rect 3798 4172 3804 4173
rect 3798 4168 3799 4172
rect 3803 4168 3804 4172
rect 1974 4167 1980 4168
rect 3798 4167 3804 4168
rect 3838 4137 3844 4138
rect 5662 4137 5668 4138
rect 3838 4133 3839 4137
rect 3843 4133 3844 4137
rect 3838 4132 3844 4133
rect 3886 4136 3892 4137
rect 3886 4132 3887 4136
rect 3891 4132 3892 4136
rect 3886 4131 3892 4132
rect 4414 4136 4420 4137
rect 4414 4132 4415 4136
rect 4419 4132 4420 4136
rect 4414 4131 4420 4132
rect 4974 4136 4980 4137
rect 4974 4132 4975 4136
rect 4979 4132 4980 4136
rect 4974 4131 4980 4132
rect 5542 4136 5548 4137
rect 5542 4132 5543 4136
rect 5547 4132 5548 4136
rect 5662 4133 5663 4137
rect 5667 4133 5668 4137
rect 5662 4132 5668 4133
rect 5542 4131 5548 4132
rect 3858 4121 3864 4122
rect 3838 4120 3844 4121
rect 3838 4116 3839 4120
rect 3843 4116 3844 4120
rect 3858 4117 3859 4121
rect 3863 4117 3864 4121
rect 3858 4116 3864 4117
rect 4386 4121 4392 4122
rect 4386 4117 4387 4121
rect 4391 4117 4392 4121
rect 4386 4116 4392 4117
rect 4946 4121 4952 4122
rect 4946 4117 4947 4121
rect 4951 4117 4952 4121
rect 4946 4116 4952 4117
rect 5514 4121 5520 4122
rect 5514 4117 5515 4121
rect 5519 4117 5520 4121
rect 5514 4116 5520 4117
rect 5662 4120 5668 4121
rect 5662 4116 5663 4120
rect 5667 4116 5668 4120
rect 3838 4115 3844 4116
rect 5662 4115 5668 4116
rect 110 4072 116 4073
rect 1934 4072 1940 4073
rect 110 4068 111 4072
rect 115 4068 116 4072
rect 110 4067 116 4068
rect 730 4071 736 4072
rect 730 4067 731 4071
rect 735 4067 736 4071
rect 730 4066 736 4067
rect 866 4071 872 4072
rect 866 4067 867 4071
rect 871 4067 872 4071
rect 866 4066 872 4067
rect 1002 4071 1008 4072
rect 1002 4067 1003 4071
rect 1007 4067 1008 4071
rect 1002 4066 1008 4067
rect 1138 4071 1144 4072
rect 1138 4067 1139 4071
rect 1143 4067 1144 4071
rect 1138 4066 1144 4067
rect 1274 4071 1280 4072
rect 1274 4067 1275 4071
rect 1279 4067 1280 4071
rect 1274 4066 1280 4067
rect 1410 4071 1416 4072
rect 1410 4067 1411 4071
rect 1415 4067 1416 4071
rect 1410 4066 1416 4067
rect 1546 4071 1552 4072
rect 1546 4067 1547 4071
rect 1551 4067 1552 4071
rect 1934 4068 1935 4072
rect 1939 4068 1940 4072
rect 1934 4067 1940 4068
rect 1546 4066 1552 4067
rect 758 4056 764 4057
rect 110 4055 116 4056
rect 110 4051 111 4055
rect 115 4051 116 4055
rect 758 4052 759 4056
rect 763 4052 764 4056
rect 758 4051 764 4052
rect 894 4056 900 4057
rect 894 4052 895 4056
rect 899 4052 900 4056
rect 894 4051 900 4052
rect 1030 4056 1036 4057
rect 1030 4052 1031 4056
rect 1035 4052 1036 4056
rect 1030 4051 1036 4052
rect 1166 4056 1172 4057
rect 1166 4052 1167 4056
rect 1171 4052 1172 4056
rect 1166 4051 1172 4052
rect 1302 4056 1308 4057
rect 1302 4052 1303 4056
rect 1307 4052 1308 4056
rect 1302 4051 1308 4052
rect 1438 4056 1444 4057
rect 1438 4052 1439 4056
rect 1443 4052 1444 4056
rect 1438 4051 1444 4052
rect 1574 4056 1580 4057
rect 1574 4052 1575 4056
rect 1579 4052 1580 4056
rect 1574 4051 1580 4052
rect 1934 4055 1940 4056
rect 1934 4051 1935 4055
rect 1939 4051 1940 4055
rect 110 4050 116 4051
rect 1934 4050 1940 4051
rect 1974 4020 1980 4021
rect 3798 4020 3804 4021
rect 1974 4016 1975 4020
rect 1979 4016 1980 4020
rect 1974 4015 1980 4016
rect 2290 4019 2296 4020
rect 2290 4015 2291 4019
rect 2295 4015 2296 4019
rect 2290 4014 2296 4015
rect 2426 4019 2432 4020
rect 2426 4015 2427 4019
rect 2431 4015 2432 4019
rect 2426 4014 2432 4015
rect 2562 4019 2568 4020
rect 2562 4015 2563 4019
rect 2567 4015 2568 4019
rect 2562 4014 2568 4015
rect 2698 4019 2704 4020
rect 2698 4015 2699 4019
rect 2703 4015 2704 4019
rect 2698 4014 2704 4015
rect 2834 4019 2840 4020
rect 2834 4015 2835 4019
rect 2839 4015 2840 4019
rect 3798 4016 3799 4020
rect 3803 4016 3804 4020
rect 3798 4015 3804 4016
rect 2834 4014 2840 4015
rect 2318 4004 2324 4005
rect 1974 4003 1980 4004
rect 1974 3999 1975 4003
rect 1979 3999 1980 4003
rect 2318 4000 2319 4004
rect 2323 4000 2324 4004
rect 2318 3999 2324 4000
rect 2454 4004 2460 4005
rect 2454 4000 2455 4004
rect 2459 4000 2460 4004
rect 2454 3999 2460 4000
rect 2590 4004 2596 4005
rect 2590 4000 2591 4004
rect 2595 4000 2596 4004
rect 2590 3999 2596 4000
rect 2726 4004 2732 4005
rect 2726 4000 2727 4004
rect 2731 4000 2732 4004
rect 2726 3999 2732 4000
rect 2862 4004 2868 4005
rect 2862 4000 2863 4004
rect 2867 4000 2868 4004
rect 2862 3999 2868 4000
rect 3798 4003 3804 4004
rect 3798 3999 3799 4003
rect 3803 3999 3804 4003
rect 1974 3998 1980 3999
rect 3798 3998 3804 3999
rect 3838 3988 3844 3989
rect 5662 3988 5668 3989
rect 3838 3984 3839 3988
rect 3843 3984 3844 3988
rect 3838 3983 3844 3984
rect 3858 3987 3864 3988
rect 3858 3983 3859 3987
rect 3863 3983 3864 3987
rect 3858 3982 3864 3983
rect 4002 3987 4008 3988
rect 4002 3983 4003 3987
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4170 3987 4176 3988
rect 4170 3983 4171 3987
rect 4175 3983 4176 3987
rect 4170 3982 4176 3983
rect 4338 3987 4344 3988
rect 4338 3983 4339 3987
rect 4343 3983 4344 3987
rect 4338 3982 4344 3983
rect 4498 3987 4504 3988
rect 4498 3983 4499 3987
rect 4503 3983 4504 3987
rect 4498 3982 4504 3983
rect 4650 3987 4656 3988
rect 4650 3983 4651 3987
rect 4655 3983 4656 3987
rect 4650 3982 4656 3983
rect 4802 3987 4808 3988
rect 4802 3983 4803 3987
rect 4807 3983 4808 3987
rect 4802 3982 4808 3983
rect 4946 3987 4952 3988
rect 4946 3983 4947 3987
rect 4951 3983 4952 3987
rect 4946 3982 4952 3983
rect 5090 3987 5096 3988
rect 5090 3983 5091 3987
rect 5095 3983 5096 3987
rect 5090 3982 5096 3983
rect 5234 3987 5240 3988
rect 5234 3983 5235 3987
rect 5239 3983 5240 3987
rect 5234 3982 5240 3983
rect 5378 3987 5384 3988
rect 5378 3983 5379 3987
rect 5383 3983 5384 3987
rect 5378 3982 5384 3983
rect 5514 3987 5520 3988
rect 5514 3983 5515 3987
rect 5519 3983 5520 3987
rect 5662 3984 5663 3988
rect 5667 3984 5668 3988
rect 5662 3983 5668 3984
rect 5514 3982 5520 3983
rect 110 3973 116 3974
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 662 3972 668 3973
rect 662 3968 663 3972
rect 667 3968 668 3972
rect 662 3967 668 3968
rect 822 3972 828 3973
rect 822 3968 823 3972
rect 827 3968 828 3972
rect 822 3967 828 3968
rect 982 3972 988 3973
rect 982 3968 983 3972
rect 987 3968 988 3972
rect 982 3967 988 3968
rect 1150 3972 1156 3973
rect 1150 3968 1151 3972
rect 1155 3968 1156 3972
rect 1150 3967 1156 3968
rect 1318 3972 1324 3973
rect 1318 3968 1319 3972
rect 1323 3968 1324 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 3886 3972 3892 3973
rect 1934 3968 1940 3969
rect 3838 3971 3844 3972
rect 1318 3967 1324 3968
rect 3838 3967 3839 3971
rect 3843 3967 3844 3971
rect 3886 3968 3887 3972
rect 3891 3968 3892 3972
rect 3886 3967 3892 3968
rect 4030 3972 4036 3973
rect 4030 3968 4031 3972
rect 4035 3968 4036 3972
rect 4030 3967 4036 3968
rect 4198 3972 4204 3973
rect 4198 3968 4199 3972
rect 4203 3968 4204 3972
rect 4198 3967 4204 3968
rect 4366 3972 4372 3973
rect 4366 3968 4367 3972
rect 4371 3968 4372 3972
rect 4366 3967 4372 3968
rect 4526 3972 4532 3973
rect 4526 3968 4527 3972
rect 4531 3968 4532 3972
rect 4526 3967 4532 3968
rect 4678 3972 4684 3973
rect 4678 3968 4679 3972
rect 4683 3968 4684 3972
rect 4678 3967 4684 3968
rect 4830 3972 4836 3973
rect 4830 3968 4831 3972
rect 4835 3968 4836 3972
rect 4830 3967 4836 3968
rect 4974 3972 4980 3973
rect 4974 3968 4975 3972
rect 4979 3968 4980 3972
rect 4974 3967 4980 3968
rect 5118 3972 5124 3973
rect 5118 3968 5119 3972
rect 5123 3968 5124 3972
rect 5118 3967 5124 3968
rect 5262 3972 5268 3973
rect 5262 3968 5263 3972
rect 5267 3968 5268 3972
rect 5262 3967 5268 3968
rect 5406 3972 5412 3973
rect 5406 3968 5407 3972
rect 5411 3968 5412 3972
rect 5406 3967 5412 3968
rect 5542 3972 5548 3973
rect 5542 3968 5543 3972
rect 5547 3968 5548 3972
rect 5542 3967 5548 3968
rect 5662 3971 5668 3972
rect 5662 3967 5663 3971
rect 5667 3967 5668 3971
rect 3838 3966 3844 3967
rect 5662 3966 5668 3967
rect 482 3957 488 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 482 3953 483 3957
rect 487 3953 488 3957
rect 482 3952 488 3953
rect 634 3957 640 3958
rect 634 3953 635 3957
rect 639 3953 640 3957
rect 634 3952 640 3953
rect 794 3957 800 3958
rect 794 3953 795 3957
rect 799 3953 800 3957
rect 794 3952 800 3953
rect 954 3957 960 3958
rect 954 3953 955 3957
rect 959 3953 960 3957
rect 954 3952 960 3953
rect 1122 3957 1128 3958
rect 1122 3953 1123 3957
rect 1127 3953 1128 3957
rect 1122 3952 1128 3953
rect 1290 3957 1296 3958
rect 1290 3953 1291 3957
rect 1295 3953 1296 3957
rect 1290 3952 1296 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 1934 3951 1940 3952
rect 1974 3941 1980 3942
rect 3798 3941 3804 3942
rect 1974 3937 1975 3941
rect 1979 3937 1980 3941
rect 1974 3936 1980 3937
rect 2118 3940 2124 3941
rect 2118 3936 2119 3940
rect 2123 3936 2124 3940
rect 2118 3935 2124 3936
rect 2326 3940 2332 3941
rect 2326 3936 2327 3940
rect 2331 3936 2332 3940
rect 2326 3935 2332 3936
rect 2534 3940 2540 3941
rect 2534 3936 2535 3940
rect 2539 3936 2540 3940
rect 2534 3935 2540 3936
rect 2742 3940 2748 3941
rect 2742 3936 2743 3940
rect 2747 3936 2748 3940
rect 2742 3935 2748 3936
rect 2942 3940 2948 3941
rect 2942 3936 2943 3940
rect 2947 3936 2948 3940
rect 2942 3935 2948 3936
rect 3134 3940 3140 3941
rect 3134 3936 3135 3940
rect 3139 3936 3140 3940
rect 3134 3935 3140 3936
rect 3318 3940 3324 3941
rect 3318 3936 3319 3940
rect 3323 3936 3324 3940
rect 3318 3935 3324 3936
rect 3510 3940 3516 3941
rect 3510 3936 3511 3940
rect 3515 3936 3516 3940
rect 3510 3935 3516 3936
rect 3678 3940 3684 3941
rect 3678 3936 3679 3940
rect 3683 3936 3684 3940
rect 3798 3937 3799 3941
rect 3803 3937 3804 3941
rect 3798 3936 3804 3937
rect 3678 3935 3684 3936
rect 2090 3925 2096 3926
rect 1974 3924 1980 3925
rect 1974 3920 1975 3924
rect 1979 3920 1980 3924
rect 2090 3921 2091 3925
rect 2095 3921 2096 3925
rect 2090 3920 2096 3921
rect 2298 3925 2304 3926
rect 2298 3921 2299 3925
rect 2303 3921 2304 3925
rect 2298 3920 2304 3921
rect 2506 3925 2512 3926
rect 2506 3921 2507 3925
rect 2511 3921 2512 3925
rect 2506 3920 2512 3921
rect 2714 3925 2720 3926
rect 2714 3921 2715 3925
rect 2719 3921 2720 3925
rect 2714 3920 2720 3921
rect 2914 3925 2920 3926
rect 2914 3921 2915 3925
rect 2919 3921 2920 3925
rect 2914 3920 2920 3921
rect 3106 3925 3112 3926
rect 3106 3921 3107 3925
rect 3111 3921 3112 3925
rect 3106 3920 3112 3921
rect 3290 3925 3296 3926
rect 3290 3921 3291 3925
rect 3295 3921 3296 3925
rect 3290 3920 3296 3921
rect 3482 3925 3488 3926
rect 3482 3921 3483 3925
rect 3487 3921 3488 3925
rect 3482 3920 3488 3921
rect 3650 3925 3656 3926
rect 3650 3921 3651 3925
rect 3655 3921 3656 3925
rect 3650 3920 3656 3921
rect 3798 3924 3804 3925
rect 3798 3920 3799 3924
rect 3803 3920 3804 3924
rect 1974 3919 1980 3920
rect 3798 3919 3804 3920
rect 3838 3889 3844 3890
rect 5662 3889 5668 3890
rect 3838 3885 3839 3889
rect 3843 3885 3844 3889
rect 3838 3884 3844 3885
rect 4382 3888 4388 3889
rect 4382 3884 4383 3888
rect 4387 3884 4388 3888
rect 4382 3883 4388 3884
rect 4598 3888 4604 3889
rect 4598 3884 4599 3888
rect 4603 3884 4604 3888
rect 4598 3883 4604 3884
rect 4822 3888 4828 3889
rect 4822 3884 4823 3888
rect 4827 3884 4828 3888
rect 4822 3883 4828 3884
rect 5062 3888 5068 3889
rect 5062 3884 5063 3888
rect 5067 3884 5068 3888
rect 5062 3883 5068 3884
rect 5310 3888 5316 3889
rect 5310 3884 5311 3888
rect 5315 3884 5316 3888
rect 5310 3883 5316 3884
rect 5542 3888 5548 3889
rect 5542 3884 5543 3888
rect 5547 3884 5548 3888
rect 5662 3885 5663 3889
rect 5667 3885 5668 3889
rect 5662 3884 5668 3885
rect 5542 3883 5548 3884
rect 4354 3873 4360 3874
rect 3838 3872 3844 3873
rect 3838 3868 3839 3872
rect 3843 3868 3844 3872
rect 4354 3869 4355 3873
rect 4359 3869 4360 3873
rect 4354 3868 4360 3869
rect 4570 3873 4576 3874
rect 4570 3869 4571 3873
rect 4575 3869 4576 3873
rect 4570 3868 4576 3869
rect 4794 3873 4800 3874
rect 4794 3869 4795 3873
rect 4799 3869 4800 3873
rect 4794 3868 4800 3869
rect 5034 3873 5040 3874
rect 5034 3869 5035 3873
rect 5039 3869 5040 3873
rect 5034 3868 5040 3869
rect 5282 3873 5288 3874
rect 5282 3869 5283 3873
rect 5287 3869 5288 3873
rect 5282 3868 5288 3869
rect 5514 3873 5520 3874
rect 5514 3869 5515 3873
rect 5519 3869 5520 3873
rect 5514 3868 5520 3869
rect 5662 3872 5668 3873
rect 5662 3868 5663 3872
rect 5667 3868 5668 3872
rect 3838 3867 3844 3868
rect 5662 3867 5668 3868
rect 110 3796 116 3797
rect 1934 3796 1940 3797
rect 110 3792 111 3796
rect 115 3792 116 3796
rect 110 3791 116 3792
rect 130 3795 136 3796
rect 130 3791 131 3795
rect 135 3791 136 3795
rect 130 3790 136 3791
rect 306 3795 312 3796
rect 306 3791 307 3795
rect 311 3791 312 3795
rect 306 3790 312 3791
rect 514 3795 520 3796
rect 514 3791 515 3795
rect 519 3791 520 3795
rect 514 3790 520 3791
rect 722 3795 728 3796
rect 722 3791 723 3795
rect 727 3791 728 3795
rect 722 3790 728 3791
rect 938 3795 944 3796
rect 938 3791 939 3795
rect 943 3791 944 3795
rect 938 3790 944 3791
rect 1162 3795 1168 3796
rect 1162 3791 1163 3795
rect 1167 3791 1168 3795
rect 1934 3792 1935 3796
rect 1939 3792 1940 3796
rect 1934 3791 1940 3792
rect 1162 3790 1168 3791
rect 158 3780 164 3781
rect 110 3779 116 3780
rect 110 3775 111 3779
rect 115 3775 116 3779
rect 158 3776 159 3780
rect 163 3776 164 3780
rect 158 3775 164 3776
rect 334 3780 340 3781
rect 334 3776 335 3780
rect 339 3776 340 3780
rect 334 3775 340 3776
rect 542 3780 548 3781
rect 542 3776 543 3780
rect 547 3776 548 3780
rect 542 3775 548 3776
rect 750 3780 756 3781
rect 750 3776 751 3780
rect 755 3776 756 3780
rect 750 3775 756 3776
rect 966 3780 972 3781
rect 966 3776 967 3780
rect 971 3776 972 3780
rect 966 3775 972 3776
rect 1190 3780 1196 3781
rect 1974 3780 1980 3781
rect 3798 3780 3804 3781
rect 1190 3776 1191 3780
rect 1195 3776 1196 3780
rect 1190 3775 1196 3776
rect 1934 3779 1940 3780
rect 1934 3775 1935 3779
rect 1939 3775 1940 3779
rect 1974 3776 1975 3780
rect 1979 3776 1980 3780
rect 1974 3775 1980 3776
rect 2138 3779 2144 3780
rect 2138 3775 2139 3779
rect 2143 3775 2144 3779
rect 110 3774 116 3775
rect 1934 3774 1940 3775
rect 2138 3774 2144 3775
rect 2370 3779 2376 3780
rect 2370 3775 2371 3779
rect 2375 3775 2376 3779
rect 2370 3774 2376 3775
rect 2586 3779 2592 3780
rect 2586 3775 2587 3779
rect 2591 3775 2592 3779
rect 2586 3774 2592 3775
rect 2794 3779 2800 3780
rect 2794 3775 2795 3779
rect 2799 3775 2800 3779
rect 2794 3774 2800 3775
rect 2994 3779 3000 3780
rect 2994 3775 2995 3779
rect 2999 3775 3000 3779
rect 2994 3774 3000 3775
rect 3194 3779 3200 3780
rect 3194 3775 3195 3779
rect 3199 3775 3200 3779
rect 3194 3774 3200 3775
rect 3402 3779 3408 3780
rect 3402 3775 3403 3779
rect 3407 3775 3408 3779
rect 3798 3776 3799 3780
rect 3803 3776 3804 3780
rect 3798 3775 3804 3776
rect 3402 3774 3408 3775
rect 2166 3764 2172 3765
rect 1974 3763 1980 3764
rect 1974 3759 1975 3763
rect 1979 3759 1980 3763
rect 2166 3760 2167 3764
rect 2171 3760 2172 3764
rect 2166 3759 2172 3760
rect 2398 3764 2404 3765
rect 2398 3760 2399 3764
rect 2403 3760 2404 3764
rect 2398 3759 2404 3760
rect 2614 3764 2620 3765
rect 2614 3760 2615 3764
rect 2619 3760 2620 3764
rect 2614 3759 2620 3760
rect 2822 3764 2828 3765
rect 2822 3760 2823 3764
rect 2827 3760 2828 3764
rect 2822 3759 2828 3760
rect 3022 3764 3028 3765
rect 3022 3760 3023 3764
rect 3027 3760 3028 3764
rect 3022 3759 3028 3760
rect 3222 3764 3228 3765
rect 3222 3760 3223 3764
rect 3227 3760 3228 3764
rect 3222 3759 3228 3760
rect 3430 3764 3436 3765
rect 3430 3760 3431 3764
rect 3435 3760 3436 3764
rect 3430 3759 3436 3760
rect 3798 3763 3804 3764
rect 3798 3759 3799 3763
rect 3803 3759 3804 3763
rect 1974 3758 1980 3759
rect 3798 3758 3804 3759
rect 3838 3724 3844 3725
rect 5662 3724 5668 3725
rect 110 3721 116 3722
rect 1934 3721 1940 3722
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 334 3720 340 3721
rect 334 3716 335 3720
rect 339 3716 340 3720
rect 334 3715 340 3716
rect 526 3720 532 3721
rect 526 3716 527 3720
rect 531 3716 532 3720
rect 526 3715 532 3716
rect 710 3720 716 3721
rect 710 3716 711 3720
rect 715 3716 716 3720
rect 710 3715 716 3716
rect 886 3720 892 3721
rect 886 3716 887 3720
rect 891 3716 892 3720
rect 886 3715 892 3716
rect 1054 3720 1060 3721
rect 1054 3716 1055 3720
rect 1059 3716 1060 3720
rect 1054 3715 1060 3716
rect 1214 3720 1220 3721
rect 1214 3716 1215 3720
rect 1219 3716 1220 3720
rect 1214 3715 1220 3716
rect 1366 3720 1372 3721
rect 1366 3716 1367 3720
rect 1371 3716 1372 3720
rect 1366 3715 1372 3716
rect 1518 3720 1524 3721
rect 1518 3716 1519 3720
rect 1523 3716 1524 3720
rect 1518 3715 1524 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1678 3715 1684 3716
rect 1814 3720 1820 3721
rect 1814 3716 1815 3720
rect 1819 3716 1820 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 3838 3720 3839 3724
rect 3843 3720 3844 3724
rect 3838 3719 3844 3720
rect 3994 3723 4000 3724
rect 3994 3719 3995 3723
rect 3999 3719 4000 3723
rect 3994 3718 4000 3719
rect 4202 3723 4208 3724
rect 4202 3719 4203 3723
rect 4207 3719 4208 3723
rect 4202 3718 4208 3719
rect 4434 3723 4440 3724
rect 4434 3719 4435 3723
rect 4439 3719 4440 3723
rect 4434 3718 4440 3719
rect 4690 3723 4696 3724
rect 4690 3719 4691 3723
rect 4695 3719 4696 3723
rect 4690 3718 4696 3719
rect 4962 3723 4968 3724
rect 4962 3719 4963 3723
rect 4967 3719 4968 3723
rect 4962 3718 4968 3719
rect 5250 3723 5256 3724
rect 5250 3719 5251 3723
rect 5255 3719 5256 3723
rect 5250 3718 5256 3719
rect 5514 3723 5520 3724
rect 5514 3719 5515 3723
rect 5519 3719 5520 3723
rect 5662 3720 5663 3724
rect 5667 3720 5668 3724
rect 5662 3719 5668 3720
rect 5514 3718 5520 3719
rect 1934 3716 1940 3717
rect 1814 3715 1820 3716
rect 4022 3708 4028 3709
rect 3838 3707 3844 3708
rect 130 3705 136 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 130 3701 131 3705
rect 135 3701 136 3705
rect 130 3700 136 3701
rect 306 3705 312 3706
rect 306 3701 307 3705
rect 311 3701 312 3705
rect 306 3700 312 3701
rect 498 3705 504 3706
rect 498 3701 499 3705
rect 503 3701 504 3705
rect 498 3700 504 3701
rect 682 3705 688 3706
rect 682 3701 683 3705
rect 687 3701 688 3705
rect 682 3700 688 3701
rect 858 3705 864 3706
rect 858 3701 859 3705
rect 863 3701 864 3705
rect 858 3700 864 3701
rect 1026 3705 1032 3706
rect 1026 3701 1027 3705
rect 1031 3701 1032 3705
rect 1026 3700 1032 3701
rect 1186 3705 1192 3706
rect 1186 3701 1187 3705
rect 1191 3701 1192 3705
rect 1186 3700 1192 3701
rect 1338 3705 1344 3706
rect 1338 3701 1339 3705
rect 1343 3701 1344 3705
rect 1338 3700 1344 3701
rect 1490 3705 1496 3706
rect 1490 3701 1491 3705
rect 1495 3701 1496 3705
rect 1490 3700 1496 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1786 3705 1792 3706
rect 1786 3701 1787 3705
rect 1791 3701 1792 3705
rect 1786 3700 1792 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 3838 3703 3839 3707
rect 3843 3703 3844 3707
rect 4022 3704 4023 3708
rect 4027 3704 4028 3708
rect 4022 3703 4028 3704
rect 4230 3708 4236 3709
rect 4230 3704 4231 3708
rect 4235 3704 4236 3708
rect 4230 3703 4236 3704
rect 4462 3708 4468 3709
rect 4462 3704 4463 3708
rect 4467 3704 4468 3708
rect 4462 3703 4468 3704
rect 4718 3708 4724 3709
rect 4718 3704 4719 3708
rect 4723 3704 4724 3708
rect 4718 3703 4724 3704
rect 4990 3708 4996 3709
rect 4990 3704 4991 3708
rect 4995 3704 4996 3708
rect 4990 3703 4996 3704
rect 5278 3708 5284 3709
rect 5278 3704 5279 3708
rect 5283 3704 5284 3708
rect 5278 3703 5284 3704
rect 5542 3708 5548 3709
rect 5542 3704 5543 3708
rect 5547 3704 5548 3708
rect 5542 3703 5548 3704
rect 5662 3707 5668 3708
rect 5662 3703 5663 3707
rect 5667 3703 5668 3707
rect 3838 3702 3844 3703
rect 5662 3702 5668 3703
rect 110 3699 116 3700
rect 1934 3699 1940 3700
rect 1974 3701 1980 3702
rect 3798 3701 3804 3702
rect 1974 3697 1975 3701
rect 1979 3697 1980 3701
rect 1974 3696 1980 3697
rect 2278 3700 2284 3701
rect 2278 3696 2279 3700
rect 2283 3696 2284 3700
rect 2278 3695 2284 3696
rect 2478 3700 2484 3701
rect 2478 3696 2479 3700
rect 2483 3696 2484 3700
rect 2478 3695 2484 3696
rect 2678 3700 2684 3701
rect 2678 3696 2679 3700
rect 2683 3696 2684 3700
rect 2678 3695 2684 3696
rect 2878 3700 2884 3701
rect 2878 3696 2879 3700
rect 2883 3696 2884 3700
rect 2878 3695 2884 3696
rect 3078 3700 3084 3701
rect 3078 3696 3079 3700
rect 3083 3696 3084 3700
rect 3078 3695 3084 3696
rect 3278 3700 3284 3701
rect 3278 3696 3279 3700
rect 3283 3696 3284 3700
rect 3798 3697 3799 3701
rect 3803 3697 3804 3701
rect 3798 3696 3804 3697
rect 3278 3695 3284 3696
rect 2250 3685 2256 3686
rect 1974 3684 1980 3685
rect 1974 3680 1975 3684
rect 1979 3680 1980 3684
rect 2250 3681 2251 3685
rect 2255 3681 2256 3685
rect 2250 3680 2256 3681
rect 2450 3685 2456 3686
rect 2450 3681 2451 3685
rect 2455 3681 2456 3685
rect 2450 3680 2456 3681
rect 2650 3685 2656 3686
rect 2650 3681 2651 3685
rect 2655 3681 2656 3685
rect 2650 3680 2656 3681
rect 2850 3685 2856 3686
rect 2850 3681 2851 3685
rect 2855 3681 2856 3685
rect 2850 3680 2856 3681
rect 3050 3685 3056 3686
rect 3050 3681 3051 3685
rect 3055 3681 3056 3685
rect 3050 3680 3056 3681
rect 3250 3685 3256 3686
rect 3250 3681 3251 3685
rect 3255 3681 3256 3685
rect 3250 3680 3256 3681
rect 3798 3684 3804 3685
rect 3798 3680 3799 3684
rect 3803 3680 3804 3684
rect 1974 3679 1980 3680
rect 3798 3679 3804 3680
rect 3838 3621 3844 3622
rect 5662 3621 5668 3622
rect 3838 3617 3839 3621
rect 3843 3617 3844 3621
rect 3838 3616 3844 3617
rect 4214 3620 4220 3621
rect 4214 3616 4215 3620
rect 4219 3616 4220 3620
rect 4214 3615 4220 3616
rect 4398 3620 4404 3621
rect 4398 3616 4399 3620
rect 4403 3616 4404 3620
rect 4398 3615 4404 3616
rect 4606 3620 4612 3621
rect 4606 3616 4607 3620
rect 4611 3616 4612 3620
rect 4606 3615 4612 3616
rect 4830 3620 4836 3621
rect 4830 3616 4831 3620
rect 4835 3616 4836 3620
rect 4830 3615 4836 3616
rect 5070 3620 5076 3621
rect 5070 3616 5071 3620
rect 5075 3616 5076 3620
rect 5070 3615 5076 3616
rect 5318 3620 5324 3621
rect 5318 3616 5319 3620
rect 5323 3616 5324 3620
rect 5318 3615 5324 3616
rect 5542 3620 5548 3621
rect 5542 3616 5543 3620
rect 5547 3616 5548 3620
rect 5662 3617 5663 3621
rect 5667 3617 5668 3621
rect 5662 3616 5668 3617
rect 5542 3615 5548 3616
rect 4186 3605 4192 3606
rect 3838 3604 3844 3605
rect 3838 3600 3839 3604
rect 3843 3600 3844 3604
rect 4186 3601 4187 3605
rect 4191 3601 4192 3605
rect 4186 3600 4192 3601
rect 4370 3605 4376 3606
rect 4370 3601 4371 3605
rect 4375 3601 4376 3605
rect 4370 3600 4376 3601
rect 4578 3605 4584 3606
rect 4578 3601 4579 3605
rect 4583 3601 4584 3605
rect 4578 3600 4584 3601
rect 4802 3605 4808 3606
rect 4802 3601 4803 3605
rect 4807 3601 4808 3605
rect 4802 3600 4808 3601
rect 5042 3605 5048 3606
rect 5042 3601 5043 3605
rect 5047 3601 5048 3605
rect 5042 3600 5048 3601
rect 5290 3605 5296 3606
rect 5290 3601 5291 3605
rect 5295 3601 5296 3605
rect 5290 3600 5296 3601
rect 5514 3605 5520 3606
rect 5514 3601 5515 3605
rect 5519 3601 5520 3605
rect 5514 3600 5520 3601
rect 5662 3604 5668 3605
rect 5662 3600 5663 3604
rect 5667 3600 5668 3604
rect 3838 3599 3844 3600
rect 5662 3599 5668 3600
rect 110 3560 116 3561
rect 1934 3560 1940 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 146 3559 152 3560
rect 146 3555 147 3559
rect 151 3555 152 3559
rect 146 3554 152 3555
rect 354 3559 360 3560
rect 354 3555 355 3559
rect 359 3555 360 3559
rect 354 3554 360 3555
rect 570 3559 576 3560
rect 570 3555 571 3559
rect 575 3555 576 3559
rect 570 3554 576 3555
rect 802 3559 808 3560
rect 802 3555 803 3559
rect 807 3555 808 3559
rect 802 3554 808 3555
rect 1042 3559 1048 3560
rect 1042 3555 1043 3559
rect 1047 3555 1048 3559
rect 1042 3554 1048 3555
rect 1290 3559 1296 3560
rect 1290 3555 1291 3559
rect 1295 3555 1296 3559
rect 1290 3554 1296 3555
rect 1546 3559 1552 3560
rect 1546 3555 1547 3559
rect 1551 3555 1552 3559
rect 1546 3554 1552 3555
rect 1786 3559 1792 3560
rect 1786 3555 1787 3559
rect 1791 3555 1792 3559
rect 1934 3556 1935 3560
rect 1939 3556 1940 3560
rect 1934 3555 1940 3556
rect 1786 3554 1792 3555
rect 174 3544 180 3545
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 174 3540 175 3544
rect 179 3540 180 3544
rect 174 3539 180 3540
rect 382 3544 388 3545
rect 382 3540 383 3544
rect 387 3540 388 3544
rect 382 3539 388 3540
rect 598 3544 604 3545
rect 598 3540 599 3544
rect 603 3540 604 3544
rect 598 3539 604 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 1070 3544 1076 3545
rect 1070 3540 1071 3544
rect 1075 3540 1076 3544
rect 1070 3539 1076 3540
rect 1318 3544 1324 3545
rect 1318 3540 1319 3544
rect 1323 3540 1324 3544
rect 1318 3539 1324 3540
rect 1574 3544 1580 3545
rect 1574 3540 1575 3544
rect 1579 3540 1580 3544
rect 1574 3539 1580 3540
rect 1814 3544 1820 3545
rect 1814 3540 1815 3544
rect 1819 3540 1820 3544
rect 1814 3539 1820 3540
rect 1934 3543 1940 3544
rect 1934 3539 1935 3543
rect 1939 3539 1940 3543
rect 110 3538 116 3539
rect 1934 3538 1940 3539
rect 1974 3540 1980 3541
rect 3798 3540 3804 3541
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 1994 3539 2000 3540
rect 1994 3535 1995 3539
rect 1999 3535 2000 3539
rect 1994 3534 2000 3535
rect 2250 3539 2256 3540
rect 2250 3535 2251 3539
rect 2255 3535 2256 3539
rect 2250 3534 2256 3535
rect 2514 3539 2520 3540
rect 2514 3535 2515 3539
rect 2519 3535 2520 3539
rect 2514 3534 2520 3535
rect 2754 3539 2760 3540
rect 2754 3535 2755 3539
rect 2759 3535 2760 3539
rect 2754 3534 2760 3535
rect 2978 3539 2984 3540
rect 2978 3535 2979 3539
rect 2983 3535 2984 3539
rect 2978 3534 2984 3535
rect 3194 3539 3200 3540
rect 3194 3535 3195 3539
rect 3199 3535 3200 3539
rect 3194 3534 3200 3535
rect 3410 3539 3416 3540
rect 3410 3535 3411 3539
rect 3415 3535 3416 3539
rect 3410 3534 3416 3535
rect 3626 3539 3632 3540
rect 3626 3535 3627 3539
rect 3631 3535 3632 3539
rect 3798 3536 3799 3540
rect 3803 3536 3804 3540
rect 3798 3535 3804 3536
rect 3626 3534 3632 3535
rect 2022 3524 2028 3525
rect 1974 3523 1980 3524
rect 1974 3519 1975 3523
rect 1979 3519 1980 3523
rect 2022 3520 2023 3524
rect 2027 3520 2028 3524
rect 2022 3519 2028 3520
rect 2278 3524 2284 3525
rect 2278 3520 2279 3524
rect 2283 3520 2284 3524
rect 2278 3519 2284 3520
rect 2542 3524 2548 3525
rect 2542 3520 2543 3524
rect 2547 3520 2548 3524
rect 2542 3519 2548 3520
rect 2782 3524 2788 3525
rect 2782 3520 2783 3524
rect 2787 3520 2788 3524
rect 2782 3519 2788 3520
rect 3006 3524 3012 3525
rect 3006 3520 3007 3524
rect 3011 3520 3012 3524
rect 3006 3519 3012 3520
rect 3222 3524 3228 3525
rect 3222 3520 3223 3524
rect 3227 3520 3228 3524
rect 3222 3519 3228 3520
rect 3438 3524 3444 3525
rect 3438 3520 3439 3524
rect 3443 3520 3444 3524
rect 3438 3519 3444 3520
rect 3654 3524 3660 3525
rect 3654 3520 3655 3524
rect 3659 3520 3660 3524
rect 3654 3519 3660 3520
rect 3798 3523 3804 3524
rect 3798 3519 3799 3523
rect 3803 3519 3804 3523
rect 1974 3518 1980 3519
rect 3798 3518 3804 3519
rect 110 3461 116 3462
rect 1934 3461 1940 3462
rect 110 3457 111 3461
rect 115 3457 116 3461
rect 110 3456 116 3457
rect 302 3460 308 3461
rect 302 3456 303 3460
rect 307 3456 308 3460
rect 302 3455 308 3456
rect 446 3460 452 3461
rect 446 3456 447 3460
rect 451 3456 452 3460
rect 446 3455 452 3456
rect 598 3460 604 3461
rect 598 3456 599 3460
rect 603 3456 604 3460
rect 598 3455 604 3456
rect 758 3460 764 3461
rect 758 3456 759 3460
rect 763 3456 764 3460
rect 758 3455 764 3456
rect 934 3460 940 3461
rect 934 3456 935 3460
rect 939 3456 940 3460
rect 934 3455 940 3456
rect 1110 3460 1116 3461
rect 1110 3456 1111 3460
rect 1115 3456 1116 3460
rect 1110 3455 1116 3456
rect 1294 3460 1300 3461
rect 1294 3456 1295 3460
rect 1299 3456 1300 3460
rect 1294 3455 1300 3456
rect 1486 3460 1492 3461
rect 1486 3456 1487 3460
rect 1491 3456 1492 3460
rect 1934 3457 1935 3461
rect 1939 3457 1940 3461
rect 1934 3456 1940 3457
rect 1974 3457 1980 3458
rect 3798 3457 3804 3458
rect 1486 3455 1492 3456
rect 1974 3453 1975 3457
rect 1979 3453 1980 3457
rect 1974 3452 1980 3453
rect 2022 3456 2028 3457
rect 2022 3452 2023 3456
rect 2027 3452 2028 3456
rect 2022 3451 2028 3452
rect 2190 3456 2196 3457
rect 2190 3452 2191 3456
rect 2195 3452 2196 3456
rect 2190 3451 2196 3452
rect 2398 3456 2404 3457
rect 2398 3452 2399 3456
rect 2403 3452 2404 3456
rect 2398 3451 2404 3452
rect 2614 3456 2620 3457
rect 2614 3452 2615 3456
rect 2619 3452 2620 3456
rect 2614 3451 2620 3452
rect 2830 3456 2836 3457
rect 2830 3452 2831 3456
rect 2835 3452 2836 3456
rect 2830 3451 2836 3452
rect 3046 3456 3052 3457
rect 3046 3452 3047 3456
rect 3051 3452 3052 3456
rect 3046 3451 3052 3452
rect 3262 3456 3268 3457
rect 3262 3452 3263 3456
rect 3267 3452 3268 3456
rect 3262 3451 3268 3452
rect 3478 3456 3484 3457
rect 3478 3452 3479 3456
rect 3483 3452 3484 3456
rect 3478 3451 3484 3452
rect 3678 3456 3684 3457
rect 3678 3452 3679 3456
rect 3683 3452 3684 3456
rect 3798 3453 3799 3457
rect 3803 3453 3804 3457
rect 3798 3452 3804 3453
rect 3678 3451 3684 3452
rect 3838 3448 3844 3449
rect 5662 3448 5668 3449
rect 274 3445 280 3446
rect 110 3444 116 3445
rect 110 3440 111 3444
rect 115 3440 116 3444
rect 274 3441 275 3445
rect 279 3441 280 3445
rect 274 3440 280 3441
rect 418 3445 424 3446
rect 418 3441 419 3445
rect 423 3441 424 3445
rect 418 3440 424 3441
rect 570 3445 576 3446
rect 570 3441 571 3445
rect 575 3441 576 3445
rect 570 3440 576 3441
rect 730 3445 736 3446
rect 730 3441 731 3445
rect 735 3441 736 3445
rect 730 3440 736 3441
rect 906 3445 912 3446
rect 906 3441 907 3445
rect 911 3441 912 3445
rect 906 3440 912 3441
rect 1082 3445 1088 3446
rect 1082 3441 1083 3445
rect 1087 3441 1088 3445
rect 1082 3440 1088 3441
rect 1266 3445 1272 3446
rect 1266 3441 1267 3445
rect 1271 3441 1272 3445
rect 1266 3440 1272 3441
rect 1458 3445 1464 3446
rect 1458 3441 1459 3445
rect 1463 3441 1464 3445
rect 1458 3440 1464 3441
rect 1934 3444 1940 3445
rect 1934 3440 1935 3444
rect 1939 3440 1940 3444
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3838 3443 3844 3444
rect 4530 3447 4536 3448
rect 4530 3443 4531 3447
rect 4535 3443 4536 3447
rect 4530 3442 4536 3443
rect 4682 3447 4688 3448
rect 4682 3443 4683 3447
rect 4687 3443 4688 3447
rect 4682 3442 4688 3443
rect 4842 3447 4848 3448
rect 4842 3443 4843 3447
rect 4847 3443 4848 3447
rect 4842 3442 4848 3443
rect 5002 3447 5008 3448
rect 5002 3443 5003 3447
rect 5007 3443 5008 3447
rect 5002 3442 5008 3443
rect 5170 3447 5176 3448
rect 5170 3443 5171 3447
rect 5175 3443 5176 3447
rect 5170 3442 5176 3443
rect 5346 3447 5352 3448
rect 5346 3443 5347 3447
rect 5351 3443 5352 3447
rect 5346 3442 5352 3443
rect 5514 3447 5520 3448
rect 5514 3443 5515 3447
rect 5519 3443 5520 3447
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 5662 3443 5668 3444
rect 5514 3442 5520 3443
rect 1994 3441 2000 3442
rect 110 3439 116 3440
rect 1934 3439 1940 3440
rect 1974 3440 1980 3441
rect 1974 3436 1975 3440
rect 1979 3436 1980 3440
rect 1994 3437 1995 3441
rect 1999 3437 2000 3441
rect 1994 3436 2000 3437
rect 2162 3441 2168 3442
rect 2162 3437 2163 3441
rect 2167 3437 2168 3441
rect 2162 3436 2168 3437
rect 2370 3441 2376 3442
rect 2370 3437 2371 3441
rect 2375 3437 2376 3441
rect 2370 3436 2376 3437
rect 2586 3441 2592 3442
rect 2586 3437 2587 3441
rect 2591 3437 2592 3441
rect 2586 3436 2592 3437
rect 2802 3441 2808 3442
rect 2802 3437 2803 3441
rect 2807 3437 2808 3441
rect 2802 3436 2808 3437
rect 3018 3441 3024 3442
rect 3018 3437 3019 3441
rect 3023 3437 3024 3441
rect 3018 3436 3024 3437
rect 3234 3441 3240 3442
rect 3234 3437 3235 3441
rect 3239 3437 3240 3441
rect 3234 3436 3240 3437
rect 3450 3441 3456 3442
rect 3450 3437 3451 3441
rect 3455 3437 3456 3441
rect 3450 3436 3456 3437
rect 3650 3441 3656 3442
rect 3650 3437 3651 3441
rect 3655 3437 3656 3441
rect 3650 3436 3656 3437
rect 3798 3440 3804 3441
rect 3798 3436 3799 3440
rect 3803 3436 3804 3440
rect 1974 3435 1980 3436
rect 3798 3435 3804 3436
rect 4558 3432 4564 3433
rect 3838 3431 3844 3432
rect 3838 3427 3839 3431
rect 3843 3427 3844 3431
rect 4558 3428 4559 3432
rect 4563 3428 4564 3432
rect 4558 3427 4564 3428
rect 4710 3432 4716 3433
rect 4710 3428 4711 3432
rect 4715 3428 4716 3432
rect 4710 3427 4716 3428
rect 4870 3432 4876 3433
rect 4870 3428 4871 3432
rect 4875 3428 4876 3432
rect 4870 3427 4876 3428
rect 5030 3432 5036 3433
rect 5030 3428 5031 3432
rect 5035 3428 5036 3432
rect 5030 3427 5036 3428
rect 5198 3432 5204 3433
rect 5198 3428 5199 3432
rect 5203 3428 5204 3432
rect 5198 3427 5204 3428
rect 5374 3432 5380 3433
rect 5374 3428 5375 3432
rect 5379 3428 5380 3432
rect 5374 3427 5380 3428
rect 5542 3432 5548 3433
rect 5542 3428 5543 3432
rect 5547 3428 5548 3432
rect 5542 3427 5548 3428
rect 5662 3431 5668 3432
rect 5662 3427 5663 3431
rect 5667 3427 5668 3431
rect 3838 3426 3844 3427
rect 5662 3426 5668 3427
rect 3838 3369 3844 3370
rect 5662 3369 5668 3370
rect 3838 3365 3839 3369
rect 3843 3365 3844 3369
rect 3838 3364 3844 3365
rect 3886 3368 3892 3369
rect 3886 3364 3887 3368
rect 3891 3364 3892 3368
rect 3886 3363 3892 3364
rect 4150 3368 4156 3369
rect 4150 3364 4151 3368
rect 4155 3364 4156 3368
rect 4150 3363 4156 3364
rect 4422 3368 4428 3369
rect 4422 3364 4423 3368
rect 4427 3364 4428 3368
rect 4422 3363 4428 3364
rect 4670 3368 4676 3369
rect 4670 3364 4671 3368
rect 4675 3364 4676 3368
rect 4670 3363 4676 3364
rect 4894 3368 4900 3369
rect 4894 3364 4895 3368
rect 4899 3364 4900 3368
rect 4894 3363 4900 3364
rect 5110 3368 5116 3369
rect 5110 3364 5111 3368
rect 5115 3364 5116 3368
rect 5110 3363 5116 3364
rect 5326 3368 5332 3369
rect 5326 3364 5327 3368
rect 5331 3364 5332 3368
rect 5326 3363 5332 3364
rect 5542 3368 5548 3369
rect 5542 3364 5543 3368
rect 5547 3364 5548 3368
rect 5662 3365 5663 3369
rect 5667 3365 5668 3369
rect 5662 3364 5668 3365
rect 5542 3363 5548 3364
rect 3858 3353 3864 3354
rect 3838 3352 3844 3353
rect 3838 3348 3839 3352
rect 3843 3348 3844 3352
rect 3858 3349 3859 3353
rect 3863 3349 3864 3353
rect 3858 3348 3864 3349
rect 4122 3353 4128 3354
rect 4122 3349 4123 3353
rect 4127 3349 4128 3353
rect 4122 3348 4128 3349
rect 4394 3353 4400 3354
rect 4394 3349 4395 3353
rect 4399 3349 4400 3353
rect 4394 3348 4400 3349
rect 4642 3353 4648 3354
rect 4642 3349 4643 3353
rect 4647 3349 4648 3353
rect 4642 3348 4648 3349
rect 4866 3353 4872 3354
rect 4866 3349 4867 3353
rect 4871 3349 4872 3353
rect 4866 3348 4872 3349
rect 5082 3353 5088 3354
rect 5082 3349 5083 3353
rect 5087 3349 5088 3353
rect 5082 3348 5088 3349
rect 5298 3353 5304 3354
rect 5298 3349 5299 3353
rect 5303 3349 5304 3353
rect 5298 3348 5304 3349
rect 5514 3353 5520 3354
rect 5514 3349 5515 3353
rect 5519 3349 5520 3353
rect 5514 3348 5520 3349
rect 5662 3352 5668 3353
rect 5662 3348 5663 3352
rect 5667 3348 5668 3352
rect 3838 3347 3844 3348
rect 5662 3347 5668 3348
rect 110 3296 116 3297
rect 1934 3296 1940 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 466 3295 472 3296
rect 466 3291 467 3295
rect 471 3291 472 3295
rect 466 3290 472 3291
rect 666 3295 672 3296
rect 666 3291 667 3295
rect 671 3291 672 3295
rect 666 3290 672 3291
rect 874 3295 880 3296
rect 874 3291 875 3295
rect 879 3291 880 3295
rect 874 3290 880 3291
rect 1090 3295 1096 3296
rect 1090 3291 1091 3295
rect 1095 3291 1096 3295
rect 1090 3290 1096 3291
rect 1314 3295 1320 3296
rect 1314 3291 1315 3295
rect 1319 3291 1320 3295
rect 1934 3292 1935 3296
rect 1939 3292 1940 3296
rect 1934 3291 1940 3292
rect 1314 3290 1320 3291
rect 494 3280 500 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 494 3276 495 3280
rect 499 3276 500 3280
rect 494 3275 500 3276
rect 694 3280 700 3281
rect 694 3276 695 3280
rect 699 3276 700 3280
rect 694 3275 700 3276
rect 902 3280 908 3281
rect 902 3276 903 3280
rect 907 3276 908 3280
rect 902 3275 908 3276
rect 1118 3280 1124 3281
rect 1118 3276 1119 3280
rect 1123 3276 1124 3280
rect 1118 3275 1124 3276
rect 1342 3280 1348 3281
rect 1342 3276 1343 3280
rect 1347 3276 1348 3280
rect 1342 3275 1348 3276
rect 1934 3279 1940 3280
rect 1934 3275 1935 3279
rect 1939 3275 1940 3279
rect 110 3274 116 3275
rect 1934 3274 1940 3275
rect 1974 3268 1980 3269
rect 3798 3268 3804 3269
rect 1974 3264 1975 3268
rect 1979 3264 1980 3268
rect 1974 3263 1980 3264
rect 1994 3267 2000 3268
rect 1994 3263 1995 3267
rect 1999 3263 2000 3267
rect 1994 3262 2000 3263
rect 2194 3267 2200 3268
rect 2194 3263 2195 3267
rect 2199 3263 2200 3267
rect 2194 3262 2200 3263
rect 2410 3267 2416 3268
rect 2410 3263 2411 3267
rect 2415 3263 2416 3267
rect 2410 3262 2416 3263
rect 2618 3267 2624 3268
rect 2618 3263 2619 3267
rect 2623 3263 2624 3267
rect 2618 3262 2624 3263
rect 2810 3267 2816 3268
rect 2810 3263 2811 3267
rect 2815 3263 2816 3267
rect 2810 3262 2816 3263
rect 3002 3267 3008 3268
rect 3002 3263 3003 3267
rect 3007 3263 3008 3267
rect 3002 3262 3008 3263
rect 3186 3267 3192 3268
rect 3186 3263 3187 3267
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3370 3267 3376 3268
rect 3370 3263 3371 3267
rect 3375 3263 3376 3267
rect 3370 3262 3376 3263
rect 3554 3267 3560 3268
rect 3554 3263 3555 3267
rect 3559 3263 3560 3267
rect 3798 3264 3799 3268
rect 3803 3264 3804 3268
rect 3798 3263 3804 3264
rect 3554 3262 3560 3263
rect 2022 3252 2028 3253
rect 1974 3251 1980 3252
rect 1974 3247 1975 3251
rect 1979 3247 1980 3251
rect 2022 3248 2023 3252
rect 2027 3248 2028 3252
rect 2022 3247 2028 3248
rect 2222 3252 2228 3253
rect 2222 3248 2223 3252
rect 2227 3248 2228 3252
rect 2222 3247 2228 3248
rect 2438 3252 2444 3253
rect 2438 3248 2439 3252
rect 2443 3248 2444 3252
rect 2438 3247 2444 3248
rect 2646 3252 2652 3253
rect 2646 3248 2647 3252
rect 2651 3248 2652 3252
rect 2646 3247 2652 3248
rect 2838 3252 2844 3253
rect 2838 3248 2839 3252
rect 2843 3248 2844 3252
rect 2838 3247 2844 3248
rect 3030 3252 3036 3253
rect 3030 3248 3031 3252
rect 3035 3248 3036 3252
rect 3030 3247 3036 3248
rect 3214 3252 3220 3253
rect 3214 3248 3215 3252
rect 3219 3248 3220 3252
rect 3214 3247 3220 3248
rect 3398 3252 3404 3253
rect 3398 3248 3399 3252
rect 3403 3248 3404 3252
rect 3398 3247 3404 3248
rect 3582 3252 3588 3253
rect 3582 3248 3583 3252
rect 3587 3248 3588 3252
rect 3582 3247 3588 3248
rect 3798 3251 3804 3252
rect 3798 3247 3799 3251
rect 3803 3247 3804 3251
rect 1974 3246 1980 3247
rect 3798 3246 3804 3247
rect 110 3221 116 3222
rect 1934 3221 1940 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 110 3216 116 3217
rect 534 3220 540 3221
rect 534 3216 535 3220
rect 539 3216 540 3220
rect 534 3215 540 3216
rect 726 3220 732 3221
rect 726 3216 727 3220
rect 731 3216 732 3220
rect 726 3215 732 3216
rect 918 3220 924 3221
rect 918 3216 919 3220
rect 923 3216 924 3220
rect 918 3215 924 3216
rect 1110 3220 1116 3221
rect 1110 3216 1111 3220
rect 1115 3216 1116 3220
rect 1110 3215 1116 3216
rect 1294 3220 1300 3221
rect 1294 3216 1295 3220
rect 1299 3216 1300 3220
rect 1294 3215 1300 3216
rect 1470 3220 1476 3221
rect 1470 3216 1471 3220
rect 1475 3216 1476 3220
rect 1470 3215 1476 3216
rect 1654 3220 1660 3221
rect 1654 3216 1655 3220
rect 1659 3216 1660 3220
rect 1654 3215 1660 3216
rect 1814 3220 1820 3221
rect 1814 3216 1815 3220
rect 1819 3216 1820 3220
rect 1934 3217 1935 3221
rect 1939 3217 1940 3221
rect 1934 3216 1940 3217
rect 3838 3220 3844 3221
rect 5662 3220 5668 3221
rect 3838 3216 3839 3220
rect 3843 3216 3844 3220
rect 1814 3215 1820 3216
rect 3838 3215 3844 3216
rect 3858 3219 3864 3220
rect 3858 3215 3859 3219
rect 3863 3215 3864 3219
rect 3858 3214 3864 3215
rect 4098 3219 4104 3220
rect 4098 3215 4099 3219
rect 4103 3215 4104 3219
rect 4098 3214 4104 3215
rect 4346 3219 4352 3220
rect 4346 3215 4347 3219
rect 4351 3215 4352 3219
rect 4346 3214 4352 3215
rect 4578 3219 4584 3220
rect 4578 3215 4579 3219
rect 4583 3215 4584 3219
rect 4578 3214 4584 3215
rect 4786 3219 4792 3220
rect 4786 3215 4787 3219
rect 4791 3215 4792 3219
rect 4786 3214 4792 3215
rect 4986 3219 4992 3220
rect 4986 3215 4987 3219
rect 4991 3215 4992 3219
rect 4986 3214 4992 3215
rect 5170 3219 5176 3220
rect 5170 3215 5171 3219
rect 5175 3215 5176 3219
rect 5170 3214 5176 3215
rect 5354 3219 5360 3220
rect 5354 3215 5355 3219
rect 5359 3215 5360 3219
rect 5354 3214 5360 3215
rect 5514 3219 5520 3220
rect 5514 3215 5515 3219
rect 5519 3215 5520 3219
rect 5662 3216 5663 3220
rect 5667 3216 5668 3220
rect 5662 3215 5668 3216
rect 5514 3214 5520 3215
rect 506 3205 512 3206
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 506 3201 507 3205
rect 511 3201 512 3205
rect 506 3200 512 3201
rect 698 3205 704 3206
rect 698 3201 699 3205
rect 703 3201 704 3205
rect 698 3200 704 3201
rect 890 3205 896 3206
rect 890 3201 891 3205
rect 895 3201 896 3205
rect 890 3200 896 3201
rect 1082 3205 1088 3206
rect 1082 3201 1083 3205
rect 1087 3201 1088 3205
rect 1082 3200 1088 3201
rect 1266 3205 1272 3206
rect 1266 3201 1267 3205
rect 1271 3201 1272 3205
rect 1266 3200 1272 3201
rect 1442 3205 1448 3206
rect 1442 3201 1443 3205
rect 1447 3201 1448 3205
rect 1442 3200 1448 3201
rect 1626 3205 1632 3206
rect 1626 3201 1627 3205
rect 1631 3201 1632 3205
rect 1626 3200 1632 3201
rect 1786 3205 1792 3206
rect 1786 3201 1787 3205
rect 1791 3201 1792 3205
rect 1786 3200 1792 3201
rect 1934 3204 1940 3205
rect 3886 3204 3892 3205
rect 1934 3200 1935 3204
rect 1939 3200 1940 3204
rect 110 3199 116 3200
rect 1934 3199 1940 3200
rect 3838 3203 3844 3204
rect 3838 3199 3839 3203
rect 3843 3199 3844 3203
rect 3886 3200 3887 3204
rect 3891 3200 3892 3204
rect 3886 3199 3892 3200
rect 4126 3204 4132 3205
rect 4126 3200 4127 3204
rect 4131 3200 4132 3204
rect 4126 3199 4132 3200
rect 4374 3204 4380 3205
rect 4374 3200 4375 3204
rect 4379 3200 4380 3204
rect 4374 3199 4380 3200
rect 4606 3204 4612 3205
rect 4606 3200 4607 3204
rect 4611 3200 4612 3204
rect 4606 3199 4612 3200
rect 4814 3204 4820 3205
rect 4814 3200 4815 3204
rect 4819 3200 4820 3204
rect 4814 3199 4820 3200
rect 5014 3204 5020 3205
rect 5014 3200 5015 3204
rect 5019 3200 5020 3204
rect 5014 3199 5020 3200
rect 5198 3204 5204 3205
rect 5198 3200 5199 3204
rect 5203 3200 5204 3204
rect 5198 3199 5204 3200
rect 5382 3204 5388 3205
rect 5382 3200 5383 3204
rect 5387 3200 5388 3204
rect 5382 3199 5388 3200
rect 5542 3204 5548 3205
rect 5542 3200 5543 3204
rect 5547 3200 5548 3204
rect 5542 3199 5548 3200
rect 5662 3203 5668 3204
rect 5662 3199 5663 3203
rect 5667 3199 5668 3203
rect 3838 3198 3844 3199
rect 5662 3198 5668 3199
rect 1974 3193 1980 3194
rect 3798 3193 3804 3194
rect 1974 3189 1975 3193
rect 1979 3189 1980 3193
rect 1974 3188 1980 3189
rect 2462 3192 2468 3193
rect 2462 3188 2463 3192
rect 2467 3188 2468 3192
rect 2462 3187 2468 3188
rect 2662 3192 2668 3193
rect 2662 3188 2663 3192
rect 2667 3188 2668 3192
rect 2662 3187 2668 3188
rect 2862 3192 2868 3193
rect 2862 3188 2863 3192
rect 2867 3188 2868 3192
rect 2862 3187 2868 3188
rect 3054 3192 3060 3193
rect 3054 3188 3055 3192
rect 3059 3188 3060 3192
rect 3054 3187 3060 3188
rect 3238 3192 3244 3193
rect 3238 3188 3239 3192
rect 3243 3188 3244 3192
rect 3238 3187 3244 3188
rect 3430 3192 3436 3193
rect 3430 3188 3431 3192
rect 3435 3188 3436 3192
rect 3430 3187 3436 3188
rect 3622 3192 3628 3193
rect 3622 3188 3623 3192
rect 3627 3188 3628 3192
rect 3798 3189 3799 3193
rect 3803 3189 3804 3193
rect 3798 3188 3804 3189
rect 3622 3187 3628 3188
rect 2434 3177 2440 3178
rect 1974 3176 1980 3177
rect 1974 3172 1975 3176
rect 1979 3172 1980 3176
rect 2434 3173 2435 3177
rect 2439 3173 2440 3177
rect 2434 3172 2440 3173
rect 2634 3177 2640 3178
rect 2634 3173 2635 3177
rect 2639 3173 2640 3177
rect 2634 3172 2640 3173
rect 2834 3177 2840 3178
rect 2834 3173 2835 3177
rect 2839 3173 2840 3177
rect 2834 3172 2840 3173
rect 3026 3177 3032 3178
rect 3026 3173 3027 3177
rect 3031 3173 3032 3177
rect 3026 3172 3032 3173
rect 3210 3177 3216 3178
rect 3210 3173 3211 3177
rect 3215 3173 3216 3177
rect 3210 3172 3216 3173
rect 3402 3177 3408 3178
rect 3402 3173 3403 3177
rect 3407 3173 3408 3177
rect 3402 3172 3408 3173
rect 3594 3177 3600 3178
rect 3594 3173 3595 3177
rect 3599 3173 3600 3177
rect 3594 3172 3600 3173
rect 3798 3176 3804 3177
rect 3798 3172 3799 3176
rect 3803 3172 3804 3176
rect 1974 3171 1980 3172
rect 3798 3171 3804 3172
rect 3838 3129 3844 3130
rect 5662 3129 5668 3130
rect 3838 3125 3839 3129
rect 3843 3125 3844 3129
rect 3838 3124 3844 3125
rect 3902 3128 3908 3129
rect 3902 3124 3903 3128
rect 3907 3124 3908 3128
rect 3902 3123 3908 3124
rect 4134 3128 4140 3129
rect 4134 3124 4135 3128
rect 4139 3124 4140 3128
rect 4134 3123 4140 3124
rect 4358 3128 4364 3129
rect 4358 3124 4359 3128
rect 4363 3124 4364 3128
rect 4358 3123 4364 3124
rect 4582 3128 4588 3129
rect 4582 3124 4583 3128
rect 4587 3124 4588 3128
rect 4582 3123 4588 3124
rect 4806 3128 4812 3129
rect 4806 3124 4807 3128
rect 4811 3124 4812 3128
rect 4806 3123 4812 3124
rect 5030 3128 5036 3129
rect 5030 3124 5031 3128
rect 5035 3124 5036 3128
rect 5662 3125 5663 3129
rect 5667 3125 5668 3129
rect 5662 3124 5668 3125
rect 5030 3123 5036 3124
rect 3874 3113 3880 3114
rect 3838 3112 3844 3113
rect 3838 3108 3839 3112
rect 3843 3108 3844 3112
rect 3874 3109 3875 3113
rect 3879 3109 3880 3113
rect 3874 3108 3880 3109
rect 4106 3113 4112 3114
rect 4106 3109 4107 3113
rect 4111 3109 4112 3113
rect 4106 3108 4112 3109
rect 4330 3113 4336 3114
rect 4330 3109 4331 3113
rect 4335 3109 4336 3113
rect 4330 3108 4336 3109
rect 4554 3113 4560 3114
rect 4554 3109 4555 3113
rect 4559 3109 4560 3113
rect 4554 3108 4560 3109
rect 4778 3113 4784 3114
rect 4778 3109 4779 3113
rect 4783 3109 4784 3113
rect 4778 3108 4784 3109
rect 5002 3113 5008 3114
rect 5002 3109 5003 3113
rect 5007 3109 5008 3113
rect 5002 3108 5008 3109
rect 5662 3112 5668 3113
rect 5662 3108 5663 3112
rect 5667 3108 5668 3112
rect 3838 3107 3844 3108
rect 5662 3107 5668 3108
rect 110 3064 116 3065
rect 1934 3064 1940 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 426 3063 432 3064
rect 426 3059 427 3063
rect 431 3059 432 3063
rect 426 3058 432 3059
rect 562 3063 568 3064
rect 562 3059 563 3063
rect 567 3059 568 3063
rect 562 3058 568 3059
rect 698 3063 704 3064
rect 698 3059 699 3063
rect 703 3059 704 3063
rect 698 3058 704 3059
rect 834 3063 840 3064
rect 834 3059 835 3063
rect 839 3059 840 3063
rect 834 3058 840 3059
rect 970 3063 976 3064
rect 970 3059 971 3063
rect 975 3059 976 3063
rect 970 3058 976 3059
rect 1106 3063 1112 3064
rect 1106 3059 1107 3063
rect 1111 3059 1112 3063
rect 1106 3058 1112 3059
rect 1242 3063 1248 3064
rect 1242 3059 1243 3063
rect 1247 3059 1248 3063
rect 1242 3058 1248 3059
rect 1378 3063 1384 3064
rect 1378 3059 1379 3063
rect 1383 3059 1384 3063
rect 1378 3058 1384 3059
rect 1514 3063 1520 3064
rect 1514 3059 1515 3063
rect 1519 3059 1520 3063
rect 1514 3058 1520 3059
rect 1650 3063 1656 3064
rect 1650 3059 1651 3063
rect 1655 3059 1656 3063
rect 1650 3058 1656 3059
rect 1786 3063 1792 3064
rect 1786 3059 1787 3063
rect 1791 3059 1792 3063
rect 1934 3060 1935 3064
rect 1939 3060 1940 3064
rect 1934 3059 1940 3060
rect 1786 3058 1792 3059
rect 454 3048 460 3049
rect 110 3047 116 3048
rect 110 3043 111 3047
rect 115 3043 116 3047
rect 454 3044 455 3048
rect 459 3044 460 3048
rect 454 3043 460 3044
rect 590 3048 596 3049
rect 590 3044 591 3048
rect 595 3044 596 3048
rect 590 3043 596 3044
rect 726 3048 732 3049
rect 726 3044 727 3048
rect 731 3044 732 3048
rect 726 3043 732 3044
rect 862 3048 868 3049
rect 862 3044 863 3048
rect 867 3044 868 3048
rect 862 3043 868 3044
rect 998 3048 1004 3049
rect 998 3044 999 3048
rect 1003 3044 1004 3048
rect 998 3043 1004 3044
rect 1134 3048 1140 3049
rect 1134 3044 1135 3048
rect 1139 3044 1140 3048
rect 1134 3043 1140 3044
rect 1270 3048 1276 3049
rect 1270 3044 1271 3048
rect 1275 3044 1276 3048
rect 1270 3043 1276 3044
rect 1406 3048 1412 3049
rect 1406 3044 1407 3048
rect 1411 3044 1412 3048
rect 1406 3043 1412 3044
rect 1542 3048 1548 3049
rect 1542 3044 1543 3048
rect 1547 3044 1548 3048
rect 1542 3043 1548 3044
rect 1678 3048 1684 3049
rect 1678 3044 1679 3048
rect 1683 3044 1684 3048
rect 1678 3043 1684 3044
rect 1814 3048 1820 3049
rect 1814 3044 1815 3048
rect 1819 3044 1820 3048
rect 1814 3043 1820 3044
rect 1934 3047 1940 3048
rect 1934 3043 1935 3047
rect 1939 3043 1940 3047
rect 110 3042 116 3043
rect 1934 3042 1940 3043
rect 1974 3032 1980 3033
rect 3798 3032 3804 3033
rect 1974 3028 1975 3032
rect 1979 3028 1980 3032
rect 1974 3027 1980 3028
rect 2330 3031 2336 3032
rect 2330 3027 2331 3031
rect 2335 3027 2336 3031
rect 2330 3026 2336 3027
rect 2554 3031 2560 3032
rect 2554 3027 2555 3031
rect 2559 3027 2560 3031
rect 2554 3026 2560 3027
rect 2778 3031 2784 3032
rect 2778 3027 2779 3031
rect 2783 3027 2784 3031
rect 2778 3026 2784 3027
rect 3002 3031 3008 3032
rect 3002 3027 3003 3031
rect 3007 3027 3008 3031
rect 3002 3026 3008 3027
rect 3234 3031 3240 3032
rect 3234 3027 3235 3031
rect 3239 3027 3240 3031
rect 3234 3026 3240 3027
rect 3466 3031 3472 3032
rect 3466 3027 3467 3031
rect 3471 3027 3472 3031
rect 3798 3028 3799 3032
rect 3803 3028 3804 3032
rect 3798 3027 3804 3028
rect 3466 3026 3472 3027
rect 2358 3016 2364 3017
rect 1974 3015 1980 3016
rect 1974 3011 1975 3015
rect 1979 3011 1980 3015
rect 2358 3012 2359 3016
rect 2363 3012 2364 3016
rect 2358 3011 2364 3012
rect 2582 3016 2588 3017
rect 2582 3012 2583 3016
rect 2587 3012 2588 3016
rect 2582 3011 2588 3012
rect 2806 3016 2812 3017
rect 2806 3012 2807 3016
rect 2811 3012 2812 3016
rect 2806 3011 2812 3012
rect 3030 3016 3036 3017
rect 3030 3012 3031 3016
rect 3035 3012 3036 3016
rect 3030 3011 3036 3012
rect 3262 3016 3268 3017
rect 3262 3012 3263 3016
rect 3267 3012 3268 3016
rect 3262 3011 3268 3012
rect 3494 3016 3500 3017
rect 3494 3012 3495 3016
rect 3499 3012 3500 3016
rect 3494 3011 3500 3012
rect 3798 3015 3804 3016
rect 3798 3011 3799 3015
rect 3803 3011 3804 3015
rect 1974 3010 1980 3011
rect 3798 3010 3804 3011
rect 3838 2980 3844 2981
rect 5662 2980 5668 2981
rect 3838 2976 3839 2980
rect 3843 2976 3844 2980
rect 3838 2975 3844 2976
rect 3906 2979 3912 2980
rect 3906 2975 3907 2979
rect 3911 2975 3912 2979
rect 3906 2974 3912 2975
rect 4074 2979 4080 2980
rect 4074 2975 4075 2979
rect 4079 2975 4080 2979
rect 4074 2974 4080 2975
rect 4242 2979 4248 2980
rect 4242 2975 4243 2979
rect 4247 2975 4248 2979
rect 4242 2974 4248 2975
rect 4410 2979 4416 2980
rect 4410 2975 4411 2979
rect 4415 2975 4416 2979
rect 4410 2974 4416 2975
rect 4578 2979 4584 2980
rect 4578 2975 4579 2979
rect 4583 2975 4584 2979
rect 4578 2974 4584 2975
rect 4754 2979 4760 2980
rect 4754 2975 4755 2979
rect 4759 2975 4760 2979
rect 5662 2976 5663 2980
rect 5667 2976 5668 2980
rect 5662 2975 5668 2976
rect 4754 2974 4760 2975
rect 3934 2964 3940 2965
rect 3838 2963 3844 2964
rect 110 2961 116 2962
rect 1934 2961 1940 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 110 2956 116 2957
rect 198 2960 204 2961
rect 198 2956 199 2960
rect 203 2956 204 2960
rect 198 2955 204 2956
rect 510 2960 516 2961
rect 510 2956 511 2960
rect 515 2956 516 2960
rect 510 2955 516 2956
rect 814 2960 820 2961
rect 814 2956 815 2960
rect 819 2956 820 2960
rect 814 2955 820 2956
rect 1110 2960 1116 2961
rect 1110 2956 1111 2960
rect 1115 2956 1116 2960
rect 1110 2955 1116 2956
rect 1414 2960 1420 2961
rect 1414 2956 1415 2960
rect 1419 2956 1420 2960
rect 1414 2955 1420 2956
rect 1718 2960 1724 2961
rect 1718 2956 1719 2960
rect 1723 2956 1724 2960
rect 1934 2957 1935 2961
rect 1939 2957 1940 2961
rect 3838 2959 3839 2963
rect 3843 2959 3844 2963
rect 3934 2960 3935 2964
rect 3939 2960 3940 2964
rect 3934 2959 3940 2960
rect 4102 2964 4108 2965
rect 4102 2960 4103 2964
rect 4107 2960 4108 2964
rect 4102 2959 4108 2960
rect 4270 2964 4276 2965
rect 4270 2960 4271 2964
rect 4275 2960 4276 2964
rect 4270 2959 4276 2960
rect 4438 2964 4444 2965
rect 4438 2960 4439 2964
rect 4443 2960 4444 2964
rect 4438 2959 4444 2960
rect 4606 2964 4612 2965
rect 4606 2960 4607 2964
rect 4611 2960 4612 2964
rect 4606 2959 4612 2960
rect 4782 2964 4788 2965
rect 4782 2960 4783 2964
rect 4787 2960 4788 2964
rect 4782 2959 4788 2960
rect 5662 2963 5668 2964
rect 5662 2959 5663 2963
rect 5667 2959 5668 2963
rect 3838 2958 3844 2959
rect 5662 2958 5668 2959
rect 1934 2956 1940 2957
rect 1718 2955 1724 2956
rect 170 2945 176 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 170 2941 171 2945
rect 175 2941 176 2945
rect 170 2940 176 2941
rect 482 2945 488 2946
rect 482 2941 483 2945
rect 487 2941 488 2945
rect 482 2940 488 2941
rect 786 2945 792 2946
rect 786 2941 787 2945
rect 791 2941 792 2945
rect 786 2940 792 2941
rect 1082 2945 1088 2946
rect 1082 2941 1083 2945
rect 1087 2941 1088 2945
rect 1082 2940 1088 2941
rect 1386 2945 1392 2946
rect 1386 2941 1387 2945
rect 1391 2941 1392 2945
rect 1386 2940 1392 2941
rect 1690 2945 1696 2946
rect 1974 2945 1980 2946
rect 3798 2945 3804 2946
rect 1690 2941 1691 2945
rect 1695 2941 1696 2945
rect 1690 2940 1696 2941
rect 1934 2944 1940 2945
rect 1934 2940 1935 2944
rect 1939 2940 1940 2944
rect 1974 2941 1975 2945
rect 1979 2941 1980 2945
rect 1974 2940 1980 2941
rect 2142 2944 2148 2945
rect 2142 2940 2143 2944
rect 2147 2940 2148 2944
rect 110 2939 116 2940
rect 1934 2939 1940 2940
rect 2142 2939 2148 2940
rect 2342 2944 2348 2945
rect 2342 2940 2343 2944
rect 2347 2940 2348 2944
rect 2342 2939 2348 2940
rect 2542 2944 2548 2945
rect 2542 2940 2543 2944
rect 2547 2940 2548 2944
rect 2542 2939 2548 2940
rect 2742 2944 2748 2945
rect 2742 2940 2743 2944
rect 2747 2940 2748 2944
rect 2742 2939 2748 2940
rect 2934 2944 2940 2945
rect 2934 2940 2935 2944
rect 2939 2940 2940 2944
rect 2934 2939 2940 2940
rect 3134 2944 3140 2945
rect 3134 2940 3135 2944
rect 3139 2940 3140 2944
rect 3134 2939 3140 2940
rect 3334 2944 3340 2945
rect 3334 2940 3335 2944
rect 3339 2940 3340 2944
rect 3798 2941 3799 2945
rect 3803 2941 3804 2945
rect 3798 2940 3804 2941
rect 3334 2939 3340 2940
rect 2114 2929 2120 2930
rect 1974 2928 1980 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 2114 2925 2115 2929
rect 2119 2925 2120 2929
rect 2114 2924 2120 2925
rect 2314 2929 2320 2930
rect 2314 2925 2315 2929
rect 2319 2925 2320 2929
rect 2314 2924 2320 2925
rect 2514 2929 2520 2930
rect 2514 2925 2515 2929
rect 2519 2925 2520 2929
rect 2514 2924 2520 2925
rect 2714 2929 2720 2930
rect 2714 2925 2715 2929
rect 2719 2925 2720 2929
rect 2714 2924 2720 2925
rect 2906 2929 2912 2930
rect 2906 2925 2907 2929
rect 2911 2925 2912 2929
rect 2906 2924 2912 2925
rect 3106 2929 3112 2930
rect 3106 2925 3107 2929
rect 3111 2925 3112 2929
rect 3106 2924 3112 2925
rect 3306 2929 3312 2930
rect 3306 2925 3307 2929
rect 3311 2925 3312 2929
rect 3306 2924 3312 2925
rect 3798 2928 3804 2929
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 1974 2923 1980 2924
rect 3798 2923 3804 2924
rect 3838 2901 3844 2902
rect 5662 2901 5668 2902
rect 3838 2897 3839 2901
rect 3843 2897 3844 2901
rect 3838 2896 3844 2897
rect 3894 2900 3900 2901
rect 3894 2896 3895 2900
rect 3899 2896 3900 2900
rect 3894 2895 3900 2896
rect 4030 2900 4036 2901
rect 4030 2896 4031 2900
rect 4035 2896 4036 2900
rect 4030 2895 4036 2896
rect 4166 2900 4172 2901
rect 4166 2896 4167 2900
rect 4171 2896 4172 2900
rect 4166 2895 4172 2896
rect 4302 2900 4308 2901
rect 4302 2896 4303 2900
rect 4307 2896 4308 2900
rect 4302 2895 4308 2896
rect 4438 2900 4444 2901
rect 4438 2896 4439 2900
rect 4443 2896 4444 2900
rect 4438 2895 4444 2896
rect 4574 2900 4580 2901
rect 4574 2896 4575 2900
rect 4579 2896 4580 2900
rect 5662 2897 5663 2901
rect 5667 2897 5668 2901
rect 5662 2896 5668 2897
rect 4574 2895 4580 2896
rect 3866 2885 3872 2886
rect 3838 2884 3844 2885
rect 3838 2880 3839 2884
rect 3843 2880 3844 2884
rect 3866 2881 3867 2885
rect 3871 2881 3872 2885
rect 3866 2880 3872 2881
rect 4002 2885 4008 2886
rect 4002 2881 4003 2885
rect 4007 2881 4008 2885
rect 4002 2880 4008 2881
rect 4138 2885 4144 2886
rect 4138 2881 4139 2885
rect 4143 2881 4144 2885
rect 4138 2880 4144 2881
rect 4274 2885 4280 2886
rect 4274 2881 4275 2885
rect 4279 2881 4280 2885
rect 4274 2880 4280 2881
rect 4410 2885 4416 2886
rect 4410 2881 4411 2885
rect 4415 2881 4416 2885
rect 4410 2880 4416 2881
rect 4546 2885 4552 2886
rect 4546 2881 4547 2885
rect 4551 2881 4552 2885
rect 4546 2880 4552 2881
rect 5662 2884 5668 2885
rect 5662 2880 5663 2884
rect 5667 2880 5668 2884
rect 3838 2879 3844 2880
rect 5662 2879 5668 2880
rect 110 2812 116 2813
rect 1934 2812 1940 2813
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 130 2811 136 2812
rect 130 2807 131 2811
rect 135 2807 136 2811
rect 130 2806 136 2807
rect 306 2811 312 2812
rect 306 2807 307 2811
rect 311 2807 312 2811
rect 306 2806 312 2807
rect 522 2811 528 2812
rect 522 2807 523 2811
rect 527 2807 528 2811
rect 522 2806 528 2807
rect 762 2811 768 2812
rect 762 2807 763 2811
rect 767 2807 768 2811
rect 762 2806 768 2807
rect 1010 2811 1016 2812
rect 1010 2807 1011 2811
rect 1015 2807 1016 2811
rect 1010 2806 1016 2807
rect 1274 2811 1280 2812
rect 1274 2807 1275 2811
rect 1279 2807 1280 2811
rect 1274 2806 1280 2807
rect 1538 2811 1544 2812
rect 1538 2807 1539 2811
rect 1543 2807 1544 2811
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 1538 2806 1544 2807
rect 158 2796 164 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 158 2792 159 2796
rect 163 2792 164 2796
rect 158 2791 164 2792
rect 334 2796 340 2797
rect 334 2792 335 2796
rect 339 2792 340 2796
rect 334 2791 340 2792
rect 550 2796 556 2797
rect 550 2792 551 2796
rect 555 2792 556 2796
rect 550 2791 556 2792
rect 790 2796 796 2797
rect 790 2792 791 2796
rect 795 2792 796 2796
rect 790 2791 796 2792
rect 1038 2796 1044 2797
rect 1038 2792 1039 2796
rect 1043 2792 1044 2796
rect 1038 2791 1044 2792
rect 1302 2796 1308 2797
rect 1302 2792 1303 2796
rect 1307 2792 1308 2796
rect 1302 2791 1308 2792
rect 1566 2796 1572 2797
rect 1566 2792 1567 2796
rect 1571 2792 1572 2796
rect 1566 2791 1572 2792
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 110 2790 116 2791
rect 1934 2790 1940 2791
rect 1974 2788 1980 2789
rect 3798 2788 3804 2789
rect 1974 2784 1975 2788
rect 1979 2784 1980 2788
rect 1974 2783 1980 2784
rect 2010 2787 2016 2788
rect 2010 2783 2011 2787
rect 2015 2783 2016 2787
rect 2010 2782 2016 2783
rect 2258 2787 2264 2788
rect 2258 2783 2259 2787
rect 2263 2783 2264 2787
rect 2258 2782 2264 2783
rect 2506 2787 2512 2788
rect 2506 2783 2507 2787
rect 2511 2783 2512 2787
rect 2506 2782 2512 2783
rect 2754 2787 2760 2788
rect 2754 2783 2755 2787
rect 2759 2783 2760 2787
rect 2754 2782 2760 2783
rect 3002 2787 3008 2788
rect 3002 2783 3003 2787
rect 3007 2783 3008 2787
rect 3798 2784 3799 2788
rect 3803 2784 3804 2788
rect 3798 2783 3804 2784
rect 3002 2782 3008 2783
rect 2038 2772 2044 2773
rect 1974 2771 1980 2772
rect 1974 2767 1975 2771
rect 1979 2767 1980 2771
rect 2038 2768 2039 2772
rect 2043 2768 2044 2772
rect 2038 2767 2044 2768
rect 2286 2772 2292 2773
rect 2286 2768 2287 2772
rect 2291 2768 2292 2772
rect 2286 2767 2292 2768
rect 2534 2772 2540 2773
rect 2534 2768 2535 2772
rect 2539 2768 2540 2772
rect 2534 2767 2540 2768
rect 2782 2772 2788 2773
rect 2782 2768 2783 2772
rect 2787 2768 2788 2772
rect 2782 2767 2788 2768
rect 3030 2772 3036 2773
rect 3030 2768 3031 2772
rect 3035 2768 3036 2772
rect 3030 2767 3036 2768
rect 3798 2771 3804 2772
rect 3798 2767 3799 2771
rect 3803 2767 3804 2771
rect 1974 2766 1980 2767
rect 3798 2766 3804 2767
rect 3838 2744 3844 2745
rect 5662 2744 5668 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4810 2738 4816 2739
rect 110 2733 116 2734
rect 1934 2733 1940 2734
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 278 2732 284 2733
rect 278 2728 279 2732
rect 283 2728 284 2732
rect 278 2727 284 2728
rect 454 2732 460 2733
rect 454 2728 455 2732
rect 459 2728 460 2732
rect 454 2727 460 2728
rect 646 2732 652 2733
rect 646 2728 647 2732
rect 651 2728 652 2732
rect 646 2727 652 2728
rect 854 2732 860 2733
rect 854 2728 855 2732
rect 859 2728 860 2732
rect 854 2727 860 2728
rect 1078 2732 1084 2733
rect 1078 2728 1079 2732
rect 1083 2728 1084 2732
rect 1078 2727 1084 2728
rect 1310 2732 1316 2733
rect 1310 2728 1311 2732
rect 1315 2728 1316 2732
rect 1310 2727 1316 2728
rect 1550 2732 1556 2733
rect 1550 2728 1551 2732
rect 1555 2728 1556 2732
rect 1550 2727 1556 2728
rect 1798 2732 1804 2733
rect 1798 2728 1799 2732
rect 1803 2728 1804 2732
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 3886 2728 3892 2729
rect 1798 2727 1804 2728
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 3838 2722 3844 2723
rect 5662 2722 5668 2723
rect 250 2717 256 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 250 2713 251 2717
rect 255 2713 256 2717
rect 250 2712 256 2713
rect 426 2717 432 2718
rect 426 2713 427 2717
rect 431 2713 432 2717
rect 426 2712 432 2713
rect 618 2717 624 2718
rect 618 2713 619 2717
rect 623 2713 624 2717
rect 618 2712 624 2713
rect 826 2717 832 2718
rect 826 2713 827 2717
rect 831 2713 832 2717
rect 826 2712 832 2713
rect 1050 2717 1056 2718
rect 1050 2713 1051 2717
rect 1055 2713 1056 2717
rect 1050 2712 1056 2713
rect 1282 2717 1288 2718
rect 1282 2713 1283 2717
rect 1287 2713 1288 2717
rect 1282 2712 1288 2713
rect 1522 2717 1528 2718
rect 1522 2713 1523 2717
rect 1527 2713 1528 2717
rect 1522 2712 1528 2713
rect 1770 2717 1776 2718
rect 1770 2713 1771 2717
rect 1775 2713 1776 2717
rect 1770 2712 1776 2713
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 110 2711 116 2712
rect 1934 2711 1940 2712
rect 1974 2709 1980 2710
rect 3798 2709 3804 2710
rect 1974 2705 1975 2709
rect 1979 2705 1980 2709
rect 1974 2704 1980 2705
rect 2022 2708 2028 2709
rect 2022 2704 2023 2708
rect 2027 2704 2028 2708
rect 2022 2703 2028 2704
rect 2246 2708 2252 2709
rect 2246 2704 2247 2708
rect 2251 2704 2252 2708
rect 2246 2703 2252 2704
rect 2502 2708 2508 2709
rect 2502 2704 2503 2708
rect 2507 2704 2508 2708
rect 2502 2703 2508 2704
rect 2758 2708 2764 2709
rect 2758 2704 2759 2708
rect 2763 2704 2764 2708
rect 2758 2703 2764 2704
rect 3014 2708 3020 2709
rect 3014 2704 3015 2708
rect 3019 2704 3020 2708
rect 3798 2705 3799 2709
rect 3803 2705 3804 2709
rect 3798 2704 3804 2705
rect 3014 2703 3020 2704
rect 1994 2693 2000 2694
rect 1974 2692 1980 2693
rect 1974 2688 1975 2692
rect 1979 2688 1980 2692
rect 1994 2689 1995 2693
rect 1999 2689 2000 2693
rect 1994 2688 2000 2689
rect 2218 2693 2224 2694
rect 2218 2689 2219 2693
rect 2223 2689 2224 2693
rect 2218 2688 2224 2689
rect 2474 2693 2480 2694
rect 2474 2689 2475 2693
rect 2479 2689 2480 2693
rect 2474 2688 2480 2689
rect 2730 2693 2736 2694
rect 2730 2689 2731 2693
rect 2735 2689 2736 2693
rect 2730 2688 2736 2689
rect 2986 2693 2992 2694
rect 2986 2689 2987 2693
rect 2991 2689 2992 2693
rect 2986 2688 2992 2689
rect 3798 2692 3804 2693
rect 3798 2688 3799 2692
rect 3803 2688 3804 2692
rect 1974 2687 1980 2688
rect 3798 2687 3804 2688
rect 3838 2669 3844 2670
rect 5662 2669 5668 2670
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 3958 2668 3964 2669
rect 3958 2664 3959 2668
rect 3963 2664 3964 2668
rect 3958 2663 3964 2664
rect 4254 2668 4260 2669
rect 4254 2664 4255 2668
rect 4259 2664 4260 2668
rect 4254 2663 4260 2664
rect 4542 2668 4548 2669
rect 4542 2664 4543 2668
rect 4547 2664 4548 2668
rect 4542 2663 4548 2664
rect 4822 2668 4828 2669
rect 4822 2664 4823 2668
rect 4827 2664 4828 2668
rect 4822 2663 4828 2664
rect 5110 2668 5116 2669
rect 5110 2664 5111 2668
rect 5115 2664 5116 2668
rect 5110 2663 5116 2664
rect 5398 2668 5404 2669
rect 5398 2664 5399 2668
rect 5403 2664 5404 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5398 2663 5404 2664
rect 3930 2653 3936 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 3930 2649 3931 2653
rect 3935 2649 3936 2653
rect 3930 2648 3936 2649
rect 4226 2653 4232 2654
rect 4226 2649 4227 2653
rect 4231 2649 4232 2653
rect 4226 2648 4232 2649
rect 4514 2653 4520 2654
rect 4514 2649 4515 2653
rect 4519 2649 4520 2653
rect 4514 2648 4520 2649
rect 4794 2653 4800 2654
rect 4794 2649 4795 2653
rect 4799 2649 4800 2653
rect 4794 2648 4800 2649
rect 5082 2653 5088 2654
rect 5082 2649 5083 2653
rect 5087 2649 5088 2653
rect 5082 2648 5088 2649
rect 5370 2653 5376 2654
rect 5370 2649 5371 2653
rect 5375 2649 5376 2653
rect 5370 2648 5376 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 3838 2647 3844 2648
rect 5662 2647 5668 2648
rect 110 2584 116 2585
rect 1934 2584 1940 2585
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 570 2583 576 2584
rect 570 2579 571 2583
rect 575 2579 576 2583
rect 570 2578 576 2579
rect 730 2583 736 2584
rect 730 2579 731 2583
rect 735 2579 736 2583
rect 730 2578 736 2579
rect 890 2583 896 2584
rect 890 2579 891 2583
rect 895 2579 896 2583
rect 890 2578 896 2579
rect 1042 2583 1048 2584
rect 1042 2579 1043 2583
rect 1047 2579 1048 2583
rect 1042 2578 1048 2579
rect 1194 2583 1200 2584
rect 1194 2579 1195 2583
rect 1199 2579 1200 2583
rect 1194 2578 1200 2579
rect 1354 2583 1360 2584
rect 1354 2579 1355 2583
rect 1359 2579 1360 2583
rect 1354 2578 1360 2579
rect 1514 2583 1520 2584
rect 1514 2579 1515 2583
rect 1519 2579 1520 2583
rect 1514 2578 1520 2579
rect 1674 2583 1680 2584
rect 1674 2579 1675 2583
rect 1679 2579 1680 2583
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1674 2578 1680 2579
rect 598 2568 604 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 598 2564 599 2568
rect 603 2564 604 2568
rect 598 2563 604 2564
rect 758 2568 764 2569
rect 758 2564 759 2568
rect 763 2564 764 2568
rect 758 2563 764 2564
rect 918 2568 924 2569
rect 918 2564 919 2568
rect 923 2564 924 2568
rect 918 2563 924 2564
rect 1070 2568 1076 2569
rect 1070 2564 1071 2568
rect 1075 2564 1076 2568
rect 1070 2563 1076 2564
rect 1222 2568 1228 2569
rect 1222 2564 1223 2568
rect 1227 2564 1228 2568
rect 1222 2563 1228 2564
rect 1382 2568 1388 2569
rect 1382 2564 1383 2568
rect 1387 2564 1388 2568
rect 1382 2563 1388 2564
rect 1542 2568 1548 2569
rect 1542 2564 1543 2568
rect 1547 2564 1548 2568
rect 1542 2563 1548 2564
rect 1702 2568 1708 2569
rect 1702 2564 1703 2568
rect 1707 2564 1708 2568
rect 1702 2563 1708 2564
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 110 2562 116 2563
rect 1934 2562 1940 2563
rect 1974 2548 1980 2549
rect 3798 2548 3804 2549
rect 1974 2544 1975 2548
rect 1979 2544 1980 2548
rect 1974 2543 1980 2544
rect 2554 2547 2560 2548
rect 2554 2543 2555 2547
rect 2559 2543 2560 2547
rect 2554 2542 2560 2543
rect 2690 2547 2696 2548
rect 2690 2543 2691 2547
rect 2695 2543 2696 2547
rect 2690 2542 2696 2543
rect 2826 2547 2832 2548
rect 2826 2543 2827 2547
rect 2831 2543 2832 2547
rect 2826 2542 2832 2543
rect 2962 2547 2968 2548
rect 2962 2543 2963 2547
rect 2967 2543 2968 2547
rect 2962 2542 2968 2543
rect 3098 2547 3104 2548
rect 3098 2543 3099 2547
rect 3103 2543 3104 2547
rect 3798 2544 3799 2548
rect 3803 2544 3804 2548
rect 3798 2543 3804 2544
rect 3098 2542 3104 2543
rect 2582 2532 2588 2533
rect 1974 2531 1980 2532
rect 1974 2527 1975 2531
rect 1979 2527 1980 2531
rect 2582 2528 2583 2532
rect 2587 2528 2588 2532
rect 2582 2527 2588 2528
rect 2718 2532 2724 2533
rect 2718 2528 2719 2532
rect 2723 2528 2724 2532
rect 2718 2527 2724 2528
rect 2854 2532 2860 2533
rect 2854 2528 2855 2532
rect 2859 2528 2860 2532
rect 2854 2527 2860 2528
rect 2990 2532 2996 2533
rect 2990 2528 2991 2532
rect 2995 2528 2996 2532
rect 2990 2527 2996 2528
rect 3126 2532 3132 2533
rect 3126 2528 3127 2532
rect 3131 2528 3132 2532
rect 3126 2527 3132 2528
rect 3798 2531 3804 2532
rect 3798 2527 3799 2531
rect 3803 2527 3804 2531
rect 1974 2526 1980 2527
rect 3798 2526 3804 2527
rect 3838 2520 3844 2521
rect 5662 2520 5668 2521
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 3838 2515 3844 2516
rect 3858 2519 3864 2520
rect 3858 2515 3859 2519
rect 3863 2515 3864 2519
rect 3858 2514 3864 2515
rect 4082 2519 4088 2520
rect 4082 2515 4083 2519
rect 4087 2515 4088 2519
rect 4082 2514 4088 2515
rect 4330 2519 4336 2520
rect 4330 2515 4331 2519
rect 4335 2515 4336 2519
rect 4330 2514 4336 2515
rect 4578 2519 4584 2520
rect 4578 2515 4579 2519
rect 4583 2515 4584 2519
rect 4578 2514 4584 2515
rect 4826 2519 4832 2520
rect 4826 2515 4827 2519
rect 4831 2515 4832 2519
rect 4826 2514 4832 2515
rect 5074 2519 5080 2520
rect 5074 2515 5075 2519
rect 5079 2515 5080 2519
rect 5074 2514 5080 2515
rect 5322 2519 5328 2520
rect 5322 2515 5323 2519
rect 5327 2515 5328 2519
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 5662 2515 5668 2516
rect 5322 2514 5328 2515
rect 110 2509 116 2510
rect 1934 2509 1940 2510
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 382 2508 388 2509
rect 382 2504 383 2508
rect 387 2504 388 2508
rect 382 2503 388 2504
rect 598 2508 604 2509
rect 598 2504 599 2508
rect 603 2504 604 2508
rect 598 2503 604 2504
rect 814 2508 820 2509
rect 814 2504 815 2508
rect 819 2504 820 2508
rect 814 2503 820 2504
rect 1022 2508 1028 2509
rect 1022 2504 1023 2508
rect 1027 2504 1028 2508
rect 1022 2503 1028 2504
rect 1230 2508 1236 2509
rect 1230 2504 1231 2508
rect 1235 2504 1236 2508
rect 1230 2503 1236 2504
rect 1430 2508 1436 2509
rect 1430 2504 1431 2508
rect 1435 2504 1436 2508
rect 1430 2503 1436 2504
rect 1630 2508 1636 2509
rect 1630 2504 1631 2508
rect 1635 2504 1636 2508
rect 1630 2503 1636 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 3886 2504 3892 2505
rect 1814 2503 1820 2504
rect 3838 2503 3844 2504
rect 3838 2499 3839 2503
rect 3843 2499 3844 2503
rect 3886 2500 3887 2504
rect 3891 2500 3892 2504
rect 3886 2499 3892 2500
rect 4110 2504 4116 2505
rect 4110 2500 4111 2504
rect 4115 2500 4116 2504
rect 4110 2499 4116 2500
rect 4358 2504 4364 2505
rect 4358 2500 4359 2504
rect 4363 2500 4364 2504
rect 4358 2499 4364 2500
rect 4606 2504 4612 2505
rect 4606 2500 4607 2504
rect 4611 2500 4612 2504
rect 4606 2499 4612 2500
rect 4854 2504 4860 2505
rect 4854 2500 4855 2504
rect 4859 2500 4860 2504
rect 4854 2499 4860 2500
rect 5102 2504 5108 2505
rect 5102 2500 5103 2504
rect 5107 2500 5108 2504
rect 5102 2499 5108 2500
rect 5350 2504 5356 2505
rect 5350 2500 5351 2504
rect 5355 2500 5356 2504
rect 5350 2499 5356 2500
rect 5662 2503 5668 2504
rect 5662 2499 5663 2503
rect 5667 2499 5668 2503
rect 3838 2498 3844 2499
rect 5662 2498 5668 2499
rect 354 2493 360 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 354 2489 355 2493
rect 359 2489 360 2493
rect 354 2488 360 2489
rect 570 2493 576 2494
rect 570 2489 571 2493
rect 575 2489 576 2493
rect 570 2488 576 2489
rect 786 2493 792 2494
rect 786 2489 787 2493
rect 791 2489 792 2493
rect 786 2488 792 2489
rect 994 2493 1000 2494
rect 994 2489 995 2493
rect 999 2489 1000 2493
rect 994 2488 1000 2489
rect 1202 2493 1208 2494
rect 1202 2489 1203 2493
rect 1207 2489 1208 2493
rect 1202 2488 1208 2489
rect 1402 2493 1408 2494
rect 1402 2489 1403 2493
rect 1407 2489 1408 2493
rect 1402 2488 1408 2489
rect 1602 2493 1608 2494
rect 1602 2489 1603 2493
rect 1607 2489 1608 2493
rect 1602 2488 1608 2489
rect 1786 2493 1792 2494
rect 1786 2489 1787 2493
rect 1791 2489 1792 2493
rect 1786 2488 1792 2489
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 110 2487 116 2488
rect 1934 2487 1940 2488
rect 1974 2449 1980 2450
rect 3798 2449 3804 2450
rect 1974 2445 1975 2449
rect 1979 2445 1980 2449
rect 1974 2444 1980 2445
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2222 2448 2228 2449
rect 2222 2444 2223 2448
rect 2227 2444 2228 2448
rect 2222 2443 2228 2444
rect 2446 2448 2452 2449
rect 2446 2444 2447 2448
rect 2451 2444 2452 2448
rect 2446 2443 2452 2444
rect 2678 2448 2684 2449
rect 2678 2444 2679 2448
rect 2683 2444 2684 2448
rect 2678 2443 2684 2444
rect 2926 2448 2932 2449
rect 2926 2444 2927 2448
rect 2931 2444 2932 2448
rect 2926 2443 2932 2444
rect 3182 2448 3188 2449
rect 3182 2444 3183 2448
rect 3187 2444 3188 2448
rect 3182 2443 3188 2444
rect 3438 2448 3444 2449
rect 3438 2444 3439 2448
rect 3443 2444 3444 2448
rect 3438 2443 3444 2444
rect 3678 2448 3684 2449
rect 3678 2444 3679 2448
rect 3683 2444 3684 2448
rect 3798 2445 3799 2449
rect 3803 2445 3804 2449
rect 3798 2444 3804 2445
rect 3678 2443 3684 2444
rect 3838 2441 3844 2442
rect 5662 2441 5668 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3886 2440 3892 2441
rect 3886 2436 3887 2440
rect 3891 2436 3892 2440
rect 3886 2435 3892 2436
rect 4086 2440 4092 2441
rect 4086 2436 4087 2440
rect 4091 2436 4092 2440
rect 4086 2435 4092 2436
rect 4326 2440 4332 2441
rect 4326 2436 4327 2440
rect 4331 2436 4332 2440
rect 4326 2435 4332 2436
rect 4582 2440 4588 2441
rect 4582 2436 4583 2440
rect 4587 2436 4588 2440
rect 4582 2435 4588 2436
rect 4846 2440 4852 2441
rect 4846 2436 4847 2440
rect 4851 2436 4852 2440
rect 4846 2435 4852 2436
rect 5118 2440 5124 2441
rect 5118 2436 5119 2440
rect 5123 2436 5124 2440
rect 5118 2435 5124 2436
rect 5398 2440 5404 2441
rect 5398 2436 5399 2440
rect 5403 2436 5404 2440
rect 5662 2437 5663 2441
rect 5667 2437 5668 2441
rect 5662 2436 5668 2437
rect 5398 2435 5404 2436
rect 1994 2433 2000 2434
rect 1974 2432 1980 2433
rect 1974 2428 1975 2432
rect 1979 2428 1980 2432
rect 1994 2429 1995 2433
rect 1999 2429 2000 2433
rect 1994 2428 2000 2429
rect 2194 2433 2200 2434
rect 2194 2429 2195 2433
rect 2199 2429 2200 2433
rect 2194 2428 2200 2429
rect 2418 2433 2424 2434
rect 2418 2429 2419 2433
rect 2423 2429 2424 2433
rect 2418 2428 2424 2429
rect 2650 2433 2656 2434
rect 2650 2429 2651 2433
rect 2655 2429 2656 2433
rect 2650 2428 2656 2429
rect 2898 2433 2904 2434
rect 2898 2429 2899 2433
rect 2903 2429 2904 2433
rect 2898 2428 2904 2429
rect 3154 2433 3160 2434
rect 3154 2429 3155 2433
rect 3159 2429 3160 2433
rect 3154 2428 3160 2429
rect 3410 2433 3416 2434
rect 3410 2429 3411 2433
rect 3415 2429 3416 2433
rect 3410 2428 3416 2429
rect 3650 2433 3656 2434
rect 3650 2429 3651 2433
rect 3655 2429 3656 2433
rect 3650 2428 3656 2429
rect 3798 2432 3804 2433
rect 3798 2428 3799 2432
rect 3803 2428 3804 2432
rect 1974 2427 1980 2428
rect 3798 2427 3804 2428
rect 3858 2425 3864 2426
rect 3838 2424 3844 2425
rect 3838 2420 3839 2424
rect 3843 2420 3844 2424
rect 3858 2421 3859 2425
rect 3863 2421 3864 2425
rect 3858 2420 3864 2421
rect 4058 2425 4064 2426
rect 4058 2421 4059 2425
rect 4063 2421 4064 2425
rect 4058 2420 4064 2421
rect 4298 2425 4304 2426
rect 4298 2421 4299 2425
rect 4303 2421 4304 2425
rect 4298 2420 4304 2421
rect 4554 2425 4560 2426
rect 4554 2421 4555 2425
rect 4559 2421 4560 2425
rect 4554 2420 4560 2421
rect 4818 2425 4824 2426
rect 4818 2421 4819 2425
rect 4823 2421 4824 2425
rect 4818 2420 4824 2421
rect 5090 2425 5096 2426
rect 5090 2421 5091 2425
rect 5095 2421 5096 2425
rect 5090 2420 5096 2421
rect 5370 2425 5376 2426
rect 5370 2421 5371 2425
rect 5375 2421 5376 2425
rect 5370 2420 5376 2421
rect 5662 2424 5668 2425
rect 5662 2420 5663 2424
rect 5667 2420 5668 2424
rect 3838 2419 3844 2420
rect 5662 2419 5668 2420
rect 110 2356 116 2357
rect 1934 2356 1940 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 226 2355 232 2356
rect 226 2351 227 2355
rect 231 2351 232 2355
rect 226 2350 232 2351
rect 522 2355 528 2356
rect 522 2351 523 2355
rect 527 2351 528 2355
rect 522 2350 528 2351
rect 834 2355 840 2356
rect 834 2351 835 2355
rect 839 2351 840 2355
rect 834 2350 840 2351
rect 1154 2355 1160 2356
rect 1154 2351 1155 2355
rect 1159 2351 1160 2355
rect 1154 2350 1160 2351
rect 1482 2355 1488 2356
rect 1482 2351 1483 2355
rect 1487 2351 1488 2355
rect 1482 2350 1488 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1934 2351 1940 2352
rect 1786 2350 1792 2351
rect 254 2340 260 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 254 2336 255 2340
rect 259 2336 260 2340
rect 254 2335 260 2336
rect 550 2340 556 2341
rect 550 2336 551 2340
rect 555 2336 556 2340
rect 550 2335 556 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 1182 2340 1188 2341
rect 1182 2336 1183 2340
rect 1187 2336 1188 2340
rect 1182 2335 1188 2336
rect 1510 2340 1516 2341
rect 1510 2336 1511 2340
rect 1515 2336 1516 2340
rect 1510 2335 1516 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 110 2334 116 2335
rect 1934 2334 1940 2335
rect 1974 2292 1980 2293
rect 3798 2292 3804 2293
rect 1974 2288 1975 2292
rect 1979 2288 1980 2292
rect 1974 2287 1980 2288
rect 1994 2291 2000 2292
rect 1994 2287 1995 2291
rect 1999 2287 2000 2291
rect 1994 2286 2000 2287
rect 2154 2291 2160 2292
rect 2154 2287 2155 2291
rect 2159 2287 2160 2291
rect 2154 2286 2160 2287
rect 2346 2291 2352 2292
rect 2346 2287 2347 2291
rect 2351 2287 2352 2291
rect 2346 2286 2352 2287
rect 2538 2291 2544 2292
rect 2538 2287 2539 2291
rect 2543 2287 2544 2291
rect 2538 2286 2544 2287
rect 2730 2291 2736 2292
rect 2730 2287 2731 2291
rect 2735 2287 2736 2291
rect 2730 2286 2736 2287
rect 2922 2291 2928 2292
rect 2922 2287 2923 2291
rect 2927 2287 2928 2291
rect 2922 2286 2928 2287
rect 3114 2291 3120 2292
rect 3114 2287 3115 2291
rect 3119 2287 3120 2291
rect 3114 2286 3120 2287
rect 3298 2291 3304 2292
rect 3298 2287 3299 2291
rect 3303 2287 3304 2291
rect 3298 2286 3304 2287
rect 3482 2291 3488 2292
rect 3482 2287 3483 2291
rect 3487 2287 3488 2291
rect 3482 2286 3488 2287
rect 3650 2291 3656 2292
rect 3650 2287 3651 2291
rect 3655 2287 3656 2291
rect 3798 2288 3799 2292
rect 3803 2288 3804 2292
rect 3798 2287 3804 2288
rect 3650 2286 3656 2287
rect 3838 2280 3844 2281
rect 5662 2280 5668 2281
rect 2022 2276 2028 2277
rect 1974 2275 1980 2276
rect 1974 2271 1975 2275
rect 1979 2271 1980 2275
rect 2022 2272 2023 2276
rect 2027 2272 2028 2276
rect 2022 2271 2028 2272
rect 2182 2276 2188 2277
rect 2182 2272 2183 2276
rect 2187 2272 2188 2276
rect 2182 2271 2188 2272
rect 2374 2276 2380 2277
rect 2374 2272 2375 2276
rect 2379 2272 2380 2276
rect 2374 2271 2380 2272
rect 2566 2276 2572 2277
rect 2566 2272 2567 2276
rect 2571 2272 2572 2276
rect 2566 2271 2572 2272
rect 2758 2276 2764 2277
rect 2758 2272 2759 2276
rect 2763 2272 2764 2276
rect 2758 2271 2764 2272
rect 2950 2276 2956 2277
rect 2950 2272 2951 2276
rect 2955 2272 2956 2276
rect 2950 2271 2956 2272
rect 3142 2276 3148 2277
rect 3142 2272 3143 2276
rect 3147 2272 3148 2276
rect 3142 2271 3148 2272
rect 3326 2276 3332 2277
rect 3326 2272 3327 2276
rect 3331 2272 3332 2276
rect 3326 2271 3332 2272
rect 3510 2276 3516 2277
rect 3510 2272 3511 2276
rect 3515 2272 3516 2276
rect 3510 2271 3516 2272
rect 3678 2276 3684 2277
rect 3838 2276 3839 2280
rect 3843 2276 3844 2280
rect 3678 2272 3679 2276
rect 3683 2272 3684 2276
rect 3678 2271 3684 2272
rect 3798 2275 3804 2276
rect 3838 2275 3844 2276
rect 4442 2279 4448 2280
rect 4442 2275 4443 2279
rect 4447 2275 4448 2279
rect 3798 2271 3799 2275
rect 3803 2271 3804 2275
rect 4442 2274 4448 2275
rect 4610 2279 4616 2280
rect 4610 2275 4611 2279
rect 4615 2275 4616 2279
rect 4610 2274 4616 2275
rect 4786 2279 4792 2280
rect 4786 2275 4787 2279
rect 4791 2275 4792 2279
rect 4786 2274 4792 2275
rect 4962 2279 4968 2280
rect 4962 2275 4963 2279
rect 4967 2275 4968 2279
rect 4962 2274 4968 2275
rect 5146 2279 5152 2280
rect 5146 2275 5147 2279
rect 5151 2275 5152 2279
rect 5146 2274 5152 2275
rect 5338 2279 5344 2280
rect 5338 2275 5339 2279
rect 5343 2275 5344 2279
rect 5338 2274 5344 2275
rect 5514 2279 5520 2280
rect 5514 2275 5515 2279
rect 5519 2275 5520 2279
rect 5662 2276 5663 2280
rect 5667 2276 5668 2280
rect 5662 2275 5668 2276
rect 5514 2274 5520 2275
rect 1974 2270 1980 2271
rect 3798 2270 3804 2271
rect 110 2265 116 2266
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 366 2264 372 2265
rect 366 2260 367 2264
rect 371 2260 372 2264
rect 366 2259 372 2260
rect 598 2264 604 2265
rect 598 2260 599 2264
rect 603 2260 604 2264
rect 598 2259 604 2260
rect 830 2264 836 2265
rect 830 2260 831 2264
rect 835 2260 836 2264
rect 830 2259 836 2260
rect 1062 2264 1068 2265
rect 1062 2260 1063 2264
rect 1067 2260 1068 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 4470 2264 4476 2265
rect 1934 2260 1940 2261
rect 3838 2263 3844 2264
rect 1062 2259 1068 2260
rect 3838 2259 3839 2263
rect 3843 2259 3844 2263
rect 4470 2260 4471 2264
rect 4475 2260 4476 2264
rect 4470 2259 4476 2260
rect 4638 2264 4644 2265
rect 4638 2260 4639 2264
rect 4643 2260 4644 2264
rect 4638 2259 4644 2260
rect 4814 2264 4820 2265
rect 4814 2260 4815 2264
rect 4819 2260 4820 2264
rect 4814 2259 4820 2260
rect 4990 2264 4996 2265
rect 4990 2260 4991 2264
rect 4995 2260 4996 2264
rect 4990 2259 4996 2260
rect 5174 2264 5180 2265
rect 5174 2260 5175 2264
rect 5179 2260 5180 2264
rect 5174 2259 5180 2260
rect 5366 2264 5372 2265
rect 5366 2260 5367 2264
rect 5371 2260 5372 2264
rect 5366 2259 5372 2260
rect 5542 2264 5548 2265
rect 5542 2260 5543 2264
rect 5547 2260 5548 2264
rect 5542 2259 5548 2260
rect 5662 2263 5668 2264
rect 5662 2259 5663 2263
rect 5667 2259 5668 2263
rect 3838 2258 3844 2259
rect 5662 2258 5668 2259
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 338 2249 344 2250
rect 338 2245 339 2249
rect 343 2245 344 2249
rect 338 2244 344 2245
rect 570 2249 576 2250
rect 570 2245 571 2249
rect 575 2245 576 2249
rect 570 2244 576 2245
rect 802 2249 808 2250
rect 802 2245 803 2249
rect 807 2245 808 2249
rect 802 2244 808 2245
rect 1034 2249 1040 2250
rect 1034 2245 1035 2249
rect 1039 2245 1040 2249
rect 1034 2244 1040 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 110 2243 116 2244
rect 1934 2243 1940 2244
rect 1974 2209 1980 2210
rect 3798 2209 3804 2210
rect 1974 2205 1975 2209
rect 1979 2205 1980 2209
rect 1974 2204 1980 2205
rect 2022 2208 2028 2209
rect 2022 2204 2023 2208
rect 2027 2204 2028 2208
rect 2022 2203 2028 2204
rect 2190 2208 2196 2209
rect 2190 2204 2191 2208
rect 2195 2204 2196 2208
rect 2190 2203 2196 2204
rect 2358 2208 2364 2209
rect 2358 2204 2359 2208
rect 2363 2204 2364 2208
rect 2358 2203 2364 2204
rect 2534 2208 2540 2209
rect 2534 2204 2535 2208
rect 2539 2204 2540 2208
rect 2534 2203 2540 2204
rect 2710 2208 2716 2209
rect 2710 2204 2711 2208
rect 2715 2204 2716 2208
rect 2710 2203 2716 2204
rect 2878 2208 2884 2209
rect 2878 2204 2879 2208
rect 2883 2204 2884 2208
rect 2878 2203 2884 2204
rect 3046 2208 3052 2209
rect 3046 2204 3047 2208
rect 3051 2204 3052 2208
rect 3046 2203 3052 2204
rect 3206 2208 3212 2209
rect 3206 2204 3207 2208
rect 3211 2204 3212 2208
rect 3206 2203 3212 2204
rect 3366 2208 3372 2209
rect 3366 2204 3367 2208
rect 3371 2204 3372 2208
rect 3366 2203 3372 2204
rect 3534 2208 3540 2209
rect 3534 2204 3535 2208
rect 3539 2204 3540 2208
rect 3534 2203 3540 2204
rect 3678 2208 3684 2209
rect 3678 2204 3679 2208
rect 3683 2204 3684 2208
rect 3798 2205 3799 2209
rect 3803 2205 3804 2209
rect 3798 2204 3804 2205
rect 3678 2203 3684 2204
rect 1994 2193 2000 2194
rect 1974 2192 1980 2193
rect 1974 2188 1975 2192
rect 1979 2188 1980 2192
rect 1994 2189 1995 2193
rect 1999 2189 2000 2193
rect 1994 2188 2000 2189
rect 2162 2193 2168 2194
rect 2162 2189 2163 2193
rect 2167 2189 2168 2193
rect 2162 2188 2168 2189
rect 2330 2193 2336 2194
rect 2330 2189 2331 2193
rect 2335 2189 2336 2193
rect 2330 2188 2336 2189
rect 2506 2193 2512 2194
rect 2506 2189 2507 2193
rect 2511 2189 2512 2193
rect 2506 2188 2512 2189
rect 2682 2193 2688 2194
rect 2682 2189 2683 2193
rect 2687 2189 2688 2193
rect 2682 2188 2688 2189
rect 2850 2193 2856 2194
rect 2850 2189 2851 2193
rect 2855 2189 2856 2193
rect 2850 2188 2856 2189
rect 3018 2193 3024 2194
rect 3018 2189 3019 2193
rect 3023 2189 3024 2193
rect 3018 2188 3024 2189
rect 3178 2193 3184 2194
rect 3178 2189 3179 2193
rect 3183 2189 3184 2193
rect 3178 2188 3184 2189
rect 3338 2193 3344 2194
rect 3338 2189 3339 2193
rect 3343 2189 3344 2193
rect 3338 2188 3344 2189
rect 3506 2193 3512 2194
rect 3506 2189 3507 2193
rect 3511 2189 3512 2193
rect 3506 2188 3512 2189
rect 3650 2193 3656 2194
rect 3838 2193 3844 2194
rect 5662 2193 5668 2194
rect 3650 2189 3651 2193
rect 3655 2189 3656 2193
rect 3650 2188 3656 2189
rect 3798 2192 3804 2193
rect 3798 2188 3799 2192
rect 3803 2188 3804 2192
rect 3838 2189 3839 2193
rect 3843 2189 3844 2193
rect 3838 2188 3844 2189
rect 4542 2192 4548 2193
rect 4542 2188 4543 2192
rect 4547 2188 4548 2192
rect 1974 2187 1980 2188
rect 3798 2187 3804 2188
rect 4542 2187 4548 2188
rect 4718 2192 4724 2193
rect 4718 2188 4719 2192
rect 4723 2188 4724 2192
rect 4718 2187 4724 2188
rect 4910 2192 4916 2193
rect 4910 2188 4911 2192
rect 4915 2188 4916 2192
rect 4910 2187 4916 2188
rect 5118 2192 5124 2193
rect 5118 2188 5119 2192
rect 5123 2188 5124 2192
rect 5118 2187 5124 2188
rect 5334 2192 5340 2193
rect 5334 2188 5335 2192
rect 5339 2188 5340 2192
rect 5334 2187 5340 2188
rect 5542 2192 5548 2193
rect 5542 2188 5543 2192
rect 5547 2188 5548 2192
rect 5662 2189 5663 2193
rect 5667 2189 5668 2193
rect 5662 2188 5668 2189
rect 5542 2187 5548 2188
rect 4514 2177 4520 2178
rect 3838 2176 3844 2177
rect 3838 2172 3839 2176
rect 3843 2172 3844 2176
rect 4514 2173 4515 2177
rect 4519 2173 4520 2177
rect 4514 2172 4520 2173
rect 4690 2177 4696 2178
rect 4690 2173 4691 2177
rect 4695 2173 4696 2177
rect 4690 2172 4696 2173
rect 4882 2177 4888 2178
rect 4882 2173 4883 2177
rect 4887 2173 4888 2177
rect 4882 2172 4888 2173
rect 5090 2177 5096 2178
rect 5090 2173 5091 2177
rect 5095 2173 5096 2177
rect 5090 2172 5096 2173
rect 5306 2177 5312 2178
rect 5306 2173 5307 2177
rect 5311 2173 5312 2177
rect 5306 2172 5312 2173
rect 5514 2177 5520 2178
rect 5514 2173 5515 2177
rect 5519 2173 5520 2177
rect 5514 2172 5520 2173
rect 5662 2176 5668 2177
rect 5662 2172 5663 2176
rect 5667 2172 5668 2176
rect 3838 2171 3844 2172
rect 5662 2171 5668 2172
rect 110 2104 116 2105
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 346 2103 352 2104
rect 346 2099 347 2103
rect 351 2099 352 2103
rect 346 2098 352 2099
rect 594 2103 600 2104
rect 594 2099 595 2103
rect 599 2099 600 2103
rect 594 2098 600 2099
rect 834 2103 840 2104
rect 834 2099 835 2103
rect 839 2099 840 2103
rect 834 2098 840 2099
rect 1074 2103 1080 2104
rect 1074 2099 1075 2103
rect 1079 2099 1080 2103
rect 1074 2098 1080 2099
rect 1314 2103 1320 2104
rect 1314 2099 1315 2103
rect 1319 2099 1320 2103
rect 1314 2098 1320 2099
rect 1562 2103 1568 2104
rect 1562 2099 1563 2103
rect 1567 2099 1568 2103
rect 1562 2098 1568 2099
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1786 2098 1792 2099
rect 158 2088 164 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 374 2088 380 2089
rect 374 2084 375 2088
rect 379 2084 380 2088
rect 374 2083 380 2084
rect 622 2088 628 2089
rect 622 2084 623 2088
rect 627 2084 628 2088
rect 622 2083 628 2084
rect 862 2088 868 2089
rect 862 2084 863 2088
rect 867 2084 868 2088
rect 862 2083 868 2084
rect 1102 2088 1108 2089
rect 1102 2084 1103 2088
rect 1107 2084 1108 2088
rect 1102 2083 1108 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1590 2088 1596 2089
rect 1590 2084 1591 2088
rect 1595 2084 1596 2088
rect 1590 2083 1596 2084
rect 1814 2088 1820 2089
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 110 2082 116 2083
rect 1934 2082 1940 2083
rect 1974 2044 1980 2045
rect 3798 2044 3804 2045
rect 1974 2040 1975 2044
rect 1979 2040 1980 2044
rect 1974 2039 1980 2040
rect 3106 2043 3112 2044
rect 3106 2039 3107 2043
rect 3111 2039 3112 2043
rect 3106 2038 3112 2039
rect 3242 2043 3248 2044
rect 3242 2039 3243 2043
rect 3247 2039 3248 2043
rect 3242 2038 3248 2039
rect 3378 2043 3384 2044
rect 3378 2039 3379 2043
rect 3383 2039 3384 2043
rect 3378 2038 3384 2039
rect 3514 2043 3520 2044
rect 3514 2039 3515 2043
rect 3519 2039 3520 2043
rect 3514 2038 3520 2039
rect 3650 2043 3656 2044
rect 3650 2039 3651 2043
rect 3655 2039 3656 2043
rect 3798 2040 3799 2044
rect 3803 2040 3804 2044
rect 3798 2039 3804 2040
rect 3838 2044 3844 2045
rect 5662 2044 5668 2045
rect 3838 2040 3839 2044
rect 3843 2040 3844 2044
rect 3838 2039 3844 2040
rect 4634 2043 4640 2044
rect 4634 2039 4635 2043
rect 4639 2039 4640 2043
rect 3650 2038 3656 2039
rect 4634 2038 4640 2039
rect 4770 2043 4776 2044
rect 4770 2039 4771 2043
rect 4775 2039 4776 2043
rect 4770 2038 4776 2039
rect 4906 2043 4912 2044
rect 4906 2039 4907 2043
rect 4911 2039 4912 2043
rect 4906 2038 4912 2039
rect 5042 2043 5048 2044
rect 5042 2039 5043 2043
rect 5047 2039 5048 2043
rect 5042 2038 5048 2039
rect 5178 2043 5184 2044
rect 5178 2039 5179 2043
rect 5183 2039 5184 2043
rect 5662 2040 5663 2044
rect 5667 2040 5668 2044
rect 5662 2039 5668 2040
rect 5178 2038 5184 2039
rect 3134 2028 3140 2029
rect 1974 2027 1980 2028
rect 110 2025 116 2026
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 270 2024 276 2025
rect 270 2020 271 2024
rect 275 2020 276 2024
rect 270 2019 276 2020
rect 406 2024 412 2025
rect 406 2020 407 2024
rect 411 2020 412 2024
rect 406 2019 412 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 686 2024 692 2025
rect 686 2020 687 2024
rect 691 2020 692 2024
rect 686 2019 692 2020
rect 830 2024 836 2025
rect 830 2020 831 2024
rect 835 2020 836 2024
rect 830 2019 836 2020
rect 974 2024 980 2025
rect 974 2020 975 2024
rect 979 2020 980 2024
rect 974 2019 980 2020
rect 1118 2024 1124 2025
rect 1118 2020 1119 2024
rect 1123 2020 1124 2024
rect 1118 2019 1124 2020
rect 1262 2024 1268 2025
rect 1262 2020 1263 2024
rect 1267 2020 1268 2024
rect 1262 2019 1268 2020
rect 1406 2024 1412 2025
rect 1406 2020 1407 2024
rect 1411 2020 1412 2024
rect 1406 2019 1412 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1974 2023 1975 2027
rect 1979 2023 1980 2027
rect 3134 2024 3135 2028
rect 3139 2024 3140 2028
rect 3134 2023 3140 2024
rect 3270 2028 3276 2029
rect 3270 2024 3271 2028
rect 3275 2024 3276 2028
rect 3270 2023 3276 2024
rect 3406 2028 3412 2029
rect 3406 2024 3407 2028
rect 3411 2024 3412 2028
rect 3406 2023 3412 2024
rect 3542 2028 3548 2029
rect 3542 2024 3543 2028
rect 3547 2024 3548 2028
rect 3542 2023 3548 2024
rect 3678 2028 3684 2029
rect 4662 2028 4668 2029
rect 3678 2024 3679 2028
rect 3683 2024 3684 2028
rect 3678 2023 3684 2024
rect 3798 2027 3804 2028
rect 3798 2023 3799 2027
rect 3803 2023 3804 2027
rect 1974 2022 1980 2023
rect 3798 2022 3804 2023
rect 3838 2027 3844 2028
rect 3838 2023 3839 2027
rect 3843 2023 3844 2027
rect 4662 2024 4663 2028
rect 4667 2024 4668 2028
rect 4662 2023 4668 2024
rect 4798 2028 4804 2029
rect 4798 2024 4799 2028
rect 4803 2024 4804 2028
rect 4798 2023 4804 2024
rect 4934 2028 4940 2029
rect 4934 2024 4935 2028
rect 4939 2024 4940 2028
rect 4934 2023 4940 2024
rect 5070 2028 5076 2029
rect 5070 2024 5071 2028
rect 5075 2024 5076 2028
rect 5070 2023 5076 2024
rect 5206 2028 5212 2029
rect 5206 2024 5207 2028
rect 5211 2024 5212 2028
rect 5206 2023 5212 2024
rect 5662 2027 5668 2028
rect 5662 2023 5663 2027
rect 5667 2023 5668 2027
rect 3838 2022 3844 2023
rect 5662 2022 5668 2023
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 242 2009 248 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 242 2005 243 2009
rect 247 2005 248 2009
rect 242 2004 248 2005
rect 378 2009 384 2010
rect 378 2005 379 2009
rect 383 2005 384 2009
rect 378 2004 384 2005
rect 514 2009 520 2010
rect 514 2005 515 2009
rect 519 2005 520 2009
rect 514 2004 520 2005
rect 658 2009 664 2010
rect 658 2005 659 2009
rect 663 2005 664 2009
rect 658 2004 664 2005
rect 802 2009 808 2010
rect 802 2005 803 2009
rect 807 2005 808 2009
rect 802 2004 808 2005
rect 946 2009 952 2010
rect 946 2005 947 2009
rect 951 2005 952 2009
rect 946 2004 952 2005
rect 1090 2009 1096 2010
rect 1090 2005 1091 2009
rect 1095 2005 1096 2009
rect 1090 2004 1096 2005
rect 1234 2009 1240 2010
rect 1234 2005 1235 2009
rect 1239 2005 1240 2009
rect 1234 2004 1240 2005
rect 1378 2009 1384 2010
rect 1378 2005 1379 2009
rect 1383 2005 1384 2009
rect 1378 2004 1384 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 110 2003 116 2004
rect 1934 2003 1940 2004
rect 1974 1969 1980 1970
rect 3798 1969 3804 1970
rect 1974 1965 1975 1969
rect 1979 1965 1980 1969
rect 1974 1964 1980 1965
rect 3126 1968 3132 1969
rect 3126 1964 3127 1968
rect 3131 1964 3132 1968
rect 3126 1963 3132 1964
rect 3262 1968 3268 1969
rect 3262 1964 3263 1968
rect 3267 1964 3268 1968
rect 3262 1963 3268 1964
rect 3398 1968 3404 1969
rect 3398 1964 3399 1968
rect 3403 1964 3404 1968
rect 3398 1963 3404 1964
rect 3534 1968 3540 1969
rect 3534 1964 3535 1968
rect 3539 1964 3540 1968
rect 3534 1963 3540 1964
rect 3670 1968 3676 1969
rect 3670 1964 3671 1968
rect 3675 1964 3676 1968
rect 3798 1965 3799 1969
rect 3803 1965 3804 1969
rect 3798 1964 3804 1965
rect 3838 1969 3844 1970
rect 5662 1969 5668 1970
rect 3838 1965 3839 1969
rect 3843 1965 3844 1969
rect 3838 1964 3844 1965
rect 4862 1968 4868 1969
rect 4862 1964 4863 1968
rect 4867 1964 4868 1968
rect 3670 1963 3676 1964
rect 4862 1963 4868 1964
rect 4998 1968 5004 1969
rect 4998 1964 4999 1968
rect 5003 1964 5004 1968
rect 4998 1963 5004 1964
rect 5134 1968 5140 1969
rect 5134 1964 5135 1968
rect 5139 1964 5140 1968
rect 5134 1963 5140 1964
rect 5270 1968 5276 1969
rect 5270 1964 5271 1968
rect 5275 1964 5276 1968
rect 5270 1963 5276 1964
rect 5406 1968 5412 1969
rect 5406 1964 5407 1968
rect 5411 1964 5412 1968
rect 5406 1963 5412 1964
rect 5542 1968 5548 1969
rect 5542 1964 5543 1968
rect 5547 1964 5548 1968
rect 5662 1965 5663 1969
rect 5667 1965 5668 1969
rect 5662 1964 5668 1965
rect 5542 1963 5548 1964
rect 3098 1953 3104 1954
rect 1974 1952 1980 1953
rect 1974 1948 1975 1952
rect 1979 1948 1980 1952
rect 3098 1949 3099 1953
rect 3103 1949 3104 1953
rect 3098 1948 3104 1949
rect 3234 1953 3240 1954
rect 3234 1949 3235 1953
rect 3239 1949 3240 1953
rect 3234 1948 3240 1949
rect 3370 1953 3376 1954
rect 3370 1949 3371 1953
rect 3375 1949 3376 1953
rect 3370 1948 3376 1949
rect 3506 1953 3512 1954
rect 3506 1949 3507 1953
rect 3511 1949 3512 1953
rect 3506 1948 3512 1949
rect 3642 1953 3648 1954
rect 4834 1953 4840 1954
rect 3642 1949 3643 1953
rect 3647 1949 3648 1953
rect 3642 1948 3648 1949
rect 3798 1952 3804 1953
rect 3798 1948 3799 1952
rect 3803 1948 3804 1952
rect 1974 1947 1980 1948
rect 3798 1947 3804 1948
rect 3838 1952 3844 1953
rect 3838 1948 3839 1952
rect 3843 1948 3844 1952
rect 4834 1949 4835 1953
rect 4839 1949 4840 1953
rect 4834 1948 4840 1949
rect 4970 1953 4976 1954
rect 4970 1949 4971 1953
rect 4975 1949 4976 1953
rect 4970 1948 4976 1949
rect 5106 1953 5112 1954
rect 5106 1949 5107 1953
rect 5111 1949 5112 1953
rect 5106 1948 5112 1949
rect 5242 1953 5248 1954
rect 5242 1949 5243 1953
rect 5247 1949 5248 1953
rect 5242 1948 5248 1949
rect 5378 1953 5384 1954
rect 5378 1949 5379 1953
rect 5383 1949 5384 1953
rect 5378 1948 5384 1949
rect 5514 1953 5520 1954
rect 5514 1949 5515 1953
rect 5519 1949 5520 1953
rect 5514 1948 5520 1949
rect 5662 1952 5668 1953
rect 5662 1948 5663 1952
rect 5667 1948 5668 1952
rect 3838 1947 3844 1948
rect 5662 1947 5668 1948
rect 110 1872 116 1873
rect 1934 1872 1940 1873
rect 110 1868 111 1872
rect 115 1868 116 1872
rect 110 1867 116 1868
rect 186 1871 192 1872
rect 186 1867 187 1871
rect 191 1867 192 1871
rect 186 1866 192 1867
rect 378 1871 384 1872
rect 378 1867 379 1871
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 586 1871 592 1872
rect 586 1867 587 1871
rect 591 1867 592 1871
rect 586 1866 592 1867
rect 810 1871 816 1872
rect 810 1867 811 1871
rect 815 1867 816 1871
rect 810 1866 816 1867
rect 1050 1871 1056 1872
rect 1050 1867 1051 1871
rect 1055 1867 1056 1871
rect 1050 1866 1056 1867
rect 1298 1871 1304 1872
rect 1298 1867 1299 1871
rect 1303 1867 1304 1871
rect 1298 1866 1304 1867
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1867 1560 1871
rect 1554 1866 1560 1867
rect 1786 1871 1792 1872
rect 1786 1867 1787 1871
rect 1791 1867 1792 1871
rect 1934 1868 1935 1872
rect 1939 1868 1940 1872
rect 1934 1867 1940 1868
rect 1786 1866 1792 1867
rect 214 1856 220 1857
rect 110 1855 116 1856
rect 110 1851 111 1855
rect 115 1851 116 1855
rect 214 1852 215 1856
rect 219 1852 220 1856
rect 214 1851 220 1852
rect 406 1856 412 1857
rect 406 1852 407 1856
rect 411 1852 412 1856
rect 406 1851 412 1852
rect 614 1856 620 1857
rect 614 1852 615 1856
rect 619 1852 620 1856
rect 614 1851 620 1852
rect 838 1856 844 1857
rect 838 1852 839 1856
rect 843 1852 844 1856
rect 838 1851 844 1852
rect 1078 1856 1084 1857
rect 1078 1852 1079 1856
rect 1083 1852 1084 1856
rect 1078 1851 1084 1852
rect 1326 1856 1332 1857
rect 1326 1852 1327 1856
rect 1331 1852 1332 1856
rect 1326 1851 1332 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1814 1856 1820 1857
rect 1814 1852 1815 1856
rect 1819 1852 1820 1856
rect 1814 1851 1820 1852
rect 1934 1855 1940 1856
rect 1934 1851 1935 1855
rect 1939 1851 1940 1855
rect 110 1850 116 1851
rect 1934 1850 1940 1851
rect 1974 1808 1980 1809
rect 3798 1808 3804 1809
rect 1974 1804 1975 1808
rect 1979 1804 1980 1808
rect 1974 1803 1980 1804
rect 1994 1807 2000 1808
rect 1994 1803 1995 1807
rect 1999 1803 2000 1807
rect 1994 1802 2000 1803
rect 2226 1807 2232 1808
rect 2226 1803 2227 1807
rect 2231 1803 2232 1807
rect 2226 1802 2232 1803
rect 2466 1807 2472 1808
rect 2466 1803 2467 1807
rect 2471 1803 2472 1807
rect 2466 1802 2472 1803
rect 2690 1807 2696 1808
rect 2690 1803 2691 1807
rect 2695 1803 2696 1807
rect 2690 1802 2696 1803
rect 2906 1807 2912 1808
rect 2906 1803 2907 1807
rect 2911 1803 2912 1807
rect 2906 1802 2912 1803
rect 3106 1807 3112 1808
rect 3106 1803 3107 1807
rect 3111 1803 3112 1807
rect 3106 1802 3112 1803
rect 3298 1807 3304 1808
rect 3298 1803 3299 1807
rect 3303 1803 3304 1807
rect 3298 1802 3304 1803
rect 3482 1807 3488 1808
rect 3482 1803 3483 1807
rect 3487 1803 3488 1807
rect 3482 1802 3488 1803
rect 3650 1807 3656 1808
rect 3650 1803 3651 1807
rect 3655 1803 3656 1807
rect 3798 1804 3799 1808
rect 3803 1804 3804 1808
rect 3798 1803 3804 1804
rect 3838 1808 3844 1809
rect 5662 1808 5668 1809
rect 3838 1804 3839 1808
rect 3843 1804 3844 1808
rect 3838 1803 3844 1804
rect 4674 1807 4680 1808
rect 4674 1803 4675 1807
rect 4679 1803 4680 1807
rect 3650 1802 3656 1803
rect 4674 1802 4680 1803
rect 4818 1807 4824 1808
rect 4818 1803 4819 1807
rect 4823 1803 4824 1807
rect 4818 1802 4824 1803
rect 4962 1807 4968 1808
rect 4962 1803 4963 1807
rect 4967 1803 4968 1807
rect 4962 1802 4968 1803
rect 5106 1807 5112 1808
rect 5106 1803 5107 1807
rect 5111 1803 5112 1807
rect 5106 1802 5112 1803
rect 5242 1807 5248 1808
rect 5242 1803 5243 1807
rect 5247 1803 5248 1807
rect 5242 1802 5248 1803
rect 5378 1807 5384 1808
rect 5378 1803 5379 1807
rect 5383 1803 5384 1807
rect 5378 1802 5384 1803
rect 5514 1807 5520 1808
rect 5514 1803 5515 1807
rect 5519 1803 5520 1807
rect 5662 1804 5663 1808
rect 5667 1804 5668 1808
rect 5662 1803 5668 1804
rect 5514 1802 5520 1803
rect 2022 1792 2028 1793
rect 1974 1791 1980 1792
rect 110 1789 116 1790
rect 1934 1789 1940 1790
rect 110 1785 111 1789
rect 115 1785 116 1789
rect 110 1784 116 1785
rect 158 1788 164 1789
rect 158 1784 159 1788
rect 163 1784 164 1788
rect 158 1783 164 1784
rect 374 1788 380 1789
rect 374 1784 375 1788
rect 379 1784 380 1788
rect 374 1783 380 1784
rect 590 1788 596 1789
rect 590 1784 591 1788
rect 595 1784 596 1788
rect 590 1783 596 1784
rect 798 1788 804 1789
rect 798 1784 799 1788
rect 803 1784 804 1788
rect 798 1783 804 1784
rect 998 1788 1004 1789
rect 998 1784 999 1788
rect 1003 1784 1004 1788
rect 998 1783 1004 1784
rect 1190 1788 1196 1789
rect 1190 1784 1191 1788
rect 1195 1784 1196 1788
rect 1190 1783 1196 1784
rect 1382 1788 1388 1789
rect 1382 1784 1383 1788
rect 1387 1784 1388 1788
rect 1382 1783 1388 1784
rect 1574 1788 1580 1789
rect 1574 1784 1575 1788
rect 1579 1784 1580 1788
rect 1934 1785 1935 1789
rect 1939 1785 1940 1789
rect 1974 1787 1975 1791
rect 1979 1787 1980 1791
rect 2022 1788 2023 1792
rect 2027 1788 2028 1792
rect 2022 1787 2028 1788
rect 2254 1792 2260 1793
rect 2254 1788 2255 1792
rect 2259 1788 2260 1792
rect 2254 1787 2260 1788
rect 2494 1792 2500 1793
rect 2494 1788 2495 1792
rect 2499 1788 2500 1792
rect 2494 1787 2500 1788
rect 2718 1792 2724 1793
rect 2718 1788 2719 1792
rect 2723 1788 2724 1792
rect 2718 1787 2724 1788
rect 2934 1792 2940 1793
rect 2934 1788 2935 1792
rect 2939 1788 2940 1792
rect 2934 1787 2940 1788
rect 3134 1792 3140 1793
rect 3134 1788 3135 1792
rect 3139 1788 3140 1792
rect 3134 1787 3140 1788
rect 3326 1792 3332 1793
rect 3326 1788 3327 1792
rect 3331 1788 3332 1792
rect 3326 1787 3332 1788
rect 3510 1792 3516 1793
rect 3510 1788 3511 1792
rect 3515 1788 3516 1792
rect 3510 1787 3516 1788
rect 3678 1792 3684 1793
rect 4702 1792 4708 1793
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3798 1791 3804 1792
rect 3798 1787 3799 1791
rect 3803 1787 3804 1791
rect 1974 1786 1980 1787
rect 3798 1786 3804 1787
rect 3838 1791 3844 1792
rect 3838 1787 3839 1791
rect 3843 1787 3844 1791
rect 4702 1788 4703 1792
rect 4707 1788 4708 1792
rect 4702 1787 4708 1788
rect 4846 1792 4852 1793
rect 4846 1788 4847 1792
rect 4851 1788 4852 1792
rect 4846 1787 4852 1788
rect 4990 1792 4996 1793
rect 4990 1788 4991 1792
rect 4995 1788 4996 1792
rect 4990 1787 4996 1788
rect 5134 1792 5140 1793
rect 5134 1788 5135 1792
rect 5139 1788 5140 1792
rect 5134 1787 5140 1788
rect 5270 1792 5276 1793
rect 5270 1788 5271 1792
rect 5275 1788 5276 1792
rect 5270 1787 5276 1788
rect 5406 1792 5412 1793
rect 5406 1788 5407 1792
rect 5411 1788 5412 1792
rect 5406 1787 5412 1788
rect 5542 1792 5548 1793
rect 5542 1788 5543 1792
rect 5547 1788 5548 1792
rect 5542 1787 5548 1788
rect 5662 1791 5668 1792
rect 5662 1787 5663 1791
rect 5667 1787 5668 1791
rect 3838 1786 3844 1787
rect 5662 1786 5668 1787
rect 1934 1784 1940 1785
rect 1574 1783 1580 1784
rect 130 1773 136 1774
rect 110 1772 116 1773
rect 110 1768 111 1772
rect 115 1768 116 1772
rect 130 1769 131 1773
rect 135 1769 136 1773
rect 130 1768 136 1769
rect 346 1773 352 1774
rect 346 1769 347 1773
rect 351 1769 352 1773
rect 346 1768 352 1769
rect 562 1773 568 1774
rect 562 1769 563 1773
rect 567 1769 568 1773
rect 562 1768 568 1769
rect 770 1773 776 1774
rect 770 1769 771 1773
rect 775 1769 776 1773
rect 770 1768 776 1769
rect 970 1773 976 1774
rect 970 1769 971 1773
rect 975 1769 976 1773
rect 970 1768 976 1769
rect 1162 1773 1168 1774
rect 1162 1769 1163 1773
rect 1167 1769 1168 1773
rect 1162 1768 1168 1769
rect 1354 1773 1360 1774
rect 1354 1769 1355 1773
rect 1359 1769 1360 1773
rect 1354 1768 1360 1769
rect 1546 1773 1552 1774
rect 1546 1769 1547 1773
rect 1551 1769 1552 1773
rect 1546 1768 1552 1769
rect 1934 1772 1940 1773
rect 1934 1768 1935 1772
rect 1939 1768 1940 1772
rect 110 1767 116 1768
rect 1934 1767 1940 1768
rect 1974 1725 1980 1726
rect 3798 1725 3804 1726
rect 1974 1721 1975 1725
rect 1979 1721 1980 1725
rect 1974 1720 1980 1721
rect 2022 1724 2028 1725
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2310 1724 2316 1725
rect 2310 1720 2311 1724
rect 2315 1720 2316 1724
rect 2310 1719 2316 1720
rect 2470 1724 2476 1725
rect 2470 1720 2471 1724
rect 2475 1720 2476 1724
rect 2470 1719 2476 1720
rect 2638 1724 2644 1725
rect 2638 1720 2639 1724
rect 2643 1720 2644 1724
rect 2638 1719 2644 1720
rect 2806 1724 2812 1725
rect 2806 1720 2807 1724
rect 2811 1720 2812 1724
rect 2806 1719 2812 1720
rect 2974 1724 2980 1725
rect 2974 1720 2975 1724
rect 2979 1720 2980 1724
rect 2974 1719 2980 1720
rect 3150 1724 3156 1725
rect 3150 1720 3151 1724
rect 3155 1720 3156 1724
rect 3798 1721 3799 1725
rect 3803 1721 3804 1725
rect 3798 1720 3804 1721
rect 3150 1719 3156 1720
rect 3838 1717 3844 1718
rect 5662 1717 5668 1718
rect 3838 1713 3839 1717
rect 3843 1713 3844 1717
rect 3838 1712 3844 1713
rect 3886 1716 3892 1717
rect 3886 1712 3887 1716
rect 3891 1712 3892 1716
rect 3886 1711 3892 1712
rect 4078 1716 4084 1717
rect 4078 1712 4079 1716
rect 4083 1712 4084 1716
rect 4078 1711 4084 1712
rect 4302 1716 4308 1717
rect 4302 1712 4303 1716
rect 4307 1712 4308 1716
rect 4302 1711 4308 1712
rect 4534 1716 4540 1717
rect 4534 1712 4535 1716
rect 4539 1712 4540 1716
rect 4534 1711 4540 1712
rect 4774 1716 4780 1717
rect 4774 1712 4775 1716
rect 4779 1712 4780 1716
rect 4774 1711 4780 1712
rect 5022 1716 5028 1717
rect 5022 1712 5023 1716
rect 5027 1712 5028 1716
rect 5022 1711 5028 1712
rect 5278 1716 5284 1717
rect 5278 1712 5279 1716
rect 5283 1712 5284 1716
rect 5278 1711 5284 1712
rect 5534 1716 5540 1717
rect 5534 1712 5535 1716
rect 5539 1712 5540 1716
rect 5662 1713 5663 1717
rect 5667 1713 5668 1717
rect 5662 1712 5668 1713
rect 5534 1711 5540 1712
rect 1994 1709 2000 1710
rect 1974 1708 1980 1709
rect 1974 1704 1975 1708
rect 1979 1704 1980 1708
rect 1994 1705 1995 1709
rect 1999 1705 2000 1709
rect 1994 1704 2000 1705
rect 2130 1709 2136 1710
rect 2130 1705 2131 1709
rect 2135 1705 2136 1709
rect 2130 1704 2136 1705
rect 2282 1709 2288 1710
rect 2282 1705 2283 1709
rect 2287 1705 2288 1709
rect 2282 1704 2288 1705
rect 2442 1709 2448 1710
rect 2442 1705 2443 1709
rect 2447 1705 2448 1709
rect 2442 1704 2448 1705
rect 2610 1709 2616 1710
rect 2610 1705 2611 1709
rect 2615 1705 2616 1709
rect 2610 1704 2616 1705
rect 2778 1709 2784 1710
rect 2778 1705 2779 1709
rect 2783 1705 2784 1709
rect 2778 1704 2784 1705
rect 2946 1709 2952 1710
rect 2946 1705 2947 1709
rect 2951 1705 2952 1709
rect 2946 1704 2952 1705
rect 3122 1709 3128 1710
rect 3122 1705 3123 1709
rect 3127 1705 3128 1709
rect 3122 1704 3128 1705
rect 3798 1708 3804 1709
rect 3798 1704 3799 1708
rect 3803 1704 3804 1708
rect 1974 1703 1980 1704
rect 3798 1703 3804 1704
rect 3858 1701 3864 1702
rect 3838 1700 3844 1701
rect 3838 1696 3839 1700
rect 3843 1696 3844 1700
rect 3858 1697 3859 1701
rect 3863 1697 3864 1701
rect 3858 1696 3864 1697
rect 4050 1701 4056 1702
rect 4050 1697 4051 1701
rect 4055 1697 4056 1701
rect 4050 1696 4056 1697
rect 4274 1701 4280 1702
rect 4274 1697 4275 1701
rect 4279 1697 4280 1701
rect 4274 1696 4280 1697
rect 4506 1701 4512 1702
rect 4506 1697 4507 1701
rect 4511 1697 4512 1701
rect 4506 1696 4512 1697
rect 4746 1701 4752 1702
rect 4746 1697 4747 1701
rect 4751 1697 4752 1701
rect 4746 1696 4752 1697
rect 4994 1701 5000 1702
rect 4994 1697 4995 1701
rect 4999 1697 5000 1701
rect 4994 1696 5000 1697
rect 5250 1701 5256 1702
rect 5250 1697 5251 1701
rect 5255 1697 5256 1701
rect 5250 1696 5256 1697
rect 5506 1701 5512 1702
rect 5506 1697 5507 1701
rect 5511 1697 5512 1701
rect 5506 1696 5512 1697
rect 5662 1700 5668 1701
rect 5662 1696 5663 1700
rect 5667 1696 5668 1700
rect 3838 1695 3844 1696
rect 5662 1695 5668 1696
rect 110 1616 116 1617
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 394 1615 400 1616
rect 394 1611 395 1615
rect 399 1611 400 1615
rect 394 1610 400 1611
rect 682 1615 688 1616
rect 682 1611 683 1615
rect 687 1611 688 1615
rect 682 1610 688 1611
rect 978 1615 984 1616
rect 978 1611 979 1615
rect 983 1611 984 1615
rect 978 1610 984 1611
rect 1274 1615 1280 1616
rect 1274 1611 1275 1615
rect 1279 1611 1280 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1274 1610 1280 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 422 1600 428 1601
rect 422 1596 423 1600
rect 427 1596 428 1600
rect 422 1595 428 1596
rect 710 1600 716 1601
rect 710 1596 711 1600
rect 715 1596 716 1600
rect 710 1595 716 1596
rect 1006 1600 1012 1601
rect 1006 1596 1007 1600
rect 1011 1596 1012 1600
rect 1006 1595 1012 1596
rect 1302 1600 1308 1601
rect 1302 1596 1303 1600
rect 1307 1596 1308 1600
rect 1302 1595 1308 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 1934 1594 1940 1595
rect 1974 1568 1980 1569
rect 3798 1568 3804 1569
rect 1974 1564 1975 1568
rect 1979 1564 1980 1568
rect 1974 1563 1980 1564
rect 2090 1567 2096 1568
rect 2090 1563 2091 1567
rect 2095 1563 2096 1567
rect 2090 1562 2096 1563
rect 2226 1567 2232 1568
rect 2226 1563 2227 1567
rect 2231 1563 2232 1567
rect 2226 1562 2232 1563
rect 2362 1567 2368 1568
rect 2362 1563 2363 1567
rect 2367 1563 2368 1567
rect 2362 1562 2368 1563
rect 2498 1567 2504 1568
rect 2498 1563 2499 1567
rect 2503 1563 2504 1567
rect 2498 1562 2504 1563
rect 2634 1567 2640 1568
rect 2634 1563 2635 1567
rect 2639 1563 2640 1567
rect 2634 1562 2640 1563
rect 2770 1567 2776 1568
rect 2770 1563 2771 1567
rect 2775 1563 2776 1567
rect 2770 1562 2776 1563
rect 2906 1567 2912 1568
rect 2906 1563 2907 1567
rect 2911 1563 2912 1567
rect 2906 1562 2912 1563
rect 3042 1567 3048 1568
rect 3042 1563 3043 1567
rect 3047 1563 3048 1567
rect 3042 1562 3048 1563
rect 3178 1567 3184 1568
rect 3178 1563 3179 1567
rect 3183 1563 3184 1567
rect 3798 1564 3799 1568
rect 3803 1564 3804 1568
rect 3798 1563 3804 1564
rect 3838 1568 3844 1569
rect 5662 1568 5668 1569
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3858 1567 3864 1568
rect 3858 1563 3859 1567
rect 3863 1563 3864 1567
rect 3178 1562 3184 1563
rect 3858 1562 3864 1563
rect 3994 1567 4000 1568
rect 3994 1563 3995 1567
rect 3999 1563 4000 1567
rect 3994 1562 4000 1563
rect 4154 1567 4160 1568
rect 4154 1563 4155 1567
rect 4159 1563 4160 1567
rect 4154 1562 4160 1563
rect 4354 1567 4360 1568
rect 4354 1563 4355 1567
rect 4359 1563 4360 1567
rect 4354 1562 4360 1563
rect 4586 1567 4592 1568
rect 4586 1563 4587 1567
rect 4591 1563 4592 1567
rect 4586 1562 4592 1563
rect 4850 1567 4856 1568
rect 4850 1563 4851 1567
rect 4855 1563 4856 1567
rect 4850 1562 4856 1563
rect 5130 1567 5136 1568
rect 5130 1563 5131 1567
rect 5135 1563 5136 1567
rect 5130 1562 5136 1563
rect 5418 1567 5424 1568
rect 5418 1563 5419 1567
rect 5423 1563 5424 1567
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5418 1562 5424 1563
rect 2118 1552 2124 1553
rect 1974 1551 1980 1552
rect 1974 1547 1975 1551
rect 1979 1547 1980 1551
rect 2118 1548 2119 1552
rect 2123 1548 2124 1552
rect 2118 1547 2124 1548
rect 2254 1552 2260 1553
rect 2254 1548 2255 1552
rect 2259 1548 2260 1552
rect 2254 1547 2260 1548
rect 2390 1552 2396 1553
rect 2390 1548 2391 1552
rect 2395 1548 2396 1552
rect 2390 1547 2396 1548
rect 2526 1552 2532 1553
rect 2526 1548 2527 1552
rect 2531 1548 2532 1552
rect 2526 1547 2532 1548
rect 2662 1552 2668 1553
rect 2662 1548 2663 1552
rect 2667 1548 2668 1552
rect 2662 1547 2668 1548
rect 2798 1552 2804 1553
rect 2798 1548 2799 1552
rect 2803 1548 2804 1552
rect 2798 1547 2804 1548
rect 2934 1552 2940 1553
rect 2934 1548 2935 1552
rect 2939 1548 2940 1552
rect 2934 1547 2940 1548
rect 3070 1552 3076 1553
rect 3070 1548 3071 1552
rect 3075 1548 3076 1552
rect 3070 1547 3076 1548
rect 3206 1552 3212 1553
rect 3886 1552 3892 1553
rect 3206 1548 3207 1552
rect 3211 1548 3212 1552
rect 3206 1547 3212 1548
rect 3798 1551 3804 1552
rect 3798 1547 3799 1551
rect 3803 1547 3804 1551
rect 1974 1546 1980 1547
rect 3798 1546 3804 1547
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3886 1548 3887 1552
rect 3891 1548 3892 1552
rect 3886 1547 3892 1548
rect 4022 1552 4028 1553
rect 4022 1548 4023 1552
rect 4027 1548 4028 1552
rect 4022 1547 4028 1548
rect 4182 1552 4188 1553
rect 4182 1548 4183 1552
rect 4187 1548 4188 1552
rect 4182 1547 4188 1548
rect 4382 1552 4388 1553
rect 4382 1548 4383 1552
rect 4387 1548 4388 1552
rect 4382 1547 4388 1548
rect 4614 1552 4620 1553
rect 4614 1548 4615 1552
rect 4619 1548 4620 1552
rect 4614 1547 4620 1548
rect 4878 1552 4884 1553
rect 4878 1548 4879 1552
rect 4883 1548 4884 1552
rect 4878 1547 4884 1548
rect 5158 1552 5164 1553
rect 5158 1548 5159 1552
rect 5163 1548 5164 1552
rect 5158 1547 5164 1548
rect 5446 1552 5452 1553
rect 5446 1548 5447 1552
rect 5451 1548 5452 1552
rect 5446 1547 5452 1548
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 3838 1546 3844 1547
rect 5662 1546 5668 1547
rect 110 1529 116 1530
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 374 1528 380 1529
rect 374 1524 375 1528
rect 379 1524 380 1528
rect 374 1523 380 1524
rect 606 1528 612 1529
rect 606 1524 607 1528
rect 611 1524 612 1528
rect 606 1523 612 1524
rect 838 1528 844 1529
rect 838 1524 839 1528
rect 843 1524 844 1528
rect 838 1523 844 1524
rect 1070 1528 1076 1529
rect 1070 1524 1071 1528
rect 1075 1524 1076 1528
rect 1070 1523 1076 1524
rect 1302 1528 1308 1529
rect 1302 1524 1303 1528
rect 1307 1524 1308 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1302 1523 1308 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 346 1513 352 1514
rect 346 1509 347 1513
rect 351 1509 352 1513
rect 346 1508 352 1509
rect 578 1513 584 1514
rect 578 1509 579 1513
rect 583 1509 584 1513
rect 578 1508 584 1509
rect 810 1513 816 1514
rect 810 1509 811 1513
rect 815 1509 816 1513
rect 810 1508 816 1509
rect 1042 1513 1048 1514
rect 1042 1509 1043 1513
rect 1047 1509 1048 1513
rect 1042 1508 1048 1509
rect 1274 1513 1280 1514
rect 1274 1509 1275 1513
rect 1279 1509 1280 1513
rect 1274 1508 1280 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 1934 1507 1940 1508
rect 3838 1493 3844 1494
rect 5662 1493 5668 1494
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 4302 1492 4308 1493
rect 4302 1488 4303 1492
rect 4307 1488 4308 1492
rect 4302 1487 4308 1488
rect 4494 1492 4500 1493
rect 4494 1488 4495 1492
rect 4499 1488 4500 1492
rect 4494 1487 4500 1488
rect 4718 1492 4724 1493
rect 4718 1488 4719 1492
rect 4723 1488 4724 1492
rect 4718 1487 4724 1488
rect 4966 1492 4972 1493
rect 4966 1488 4967 1492
rect 4971 1488 4972 1492
rect 4966 1487 4972 1488
rect 5222 1492 5228 1493
rect 5222 1488 5223 1492
rect 5227 1488 5228 1492
rect 5222 1487 5228 1488
rect 5486 1492 5492 1493
rect 5486 1488 5487 1492
rect 5491 1488 5492 1492
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5486 1487 5492 1488
rect 3858 1477 3864 1478
rect 3838 1476 3844 1477
rect 1974 1473 1980 1474
rect 3798 1473 3804 1474
rect 1974 1469 1975 1473
rect 1979 1469 1980 1473
rect 1974 1468 1980 1469
rect 2022 1472 2028 1473
rect 2022 1468 2023 1472
rect 2027 1468 2028 1472
rect 2022 1467 2028 1468
rect 2158 1472 2164 1473
rect 2158 1468 2159 1472
rect 2163 1468 2164 1472
rect 2158 1467 2164 1468
rect 2294 1472 2300 1473
rect 2294 1468 2295 1472
rect 2299 1468 2300 1472
rect 2294 1467 2300 1468
rect 2430 1472 2436 1473
rect 2430 1468 2431 1472
rect 2435 1468 2436 1472
rect 2430 1467 2436 1468
rect 2566 1472 2572 1473
rect 2566 1468 2567 1472
rect 2571 1468 2572 1472
rect 2566 1467 2572 1468
rect 2702 1472 2708 1473
rect 2702 1468 2703 1472
rect 2707 1468 2708 1472
rect 2702 1467 2708 1468
rect 2838 1472 2844 1473
rect 2838 1468 2839 1472
rect 2843 1468 2844 1472
rect 2838 1467 2844 1468
rect 2974 1472 2980 1473
rect 2974 1468 2975 1472
rect 2979 1468 2980 1472
rect 3798 1469 3799 1473
rect 3803 1469 3804 1473
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 4274 1477 4280 1478
rect 4274 1473 4275 1477
rect 4279 1473 4280 1477
rect 4274 1472 4280 1473
rect 4466 1477 4472 1478
rect 4466 1473 4467 1477
rect 4471 1473 4472 1477
rect 4466 1472 4472 1473
rect 4690 1477 4696 1478
rect 4690 1473 4691 1477
rect 4695 1473 4696 1477
rect 4690 1472 4696 1473
rect 4938 1477 4944 1478
rect 4938 1473 4939 1477
rect 4943 1473 4944 1477
rect 4938 1472 4944 1473
rect 5194 1477 5200 1478
rect 5194 1473 5195 1477
rect 5199 1473 5200 1477
rect 5194 1472 5200 1473
rect 5458 1477 5464 1478
rect 5458 1473 5459 1477
rect 5463 1473 5464 1477
rect 5458 1472 5464 1473
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 3838 1471 3844 1472
rect 5662 1471 5668 1472
rect 3798 1468 3804 1469
rect 2974 1467 2980 1468
rect 1994 1457 2000 1458
rect 1974 1456 1980 1457
rect 1974 1452 1975 1456
rect 1979 1452 1980 1456
rect 1994 1453 1995 1457
rect 1999 1453 2000 1457
rect 1994 1452 2000 1453
rect 2130 1457 2136 1458
rect 2130 1453 2131 1457
rect 2135 1453 2136 1457
rect 2130 1452 2136 1453
rect 2266 1457 2272 1458
rect 2266 1453 2267 1457
rect 2271 1453 2272 1457
rect 2266 1452 2272 1453
rect 2402 1457 2408 1458
rect 2402 1453 2403 1457
rect 2407 1453 2408 1457
rect 2402 1452 2408 1453
rect 2538 1457 2544 1458
rect 2538 1453 2539 1457
rect 2543 1453 2544 1457
rect 2538 1452 2544 1453
rect 2674 1457 2680 1458
rect 2674 1453 2675 1457
rect 2679 1453 2680 1457
rect 2674 1452 2680 1453
rect 2810 1457 2816 1458
rect 2810 1453 2811 1457
rect 2815 1453 2816 1457
rect 2810 1452 2816 1453
rect 2946 1457 2952 1458
rect 2946 1453 2947 1457
rect 2951 1453 2952 1457
rect 2946 1452 2952 1453
rect 3798 1456 3804 1457
rect 3798 1452 3799 1456
rect 3803 1452 3804 1456
rect 1974 1451 1980 1452
rect 3798 1451 3804 1452
rect 110 1368 116 1369
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 410 1367 416 1368
rect 410 1363 411 1367
rect 415 1363 416 1367
rect 410 1362 416 1363
rect 738 1367 744 1368
rect 738 1363 739 1367
rect 743 1363 744 1367
rect 738 1362 744 1363
rect 1090 1367 1096 1368
rect 1090 1363 1091 1367
rect 1095 1363 1096 1367
rect 1090 1362 1096 1363
rect 1450 1367 1456 1368
rect 1450 1363 1451 1367
rect 1455 1363 1456 1367
rect 1450 1362 1456 1363
rect 1786 1367 1792 1368
rect 1786 1363 1787 1367
rect 1791 1363 1792 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1786 1362 1792 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 438 1352 444 1353
rect 438 1348 439 1352
rect 443 1348 444 1352
rect 438 1347 444 1348
rect 766 1352 772 1353
rect 766 1348 767 1352
rect 771 1348 772 1352
rect 766 1347 772 1348
rect 1118 1352 1124 1353
rect 1118 1348 1119 1352
rect 1123 1348 1124 1352
rect 1118 1347 1124 1348
rect 1478 1352 1484 1353
rect 1478 1348 1479 1352
rect 1483 1348 1484 1352
rect 1478 1347 1484 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 1934 1346 1940 1347
rect 3838 1340 3844 1341
rect 5662 1340 5668 1341
rect 3838 1336 3839 1340
rect 3843 1336 3844 1340
rect 3838 1335 3844 1336
rect 3858 1339 3864 1340
rect 3858 1335 3859 1339
rect 3863 1335 3864 1339
rect 3858 1334 3864 1335
rect 4058 1339 4064 1340
rect 4058 1335 4059 1339
rect 4063 1335 4064 1339
rect 4058 1334 4064 1335
rect 4306 1339 4312 1340
rect 4306 1335 4307 1339
rect 4311 1335 4312 1339
rect 4306 1334 4312 1335
rect 4578 1339 4584 1340
rect 4578 1335 4579 1339
rect 4583 1335 4584 1339
rect 4578 1334 4584 1335
rect 4874 1339 4880 1340
rect 4874 1335 4875 1339
rect 4879 1335 4880 1339
rect 4874 1334 4880 1335
rect 5186 1339 5192 1340
rect 5186 1335 5187 1339
rect 5191 1335 5192 1339
rect 5186 1334 5192 1335
rect 5498 1339 5504 1340
rect 5498 1335 5499 1339
rect 5503 1335 5504 1339
rect 5662 1336 5663 1340
rect 5667 1336 5668 1340
rect 5662 1335 5668 1336
rect 5498 1334 5504 1335
rect 3886 1324 3892 1325
rect 3838 1323 3844 1324
rect 3838 1319 3839 1323
rect 3843 1319 3844 1323
rect 3886 1320 3887 1324
rect 3891 1320 3892 1324
rect 3886 1319 3892 1320
rect 4086 1324 4092 1325
rect 4086 1320 4087 1324
rect 4091 1320 4092 1324
rect 4086 1319 4092 1320
rect 4334 1324 4340 1325
rect 4334 1320 4335 1324
rect 4339 1320 4340 1324
rect 4334 1319 4340 1320
rect 4606 1324 4612 1325
rect 4606 1320 4607 1324
rect 4611 1320 4612 1324
rect 4606 1319 4612 1320
rect 4902 1324 4908 1325
rect 4902 1320 4903 1324
rect 4907 1320 4908 1324
rect 4902 1319 4908 1320
rect 5214 1324 5220 1325
rect 5214 1320 5215 1324
rect 5219 1320 5220 1324
rect 5214 1319 5220 1320
rect 5526 1324 5532 1325
rect 5526 1320 5527 1324
rect 5531 1320 5532 1324
rect 5526 1319 5532 1320
rect 5662 1323 5668 1324
rect 5662 1319 5663 1323
rect 5667 1319 5668 1323
rect 3838 1318 3844 1319
rect 5662 1318 5668 1319
rect 1974 1316 1980 1317
rect 3798 1316 3804 1317
rect 1974 1312 1975 1316
rect 1979 1312 1980 1316
rect 1974 1311 1980 1312
rect 1994 1315 2000 1316
rect 1994 1311 1995 1315
rect 1999 1311 2000 1315
rect 1994 1310 2000 1311
rect 2274 1315 2280 1316
rect 2274 1311 2275 1315
rect 2279 1311 2280 1315
rect 2274 1310 2280 1311
rect 2562 1315 2568 1316
rect 2562 1311 2563 1315
rect 2567 1311 2568 1315
rect 2562 1310 2568 1311
rect 2842 1315 2848 1316
rect 2842 1311 2843 1315
rect 2847 1311 2848 1315
rect 2842 1310 2848 1311
rect 3122 1315 3128 1316
rect 3122 1311 3123 1315
rect 3127 1311 3128 1315
rect 3122 1310 3128 1311
rect 3394 1315 3400 1316
rect 3394 1311 3395 1315
rect 3399 1311 3400 1315
rect 3394 1310 3400 1311
rect 3650 1315 3656 1316
rect 3650 1311 3651 1315
rect 3655 1311 3656 1315
rect 3798 1312 3799 1316
rect 3803 1312 3804 1316
rect 3798 1311 3804 1312
rect 3650 1310 3656 1311
rect 2022 1300 2028 1301
rect 1974 1299 1980 1300
rect 1974 1295 1975 1299
rect 1979 1295 1980 1299
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2302 1300 2308 1301
rect 2302 1296 2303 1300
rect 2307 1296 2308 1300
rect 2302 1295 2308 1296
rect 2590 1300 2596 1301
rect 2590 1296 2591 1300
rect 2595 1296 2596 1300
rect 2590 1295 2596 1296
rect 2870 1300 2876 1301
rect 2870 1296 2871 1300
rect 2875 1296 2876 1300
rect 2870 1295 2876 1296
rect 3150 1300 3156 1301
rect 3150 1296 3151 1300
rect 3155 1296 3156 1300
rect 3150 1295 3156 1296
rect 3422 1300 3428 1301
rect 3422 1296 3423 1300
rect 3427 1296 3428 1300
rect 3422 1295 3428 1296
rect 3678 1300 3684 1301
rect 3678 1296 3679 1300
rect 3683 1296 3684 1300
rect 3678 1295 3684 1296
rect 3798 1299 3804 1300
rect 3798 1295 3799 1299
rect 3803 1295 3804 1299
rect 1974 1294 1980 1295
rect 3798 1294 3804 1295
rect 110 1293 116 1294
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 358 1292 364 1293
rect 358 1288 359 1292
rect 363 1288 364 1292
rect 358 1287 364 1288
rect 574 1292 580 1293
rect 574 1288 575 1292
rect 579 1288 580 1292
rect 574 1287 580 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 966 1292 972 1293
rect 966 1288 967 1292
rect 971 1288 972 1292
rect 966 1287 972 1288
rect 1150 1292 1156 1293
rect 1150 1288 1151 1292
rect 1155 1288 1156 1292
rect 1150 1287 1156 1288
rect 1326 1292 1332 1293
rect 1326 1288 1327 1292
rect 1331 1288 1332 1292
rect 1326 1287 1332 1288
rect 1494 1292 1500 1293
rect 1494 1288 1495 1292
rect 1499 1288 1500 1292
rect 1494 1287 1500 1288
rect 1662 1292 1668 1293
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 330 1277 336 1278
rect 330 1273 331 1277
rect 335 1273 336 1277
rect 330 1272 336 1273
rect 546 1277 552 1278
rect 546 1273 547 1277
rect 551 1273 552 1277
rect 546 1272 552 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 938 1277 944 1278
rect 938 1273 939 1277
rect 943 1273 944 1277
rect 938 1272 944 1273
rect 1122 1277 1128 1278
rect 1122 1273 1123 1277
rect 1127 1273 1128 1277
rect 1122 1272 1128 1273
rect 1298 1277 1304 1278
rect 1298 1273 1299 1277
rect 1303 1273 1304 1277
rect 1298 1272 1304 1273
rect 1466 1277 1472 1278
rect 1466 1273 1467 1277
rect 1471 1273 1472 1277
rect 1466 1272 1472 1273
rect 1634 1277 1640 1278
rect 1634 1273 1635 1277
rect 1639 1273 1640 1277
rect 1634 1272 1640 1273
rect 1786 1277 1792 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 1934 1271 1940 1272
rect 3838 1257 3844 1258
rect 5662 1257 5668 1258
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4614 1256 4620 1257
rect 4614 1252 4615 1256
rect 4619 1252 4620 1256
rect 4614 1251 4620 1252
rect 4790 1256 4796 1257
rect 4790 1252 4791 1256
rect 4795 1252 4796 1256
rect 4790 1251 4796 1252
rect 4974 1256 4980 1257
rect 4974 1252 4975 1256
rect 4979 1252 4980 1256
rect 4974 1251 4980 1252
rect 5166 1256 5172 1257
rect 5166 1252 5167 1256
rect 5171 1252 5172 1256
rect 5166 1251 5172 1252
rect 5366 1256 5372 1257
rect 5366 1252 5367 1256
rect 5371 1252 5372 1256
rect 5366 1251 5372 1252
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5542 1251 5548 1252
rect 4586 1241 4592 1242
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4586 1237 4587 1241
rect 4591 1237 4592 1241
rect 4586 1236 4592 1237
rect 4762 1241 4768 1242
rect 4762 1237 4763 1241
rect 4767 1237 4768 1241
rect 4762 1236 4768 1237
rect 4946 1241 4952 1242
rect 4946 1237 4947 1241
rect 4951 1237 4952 1241
rect 4946 1236 4952 1237
rect 5138 1241 5144 1242
rect 5138 1237 5139 1241
rect 5143 1237 5144 1241
rect 5138 1236 5144 1237
rect 5338 1241 5344 1242
rect 5338 1237 5339 1241
rect 5343 1237 5344 1241
rect 5338 1236 5344 1237
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 5662 1235 5668 1236
rect 1974 1217 1980 1218
rect 3798 1217 3804 1218
rect 1974 1213 1975 1217
rect 1979 1213 1980 1217
rect 1974 1212 1980 1213
rect 2654 1216 2660 1217
rect 2654 1212 2655 1216
rect 2659 1212 2660 1216
rect 2654 1211 2660 1212
rect 2830 1216 2836 1217
rect 2830 1212 2831 1216
rect 2835 1212 2836 1216
rect 2830 1211 2836 1212
rect 3006 1216 3012 1217
rect 3006 1212 3007 1216
rect 3011 1212 3012 1216
rect 3006 1211 3012 1212
rect 3182 1216 3188 1217
rect 3182 1212 3183 1216
rect 3187 1212 3188 1216
rect 3182 1211 3188 1212
rect 3358 1216 3364 1217
rect 3358 1212 3359 1216
rect 3363 1212 3364 1216
rect 3358 1211 3364 1212
rect 3542 1216 3548 1217
rect 3542 1212 3543 1216
rect 3547 1212 3548 1216
rect 3798 1213 3799 1217
rect 3803 1213 3804 1217
rect 3798 1212 3804 1213
rect 3542 1211 3548 1212
rect 2626 1201 2632 1202
rect 1974 1200 1980 1201
rect 1974 1196 1975 1200
rect 1979 1196 1980 1200
rect 2626 1197 2627 1201
rect 2631 1197 2632 1201
rect 2626 1196 2632 1197
rect 2802 1201 2808 1202
rect 2802 1197 2803 1201
rect 2807 1197 2808 1201
rect 2802 1196 2808 1197
rect 2978 1201 2984 1202
rect 2978 1197 2979 1201
rect 2983 1197 2984 1201
rect 2978 1196 2984 1197
rect 3154 1201 3160 1202
rect 3154 1197 3155 1201
rect 3159 1197 3160 1201
rect 3154 1196 3160 1197
rect 3330 1201 3336 1202
rect 3330 1197 3331 1201
rect 3335 1197 3336 1201
rect 3330 1196 3336 1197
rect 3514 1201 3520 1202
rect 3514 1197 3515 1201
rect 3519 1197 3520 1201
rect 3514 1196 3520 1197
rect 3798 1200 3804 1201
rect 3798 1196 3799 1200
rect 3803 1196 3804 1200
rect 1974 1195 1980 1196
rect 3798 1195 3804 1196
rect 110 1132 116 1133
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 290 1131 296 1132
rect 290 1127 291 1131
rect 295 1127 296 1131
rect 290 1126 296 1127
rect 474 1131 480 1132
rect 474 1127 475 1131
rect 479 1127 480 1131
rect 474 1126 480 1127
rect 658 1131 664 1132
rect 658 1127 659 1131
rect 663 1127 664 1131
rect 658 1126 664 1127
rect 834 1131 840 1132
rect 834 1127 835 1131
rect 839 1127 840 1131
rect 834 1126 840 1127
rect 1002 1131 1008 1132
rect 1002 1127 1003 1131
rect 1007 1127 1008 1131
rect 1002 1126 1008 1127
rect 1170 1131 1176 1132
rect 1170 1127 1171 1131
rect 1175 1127 1176 1131
rect 1170 1126 1176 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1490 1131 1496 1132
rect 1490 1127 1491 1131
rect 1495 1127 1496 1131
rect 1490 1126 1496 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 158 1116 164 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 318 1116 324 1117
rect 318 1112 319 1116
rect 323 1112 324 1116
rect 318 1111 324 1112
rect 502 1116 508 1117
rect 502 1112 503 1116
rect 507 1112 508 1116
rect 502 1111 508 1112
rect 686 1116 692 1117
rect 686 1112 687 1116
rect 691 1112 692 1116
rect 686 1111 692 1112
rect 862 1116 868 1117
rect 862 1112 863 1116
rect 867 1112 868 1116
rect 862 1111 868 1112
rect 1030 1116 1036 1117
rect 1030 1112 1031 1116
rect 1035 1112 1036 1116
rect 1030 1111 1036 1112
rect 1198 1116 1204 1117
rect 1198 1112 1199 1116
rect 1203 1112 1204 1116
rect 1198 1111 1204 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1518 1116 1524 1117
rect 1518 1112 1519 1116
rect 1523 1112 1524 1116
rect 1518 1111 1524 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 110 1110 116 1111
rect 1934 1110 1940 1111
rect 3838 1104 3844 1105
rect 5662 1104 5668 1105
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4834 1103 4840 1104
rect 4834 1099 4835 1103
rect 4839 1099 4840 1103
rect 4834 1098 4840 1099
rect 4970 1103 4976 1104
rect 4970 1099 4971 1103
rect 4975 1099 4976 1103
rect 4970 1098 4976 1099
rect 5106 1103 5112 1104
rect 5106 1099 5107 1103
rect 5111 1099 5112 1103
rect 5106 1098 5112 1099
rect 5242 1103 5248 1104
rect 5242 1099 5243 1103
rect 5247 1099 5248 1103
rect 5242 1098 5248 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5514 1098 5520 1099
rect 4862 1088 4868 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4862 1084 4863 1088
rect 4867 1084 4868 1088
rect 4862 1083 4868 1084
rect 4998 1088 5004 1089
rect 4998 1084 4999 1088
rect 5003 1084 5004 1088
rect 4998 1083 5004 1084
rect 5134 1088 5140 1089
rect 5134 1084 5135 1088
rect 5139 1084 5140 1088
rect 5134 1083 5140 1084
rect 5270 1088 5276 1089
rect 5270 1084 5271 1088
rect 5275 1084 5276 1088
rect 5270 1083 5276 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 3838 1082 3844 1083
rect 5662 1082 5668 1083
rect 1974 1052 1980 1053
rect 3798 1052 3804 1053
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 1994 1051 2000 1052
rect 1994 1047 1995 1051
rect 1999 1047 2000 1051
rect 1994 1046 2000 1047
rect 2170 1051 2176 1052
rect 2170 1047 2171 1051
rect 2175 1047 2176 1051
rect 2170 1046 2176 1047
rect 2362 1051 2368 1052
rect 2362 1047 2363 1051
rect 2367 1047 2368 1051
rect 2362 1046 2368 1047
rect 2546 1051 2552 1052
rect 2546 1047 2547 1051
rect 2551 1047 2552 1051
rect 2546 1046 2552 1047
rect 2722 1051 2728 1052
rect 2722 1047 2723 1051
rect 2727 1047 2728 1051
rect 2722 1046 2728 1047
rect 2890 1051 2896 1052
rect 2890 1047 2891 1051
rect 2895 1047 2896 1051
rect 2890 1046 2896 1047
rect 3058 1051 3064 1052
rect 3058 1047 3059 1051
rect 3063 1047 3064 1051
rect 3058 1046 3064 1047
rect 3218 1051 3224 1052
rect 3218 1047 3219 1051
rect 3223 1047 3224 1051
rect 3218 1046 3224 1047
rect 3386 1051 3392 1052
rect 3386 1047 3387 1051
rect 3391 1047 3392 1051
rect 3798 1048 3799 1052
rect 3803 1048 3804 1052
rect 3798 1047 3804 1048
rect 3386 1046 3392 1047
rect 110 1045 116 1046
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 174 1044 180 1045
rect 174 1040 175 1044
rect 179 1040 180 1044
rect 174 1039 180 1040
rect 430 1044 436 1045
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 686 1044 692 1045
rect 686 1040 687 1044
rect 691 1040 692 1044
rect 686 1039 692 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1214 1044 1220 1045
rect 1214 1040 1215 1044
rect 1219 1040 1220 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1214 1039 1220 1040
rect 2022 1036 2028 1037
rect 1974 1035 1980 1036
rect 1974 1031 1975 1035
rect 1979 1031 1980 1035
rect 2022 1032 2023 1036
rect 2027 1032 2028 1036
rect 2022 1031 2028 1032
rect 2198 1036 2204 1037
rect 2198 1032 2199 1036
rect 2203 1032 2204 1036
rect 2198 1031 2204 1032
rect 2390 1036 2396 1037
rect 2390 1032 2391 1036
rect 2395 1032 2396 1036
rect 2390 1031 2396 1032
rect 2574 1036 2580 1037
rect 2574 1032 2575 1036
rect 2579 1032 2580 1036
rect 2574 1031 2580 1032
rect 2750 1036 2756 1037
rect 2750 1032 2751 1036
rect 2755 1032 2756 1036
rect 2750 1031 2756 1032
rect 2918 1036 2924 1037
rect 2918 1032 2919 1036
rect 2923 1032 2924 1036
rect 2918 1031 2924 1032
rect 3086 1036 3092 1037
rect 3086 1032 3087 1036
rect 3091 1032 3092 1036
rect 3086 1031 3092 1032
rect 3246 1036 3252 1037
rect 3246 1032 3247 1036
rect 3251 1032 3252 1036
rect 3246 1031 3252 1032
rect 3414 1036 3420 1037
rect 3414 1032 3415 1036
rect 3419 1032 3420 1036
rect 3414 1031 3420 1032
rect 3798 1035 3804 1036
rect 3798 1031 3799 1035
rect 3803 1031 3804 1035
rect 1974 1030 1980 1031
rect 3798 1030 3804 1031
rect 146 1029 152 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 146 1025 147 1029
rect 151 1025 152 1029
rect 146 1024 152 1025
rect 402 1029 408 1030
rect 402 1025 403 1029
rect 407 1025 408 1029
rect 402 1024 408 1025
rect 658 1029 664 1030
rect 658 1025 659 1029
rect 663 1025 664 1029
rect 658 1024 664 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1186 1029 1192 1030
rect 1186 1025 1187 1029
rect 1191 1025 1192 1029
rect 1186 1024 1192 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 1934 1023 1940 1024
rect 3838 1025 3844 1026
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5486 1019 5492 1020
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 5662 1003 5668 1004
rect 1974 977 1980 978
rect 3798 977 3804 978
rect 1974 973 1975 977
rect 1979 973 1980 977
rect 1974 972 1980 973
rect 2022 976 2028 977
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 2190 976 2196 977
rect 2190 972 2191 976
rect 2195 972 2196 976
rect 2190 971 2196 972
rect 2374 976 2380 977
rect 2374 972 2375 976
rect 2379 972 2380 976
rect 2374 971 2380 972
rect 2566 976 2572 977
rect 2566 972 2567 976
rect 2571 972 2572 976
rect 2566 971 2572 972
rect 2758 976 2764 977
rect 2758 972 2759 976
rect 2763 972 2764 976
rect 2758 971 2764 972
rect 2942 976 2948 977
rect 2942 972 2943 976
rect 2947 972 2948 976
rect 2942 971 2948 972
rect 3126 976 3132 977
rect 3126 972 3127 976
rect 3131 972 3132 976
rect 3126 971 3132 972
rect 3310 976 3316 977
rect 3310 972 3311 976
rect 3315 972 3316 976
rect 3310 971 3316 972
rect 3494 976 3500 977
rect 3494 972 3495 976
rect 3499 972 3500 976
rect 3494 971 3500 972
rect 3678 976 3684 977
rect 3678 972 3679 976
rect 3683 972 3684 976
rect 3798 973 3799 977
rect 3803 973 3804 977
rect 3798 972 3804 973
rect 3678 971 3684 972
rect 1994 961 2000 962
rect 1974 960 1980 961
rect 1974 956 1975 960
rect 1979 956 1980 960
rect 1994 957 1995 961
rect 1999 957 2000 961
rect 1994 956 2000 957
rect 2162 961 2168 962
rect 2162 957 2163 961
rect 2167 957 2168 961
rect 2162 956 2168 957
rect 2346 961 2352 962
rect 2346 957 2347 961
rect 2351 957 2352 961
rect 2346 956 2352 957
rect 2538 961 2544 962
rect 2538 957 2539 961
rect 2543 957 2544 961
rect 2538 956 2544 957
rect 2730 961 2736 962
rect 2730 957 2731 961
rect 2735 957 2736 961
rect 2730 956 2736 957
rect 2914 961 2920 962
rect 2914 957 2915 961
rect 2919 957 2920 961
rect 2914 956 2920 957
rect 3098 961 3104 962
rect 3098 957 3099 961
rect 3103 957 3104 961
rect 3098 956 3104 957
rect 3282 961 3288 962
rect 3282 957 3283 961
rect 3287 957 3288 961
rect 3282 956 3288 957
rect 3466 961 3472 962
rect 3466 957 3467 961
rect 3471 957 3472 961
rect 3466 956 3472 957
rect 3650 961 3656 962
rect 3650 957 3651 961
rect 3655 957 3656 961
rect 3650 956 3656 957
rect 3798 960 3804 961
rect 3798 956 3799 960
rect 3803 956 3804 960
rect 1974 955 1980 956
rect 3798 955 3804 956
rect 110 884 116 885
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 234 883 240 884
rect 234 879 235 883
rect 239 879 240 883
rect 234 878 240 879
rect 458 883 464 884
rect 458 879 459 883
rect 463 879 464 883
rect 458 878 464 879
rect 682 883 688 884
rect 682 879 683 883
rect 687 879 688 883
rect 682 878 688 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1130 883 1136 884
rect 1130 879 1131 883
rect 1135 879 1136 883
rect 1130 878 1136 879
rect 1362 883 1368 884
rect 1362 879 1363 883
rect 1367 879 1368 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1362 878 1368 879
rect 3838 872 3844 873
rect 5662 872 5668 873
rect 262 868 268 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 262 864 263 868
rect 267 864 268 868
rect 262 863 268 864
rect 486 868 492 869
rect 486 864 487 868
rect 491 864 492 868
rect 486 863 492 864
rect 710 868 716 869
rect 710 864 711 868
rect 715 864 716 868
rect 710 863 716 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1158 868 1164 869
rect 1158 864 1159 868
rect 1163 864 1164 868
rect 1158 863 1164 864
rect 1390 868 1396 869
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 1390 864 1391 868
rect 1395 864 1396 868
rect 1390 863 1396 864
rect 1934 867 1940 868
rect 3838 867 3844 868
rect 3858 871 3864 872
rect 3858 867 3859 871
rect 3863 867 3864 871
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 3858 866 3864 867
rect 3994 871 4000 872
rect 3994 867 3995 871
rect 3999 867 4000 871
rect 3994 866 4000 867
rect 4170 871 4176 872
rect 4170 867 4171 871
rect 4175 867 4176 871
rect 4170 866 4176 867
rect 4386 871 4392 872
rect 4386 867 4387 871
rect 4391 867 4392 871
rect 4386 866 4392 867
rect 4642 871 4648 872
rect 4642 867 4643 871
rect 4647 867 4648 871
rect 4642 866 4648 867
rect 4930 871 4936 872
rect 4930 867 4931 871
rect 4935 867 4936 871
rect 4930 866 4936 867
rect 5234 871 5240 872
rect 5234 867 5235 871
rect 5239 867 5240 871
rect 5234 866 5240 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5514 866 5520 867
rect 110 862 116 863
rect 1934 862 1940 863
rect 3886 856 3892 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 3886 852 3887 856
rect 3891 852 3892 856
rect 3886 851 3892 852
rect 4022 856 4028 857
rect 4022 852 4023 856
rect 4027 852 4028 856
rect 4022 851 4028 852
rect 4198 856 4204 857
rect 4198 852 4199 856
rect 4203 852 4204 856
rect 4198 851 4204 852
rect 4414 856 4420 857
rect 4414 852 4415 856
rect 4419 852 4420 856
rect 4414 851 4420 852
rect 4670 856 4676 857
rect 4670 852 4671 856
rect 4675 852 4676 856
rect 4670 851 4676 852
rect 4958 856 4964 857
rect 4958 852 4959 856
rect 4963 852 4964 856
rect 4958 851 4964 852
rect 5262 856 5268 857
rect 5262 852 5263 856
rect 5267 852 5268 856
rect 5262 851 5268 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 3838 850 3844 851
rect 5662 850 5668 851
rect 1974 824 1980 825
rect 3798 824 3804 825
rect 1974 820 1975 824
rect 1979 820 1980 824
rect 1974 819 1980 820
rect 1994 823 2000 824
rect 1994 819 1995 823
rect 1999 819 2000 823
rect 1994 818 2000 819
rect 2178 823 2184 824
rect 2178 819 2179 823
rect 2183 819 2184 823
rect 2178 818 2184 819
rect 2402 823 2408 824
rect 2402 819 2403 823
rect 2407 819 2408 823
rect 2402 818 2408 819
rect 2674 823 2680 824
rect 2674 819 2675 823
rect 2679 819 2680 823
rect 2674 818 2680 819
rect 2986 823 2992 824
rect 2986 819 2987 823
rect 2991 819 2992 823
rect 2986 818 2992 819
rect 3322 823 3328 824
rect 3322 819 3323 823
rect 3327 819 3328 823
rect 3322 818 3328 819
rect 3650 823 3656 824
rect 3650 819 3651 823
rect 3655 819 3656 823
rect 3798 820 3799 824
rect 3803 820 3804 824
rect 3798 819 3804 820
rect 3650 818 3656 819
rect 2022 808 2028 809
rect 1974 807 1980 808
rect 1974 803 1975 807
rect 1979 803 1980 807
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2430 808 2436 809
rect 2430 804 2431 808
rect 2435 804 2436 808
rect 2430 803 2436 804
rect 2702 808 2708 809
rect 2702 804 2703 808
rect 2707 804 2708 808
rect 2702 803 2708 804
rect 3014 808 3020 809
rect 3014 804 3015 808
rect 3019 804 3020 808
rect 3014 803 3020 804
rect 3350 808 3356 809
rect 3350 804 3351 808
rect 3355 804 3356 808
rect 3350 803 3356 804
rect 3678 808 3684 809
rect 3678 804 3679 808
rect 3683 804 3684 808
rect 3678 803 3684 804
rect 3798 807 3804 808
rect 3798 803 3799 807
rect 3803 803 3804 807
rect 1974 802 1980 803
rect 3798 802 3804 803
rect 3838 797 3844 798
rect 5662 797 5668 798
rect 110 793 116 794
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 174 792 180 793
rect 174 788 175 792
rect 179 788 180 792
rect 174 787 180 788
rect 430 792 436 793
rect 430 788 431 792
rect 435 788 436 792
rect 430 787 436 788
rect 670 792 676 793
rect 670 788 671 792
rect 675 788 676 792
rect 670 787 676 788
rect 902 792 908 793
rect 902 788 903 792
rect 907 788 908 792
rect 902 787 908 788
rect 1126 792 1132 793
rect 1126 788 1127 792
rect 1131 788 1132 792
rect 1126 787 1132 788
rect 1350 792 1356 793
rect 1350 788 1351 792
rect 1355 788 1356 792
rect 1350 787 1356 788
rect 1574 792 1580 793
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3886 796 3892 797
rect 3886 792 3887 796
rect 3891 792 3892 796
rect 3886 791 3892 792
rect 4022 796 4028 797
rect 4022 792 4023 796
rect 4027 792 4028 796
rect 4022 791 4028 792
rect 4158 796 4164 797
rect 4158 792 4159 796
rect 4163 792 4164 796
rect 4158 791 4164 792
rect 4294 796 4300 797
rect 4294 792 4295 796
rect 4299 792 4300 796
rect 4294 791 4300 792
rect 4430 796 4436 797
rect 4430 792 4431 796
rect 4435 792 4436 796
rect 4430 791 4436 792
rect 4566 796 4572 797
rect 4566 792 4567 796
rect 4571 792 4572 796
rect 4566 791 4572 792
rect 4718 796 4724 797
rect 4718 792 4719 796
rect 4723 792 4724 796
rect 4718 791 4724 792
rect 4894 796 4900 797
rect 4894 792 4895 796
rect 4899 792 4900 796
rect 4894 791 4900 792
rect 5086 796 5092 797
rect 5086 792 5087 796
rect 5091 792 5092 796
rect 5086 791 5092 792
rect 5286 796 5292 797
rect 5286 792 5287 796
rect 5291 792 5292 796
rect 5286 791 5292 792
rect 5486 796 5492 797
rect 5486 792 5487 796
rect 5491 792 5492 796
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5486 791 5492 792
rect 1934 788 1940 789
rect 1574 787 1580 788
rect 3858 781 3864 782
rect 3838 780 3844 781
rect 146 777 152 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 146 773 147 777
rect 151 773 152 777
rect 146 772 152 773
rect 402 777 408 778
rect 402 773 403 777
rect 407 773 408 777
rect 402 772 408 773
rect 642 777 648 778
rect 642 773 643 777
rect 647 773 648 777
rect 642 772 648 773
rect 874 777 880 778
rect 874 773 875 777
rect 879 773 880 777
rect 874 772 880 773
rect 1098 777 1104 778
rect 1098 773 1099 777
rect 1103 773 1104 777
rect 1098 772 1104 773
rect 1322 777 1328 778
rect 1322 773 1323 777
rect 1327 773 1328 777
rect 1322 772 1328 773
rect 1546 777 1552 778
rect 1546 773 1547 777
rect 1551 773 1552 777
rect 1546 772 1552 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3858 777 3859 781
rect 3863 777 3864 781
rect 3858 776 3864 777
rect 3994 781 4000 782
rect 3994 777 3995 781
rect 3999 777 4000 781
rect 3994 776 4000 777
rect 4130 781 4136 782
rect 4130 777 4131 781
rect 4135 777 4136 781
rect 4130 776 4136 777
rect 4266 781 4272 782
rect 4266 777 4267 781
rect 4271 777 4272 781
rect 4266 776 4272 777
rect 4402 781 4408 782
rect 4402 777 4403 781
rect 4407 777 4408 781
rect 4402 776 4408 777
rect 4538 781 4544 782
rect 4538 777 4539 781
rect 4543 777 4544 781
rect 4538 776 4544 777
rect 4690 781 4696 782
rect 4690 777 4691 781
rect 4695 777 4696 781
rect 4690 776 4696 777
rect 4866 781 4872 782
rect 4866 777 4867 781
rect 4871 777 4872 781
rect 4866 776 4872 777
rect 5058 781 5064 782
rect 5058 777 5059 781
rect 5063 777 5064 781
rect 5058 776 5064 777
rect 5258 781 5264 782
rect 5258 777 5259 781
rect 5263 777 5264 781
rect 5258 776 5264 777
rect 5458 781 5464 782
rect 5458 777 5459 781
rect 5463 777 5464 781
rect 5458 776 5464 777
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 3838 775 3844 776
rect 5662 775 5668 776
rect 110 771 116 772
rect 1934 771 1940 772
rect 110 644 116 645
rect 1934 644 1940 645
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 314 643 320 644
rect 314 639 315 643
rect 319 639 320 643
rect 314 638 320 639
rect 522 643 528 644
rect 522 639 523 643
rect 527 639 528 643
rect 522 638 528 639
rect 722 643 728 644
rect 722 639 723 643
rect 727 639 728 643
rect 722 638 728 639
rect 906 643 912 644
rect 906 639 907 643
rect 911 639 912 643
rect 906 638 912 639
rect 1082 643 1088 644
rect 1082 639 1083 643
rect 1087 639 1088 643
rect 1082 638 1088 639
rect 1258 643 1264 644
rect 1258 639 1259 643
rect 1263 639 1264 643
rect 1258 638 1264 639
rect 1426 643 1432 644
rect 1426 639 1427 643
rect 1431 639 1432 643
rect 1426 638 1432 639
rect 1594 643 1600 644
rect 1594 639 1595 643
rect 1599 639 1600 643
rect 1594 638 1600 639
rect 1770 643 1776 644
rect 1770 639 1771 643
rect 1775 639 1776 643
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 3838 644 3844 645
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 1770 638 1776 639
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4698 643 4704 644
rect 4698 639 4699 643
rect 4703 639 4704 643
rect 4698 638 4704 639
rect 4890 643 4896 644
rect 4890 639 4891 643
rect 4895 639 4896 643
rect 4890 638 4896 639
rect 5098 643 5104 644
rect 5098 639 5099 643
rect 5103 639 5104 643
rect 5098 638 5104 639
rect 5314 643 5320 644
rect 5314 639 5315 643
rect 5319 639 5320 643
rect 5314 638 5320 639
rect 5514 643 5520 644
rect 5514 639 5515 643
rect 5519 639 5520 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5514 638 5520 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 342 628 348 629
rect 342 624 343 628
rect 347 624 348 628
rect 342 623 348 624
rect 550 628 556 629
rect 550 624 551 628
rect 555 624 556 628
rect 550 623 556 624
rect 750 628 756 629
rect 750 624 751 628
rect 755 624 756 628
rect 750 623 756 624
rect 934 628 940 629
rect 934 624 935 628
rect 939 624 940 628
rect 934 623 940 624
rect 1110 628 1116 629
rect 1110 624 1111 628
rect 1115 624 1116 628
rect 1110 623 1116 624
rect 1286 628 1292 629
rect 1286 624 1287 628
rect 1291 624 1292 628
rect 1286 623 1292 624
rect 1454 628 1460 629
rect 1454 624 1455 628
rect 1459 624 1460 628
rect 1454 623 1460 624
rect 1622 628 1628 629
rect 1622 624 1623 628
rect 1627 624 1628 628
rect 1622 623 1628 624
rect 1798 628 1804 629
rect 3886 628 3892 629
rect 1798 624 1799 628
rect 1803 624 1804 628
rect 1798 623 1804 624
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 110 622 116 623
rect 1934 622 1940 623
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4726 628 4732 629
rect 4726 624 4727 628
rect 4731 624 4732 628
rect 4726 623 4732 624
rect 4918 628 4924 629
rect 4918 624 4919 628
rect 4923 624 4924 628
rect 4918 623 4924 624
rect 5126 628 5132 629
rect 5126 624 5127 628
rect 5131 624 5132 628
rect 5126 623 5132 624
rect 5342 628 5348 629
rect 5342 624 5343 628
rect 5347 624 5348 628
rect 5342 623 5348 624
rect 5542 628 5548 629
rect 5542 624 5543 628
rect 5547 624 5548 628
rect 5542 623 5548 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 5662 622 5668 623
rect 110 569 116 570
rect 1934 569 1940 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 374 568 380 569
rect 374 564 375 568
rect 379 564 380 568
rect 374 563 380 564
rect 598 568 604 569
rect 598 564 599 568
rect 603 564 604 568
rect 598 563 604 564
rect 806 568 812 569
rect 806 564 807 568
rect 811 564 812 568
rect 806 563 812 564
rect 998 568 1004 569
rect 998 564 999 568
rect 1003 564 1004 568
rect 998 563 1004 564
rect 1174 568 1180 569
rect 1174 564 1175 568
rect 1179 564 1180 568
rect 1174 563 1180 564
rect 1342 568 1348 569
rect 1342 564 1343 568
rect 1347 564 1348 568
rect 1342 563 1348 564
rect 1510 568 1516 569
rect 1510 564 1511 568
rect 1515 564 1516 568
rect 1510 563 1516 564
rect 1670 568 1676 569
rect 1670 564 1671 568
rect 1675 564 1676 568
rect 1670 563 1676 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 3838 569 3844 570
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 1814 563 1820 564
rect 3886 563 3892 564
rect 4070 568 4076 569
rect 4070 564 4071 568
rect 4075 564 4076 568
rect 4070 563 4076 564
rect 4310 568 4316 569
rect 4310 564 4311 568
rect 4315 564 4316 568
rect 4310 563 4316 564
rect 4574 568 4580 569
rect 4574 564 4575 568
rect 4579 564 4580 568
rect 4574 563 4580 564
rect 4854 568 4860 569
rect 4854 564 4855 568
rect 4859 564 4860 568
rect 4854 563 4860 564
rect 5150 568 5156 569
rect 5150 564 5151 568
rect 5155 564 5156 568
rect 5150 563 5156 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 346 553 352 554
rect 346 549 347 553
rect 351 549 352 553
rect 346 548 352 549
rect 570 553 576 554
rect 570 549 571 553
rect 575 549 576 553
rect 570 548 576 549
rect 778 553 784 554
rect 778 549 779 553
rect 783 549 784 553
rect 778 548 784 549
rect 970 553 976 554
rect 970 549 971 553
rect 975 549 976 553
rect 970 548 976 549
rect 1146 553 1152 554
rect 1146 549 1147 553
rect 1151 549 1152 553
rect 1146 548 1152 549
rect 1314 553 1320 554
rect 1314 549 1315 553
rect 1319 549 1320 553
rect 1314 548 1320 549
rect 1482 553 1488 554
rect 1482 549 1483 553
rect 1487 549 1488 553
rect 1482 548 1488 549
rect 1642 553 1648 554
rect 1642 549 1643 553
rect 1647 549 1648 553
rect 1642 548 1648 549
rect 1786 553 1792 554
rect 3858 553 3864 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 3838 552 3844 553
rect 110 547 116 548
rect 1934 547 1940 548
rect 1974 549 1980 550
rect 3798 549 3804 550
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3134 548 3140 549
rect 3134 544 3135 548
rect 3139 544 3140 548
rect 3134 543 3140 544
rect 3270 548 3276 549
rect 3270 544 3271 548
rect 3275 544 3276 548
rect 3270 543 3276 544
rect 3406 548 3412 549
rect 3406 544 3407 548
rect 3411 544 3412 548
rect 3406 543 3412 544
rect 3542 548 3548 549
rect 3542 544 3543 548
rect 3547 544 3548 548
rect 3542 543 3548 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 4042 553 4048 554
rect 4042 549 4043 553
rect 4047 549 4048 553
rect 4042 548 4048 549
rect 4282 553 4288 554
rect 4282 549 4283 553
rect 4287 549 4288 553
rect 4282 548 4288 549
rect 4546 553 4552 554
rect 4546 549 4547 553
rect 4551 549 4552 553
rect 4546 548 4552 549
rect 4826 553 4832 554
rect 4826 549 4827 553
rect 4831 549 4832 553
rect 4826 548 4832 549
rect 5122 553 5128 554
rect 5122 549 5123 553
rect 5127 549 5128 553
rect 5122 548 5128 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 5662 547 5668 548
rect 3798 544 3804 545
rect 3678 543 3684 544
rect 3106 533 3112 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3106 529 3107 533
rect 3111 529 3112 533
rect 3106 528 3112 529
rect 3242 533 3248 534
rect 3242 529 3243 533
rect 3247 529 3248 533
rect 3242 528 3248 529
rect 3378 533 3384 534
rect 3378 529 3379 533
rect 3383 529 3384 533
rect 3378 528 3384 529
rect 3514 533 3520 534
rect 3514 529 3515 533
rect 3519 529 3520 533
rect 3514 528 3520 529
rect 3650 533 3656 534
rect 3650 529 3651 533
rect 3655 529 3656 533
rect 3650 528 3656 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 3798 527 3804 528
rect 110 420 116 421
rect 1934 420 1940 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 154 419 160 420
rect 154 415 155 419
rect 159 415 160 419
rect 154 414 160 415
rect 482 419 488 420
rect 482 415 483 419
rect 487 415 488 419
rect 482 414 488 415
rect 810 419 816 420
rect 810 415 811 419
rect 815 415 816 419
rect 810 414 816 415
rect 1138 419 1144 420
rect 1138 415 1139 419
rect 1143 415 1144 419
rect 1138 414 1144 415
rect 1474 419 1480 420
rect 1474 415 1475 419
rect 1479 415 1480 419
rect 1474 414 1480 415
rect 1786 419 1792 420
rect 1786 415 1787 419
rect 1791 415 1792 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 1786 414 1792 415
rect 3838 408 3844 409
rect 5662 408 5668 409
rect 182 404 188 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 182 400 183 404
rect 187 400 188 404
rect 182 399 188 400
rect 510 404 516 405
rect 510 400 511 404
rect 515 400 516 404
rect 510 399 516 400
rect 838 404 844 405
rect 838 400 839 404
rect 843 400 844 404
rect 838 399 844 400
rect 1166 404 1172 405
rect 1166 400 1167 404
rect 1171 400 1172 404
rect 1166 399 1172 400
rect 1502 404 1508 405
rect 1502 400 1503 404
rect 1507 400 1508 404
rect 1502 399 1508 400
rect 1814 404 1820 405
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 1814 400 1815 404
rect 1819 400 1820 404
rect 1814 399 1820 400
rect 1934 403 1940 404
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 4450 402 4456 403
rect 4642 407 4648 408
rect 4642 403 4643 407
rect 4647 403 4648 407
rect 4642 402 4648 403
rect 4842 407 4848 408
rect 4842 403 4843 407
rect 4847 403 4848 407
rect 4842 402 4848 403
rect 5050 407 5056 408
rect 5050 403 5051 407
rect 5055 403 5056 407
rect 5050 402 5056 403
rect 5266 407 5272 408
rect 5266 403 5267 407
rect 5271 403 5272 407
rect 5266 402 5272 403
rect 5482 407 5488 408
rect 5482 403 5483 407
rect 5487 403 5488 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5482 402 5488 403
rect 110 398 116 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 3798 400 3804 401
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2858 399 2864 400
rect 2858 395 2859 399
rect 2863 395 2864 399
rect 2858 394 2864 395
rect 3066 399 3072 400
rect 3066 395 3067 399
rect 3071 395 3072 399
rect 3066 394 3072 395
rect 3266 399 3272 400
rect 3266 395 3267 399
rect 3271 395 3272 399
rect 3266 394 3272 395
rect 3466 399 3472 400
rect 3466 395 3467 399
rect 3471 395 3472 399
rect 3466 394 3472 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4670 392 4676 393
rect 4670 388 4671 392
rect 4675 388 4676 392
rect 4670 387 4676 388
rect 4870 392 4876 393
rect 4870 388 4871 392
rect 4875 388 4876 392
rect 4870 387 4876 388
rect 5078 392 5084 393
rect 5078 388 5079 392
rect 5083 388 5084 392
rect 5078 387 5084 388
rect 5294 392 5300 393
rect 5294 388 5295 392
rect 5299 388 5300 392
rect 5294 387 5300 388
rect 5510 392 5516 393
rect 5510 388 5511 392
rect 5515 388 5516 392
rect 5510 387 5516 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 5662 386 5668 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 2886 384 2892 385
rect 2886 380 2887 384
rect 2891 380 2892 384
rect 2886 379 2892 380
rect 3094 384 3100 385
rect 3094 380 3095 384
rect 3099 380 3100 384
rect 3094 379 3100 380
rect 3294 384 3300 385
rect 3294 380 3295 384
rect 3299 380 3300 384
rect 3294 379 3300 380
rect 3494 384 3500 385
rect 3494 380 3495 384
rect 3499 380 3500 384
rect 3494 379 3500 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 3798 378 3804 379
rect 110 333 116 334
rect 1934 333 1940 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 278 332 284 333
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 486 332 492 333
rect 486 328 487 332
rect 491 328 492 332
rect 486 327 492 328
rect 702 332 708 333
rect 702 328 703 332
rect 707 328 708 332
rect 702 327 708 328
rect 918 332 924 333
rect 918 328 919 332
rect 923 328 924 332
rect 918 327 924 328
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 3838 329 3844 330
rect 5662 329 5668 330
rect 1134 327 1140 328
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4614 328 4620 329
rect 4614 324 4615 328
rect 4619 324 4620 328
rect 4614 323 4620 324
rect 4774 328 4780 329
rect 4774 324 4775 328
rect 4779 324 4780 328
rect 4774 323 4780 324
rect 4950 328 4956 329
rect 4950 324 4951 328
rect 4955 324 4956 328
rect 4950 323 4956 324
rect 5134 328 5140 329
rect 5134 324 5135 328
rect 5139 324 5140 328
rect 5134 323 5140 324
rect 5326 328 5332 329
rect 5326 324 5327 328
rect 5331 324 5332 328
rect 5326 323 5332 324
rect 5526 328 5532 329
rect 5526 324 5527 328
rect 5531 324 5532 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5526 323 5532 324
rect 250 317 256 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 250 313 251 317
rect 255 313 256 317
rect 250 312 256 313
rect 458 317 464 318
rect 458 313 459 317
rect 463 313 464 317
rect 458 312 464 313
rect 674 317 680 318
rect 674 313 675 317
rect 679 313 680 317
rect 674 312 680 313
rect 890 317 896 318
rect 890 313 891 317
rect 895 313 896 317
rect 890 312 896 313
rect 1106 317 1112 318
rect 1106 313 1107 317
rect 1111 313 1112 317
rect 1106 312 1112 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 4586 313 4592 314
rect 110 311 116 312
rect 1934 311 1940 312
rect 3838 312 3844 313
rect 1974 309 1980 310
rect 3798 309 3804 310
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4586 309 4587 313
rect 4591 309 4592 313
rect 4586 308 4592 309
rect 4746 313 4752 314
rect 4746 309 4747 313
rect 4751 309 4752 313
rect 4746 308 4752 309
rect 4922 313 4928 314
rect 4922 309 4923 313
rect 4927 309 4928 313
rect 4922 308 4928 309
rect 5106 313 5112 314
rect 5106 309 5107 313
rect 5111 309 5112 313
rect 5106 308 5112 309
rect 5298 313 5304 314
rect 5298 309 5299 313
rect 5303 309 5304 313
rect 5298 308 5304 309
rect 5498 313 5504 314
rect 5498 309 5499 313
rect 5503 309 5504 313
rect 5498 308 5504 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 5662 307 5668 308
rect 3798 304 3804 305
rect 3654 303 3660 304
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 1974 287 1980 288
rect 3798 287 3804 288
rect 110 144 116 145
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 3838 140 3844 141
rect 5662 140 5668 141
rect 1082 138 1088 139
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 110 122 116 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 3798 124 3804 125
rect 4318 124 4324 125
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3626 118 3632 119
rect 3838 118 3844 119
rect 5662 118 5668 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 3798 102 3804 103
<< m3c >>
rect 111 5725 115 5729
rect 159 5724 163 5728
rect 295 5724 299 5728
rect 1935 5725 1939 5729
rect 111 5708 115 5712
rect 131 5709 135 5713
rect 267 5709 271 5713
rect 1935 5708 1939 5712
rect 1975 5625 1979 5629
rect 2023 5624 2027 5628
rect 2183 5624 2187 5628
rect 2367 5624 2371 5628
rect 2551 5624 2555 5628
rect 2727 5624 2731 5628
rect 2895 5624 2899 5628
rect 3063 5624 3067 5628
rect 3223 5624 3227 5628
rect 3383 5624 3387 5628
rect 3543 5624 3547 5628
rect 3679 5624 3683 5628
rect 3799 5625 3803 5629
rect 3839 5621 3843 5625
rect 4335 5620 4339 5624
rect 4471 5620 4475 5624
rect 4607 5620 4611 5624
rect 4743 5620 4747 5624
rect 4879 5620 4883 5624
rect 5015 5620 5019 5624
rect 5663 5621 5667 5625
rect 1975 5608 1979 5612
rect 1995 5609 1999 5613
rect 2155 5609 2159 5613
rect 2339 5609 2343 5613
rect 2523 5609 2527 5613
rect 2699 5609 2703 5613
rect 2867 5609 2871 5613
rect 3035 5609 3039 5613
rect 3195 5609 3199 5613
rect 3355 5609 3359 5613
rect 3515 5609 3519 5613
rect 3651 5609 3655 5613
rect 3799 5608 3803 5612
rect 3839 5604 3843 5608
rect 4307 5605 4311 5609
rect 4443 5605 4447 5609
rect 4579 5605 4583 5609
rect 4715 5605 4719 5609
rect 4851 5605 4855 5609
rect 4987 5605 4991 5609
rect 5663 5604 5667 5608
rect 111 5576 115 5580
rect 131 5575 135 5579
rect 275 5575 279 5579
rect 475 5575 479 5579
rect 699 5575 703 5579
rect 955 5575 959 5579
rect 1227 5575 1231 5579
rect 1515 5575 1519 5579
rect 1787 5575 1791 5579
rect 1935 5576 1939 5580
rect 111 5559 115 5563
rect 159 5560 163 5564
rect 303 5560 307 5564
rect 503 5560 507 5564
rect 727 5560 731 5564
rect 983 5560 987 5564
rect 1255 5560 1259 5564
rect 1543 5560 1547 5564
rect 1815 5560 1819 5564
rect 1935 5559 1939 5563
rect 111 5501 115 5505
rect 279 5500 283 5504
rect 519 5500 523 5504
rect 767 5500 771 5504
rect 1015 5500 1019 5504
rect 1263 5500 1267 5504
rect 1511 5500 1515 5504
rect 1767 5500 1771 5504
rect 1935 5501 1939 5505
rect 111 5484 115 5488
rect 251 5485 255 5489
rect 491 5485 495 5489
rect 739 5485 743 5489
rect 987 5485 991 5489
rect 1235 5485 1239 5489
rect 1483 5485 1487 5489
rect 1739 5485 1743 5489
rect 1935 5484 1939 5488
rect 1975 5476 1979 5480
rect 2139 5475 2143 5479
rect 2355 5475 2359 5479
rect 2563 5475 2567 5479
rect 2755 5475 2759 5479
rect 2939 5475 2943 5479
rect 3115 5475 3119 5479
rect 3291 5475 3295 5479
rect 3467 5475 3471 5479
rect 3643 5475 3647 5479
rect 3799 5476 3803 5480
rect 3839 5472 3843 5476
rect 4251 5471 4255 5475
rect 4403 5471 4407 5475
rect 4555 5471 4559 5475
rect 4707 5471 4711 5475
rect 4859 5471 4863 5475
rect 5019 5471 5023 5475
rect 5663 5472 5667 5476
rect 1975 5459 1979 5463
rect 2167 5460 2171 5464
rect 2383 5460 2387 5464
rect 2591 5460 2595 5464
rect 2783 5460 2787 5464
rect 2967 5460 2971 5464
rect 3143 5460 3147 5464
rect 3319 5460 3323 5464
rect 3495 5460 3499 5464
rect 3671 5460 3675 5464
rect 3799 5459 3803 5463
rect 3839 5455 3843 5459
rect 4279 5456 4283 5460
rect 4431 5456 4435 5460
rect 4583 5456 4587 5460
rect 4735 5456 4739 5460
rect 4887 5456 4891 5460
rect 5047 5456 5051 5460
rect 5663 5455 5667 5459
rect 1975 5393 1979 5397
rect 2311 5392 2315 5396
rect 2511 5392 2515 5396
rect 2703 5392 2707 5396
rect 2887 5392 2891 5396
rect 3071 5392 3075 5396
rect 3247 5392 3251 5396
rect 3423 5392 3427 5396
rect 3607 5392 3611 5396
rect 3799 5393 3803 5397
rect 1975 5376 1979 5380
rect 2283 5377 2287 5381
rect 2483 5377 2487 5381
rect 2675 5377 2679 5381
rect 2859 5377 2863 5381
rect 3043 5377 3047 5381
rect 3219 5377 3223 5381
rect 3395 5377 3399 5381
rect 3579 5377 3583 5381
rect 3799 5376 3803 5380
rect 3839 5377 3843 5381
rect 4279 5376 4283 5380
rect 4487 5376 4491 5380
rect 4695 5376 4699 5380
rect 4911 5376 4915 5380
rect 5127 5376 5131 5380
rect 5663 5377 5667 5381
rect 3839 5360 3843 5364
rect 4251 5361 4255 5365
rect 4459 5361 4463 5365
rect 4667 5361 4671 5365
rect 4883 5361 4887 5365
rect 5099 5361 5103 5365
rect 5663 5360 5667 5364
rect 111 5352 115 5356
rect 411 5351 415 5355
rect 611 5351 615 5355
rect 819 5351 823 5355
rect 1035 5351 1039 5355
rect 1259 5351 1263 5355
rect 1491 5351 1495 5355
rect 1935 5352 1939 5356
rect 111 5335 115 5339
rect 439 5336 443 5340
rect 639 5336 643 5340
rect 847 5336 851 5340
rect 1063 5336 1067 5340
rect 1287 5336 1291 5340
rect 1519 5336 1523 5340
rect 1935 5335 1939 5339
rect 111 5277 115 5281
rect 591 5276 595 5280
rect 727 5276 731 5280
rect 863 5276 867 5280
rect 999 5276 1003 5280
rect 1135 5276 1139 5280
rect 1271 5276 1275 5280
rect 1407 5276 1411 5280
rect 1543 5276 1547 5280
rect 1935 5277 1939 5281
rect 111 5260 115 5264
rect 563 5261 567 5265
rect 699 5261 703 5265
rect 835 5261 839 5265
rect 971 5261 975 5265
rect 1107 5261 1111 5265
rect 1243 5261 1247 5265
rect 1379 5261 1383 5265
rect 1515 5261 1519 5265
rect 1935 5260 1939 5264
rect 1975 5244 1979 5248
rect 2195 5243 2199 5247
rect 2339 5243 2343 5247
rect 2491 5243 2495 5247
rect 2651 5243 2655 5247
rect 2819 5243 2823 5247
rect 3003 5243 3007 5247
rect 3187 5243 3191 5247
rect 3379 5243 3383 5247
rect 3579 5243 3583 5247
rect 3799 5244 3803 5248
rect 1975 5227 1979 5231
rect 2223 5228 2227 5232
rect 2367 5228 2371 5232
rect 2519 5228 2523 5232
rect 2679 5228 2683 5232
rect 2847 5228 2851 5232
rect 3031 5228 3035 5232
rect 3215 5228 3219 5232
rect 3407 5228 3411 5232
rect 3607 5228 3611 5232
rect 3799 5227 3803 5231
rect 3839 5212 3843 5216
rect 4251 5211 4255 5215
rect 4483 5211 4487 5215
rect 4715 5211 4719 5215
rect 4947 5211 4951 5215
rect 5187 5211 5191 5215
rect 5663 5212 5667 5216
rect 3839 5195 3843 5199
rect 4279 5196 4283 5200
rect 4511 5196 4515 5200
rect 4743 5196 4747 5200
rect 4975 5196 4979 5200
rect 5215 5196 5219 5200
rect 5663 5195 5667 5199
rect 1975 5169 1979 5173
rect 2023 5168 2027 5172
rect 2159 5168 2163 5172
rect 2327 5168 2331 5172
rect 2511 5168 2515 5172
rect 2695 5168 2699 5172
rect 2887 5168 2891 5172
rect 3087 5168 3091 5172
rect 3287 5168 3291 5172
rect 3495 5168 3499 5172
rect 3679 5168 3683 5172
rect 3799 5169 3803 5173
rect 1975 5152 1979 5156
rect 1995 5153 1999 5157
rect 2131 5153 2135 5157
rect 2299 5153 2303 5157
rect 2483 5153 2487 5157
rect 2667 5153 2671 5157
rect 2859 5153 2863 5157
rect 3059 5153 3063 5157
rect 3259 5153 3263 5157
rect 3467 5153 3471 5157
rect 3651 5153 3655 5157
rect 3799 5152 3803 5156
rect 3839 5109 3843 5113
rect 3887 5108 3891 5112
rect 4135 5108 4139 5112
rect 4407 5108 4411 5112
rect 4679 5108 4683 5112
rect 4959 5108 4963 5112
rect 5239 5108 5243 5112
rect 5663 5109 5667 5113
rect 3839 5092 3843 5096
rect 3859 5093 3863 5097
rect 4107 5093 4111 5097
rect 4379 5093 4383 5097
rect 4651 5093 4655 5097
rect 4931 5093 4935 5097
rect 5211 5093 5215 5097
rect 5663 5092 5667 5096
rect 111 5024 115 5028
rect 347 5023 351 5027
rect 483 5023 487 5027
rect 619 5023 623 5027
rect 755 5023 759 5027
rect 891 5023 895 5027
rect 1035 5023 1039 5027
rect 1187 5023 1191 5027
rect 1339 5023 1343 5027
rect 1491 5023 1495 5027
rect 1651 5023 1655 5027
rect 1787 5023 1791 5027
rect 1935 5024 1939 5028
rect 1975 5020 1979 5024
rect 1995 5019 1999 5023
rect 2531 5019 2535 5023
rect 3099 5019 3103 5023
rect 3651 5019 3655 5023
rect 3799 5020 3803 5024
rect 111 5007 115 5011
rect 375 5008 379 5012
rect 511 5008 515 5012
rect 647 5008 651 5012
rect 783 5008 787 5012
rect 919 5008 923 5012
rect 1063 5008 1067 5012
rect 1215 5008 1219 5012
rect 1367 5008 1371 5012
rect 1519 5008 1523 5012
rect 1679 5008 1683 5012
rect 1815 5008 1819 5012
rect 1935 5007 1939 5011
rect 1975 5003 1979 5007
rect 2023 5004 2027 5008
rect 2559 5004 2563 5008
rect 3127 5004 3131 5008
rect 3679 5004 3683 5008
rect 3799 5003 3803 5007
rect 111 4949 115 4953
rect 159 4948 163 4952
rect 343 4948 347 4952
rect 551 4948 555 4952
rect 751 4948 755 4952
rect 943 4948 947 4952
rect 1127 4948 1131 4952
rect 1311 4948 1315 4952
rect 1487 4948 1491 4952
rect 1663 4948 1667 4952
rect 1815 4948 1819 4952
rect 1935 4949 1939 4953
rect 3839 4948 3843 4952
rect 3859 4947 3863 4951
rect 4019 4947 4023 4951
rect 4211 4947 4215 4951
rect 4411 4947 4415 4951
rect 4627 4947 4631 4951
rect 4843 4947 4847 4951
rect 5067 4947 5071 4951
rect 5299 4947 5303 4951
rect 5663 4948 5667 4952
rect 111 4932 115 4936
rect 131 4933 135 4937
rect 315 4933 319 4937
rect 523 4933 527 4937
rect 723 4933 727 4937
rect 915 4933 919 4937
rect 1099 4933 1103 4937
rect 1283 4933 1287 4937
rect 1459 4933 1463 4937
rect 1635 4933 1639 4937
rect 1787 4933 1791 4937
rect 1935 4932 1939 4936
rect 3839 4931 3843 4935
rect 3887 4932 3891 4936
rect 4047 4932 4051 4936
rect 4239 4932 4243 4936
rect 4439 4932 4443 4936
rect 4655 4932 4659 4936
rect 4871 4932 4875 4936
rect 5095 4932 5099 4936
rect 5327 4932 5331 4936
rect 5663 4931 5667 4935
rect 1975 4913 1979 4917
rect 2871 4912 2875 4916
rect 3007 4912 3011 4916
rect 3799 4913 3803 4917
rect 1975 4896 1979 4900
rect 2843 4897 2847 4901
rect 2979 4897 2983 4901
rect 3799 4896 3803 4900
rect 3839 4853 3843 4857
rect 3887 4852 3891 4856
rect 4071 4852 4075 4856
rect 4287 4852 4291 4856
rect 4511 4852 4515 4856
rect 4735 4852 4739 4856
rect 4959 4852 4963 4856
rect 5183 4852 5187 4856
rect 5407 4852 5411 4856
rect 5663 4853 5667 4857
rect 3839 4836 3843 4840
rect 3859 4837 3863 4841
rect 4043 4837 4047 4841
rect 4259 4837 4263 4841
rect 4483 4837 4487 4841
rect 4707 4837 4711 4841
rect 4931 4837 4935 4841
rect 5155 4837 5159 4841
rect 5379 4837 5383 4841
rect 5663 4836 5667 4840
rect 111 4792 115 4796
rect 131 4791 135 4795
rect 267 4791 271 4795
rect 403 4791 407 4795
rect 539 4791 543 4795
rect 675 4791 679 4795
rect 1935 4792 1939 4796
rect 111 4775 115 4779
rect 159 4776 163 4780
rect 295 4776 299 4780
rect 431 4776 435 4780
rect 567 4776 571 4780
rect 703 4776 707 4780
rect 1935 4775 1939 4779
rect 1975 4740 1979 4744
rect 1995 4739 1999 4743
rect 2155 4739 2159 4743
rect 2347 4739 2351 4743
rect 2539 4739 2543 4743
rect 2731 4739 2735 4743
rect 2931 4739 2935 4743
rect 3131 4739 3135 4743
rect 3799 4740 3803 4744
rect 1975 4723 1979 4727
rect 2023 4724 2027 4728
rect 2183 4724 2187 4728
rect 2375 4724 2379 4728
rect 2567 4724 2571 4728
rect 2759 4724 2763 4728
rect 2959 4724 2963 4728
rect 3159 4724 3163 4728
rect 3799 4723 3803 4727
rect 111 4709 115 4713
rect 159 4708 163 4712
rect 343 4708 347 4712
rect 567 4708 571 4712
rect 807 4708 811 4712
rect 1055 4708 1059 4712
rect 1311 4708 1315 4712
rect 1575 4708 1579 4712
rect 1815 4708 1819 4712
rect 1935 4709 1939 4713
rect 3839 4700 3843 4704
rect 3915 4699 3919 4703
rect 4187 4699 4191 4703
rect 4467 4699 4471 4703
rect 4763 4699 4767 4703
rect 5067 4699 5071 4703
rect 5371 4699 5375 4703
rect 5663 4700 5667 4704
rect 111 4692 115 4696
rect 131 4693 135 4697
rect 315 4693 319 4697
rect 539 4693 543 4697
rect 779 4693 783 4697
rect 1027 4693 1031 4697
rect 1283 4693 1287 4697
rect 1547 4693 1551 4697
rect 1787 4693 1791 4697
rect 1935 4692 1939 4696
rect 3839 4683 3843 4687
rect 3943 4684 3947 4688
rect 4215 4684 4219 4688
rect 4495 4684 4499 4688
rect 4791 4684 4795 4688
rect 5095 4684 5099 4688
rect 5399 4684 5403 4688
rect 5663 4683 5667 4687
rect 1975 4661 1979 4665
rect 2023 4660 2027 4664
rect 2239 4660 2243 4664
rect 2471 4660 2475 4664
rect 2695 4660 2699 4664
rect 2919 4660 2923 4664
rect 3143 4660 3147 4664
rect 3367 4660 3371 4664
rect 3799 4661 3803 4665
rect 1975 4644 1979 4648
rect 1995 4645 1999 4649
rect 2211 4645 2215 4649
rect 2443 4645 2447 4649
rect 2667 4645 2671 4649
rect 2891 4645 2895 4649
rect 3115 4645 3119 4649
rect 3339 4645 3343 4649
rect 3799 4644 3803 4648
rect 3839 4625 3843 4629
rect 4063 4624 4067 4628
rect 4327 4624 4331 4628
rect 4599 4624 4603 4628
rect 4871 4624 4875 4628
rect 5151 4624 5155 4628
rect 5439 4624 5443 4628
rect 5663 4625 5667 4629
rect 3839 4608 3843 4612
rect 4035 4609 4039 4613
rect 4299 4609 4303 4613
rect 4571 4609 4575 4613
rect 4843 4609 4847 4613
rect 5123 4609 5127 4613
rect 5411 4609 5415 4613
rect 5663 4608 5667 4612
rect 111 4544 115 4548
rect 171 4543 175 4547
rect 395 4543 399 4547
rect 643 4543 647 4547
rect 907 4543 911 4547
rect 1195 4543 1199 4547
rect 1491 4543 1495 4547
rect 1787 4543 1791 4547
rect 1935 4544 1939 4548
rect 111 4527 115 4531
rect 199 4528 203 4532
rect 423 4528 427 4532
rect 671 4528 675 4532
rect 935 4528 939 4532
rect 1223 4528 1227 4532
rect 1519 4528 1523 4532
rect 1815 4528 1819 4532
rect 1935 4527 1939 4531
rect 1975 4508 1979 4512
rect 2099 4507 2103 4511
rect 2347 4507 2351 4511
rect 2579 4507 2583 4511
rect 2795 4507 2799 4511
rect 3003 4507 3007 4511
rect 3203 4507 3207 4511
rect 3403 4507 3407 4511
rect 3611 4507 3615 4511
rect 3799 4508 3803 4512
rect 1975 4491 1979 4495
rect 2127 4492 2131 4496
rect 2375 4492 2379 4496
rect 2607 4492 2611 4496
rect 2823 4492 2827 4496
rect 3031 4492 3035 4496
rect 3231 4492 3235 4496
rect 3431 4492 3435 4496
rect 3639 4492 3643 4496
rect 3799 4491 3803 4495
rect 3839 4476 3843 4480
rect 4179 4475 4183 4479
rect 4411 4475 4415 4479
rect 4659 4475 4663 4479
rect 4915 4475 4919 4479
rect 5179 4475 5183 4479
rect 5443 4475 5447 4479
rect 5663 4476 5667 4480
rect 111 4465 115 4469
rect 447 4464 451 4468
rect 655 4464 659 4468
rect 887 4464 891 4468
rect 1143 4464 1147 4468
rect 1407 4464 1411 4468
rect 1679 4464 1683 4468
rect 1935 4465 1939 4469
rect 3839 4459 3843 4463
rect 4207 4460 4211 4464
rect 4439 4460 4443 4464
rect 4687 4460 4691 4464
rect 4943 4460 4947 4464
rect 5207 4460 5211 4464
rect 5471 4460 5475 4464
rect 5663 4459 5667 4463
rect 111 4448 115 4452
rect 419 4449 423 4453
rect 627 4449 631 4453
rect 859 4449 863 4453
rect 1115 4449 1119 4453
rect 1379 4449 1383 4453
rect 1651 4449 1655 4453
rect 1935 4448 1939 4452
rect 1975 4425 1979 4429
rect 2231 4424 2235 4428
rect 2447 4424 2451 4428
rect 2663 4424 2667 4428
rect 2871 4424 2875 4428
rect 3079 4424 3083 4428
rect 3287 4424 3291 4428
rect 3495 4424 3499 4428
rect 3679 4424 3683 4428
rect 3799 4425 3803 4429
rect 1975 4408 1979 4412
rect 2203 4409 2207 4413
rect 2419 4409 2423 4413
rect 2635 4409 2639 4413
rect 2843 4409 2847 4413
rect 3051 4409 3055 4413
rect 3259 4409 3263 4413
rect 3467 4409 3471 4413
rect 3651 4409 3655 4413
rect 3799 4408 3803 4412
rect 3839 4393 3843 4397
rect 4359 4392 4363 4396
rect 4519 4392 4523 4396
rect 4687 4392 4691 4396
rect 4879 4392 4883 4396
rect 5079 4392 5083 4396
rect 5287 4392 5291 4396
rect 5503 4392 5507 4396
rect 5663 4393 5667 4397
rect 3839 4376 3843 4380
rect 4331 4377 4335 4381
rect 4491 4377 4495 4381
rect 4659 4377 4663 4381
rect 4851 4377 4855 4381
rect 5051 4377 5055 4381
rect 5259 4377 5263 4381
rect 5475 4377 5479 4381
rect 5663 4376 5667 4380
rect 111 4312 115 4316
rect 667 4311 671 4315
rect 811 4311 815 4315
rect 963 4311 967 4315
rect 1123 4311 1127 4315
rect 1291 4311 1295 4315
rect 1467 4311 1471 4315
rect 1651 4311 1655 4315
rect 1935 4312 1939 4316
rect 111 4295 115 4299
rect 695 4296 699 4300
rect 839 4296 843 4300
rect 991 4296 995 4300
rect 1151 4296 1155 4300
rect 1319 4296 1323 4300
rect 1495 4296 1499 4300
rect 1679 4296 1683 4300
rect 1935 4295 1939 4299
rect 1975 4268 1979 4272
rect 2307 4267 2311 4271
rect 2459 4267 2463 4271
rect 2627 4267 2631 4271
rect 2811 4267 2815 4271
rect 3011 4267 3015 4271
rect 3227 4267 3231 4271
rect 3451 4267 3455 4271
rect 3651 4267 3655 4271
rect 3799 4268 3803 4272
rect 1975 4251 1979 4255
rect 2335 4252 2339 4256
rect 2487 4252 2491 4256
rect 2655 4252 2659 4256
rect 2839 4252 2843 4256
rect 3039 4252 3043 4256
rect 3255 4252 3259 4256
rect 3479 4252 3483 4256
rect 3679 4252 3683 4256
rect 3799 4251 3803 4255
rect 3839 4244 3843 4248
rect 3859 4243 3863 4247
rect 4043 4243 4047 4247
rect 4251 4243 4255 4247
rect 4475 4243 4479 4247
rect 4715 4243 4719 4247
rect 4971 4243 4975 4247
rect 5235 4243 5239 4247
rect 5499 4243 5503 4247
rect 5663 4244 5667 4248
rect 3839 4227 3843 4231
rect 3887 4228 3891 4232
rect 4071 4228 4075 4232
rect 4279 4228 4283 4232
rect 4503 4228 4507 4232
rect 4743 4228 4747 4232
rect 4999 4228 5003 4232
rect 5263 4228 5267 4232
rect 5527 4228 5531 4232
rect 5663 4227 5667 4231
rect 111 4221 115 4225
rect 815 4220 819 4224
rect 951 4220 955 4224
rect 1087 4220 1091 4224
rect 1223 4220 1227 4224
rect 1359 4220 1363 4224
rect 1495 4220 1499 4224
rect 1631 4220 1635 4224
rect 1767 4220 1771 4224
rect 1935 4221 1939 4225
rect 111 4204 115 4208
rect 787 4205 791 4209
rect 923 4205 927 4209
rect 1059 4205 1063 4209
rect 1195 4205 1199 4209
rect 1331 4205 1335 4209
rect 1467 4205 1471 4209
rect 1603 4205 1607 4209
rect 1739 4205 1743 4209
rect 1935 4204 1939 4208
rect 1975 4185 1979 4189
rect 2567 4184 2571 4188
rect 2703 4184 2707 4188
rect 2839 4184 2843 4188
rect 2975 4184 2979 4188
rect 3799 4185 3803 4189
rect 1975 4168 1979 4172
rect 2539 4169 2543 4173
rect 2675 4169 2679 4173
rect 2811 4169 2815 4173
rect 2947 4169 2951 4173
rect 3799 4168 3803 4172
rect 3839 4133 3843 4137
rect 3887 4132 3891 4136
rect 4415 4132 4419 4136
rect 4975 4132 4979 4136
rect 5543 4132 5547 4136
rect 5663 4133 5667 4137
rect 3839 4116 3843 4120
rect 3859 4117 3863 4121
rect 4387 4117 4391 4121
rect 4947 4117 4951 4121
rect 5515 4117 5519 4121
rect 5663 4116 5667 4120
rect 111 4068 115 4072
rect 731 4067 735 4071
rect 867 4067 871 4071
rect 1003 4067 1007 4071
rect 1139 4067 1143 4071
rect 1275 4067 1279 4071
rect 1411 4067 1415 4071
rect 1547 4067 1551 4071
rect 1935 4068 1939 4072
rect 111 4051 115 4055
rect 759 4052 763 4056
rect 895 4052 899 4056
rect 1031 4052 1035 4056
rect 1167 4052 1171 4056
rect 1303 4052 1307 4056
rect 1439 4052 1443 4056
rect 1575 4052 1579 4056
rect 1935 4051 1939 4055
rect 1975 4016 1979 4020
rect 2291 4015 2295 4019
rect 2427 4015 2431 4019
rect 2563 4015 2567 4019
rect 2699 4015 2703 4019
rect 2835 4015 2839 4019
rect 3799 4016 3803 4020
rect 1975 3999 1979 4003
rect 2319 4000 2323 4004
rect 2455 4000 2459 4004
rect 2591 4000 2595 4004
rect 2727 4000 2731 4004
rect 2863 4000 2867 4004
rect 3799 3999 3803 4003
rect 3839 3984 3843 3988
rect 3859 3983 3863 3987
rect 4003 3983 4007 3987
rect 4171 3983 4175 3987
rect 4339 3983 4343 3987
rect 4499 3983 4503 3987
rect 4651 3983 4655 3987
rect 4803 3983 4807 3987
rect 4947 3983 4951 3987
rect 5091 3983 5095 3987
rect 5235 3983 5239 3987
rect 5379 3983 5383 3987
rect 5515 3983 5519 3987
rect 5663 3984 5667 3988
rect 111 3969 115 3973
rect 511 3968 515 3972
rect 663 3968 667 3972
rect 823 3968 827 3972
rect 983 3968 987 3972
rect 1151 3968 1155 3972
rect 1319 3968 1323 3972
rect 1935 3969 1939 3973
rect 3839 3967 3843 3971
rect 3887 3968 3891 3972
rect 4031 3968 4035 3972
rect 4199 3968 4203 3972
rect 4367 3968 4371 3972
rect 4527 3968 4531 3972
rect 4679 3968 4683 3972
rect 4831 3968 4835 3972
rect 4975 3968 4979 3972
rect 5119 3968 5123 3972
rect 5263 3968 5267 3972
rect 5407 3968 5411 3972
rect 5543 3968 5547 3972
rect 5663 3967 5667 3971
rect 111 3952 115 3956
rect 483 3953 487 3957
rect 635 3953 639 3957
rect 795 3953 799 3957
rect 955 3953 959 3957
rect 1123 3953 1127 3957
rect 1291 3953 1295 3957
rect 1935 3952 1939 3956
rect 1975 3937 1979 3941
rect 2119 3936 2123 3940
rect 2327 3936 2331 3940
rect 2535 3936 2539 3940
rect 2743 3936 2747 3940
rect 2943 3936 2947 3940
rect 3135 3936 3139 3940
rect 3319 3936 3323 3940
rect 3511 3936 3515 3940
rect 3679 3936 3683 3940
rect 3799 3937 3803 3941
rect 1975 3920 1979 3924
rect 2091 3921 2095 3925
rect 2299 3921 2303 3925
rect 2507 3921 2511 3925
rect 2715 3921 2719 3925
rect 2915 3921 2919 3925
rect 3107 3921 3111 3925
rect 3291 3921 3295 3925
rect 3483 3921 3487 3925
rect 3651 3921 3655 3925
rect 3799 3920 3803 3924
rect 3839 3885 3843 3889
rect 4383 3884 4387 3888
rect 4599 3884 4603 3888
rect 4823 3884 4827 3888
rect 5063 3884 5067 3888
rect 5311 3884 5315 3888
rect 5543 3884 5547 3888
rect 5663 3885 5667 3889
rect 3839 3868 3843 3872
rect 4355 3869 4359 3873
rect 4571 3869 4575 3873
rect 4795 3869 4799 3873
rect 5035 3869 5039 3873
rect 5283 3869 5287 3873
rect 5515 3869 5519 3873
rect 5663 3868 5667 3872
rect 111 3792 115 3796
rect 131 3791 135 3795
rect 307 3791 311 3795
rect 515 3791 519 3795
rect 723 3791 727 3795
rect 939 3791 943 3795
rect 1163 3791 1167 3795
rect 1935 3792 1939 3796
rect 111 3775 115 3779
rect 159 3776 163 3780
rect 335 3776 339 3780
rect 543 3776 547 3780
rect 751 3776 755 3780
rect 967 3776 971 3780
rect 1191 3776 1195 3780
rect 1935 3775 1939 3779
rect 1975 3776 1979 3780
rect 2139 3775 2143 3779
rect 2371 3775 2375 3779
rect 2587 3775 2591 3779
rect 2795 3775 2799 3779
rect 2995 3775 2999 3779
rect 3195 3775 3199 3779
rect 3403 3775 3407 3779
rect 3799 3776 3803 3780
rect 1975 3759 1979 3763
rect 2167 3760 2171 3764
rect 2399 3760 2403 3764
rect 2615 3760 2619 3764
rect 2823 3760 2827 3764
rect 3023 3760 3027 3764
rect 3223 3760 3227 3764
rect 3431 3760 3435 3764
rect 3799 3759 3803 3763
rect 111 3717 115 3721
rect 159 3716 163 3720
rect 335 3716 339 3720
rect 527 3716 531 3720
rect 711 3716 715 3720
rect 887 3716 891 3720
rect 1055 3716 1059 3720
rect 1215 3716 1219 3720
rect 1367 3716 1371 3720
rect 1519 3716 1523 3720
rect 1679 3716 1683 3720
rect 1815 3716 1819 3720
rect 1935 3717 1939 3721
rect 3839 3720 3843 3724
rect 3995 3719 3999 3723
rect 4203 3719 4207 3723
rect 4435 3719 4439 3723
rect 4691 3719 4695 3723
rect 4963 3719 4967 3723
rect 5251 3719 5255 3723
rect 5515 3719 5519 3723
rect 5663 3720 5667 3724
rect 111 3700 115 3704
rect 131 3701 135 3705
rect 307 3701 311 3705
rect 499 3701 503 3705
rect 683 3701 687 3705
rect 859 3701 863 3705
rect 1027 3701 1031 3705
rect 1187 3701 1191 3705
rect 1339 3701 1343 3705
rect 1491 3701 1495 3705
rect 1651 3701 1655 3705
rect 1787 3701 1791 3705
rect 1935 3700 1939 3704
rect 3839 3703 3843 3707
rect 4023 3704 4027 3708
rect 4231 3704 4235 3708
rect 4463 3704 4467 3708
rect 4719 3704 4723 3708
rect 4991 3704 4995 3708
rect 5279 3704 5283 3708
rect 5543 3704 5547 3708
rect 5663 3703 5667 3707
rect 1975 3697 1979 3701
rect 2279 3696 2283 3700
rect 2479 3696 2483 3700
rect 2679 3696 2683 3700
rect 2879 3696 2883 3700
rect 3079 3696 3083 3700
rect 3279 3696 3283 3700
rect 3799 3697 3803 3701
rect 1975 3680 1979 3684
rect 2251 3681 2255 3685
rect 2451 3681 2455 3685
rect 2651 3681 2655 3685
rect 2851 3681 2855 3685
rect 3051 3681 3055 3685
rect 3251 3681 3255 3685
rect 3799 3680 3803 3684
rect 3839 3617 3843 3621
rect 4215 3616 4219 3620
rect 4399 3616 4403 3620
rect 4607 3616 4611 3620
rect 4831 3616 4835 3620
rect 5071 3616 5075 3620
rect 5319 3616 5323 3620
rect 5543 3616 5547 3620
rect 5663 3617 5667 3621
rect 3839 3600 3843 3604
rect 4187 3601 4191 3605
rect 4371 3601 4375 3605
rect 4579 3601 4583 3605
rect 4803 3601 4807 3605
rect 5043 3601 5047 3605
rect 5291 3601 5295 3605
rect 5515 3601 5519 3605
rect 5663 3600 5667 3604
rect 111 3556 115 3560
rect 147 3555 151 3559
rect 355 3555 359 3559
rect 571 3555 575 3559
rect 803 3555 807 3559
rect 1043 3555 1047 3559
rect 1291 3555 1295 3559
rect 1547 3555 1551 3559
rect 1787 3555 1791 3559
rect 1935 3556 1939 3560
rect 111 3539 115 3543
rect 175 3540 179 3544
rect 383 3540 387 3544
rect 599 3540 603 3544
rect 831 3540 835 3544
rect 1071 3540 1075 3544
rect 1319 3540 1323 3544
rect 1575 3540 1579 3544
rect 1815 3540 1819 3544
rect 1935 3539 1939 3543
rect 1975 3536 1979 3540
rect 1995 3535 1999 3539
rect 2251 3535 2255 3539
rect 2515 3535 2519 3539
rect 2755 3535 2759 3539
rect 2979 3535 2983 3539
rect 3195 3535 3199 3539
rect 3411 3535 3415 3539
rect 3627 3535 3631 3539
rect 3799 3536 3803 3540
rect 1975 3519 1979 3523
rect 2023 3520 2027 3524
rect 2279 3520 2283 3524
rect 2543 3520 2547 3524
rect 2783 3520 2787 3524
rect 3007 3520 3011 3524
rect 3223 3520 3227 3524
rect 3439 3520 3443 3524
rect 3655 3520 3659 3524
rect 3799 3519 3803 3523
rect 111 3457 115 3461
rect 303 3456 307 3460
rect 447 3456 451 3460
rect 599 3456 603 3460
rect 759 3456 763 3460
rect 935 3456 939 3460
rect 1111 3456 1115 3460
rect 1295 3456 1299 3460
rect 1487 3456 1491 3460
rect 1935 3457 1939 3461
rect 1975 3453 1979 3457
rect 2023 3452 2027 3456
rect 2191 3452 2195 3456
rect 2399 3452 2403 3456
rect 2615 3452 2619 3456
rect 2831 3452 2835 3456
rect 3047 3452 3051 3456
rect 3263 3452 3267 3456
rect 3479 3452 3483 3456
rect 3679 3452 3683 3456
rect 3799 3453 3803 3457
rect 111 3440 115 3444
rect 275 3441 279 3445
rect 419 3441 423 3445
rect 571 3441 575 3445
rect 731 3441 735 3445
rect 907 3441 911 3445
rect 1083 3441 1087 3445
rect 1267 3441 1271 3445
rect 1459 3441 1463 3445
rect 1935 3440 1939 3444
rect 3839 3444 3843 3448
rect 4531 3443 4535 3447
rect 4683 3443 4687 3447
rect 4843 3443 4847 3447
rect 5003 3443 5007 3447
rect 5171 3443 5175 3447
rect 5347 3443 5351 3447
rect 5515 3443 5519 3447
rect 5663 3444 5667 3448
rect 1975 3436 1979 3440
rect 1995 3437 1999 3441
rect 2163 3437 2167 3441
rect 2371 3437 2375 3441
rect 2587 3437 2591 3441
rect 2803 3437 2807 3441
rect 3019 3437 3023 3441
rect 3235 3437 3239 3441
rect 3451 3437 3455 3441
rect 3651 3437 3655 3441
rect 3799 3436 3803 3440
rect 3839 3427 3843 3431
rect 4559 3428 4563 3432
rect 4711 3428 4715 3432
rect 4871 3428 4875 3432
rect 5031 3428 5035 3432
rect 5199 3428 5203 3432
rect 5375 3428 5379 3432
rect 5543 3428 5547 3432
rect 5663 3427 5667 3431
rect 3839 3365 3843 3369
rect 3887 3364 3891 3368
rect 4151 3364 4155 3368
rect 4423 3364 4427 3368
rect 4671 3364 4675 3368
rect 4895 3364 4899 3368
rect 5111 3364 5115 3368
rect 5327 3364 5331 3368
rect 5543 3364 5547 3368
rect 5663 3365 5667 3369
rect 3839 3348 3843 3352
rect 3859 3349 3863 3353
rect 4123 3349 4127 3353
rect 4395 3349 4399 3353
rect 4643 3349 4647 3353
rect 4867 3349 4871 3353
rect 5083 3349 5087 3353
rect 5299 3349 5303 3353
rect 5515 3349 5519 3353
rect 5663 3348 5667 3352
rect 111 3292 115 3296
rect 467 3291 471 3295
rect 667 3291 671 3295
rect 875 3291 879 3295
rect 1091 3291 1095 3295
rect 1315 3291 1319 3295
rect 1935 3292 1939 3296
rect 111 3275 115 3279
rect 495 3276 499 3280
rect 695 3276 699 3280
rect 903 3276 907 3280
rect 1119 3276 1123 3280
rect 1343 3276 1347 3280
rect 1935 3275 1939 3279
rect 1975 3264 1979 3268
rect 1995 3263 1999 3267
rect 2195 3263 2199 3267
rect 2411 3263 2415 3267
rect 2619 3263 2623 3267
rect 2811 3263 2815 3267
rect 3003 3263 3007 3267
rect 3187 3263 3191 3267
rect 3371 3263 3375 3267
rect 3555 3263 3559 3267
rect 3799 3264 3803 3268
rect 1975 3247 1979 3251
rect 2023 3248 2027 3252
rect 2223 3248 2227 3252
rect 2439 3248 2443 3252
rect 2647 3248 2651 3252
rect 2839 3248 2843 3252
rect 3031 3248 3035 3252
rect 3215 3248 3219 3252
rect 3399 3248 3403 3252
rect 3583 3248 3587 3252
rect 3799 3247 3803 3251
rect 111 3217 115 3221
rect 535 3216 539 3220
rect 727 3216 731 3220
rect 919 3216 923 3220
rect 1111 3216 1115 3220
rect 1295 3216 1299 3220
rect 1471 3216 1475 3220
rect 1655 3216 1659 3220
rect 1815 3216 1819 3220
rect 1935 3217 1939 3221
rect 3839 3216 3843 3220
rect 3859 3215 3863 3219
rect 4099 3215 4103 3219
rect 4347 3215 4351 3219
rect 4579 3215 4583 3219
rect 4787 3215 4791 3219
rect 4987 3215 4991 3219
rect 5171 3215 5175 3219
rect 5355 3215 5359 3219
rect 5515 3215 5519 3219
rect 5663 3216 5667 3220
rect 111 3200 115 3204
rect 507 3201 511 3205
rect 699 3201 703 3205
rect 891 3201 895 3205
rect 1083 3201 1087 3205
rect 1267 3201 1271 3205
rect 1443 3201 1447 3205
rect 1627 3201 1631 3205
rect 1787 3201 1791 3205
rect 1935 3200 1939 3204
rect 3839 3199 3843 3203
rect 3887 3200 3891 3204
rect 4127 3200 4131 3204
rect 4375 3200 4379 3204
rect 4607 3200 4611 3204
rect 4815 3200 4819 3204
rect 5015 3200 5019 3204
rect 5199 3200 5203 3204
rect 5383 3200 5387 3204
rect 5543 3200 5547 3204
rect 5663 3199 5667 3203
rect 1975 3189 1979 3193
rect 2463 3188 2467 3192
rect 2663 3188 2667 3192
rect 2863 3188 2867 3192
rect 3055 3188 3059 3192
rect 3239 3188 3243 3192
rect 3431 3188 3435 3192
rect 3623 3188 3627 3192
rect 3799 3189 3803 3193
rect 1975 3172 1979 3176
rect 2435 3173 2439 3177
rect 2635 3173 2639 3177
rect 2835 3173 2839 3177
rect 3027 3173 3031 3177
rect 3211 3173 3215 3177
rect 3403 3173 3407 3177
rect 3595 3173 3599 3177
rect 3799 3172 3803 3176
rect 3839 3125 3843 3129
rect 3903 3124 3907 3128
rect 4135 3124 4139 3128
rect 4359 3124 4363 3128
rect 4583 3124 4587 3128
rect 4807 3124 4811 3128
rect 5031 3124 5035 3128
rect 5663 3125 5667 3129
rect 3839 3108 3843 3112
rect 3875 3109 3879 3113
rect 4107 3109 4111 3113
rect 4331 3109 4335 3113
rect 4555 3109 4559 3113
rect 4779 3109 4783 3113
rect 5003 3109 5007 3113
rect 5663 3108 5667 3112
rect 111 3060 115 3064
rect 427 3059 431 3063
rect 563 3059 567 3063
rect 699 3059 703 3063
rect 835 3059 839 3063
rect 971 3059 975 3063
rect 1107 3059 1111 3063
rect 1243 3059 1247 3063
rect 1379 3059 1383 3063
rect 1515 3059 1519 3063
rect 1651 3059 1655 3063
rect 1787 3059 1791 3063
rect 1935 3060 1939 3064
rect 111 3043 115 3047
rect 455 3044 459 3048
rect 591 3044 595 3048
rect 727 3044 731 3048
rect 863 3044 867 3048
rect 999 3044 1003 3048
rect 1135 3044 1139 3048
rect 1271 3044 1275 3048
rect 1407 3044 1411 3048
rect 1543 3044 1547 3048
rect 1679 3044 1683 3048
rect 1815 3044 1819 3048
rect 1935 3043 1939 3047
rect 1975 3028 1979 3032
rect 2331 3027 2335 3031
rect 2555 3027 2559 3031
rect 2779 3027 2783 3031
rect 3003 3027 3007 3031
rect 3235 3027 3239 3031
rect 3467 3027 3471 3031
rect 3799 3028 3803 3032
rect 1975 3011 1979 3015
rect 2359 3012 2363 3016
rect 2583 3012 2587 3016
rect 2807 3012 2811 3016
rect 3031 3012 3035 3016
rect 3263 3012 3267 3016
rect 3495 3012 3499 3016
rect 3799 3011 3803 3015
rect 3839 2976 3843 2980
rect 3907 2975 3911 2979
rect 4075 2975 4079 2979
rect 4243 2975 4247 2979
rect 4411 2975 4415 2979
rect 4579 2975 4583 2979
rect 4755 2975 4759 2979
rect 5663 2976 5667 2980
rect 111 2957 115 2961
rect 199 2956 203 2960
rect 511 2956 515 2960
rect 815 2956 819 2960
rect 1111 2956 1115 2960
rect 1415 2956 1419 2960
rect 1719 2956 1723 2960
rect 1935 2957 1939 2961
rect 3839 2959 3843 2963
rect 3935 2960 3939 2964
rect 4103 2960 4107 2964
rect 4271 2960 4275 2964
rect 4439 2960 4443 2964
rect 4607 2960 4611 2964
rect 4783 2960 4787 2964
rect 5663 2959 5667 2963
rect 111 2940 115 2944
rect 171 2941 175 2945
rect 483 2941 487 2945
rect 787 2941 791 2945
rect 1083 2941 1087 2945
rect 1387 2941 1391 2945
rect 1691 2941 1695 2945
rect 1935 2940 1939 2944
rect 1975 2941 1979 2945
rect 2143 2940 2147 2944
rect 2343 2940 2347 2944
rect 2543 2940 2547 2944
rect 2743 2940 2747 2944
rect 2935 2940 2939 2944
rect 3135 2940 3139 2944
rect 3335 2940 3339 2944
rect 3799 2941 3803 2945
rect 1975 2924 1979 2928
rect 2115 2925 2119 2929
rect 2315 2925 2319 2929
rect 2515 2925 2519 2929
rect 2715 2925 2719 2929
rect 2907 2925 2911 2929
rect 3107 2925 3111 2929
rect 3307 2925 3311 2929
rect 3799 2924 3803 2928
rect 3839 2897 3843 2901
rect 3895 2896 3899 2900
rect 4031 2896 4035 2900
rect 4167 2896 4171 2900
rect 4303 2896 4307 2900
rect 4439 2896 4443 2900
rect 4575 2896 4579 2900
rect 5663 2897 5667 2901
rect 3839 2880 3843 2884
rect 3867 2881 3871 2885
rect 4003 2881 4007 2885
rect 4139 2881 4143 2885
rect 4275 2881 4279 2885
rect 4411 2881 4415 2885
rect 4547 2881 4551 2885
rect 5663 2880 5667 2884
rect 111 2808 115 2812
rect 131 2807 135 2811
rect 307 2807 311 2811
rect 523 2807 527 2811
rect 763 2807 767 2811
rect 1011 2807 1015 2811
rect 1275 2807 1279 2811
rect 1539 2807 1543 2811
rect 1935 2808 1939 2812
rect 111 2791 115 2795
rect 159 2792 163 2796
rect 335 2792 339 2796
rect 551 2792 555 2796
rect 791 2792 795 2796
rect 1039 2792 1043 2796
rect 1303 2792 1307 2796
rect 1567 2792 1571 2796
rect 1935 2791 1939 2795
rect 1975 2784 1979 2788
rect 2011 2783 2015 2787
rect 2259 2783 2263 2787
rect 2507 2783 2511 2787
rect 2755 2783 2759 2787
rect 3003 2783 3007 2787
rect 3799 2784 3803 2788
rect 1975 2767 1979 2771
rect 2039 2768 2043 2772
rect 2287 2768 2291 2772
rect 2535 2768 2539 2772
rect 2783 2768 2787 2772
rect 3031 2768 3035 2772
rect 3799 2767 3803 2771
rect 3839 2740 3843 2744
rect 3859 2739 3863 2743
rect 3995 2739 3999 2743
rect 4131 2739 4135 2743
rect 4267 2739 4271 2743
rect 4403 2739 4407 2743
rect 4539 2739 4543 2743
rect 4675 2739 4679 2743
rect 4811 2739 4815 2743
rect 5663 2740 5667 2744
rect 111 2729 115 2733
rect 279 2728 283 2732
rect 455 2728 459 2732
rect 647 2728 651 2732
rect 855 2728 859 2732
rect 1079 2728 1083 2732
rect 1311 2728 1315 2732
rect 1551 2728 1555 2732
rect 1799 2728 1803 2732
rect 1935 2729 1939 2733
rect 3839 2723 3843 2727
rect 3887 2724 3891 2728
rect 4023 2724 4027 2728
rect 4159 2724 4163 2728
rect 4295 2724 4299 2728
rect 4431 2724 4435 2728
rect 4567 2724 4571 2728
rect 4703 2724 4707 2728
rect 4839 2724 4843 2728
rect 5663 2723 5667 2727
rect 111 2712 115 2716
rect 251 2713 255 2717
rect 427 2713 431 2717
rect 619 2713 623 2717
rect 827 2713 831 2717
rect 1051 2713 1055 2717
rect 1283 2713 1287 2717
rect 1523 2713 1527 2717
rect 1771 2713 1775 2717
rect 1935 2712 1939 2716
rect 1975 2705 1979 2709
rect 2023 2704 2027 2708
rect 2247 2704 2251 2708
rect 2503 2704 2507 2708
rect 2759 2704 2763 2708
rect 3015 2704 3019 2708
rect 3799 2705 3803 2709
rect 1975 2688 1979 2692
rect 1995 2689 1999 2693
rect 2219 2689 2223 2693
rect 2475 2689 2479 2693
rect 2731 2689 2735 2693
rect 2987 2689 2991 2693
rect 3799 2688 3803 2692
rect 3839 2665 3843 2669
rect 3959 2664 3963 2668
rect 4255 2664 4259 2668
rect 4543 2664 4547 2668
rect 4823 2664 4827 2668
rect 5111 2664 5115 2668
rect 5399 2664 5403 2668
rect 5663 2665 5667 2669
rect 3839 2648 3843 2652
rect 3931 2649 3935 2653
rect 4227 2649 4231 2653
rect 4515 2649 4519 2653
rect 4795 2649 4799 2653
rect 5083 2649 5087 2653
rect 5371 2649 5375 2653
rect 5663 2648 5667 2652
rect 111 2580 115 2584
rect 571 2579 575 2583
rect 731 2579 735 2583
rect 891 2579 895 2583
rect 1043 2579 1047 2583
rect 1195 2579 1199 2583
rect 1355 2579 1359 2583
rect 1515 2579 1519 2583
rect 1675 2579 1679 2583
rect 1935 2580 1939 2584
rect 111 2563 115 2567
rect 599 2564 603 2568
rect 759 2564 763 2568
rect 919 2564 923 2568
rect 1071 2564 1075 2568
rect 1223 2564 1227 2568
rect 1383 2564 1387 2568
rect 1543 2564 1547 2568
rect 1703 2564 1707 2568
rect 1935 2563 1939 2567
rect 1975 2544 1979 2548
rect 2555 2543 2559 2547
rect 2691 2543 2695 2547
rect 2827 2543 2831 2547
rect 2963 2543 2967 2547
rect 3099 2543 3103 2547
rect 3799 2544 3803 2548
rect 1975 2527 1979 2531
rect 2583 2528 2587 2532
rect 2719 2528 2723 2532
rect 2855 2528 2859 2532
rect 2991 2528 2995 2532
rect 3127 2528 3131 2532
rect 3799 2527 3803 2531
rect 3839 2516 3843 2520
rect 3859 2515 3863 2519
rect 4083 2515 4087 2519
rect 4331 2515 4335 2519
rect 4579 2515 4583 2519
rect 4827 2515 4831 2519
rect 5075 2515 5079 2519
rect 5323 2515 5327 2519
rect 5663 2516 5667 2520
rect 111 2505 115 2509
rect 383 2504 387 2508
rect 599 2504 603 2508
rect 815 2504 819 2508
rect 1023 2504 1027 2508
rect 1231 2504 1235 2508
rect 1431 2504 1435 2508
rect 1631 2504 1635 2508
rect 1815 2504 1819 2508
rect 1935 2505 1939 2509
rect 3839 2499 3843 2503
rect 3887 2500 3891 2504
rect 4111 2500 4115 2504
rect 4359 2500 4363 2504
rect 4607 2500 4611 2504
rect 4855 2500 4859 2504
rect 5103 2500 5107 2504
rect 5351 2500 5355 2504
rect 5663 2499 5667 2503
rect 111 2488 115 2492
rect 355 2489 359 2493
rect 571 2489 575 2493
rect 787 2489 791 2493
rect 995 2489 999 2493
rect 1203 2489 1207 2493
rect 1403 2489 1407 2493
rect 1603 2489 1607 2493
rect 1787 2489 1791 2493
rect 1935 2488 1939 2492
rect 1975 2445 1979 2449
rect 2023 2444 2027 2448
rect 2223 2444 2227 2448
rect 2447 2444 2451 2448
rect 2679 2444 2683 2448
rect 2927 2444 2931 2448
rect 3183 2444 3187 2448
rect 3439 2444 3443 2448
rect 3679 2444 3683 2448
rect 3799 2445 3803 2449
rect 3839 2437 3843 2441
rect 3887 2436 3891 2440
rect 4087 2436 4091 2440
rect 4327 2436 4331 2440
rect 4583 2436 4587 2440
rect 4847 2436 4851 2440
rect 5119 2436 5123 2440
rect 5399 2436 5403 2440
rect 5663 2437 5667 2441
rect 1975 2428 1979 2432
rect 1995 2429 1999 2433
rect 2195 2429 2199 2433
rect 2419 2429 2423 2433
rect 2651 2429 2655 2433
rect 2899 2429 2903 2433
rect 3155 2429 3159 2433
rect 3411 2429 3415 2433
rect 3651 2429 3655 2433
rect 3799 2428 3803 2432
rect 3839 2420 3843 2424
rect 3859 2421 3863 2425
rect 4059 2421 4063 2425
rect 4299 2421 4303 2425
rect 4555 2421 4559 2425
rect 4819 2421 4823 2425
rect 5091 2421 5095 2425
rect 5371 2421 5375 2425
rect 5663 2420 5667 2424
rect 111 2352 115 2356
rect 227 2351 231 2355
rect 523 2351 527 2355
rect 835 2351 839 2355
rect 1155 2351 1159 2355
rect 1483 2351 1487 2355
rect 1787 2351 1791 2355
rect 1935 2352 1939 2356
rect 111 2335 115 2339
rect 255 2336 259 2340
rect 551 2336 555 2340
rect 863 2336 867 2340
rect 1183 2336 1187 2340
rect 1511 2336 1515 2340
rect 1815 2336 1819 2340
rect 1935 2335 1939 2339
rect 1975 2288 1979 2292
rect 1995 2287 1999 2291
rect 2155 2287 2159 2291
rect 2347 2287 2351 2291
rect 2539 2287 2543 2291
rect 2731 2287 2735 2291
rect 2923 2287 2927 2291
rect 3115 2287 3119 2291
rect 3299 2287 3303 2291
rect 3483 2287 3487 2291
rect 3651 2287 3655 2291
rect 3799 2288 3803 2292
rect 1975 2271 1979 2275
rect 2023 2272 2027 2276
rect 2183 2272 2187 2276
rect 2375 2272 2379 2276
rect 2567 2272 2571 2276
rect 2759 2272 2763 2276
rect 2951 2272 2955 2276
rect 3143 2272 3147 2276
rect 3327 2272 3331 2276
rect 3511 2272 3515 2276
rect 3839 2276 3843 2280
rect 3679 2272 3683 2276
rect 4443 2275 4447 2279
rect 3799 2271 3803 2275
rect 4611 2275 4615 2279
rect 4787 2275 4791 2279
rect 4963 2275 4967 2279
rect 5147 2275 5151 2279
rect 5339 2275 5343 2279
rect 5515 2275 5519 2279
rect 5663 2276 5667 2280
rect 111 2261 115 2265
rect 159 2260 163 2264
rect 367 2260 371 2264
rect 599 2260 603 2264
rect 831 2260 835 2264
rect 1063 2260 1067 2264
rect 1935 2261 1939 2265
rect 3839 2259 3843 2263
rect 4471 2260 4475 2264
rect 4639 2260 4643 2264
rect 4815 2260 4819 2264
rect 4991 2260 4995 2264
rect 5175 2260 5179 2264
rect 5367 2260 5371 2264
rect 5543 2260 5547 2264
rect 5663 2259 5667 2263
rect 111 2244 115 2248
rect 131 2245 135 2249
rect 339 2245 343 2249
rect 571 2245 575 2249
rect 803 2245 807 2249
rect 1035 2245 1039 2249
rect 1935 2244 1939 2248
rect 1975 2205 1979 2209
rect 2023 2204 2027 2208
rect 2191 2204 2195 2208
rect 2359 2204 2363 2208
rect 2535 2204 2539 2208
rect 2711 2204 2715 2208
rect 2879 2204 2883 2208
rect 3047 2204 3051 2208
rect 3207 2204 3211 2208
rect 3367 2204 3371 2208
rect 3535 2204 3539 2208
rect 3679 2204 3683 2208
rect 3799 2205 3803 2209
rect 1975 2188 1979 2192
rect 1995 2189 1999 2193
rect 2163 2189 2167 2193
rect 2331 2189 2335 2193
rect 2507 2189 2511 2193
rect 2683 2189 2687 2193
rect 2851 2189 2855 2193
rect 3019 2189 3023 2193
rect 3179 2189 3183 2193
rect 3339 2189 3343 2193
rect 3507 2189 3511 2193
rect 3651 2189 3655 2193
rect 3799 2188 3803 2192
rect 3839 2189 3843 2193
rect 4543 2188 4547 2192
rect 4719 2188 4723 2192
rect 4911 2188 4915 2192
rect 5119 2188 5123 2192
rect 5335 2188 5339 2192
rect 5543 2188 5547 2192
rect 5663 2189 5667 2193
rect 3839 2172 3843 2176
rect 4515 2173 4519 2177
rect 4691 2173 4695 2177
rect 4883 2173 4887 2177
rect 5091 2173 5095 2177
rect 5307 2173 5311 2177
rect 5515 2173 5519 2177
rect 5663 2172 5667 2176
rect 111 2100 115 2104
rect 131 2099 135 2103
rect 347 2099 351 2103
rect 595 2099 599 2103
rect 835 2099 839 2103
rect 1075 2099 1079 2103
rect 1315 2099 1319 2103
rect 1563 2099 1567 2103
rect 1787 2099 1791 2103
rect 1935 2100 1939 2104
rect 111 2083 115 2087
rect 159 2084 163 2088
rect 375 2084 379 2088
rect 623 2084 627 2088
rect 863 2084 867 2088
rect 1103 2084 1107 2088
rect 1343 2084 1347 2088
rect 1591 2084 1595 2088
rect 1815 2084 1819 2088
rect 1935 2083 1939 2087
rect 1975 2040 1979 2044
rect 3107 2039 3111 2043
rect 3243 2039 3247 2043
rect 3379 2039 3383 2043
rect 3515 2039 3519 2043
rect 3651 2039 3655 2043
rect 3799 2040 3803 2044
rect 3839 2040 3843 2044
rect 4635 2039 4639 2043
rect 4771 2039 4775 2043
rect 4907 2039 4911 2043
rect 5043 2039 5047 2043
rect 5179 2039 5183 2043
rect 5663 2040 5667 2044
rect 111 2021 115 2025
rect 271 2020 275 2024
rect 407 2020 411 2024
rect 543 2020 547 2024
rect 687 2020 691 2024
rect 831 2020 835 2024
rect 975 2020 979 2024
rect 1119 2020 1123 2024
rect 1263 2020 1267 2024
rect 1407 2020 1411 2024
rect 1543 2020 1547 2024
rect 1679 2020 1683 2024
rect 1815 2020 1819 2024
rect 1935 2021 1939 2025
rect 1975 2023 1979 2027
rect 3135 2024 3139 2028
rect 3271 2024 3275 2028
rect 3407 2024 3411 2028
rect 3543 2024 3547 2028
rect 3679 2024 3683 2028
rect 3799 2023 3803 2027
rect 3839 2023 3843 2027
rect 4663 2024 4667 2028
rect 4799 2024 4803 2028
rect 4935 2024 4939 2028
rect 5071 2024 5075 2028
rect 5207 2024 5211 2028
rect 5663 2023 5667 2027
rect 111 2004 115 2008
rect 243 2005 247 2009
rect 379 2005 383 2009
rect 515 2005 519 2009
rect 659 2005 663 2009
rect 803 2005 807 2009
rect 947 2005 951 2009
rect 1091 2005 1095 2009
rect 1235 2005 1239 2009
rect 1379 2005 1383 2009
rect 1515 2005 1519 2009
rect 1651 2005 1655 2009
rect 1787 2005 1791 2009
rect 1935 2004 1939 2008
rect 1975 1965 1979 1969
rect 3127 1964 3131 1968
rect 3263 1964 3267 1968
rect 3399 1964 3403 1968
rect 3535 1964 3539 1968
rect 3671 1964 3675 1968
rect 3799 1965 3803 1969
rect 3839 1965 3843 1969
rect 4863 1964 4867 1968
rect 4999 1964 5003 1968
rect 5135 1964 5139 1968
rect 5271 1964 5275 1968
rect 5407 1964 5411 1968
rect 5543 1964 5547 1968
rect 5663 1965 5667 1969
rect 1975 1948 1979 1952
rect 3099 1949 3103 1953
rect 3235 1949 3239 1953
rect 3371 1949 3375 1953
rect 3507 1949 3511 1953
rect 3643 1949 3647 1953
rect 3799 1948 3803 1952
rect 3839 1948 3843 1952
rect 4835 1949 4839 1953
rect 4971 1949 4975 1953
rect 5107 1949 5111 1953
rect 5243 1949 5247 1953
rect 5379 1949 5383 1953
rect 5515 1949 5519 1953
rect 5663 1948 5667 1952
rect 111 1868 115 1872
rect 187 1867 191 1871
rect 379 1867 383 1871
rect 587 1867 591 1871
rect 811 1867 815 1871
rect 1051 1867 1055 1871
rect 1299 1867 1303 1871
rect 1555 1867 1559 1871
rect 1787 1867 1791 1871
rect 1935 1868 1939 1872
rect 111 1851 115 1855
rect 215 1852 219 1856
rect 407 1852 411 1856
rect 615 1852 619 1856
rect 839 1852 843 1856
rect 1079 1852 1083 1856
rect 1327 1852 1331 1856
rect 1583 1852 1587 1856
rect 1815 1852 1819 1856
rect 1935 1851 1939 1855
rect 1975 1804 1979 1808
rect 1995 1803 1999 1807
rect 2227 1803 2231 1807
rect 2467 1803 2471 1807
rect 2691 1803 2695 1807
rect 2907 1803 2911 1807
rect 3107 1803 3111 1807
rect 3299 1803 3303 1807
rect 3483 1803 3487 1807
rect 3651 1803 3655 1807
rect 3799 1804 3803 1808
rect 3839 1804 3843 1808
rect 4675 1803 4679 1807
rect 4819 1803 4823 1807
rect 4963 1803 4967 1807
rect 5107 1803 5111 1807
rect 5243 1803 5247 1807
rect 5379 1803 5383 1807
rect 5515 1803 5519 1807
rect 5663 1804 5667 1808
rect 111 1785 115 1789
rect 159 1784 163 1788
rect 375 1784 379 1788
rect 591 1784 595 1788
rect 799 1784 803 1788
rect 999 1784 1003 1788
rect 1191 1784 1195 1788
rect 1383 1784 1387 1788
rect 1575 1784 1579 1788
rect 1935 1785 1939 1789
rect 1975 1787 1979 1791
rect 2023 1788 2027 1792
rect 2255 1788 2259 1792
rect 2495 1788 2499 1792
rect 2719 1788 2723 1792
rect 2935 1788 2939 1792
rect 3135 1788 3139 1792
rect 3327 1788 3331 1792
rect 3511 1788 3515 1792
rect 3679 1788 3683 1792
rect 3799 1787 3803 1791
rect 3839 1787 3843 1791
rect 4703 1788 4707 1792
rect 4847 1788 4851 1792
rect 4991 1788 4995 1792
rect 5135 1788 5139 1792
rect 5271 1788 5275 1792
rect 5407 1788 5411 1792
rect 5543 1788 5547 1792
rect 5663 1787 5667 1791
rect 111 1768 115 1772
rect 131 1769 135 1773
rect 347 1769 351 1773
rect 563 1769 567 1773
rect 771 1769 775 1773
rect 971 1769 975 1773
rect 1163 1769 1167 1773
rect 1355 1769 1359 1773
rect 1547 1769 1551 1773
rect 1935 1768 1939 1772
rect 1975 1721 1979 1725
rect 2023 1720 2027 1724
rect 2159 1720 2163 1724
rect 2311 1720 2315 1724
rect 2471 1720 2475 1724
rect 2639 1720 2643 1724
rect 2807 1720 2811 1724
rect 2975 1720 2979 1724
rect 3151 1720 3155 1724
rect 3799 1721 3803 1725
rect 3839 1713 3843 1717
rect 3887 1712 3891 1716
rect 4079 1712 4083 1716
rect 4303 1712 4307 1716
rect 4535 1712 4539 1716
rect 4775 1712 4779 1716
rect 5023 1712 5027 1716
rect 5279 1712 5283 1716
rect 5535 1712 5539 1716
rect 5663 1713 5667 1717
rect 1975 1704 1979 1708
rect 1995 1705 1999 1709
rect 2131 1705 2135 1709
rect 2283 1705 2287 1709
rect 2443 1705 2447 1709
rect 2611 1705 2615 1709
rect 2779 1705 2783 1709
rect 2947 1705 2951 1709
rect 3123 1705 3127 1709
rect 3799 1704 3803 1708
rect 3839 1696 3843 1700
rect 3859 1697 3863 1701
rect 4051 1697 4055 1701
rect 4275 1697 4279 1701
rect 4507 1697 4511 1701
rect 4747 1697 4751 1701
rect 4995 1697 4999 1701
rect 5251 1697 5255 1701
rect 5507 1697 5511 1701
rect 5663 1696 5667 1700
rect 111 1612 115 1616
rect 131 1611 135 1615
rect 395 1611 399 1615
rect 683 1611 687 1615
rect 979 1611 983 1615
rect 1275 1611 1279 1615
rect 1935 1612 1939 1616
rect 111 1595 115 1599
rect 159 1596 163 1600
rect 423 1596 427 1600
rect 711 1596 715 1600
rect 1007 1596 1011 1600
rect 1303 1596 1307 1600
rect 1935 1595 1939 1599
rect 1975 1564 1979 1568
rect 2091 1563 2095 1567
rect 2227 1563 2231 1567
rect 2363 1563 2367 1567
rect 2499 1563 2503 1567
rect 2635 1563 2639 1567
rect 2771 1563 2775 1567
rect 2907 1563 2911 1567
rect 3043 1563 3047 1567
rect 3179 1563 3183 1567
rect 3799 1564 3803 1568
rect 3839 1564 3843 1568
rect 3859 1563 3863 1567
rect 3995 1563 3999 1567
rect 4155 1563 4159 1567
rect 4355 1563 4359 1567
rect 4587 1563 4591 1567
rect 4851 1563 4855 1567
rect 5131 1563 5135 1567
rect 5419 1563 5423 1567
rect 5663 1564 5667 1568
rect 1975 1547 1979 1551
rect 2119 1548 2123 1552
rect 2255 1548 2259 1552
rect 2391 1548 2395 1552
rect 2527 1548 2531 1552
rect 2663 1548 2667 1552
rect 2799 1548 2803 1552
rect 2935 1548 2939 1552
rect 3071 1548 3075 1552
rect 3207 1548 3211 1552
rect 3799 1547 3803 1551
rect 3839 1547 3843 1551
rect 3887 1548 3891 1552
rect 4023 1548 4027 1552
rect 4183 1548 4187 1552
rect 4383 1548 4387 1552
rect 4615 1548 4619 1552
rect 4879 1548 4883 1552
rect 5159 1548 5163 1552
rect 5447 1548 5451 1552
rect 5663 1547 5667 1551
rect 111 1525 115 1529
rect 159 1524 163 1528
rect 375 1524 379 1528
rect 607 1524 611 1528
rect 839 1524 843 1528
rect 1071 1524 1075 1528
rect 1303 1524 1307 1528
rect 1935 1525 1939 1529
rect 111 1508 115 1512
rect 131 1509 135 1513
rect 347 1509 351 1513
rect 579 1509 583 1513
rect 811 1509 815 1513
rect 1043 1509 1047 1513
rect 1275 1509 1279 1513
rect 1935 1508 1939 1512
rect 3839 1489 3843 1493
rect 3887 1488 3891 1492
rect 4023 1488 4027 1492
rect 4159 1488 4163 1492
rect 4303 1488 4307 1492
rect 4495 1488 4499 1492
rect 4719 1488 4723 1492
rect 4967 1488 4971 1492
rect 5223 1488 5227 1492
rect 5487 1488 5491 1492
rect 5663 1489 5667 1493
rect 1975 1469 1979 1473
rect 2023 1468 2027 1472
rect 2159 1468 2163 1472
rect 2295 1468 2299 1472
rect 2431 1468 2435 1472
rect 2567 1468 2571 1472
rect 2703 1468 2707 1472
rect 2839 1468 2843 1472
rect 2975 1468 2979 1472
rect 3799 1469 3803 1473
rect 3839 1472 3843 1476
rect 3859 1473 3863 1477
rect 3995 1473 3999 1477
rect 4131 1473 4135 1477
rect 4275 1473 4279 1477
rect 4467 1473 4471 1477
rect 4691 1473 4695 1477
rect 4939 1473 4943 1477
rect 5195 1473 5199 1477
rect 5459 1473 5463 1477
rect 5663 1472 5667 1476
rect 1975 1452 1979 1456
rect 1995 1453 1999 1457
rect 2131 1453 2135 1457
rect 2267 1453 2271 1457
rect 2403 1453 2407 1457
rect 2539 1453 2543 1457
rect 2675 1453 2679 1457
rect 2811 1453 2815 1457
rect 2947 1453 2951 1457
rect 3799 1452 3803 1456
rect 111 1364 115 1368
rect 131 1363 135 1367
rect 411 1363 415 1367
rect 739 1363 743 1367
rect 1091 1363 1095 1367
rect 1451 1363 1455 1367
rect 1787 1363 1791 1367
rect 1935 1364 1939 1368
rect 111 1347 115 1351
rect 159 1348 163 1352
rect 439 1348 443 1352
rect 767 1348 771 1352
rect 1119 1348 1123 1352
rect 1479 1348 1483 1352
rect 1815 1348 1819 1352
rect 1935 1347 1939 1351
rect 3839 1336 3843 1340
rect 3859 1335 3863 1339
rect 4059 1335 4063 1339
rect 4307 1335 4311 1339
rect 4579 1335 4583 1339
rect 4875 1335 4879 1339
rect 5187 1335 5191 1339
rect 5499 1335 5503 1339
rect 5663 1336 5667 1340
rect 3839 1319 3843 1323
rect 3887 1320 3891 1324
rect 4087 1320 4091 1324
rect 4335 1320 4339 1324
rect 4607 1320 4611 1324
rect 4903 1320 4907 1324
rect 5215 1320 5219 1324
rect 5527 1320 5531 1324
rect 5663 1319 5667 1323
rect 1975 1312 1979 1316
rect 1995 1311 1999 1315
rect 2275 1311 2279 1315
rect 2563 1311 2567 1315
rect 2843 1311 2847 1315
rect 3123 1311 3127 1315
rect 3395 1311 3399 1315
rect 3651 1311 3655 1315
rect 3799 1312 3803 1316
rect 1975 1295 1979 1299
rect 2023 1296 2027 1300
rect 2303 1296 2307 1300
rect 2591 1296 2595 1300
rect 2871 1296 2875 1300
rect 3151 1296 3155 1300
rect 3423 1296 3427 1300
rect 3679 1296 3683 1300
rect 3799 1295 3803 1299
rect 111 1289 115 1293
rect 159 1288 163 1292
rect 359 1288 363 1292
rect 575 1288 579 1292
rect 775 1288 779 1292
rect 967 1288 971 1292
rect 1151 1288 1155 1292
rect 1327 1288 1331 1292
rect 1495 1288 1499 1292
rect 1663 1288 1667 1292
rect 1815 1288 1819 1292
rect 1935 1289 1939 1293
rect 111 1272 115 1276
rect 131 1273 135 1277
rect 331 1273 335 1277
rect 547 1273 551 1277
rect 747 1273 751 1277
rect 939 1273 943 1277
rect 1123 1273 1127 1277
rect 1299 1273 1303 1277
rect 1467 1273 1471 1277
rect 1635 1273 1639 1277
rect 1787 1273 1791 1277
rect 1935 1272 1939 1276
rect 3839 1253 3843 1257
rect 4615 1252 4619 1256
rect 4791 1252 4795 1256
rect 4975 1252 4979 1256
rect 5167 1252 5171 1256
rect 5367 1252 5371 1256
rect 5543 1252 5547 1256
rect 5663 1253 5667 1257
rect 3839 1236 3843 1240
rect 4587 1237 4591 1241
rect 4763 1237 4767 1241
rect 4947 1237 4951 1241
rect 5139 1237 5143 1241
rect 5339 1237 5343 1241
rect 5515 1237 5519 1241
rect 5663 1236 5667 1240
rect 1975 1213 1979 1217
rect 2655 1212 2659 1216
rect 2831 1212 2835 1216
rect 3007 1212 3011 1216
rect 3183 1212 3187 1216
rect 3359 1212 3363 1216
rect 3543 1212 3547 1216
rect 3799 1213 3803 1217
rect 1975 1196 1979 1200
rect 2627 1197 2631 1201
rect 2803 1197 2807 1201
rect 2979 1197 2983 1201
rect 3155 1197 3159 1201
rect 3331 1197 3335 1201
rect 3515 1197 3519 1201
rect 3799 1196 3803 1200
rect 111 1128 115 1132
rect 131 1127 135 1131
rect 291 1127 295 1131
rect 475 1127 479 1131
rect 659 1127 663 1131
rect 835 1127 839 1131
rect 1003 1127 1007 1131
rect 1171 1127 1175 1131
rect 1331 1127 1335 1131
rect 1491 1127 1495 1131
rect 1651 1127 1655 1131
rect 1787 1127 1791 1131
rect 1935 1128 1939 1132
rect 111 1111 115 1115
rect 159 1112 163 1116
rect 319 1112 323 1116
rect 503 1112 507 1116
rect 687 1112 691 1116
rect 863 1112 867 1116
rect 1031 1112 1035 1116
rect 1199 1112 1203 1116
rect 1359 1112 1363 1116
rect 1519 1112 1523 1116
rect 1679 1112 1683 1116
rect 1815 1112 1819 1116
rect 1935 1111 1939 1115
rect 3839 1100 3843 1104
rect 4835 1099 4839 1103
rect 4971 1099 4975 1103
rect 5107 1099 5111 1103
rect 5243 1099 5247 1103
rect 5379 1099 5383 1103
rect 5515 1099 5519 1103
rect 5663 1100 5667 1104
rect 3839 1083 3843 1087
rect 4863 1084 4867 1088
rect 4999 1084 5003 1088
rect 5135 1084 5139 1088
rect 5271 1084 5275 1088
rect 5407 1084 5411 1088
rect 5543 1084 5547 1088
rect 5663 1083 5667 1087
rect 1975 1048 1979 1052
rect 1995 1047 1999 1051
rect 2171 1047 2175 1051
rect 2363 1047 2367 1051
rect 2547 1047 2551 1051
rect 2723 1047 2727 1051
rect 2891 1047 2895 1051
rect 3059 1047 3063 1051
rect 3219 1047 3223 1051
rect 3387 1047 3391 1051
rect 3799 1048 3803 1052
rect 111 1041 115 1045
rect 175 1040 179 1044
rect 431 1040 435 1044
rect 687 1040 691 1044
rect 951 1040 955 1044
rect 1215 1040 1219 1044
rect 1935 1041 1939 1045
rect 1975 1031 1979 1035
rect 2023 1032 2027 1036
rect 2199 1032 2203 1036
rect 2391 1032 2395 1036
rect 2575 1032 2579 1036
rect 2751 1032 2755 1036
rect 2919 1032 2923 1036
rect 3087 1032 3091 1036
rect 3247 1032 3251 1036
rect 3415 1032 3419 1036
rect 3799 1031 3803 1035
rect 111 1024 115 1028
rect 147 1025 151 1029
rect 403 1025 407 1029
rect 659 1025 663 1029
rect 923 1025 927 1029
rect 1187 1025 1191 1029
rect 1935 1024 1939 1028
rect 3839 1021 3843 1025
rect 4807 1020 4811 1024
rect 4943 1020 4947 1024
rect 5079 1020 5083 1024
rect 5215 1020 5219 1024
rect 5351 1020 5355 1024
rect 5487 1020 5491 1024
rect 5663 1021 5667 1025
rect 3839 1004 3843 1008
rect 4779 1005 4783 1009
rect 4915 1005 4919 1009
rect 5051 1005 5055 1009
rect 5187 1005 5191 1009
rect 5323 1005 5327 1009
rect 5459 1005 5463 1009
rect 5663 1004 5667 1008
rect 1975 973 1979 977
rect 2023 972 2027 976
rect 2191 972 2195 976
rect 2375 972 2379 976
rect 2567 972 2571 976
rect 2759 972 2763 976
rect 2943 972 2947 976
rect 3127 972 3131 976
rect 3311 972 3315 976
rect 3495 972 3499 976
rect 3679 972 3683 976
rect 3799 973 3803 977
rect 1975 956 1979 960
rect 1995 957 1999 961
rect 2163 957 2167 961
rect 2347 957 2351 961
rect 2539 957 2543 961
rect 2731 957 2735 961
rect 2915 957 2919 961
rect 3099 957 3103 961
rect 3283 957 3287 961
rect 3467 957 3471 961
rect 3651 957 3655 961
rect 3799 956 3803 960
rect 111 880 115 884
rect 235 879 239 883
rect 459 879 463 883
rect 683 879 687 883
rect 907 879 911 883
rect 1131 879 1135 883
rect 1363 879 1367 883
rect 1935 880 1939 884
rect 111 863 115 867
rect 263 864 267 868
rect 487 864 491 868
rect 711 864 715 868
rect 935 864 939 868
rect 1159 864 1163 868
rect 3839 868 3843 872
rect 1391 864 1395 868
rect 3859 867 3863 871
rect 1935 863 1939 867
rect 3995 867 3999 871
rect 4171 867 4175 871
rect 4387 867 4391 871
rect 4643 867 4647 871
rect 4931 867 4935 871
rect 5235 867 5239 871
rect 5515 867 5519 871
rect 5663 868 5667 872
rect 3839 851 3843 855
rect 3887 852 3891 856
rect 4023 852 4027 856
rect 4199 852 4203 856
rect 4415 852 4419 856
rect 4671 852 4675 856
rect 4959 852 4963 856
rect 5263 852 5267 856
rect 5543 852 5547 856
rect 5663 851 5667 855
rect 1975 820 1979 824
rect 1995 819 1999 823
rect 2179 819 2183 823
rect 2403 819 2407 823
rect 2675 819 2679 823
rect 2987 819 2991 823
rect 3323 819 3327 823
rect 3651 819 3655 823
rect 3799 820 3803 824
rect 1975 803 1979 807
rect 2023 804 2027 808
rect 2207 804 2211 808
rect 2431 804 2435 808
rect 2703 804 2707 808
rect 3015 804 3019 808
rect 3351 804 3355 808
rect 3679 804 3683 808
rect 3799 803 3803 807
rect 111 789 115 793
rect 175 788 179 792
rect 431 788 435 792
rect 671 788 675 792
rect 903 788 907 792
rect 1127 788 1131 792
rect 1351 788 1355 792
rect 1575 788 1579 792
rect 1935 789 1939 793
rect 3839 793 3843 797
rect 3887 792 3891 796
rect 4023 792 4027 796
rect 4159 792 4163 796
rect 4295 792 4299 796
rect 4431 792 4435 796
rect 4567 792 4571 796
rect 4719 792 4723 796
rect 4895 792 4899 796
rect 5087 792 5091 796
rect 5287 792 5291 796
rect 5487 792 5491 796
rect 5663 793 5667 797
rect 111 772 115 776
rect 147 773 151 777
rect 403 773 407 777
rect 643 773 647 777
rect 875 773 879 777
rect 1099 773 1103 777
rect 1323 773 1327 777
rect 1547 773 1551 777
rect 1935 772 1939 776
rect 3839 776 3843 780
rect 3859 777 3863 781
rect 3995 777 3999 781
rect 4131 777 4135 781
rect 4267 777 4271 781
rect 4403 777 4407 781
rect 4539 777 4543 781
rect 4691 777 4695 781
rect 4867 777 4871 781
rect 5059 777 5063 781
rect 5259 777 5263 781
rect 5459 777 5463 781
rect 5663 776 5667 780
rect 111 640 115 644
rect 131 639 135 643
rect 315 639 319 643
rect 523 639 527 643
rect 723 639 727 643
rect 907 639 911 643
rect 1083 639 1087 643
rect 1259 639 1263 643
rect 1427 639 1431 643
rect 1595 639 1599 643
rect 1771 639 1775 643
rect 1935 640 1939 644
rect 3839 640 3843 644
rect 3859 639 3863 643
rect 3995 639 3999 643
rect 4131 639 4135 643
rect 4267 639 4271 643
rect 4403 639 4407 643
rect 4539 639 4543 643
rect 4699 639 4703 643
rect 4891 639 4895 643
rect 5099 639 5103 643
rect 5315 639 5319 643
rect 5515 639 5519 643
rect 5663 640 5667 644
rect 111 623 115 627
rect 159 624 163 628
rect 343 624 347 628
rect 551 624 555 628
rect 751 624 755 628
rect 935 624 939 628
rect 1111 624 1115 628
rect 1287 624 1291 628
rect 1455 624 1459 628
rect 1623 624 1627 628
rect 1799 624 1803 628
rect 1935 623 1939 627
rect 3839 623 3843 627
rect 3887 624 3891 628
rect 4023 624 4027 628
rect 4159 624 4163 628
rect 4295 624 4299 628
rect 4431 624 4435 628
rect 4567 624 4571 628
rect 4727 624 4731 628
rect 4919 624 4923 628
rect 5127 624 5131 628
rect 5343 624 5347 628
rect 5543 624 5547 628
rect 5663 623 5667 627
rect 111 565 115 569
rect 159 564 163 568
rect 375 564 379 568
rect 599 564 603 568
rect 807 564 811 568
rect 999 564 1003 568
rect 1175 564 1179 568
rect 1343 564 1347 568
rect 1511 564 1515 568
rect 1671 564 1675 568
rect 1815 564 1819 568
rect 1935 565 1939 569
rect 3839 565 3843 569
rect 3887 564 3891 568
rect 4071 564 4075 568
rect 4311 564 4315 568
rect 4575 564 4579 568
rect 4855 564 4859 568
rect 5151 564 5155 568
rect 5447 564 5451 568
rect 5663 565 5667 569
rect 111 548 115 552
rect 131 549 135 553
rect 347 549 351 553
rect 571 549 575 553
rect 779 549 783 553
rect 971 549 975 553
rect 1147 549 1151 553
rect 1315 549 1319 553
rect 1483 549 1487 553
rect 1643 549 1647 553
rect 1787 549 1791 553
rect 1935 548 1939 552
rect 1975 545 1979 549
rect 3135 544 3139 548
rect 3271 544 3275 548
rect 3407 544 3411 548
rect 3543 544 3547 548
rect 3679 544 3683 548
rect 3799 545 3803 549
rect 3839 548 3843 552
rect 3859 549 3863 553
rect 4043 549 4047 553
rect 4283 549 4287 553
rect 4547 549 4551 553
rect 4827 549 4831 553
rect 5123 549 5127 553
rect 5419 549 5423 553
rect 5663 548 5667 552
rect 1975 528 1979 532
rect 3107 529 3111 533
rect 3243 529 3247 533
rect 3379 529 3383 533
rect 3515 529 3519 533
rect 3651 529 3655 533
rect 3799 528 3803 532
rect 111 416 115 420
rect 155 415 159 419
rect 483 415 487 419
rect 811 415 815 419
rect 1139 415 1143 419
rect 1475 415 1479 419
rect 1787 415 1791 419
rect 1935 416 1939 420
rect 111 399 115 403
rect 183 400 187 404
rect 511 400 515 404
rect 839 400 843 404
rect 1167 400 1171 404
rect 1503 400 1507 404
rect 3839 404 3843 408
rect 1815 400 1819 404
rect 4451 403 4455 407
rect 1935 399 1939 403
rect 4643 403 4647 407
rect 4843 403 4847 407
rect 5051 403 5055 407
rect 5267 403 5271 407
rect 5483 403 5487 407
rect 5663 404 5667 408
rect 1975 396 1979 400
rect 1995 395 1999 399
rect 2203 395 2207 399
rect 2427 395 2431 399
rect 2651 395 2655 399
rect 2859 395 2863 399
rect 3067 395 3071 399
rect 3267 395 3271 399
rect 3467 395 3471 399
rect 3651 395 3655 399
rect 3799 396 3803 400
rect 3839 387 3843 391
rect 4479 388 4483 392
rect 4671 388 4675 392
rect 4871 388 4875 392
rect 5079 388 5083 392
rect 5295 388 5299 392
rect 5511 388 5515 392
rect 5663 387 5667 391
rect 1975 379 1979 383
rect 2023 380 2027 384
rect 2231 380 2235 384
rect 2455 380 2459 384
rect 2679 380 2683 384
rect 2887 380 2891 384
rect 3095 380 3099 384
rect 3295 380 3299 384
rect 3495 380 3499 384
rect 3679 380 3683 384
rect 3799 379 3803 383
rect 111 329 115 333
rect 279 328 283 332
rect 487 328 491 332
rect 703 328 707 332
rect 919 328 923 332
rect 1135 328 1139 332
rect 1935 329 1939 333
rect 3839 325 3843 329
rect 4615 324 4619 328
rect 4775 324 4779 328
rect 4951 324 4955 328
rect 5135 324 5139 328
rect 5327 324 5331 328
rect 5527 324 5531 328
rect 5663 325 5667 329
rect 111 312 115 316
rect 251 313 255 317
rect 459 313 463 317
rect 675 313 679 317
rect 891 313 895 317
rect 1107 313 1111 317
rect 1935 312 1939 316
rect 1975 305 1979 309
rect 2023 304 2027 308
rect 2159 304 2163 308
rect 2295 304 2299 308
rect 2431 304 2435 308
rect 2567 304 2571 308
rect 2703 304 2707 308
rect 2839 304 2843 308
rect 2975 304 2979 308
rect 3111 304 3115 308
rect 3247 304 3251 308
rect 3383 304 3387 308
rect 3519 304 3523 308
rect 3655 304 3659 308
rect 3799 305 3803 309
rect 3839 308 3843 312
rect 4587 309 4591 313
rect 4747 309 4751 313
rect 4923 309 4927 313
rect 5107 309 5111 313
rect 5299 309 5303 313
rect 5499 309 5503 313
rect 5663 308 5667 312
rect 1975 288 1979 292
rect 1995 289 1999 293
rect 2131 289 2135 293
rect 2267 289 2271 293
rect 2403 289 2407 293
rect 2539 289 2543 293
rect 2675 289 2679 293
rect 2811 289 2815 293
rect 2947 289 2951 293
rect 3083 289 3087 293
rect 3219 289 3223 293
rect 3355 289 3359 293
rect 3491 289 3495 293
rect 3627 289 3631 293
rect 3799 288 3803 292
rect 111 140 115 144
rect 131 139 135 143
rect 267 139 271 143
rect 403 139 407 143
rect 539 139 543 143
rect 675 139 679 143
rect 811 139 815 143
rect 947 139 951 143
rect 1083 139 1087 143
rect 1935 140 1939 144
rect 3839 136 3843 140
rect 4291 135 4295 139
rect 4427 135 4431 139
rect 4563 135 4567 139
rect 4699 135 4703 139
rect 4835 135 4839 139
rect 4971 135 4975 139
rect 5107 135 5111 139
rect 5243 135 5247 139
rect 5379 135 5383 139
rect 5515 135 5519 139
rect 5663 136 5667 140
rect 111 123 115 127
rect 159 124 163 128
rect 295 124 299 128
rect 431 124 435 128
rect 567 124 571 128
rect 703 124 707 128
rect 839 124 843 128
rect 975 124 979 128
rect 1111 124 1115 128
rect 1935 123 1939 127
rect 1975 120 1979 124
rect 1995 119 1999 123
rect 2131 119 2135 123
rect 2267 119 2271 123
rect 2403 119 2407 123
rect 2539 119 2543 123
rect 2675 119 2679 123
rect 2811 119 2815 123
rect 2947 119 2951 123
rect 3083 119 3087 123
rect 3219 119 3223 123
rect 3355 119 3359 123
rect 3491 119 3495 123
rect 3627 119 3631 123
rect 3799 120 3803 124
rect 3839 119 3843 123
rect 4319 120 4323 124
rect 4455 120 4459 124
rect 4591 120 4595 124
rect 4727 120 4731 124
rect 4863 120 4867 124
rect 4999 120 5003 124
rect 5135 120 5139 124
rect 5271 120 5275 124
rect 5407 120 5411 124
rect 5543 120 5547 124
rect 5663 119 5667 123
rect 1975 103 1979 107
rect 2023 104 2027 108
rect 2159 104 2163 108
rect 2295 104 2299 108
rect 2431 104 2435 108
rect 2567 104 2571 108
rect 2703 104 2707 108
rect 2839 104 2843 108
rect 2975 104 2979 108
rect 3111 104 3115 108
rect 3247 104 3251 108
rect 3383 104 3387 108
rect 3519 104 3523 108
rect 3655 104 3659 108
rect 3799 103 3803 107
<< m3 >>
rect 111 5758 115 5759
rect 111 5753 115 5754
rect 159 5758 163 5759
rect 159 5753 163 5754
rect 295 5758 299 5759
rect 295 5753 299 5754
rect 1935 5758 1939 5759
rect 1935 5753 1939 5754
rect 112 5730 114 5753
rect 110 5729 116 5730
rect 160 5729 162 5753
rect 296 5729 298 5753
rect 1936 5730 1938 5753
rect 1934 5729 1940 5730
rect 110 5725 111 5729
rect 115 5725 116 5729
rect 110 5724 116 5725
rect 158 5728 164 5729
rect 158 5724 159 5728
rect 163 5724 164 5728
rect 158 5723 164 5724
rect 294 5728 300 5729
rect 294 5724 295 5728
rect 299 5724 300 5728
rect 1934 5725 1935 5729
rect 1939 5725 1940 5729
rect 1934 5724 1940 5725
rect 294 5723 300 5724
rect 130 5713 136 5714
rect 110 5712 116 5713
rect 110 5708 111 5712
rect 115 5708 116 5712
rect 130 5709 131 5713
rect 135 5709 136 5713
rect 130 5708 136 5709
rect 266 5713 272 5714
rect 266 5709 267 5713
rect 271 5709 272 5713
rect 266 5708 272 5709
rect 1934 5712 1940 5713
rect 1934 5708 1935 5712
rect 1939 5708 1940 5712
rect 110 5707 116 5708
rect 112 5647 114 5707
rect 132 5647 134 5708
rect 268 5647 270 5708
rect 1934 5707 1940 5708
rect 1936 5647 1938 5707
rect 1975 5658 1979 5659
rect 1975 5653 1979 5654
rect 2023 5658 2027 5659
rect 2023 5653 2027 5654
rect 2183 5658 2187 5659
rect 2183 5653 2187 5654
rect 2367 5658 2371 5659
rect 2367 5653 2371 5654
rect 2551 5658 2555 5659
rect 2551 5653 2555 5654
rect 2727 5658 2731 5659
rect 2727 5653 2731 5654
rect 2895 5658 2899 5659
rect 2895 5653 2899 5654
rect 3063 5658 3067 5659
rect 3063 5653 3067 5654
rect 3223 5658 3227 5659
rect 3223 5653 3227 5654
rect 3383 5658 3387 5659
rect 3383 5653 3387 5654
rect 3543 5658 3547 5659
rect 3543 5653 3547 5654
rect 3679 5658 3683 5659
rect 3679 5653 3683 5654
rect 3799 5658 3803 5659
rect 3799 5653 3803 5654
rect 3839 5654 3843 5655
rect 111 5646 115 5647
rect 111 5641 115 5642
rect 131 5646 135 5647
rect 131 5641 135 5642
rect 267 5646 271 5647
rect 267 5641 271 5642
rect 275 5646 279 5647
rect 275 5641 279 5642
rect 475 5646 479 5647
rect 475 5641 479 5642
rect 699 5646 703 5647
rect 699 5641 703 5642
rect 955 5646 959 5647
rect 955 5641 959 5642
rect 1227 5646 1231 5647
rect 1227 5641 1231 5642
rect 1515 5646 1519 5647
rect 1515 5641 1519 5642
rect 1787 5646 1791 5647
rect 1787 5641 1791 5642
rect 1935 5646 1939 5647
rect 1935 5641 1939 5642
rect 112 5581 114 5641
rect 110 5580 116 5581
rect 132 5580 134 5641
rect 276 5580 278 5641
rect 476 5580 478 5641
rect 700 5580 702 5641
rect 956 5580 958 5641
rect 1228 5580 1230 5641
rect 1516 5580 1518 5641
rect 1788 5580 1790 5641
rect 1936 5581 1938 5641
rect 1976 5630 1978 5653
rect 1974 5629 1980 5630
rect 2024 5629 2026 5653
rect 2184 5629 2186 5653
rect 2368 5629 2370 5653
rect 2552 5629 2554 5653
rect 2728 5629 2730 5653
rect 2896 5629 2898 5653
rect 3064 5629 3066 5653
rect 3224 5629 3226 5653
rect 3384 5629 3386 5653
rect 3544 5629 3546 5653
rect 3680 5629 3682 5653
rect 3800 5630 3802 5653
rect 3839 5649 3843 5650
rect 4335 5654 4339 5655
rect 4335 5649 4339 5650
rect 4471 5654 4475 5655
rect 4471 5649 4475 5650
rect 4607 5654 4611 5655
rect 4607 5649 4611 5650
rect 4743 5654 4747 5655
rect 4743 5649 4747 5650
rect 4879 5654 4883 5655
rect 4879 5649 4883 5650
rect 5015 5654 5019 5655
rect 5015 5649 5019 5650
rect 5663 5654 5667 5655
rect 5663 5649 5667 5650
rect 3798 5629 3804 5630
rect 1974 5625 1975 5629
rect 1979 5625 1980 5629
rect 1974 5624 1980 5625
rect 2022 5628 2028 5629
rect 2022 5624 2023 5628
rect 2027 5624 2028 5628
rect 2022 5623 2028 5624
rect 2182 5628 2188 5629
rect 2182 5624 2183 5628
rect 2187 5624 2188 5628
rect 2182 5623 2188 5624
rect 2366 5628 2372 5629
rect 2366 5624 2367 5628
rect 2371 5624 2372 5628
rect 2366 5623 2372 5624
rect 2550 5628 2556 5629
rect 2550 5624 2551 5628
rect 2555 5624 2556 5628
rect 2550 5623 2556 5624
rect 2726 5628 2732 5629
rect 2726 5624 2727 5628
rect 2731 5624 2732 5628
rect 2726 5623 2732 5624
rect 2894 5628 2900 5629
rect 2894 5624 2895 5628
rect 2899 5624 2900 5628
rect 2894 5623 2900 5624
rect 3062 5628 3068 5629
rect 3062 5624 3063 5628
rect 3067 5624 3068 5628
rect 3062 5623 3068 5624
rect 3222 5628 3228 5629
rect 3222 5624 3223 5628
rect 3227 5624 3228 5628
rect 3222 5623 3228 5624
rect 3382 5628 3388 5629
rect 3382 5624 3383 5628
rect 3387 5624 3388 5628
rect 3382 5623 3388 5624
rect 3542 5628 3548 5629
rect 3542 5624 3543 5628
rect 3547 5624 3548 5628
rect 3542 5623 3548 5624
rect 3678 5628 3684 5629
rect 3678 5624 3679 5628
rect 3683 5624 3684 5628
rect 3798 5625 3799 5629
rect 3803 5625 3804 5629
rect 3840 5626 3842 5649
rect 3798 5624 3804 5625
rect 3838 5625 3844 5626
rect 4336 5625 4338 5649
rect 4472 5625 4474 5649
rect 4608 5625 4610 5649
rect 4744 5625 4746 5649
rect 4880 5625 4882 5649
rect 5016 5625 5018 5649
rect 5664 5626 5666 5649
rect 5662 5625 5668 5626
rect 3678 5623 3684 5624
rect 3838 5621 3839 5625
rect 3843 5621 3844 5625
rect 3838 5620 3844 5621
rect 4334 5624 4340 5625
rect 4334 5620 4335 5624
rect 4339 5620 4340 5624
rect 4334 5619 4340 5620
rect 4470 5624 4476 5625
rect 4470 5620 4471 5624
rect 4475 5620 4476 5624
rect 4470 5619 4476 5620
rect 4606 5624 4612 5625
rect 4606 5620 4607 5624
rect 4611 5620 4612 5624
rect 4606 5619 4612 5620
rect 4742 5624 4748 5625
rect 4742 5620 4743 5624
rect 4747 5620 4748 5624
rect 4742 5619 4748 5620
rect 4878 5624 4884 5625
rect 4878 5620 4879 5624
rect 4883 5620 4884 5624
rect 4878 5619 4884 5620
rect 5014 5624 5020 5625
rect 5014 5620 5015 5624
rect 5019 5620 5020 5624
rect 5662 5621 5663 5625
rect 5667 5621 5668 5625
rect 5662 5620 5668 5621
rect 5014 5619 5020 5620
rect 1994 5613 2000 5614
rect 1974 5612 1980 5613
rect 1974 5608 1975 5612
rect 1979 5608 1980 5612
rect 1994 5609 1995 5613
rect 1999 5609 2000 5613
rect 1994 5608 2000 5609
rect 2154 5613 2160 5614
rect 2154 5609 2155 5613
rect 2159 5609 2160 5613
rect 2154 5608 2160 5609
rect 2338 5613 2344 5614
rect 2338 5609 2339 5613
rect 2343 5609 2344 5613
rect 2338 5608 2344 5609
rect 2522 5613 2528 5614
rect 2522 5609 2523 5613
rect 2527 5609 2528 5613
rect 2522 5608 2528 5609
rect 2698 5613 2704 5614
rect 2698 5609 2699 5613
rect 2703 5609 2704 5613
rect 2698 5608 2704 5609
rect 2866 5613 2872 5614
rect 2866 5609 2867 5613
rect 2871 5609 2872 5613
rect 2866 5608 2872 5609
rect 3034 5613 3040 5614
rect 3034 5609 3035 5613
rect 3039 5609 3040 5613
rect 3034 5608 3040 5609
rect 3194 5613 3200 5614
rect 3194 5609 3195 5613
rect 3199 5609 3200 5613
rect 3194 5608 3200 5609
rect 3354 5613 3360 5614
rect 3354 5609 3355 5613
rect 3359 5609 3360 5613
rect 3354 5608 3360 5609
rect 3514 5613 3520 5614
rect 3514 5609 3515 5613
rect 3519 5609 3520 5613
rect 3514 5608 3520 5609
rect 3650 5613 3656 5614
rect 3650 5609 3651 5613
rect 3655 5609 3656 5613
rect 3650 5608 3656 5609
rect 3798 5612 3804 5613
rect 3798 5608 3799 5612
rect 3803 5608 3804 5612
rect 4306 5609 4312 5610
rect 1974 5607 1980 5608
rect 1934 5580 1940 5581
rect 110 5576 111 5580
rect 115 5576 116 5580
rect 110 5575 116 5576
rect 130 5579 136 5580
rect 130 5575 131 5579
rect 135 5575 136 5579
rect 130 5574 136 5575
rect 274 5579 280 5580
rect 274 5575 275 5579
rect 279 5575 280 5579
rect 274 5574 280 5575
rect 474 5579 480 5580
rect 474 5575 475 5579
rect 479 5575 480 5579
rect 474 5574 480 5575
rect 698 5579 704 5580
rect 698 5575 699 5579
rect 703 5575 704 5579
rect 698 5574 704 5575
rect 954 5579 960 5580
rect 954 5575 955 5579
rect 959 5575 960 5579
rect 954 5574 960 5575
rect 1226 5579 1232 5580
rect 1226 5575 1227 5579
rect 1231 5575 1232 5579
rect 1226 5574 1232 5575
rect 1514 5579 1520 5580
rect 1514 5575 1515 5579
rect 1519 5575 1520 5579
rect 1514 5574 1520 5575
rect 1786 5579 1792 5580
rect 1786 5575 1787 5579
rect 1791 5575 1792 5579
rect 1934 5576 1935 5580
rect 1939 5576 1940 5580
rect 1934 5575 1940 5576
rect 1786 5574 1792 5575
rect 158 5564 164 5565
rect 110 5563 116 5564
rect 110 5559 111 5563
rect 115 5559 116 5563
rect 158 5560 159 5564
rect 163 5560 164 5564
rect 158 5559 164 5560
rect 302 5564 308 5565
rect 302 5560 303 5564
rect 307 5560 308 5564
rect 302 5559 308 5560
rect 502 5564 508 5565
rect 502 5560 503 5564
rect 507 5560 508 5564
rect 502 5559 508 5560
rect 726 5564 732 5565
rect 726 5560 727 5564
rect 731 5560 732 5564
rect 726 5559 732 5560
rect 982 5564 988 5565
rect 982 5560 983 5564
rect 987 5560 988 5564
rect 982 5559 988 5560
rect 1254 5564 1260 5565
rect 1254 5560 1255 5564
rect 1259 5560 1260 5564
rect 1254 5559 1260 5560
rect 1542 5564 1548 5565
rect 1542 5560 1543 5564
rect 1547 5560 1548 5564
rect 1542 5559 1548 5560
rect 1814 5564 1820 5565
rect 1814 5560 1815 5564
rect 1819 5560 1820 5564
rect 1814 5559 1820 5560
rect 1934 5563 1940 5564
rect 1934 5559 1935 5563
rect 1939 5559 1940 5563
rect 110 5558 116 5559
rect 112 5535 114 5558
rect 160 5535 162 5559
rect 304 5535 306 5559
rect 504 5535 506 5559
rect 728 5535 730 5559
rect 984 5535 986 5559
rect 1256 5535 1258 5559
rect 1544 5535 1546 5559
rect 1816 5535 1818 5559
rect 1934 5558 1940 5559
rect 1936 5535 1938 5558
rect 1976 5547 1978 5607
rect 1996 5547 1998 5608
rect 2156 5547 2158 5608
rect 2340 5547 2342 5608
rect 2524 5547 2526 5608
rect 2700 5547 2702 5608
rect 2868 5547 2870 5608
rect 3036 5547 3038 5608
rect 3196 5547 3198 5608
rect 3356 5547 3358 5608
rect 3516 5547 3518 5608
rect 3652 5547 3654 5608
rect 3798 5607 3804 5608
rect 3838 5608 3844 5609
rect 3800 5547 3802 5607
rect 3838 5604 3839 5608
rect 3843 5604 3844 5608
rect 4306 5605 4307 5609
rect 4311 5605 4312 5609
rect 4306 5604 4312 5605
rect 4442 5609 4448 5610
rect 4442 5605 4443 5609
rect 4447 5605 4448 5609
rect 4442 5604 4448 5605
rect 4578 5609 4584 5610
rect 4578 5605 4579 5609
rect 4583 5605 4584 5609
rect 4578 5604 4584 5605
rect 4714 5609 4720 5610
rect 4714 5605 4715 5609
rect 4719 5605 4720 5609
rect 4714 5604 4720 5605
rect 4850 5609 4856 5610
rect 4850 5605 4851 5609
rect 4855 5605 4856 5609
rect 4850 5604 4856 5605
rect 4986 5609 4992 5610
rect 4986 5605 4987 5609
rect 4991 5605 4992 5609
rect 4986 5604 4992 5605
rect 5662 5608 5668 5609
rect 5662 5604 5663 5608
rect 5667 5604 5668 5608
rect 3838 5603 3844 5604
rect 1975 5546 1979 5547
rect 1975 5541 1979 5542
rect 1995 5546 1999 5547
rect 1995 5541 1999 5542
rect 2139 5546 2143 5547
rect 2139 5541 2143 5542
rect 2155 5546 2159 5547
rect 2155 5541 2159 5542
rect 2339 5546 2343 5547
rect 2339 5541 2343 5542
rect 2355 5546 2359 5547
rect 2355 5541 2359 5542
rect 2523 5546 2527 5547
rect 2523 5541 2527 5542
rect 2563 5546 2567 5547
rect 2563 5541 2567 5542
rect 2699 5546 2703 5547
rect 2699 5541 2703 5542
rect 2755 5546 2759 5547
rect 2755 5541 2759 5542
rect 2867 5546 2871 5547
rect 2867 5541 2871 5542
rect 2939 5546 2943 5547
rect 2939 5541 2943 5542
rect 3035 5546 3039 5547
rect 3035 5541 3039 5542
rect 3115 5546 3119 5547
rect 3115 5541 3119 5542
rect 3195 5546 3199 5547
rect 3195 5541 3199 5542
rect 3291 5546 3295 5547
rect 3291 5541 3295 5542
rect 3355 5546 3359 5547
rect 3355 5541 3359 5542
rect 3467 5546 3471 5547
rect 3467 5541 3471 5542
rect 3515 5546 3519 5547
rect 3515 5541 3519 5542
rect 3643 5546 3647 5547
rect 3643 5541 3647 5542
rect 3651 5546 3655 5547
rect 3651 5541 3655 5542
rect 3799 5546 3803 5547
rect 3840 5543 3842 5603
rect 4308 5543 4310 5604
rect 4444 5543 4446 5604
rect 4580 5543 4582 5604
rect 4716 5543 4718 5604
rect 4852 5543 4854 5604
rect 4988 5543 4990 5604
rect 5662 5603 5668 5604
rect 5664 5543 5666 5603
rect 3799 5541 3803 5542
rect 3839 5542 3843 5543
rect 111 5534 115 5535
rect 111 5529 115 5530
rect 159 5534 163 5535
rect 159 5529 163 5530
rect 279 5534 283 5535
rect 279 5529 283 5530
rect 303 5534 307 5535
rect 303 5529 307 5530
rect 503 5534 507 5535
rect 503 5529 507 5530
rect 519 5534 523 5535
rect 519 5529 523 5530
rect 727 5534 731 5535
rect 727 5529 731 5530
rect 767 5534 771 5535
rect 767 5529 771 5530
rect 983 5534 987 5535
rect 983 5529 987 5530
rect 1015 5534 1019 5535
rect 1015 5529 1019 5530
rect 1255 5534 1259 5535
rect 1255 5529 1259 5530
rect 1263 5534 1267 5535
rect 1263 5529 1267 5530
rect 1511 5534 1515 5535
rect 1511 5529 1515 5530
rect 1543 5534 1547 5535
rect 1543 5529 1547 5530
rect 1767 5534 1771 5535
rect 1767 5529 1771 5530
rect 1815 5534 1819 5535
rect 1815 5529 1819 5530
rect 1935 5534 1939 5535
rect 1935 5529 1939 5530
rect 112 5506 114 5529
rect 110 5505 116 5506
rect 280 5505 282 5529
rect 520 5505 522 5529
rect 768 5505 770 5529
rect 1016 5505 1018 5529
rect 1264 5505 1266 5529
rect 1512 5505 1514 5529
rect 1768 5505 1770 5529
rect 1936 5506 1938 5529
rect 1934 5505 1940 5506
rect 110 5501 111 5505
rect 115 5501 116 5505
rect 110 5500 116 5501
rect 278 5504 284 5505
rect 278 5500 279 5504
rect 283 5500 284 5504
rect 278 5499 284 5500
rect 518 5504 524 5505
rect 518 5500 519 5504
rect 523 5500 524 5504
rect 518 5499 524 5500
rect 766 5504 772 5505
rect 766 5500 767 5504
rect 771 5500 772 5504
rect 766 5499 772 5500
rect 1014 5504 1020 5505
rect 1014 5500 1015 5504
rect 1019 5500 1020 5504
rect 1014 5499 1020 5500
rect 1262 5504 1268 5505
rect 1262 5500 1263 5504
rect 1267 5500 1268 5504
rect 1262 5499 1268 5500
rect 1510 5504 1516 5505
rect 1510 5500 1511 5504
rect 1515 5500 1516 5504
rect 1510 5499 1516 5500
rect 1766 5504 1772 5505
rect 1766 5500 1767 5504
rect 1771 5500 1772 5504
rect 1934 5501 1935 5505
rect 1939 5501 1940 5505
rect 1934 5500 1940 5501
rect 1766 5499 1772 5500
rect 250 5489 256 5490
rect 110 5488 116 5489
rect 110 5484 111 5488
rect 115 5484 116 5488
rect 250 5485 251 5489
rect 255 5485 256 5489
rect 250 5484 256 5485
rect 490 5489 496 5490
rect 490 5485 491 5489
rect 495 5485 496 5489
rect 490 5484 496 5485
rect 738 5489 744 5490
rect 738 5485 739 5489
rect 743 5485 744 5489
rect 738 5484 744 5485
rect 986 5489 992 5490
rect 986 5485 987 5489
rect 991 5485 992 5489
rect 986 5484 992 5485
rect 1234 5489 1240 5490
rect 1234 5485 1235 5489
rect 1239 5485 1240 5489
rect 1234 5484 1240 5485
rect 1482 5489 1488 5490
rect 1482 5485 1483 5489
rect 1487 5485 1488 5489
rect 1482 5484 1488 5485
rect 1738 5489 1744 5490
rect 1738 5485 1739 5489
rect 1743 5485 1744 5489
rect 1738 5484 1744 5485
rect 1934 5488 1940 5489
rect 1934 5484 1935 5488
rect 1939 5484 1940 5488
rect 110 5483 116 5484
rect 112 5423 114 5483
rect 252 5423 254 5484
rect 492 5423 494 5484
rect 740 5423 742 5484
rect 988 5423 990 5484
rect 1236 5423 1238 5484
rect 1484 5423 1486 5484
rect 1740 5423 1742 5484
rect 1934 5483 1940 5484
rect 1936 5423 1938 5483
rect 1976 5481 1978 5541
rect 1974 5480 1980 5481
rect 2140 5480 2142 5541
rect 2356 5480 2358 5541
rect 2564 5480 2566 5541
rect 2756 5480 2758 5541
rect 2940 5480 2942 5541
rect 3116 5480 3118 5541
rect 3292 5480 3294 5541
rect 3468 5480 3470 5541
rect 3644 5480 3646 5541
rect 3800 5481 3802 5541
rect 3839 5537 3843 5538
rect 4251 5542 4255 5543
rect 4251 5537 4255 5538
rect 4307 5542 4311 5543
rect 4307 5537 4311 5538
rect 4403 5542 4407 5543
rect 4403 5537 4407 5538
rect 4443 5542 4447 5543
rect 4443 5537 4447 5538
rect 4555 5542 4559 5543
rect 4555 5537 4559 5538
rect 4579 5542 4583 5543
rect 4579 5537 4583 5538
rect 4707 5542 4711 5543
rect 4707 5537 4711 5538
rect 4715 5542 4719 5543
rect 4715 5537 4719 5538
rect 4851 5542 4855 5543
rect 4851 5537 4855 5538
rect 4859 5542 4863 5543
rect 4859 5537 4863 5538
rect 4987 5542 4991 5543
rect 4987 5537 4991 5538
rect 5019 5542 5023 5543
rect 5019 5537 5023 5538
rect 5663 5542 5667 5543
rect 5663 5537 5667 5538
rect 3798 5480 3804 5481
rect 1974 5476 1975 5480
rect 1979 5476 1980 5480
rect 1974 5475 1980 5476
rect 2138 5479 2144 5480
rect 2138 5475 2139 5479
rect 2143 5475 2144 5479
rect 2138 5474 2144 5475
rect 2354 5479 2360 5480
rect 2354 5475 2355 5479
rect 2359 5475 2360 5479
rect 2354 5474 2360 5475
rect 2562 5479 2568 5480
rect 2562 5475 2563 5479
rect 2567 5475 2568 5479
rect 2562 5474 2568 5475
rect 2754 5479 2760 5480
rect 2754 5475 2755 5479
rect 2759 5475 2760 5479
rect 2754 5474 2760 5475
rect 2938 5479 2944 5480
rect 2938 5475 2939 5479
rect 2943 5475 2944 5479
rect 2938 5474 2944 5475
rect 3114 5479 3120 5480
rect 3114 5475 3115 5479
rect 3119 5475 3120 5479
rect 3114 5474 3120 5475
rect 3290 5479 3296 5480
rect 3290 5475 3291 5479
rect 3295 5475 3296 5479
rect 3290 5474 3296 5475
rect 3466 5479 3472 5480
rect 3466 5475 3467 5479
rect 3471 5475 3472 5479
rect 3466 5474 3472 5475
rect 3642 5479 3648 5480
rect 3642 5475 3643 5479
rect 3647 5475 3648 5479
rect 3798 5476 3799 5480
rect 3803 5476 3804 5480
rect 3840 5477 3842 5537
rect 3798 5475 3804 5476
rect 3838 5476 3844 5477
rect 4252 5476 4254 5537
rect 4404 5476 4406 5537
rect 4556 5476 4558 5537
rect 4708 5476 4710 5537
rect 4860 5476 4862 5537
rect 5020 5476 5022 5537
rect 5664 5477 5666 5537
rect 5662 5476 5668 5477
rect 3642 5474 3648 5475
rect 3838 5472 3839 5476
rect 3843 5472 3844 5476
rect 3838 5471 3844 5472
rect 4250 5475 4256 5476
rect 4250 5471 4251 5475
rect 4255 5471 4256 5475
rect 4250 5470 4256 5471
rect 4402 5475 4408 5476
rect 4402 5471 4403 5475
rect 4407 5471 4408 5475
rect 4402 5470 4408 5471
rect 4554 5475 4560 5476
rect 4554 5471 4555 5475
rect 4559 5471 4560 5475
rect 4554 5470 4560 5471
rect 4706 5475 4712 5476
rect 4706 5471 4707 5475
rect 4711 5471 4712 5475
rect 4706 5470 4712 5471
rect 4858 5475 4864 5476
rect 4858 5471 4859 5475
rect 4863 5471 4864 5475
rect 4858 5470 4864 5471
rect 5018 5475 5024 5476
rect 5018 5471 5019 5475
rect 5023 5471 5024 5475
rect 5662 5472 5663 5476
rect 5667 5472 5668 5476
rect 5662 5471 5668 5472
rect 5018 5470 5024 5471
rect 2166 5464 2172 5465
rect 1974 5463 1980 5464
rect 1974 5459 1975 5463
rect 1979 5459 1980 5463
rect 2166 5460 2167 5464
rect 2171 5460 2172 5464
rect 2166 5459 2172 5460
rect 2382 5464 2388 5465
rect 2382 5460 2383 5464
rect 2387 5460 2388 5464
rect 2382 5459 2388 5460
rect 2590 5464 2596 5465
rect 2590 5460 2591 5464
rect 2595 5460 2596 5464
rect 2590 5459 2596 5460
rect 2782 5464 2788 5465
rect 2782 5460 2783 5464
rect 2787 5460 2788 5464
rect 2782 5459 2788 5460
rect 2966 5464 2972 5465
rect 2966 5460 2967 5464
rect 2971 5460 2972 5464
rect 2966 5459 2972 5460
rect 3142 5464 3148 5465
rect 3142 5460 3143 5464
rect 3147 5460 3148 5464
rect 3142 5459 3148 5460
rect 3318 5464 3324 5465
rect 3318 5460 3319 5464
rect 3323 5460 3324 5464
rect 3318 5459 3324 5460
rect 3494 5464 3500 5465
rect 3494 5460 3495 5464
rect 3499 5460 3500 5464
rect 3494 5459 3500 5460
rect 3670 5464 3676 5465
rect 3670 5460 3671 5464
rect 3675 5460 3676 5464
rect 3670 5459 3676 5460
rect 3798 5463 3804 5464
rect 3798 5459 3799 5463
rect 3803 5459 3804 5463
rect 4278 5460 4284 5461
rect 1974 5458 1980 5459
rect 1976 5427 1978 5458
rect 2168 5427 2170 5459
rect 2384 5427 2386 5459
rect 2592 5427 2594 5459
rect 2784 5427 2786 5459
rect 2968 5427 2970 5459
rect 3144 5427 3146 5459
rect 3320 5427 3322 5459
rect 3496 5427 3498 5459
rect 3672 5427 3674 5459
rect 3798 5458 3804 5459
rect 3838 5459 3844 5460
rect 3800 5427 3802 5458
rect 3838 5455 3839 5459
rect 3843 5455 3844 5459
rect 4278 5456 4279 5460
rect 4283 5456 4284 5460
rect 4278 5455 4284 5456
rect 4430 5460 4436 5461
rect 4430 5456 4431 5460
rect 4435 5456 4436 5460
rect 4430 5455 4436 5456
rect 4582 5460 4588 5461
rect 4582 5456 4583 5460
rect 4587 5456 4588 5460
rect 4582 5455 4588 5456
rect 4734 5460 4740 5461
rect 4734 5456 4735 5460
rect 4739 5456 4740 5460
rect 4734 5455 4740 5456
rect 4886 5460 4892 5461
rect 4886 5456 4887 5460
rect 4891 5456 4892 5460
rect 4886 5455 4892 5456
rect 5046 5460 5052 5461
rect 5046 5456 5047 5460
rect 5051 5456 5052 5460
rect 5046 5455 5052 5456
rect 5662 5459 5668 5460
rect 5662 5455 5663 5459
rect 5667 5455 5668 5459
rect 3838 5454 3844 5455
rect 1975 5426 1979 5427
rect 111 5422 115 5423
rect 111 5417 115 5418
rect 251 5422 255 5423
rect 251 5417 255 5418
rect 411 5422 415 5423
rect 411 5417 415 5418
rect 491 5422 495 5423
rect 491 5417 495 5418
rect 611 5422 615 5423
rect 611 5417 615 5418
rect 739 5422 743 5423
rect 739 5417 743 5418
rect 819 5422 823 5423
rect 819 5417 823 5418
rect 987 5422 991 5423
rect 987 5417 991 5418
rect 1035 5422 1039 5423
rect 1035 5417 1039 5418
rect 1235 5422 1239 5423
rect 1235 5417 1239 5418
rect 1259 5422 1263 5423
rect 1259 5417 1263 5418
rect 1483 5422 1487 5423
rect 1483 5417 1487 5418
rect 1491 5422 1495 5423
rect 1491 5417 1495 5418
rect 1739 5422 1743 5423
rect 1739 5417 1743 5418
rect 1935 5422 1939 5423
rect 1975 5421 1979 5422
rect 2167 5426 2171 5427
rect 2167 5421 2171 5422
rect 2311 5426 2315 5427
rect 2311 5421 2315 5422
rect 2383 5426 2387 5427
rect 2383 5421 2387 5422
rect 2511 5426 2515 5427
rect 2511 5421 2515 5422
rect 2591 5426 2595 5427
rect 2591 5421 2595 5422
rect 2703 5426 2707 5427
rect 2703 5421 2707 5422
rect 2783 5426 2787 5427
rect 2783 5421 2787 5422
rect 2887 5426 2891 5427
rect 2887 5421 2891 5422
rect 2967 5426 2971 5427
rect 2967 5421 2971 5422
rect 3071 5426 3075 5427
rect 3071 5421 3075 5422
rect 3143 5426 3147 5427
rect 3143 5421 3147 5422
rect 3247 5426 3251 5427
rect 3247 5421 3251 5422
rect 3319 5426 3323 5427
rect 3319 5421 3323 5422
rect 3423 5426 3427 5427
rect 3423 5421 3427 5422
rect 3495 5426 3499 5427
rect 3495 5421 3499 5422
rect 3607 5426 3611 5427
rect 3607 5421 3611 5422
rect 3671 5426 3675 5427
rect 3671 5421 3675 5422
rect 3799 5426 3803 5427
rect 3799 5421 3803 5422
rect 1935 5417 1939 5418
rect 112 5357 114 5417
rect 110 5356 116 5357
rect 412 5356 414 5417
rect 612 5356 614 5417
rect 820 5356 822 5417
rect 1036 5356 1038 5417
rect 1260 5356 1262 5417
rect 1492 5356 1494 5417
rect 1936 5357 1938 5417
rect 1976 5398 1978 5421
rect 1974 5397 1980 5398
rect 2312 5397 2314 5421
rect 2512 5397 2514 5421
rect 2704 5397 2706 5421
rect 2888 5397 2890 5421
rect 3072 5397 3074 5421
rect 3248 5397 3250 5421
rect 3424 5397 3426 5421
rect 3608 5397 3610 5421
rect 3800 5398 3802 5421
rect 3840 5411 3842 5454
rect 4280 5411 4282 5455
rect 4432 5411 4434 5455
rect 4584 5411 4586 5455
rect 4736 5411 4738 5455
rect 4888 5411 4890 5455
rect 5048 5411 5050 5455
rect 5662 5454 5668 5455
rect 5664 5411 5666 5454
rect 3839 5410 3843 5411
rect 3839 5405 3843 5406
rect 4279 5410 4283 5411
rect 4279 5405 4283 5406
rect 4431 5410 4435 5411
rect 4431 5405 4435 5406
rect 4487 5410 4491 5411
rect 4487 5405 4491 5406
rect 4583 5410 4587 5411
rect 4583 5405 4587 5406
rect 4695 5410 4699 5411
rect 4695 5405 4699 5406
rect 4735 5410 4739 5411
rect 4735 5405 4739 5406
rect 4887 5410 4891 5411
rect 4887 5405 4891 5406
rect 4911 5410 4915 5411
rect 4911 5405 4915 5406
rect 5047 5410 5051 5411
rect 5047 5405 5051 5406
rect 5127 5410 5131 5411
rect 5127 5405 5131 5406
rect 5663 5410 5667 5411
rect 5663 5405 5667 5406
rect 3798 5397 3804 5398
rect 1974 5393 1975 5397
rect 1979 5393 1980 5397
rect 1974 5392 1980 5393
rect 2310 5396 2316 5397
rect 2310 5392 2311 5396
rect 2315 5392 2316 5396
rect 2310 5391 2316 5392
rect 2510 5396 2516 5397
rect 2510 5392 2511 5396
rect 2515 5392 2516 5396
rect 2510 5391 2516 5392
rect 2702 5396 2708 5397
rect 2702 5392 2703 5396
rect 2707 5392 2708 5396
rect 2702 5391 2708 5392
rect 2886 5396 2892 5397
rect 2886 5392 2887 5396
rect 2891 5392 2892 5396
rect 2886 5391 2892 5392
rect 3070 5396 3076 5397
rect 3070 5392 3071 5396
rect 3075 5392 3076 5396
rect 3070 5391 3076 5392
rect 3246 5396 3252 5397
rect 3246 5392 3247 5396
rect 3251 5392 3252 5396
rect 3246 5391 3252 5392
rect 3422 5396 3428 5397
rect 3422 5392 3423 5396
rect 3427 5392 3428 5396
rect 3422 5391 3428 5392
rect 3606 5396 3612 5397
rect 3606 5392 3607 5396
rect 3611 5392 3612 5396
rect 3798 5393 3799 5397
rect 3803 5393 3804 5397
rect 3798 5392 3804 5393
rect 3606 5391 3612 5392
rect 3840 5382 3842 5405
rect 2282 5381 2288 5382
rect 1974 5380 1980 5381
rect 1974 5376 1975 5380
rect 1979 5376 1980 5380
rect 2282 5377 2283 5381
rect 2287 5377 2288 5381
rect 2282 5376 2288 5377
rect 2482 5381 2488 5382
rect 2482 5377 2483 5381
rect 2487 5377 2488 5381
rect 2482 5376 2488 5377
rect 2674 5381 2680 5382
rect 2674 5377 2675 5381
rect 2679 5377 2680 5381
rect 2674 5376 2680 5377
rect 2858 5381 2864 5382
rect 2858 5377 2859 5381
rect 2863 5377 2864 5381
rect 2858 5376 2864 5377
rect 3042 5381 3048 5382
rect 3042 5377 3043 5381
rect 3047 5377 3048 5381
rect 3042 5376 3048 5377
rect 3218 5381 3224 5382
rect 3218 5377 3219 5381
rect 3223 5377 3224 5381
rect 3218 5376 3224 5377
rect 3394 5381 3400 5382
rect 3394 5377 3395 5381
rect 3399 5377 3400 5381
rect 3394 5376 3400 5377
rect 3578 5381 3584 5382
rect 3838 5381 3844 5382
rect 4280 5381 4282 5405
rect 4488 5381 4490 5405
rect 4696 5381 4698 5405
rect 4912 5381 4914 5405
rect 5128 5381 5130 5405
rect 5664 5382 5666 5405
rect 5662 5381 5668 5382
rect 3578 5377 3579 5381
rect 3583 5377 3584 5381
rect 3578 5376 3584 5377
rect 3798 5380 3804 5381
rect 3798 5376 3799 5380
rect 3803 5376 3804 5380
rect 3838 5377 3839 5381
rect 3843 5377 3844 5381
rect 3838 5376 3844 5377
rect 4278 5380 4284 5381
rect 4278 5376 4279 5380
rect 4283 5376 4284 5380
rect 1974 5375 1980 5376
rect 1934 5356 1940 5357
rect 110 5352 111 5356
rect 115 5352 116 5356
rect 110 5351 116 5352
rect 410 5355 416 5356
rect 410 5351 411 5355
rect 415 5351 416 5355
rect 410 5350 416 5351
rect 610 5355 616 5356
rect 610 5351 611 5355
rect 615 5351 616 5355
rect 610 5350 616 5351
rect 818 5355 824 5356
rect 818 5351 819 5355
rect 823 5351 824 5355
rect 818 5350 824 5351
rect 1034 5355 1040 5356
rect 1034 5351 1035 5355
rect 1039 5351 1040 5355
rect 1034 5350 1040 5351
rect 1258 5355 1264 5356
rect 1258 5351 1259 5355
rect 1263 5351 1264 5355
rect 1258 5350 1264 5351
rect 1490 5355 1496 5356
rect 1490 5351 1491 5355
rect 1495 5351 1496 5355
rect 1934 5352 1935 5356
rect 1939 5352 1940 5356
rect 1934 5351 1940 5352
rect 1490 5350 1496 5351
rect 438 5340 444 5341
rect 110 5339 116 5340
rect 110 5335 111 5339
rect 115 5335 116 5339
rect 438 5336 439 5340
rect 443 5336 444 5340
rect 438 5335 444 5336
rect 638 5340 644 5341
rect 638 5336 639 5340
rect 643 5336 644 5340
rect 638 5335 644 5336
rect 846 5340 852 5341
rect 846 5336 847 5340
rect 851 5336 852 5340
rect 846 5335 852 5336
rect 1062 5340 1068 5341
rect 1062 5336 1063 5340
rect 1067 5336 1068 5340
rect 1062 5335 1068 5336
rect 1286 5340 1292 5341
rect 1286 5336 1287 5340
rect 1291 5336 1292 5340
rect 1286 5335 1292 5336
rect 1518 5340 1524 5341
rect 1518 5336 1519 5340
rect 1523 5336 1524 5340
rect 1518 5335 1524 5336
rect 1934 5339 1940 5340
rect 1934 5335 1935 5339
rect 1939 5335 1940 5339
rect 110 5334 116 5335
rect 112 5311 114 5334
rect 440 5311 442 5335
rect 640 5311 642 5335
rect 848 5311 850 5335
rect 1064 5311 1066 5335
rect 1288 5311 1290 5335
rect 1520 5311 1522 5335
rect 1934 5334 1940 5335
rect 1936 5311 1938 5334
rect 1976 5315 1978 5375
rect 2284 5315 2286 5376
rect 2484 5315 2486 5376
rect 2676 5315 2678 5376
rect 2860 5315 2862 5376
rect 3044 5315 3046 5376
rect 3220 5315 3222 5376
rect 3396 5315 3398 5376
rect 3580 5315 3582 5376
rect 3798 5375 3804 5376
rect 4278 5375 4284 5376
rect 4486 5380 4492 5381
rect 4486 5376 4487 5380
rect 4491 5376 4492 5380
rect 4486 5375 4492 5376
rect 4694 5380 4700 5381
rect 4694 5376 4695 5380
rect 4699 5376 4700 5380
rect 4694 5375 4700 5376
rect 4910 5380 4916 5381
rect 4910 5376 4911 5380
rect 4915 5376 4916 5380
rect 4910 5375 4916 5376
rect 5126 5380 5132 5381
rect 5126 5376 5127 5380
rect 5131 5376 5132 5380
rect 5662 5377 5663 5381
rect 5667 5377 5668 5381
rect 5662 5376 5668 5377
rect 5126 5375 5132 5376
rect 3800 5315 3802 5375
rect 4250 5365 4256 5366
rect 3838 5364 3844 5365
rect 3838 5360 3839 5364
rect 3843 5360 3844 5364
rect 4250 5361 4251 5365
rect 4255 5361 4256 5365
rect 4250 5360 4256 5361
rect 4458 5365 4464 5366
rect 4458 5361 4459 5365
rect 4463 5361 4464 5365
rect 4458 5360 4464 5361
rect 4666 5365 4672 5366
rect 4666 5361 4667 5365
rect 4671 5361 4672 5365
rect 4666 5360 4672 5361
rect 4882 5365 4888 5366
rect 4882 5361 4883 5365
rect 4887 5361 4888 5365
rect 4882 5360 4888 5361
rect 5098 5365 5104 5366
rect 5098 5361 5099 5365
rect 5103 5361 5104 5365
rect 5098 5360 5104 5361
rect 5662 5364 5668 5365
rect 5662 5360 5663 5364
rect 5667 5360 5668 5364
rect 3838 5359 3844 5360
rect 1975 5314 1979 5315
rect 111 5310 115 5311
rect 111 5305 115 5306
rect 439 5310 443 5311
rect 439 5305 443 5306
rect 591 5310 595 5311
rect 591 5305 595 5306
rect 639 5310 643 5311
rect 639 5305 643 5306
rect 727 5310 731 5311
rect 727 5305 731 5306
rect 847 5310 851 5311
rect 847 5305 851 5306
rect 863 5310 867 5311
rect 863 5305 867 5306
rect 999 5310 1003 5311
rect 999 5305 1003 5306
rect 1063 5310 1067 5311
rect 1063 5305 1067 5306
rect 1135 5310 1139 5311
rect 1135 5305 1139 5306
rect 1271 5310 1275 5311
rect 1271 5305 1275 5306
rect 1287 5310 1291 5311
rect 1287 5305 1291 5306
rect 1407 5310 1411 5311
rect 1407 5305 1411 5306
rect 1519 5310 1523 5311
rect 1519 5305 1523 5306
rect 1543 5310 1547 5311
rect 1543 5305 1547 5306
rect 1935 5310 1939 5311
rect 1975 5309 1979 5310
rect 2195 5314 2199 5315
rect 2195 5309 2199 5310
rect 2283 5314 2287 5315
rect 2283 5309 2287 5310
rect 2339 5314 2343 5315
rect 2339 5309 2343 5310
rect 2483 5314 2487 5315
rect 2483 5309 2487 5310
rect 2491 5314 2495 5315
rect 2491 5309 2495 5310
rect 2651 5314 2655 5315
rect 2651 5309 2655 5310
rect 2675 5314 2679 5315
rect 2675 5309 2679 5310
rect 2819 5314 2823 5315
rect 2819 5309 2823 5310
rect 2859 5314 2863 5315
rect 2859 5309 2863 5310
rect 3003 5314 3007 5315
rect 3003 5309 3007 5310
rect 3043 5314 3047 5315
rect 3043 5309 3047 5310
rect 3187 5314 3191 5315
rect 3187 5309 3191 5310
rect 3219 5314 3223 5315
rect 3219 5309 3223 5310
rect 3379 5314 3383 5315
rect 3379 5309 3383 5310
rect 3395 5314 3399 5315
rect 3395 5309 3399 5310
rect 3579 5314 3583 5315
rect 3579 5309 3583 5310
rect 3799 5314 3803 5315
rect 3799 5309 3803 5310
rect 1935 5305 1939 5306
rect 112 5282 114 5305
rect 110 5281 116 5282
rect 592 5281 594 5305
rect 728 5281 730 5305
rect 864 5281 866 5305
rect 1000 5281 1002 5305
rect 1136 5281 1138 5305
rect 1272 5281 1274 5305
rect 1408 5281 1410 5305
rect 1544 5281 1546 5305
rect 1936 5282 1938 5305
rect 1934 5281 1940 5282
rect 110 5277 111 5281
rect 115 5277 116 5281
rect 110 5276 116 5277
rect 590 5280 596 5281
rect 590 5276 591 5280
rect 595 5276 596 5280
rect 590 5275 596 5276
rect 726 5280 732 5281
rect 726 5276 727 5280
rect 731 5276 732 5280
rect 726 5275 732 5276
rect 862 5280 868 5281
rect 862 5276 863 5280
rect 867 5276 868 5280
rect 862 5275 868 5276
rect 998 5280 1004 5281
rect 998 5276 999 5280
rect 1003 5276 1004 5280
rect 998 5275 1004 5276
rect 1134 5280 1140 5281
rect 1134 5276 1135 5280
rect 1139 5276 1140 5280
rect 1134 5275 1140 5276
rect 1270 5280 1276 5281
rect 1270 5276 1271 5280
rect 1275 5276 1276 5280
rect 1270 5275 1276 5276
rect 1406 5280 1412 5281
rect 1406 5276 1407 5280
rect 1411 5276 1412 5280
rect 1406 5275 1412 5276
rect 1542 5280 1548 5281
rect 1542 5276 1543 5280
rect 1547 5276 1548 5280
rect 1934 5277 1935 5281
rect 1939 5277 1940 5281
rect 1934 5276 1940 5277
rect 1542 5275 1548 5276
rect 562 5265 568 5266
rect 110 5264 116 5265
rect 110 5260 111 5264
rect 115 5260 116 5264
rect 562 5261 563 5265
rect 567 5261 568 5265
rect 562 5260 568 5261
rect 698 5265 704 5266
rect 698 5261 699 5265
rect 703 5261 704 5265
rect 698 5260 704 5261
rect 834 5265 840 5266
rect 834 5261 835 5265
rect 839 5261 840 5265
rect 834 5260 840 5261
rect 970 5265 976 5266
rect 970 5261 971 5265
rect 975 5261 976 5265
rect 970 5260 976 5261
rect 1106 5265 1112 5266
rect 1106 5261 1107 5265
rect 1111 5261 1112 5265
rect 1106 5260 1112 5261
rect 1242 5265 1248 5266
rect 1242 5261 1243 5265
rect 1247 5261 1248 5265
rect 1242 5260 1248 5261
rect 1378 5265 1384 5266
rect 1378 5261 1379 5265
rect 1383 5261 1384 5265
rect 1378 5260 1384 5261
rect 1514 5265 1520 5266
rect 1514 5261 1515 5265
rect 1519 5261 1520 5265
rect 1514 5260 1520 5261
rect 1934 5264 1940 5265
rect 1934 5260 1935 5264
rect 1939 5260 1940 5264
rect 110 5259 116 5260
rect 112 5095 114 5259
rect 564 5095 566 5260
rect 700 5095 702 5260
rect 836 5095 838 5260
rect 972 5095 974 5260
rect 1108 5095 1110 5260
rect 1244 5095 1246 5260
rect 1380 5095 1382 5260
rect 1516 5095 1518 5260
rect 1934 5259 1940 5260
rect 1936 5095 1938 5259
rect 1976 5249 1978 5309
rect 1974 5248 1980 5249
rect 2196 5248 2198 5309
rect 2340 5248 2342 5309
rect 2492 5248 2494 5309
rect 2652 5248 2654 5309
rect 2820 5248 2822 5309
rect 3004 5248 3006 5309
rect 3188 5248 3190 5309
rect 3380 5248 3382 5309
rect 3580 5248 3582 5309
rect 3800 5249 3802 5309
rect 3840 5283 3842 5359
rect 4252 5283 4254 5360
rect 4460 5283 4462 5360
rect 4668 5283 4670 5360
rect 4884 5283 4886 5360
rect 5100 5283 5102 5360
rect 5662 5359 5668 5360
rect 5664 5283 5666 5359
rect 3839 5282 3843 5283
rect 3839 5277 3843 5278
rect 4251 5282 4255 5283
rect 4251 5277 4255 5278
rect 4459 5282 4463 5283
rect 4459 5277 4463 5278
rect 4483 5282 4487 5283
rect 4483 5277 4487 5278
rect 4667 5282 4671 5283
rect 4667 5277 4671 5278
rect 4715 5282 4719 5283
rect 4715 5277 4719 5278
rect 4883 5282 4887 5283
rect 4883 5277 4887 5278
rect 4947 5282 4951 5283
rect 4947 5277 4951 5278
rect 5099 5282 5103 5283
rect 5099 5277 5103 5278
rect 5187 5282 5191 5283
rect 5187 5277 5191 5278
rect 5663 5282 5667 5283
rect 5663 5277 5667 5278
rect 3798 5248 3804 5249
rect 1974 5244 1975 5248
rect 1979 5244 1980 5248
rect 1974 5243 1980 5244
rect 2194 5247 2200 5248
rect 2194 5243 2195 5247
rect 2199 5243 2200 5247
rect 2194 5242 2200 5243
rect 2338 5247 2344 5248
rect 2338 5243 2339 5247
rect 2343 5243 2344 5247
rect 2338 5242 2344 5243
rect 2490 5247 2496 5248
rect 2490 5243 2491 5247
rect 2495 5243 2496 5247
rect 2490 5242 2496 5243
rect 2650 5247 2656 5248
rect 2650 5243 2651 5247
rect 2655 5243 2656 5247
rect 2650 5242 2656 5243
rect 2818 5247 2824 5248
rect 2818 5243 2819 5247
rect 2823 5243 2824 5247
rect 2818 5242 2824 5243
rect 3002 5247 3008 5248
rect 3002 5243 3003 5247
rect 3007 5243 3008 5247
rect 3002 5242 3008 5243
rect 3186 5247 3192 5248
rect 3186 5243 3187 5247
rect 3191 5243 3192 5247
rect 3186 5242 3192 5243
rect 3378 5247 3384 5248
rect 3378 5243 3379 5247
rect 3383 5243 3384 5247
rect 3378 5242 3384 5243
rect 3578 5247 3584 5248
rect 3578 5243 3579 5247
rect 3583 5243 3584 5247
rect 3798 5244 3799 5248
rect 3803 5244 3804 5248
rect 3798 5243 3804 5244
rect 3578 5242 3584 5243
rect 2222 5232 2228 5233
rect 1974 5231 1980 5232
rect 1974 5227 1975 5231
rect 1979 5227 1980 5231
rect 2222 5228 2223 5232
rect 2227 5228 2228 5232
rect 2222 5227 2228 5228
rect 2366 5232 2372 5233
rect 2366 5228 2367 5232
rect 2371 5228 2372 5232
rect 2366 5227 2372 5228
rect 2518 5232 2524 5233
rect 2518 5228 2519 5232
rect 2523 5228 2524 5232
rect 2518 5227 2524 5228
rect 2678 5232 2684 5233
rect 2678 5228 2679 5232
rect 2683 5228 2684 5232
rect 2678 5227 2684 5228
rect 2846 5232 2852 5233
rect 2846 5228 2847 5232
rect 2851 5228 2852 5232
rect 2846 5227 2852 5228
rect 3030 5232 3036 5233
rect 3030 5228 3031 5232
rect 3035 5228 3036 5232
rect 3030 5227 3036 5228
rect 3214 5232 3220 5233
rect 3214 5228 3215 5232
rect 3219 5228 3220 5232
rect 3214 5227 3220 5228
rect 3406 5232 3412 5233
rect 3406 5228 3407 5232
rect 3411 5228 3412 5232
rect 3406 5227 3412 5228
rect 3606 5232 3612 5233
rect 3606 5228 3607 5232
rect 3611 5228 3612 5232
rect 3606 5227 3612 5228
rect 3798 5231 3804 5232
rect 3798 5227 3799 5231
rect 3803 5227 3804 5231
rect 1974 5226 1980 5227
rect 1976 5203 1978 5226
rect 2224 5203 2226 5227
rect 2368 5203 2370 5227
rect 2520 5203 2522 5227
rect 2680 5203 2682 5227
rect 2848 5203 2850 5227
rect 3032 5203 3034 5227
rect 3216 5203 3218 5227
rect 3408 5203 3410 5227
rect 3608 5203 3610 5227
rect 3798 5226 3804 5227
rect 3800 5203 3802 5226
rect 3840 5217 3842 5277
rect 3838 5216 3844 5217
rect 4252 5216 4254 5277
rect 4484 5216 4486 5277
rect 4716 5216 4718 5277
rect 4948 5216 4950 5277
rect 5188 5216 5190 5277
rect 5664 5217 5666 5277
rect 5662 5216 5668 5217
rect 3838 5212 3839 5216
rect 3843 5212 3844 5216
rect 3838 5211 3844 5212
rect 4250 5215 4256 5216
rect 4250 5211 4251 5215
rect 4255 5211 4256 5215
rect 4250 5210 4256 5211
rect 4482 5215 4488 5216
rect 4482 5211 4483 5215
rect 4487 5211 4488 5215
rect 4482 5210 4488 5211
rect 4714 5215 4720 5216
rect 4714 5211 4715 5215
rect 4719 5211 4720 5215
rect 4714 5210 4720 5211
rect 4946 5215 4952 5216
rect 4946 5211 4947 5215
rect 4951 5211 4952 5215
rect 4946 5210 4952 5211
rect 5186 5215 5192 5216
rect 5186 5211 5187 5215
rect 5191 5211 5192 5215
rect 5662 5212 5663 5216
rect 5667 5212 5668 5216
rect 5662 5211 5668 5212
rect 5186 5210 5192 5211
rect 1975 5202 1979 5203
rect 1975 5197 1979 5198
rect 2023 5202 2027 5203
rect 2023 5197 2027 5198
rect 2159 5202 2163 5203
rect 2159 5197 2163 5198
rect 2223 5202 2227 5203
rect 2223 5197 2227 5198
rect 2327 5202 2331 5203
rect 2327 5197 2331 5198
rect 2367 5202 2371 5203
rect 2367 5197 2371 5198
rect 2511 5202 2515 5203
rect 2511 5197 2515 5198
rect 2519 5202 2523 5203
rect 2519 5197 2523 5198
rect 2679 5202 2683 5203
rect 2679 5197 2683 5198
rect 2695 5202 2699 5203
rect 2695 5197 2699 5198
rect 2847 5202 2851 5203
rect 2847 5197 2851 5198
rect 2887 5202 2891 5203
rect 2887 5197 2891 5198
rect 3031 5202 3035 5203
rect 3031 5197 3035 5198
rect 3087 5202 3091 5203
rect 3087 5197 3091 5198
rect 3215 5202 3219 5203
rect 3215 5197 3219 5198
rect 3287 5202 3291 5203
rect 3287 5197 3291 5198
rect 3407 5202 3411 5203
rect 3407 5197 3411 5198
rect 3495 5202 3499 5203
rect 3495 5197 3499 5198
rect 3607 5202 3611 5203
rect 3607 5197 3611 5198
rect 3679 5202 3683 5203
rect 3679 5197 3683 5198
rect 3799 5202 3803 5203
rect 4278 5200 4284 5201
rect 3799 5197 3803 5198
rect 3838 5199 3844 5200
rect 1976 5174 1978 5197
rect 1974 5173 1980 5174
rect 2024 5173 2026 5197
rect 2160 5173 2162 5197
rect 2328 5173 2330 5197
rect 2512 5173 2514 5197
rect 2696 5173 2698 5197
rect 2888 5173 2890 5197
rect 3088 5173 3090 5197
rect 3288 5173 3290 5197
rect 3496 5173 3498 5197
rect 3680 5173 3682 5197
rect 3800 5174 3802 5197
rect 3838 5195 3839 5199
rect 3843 5195 3844 5199
rect 4278 5196 4279 5200
rect 4283 5196 4284 5200
rect 4278 5195 4284 5196
rect 4510 5200 4516 5201
rect 4510 5196 4511 5200
rect 4515 5196 4516 5200
rect 4510 5195 4516 5196
rect 4742 5200 4748 5201
rect 4742 5196 4743 5200
rect 4747 5196 4748 5200
rect 4742 5195 4748 5196
rect 4974 5200 4980 5201
rect 4974 5196 4975 5200
rect 4979 5196 4980 5200
rect 4974 5195 4980 5196
rect 5214 5200 5220 5201
rect 5214 5196 5215 5200
rect 5219 5196 5220 5200
rect 5214 5195 5220 5196
rect 5662 5199 5668 5200
rect 5662 5195 5663 5199
rect 5667 5195 5668 5199
rect 3838 5194 3844 5195
rect 3798 5173 3804 5174
rect 1974 5169 1975 5173
rect 1979 5169 1980 5173
rect 1974 5168 1980 5169
rect 2022 5172 2028 5173
rect 2022 5168 2023 5172
rect 2027 5168 2028 5172
rect 2022 5167 2028 5168
rect 2158 5172 2164 5173
rect 2158 5168 2159 5172
rect 2163 5168 2164 5172
rect 2158 5167 2164 5168
rect 2326 5172 2332 5173
rect 2326 5168 2327 5172
rect 2331 5168 2332 5172
rect 2326 5167 2332 5168
rect 2510 5172 2516 5173
rect 2510 5168 2511 5172
rect 2515 5168 2516 5172
rect 2510 5167 2516 5168
rect 2694 5172 2700 5173
rect 2694 5168 2695 5172
rect 2699 5168 2700 5172
rect 2694 5167 2700 5168
rect 2886 5172 2892 5173
rect 2886 5168 2887 5172
rect 2891 5168 2892 5172
rect 2886 5167 2892 5168
rect 3086 5172 3092 5173
rect 3086 5168 3087 5172
rect 3091 5168 3092 5172
rect 3086 5167 3092 5168
rect 3286 5172 3292 5173
rect 3286 5168 3287 5172
rect 3291 5168 3292 5172
rect 3286 5167 3292 5168
rect 3494 5172 3500 5173
rect 3494 5168 3495 5172
rect 3499 5168 3500 5172
rect 3494 5167 3500 5168
rect 3678 5172 3684 5173
rect 3678 5168 3679 5172
rect 3683 5168 3684 5172
rect 3798 5169 3799 5173
rect 3803 5169 3804 5173
rect 3798 5168 3804 5169
rect 3678 5167 3684 5168
rect 1994 5157 2000 5158
rect 1974 5156 1980 5157
rect 1974 5152 1975 5156
rect 1979 5152 1980 5156
rect 1994 5153 1995 5157
rect 1999 5153 2000 5157
rect 1994 5152 2000 5153
rect 2130 5157 2136 5158
rect 2130 5153 2131 5157
rect 2135 5153 2136 5157
rect 2130 5152 2136 5153
rect 2298 5157 2304 5158
rect 2298 5153 2299 5157
rect 2303 5153 2304 5157
rect 2298 5152 2304 5153
rect 2482 5157 2488 5158
rect 2482 5153 2483 5157
rect 2487 5153 2488 5157
rect 2482 5152 2488 5153
rect 2666 5157 2672 5158
rect 2666 5153 2667 5157
rect 2671 5153 2672 5157
rect 2666 5152 2672 5153
rect 2858 5157 2864 5158
rect 2858 5153 2859 5157
rect 2863 5153 2864 5157
rect 2858 5152 2864 5153
rect 3058 5157 3064 5158
rect 3058 5153 3059 5157
rect 3063 5153 3064 5157
rect 3058 5152 3064 5153
rect 3258 5157 3264 5158
rect 3258 5153 3259 5157
rect 3263 5153 3264 5157
rect 3258 5152 3264 5153
rect 3466 5157 3472 5158
rect 3466 5153 3467 5157
rect 3471 5153 3472 5157
rect 3466 5152 3472 5153
rect 3650 5157 3656 5158
rect 3650 5153 3651 5157
rect 3655 5153 3656 5157
rect 3650 5152 3656 5153
rect 3798 5156 3804 5157
rect 3798 5152 3799 5156
rect 3803 5152 3804 5156
rect 1974 5151 1980 5152
rect 111 5094 115 5095
rect 111 5089 115 5090
rect 347 5094 351 5095
rect 347 5089 351 5090
rect 483 5094 487 5095
rect 483 5089 487 5090
rect 563 5094 567 5095
rect 563 5089 567 5090
rect 619 5094 623 5095
rect 619 5089 623 5090
rect 699 5094 703 5095
rect 699 5089 703 5090
rect 755 5094 759 5095
rect 755 5089 759 5090
rect 835 5094 839 5095
rect 835 5089 839 5090
rect 891 5094 895 5095
rect 891 5089 895 5090
rect 971 5094 975 5095
rect 971 5089 975 5090
rect 1035 5094 1039 5095
rect 1035 5089 1039 5090
rect 1107 5094 1111 5095
rect 1107 5089 1111 5090
rect 1187 5094 1191 5095
rect 1187 5089 1191 5090
rect 1243 5094 1247 5095
rect 1243 5089 1247 5090
rect 1339 5094 1343 5095
rect 1339 5089 1343 5090
rect 1379 5094 1383 5095
rect 1379 5089 1383 5090
rect 1491 5094 1495 5095
rect 1491 5089 1495 5090
rect 1515 5094 1519 5095
rect 1515 5089 1519 5090
rect 1651 5094 1655 5095
rect 1651 5089 1655 5090
rect 1787 5094 1791 5095
rect 1787 5089 1791 5090
rect 1935 5094 1939 5095
rect 1976 5091 1978 5151
rect 1996 5091 1998 5152
rect 2132 5091 2134 5152
rect 2300 5091 2302 5152
rect 2484 5091 2486 5152
rect 2668 5091 2670 5152
rect 2860 5091 2862 5152
rect 3060 5091 3062 5152
rect 3260 5091 3262 5152
rect 3468 5091 3470 5152
rect 3652 5091 3654 5152
rect 3798 5151 3804 5152
rect 3800 5091 3802 5151
rect 3840 5143 3842 5194
rect 4280 5143 4282 5195
rect 4512 5143 4514 5195
rect 4744 5143 4746 5195
rect 4976 5143 4978 5195
rect 5216 5143 5218 5195
rect 5662 5194 5668 5195
rect 5664 5143 5666 5194
rect 3839 5142 3843 5143
rect 3839 5137 3843 5138
rect 3887 5142 3891 5143
rect 3887 5137 3891 5138
rect 4135 5142 4139 5143
rect 4135 5137 4139 5138
rect 4279 5142 4283 5143
rect 4279 5137 4283 5138
rect 4407 5142 4411 5143
rect 4407 5137 4411 5138
rect 4511 5142 4515 5143
rect 4511 5137 4515 5138
rect 4679 5142 4683 5143
rect 4679 5137 4683 5138
rect 4743 5142 4747 5143
rect 4743 5137 4747 5138
rect 4959 5142 4963 5143
rect 4959 5137 4963 5138
rect 4975 5142 4979 5143
rect 4975 5137 4979 5138
rect 5215 5142 5219 5143
rect 5215 5137 5219 5138
rect 5239 5142 5243 5143
rect 5239 5137 5243 5138
rect 5663 5142 5667 5143
rect 5663 5137 5667 5138
rect 3840 5114 3842 5137
rect 3838 5113 3844 5114
rect 3888 5113 3890 5137
rect 4136 5113 4138 5137
rect 4408 5113 4410 5137
rect 4680 5113 4682 5137
rect 4960 5113 4962 5137
rect 5240 5113 5242 5137
rect 5664 5114 5666 5137
rect 5662 5113 5668 5114
rect 3838 5109 3839 5113
rect 3843 5109 3844 5113
rect 3838 5108 3844 5109
rect 3886 5112 3892 5113
rect 3886 5108 3887 5112
rect 3891 5108 3892 5112
rect 3886 5107 3892 5108
rect 4134 5112 4140 5113
rect 4134 5108 4135 5112
rect 4139 5108 4140 5112
rect 4134 5107 4140 5108
rect 4406 5112 4412 5113
rect 4406 5108 4407 5112
rect 4411 5108 4412 5112
rect 4406 5107 4412 5108
rect 4678 5112 4684 5113
rect 4678 5108 4679 5112
rect 4683 5108 4684 5112
rect 4678 5107 4684 5108
rect 4958 5112 4964 5113
rect 4958 5108 4959 5112
rect 4963 5108 4964 5112
rect 4958 5107 4964 5108
rect 5238 5112 5244 5113
rect 5238 5108 5239 5112
rect 5243 5108 5244 5112
rect 5662 5109 5663 5113
rect 5667 5109 5668 5113
rect 5662 5108 5668 5109
rect 5238 5107 5244 5108
rect 3858 5097 3864 5098
rect 3838 5096 3844 5097
rect 3838 5092 3839 5096
rect 3843 5092 3844 5096
rect 3858 5093 3859 5097
rect 3863 5093 3864 5097
rect 3858 5092 3864 5093
rect 4106 5097 4112 5098
rect 4106 5093 4107 5097
rect 4111 5093 4112 5097
rect 4106 5092 4112 5093
rect 4378 5097 4384 5098
rect 4378 5093 4379 5097
rect 4383 5093 4384 5097
rect 4378 5092 4384 5093
rect 4650 5097 4656 5098
rect 4650 5093 4651 5097
rect 4655 5093 4656 5097
rect 4650 5092 4656 5093
rect 4930 5097 4936 5098
rect 4930 5093 4931 5097
rect 4935 5093 4936 5097
rect 4930 5092 4936 5093
rect 5210 5097 5216 5098
rect 5210 5093 5211 5097
rect 5215 5093 5216 5097
rect 5210 5092 5216 5093
rect 5662 5096 5668 5097
rect 5662 5092 5663 5096
rect 5667 5092 5668 5096
rect 3838 5091 3844 5092
rect 1935 5089 1939 5090
rect 1975 5090 1979 5091
rect 112 5029 114 5089
rect 110 5028 116 5029
rect 348 5028 350 5089
rect 484 5028 486 5089
rect 620 5028 622 5089
rect 756 5028 758 5089
rect 892 5028 894 5089
rect 1036 5028 1038 5089
rect 1188 5028 1190 5089
rect 1340 5028 1342 5089
rect 1492 5028 1494 5089
rect 1652 5028 1654 5089
rect 1788 5028 1790 5089
rect 1936 5029 1938 5089
rect 1975 5085 1979 5086
rect 1995 5090 1999 5091
rect 1995 5085 1999 5086
rect 2131 5090 2135 5091
rect 2131 5085 2135 5086
rect 2299 5090 2303 5091
rect 2299 5085 2303 5086
rect 2483 5090 2487 5091
rect 2483 5085 2487 5086
rect 2531 5090 2535 5091
rect 2531 5085 2535 5086
rect 2667 5090 2671 5091
rect 2667 5085 2671 5086
rect 2859 5090 2863 5091
rect 2859 5085 2863 5086
rect 3059 5090 3063 5091
rect 3059 5085 3063 5086
rect 3099 5090 3103 5091
rect 3099 5085 3103 5086
rect 3259 5090 3263 5091
rect 3259 5085 3263 5086
rect 3467 5090 3471 5091
rect 3467 5085 3471 5086
rect 3651 5090 3655 5091
rect 3651 5085 3655 5086
rect 3799 5090 3803 5091
rect 3799 5085 3803 5086
rect 1934 5028 1940 5029
rect 110 5024 111 5028
rect 115 5024 116 5028
rect 110 5023 116 5024
rect 346 5027 352 5028
rect 346 5023 347 5027
rect 351 5023 352 5027
rect 346 5022 352 5023
rect 482 5027 488 5028
rect 482 5023 483 5027
rect 487 5023 488 5027
rect 482 5022 488 5023
rect 618 5027 624 5028
rect 618 5023 619 5027
rect 623 5023 624 5027
rect 618 5022 624 5023
rect 754 5027 760 5028
rect 754 5023 755 5027
rect 759 5023 760 5027
rect 754 5022 760 5023
rect 890 5027 896 5028
rect 890 5023 891 5027
rect 895 5023 896 5027
rect 890 5022 896 5023
rect 1034 5027 1040 5028
rect 1034 5023 1035 5027
rect 1039 5023 1040 5027
rect 1034 5022 1040 5023
rect 1186 5027 1192 5028
rect 1186 5023 1187 5027
rect 1191 5023 1192 5027
rect 1186 5022 1192 5023
rect 1338 5027 1344 5028
rect 1338 5023 1339 5027
rect 1343 5023 1344 5027
rect 1338 5022 1344 5023
rect 1490 5027 1496 5028
rect 1490 5023 1491 5027
rect 1495 5023 1496 5027
rect 1490 5022 1496 5023
rect 1650 5027 1656 5028
rect 1650 5023 1651 5027
rect 1655 5023 1656 5027
rect 1650 5022 1656 5023
rect 1786 5027 1792 5028
rect 1786 5023 1787 5027
rect 1791 5023 1792 5027
rect 1934 5024 1935 5028
rect 1939 5024 1940 5028
rect 1976 5025 1978 5085
rect 1934 5023 1940 5024
rect 1974 5024 1980 5025
rect 1996 5024 1998 5085
rect 2532 5024 2534 5085
rect 3100 5024 3102 5085
rect 3652 5024 3654 5085
rect 3800 5025 3802 5085
rect 3798 5024 3804 5025
rect 1786 5022 1792 5023
rect 1974 5020 1975 5024
rect 1979 5020 1980 5024
rect 1974 5019 1980 5020
rect 1994 5023 2000 5024
rect 1994 5019 1995 5023
rect 1999 5019 2000 5023
rect 1994 5018 2000 5019
rect 2530 5023 2536 5024
rect 2530 5019 2531 5023
rect 2535 5019 2536 5023
rect 2530 5018 2536 5019
rect 3098 5023 3104 5024
rect 3098 5019 3099 5023
rect 3103 5019 3104 5023
rect 3098 5018 3104 5019
rect 3650 5023 3656 5024
rect 3650 5019 3651 5023
rect 3655 5019 3656 5023
rect 3798 5020 3799 5024
rect 3803 5020 3804 5024
rect 3798 5019 3804 5020
rect 3840 5019 3842 5091
rect 3860 5019 3862 5092
rect 4108 5019 4110 5092
rect 4380 5019 4382 5092
rect 4652 5019 4654 5092
rect 4932 5019 4934 5092
rect 5212 5019 5214 5092
rect 5662 5091 5668 5092
rect 5664 5019 5666 5091
rect 3650 5018 3656 5019
rect 3839 5018 3843 5019
rect 3839 5013 3843 5014
rect 3859 5018 3863 5019
rect 3859 5013 3863 5014
rect 4019 5018 4023 5019
rect 4019 5013 4023 5014
rect 4107 5018 4111 5019
rect 4107 5013 4111 5014
rect 4211 5018 4215 5019
rect 4211 5013 4215 5014
rect 4379 5018 4383 5019
rect 4379 5013 4383 5014
rect 4411 5018 4415 5019
rect 4411 5013 4415 5014
rect 4627 5018 4631 5019
rect 4627 5013 4631 5014
rect 4651 5018 4655 5019
rect 4651 5013 4655 5014
rect 4843 5018 4847 5019
rect 4843 5013 4847 5014
rect 4931 5018 4935 5019
rect 4931 5013 4935 5014
rect 5067 5018 5071 5019
rect 5067 5013 5071 5014
rect 5211 5018 5215 5019
rect 5211 5013 5215 5014
rect 5299 5018 5303 5019
rect 5299 5013 5303 5014
rect 5663 5018 5667 5019
rect 5663 5013 5667 5014
rect 374 5012 380 5013
rect 110 5011 116 5012
rect 110 5007 111 5011
rect 115 5007 116 5011
rect 374 5008 375 5012
rect 379 5008 380 5012
rect 374 5007 380 5008
rect 510 5012 516 5013
rect 510 5008 511 5012
rect 515 5008 516 5012
rect 510 5007 516 5008
rect 646 5012 652 5013
rect 646 5008 647 5012
rect 651 5008 652 5012
rect 646 5007 652 5008
rect 782 5012 788 5013
rect 782 5008 783 5012
rect 787 5008 788 5012
rect 782 5007 788 5008
rect 918 5012 924 5013
rect 918 5008 919 5012
rect 923 5008 924 5012
rect 918 5007 924 5008
rect 1062 5012 1068 5013
rect 1062 5008 1063 5012
rect 1067 5008 1068 5012
rect 1062 5007 1068 5008
rect 1214 5012 1220 5013
rect 1214 5008 1215 5012
rect 1219 5008 1220 5012
rect 1214 5007 1220 5008
rect 1366 5012 1372 5013
rect 1366 5008 1367 5012
rect 1371 5008 1372 5012
rect 1366 5007 1372 5008
rect 1518 5012 1524 5013
rect 1518 5008 1519 5012
rect 1523 5008 1524 5012
rect 1518 5007 1524 5008
rect 1678 5012 1684 5013
rect 1678 5008 1679 5012
rect 1683 5008 1684 5012
rect 1678 5007 1684 5008
rect 1814 5012 1820 5013
rect 1814 5008 1815 5012
rect 1819 5008 1820 5012
rect 1814 5007 1820 5008
rect 1934 5011 1940 5012
rect 1934 5007 1935 5011
rect 1939 5007 1940 5011
rect 2022 5008 2028 5009
rect 110 5006 116 5007
rect 112 4983 114 5006
rect 376 4983 378 5007
rect 512 4983 514 5007
rect 648 4983 650 5007
rect 784 4983 786 5007
rect 920 4983 922 5007
rect 1064 4983 1066 5007
rect 1216 4983 1218 5007
rect 1368 4983 1370 5007
rect 1520 4983 1522 5007
rect 1680 4983 1682 5007
rect 1816 4983 1818 5007
rect 1934 5006 1940 5007
rect 1974 5007 1980 5008
rect 1936 4983 1938 5006
rect 1974 5003 1975 5007
rect 1979 5003 1980 5007
rect 2022 5004 2023 5008
rect 2027 5004 2028 5008
rect 2022 5003 2028 5004
rect 2558 5008 2564 5009
rect 2558 5004 2559 5008
rect 2563 5004 2564 5008
rect 2558 5003 2564 5004
rect 3126 5008 3132 5009
rect 3126 5004 3127 5008
rect 3131 5004 3132 5008
rect 3126 5003 3132 5004
rect 3678 5008 3684 5009
rect 3678 5004 3679 5008
rect 3683 5004 3684 5008
rect 3678 5003 3684 5004
rect 3798 5007 3804 5008
rect 3798 5003 3799 5007
rect 3803 5003 3804 5007
rect 1974 5002 1980 5003
rect 111 4982 115 4983
rect 111 4977 115 4978
rect 159 4982 163 4983
rect 159 4977 163 4978
rect 343 4982 347 4983
rect 343 4977 347 4978
rect 375 4982 379 4983
rect 375 4977 379 4978
rect 511 4982 515 4983
rect 511 4977 515 4978
rect 551 4982 555 4983
rect 551 4977 555 4978
rect 647 4982 651 4983
rect 647 4977 651 4978
rect 751 4982 755 4983
rect 751 4977 755 4978
rect 783 4982 787 4983
rect 783 4977 787 4978
rect 919 4982 923 4983
rect 919 4977 923 4978
rect 943 4982 947 4983
rect 943 4977 947 4978
rect 1063 4982 1067 4983
rect 1063 4977 1067 4978
rect 1127 4982 1131 4983
rect 1127 4977 1131 4978
rect 1215 4982 1219 4983
rect 1215 4977 1219 4978
rect 1311 4982 1315 4983
rect 1311 4977 1315 4978
rect 1367 4982 1371 4983
rect 1367 4977 1371 4978
rect 1487 4982 1491 4983
rect 1487 4977 1491 4978
rect 1519 4982 1523 4983
rect 1519 4977 1523 4978
rect 1663 4982 1667 4983
rect 1663 4977 1667 4978
rect 1679 4982 1683 4983
rect 1679 4977 1683 4978
rect 1815 4982 1819 4983
rect 1815 4977 1819 4978
rect 1935 4982 1939 4983
rect 1935 4977 1939 4978
rect 112 4954 114 4977
rect 110 4953 116 4954
rect 160 4953 162 4977
rect 344 4953 346 4977
rect 552 4953 554 4977
rect 752 4953 754 4977
rect 944 4953 946 4977
rect 1128 4953 1130 4977
rect 1312 4953 1314 4977
rect 1488 4953 1490 4977
rect 1664 4953 1666 4977
rect 1816 4953 1818 4977
rect 1936 4954 1938 4977
rect 1934 4953 1940 4954
rect 110 4949 111 4953
rect 115 4949 116 4953
rect 110 4948 116 4949
rect 158 4952 164 4953
rect 158 4948 159 4952
rect 163 4948 164 4952
rect 158 4947 164 4948
rect 342 4952 348 4953
rect 342 4948 343 4952
rect 347 4948 348 4952
rect 342 4947 348 4948
rect 550 4952 556 4953
rect 550 4948 551 4952
rect 555 4948 556 4952
rect 550 4947 556 4948
rect 750 4952 756 4953
rect 750 4948 751 4952
rect 755 4948 756 4952
rect 750 4947 756 4948
rect 942 4952 948 4953
rect 942 4948 943 4952
rect 947 4948 948 4952
rect 942 4947 948 4948
rect 1126 4952 1132 4953
rect 1126 4948 1127 4952
rect 1131 4948 1132 4952
rect 1126 4947 1132 4948
rect 1310 4952 1316 4953
rect 1310 4948 1311 4952
rect 1315 4948 1316 4952
rect 1310 4947 1316 4948
rect 1486 4952 1492 4953
rect 1486 4948 1487 4952
rect 1491 4948 1492 4952
rect 1486 4947 1492 4948
rect 1662 4952 1668 4953
rect 1662 4948 1663 4952
rect 1667 4948 1668 4952
rect 1662 4947 1668 4948
rect 1814 4952 1820 4953
rect 1814 4948 1815 4952
rect 1819 4948 1820 4952
rect 1934 4949 1935 4953
rect 1939 4949 1940 4953
rect 1934 4948 1940 4949
rect 1814 4947 1820 4948
rect 1976 4947 1978 5002
rect 2024 4947 2026 5003
rect 2560 4947 2562 5003
rect 3128 4947 3130 5003
rect 3680 4947 3682 5003
rect 3798 5002 3804 5003
rect 3800 4947 3802 5002
rect 3840 4953 3842 5013
rect 3838 4952 3844 4953
rect 3860 4952 3862 5013
rect 4020 4952 4022 5013
rect 4212 4952 4214 5013
rect 4412 4952 4414 5013
rect 4628 4952 4630 5013
rect 4844 4952 4846 5013
rect 5068 4952 5070 5013
rect 5300 4952 5302 5013
rect 5664 4953 5666 5013
rect 5662 4952 5668 4953
rect 3838 4948 3839 4952
rect 3843 4948 3844 4952
rect 3838 4947 3844 4948
rect 3858 4951 3864 4952
rect 3858 4947 3859 4951
rect 3863 4947 3864 4951
rect 1975 4946 1979 4947
rect 1975 4941 1979 4942
rect 2023 4946 2027 4947
rect 2023 4941 2027 4942
rect 2559 4946 2563 4947
rect 2559 4941 2563 4942
rect 2871 4946 2875 4947
rect 2871 4941 2875 4942
rect 3007 4946 3011 4947
rect 3007 4941 3011 4942
rect 3127 4946 3131 4947
rect 3127 4941 3131 4942
rect 3679 4946 3683 4947
rect 3679 4941 3683 4942
rect 3799 4946 3803 4947
rect 3858 4946 3864 4947
rect 4018 4951 4024 4952
rect 4018 4947 4019 4951
rect 4023 4947 4024 4951
rect 4018 4946 4024 4947
rect 4210 4951 4216 4952
rect 4210 4947 4211 4951
rect 4215 4947 4216 4951
rect 4210 4946 4216 4947
rect 4410 4951 4416 4952
rect 4410 4947 4411 4951
rect 4415 4947 4416 4951
rect 4410 4946 4416 4947
rect 4626 4951 4632 4952
rect 4626 4947 4627 4951
rect 4631 4947 4632 4951
rect 4626 4946 4632 4947
rect 4842 4951 4848 4952
rect 4842 4947 4843 4951
rect 4847 4947 4848 4951
rect 4842 4946 4848 4947
rect 5066 4951 5072 4952
rect 5066 4947 5067 4951
rect 5071 4947 5072 4951
rect 5066 4946 5072 4947
rect 5298 4951 5304 4952
rect 5298 4947 5299 4951
rect 5303 4947 5304 4951
rect 5662 4948 5663 4952
rect 5667 4948 5668 4952
rect 5662 4947 5668 4948
rect 5298 4946 5304 4947
rect 3799 4941 3803 4942
rect 130 4937 136 4938
rect 110 4936 116 4937
rect 110 4932 111 4936
rect 115 4932 116 4936
rect 130 4933 131 4937
rect 135 4933 136 4937
rect 130 4932 136 4933
rect 314 4937 320 4938
rect 314 4933 315 4937
rect 319 4933 320 4937
rect 314 4932 320 4933
rect 522 4937 528 4938
rect 522 4933 523 4937
rect 527 4933 528 4937
rect 522 4932 528 4933
rect 722 4937 728 4938
rect 722 4933 723 4937
rect 727 4933 728 4937
rect 722 4932 728 4933
rect 914 4937 920 4938
rect 914 4933 915 4937
rect 919 4933 920 4937
rect 914 4932 920 4933
rect 1098 4937 1104 4938
rect 1098 4933 1099 4937
rect 1103 4933 1104 4937
rect 1098 4932 1104 4933
rect 1282 4937 1288 4938
rect 1282 4933 1283 4937
rect 1287 4933 1288 4937
rect 1282 4932 1288 4933
rect 1458 4937 1464 4938
rect 1458 4933 1459 4937
rect 1463 4933 1464 4937
rect 1458 4932 1464 4933
rect 1634 4937 1640 4938
rect 1634 4933 1635 4937
rect 1639 4933 1640 4937
rect 1634 4932 1640 4933
rect 1786 4937 1792 4938
rect 1786 4933 1787 4937
rect 1791 4933 1792 4937
rect 1786 4932 1792 4933
rect 1934 4936 1940 4937
rect 1934 4932 1935 4936
rect 1939 4932 1940 4936
rect 110 4931 116 4932
rect 112 4863 114 4931
rect 132 4863 134 4932
rect 316 4863 318 4932
rect 524 4863 526 4932
rect 724 4863 726 4932
rect 916 4863 918 4932
rect 1100 4863 1102 4932
rect 1284 4863 1286 4932
rect 1460 4863 1462 4932
rect 1636 4863 1638 4932
rect 1788 4863 1790 4932
rect 1934 4931 1940 4932
rect 1936 4863 1938 4931
rect 1976 4918 1978 4941
rect 1974 4917 1980 4918
rect 2872 4917 2874 4941
rect 3008 4917 3010 4941
rect 3800 4918 3802 4941
rect 3886 4936 3892 4937
rect 3838 4935 3844 4936
rect 3838 4931 3839 4935
rect 3843 4931 3844 4935
rect 3886 4932 3887 4936
rect 3891 4932 3892 4936
rect 3886 4931 3892 4932
rect 4046 4936 4052 4937
rect 4046 4932 4047 4936
rect 4051 4932 4052 4936
rect 4046 4931 4052 4932
rect 4238 4936 4244 4937
rect 4238 4932 4239 4936
rect 4243 4932 4244 4936
rect 4238 4931 4244 4932
rect 4438 4936 4444 4937
rect 4438 4932 4439 4936
rect 4443 4932 4444 4936
rect 4438 4931 4444 4932
rect 4654 4936 4660 4937
rect 4654 4932 4655 4936
rect 4659 4932 4660 4936
rect 4654 4931 4660 4932
rect 4870 4936 4876 4937
rect 4870 4932 4871 4936
rect 4875 4932 4876 4936
rect 4870 4931 4876 4932
rect 5094 4936 5100 4937
rect 5094 4932 5095 4936
rect 5099 4932 5100 4936
rect 5094 4931 5100 4932
rect 5326 4936 5332 4937
rect 5326 4932 5327 4936
rect 5331 4932 5332 4936
rect 5326 4931 5332 4932
rect 5662 4935 5668 4936
rect 5662 4931 5663 4935
rect 5667 4931 5668 4935
rect 3838 4930 3844 4931
rect 3798 4917 3804 4918
rect 1974 4913 1975 4917
rect 1979 4913 1980 4917
rect 1974 4912 1980 4913
rect 2870 4916 2876 4917
rect 2870 4912 2871 4916
rect 2875 4912 2876 4916
rect 2870 4911 2876 4912
rect 3006 4916 3012 4917
rect 3006 4912 3007 4916
rect 3011 4912 3012 4916
rect 3798 4913 3799 4917
rect 3803 4913 3804 4917
rect 3798 4912 3804 4913
rect 3006 4911 3012 4912
rect 2842 4901 2848 4902
rect 1974 4900 1980 4901
rect 1974 4896 1975 4900
rect 1979 4896 1980 4900
rect 2842 4897 2843 4901
rect 2847 4897 2848 4901
rect 2842 4896 2848 4897
rect 2978 4901 2984 4902
rect 2978 4897 2979 4901
rect 2983 4897 2984 4901
rect 2978 4896 2984 4897
rect 3798 4900 3804 4901
rect 3798 4896 3799 4900
rect 3803 4896 3804 4900
rect 1974 4895 1980 4896
rect 111 4862 115 4863
rect 111 4857 115 4858
rect 131 4862 135 4863
rect 131 4857 135 4858
rect 267 4862 271 4863
rect 267 4857 271 4858
rect 315 4862 319 4863
rect 315 4857 319 4858
rect 403 4862 407 4863
rect 403 4857 407 4858
rect 523 4862 527 4863
rect 523 4857 527 4858
rect 539 4862 543 4863
rect 539 4857 543 4858
rect 675 4862 679 4863
rect 675 4857 679 4858
rect 723 4862 727 4863
rect 723 4857 727 4858
rect 915 4862 919 4863
rect 915 4857 919 4858
rect 1099 4862 1103 4863
rect 1099 4857 1103 4858
rect 1283 4862 1287 4863
rect 1283 4857 1287 4858
rect 1459 4862 1463 4863
rect 1459 4857 1463 4858
rect 1635 4862 1639 4863
rect 1635 4857 1639 4858
rect 1787 4862 1791 4863
rect 1787 4857 1791 4858
rect 1935 4862 1939 4863
rect 1935 4857 1939 4858
rect 112 4797 114 4857
rect 110 4796 116 4797
rect 132 4796 134 4857
rect 268 4796 270 4857
rect 404 4796 406 4857
rect 540 4796 542 4857
rect 676 4796 678 4857
rect 1936 4797 1938 4857
rect 1976 4811 1978 4895
rect 2844 4811 2846 4896
rect 2980 4811 2982 4896
rect 3798 4895 3804 4896
rect 3800 4811 3802 4895
rect 3840 4887 3842 4930
rect 3888 4887 3890 4931
rect 4048 4887 4050 4931
rect 4240 4887 4242 4931
rect 4440 4887 4442 4931
rect 4656 4887 4658 4931
rect 4872 4887 4874 4931
rect 5096 4887 5098 4931
rect 5328 4887 5330 4931
rect 5662 4930 5668 4931
rect 5664 4887 5666 4930
rect 3839 4886 3843 4887
rect 3839 4881 3843 4882
rect 3887 4886 3891 4887
rect 3887 4881 3891 4882
rect 4047 4886 4051 4887
rect 4047 4881 4051 4882
rect 4071 4886 4075 4887
rect 4071 4881 4075 4882
rect 4239 4886 4243 4887
rect 4239 4881 4243 4882
rect 4287 4886 4291 4887
rect 4287 4881 4291 4882
rect 4439 4886 4443 4887
rect 4439 4881 4443 4882
rect 4511 4886 4515 4887
rect 4511 4881 4515 4882
rect 4655 4886 4659 4887
rect 4655 4881 4659 4882
rect 4735 4886 4739 4887
rect 4735 4881 4739 4882
rect 4871 4886 4875 4887
rect 4871 4881 4875 4882
rect 4959 4886 4963 4887
rect 4959 4881 4963 4882
rect 5095 4886 5099 4887
rect 5095 4881 5099 4882
rect 5183 4886 5187 4887
rect 5183 4881 5187 4882
rect 5327 4886 5331 4887
rect 5327 4881 5331 4882
rect 5407 4886 5411 4887
rect 5407 4881 5411 4882
rect 5663 4886 5667 4887
rect 5663 4881 5667 4882
rect 3840 4858 3842 4881
rect 3838 4857 3844 4858
rect 3888 4857 3890 4881
rect 4072 4857 4074 4881
rect 4288 4857 4290 4881
rect 4512 4857 4514 4881
rect 4736 4857 4738 4881
rect 4960 4857 4962 4881
rect 5184 4857 5186 4881
rect 5408 4857 5410 4881
rect 5664 4858 5666 4881
rect 5662 4857 5668 4858
rect 3838 4853 3839 4857
rect 3843 4853 3844 4857
rect 3838 4852 3844 4853
rect 3886 4856 3892 4857
rect 3886 4852 3887 4856
rect 3891 4852 3892 4856
rect 3886 4851 3892 4852
rect 4070 4856 4076 4857
rect 4070 4852 4071 4856
rect 4075 4852 4076 4856
rect 4070 4851 4076 4852
rect 4286 4856 4292 4857
rect 4286 4852 4287 4856
rect 4291 4852 4292 4856
rect 4286 4851 4292 4852
rect 4510 4856 4516 4857
rect 4510 4852 4511 4856
rect 4515 4852 4516 4856
rect 4510 4851 4516 4852
rect 4734 4856 4740 4857
rect 4734 4852 4735 4856
rect 4739 4852 4740 4856
rect 4734 4851 4740 4852
rect 4958 4856 4964 4857
rect 4958 4852 4959 4856
rect 4963 4852 4964 4856
rect 4958 4851 4964 4852
rect 5182 4856 5188 4857
rect 5182 4852 5183 4856
rect 5187 4852 5188 4856
rect 5182 4851 5188 4852
rect 5406 4856 5412 4857
rect 5406 4852 5407 4856
rect 5411 4852 5412 4856
rect 5662 4853 5663 4857
rect 5667 4853 5668 4857
rect 5662 4852 5668 4853
rect 5406 4851 5412 4852
rect 3858 4841 3864 4842
rect 3838 4840 3844 4841
rect 3838 4836 3839 4840
rect 3843 4836 3844 4840
rect 3858 4837 3859 4841
rect 3863 4837 3864 4841
rect 3858 4836 3864 4837
rect 4042 4841 4048 4842
rect 4042 4837 4043 4841
rect 4047 4837 4048 4841
rect 4042 4836 4048 4837
rect 4258 4841 4264 4842
rect 4258 4837 4259 4841
rect 4263 4837 4264 4841
rect 4258 4836 4264 4837
rect 4482 4841 4488 4842
rect 4482 4837 4483 4841
rect 4487 4837 4488 4841
rect 4482 4836 4488 4837
rect 4706 4841 4712 4842
rect 4706 4837 4707 4841
rect 4711 4837 4712 4841
rect 4706 4836 4712 4837
rect 4930 4841 4936 4842
rect 4930 4837 4931 4841
rect 4935 4837 4936 4841
rect 4930 4836 4936 4837
rect 5154 4841 5160 4842
rect 5154 4837 5155 4841
rect 5159 4837 5160 4841
rect 5154 4836 5160 4837
rect 5378 4841 5384 4842
rect 5378 4837 5379 4841
rect 5383 4837 5384 4841
rect 5378 4836 5384 4837
rect 5662 4840 5668 4841
rect 5662 4836 5663 4840
rect 5667 4836 5668 4840
rect 3838 4835 3844 4836
rect 1975 4810 1979 4811
rect 1975 4805 1979 4806
rect 1995 4810 1999 4811
rect 1995 4805 1999 4806
rect 2155 4810 2159 4811
rect 2155 4805 2159 4806
rect 2347 4810 2351 4811
rect 2347 4805 2351 4806
rect 2539 4810 2543 4811
rect 2539 4805 2543 4806
rect 2731 4810 2735 4811
rect 2731 4805 2735 4806
rect 2843 4810 2847 4811
rect 2843 4805 2847 4806
rect 2931 4810 2935 4811
rect 2931 4805 2935 4806
rect 2979 4810 2983 4811
rect 2979 4805 2983 4806
rect 3131 4810 3135 4811
rect 3131 4805 3135 4806
rect 3799 4810 3803 4811
rect 3799 4805 3803 4806
rect 1934 4796 1940 4797
rect 110 4792 111 4796
rect 115 4792 116 4796
rect 110 4791 116 4792
rect 130 4795 136 4796
rect 130 4791 131 4795
rect 135 4791 136 4795
rect 130 4790 136 4791
rect 266 4795 272 4796
rect 266 4791 267 4795
rect 271 4791 272 4795
rect 266 4790 272 4791
rect 402 4795 408 4796
rect 402 4791 403 4795
rect 407 4791 408 4795
rect 402 4790 408 4791
rect 538 4795 544 4796
rect 538 4791 539 4795
rect 543 4791 544 4795
rect 538 4790 544 4791
rect 674 4795 680 4796
rect 674 4791 675 4795
rect 679 4791 680 4795
rect 1934 4792 1935 4796
rect 1939 4792 1940 4796
rect 1934 4791 1940 4792
rect 674 4790 680 4791
rect 158 4780 164 4781
rect 110 4779 116 4780
rect 110 4775 111 4779
rect 115 4775 116 4779
rect 158 4776 159 4780
rect 163 4776 164 4780
rect 158 4775 164 4776
rect 294 4780 300 4781
rect 294 4776 295 4780
rect 299 4776 300 4780
rect 294 4775 300 4776
rect 430 4780 436 4781
rect 430 4776 431 4780
rect 435 4776 436 4780
rect 430 4775 436 4776
rect 566 4780 572 4781
rect 566 4776 567 4780
rect 571 4776 572 4780
rect 566 4775 572 4776
rect 702 4780 708 4781
rect 702 4776 703 4780
rect 707 4776 708 4780
rect 702 4775 708 4776
rect 1934 4779 1940 4780
rect 1934 4775 1935 4779
rect 1939 4775 1940 4779
rect 110 4774 116 4775
rect 112 4743 114 4774
rect 160 4743 162 4775
rect 296 4743 298 4775
rect 432 4743 434 4775
rect 568 4743 570 4775
rect 704 4743 706 4775
rect 1934 4774 1940 4775
rect 1936 4743 1938 4774
rect 1976 4745 1978 4805
rect 1974 4744 1980 4745
rect 1996 4744 1998 4805
rect 2156 4744 2158 4805
rect 2348 4744 2350 4805
rect 2540 4744 2542 4805
rect 2732 4744 2734 4805
rect 2932 4744 2934 4805
rect 3132 4744 3134 4805
rect 3800 4745 3802 4805
rect 3840 4771 3842 4835
rect 3860 4771 3862 4836
rect 4044 4771 4046 4836
rect 4260 4771 4262 4836
rect 4484 4771 4486 4836
rect 4708 4771 4710 4836
rect 4932 4771 4934 4836
rect 5156 4771 5158 4836
rect 5380 4771 5382 4836
rect 5662 4835 5668 4836
rect 5664 4771 5666 4835
rect 3839 4770 3843 4771
rect 3839 4765 3843 4766
rect 3859 4770 3863 4771
rect 3859 4765 3863 4766
rect 3915 4770 3919 4771
rect 3915 4765 3919 4766
rect 4043 4770 4047 4771
rect 4043 4765 4047 4766
rect 4187 4770 4191 4771
rect 4187 4765 4191 4766
rect 4259 4770 4263 4771
rect 4259 4765 4263 4766
rect 4467 4770 4471 4771
rect 4467 4765 4471 4766
rect 4483 4770 4487 4771
rect 4483 4765 4487 4766
rect 4707 4770 4711 4771
rect 4707 4765 4711 4766
rect 4763 4770 4767 4771
rect 4763 4765 4767 4766
rect 4931 4770 4935 4771
rect 4931 4765 4935 4766
rect 5067 4770 5071 4771
rect 5067 4765 5071 4766
rect 5155 4770 5159 4771
rect 5155 4765 5159 4766
rect 5371 4770 5375 4771
rect 5371 4765 5375 4766
rect 5379 4770 5383 4771
rect 5379 4765 5383 4766
rect 5663 4770 5667 4771
rect 5663 4765 5667 4766
rect 3798 4744 3804 4745
rect 111 4742 115 4743
rect 111 4737 115 4738
rect 159 4742 163 4743
rect 159 4737 163 4738
rect 295 4742 299 4743
rect 295 4737 299 4738
rect 343 4742 347 4743
rect 343 4737 347 4738
rect 431 4742 435 4743
rect 431 4737 435 4738
rect 567 4742 571 4743
rect 567 4737 571 4738
rect 703 4742 707 4743
rect 703 4737 707 4738
rect 807 4742 811 4743
rect 807 4737 811 4738
rect 1055 4742 1059 4743
rect 1055 4737 1059 4738
rect 1311 4742 1315 4743
rect 1311 4737 1315 4738
rect 1575 4742 1579 4743
rect 1575 4737 1579 4738
rect 1815 4742 1819 4743
rect 1815 4737 1819 4738
rect 1935 4742 1939 4743
rect 1974 4740 1975 4744
rect 1979 4740 1980 4744
rect 1974 4739 1980 4740
rect 1994 4743 2000 4744
rect 1994 4739 1995 4743
rect 1999 4739 2000 4743
rect 1994 4738 2000 4739
rect 2154 4743 2160 4744
rect 2154 4739 2155 4743
rect 2159 4739 2160 4743
rect 2154 4738 2160 4739
rect 2346 4743 2352 4744
rect 2346 4739 2347 4743
rect 2351 4739 2352 4743
rect 2346 4738 2352 4739
rect 2538 4743 2544 4744
rect 2538 4739 2539 4743
rect 2543 4739 2544 4743
rect 2538 4738 2544 4739
rect 2730 4743 2736 4744
rect 2730 4739 2731 4743
rect 2735 4739 2736 4743
rect 2730 4738 2736 4739
rect 2930 4743 2936 4744
rect 2930 4739 2931 4743
rect 2935 4739 2936 4743
rect 2930 4738 2936 4739
rect 3130 4743 3136 4744
rect 3130 4739 3131 4743
rect 3135 4739 3136 4743
rect 3798 4740 3799 4744
rect 3803 4740 3804 4744
rect 3798 4739 3804 4740
rect 3130 4738 3136 4739
rect 1935 4737 1939 4738
rect 112 4714 114 4737
rect 110 4713 116 4714
rect 160 4713 162 4737
rect 344 4713 346 4737
rect 568 4713 570 4737
rect 808 4713 810 4737
rect 1056 4713 1058 4737
rect 1312 4713 1314 4737
rect 1576 4713 1578 4737
rect 1816 4713 1818 4737
rect 1936 4714 1938 4737
rect 2022 4728 2028 4729
rect 1974 4727 1980 4728
rect 1974 4723 1975 4727
rect 1979 4723 1980 4727
rect 2022 4724 2023 4728
rect 2027 4724 2028 4728
rect 2022 4723 2028 4724
rect 2182 4728 2188 4729
rect 2182 4724 2183 4728
rect 2187 4724 2188 4728
rect 2182 4723 2188 4724
rect 2374 4728 2380 4729
rect 2374 4724 2375 4728
rect 2379 4724 2380 4728
rect 2374 4723 2380 4724
rect 2566 4728 2572 4729
rect 2566 4724 2567 4728
rect 2571 4724 2572 4728
rect 2566 4723 2572 4724
rect 2758 4728 2764 4729
rect 2758 4724 2759 4728
rect 2763 4724 2764 4728
rect 2758 4723 2764 4724
rect 2958 4728 2964 4729
rect 2958 4724 2959 4728
rect 2963 4724 2964 4728
rect 2958 4723 2964 4724
rect 3158 4728 3164 4729
rect 3158 4724 3159 4728
rect 3163 4724 3164 4728
rect 3158 4723 3164 4724
rect 3798 4727 3804 4728
rect 3798 4723 3799 4727
rect 3803 4723 3804 4727
rect 1974 4722 1980 4723
rect 1934 4713 1940 4714
rect 110 4709 111 4713
rect 115 4709 116 4713
rect 110 4708 116 4709
rect 158 4712 164 4713
rect 158 4708 159 4712
rect 163 4708 164 4712
rect 158 4707 164 4708
rect 342 4712 348 4713
rect 342 4708 343 4712
rect 347 4708 348 4712
rect 342 4707 348 4708
rect 566 4712 572 4713
rect 566 4708 567 4712
rect 571 4708 572 4712
rect 566 4707 572 4708
rect 806 4712 812 4713
rect 806 4708 807 4712
rect 811 4708 812 4712
rect 806 4707 812 4708
rect 1054 4712 1060 4713
rect 1054 4708 1055 4712
rect 1059 4708 1060 4712
rect 1054 4707 1060 4708
rect 1310 4712 1316 4713
rect 1310 4708 1311 4712
rect 1315 4708 1316 4712
rect 1310 4707 1316 4708
rect 1574 4712 1580 4713
rect 1574 4708 1575 4712
rect 1579 4708 1580 4712
rect 1574 4707 1580 4708
rect 1814 4712 1820 4713
rect 1814 4708 1815 4712
rect 1819 4708 1820 4712
rect 1934 4709 1935 4713
rect 1939 4709 1940 4713
rect 1934 4708 1940 4709
rect 1814 4707 1820 4708
rect 130 4697 136 4698
rect 110 4696 116 4697
rect 110 4692 111 4696
rect 115 4692 116 4696
rect 130 4693 131 4697
rect 135 4693 136 4697
rect 130 4692 136 4693
rect 314 4697 320 4698
rect 314 4693 315 4697
rect 319 4693 320 4697
rect 314 4692 320 4693
rect 538 4697 544 4698
rect 538 4693 539 4697
rect 543 4693 544 4697
rect 538 4692 544 4693
rect 778 4697 784 4698
rect 778 4693 779 4697
rect 783 4693 784 4697
rect 778 4692 784 4693
rect 1026 4697 1032 4698
rect 1026 4693 1027 4697
rect 1031 4693 1032 4697
rect 1026 4692 1032 4693
rect 1282 4697 1288 4698
rect 1282 4693 1283 4697
rect 1287 4693 1288 4697
rect 1282 4692 1288 4693
rect 1546 4697 1552 4698
rect 1546 4693 1547 4697
rect 1551 4693 1552 4697
rect 1546 4692 1552 4693
rect 1786 4697 1792 4698
rect 1786 4693 1787 4697
rect 1791 4693 1792 4697
rect 1786 4692 1792 4693
rect 1934 4696 1940 4697
rect 1934 4692 1935 4696
rect 1939 4692 1940 4696
rect 1976 4695 1978 4722
rect 2024 4695 2026 4723
rect 2184 4695 2186 4723
rect 2376 4695 2378 4723
rect 2568 4695 2570 4723
rect 2760 4695 2762 4723
rect 2960 4695 2962 4723
rect 3160 4695 3162 4723
rect 3798 4722 3804 4723
rect 3800 4695 3802 4722
rect 3840 4705 3842 4765
rect 3838 4704 3844 4705
rect 3916 4704 3918 4765
rect 4188 4704 4190 4765
rect 4468 4704 4470 4765
rect 4764 4704 4766 4765
rect 5068 4704 5070 4765
rect 5372 4704 5374 4765
rect 5664 4705 5666 4765
rect 5662 4704 5668 4705
rect 3838 4700 3839 4704
rect 3843 4700 3844 4704
rect 3838 4699 3844 4700
rect 3914 4703 3920 4704
rect 3914 4699 3915 4703
rect 3919 4699 3920 4703
rect 3914 4698 3920 4699
rect 4186 4703 4192 4704
rect 4186 4699 4187 4703
rect 4191 4699 4192 4703
rect 4186 4698 4192 4699
rect 4466 4703 4472 4704
rect 4466 4699 4467 4703
rect 4471 4699 4472 4703
rect 4466 4698 4472 4699
rect 4762 4703 4768 4704
rect 4762 4699 4763 4703
rect 4767 4699 4768 4703
rect 4762 4698 4768 4699
rect 5066 4703 5072 4704
rect 5066 4699 5067 4703
rect 5071 4699 5072 4703
rect 5066 4698 5072 4699
rect 5370 4703 5376 4704
rect 5370 4699 5371 4703
rect 5375 4699 5376 4703
rect 5662 4700 5663 4704
rect 5667 4700 5668 4704
rect 5662 4699 5668 4700
rect 5370 4698 5376 4699
rect 110 4691 116 4692
rect 112 4615 114 4691
rect 132 4615 134 4692
rect 316 4615 318 4692
rect 540 4615 542 4692
rect 780 4615 782 4692
rect 1028 4615 1030 4692
rect 1284 4615 1286 4692
rect 1548 4615 1550 4692
rect 1788 4615 1790 4692
rect 1934 4691 1940 4692
rect 1975 4694 1979 4695
rect 1936 4615 1938 4691
rect 1975 4689 1979 4690
rect 2023 4694 2027 4695
rect 2023 4689 2027 4690
rect 2183 4694 2187 4695
rect 2183 4689 2187 4690
rect 2239 4694 2243 4695
rect 2239 4689 2243 4690
rect 2375 4694 2379 4695
rect 2375 4689 2379 4690
rect 2471 4694 2475 4695
rect 2471 4689 2475 4690
rect 2567 4694 2571 4695
rect 2567 4689 2571 4690
rect 2695 4694 2699 4695
rect 2695 4689 2699 4690
rect 2759 4694 2763 4695
rect 2759 4689 2763 4690
rect 2919 4694 2923 4695
rect 2919 4689 2923 4690
rect 2959 4694 2963 4695
rect 2959 4689 2963 4690
rect 3143 4694 3147 4695
rect 3143 4689 3147 4690
rect 3159 4694 3163 4695
rect 3159 4689 3163 4690
rect 3367 4694 3371 4695
rect 3367 4689 3371 4690
rect 3799 4694 3803 4695
rect 3799 4689 3803 4690
rect 1976 4666 1978 4689
rect 1974 4665 1980 4666
rect 2024 4665 2026 4689
rect 2240 4665 2242 4689
rect 2472 4665 2474 4689
rect 2696 4665 2698 4689
rect 2920 4665 2922 4689
rect 3144 4665 3146 4689
rect 3368 4665 3370 4689
rect 3800 4666 3802 4689
rect 3942 4688 3948 4689
rect 3838 4687 3844 4688
rect 3838 4683 3839 4687
rect 3843 4683 3844 4687
rect 3942 4684 3943 4688
rect 3947 4684 3948 4688
rect 3942 4683 3948 4684
rect 4214 4688 4220 4689
rect 4214 4684 4215 4688
rect 4219 4684 4220 4688
rect 4214 4683 4220 4684
rect 4494 4688 4500 4689
rect 4494 4684 4495 4688
rect 4499 4684 4500 4688
rect 4494 4683 4500 4684
rect 4790 4688 4796 4689
rect 4790 4684 4791 4688
rect 4795 4684 4796 4688
rect 4790 4683 4796 4684
rect 5094 4688 5100 4689
rect 5094 4684 5095 4688
rect 5099 4684 5100 4688
rect 5094 4683 5100 4684
rect 5398 4688 5404 4689
rect 5398 4684 5399 4688
rect 5403 4684 5404 4688
rect 5398 4683 5404 4684
rect 5662 4687 5668 4688
rect 5662 4683 5663 4687
rect 5667 4683 5668 4687
rect 3838 4682 3844 4683
rect 3798 4665 3804 4666
rect 1974 4661 1975 4665
rect 1979 4661 1980 4665
rect 1974 4660 1980 4661
rect 2022 4664 2028 4665
rect 2022 4660 2023 4664
rect 2027 4660 2028 4664
rect 2022 4659 2028 4660
rect 2238 4664 2244 4665
rect 2238 4660 2239 4664
rect 2243 4660 2244 4664
rect 2238 4659 2244 4660
rect 2470 4664 2476 4665
rect 2470 4660 2471 4664
rect 2475 4660 2476 4664
rect 2470 4659 2476 4660
rect 2694 4664 2700 4665
rect 2694 4660 2695 4664
rect 2699 4660 2700 4664
rect 2694 4659 2700 4660
rect 2918 4664 2924 4665
rect 2918 4660 2919 4664
rect 2923 4660 2924 4664
rect 2918 4659 2924 4660
rect 3142 4664 3148 4665
rect 3142 4660 3143 4664
rect 3147 4660 3148 4664
rect 3142 4659 3148 4660
rect 3366 4664 3372 4665
rect 3366 4660 3367 4664
rect 3371 4660 3372 4664
rect 3798 4661 3799 4665
rect 3803 4661 3804 4665
rect 3798 4660 3804 4661
rect 3366 4659 3372 4660
rect 3840 4659 3842 4682
rect 3944 4659 3946 4683
rect 4216 4659 4218 4683
rect 4496 4659 4498 4683
rect 4792 4659 4794 4683
rect 5096 4659 5098 4683
rect 5400 4659 5402 4683
rect 5662 4682 5668 4683
rect 5664 4659 5666 4682
rect 3839 4658 3843 4659
rect 3839 4653 3843 4654
rect 3943 4658 3947 4659
rect 3943 4653 3947 4654
rect 4063 4658 4067 4659
rect 4063 4653 4067 4654
rect 4215 4658 4219 4659
rect 4215 4653 4219 4654
rect 4327 4658 4331 4659
rect 4327 4653 4331 4654
rect 4495 4658 4499 4659
rect 4495 4653 4499 4654
rect 4599 4658 4603 4659
rect 4599 4653 4603 4654
rect 4791 4658 4795 4659
rect 4791 4653 4795 4654
rect 4871 4658 4875 4659
rect 4871 4653 4875 4654
rect 5095 4658 5099 4659
rect 5095 4653 5099 4654
rect 5151 4658 5155 4659
rect 5151 4653 5155 4654
rect 5399 4658 5403 4659
rect 5399 4653 5403 4654
rect 5439 4658 5443 4659
rect 5439 4653 5443 4654
rect 5663 4658 5667 4659
rect 5663 4653 5667 4654
rect 1994 4649 2000 4650
rect 1974 4648 1980 4649
rect 1974 4644 1975 4648
rect 1979 4644 1980 4648
rect 1994 4645 1995 4649
rect 1999 4645 2000 4649
rect 1994 4644 2000 4645
rect 2210 4649 2216 4650
rect 2210 4645 2211 4649
rect 2215 4645 2216 4649
rect 2210 4644 2216 4645
rect 2442 4649 2448 4650
rect 2442 4645 2443 4649
rect 2447 4645 2448 4649
rect 2442 4644 2448 4645
rect 2666 4649 2672 4650
rect 2666 4645 2667 4649
rect 2671 4645 2672 4649
rect 2666 4644 2672 4645
rect 2890 4649 2896 4650
rect 2890 4645 2891 4649
rect 2895 4645 2896 4649
rect 2890 4644 2896 4645
rect 3114 4649 3120 4650
rect 3114 4645 3115 4649
rect 3119 4645 3120 4649
rect 3114 4644 3120 4645
rect 3338 4649 3344 4650
rect 3338 4645 3339 4649
rect 3343 4645 3344 4649
rect 3338 4644 3344 4645
rect 3798 4648 3804 4649
rect 3798 4644 3799 4648
rect 3803 4644 3804 4648
rect 1974 4643 1980 4644
rect 111 4614 115 4615
rect 111 4609 115 4610
rect 131 4614 135 4615
rect 131 4609 135 4610
rect 171 4614 175 4615
rect 171 4609 175 4610
rect 315 4614 319 4615
rect 315 4609 319 4610
rect 395 4614 399 4615
rect 395 4609 399 4610
rect 539 4614 543 4615
rect 539 4609 543 4610
rect 643 4614 647 4615
rect 643 4609 647 4610
rect 779 4614 783 4615
rect 779 4609 783 4610
rect 907 4614 911 4615
rect 907 4609 911 4610
rect 1027 4614 1031 4615
rect 1027 4609 1031 4610
rect 1195 4614 1199 4615
rect 1195 4609 1199 4610
rect 1283 4614 1287 4615
rect 1283 4609 1287 4610
rect 1491 4614 1495 4615
rect 1491 4609 1495 4610
rect 1547 4614 1551 4615
rect 1547 4609 1551 4610
rect 1787 4614 1791 4615
rect 1787 4609 1791 4610
rect 1935 4614 1939 4615
rect 1935 4609 1939 4610
rect 112 4549 114 4609
rect 110 4548 116 4549
rect 172 4548 174 4609
rect 396 4548 398 4609
rect 644 4548 646 4609
rect 908 4548 910 4609
rect 1196 4548 1198 4609
rect 1492 4548 1494 4609
rect 1788 4548 1790 4609
rect 1936 4549 1938 4609
rect 1976 4579 1978 4643
rect 1996 4579 1998 4644
rect 2212 4579 2214 4644
rect 2444 4579 2446 4644
rect 2668 4579 2670 4644
rect 2892 4579 2894 4644
rect 3116 4579 3118 4644
rect 3340 4579 3342 4644
rect 3798 4643 3804 4644
rect 3800 4579 3802 4643
rect 3840 4630 3842 4653
rect 3838 4629 3844 4630
rect 4064 4629 4066 4653
rect 4328 4629 4330 4653
rect 4600 4629 4602 4653
rect 4872 4629 4874 4653
rect 5152 4629 5154 4653
rect 5440 4629 5442 4653
rect 5664 4630 5666 4653
rect 5662 4629 5668 4630
rect 3838 4625 3839 4629
rect 3843 4625 3844 4629
rect 3838 4624 3844 4625
rect 4062 4628 4068 4629
rect 4062 4624 4063 4628
rect 4067 4624 4068 4628
rect 4062 4623 4068 4624
rect 4326 4628 4332 4629
rect 4326 4624 4327 4628
rect 4331 4624 4332 4628
rect 4326 4623 4332 4624
rect 4598 4628 4604 4629
rect 4598 4624 4599 4628
rect 4603 4624 4604 4628
rect 4598 4623 4604 4624
rect 4870 4628 4876 4629
rect 4870 4624 4871 4628
rect 4875 4624 4876 4628
rect 4870 4623 4876 4624
rect 5150 4628 5156 4629
rect 5150 4624 5151 4628
rect 5155 4624 5156 4628
rect 5150 4623 5156 4624
rect 5438 4628 5444 4629
rect 5438 4624 5439 4628
rect 5443 4624 5444 4628
rect 5662 4625 5663 4629
rect 5667 4625 5668 4629
rect 5662 4624 5668 4625
rect 5438 4623 5444 4624
rect 4034 4613 4040 4614
rect 3838 4612 3844 4613
rect 3838 4608 3839 4612
rect 3843 4608 3844 4612
rect 4034 4609 4035 4613
rect 4039 4609 4040 4613
rect 4034 4608 4040 4609
rect 4298 4613 4304 4614
rect 4298 4609 4299 4613
rect 4303 4609 4304 4613
rect 4298 4608 4304 4609
rect 4570 4613 4576 4614
rect 4570 4609 4571 4613
rect 4575 4609 4576 4613
rect 4570 4608 4576 4609
rect 4842 4613 4848 4614
rect 4842 4609 4843 4613
rect 4847 4609 4848 4613
rect 4842 4608 4848 4609
rect 5122 4613 5128 4614
rect 5122 4609 5123 4613
rect 5127 4609 5128 4613
rect 5122 4608 5128 4609
rect 5410 4613 5416 4614
rect 5410 4609 5411 4613
rect 5415 4609 5416 4613
rect 5410 4608 5416 4609
rect 5662 4612 5668 4613
rect 5662 4608 5663 4612
rect 5667 4608 5668 4612
rect 3838 4607 3844 4608
rect 1975 4578 1979 4579
rect 1975 4573 1979 4574
rect 1995 4578 1999 4579
rect 1995 4573 1999 4574
rect 2099 4578 2103 4579
rect 2099 4573 2103 4574
rect 2211 4578 2215 4579
rect 2211 4573 2215 4574
rect 2347 4578 2351 4579
rect 2347 4573 2351 4574
rect 2443 4578 2447 4579
rect 2443 4573 2447 4574
rect 2579 4578 2583 4579
rect 2579 4573 2583 4574
rect 2667 4578 2671 4579
rect 2667 4573 2671 4574
rect 2795 4578 2799 4579
rect 2795 4573 2799 4574
rect 2891 4578 2895 4579
rect 2891 4573 2895 4574
rect 3003 4578 3007 4579
rect 3003 4573 3007 4574
rect 3115 4578 3119 4579
rect 3115 4573 3119 4574
rect 3203 4578 3207 4579
rect 3203 4573 3207 4574
rect 3339 4578 3343 4579
rect 3339 4573 3343 4574
rect 3403 4578 3407 4579
rect 3403 4573 3407 4574
rect 3611 4578 3615 4579
rect 3611 4573 3615 4574
rect 3799 4578 3803 4579
rect 3799 4573 3803 4574
rect 1934 4548 1940 4549
rect 110 4544 111 4548
rect 115 4544 116 4548
rect 110 4543 116 4544
rect 170 4547 176 4548
rect 170 4543 171 4547
rect 175 4543 176 4547
rect 170 4542 176 4543
rect 394 4547 400 4548
rect 394 4543 395 4547
rect 399 4543 400 4547
rect 394 4542 400 4543
rect 642 4547 648 4548
rect 642 4543 643 4547
rect 647 4543 648 4547
rect 642 4542 648 4543
rect 906 4547 912 4548
rect 906 4543 907 4547
rect 911 4543 912 4547
rect 906 4542 912 4543
rect 1194 4547 1200 4548
rect 1194 4543 1195 4547
rect 1199 4543 1200 4547
rect 1194 4542 1200 4543
rect 1490 4547 1496 4548
rect 1490 4543 1491 4547
rect 1495 4543 1496 4547
rect 1490 4542 1496 4543
rect 1786 4547 1792 4548
rect 1786 4543 1787 4547
rect 1791 4543 1792 4547
rect 1934 4544 1935 4548
rect 1939 4544 1940 4548
rect 1934 4543 1940 4544
rect 1786 4542 1792 4543
rect 198 4532 204 4533
rect 110 4531 116 4532
rect 110 4527 111 4531
rect 115 4527 116 4531
rect 198 4528 199 4532
rect 203 4528 204 4532
rect 198 4527 204 4528
rect 422 4532 428 4533
rect 422 4528 423 4532
rect 427 4528 428 4532
rect 422 4527 428 4528
rect 670 4532 676 4533
rect 670 4528 671 4532
rect 675 4528 676 4532
rect 670 4527 676 4528
rect 934 4532 940 4533
rect 934 4528 935 4532
rect 939 4528 940 4532
rect 934 4527 940 4528
rect 1222 4532 1228 4533
rect 1222 4528 1223 4532
rect 1227 4528 1228 4532
rect 1222 4527 1228 4528
rect 1518 4532 1524 4533
rect 1518 4528 1519 4532
rect 1523 4528 1524 4532
rect 1518 4527 1524 4528
rect 1814 4532 1820 4533
rect 1814 4528 1815 4532
rect 1819 4528 1820 4532
rect 1814 4527 1820 4528
rect 1934 4531 1940 4532
rect 1934 4527 1935 4531
rect 1939 4527 1940 4531
rect 110 4526 116 4527
rect 112 4499 114 4526
rect 200 4499 202 4527
rect 424 4499 426 4527
rect 672 4499 674 4527
rect 936 4499 938 4527
rect 1224 4499 1226 4527
rect 1520 4499 1522 4527
rect 1816 4499 1818 4527
rect 1934 4526 1940 4527
rect 1936 4499 1938 4526
rect 1976 4513 1978 4573
rect 1974 4512 1980 4513
rect 2100 4512 2102 4573
rect 2348 4512 2350 4573
rect 2580 4512 2582 4573
rect 2796 4512 2798 4573
rect 3004 4512 3006 4573
rect 3204 4512 3206 4573
rect 3404 4512 3406 4573
rect 3612 4512 3614 4573
rect 3800 4513 3802 4573
rect 3840 4547 3842 4607
rect 4036 4547 4038 4608
rect 4300 4547 4302 4608
rect 4572 4547 4574 4608
rect 4844 4547 4846 4608
rect 5124 4547 5126 4608
rect 5412 4547 5414 4608
rect 5662 4607 5668 4608
rect 5664 4547 5666 4607
rect 3839 4546 3843 4547
rect 3839 4541 3843 4542
rect 4035 4546 4039 4547
rect 4035 4541 4039 4542
rect 4179 4546 4183 4547
rect 4179 4541 4183 4542
rect 4299 4546 4303 4547
rect 4299 4541 4303 4542
rect 4411 4546 4415 4547
rect 4411 4541 4415 4542
rect 4571 4546 4575 4547
rect 4571 4541 4575 4542
rect 4659 4546 4663 4547
rect 4659 4541 4663 4542
rect 4843 4546 4847 4547
rect 4843 4541 4847 4542
rect 4915 4546 4919 4547
rect 4915 4541 4919 4542
rect 5123 4546 5127 4547
rect 5123 4541 5127 4542
rect 5179 4546 5183 4547
rect 5179 4541 5183 4542
rect 5411 4546 5415 4547
rect 5411 4541 5415 4542
rect 5443 4546 5447 4547
rect 5443 4541 5447 4542
rect 5663 4546 5667 4547
rect 5663 4541 5667 4542
rect 3798 4512 3804 4513
rect 1974 4508 1975 4512
rect 1979 4508 1980 4512
rect 1974 4507 1980 4508
rect 2098 4511 2104 4512
rect 2098 4507 2099 4511
rect 2103 4507 2104 4511
rect 2098 4506 2104 4507
rect 2346 4511 2352 4512
rect 2346 4507 2347 4511
rect 2351 4507 2352 4511
rect 2346 4506 2352 4507
rect 2578 4511 2584 4512
rect 2578 4507 2579 4511
rect 2583 4507 2584 4511
rect 2578 4506 2584 4507
rect 2794 4511 2800 4512
rect 2794 4507 2795 4511
rect 2799 4507 2800 4511
rect 2794 4506 2800 4507
rect 3002 4511 3008 4512
rect 3002 4507 3003 4511
rect 3007 4507 3008 4511
rect 3002 4506 3008 4507
rect 3202 4511 3208 4512
rect 3202 4507 3203 4511
rect 3207 4507 3208 4511
rect 3202 4506 3208 4507
rect 3402 4511 3408 4512
rect 3402 4507 3403 4511
rect 3407 4507 3408 4511
rect 3402 4506 3408 4507
rect 3610 4511 3616 4512
rect 3610 4507 3611 4511
rect 3615 4507 3616 4511
rect 3798 4508 3799 4512
rect 3803 4508 3804 4512
rect 3798 4507 3804 4508
rect 3610 4506 3616 4507
rect 111 4498 115 4499
rect 111 4493 115 4494
rect 199 4498 203 4499
rect 199 4493 203 4494
rect 423 4498 427 4499
rect 423 4493 427 4494
rect 447 4498 451 4499
rect 447 4493 451 4494
rect 655 4498 659 4499
rect 655 4493 659 4494
rect 671 4498 675 4499
rect 671 4493 675 4494
rect 887 4498 891 4499
rect 887 4493 891 4494
rect 935 4498 939 4499
rect 935 4493 939 4494
rect 1143 4498 1147 4499
rect 1143 4493 1147 4494
rect 1223 4498 1227 4499
rect 1223 4493 1227 4494
rect 1407 4498 1411 4499
rect 1407 4493 1411 4494
rect 1519 4498 1523 4499
rect 1519 4493 1523 4494
rect 1679 4498 1683 4499
rect 1679 4493 1683 4494
rect 1815 4498 1819 4499
rect 1815 4493 1819 4494
rect 1935 4498 1939 4499
rect 2126 4496 2132 4497
rect 1935 4493 1939 4494
rect 1974 4495 1980 4496
rect 112 4470 114 4493
rect 110 4469 116 4470
rect 448 4469 450 4493
rect 656 4469 658 4493
rect 888 4469 890 4493
rect 1144 4469 1146 4493
rect 1408 4469 1410 4493
rect 1680 4469 1682 4493
rect 1936 4470 1938 4493
rect 1974 4491 1975 4495
rect 1979 4491 1980 4495
rect 2126 4492 2127 4496
rect 2131 4492 2132 4496
rect 2126 4491 2132 4492
rect 2374 4496 2380 4497
rect 2374 4492 2375 4496
rect 2379 4492 2380 4496
rect 2374 4491 2380 4492
rect 2606 4496 2612 4497
rect 2606 4492 2607 4496
rect 2611 4492 2612 4496
rect 2606 4491 2612 4492
rect 2822 4496 2828 4497
rect 2822 4492 2823 4496
rect 2827 4492 2828 4496
rect 2822 4491 2828 4492
rect 3030 4496 3036 4497
rect 3030 4492 3031 4496
rect 3035 4492 3036 4496
rect 3030 4491 3036 4492
rect 3230 4496 3236 4497
rect 3230 4492 3231 4496
rect 3235 4492 3236 4496
rect 3230 4491 3236 4492
rect 3430 4496 3436 4497
rect 3430 4492 3431 4496
rect 3435 4492 3436 4496
rect 3430 4491 3436 4492
rect 3638 4496 3644 4497
rect 3638 4492 3639 4496
rect 3643 4492 3644 4496
rect 3638 4491 3644 4492
rect 3798 4495 3804 4496
rect 3798 4491 3799 4495
rect 3803 4491 3804 4495
rect 1974 4490 1980 4491
rect 1934 4469 1940 4470
rect 110 4465 111 4469
rect 115 4465 116 4469
rect 110 4464 116 4465
rect 446 4468 452 4469
rect 446 4464 447 4468
rect 451 4464 452 4468
rect 446 4463 452 4464
rect 654 4468 660 4469
rect 654 4464 655 4468
rect 659 4464 660 4468
rect 654 4463 660 4464
rect 886 4468 892 4469
rect 886 4464 887 4468
rect 891 4464 892 4468
rect 886 4463 892 4464
rect 1142 4468 1148 4469
rect 1142 4464 1143 4468
rect 1147 4464 1148 4468
rect 1142 4463 1148 4464
rect 1406 4468 1412 4469
rect 1406 4464 1407 4468
rect 1411 4464 1412 4468
rect 1406 4463 1412 4464
rect 1678 4468 1684 4469
rect 1678 4464 1679 4468
rect 1683 4464 1684 4468
rect 1934 4465 1935 4469
rect 1939 4465 1940 4469
rect 1934 4464 1940 4465
rect 1678 4463 1684 4464
rect 1976 4459 1978 4490
rect 2128 4459 2130 4491
rect 2376 4459 2378 4491
rect 2608 4459 2610 4491
rect 2824 4459 2826 4491
rect 3032 4459 3034 4491
rect 3232 4459 3234 4491
rect 3432 4459 3434 4491
rect 3640 4459 3642 4491
rect 3798 4490 3804 4491
rect 3800 4459 3802 4490
rect 3840 4481 3842 4541
rect 3838 4480 3844 4481
rect 4180 4480 4182 4541
rect 4412 4480 4414 4541
rect 4660 4480 4662 4541
rect 4916 4480 4918 4541
rect 5180 4480 5182 4541
rect 5444 4480 5446 4541
rect 5664 4481 5666 4541
rect 5662 4480 5668 4481
rect 3838 4476 3839 4480
rect 3843 4476 3844 4480
rect 3838 4475 3844 4476
rect 4178 4479 4184 4480
rect 4178 4475 4179 4479
rect 4183 4475 4184 4479
rect 4178 4474 4184 4475
rect 4410 4479 4416 4480
rect 4410 4475 4411 4479
rect 4415 4475 4416 4479
rect 4410 4474 4416 4475
rect 4658 4479 4664 4480
rect 4658 4475 4659 4479
rect 4663 4475 4664 4479
rect 4658 4474 4664 4475
rect 4914 4479 4920 4480
rect 4914 4475 4915 4479
rect 4919 4475 4920 4479
rect 4914 4474 4920 4475
rect 5178 4479 5184 4480
rect 5178 4475 5179 4479
rect 5183 4475 5184 4479
rect 5178 4474 5184 4475
rect 5442 4479 5448 4480
rect 5442 4475 5443 4479
rect 5447 4475 5448 4479
rect 5662 4476 5663 4480
rect 5667 4476 5668 4480
rect 5662 4475 5668 4476
rect 5442 4474 5448 4475
rect 4206 4464 4212 4465
rect 3838 4463 3844 4464
rect 3838 4459 3839 4463
rect 3843 4459 3844 4463
rect 4206 4460 4207 4464
rect 4211 4460 4212 4464
rect 4206 4459 4212 4460
rect 4438 4464 4444 4465
rect 4438 4460 4439 4464
rect 4443 4460 4444 4464
rect 4438 4459 4444 4460
rect 4686 4464 4692 4465
rect 4686 4460 4687 4464
rect 4691 4460 4692 4464
rect 4686 4459 4692 4460
rect 4942 4464 4948 4465
rect 4942 4460 4943 4464
rect 4947 4460 4948 4464
rect 4942 4459 4948 4460
rect 5206 4464 5212 4465
rect 5206 4460 5207 4464
rect 5211 4460 5212 4464
rect 5206 4459 5212 4460
rect 5470 4464 5476 4465
rect 5470 4460 5471 4464
rect 5475 4460 5476 4464
rect 5470 4459 5476 4460
rect 5662 4463 5668 4464
rect 5662 4459 5663 4463
rect 5667 4459 5668 4463
rect 1975 4458 1979 4459
rect 418 4453 424 4454
rect 110 4452 116 4453
rect 110 4448 111 4452
rect 115 4448 116 4452
rect 418 4449 419 4453
rect 423 4449 424 4453
rect 418 4448 424 4449
rect 626 4453 632 4454
rect 626 4449 627 4453
rect 631 4449 632 4453
rect 626 4448 632 4449
rect 858 4453 864 4454
rect 858 4449 859 4453
rect 863 4449 864 4453
rect 858 4448 864 4449
rect 1114 4453 1120 4454
rect 1114 4449 1115 4453
rect 1119 4449 1120 4453
rect 1114 4448 1120 4449
rect 1378 4453 1384 4454
rect 1378 4449 1379 4453
rect 1383 4449 1384 4453
rect 1378 4448 1384 4449
rect 1650 4453 1656 4454
rect 1975 4453 1979 4454
rect 2127 4458 2131 4459
rect 2127 4453 2131 4454
rect 2231 4458 2235 4459
rect 2231 4453 2235 4454
rect 2375 4458 2379 4459
rect 2375 4453 2379 4454
rect 2447 4458 2451 4459
rect 2447 4453 2451 4454
rect 2607 4458 2611 4459
rect 2607 4453 2611 4454
rect 2663 4458 2667 4459
rect 2663 4453 2667 4454
rect 2823 4458 2827 4459
rect 2823 4453 2827 4454
rect 2871 4458 2875 4459
rect 2871 4453 2875 4454
rect 3031 4458 3035 4459
rect 3031 4453 3035 4454
rect 3079 4458 3083 4459
rect 3079 4453 3083 4454
rect 3231 4458 3235 4459
rect 3231 4453 3235 4454
rect 3287 4458 3291 4459
rect 3287 4453 3291 4454
rect 3431 4458 3435 4459
rect 3431 4453 3435 4454
rect 3495 4458 3499 4459
rect 3495 4453 3499 4454
rect 3639 4458 3643 4459
rect 3639 4453 3643 4454
rect 3679 4458 3683 4459
rect 3679 4453 3683 4454
rect 3799 4458 3803 4459
rect 3838 4458 3844 4459
rect 3799 4453 3803 4454
rect 1650 4449 1651 4453
rect 1655 4449 1656 4453
rect 1650 4448 1656 4449
rect 1934 4452 1940 4453
rect 1934 4448 1935 4452
rect 1939 4448 1940 4452
rect 110 4447 116 4448
rect 112 4383 114 4447
rect 420 4383 422 4448
rect 628 4383 630 4448
rect 860 4383 862 4448
rect 1116 4383 1118 4448
rect 1380 4383 1382 4448
rect 1652 4383 1654 4448
rect 1934 4447 1940 4448
rect 1936 4383 1938 4447
rect 1976 4430 1978 4453
rect 1974 4429 1980 4430
rect 2232 4429 2234 4453
rect 2448 4429 2450 4453
rect 2664 4429 2666 4453
rect 2872 4429 2874 4453
rect 3080 4429 3082 4453
rect 3288 4429 3290 4453
rect 3496 4429 3498 4453
rect 3680 4429 3682 4453
rect 3800 4430 3802 4453
rect 3798 4429 3804 4430
rect 1974 4425 1975 4429
rect 1979 4425 1980 4429
rect 1974 4424 1980 4425
rect 2230 4428 2236 4429
rect 2230 4424 2231 4428
rect 2235 4424 2236 4428
rect 2230 4423 2236 4424
rect 2446 4428 2452 4429
rect 2446 4424 2447 4428
rect 2451 4424 2452 4428
rect 2446 4423 2452 4424
rect 2662 4428 2668 4429
rect 2662 4424 2663 4428
rect 2667 4424 2668 4428
rect 2662 4423 2668 4424
rect 2870 4428 2876 4429
rect 2870 4424 2871 4428
rect 2875 4424 2876 4428
rect 2870 4423 2876 4424
rect 3078 4428 3084 4429
rect 3078 4424 3079 4428
rect 3083 4424 3084 4428
rect 3078 4423 3084 4424
rect 3286 4428 3292 4429
rect 3286 4424 3287 4428
rect 3291 4424 3292 4428
rect 3286 4423 3292 4424
rect 3494 4428 3500 4429
rect 3494 4424 3495 4428
rect 3499 4424 3500 4428
rect 3494 4423 3500 4424
rect 3678 4428 3684 4429
rect 3678 4424 3679 4428
rect 3683 4424 3684 4428
rect 3798 4425 3799 4429
rect 3803 4425 3804 4429
rect 3840 4427 3842 4458
rect 4208 4427 4210 4459
rect 4440 4427 4442 4459
rect 4688 4427 4690 4459
rect 4944 4427 4946 4459
rect 5208 4427 5210 4459
rect 5472 4427 5474 4459
rect 5662 4458 5668 4459
rect 5664 4427 5666 4458
rect 3798 4424 3804 4425
rect 3839 4426 3843 4427
rect 3678 4423 3684 4424
rect 3839 4421 3843 4422
rect 4207 4426 4211 4427
rect 4207 4421 4211 4422
rect 4359 4426 4363 4427
rect 4359 4421 4363 4422
rect 4439 4426 4443 4427
rect 4439 4421 4443 4422
rect 4519 4426 4523 4427
rect 4519 4421 4523 4422
rect 4687 4426 4691 4427
rect 4687 4421 4691 4422
rect 4879 4426 4883 4427
rect 4879 4421 4883 4422
rect 4943 4426 4947 4427
rect 4943 4421 4947 4422
rect 5079 4426 5083 4427
rect 5079 4421 5083 4422
rect 5207 4426 5211 4427
rect 5207 4421 5211 4422
rect 5287 4426 5291 4427
rect 5287 4421 5291 4422
rect 5471 4426 5475 4427
rect 5471 4421 5475 4422
rect 5503 4426 5507 4427
rect 5503 4421 5507 4422
rect 5663 4426 5667 4427
rect 5663 4421 5667 4422
rect 2202 4413 2208 4414
rect 1974 4412 1980 4413
rect 1974 4408 1975 4412
rect 1979 4408 1980 4412
rect 2202 4409 2203 4413
rect 2207 4409 2208 4413
rect 2202 4408 2208 4409
rect 2418 4413 2424 4414
rect 2418 4409 2419 4413
rect 2423 4409 2424 4413
rect 2418 4408 2424 4409
rect 2634 4413 2640 4414
rect 2634 4409 2635 4413
rect 2639 4409 2640 4413
rect 2634 4408 2640 4409
rect 2842 4413 2848 4414
rect 2842 4409 2843 4413
rect 2847 4409 2848 4413
rect 2842 4408 2848 4409
rect 3050 4413 3056 4414
rect 3050 4409 3051 4413
rect 3055 4409 3056 4413
rect 3050 4408 3056 4409
rect 3258 4413 3264 4414
rect 3258 4409 3259 4413
rect 3263 4409 3264 4413
rect 3258 4408 3264 4409
rect 3466 4413 3472 4414
rect 3466 4409 3467 4413
rect 3471 4409 3472 4413
rect 3466 4408 3472 4409
rect 3650 4413 3656 4414
rect 3650 4409 3651 4413
rect 3655 4409 3656 4413
rect 3650 4408 3656 4409
rect 3798 4412 3804 4413
rect 3798 4408 3799 4412
rect 3803 4408 3804 4412
rect 1974 4407 1980 4408
rect 111 4382 115 4383
rect 111 4377 115 4378
rect 419 4382 423 4383
rect 419 4377 423 4378
rect 627 4382 631 4383
rect 627 4377 631 4378
rect 667 4382 671 4383
rect 667 4377 671 4378
rect 811 4382 815 4383
rect 811 4377 815 4378
rect 859 4382 863 4383
rect 859 4377 863 4378
rect 963 4382 967 4383
rect 963 4377 967 4378
rect 1115 4382 1119 4383
rect 1115 4377 1119 4378
rect 1123 4382 1127 4383
rect 1123 4377 1127 4378
rect 1291 4382 1295 4383
rect 1291 4377 1295 4378
rect 1379 4382 1383 4383
rect 1379 4377 1383 4378
rect 1467 4382 1471 4383
rect 1467 4377 1471 4378
rect 1651 4382 1655 4383
rect 1651 4377 1655 4378
rect 1935 4382 1939 4383
rect 1935 4377 1939 4378
rect 112 4317 114 4377
rect 110 4316 116 4317
rect 668 4316 670 4377
rect 812 4316 814 4377
rect 964 4316 966 4377
rect 1124 4316 1126 4377
rect 1292 4316 1294 4377
rect 1468 4316 1470 4377
rect 1652 4316 1654 4377
rect 1936 4317 1938 4377
rect 1976 4339 1978 4407
rect 2204 4339 2206 4408
rect 2420 4339 2422 4408
rect 2636 4339 2638 4408
rect 2844 4339 2846 4408
rect 3052 4339 3054 4408
rect 3260 4339 3262 4408
rect 3468 4339 3470 4408
rect 3652 4339 3654 4408
rect 3798 4407 3804 4408
rect 3800 4339 3802 4407
rect 3840 4398 3842 4421
rect 3838 4397 3844 4398
rect 4360 4397 4362 4421
rect 4520 4397 4522 4421
rect 4688 4397 4690 4421
rect 4880 4397 4882 4421
rect 5080 4397 5082 4421
rect 5288 4397 5290 4421
rect 5504 4397 5506 4421
rect 5664 4398 5666 4421
rect 5662 4397 5668 4398
rect 3838 4393 3839 4397
rect 3843 4393 3844 4397
rect 3838 4392 3844 4393
rect 4358 4396 4364 4397
rect 4358 4392 4359 4396
rect 4363 4392 4364 4396
rect 4358 4391 4364 4392
rect 4518 4396 4524 4397
rect 4518 4392 4519 4396
rect 4523 4392 4524 4396
rect 4518 4391 4524 4392
rect 4686 4396 4692 4397
rect 4686 4392 4687 4396
rect 4691 4392 4692 4396
rect 4686 4391 4692 4392
rect 4878 4396 4884 4397
rect 4878 4392 4879 4396
rect 4883 4392 4884 4396
rect 4878 4391 4884 4392
rect 5078 4396 5084 4397
rect 5078 4392 5079 4396
rect 5083 4392 5084 4396
rect 5078 4391 5084 4392
rect 5286 4396 5292 4397
rect 5286 4392 5287 4396
rect 5291 4392 5292 4396
rect 5286 4391 5292 4392
rect 5502 4396 5508 4397
rect 5502 4392 5503 4396
rect 5507 4392 5508 4396
rect 5662 4393 5663 4397
rect 5667 4393 5668 4397
rect 5662 4392 5668 4393
rect 5502 4391 5508 4392
rect 4330 4381 4336 4382
rect 3838 4380 3844 4381
rect 3838 4376 3839 4380
rect 3843 4376 3844 4380
rect 4330 4377 4331 4381
rect 4335 4377 4336 4381
rect 4330 4376 4336 4377
rect 4490 4381 4496 4382
rect 4490 4377 4491 4381
rect 4495 4377 4496 4381
rect 4490 4376 4496 4377
rect 4658 4381 4664 4382
rect 4658 4377 4659 4381
rect 4663 4377 4664 4381
rect 4658 4376 4664 4377
rect 4850 4381 4856 4382
rect 4850 4377 4851 4381
rect 4855 4377 4856 4381
rect 4850 4376 4856 4377
rect 5050 4381 5056 4382
rect 5050 4377 5051 4381
rect 5055 4377 5056 4381
rect 5050 4376 5056 4377
rect 5258 4381 5264 4382
rect 5258 4377 5259 4381
rect 5263 4377 5264 4381
rect 5258 4376 5264 4377
rect 5474 4381 5480 4382
rect 5474 4377 5475 4381
rect 5479 4377 5480 4381
rect 5474 4376 5480 4377
rect 5662 4380 5668 4381
rect 5662 4376 5663 4380
rect 5667 4376 5668 4380
rect 3838 4375 3844 4376
rect 1975 4338 1979 4339
rect 1975 4333 1979 4334
rect 2203 4338 2207 4339
rect 2203 4333 2207 4334
rect 2307 4338 2311 4339
rect 2307 4333 2311 4334
rect 2419 4338 2423 4339
rect 2419 4333 2423 4334
rect 2459 4338 2463 4339
rect 2459 4333 2463 4334
rect 2627 4338 2631 4339
rect 2627 4333 2631 4334
rect 2635 4338 2639 4339
rect 2635 4333 2639 4334
rect 2811 4338 2815 4339
rect 2811 4333 2815 4334
rect 2843 4338 2847 4339
rect 2843 4333 2847 4334
rect 3011 4338 3015 4339
rect 3011 4333 3015 4334
rect 3051 4338 3055 4339
rect 3051 4333 3055 4334
rect 3227 4338 3231 4339
rect 3227 4333 3231 4334
rect 3259 4338 3263 4339
rect 3259 4333 3263 4334
rect 3451 4338 3455 4339
rect 3451 4333 3455 4334
rect 3467 4338 3471 4339
rect 3467 4333 3471 4334
rect 3651 4338 3655 4339
rect 3651 4333 3655 4334
rect 3799 4338 3803 4339
rect 3799 4333 3803 4334
rect 1934 4316 1940 4317
rect 110 4312 111 4316
rect 115 4312 116 4316
rect 110 4311 116 4312
rect 666 4315 672 4316
rect 666 4311 667 4315
rect 671 4311 672 4315
rect 666 4310 672 4311
rect 810 4315 816 4316
rect 810 4311 811 4315
rect 815 4311 816 4315
rect 810 4310 816 4311
rect 962 4315 968 4316
rect 962 4311 963 4315
rect 967 4311 968 4315
rect 962 4310 968 4311
rect 1122 4315 1128 4316
rect 1122 4311 1123 4315
rect 1127 4311 1128 4315
rect 1122 4310 1128 4311
rect 1290 4315 1296 4316
rect 1290 4311 1291 4315
rect 1295 4311 1296 4315
rect 1290 4310 1296 4311
rect 1466 4315 1472 4316
rect 1466 4311 1467 4315
rect 1471 4311 1472 4315
rect 1466 4310 1472 4311
rect 1650 4315 1656 4316
rect 1650 4311 1651 4315
rect 1655 4311 1656 4315
rect 1934 4312 1935 4316
rect 1939 4312 1940 4316
rect 1934 4311 1940 4312
rect 1650 4310 1656 4311
rect 694 4300 700 4301
rect 110 4299 116 4300
rect 110 4295 111 4299
rect 115 4295 116 4299
rect 694 4296 695 4300
rect 699 4296 700 4300
rect 694 4295 700 4296
rect 838 4300 844 4301
rect 838 4296 839 4300
rect 843 4296 844 4300
rect 838 4295 844 4296
rect 990 4300 996 4301
rect 990 4296 991 4300
rect 995 4296 996 4300
rect 990 4295 996 4296
rect 1150 4300 1156 4301
rect 1150 4296 1151 4300
rect 1155 4296 1156 4300
rect 1150 4295 1156 4296
rect 1318 4300 1324 4301
rect 1318 4296 1319 4300
rect 1323 4296 1324 4300
rect 1318 4295 1324 4296
rect 1494 4300 1500 4301
rect 1494 4296 1495 4300
rect 1499 4296 1500 4300
rect 1494 4295 1500 4296
rect 1678 4300 1684 4301
rect 1678 4296 1679 4300
rect 1683 4296 1684 4300
rect 1678 4295 1684 4296
rect 1934 4299 1940 4300
rect 1934 4295 1935 4299
rect 1939 4295 1940 4299
rect 110 4294 116 4295
rect 112 4255 114 4294
rect 696 4255 698 4295
rect 840 4255 842 4295
rect 992 4255 994 4295
rect 1152 4255 1154 4295
rect 1320 4255 1322 4295
rect 1496 4255 1498 4295
rect 1680 4255 1682 4295
rect 1934 4294 1940 4295
rect 1936 4255 1938 4294
rect 1976 4273 1978 4333
rect 1974 4272 1980 4273
rect 2308 4272 2310 4333
rect 2460 4272 2462 4333
rect 2628 4272 2630 4333
rect 2812 4272 2814 4333
rect 3012 4272 3014 4333
rect 3228 4272 3230 4333
rect 3452 4272 3454 4333
rect 3652 4272 3654 4333
rect 3800 4273 3802 4333
rect 3840 4315 3842 4375
rect 4332 4315 4334 4376
rect 4492 4315 4494 4376
rect 4660 4315 4662 4376
rect 4852 4315 4854 4376
rect 5052 4315 5054 4376
rect 5260 4315 5262 4376
rect 5476 4315 5478 4376
rect 5662 4375 5668 4376
rect 5664 4315 5666 4375
rect 3839 4314 3843 4315
rect 3839 4309 3843 4310
rect 3859 4314 3863 4315
rect 3859 4309 3863 4310
rect 4043 4314 4047 4315
rect 4043 4309 4047 4310
rect 4251 4314 4255 4315
rect 4251 4309 4255 4310
rect 4331 4314 4335 4315
rect 4331 4309 4335 4310
rect 4475 4314 4479 4315
rect 4475 4309 4479 4310
rect 4491 4314 4495 4315
rect 4491 4309 4495 4310
rect 4659 4314 4663 4315
rect 4659 4309 4663 4310
rect 4715 4314 4719 4315
rect 4715 4309 4719 4310
rect 4851 4314 4855 4315
rect 4851 4309 4855 4310
rect 4971 4314 4975 4315
rect 4971 4309 4975 4310
rect 5051 4314 5055 4315
rect 5051 4309 5055 4310
rect 5235 4314 5239 4315
rect 5235 4309 5239 4310
rect 5259 4314 5263 4315
rect 5259 4309 5263 4310
rect 5475 4314 5479 4315
rect 5475 4309 5479 4310
rect 5499 4314 5503 4315
rect 5499 4309 5503 4310
rect 5663 4314 5667 4315
rect 5663 4309 5667 4310
rect 3798 4272 3804 4273
rect 1974 4268 1975 4272
rect 1979 4268 1980 4272
rect 1974 4267 1980 4268
rect 2306 4271 2312 4272
rect 2306 4267 2307 4271
rect 2311 4267 2312 4271
rect 2306 4266 2312 4267
rect 2458 4271 2464 4272
rect 2458 4267 2459 4271
rect 2463 4267 2464 4271
rect 2458 4266 2464 4267
rect 2626 4271 2632 4272
rect 2626 4267 2627 4271
rect 2631 4267 2632 4271
rect 2626 4266 2632 4267
rect 2810 4271 2816 4272
rect 2810 4267 2811 4271
rect 2815 4267 2816 4271
rect 2810 4266 2816 4267
rect 3010 4271 3016 4272
rect 3010 4267 3011 4271
rect 3015 4267 3016 4271
rect 3010 4266 3016 4267
rect 3226 4271 3232 4272
rect 3226 4267 3227 4271
rect 3231 4267 3232 4271
rect 3226 4266 3232 4267
rect 3450 4271 3456 4272
rect 3450 4267 3451 4271
rect 3455 4267 3456 4271
rect 3450 4266 3456 4267
rect 3650 4271 3656 4272
rect 3650 4267 3651 4271
rect 3655 4267 3656 4271
rect 3798 4268 3799 4272
rect 3803 4268 3804 4272
rect 3798 4267 3804 4268
rect 3650 4266 3656 4267
rect 2334 4256 2340 4257
rect 1974 4255 1980 4256
rect 111 4254 115 4255
rect 111 4249 115 4250
rect 695 4254 699 4255
rect 695 4249 699 4250
rect 815 4254 819 4255
rect 815 4249 819 4250
rect 839 4254 843 4255
rect 839 4249 843 4250
rect 951 4254 955 4255
rect 951 4249 955 4250
rect 991 4254 995 4255
rect 991 4249 995 4250
rect 1087 4254 1091 4255
rect 1087 4249 1091 4250
rect 1151 4254 1155 4255
rect 1151 4249 1155 4250
rect 1223 4254 1227 4255
rect 1223 4249 1227 4250
rect 1319 4254 1323 4255
rect 1319 4249 1323 4250
rect 1359 4254 1363 4255
rect 1359 4249 1363 4250
rect 1495 4254 1499 4255
rect 1495 4249 1499 4250
rect 1631 4254 1635 4255
rect 1631 4249 1635 4250
rect 1679 4254 1683 4255
rect 1679 4249 1683 4250
rect 1767 4254 1771 4255
rect 1767 4249 1771 4250
rect 1935 4254 1939 4255
rect 1974 4251 1975 4255
rect 1979 4251 1980 4255
rect 2334 4252 2335 4256
rect 2339 4252 2340 4256
rect 2334 4251 2340 4252
rect 2486 4256 2492 4257
rect 2486 4252 2487 4256
rect 2491 4252 2492 4256
rect 2486 4251 2492 4252
rect 2654 4256 2660 4257
rect 2654 4252 2655 4256
rect 2659 4252 2660 4256
rect 2654 4251 2660 4252
rect 2838 4256 2844 4257
rect 2838 4252 2839 4256
rect 2843 4252 2844 4256
rect 2838 4251 2844 4252
rect 3038 4256 3044 4257
rect 3038 4252 3039 4256
rect 3043 4252 3044 4256
rect 3038 4251 3044 4252
rect 3254 4256 3260 4257
rect 3254 4252 3255 4256
rect 3259 4252 3260 4256
rect 3254 4251 3260 4252
rect 3478 4256 3484 4257
rect 3478 4252 3479 4256
rect 3483 4252 3484 4256
rect 3478 4251 3484 4252
rect 3678 4256 3684 4257
rect 3678 4252 3679 4256
rect 3683 4252 3684 4256
rect 3678 4251 3684 4252
rect 3798 4255 3804 4256
rect 3798 4251 3799 4255
rect 3803 4251 3804 4255
rect 1974 4250 1980 4251
rect 1935 4249 1939 4250
rect 112 4226 114 4249
rect 110 4225 116 4226
rect 816 4225 818 4249
rect 952 4225 954 4249
rect 1088 4225 1090 4249
rect 1224 4225 1226 4249
rect 1360 4225 1362 4249
rect 1496 4225 1498 4249
rect 1632 4225 1634 4249
rect 1768 4225 1770 4249
rect 1936 4226 1938 4249
rect 1934 4225 1940 4226
rect 110 4221 111 4225
rect 115 4221 116 4225
rect 110 4220 116 4221
rect 814 4224 820 4225
rect 814 4220 815 4224
rect 819 4220 820 4224
rect 814 4219 820 4220
rect 950 4224 956 4225
rect 950 4220 951 4224
rect 955 4220 956 4224
rect 950 4219 956 4220
rect 1086 4224 1092 4225
rect 1086 4220 1087 4224
rect 1091 4220 1092 4224
rect 1086 4219 1092 4220
rect 1222 4224 1228 4225
rect 1222 4220 1223 4224
rect 1227 4220 1228 4224
rect 1222 4219 1228 4220
rect 1358 4224 1364 4225
rect 1358 4220 1359 4224
rect 1363 4220 1364 4224
rect 1358 4219 1364 4220
rect 1494 4224 1500 4225
rect 1494 4220 1495 4224
rect 1499 4220 1500 4224
rect 1494 4219 1500 4220
rect 1630 4224 1636 4225
rect 1630 4220 1631 4224
rect 1635 4220 1636 4224
rect 1630 4219 1636 4220
rect 1766 4224 1772 4225
rect 1766 4220 1767 4224
rect 1771 4220 1772 4224
rect 1934 4221 1935 4225
rect 1939 4221 1940 4225
rect 1934 4220 1940 4221
rect 1766 4219 1772 4220
rect 1976 4219 1978 4250
rect 2336 4219 2338 4251
rect 2488 4219 2490 4251
rect 2656 4219 2658 4251
rect 2840 4219 2842 4251
rect 3040 4219 3042 4251
rect 3256 4219 3258 4251
rect 3480 4219 3482 4251
rect 3680 4219 3682 4251
rect 3798 4250 3804 4251
rect 3800 4219 3802 4250
rect 3840 4249 3842 4309
rect 3838 4248 3844 4249
rect 3860 4248 3862 4309
rect 4044 4248 4046 4309
rect 4252 4248 4254 4309
rect 4476 4248 4478 4309
rect 4716 4248 4718 4309
rect 4972 4248 4974 4309
rect 5236 4248 5238 4309
rect 5500 4248 5502 4309
rect 5664 4249 5666 4309
rect 5662 4248 5668 4249
rect 3838 4244 3839 4248
rect 3843 4244 3844 4248
rect 3838 4243 3844 4244
rect 3858 4247 3864 4248
rect 3858 4243 3859 4247
rect 3863 4243 3864 4247
rect 3858 4242 3864 4243
rect 4042 4247 4048 4248
rect 4042 4243 4043 4247
rect 4047 4243 4048 4247
rect 4042 4242 4048 4243
rect 4250 4247 4256 4248
rect 4250 4243 4251 4247
rect 4255 4243 4256 4247
rect 4250 4242 4256 4243
rect 4474 4247 4480 4248
rect 4474 4243 4475 4247
rect 4479 4243 4480 4247
rect 4474 4242 4480 4243
rect 4714 4247 4720 4248
rect 4714 4243 4715 4247
rect 4719 4243 4720 4247
rect 4714 4242 4720 4243
rect 4970 4247 4976 4248
rect 4970 4243 4971 4247
rect 4975 4243 4976 4247
rect 4970 4242 4976 4243
rect 5234 4247 5240 4248
rect 5234 4243 5235 4247
rect 5239 4243 5240 4247
rect 5234 4242 5240 4243
rect 5498 4247 5504 4248
rect 5498 4243 5499 4247
rect 5503 4243 5504 4247
rect 5662 4244 5663 4248
rect 5667 4244 5668 4248
rect 5662 4243 5668 4244
rect 5498 4242 5504 4243
rect 3886 4232 3892 4233
rect 3838 4231 3844 4232
rect 3838 4227 3839 4231
rect 3843 4227 3844 4231
rect 3886 4228 3887 4232
rect 3891 4228 3892 4232
rect 3886 4227 3892 4228
rect 4070 4232 4076 4233
rect 4070 4228 4071 4232
rect 4075 4228 4076 4232
rect 4070 4227 4076 4228
rect 4278 4232 4284 4233
rect 4278 4228 4279 4232
rect 4283 4228 4284 4232
rect 4278 4227 4284 4228
rect 4502 4232 4508 4233
rect 4502 4228 4503 4232
rect 4507 4228 4508 4232
rect 4502 4227 4508 4228
rect 4742 4232 4748 4233
rect 4742 4228 4743 4232
rect 4747 4228 4748 4232
rect 4742 4227 4748 4228
rect 4998 4232 5004 4233
rect 4998 4228 4999 4232
rect 5003 4228 5004 4232
rect 4998 4227 5004 4228
rect 5262 4232 5268 4233
rect 5262 4228 5263 4232
rect 5267 4228 5268 4232
rect 5262 4227 5268 4228
rect 5526 4232 5532 4233
rect 5526 4228 5527 4232
rect 5531 4228 5532 4232
rect 5526 4227 5532 4228
rect 5662 4231 5668 4232
rect 5662 4227 5663 4231
rect 5667 4227 5668 4231
rect 3838 4226 3844 4227
rect 1975 4218 1979 4219
rect 1975 4213 1979 4214
rect 2335 4218 2339 4219
rect 2335 4213 2339 4214
rect 2487 4218 2491 4219
rect 2487 4213 2491 4214
rect 2567 4218 2571 4219
rect 2567 4213 2571 4214
rect 2655 4218 2659 4219
rect 2655 4213 2659 4214
rect 2703 4218 2707 4219
rect 2703 4213 2707 4214
rect 2839 4218 2843 4219
rect 2839 4213 2843 4214
rect 2975 4218 2979 4219
rect 2975 4213 2979 4214
rect 3039 4218 3043 4219
rect 3039 4213 3043 4214
rect 3255 4218 3259 4219
rect 3255 4213 3259 4214
rect 3479 4218 3483 4219
rect 3479 4213 3483 4214
rect 3679 4218 3683 4219
rect 3679 4213 3683 4214
rect 3799 4218 3803 4219
rect 3799 4213 3803 4214
rect 786 4209 792 4210
rect 110 4208 116 4209
rect 110 4204 111 4208
rect 115 4204 116 4208
rect 786 4205 787 4209
rect 791 4205 792 4209
rect 786 4204 792 4205
rect 922 4209 928 4210
rect 922 4205 923 4209
rect 927 4205 928 4209
rect 922 4204 928 4205
rect 1058 4209 1064 4210
rect 1058 4205 1059 4209
rect 1063 4205 1064 4209
rect 1058 4204 1064 4205
rect 1194 4209 1200 4210
rect 1194 4205 1195 4209
rect 1199 4205 1200 4209
rect 1194 4204 1200 4205
rect 1330 4209 1336 4210
rect 1330 4205 1331 4209
rect 1335 4205 1336 4209
rect 1330 4204 1336 4205
rect 1466 4209 1472 4210
rect 1466 4205 1467 4209
rect 1471 4205 1472 4209
rect 1466 4204 1472 4205
rect 1602 4209 1608 4210
rect 1602 4205 1603 4209
rect 1607 4205 1608 4209
rect 1602 4204 1608 4205
rect 1738 4209 1744 4210
rect 1738 4205 1739 4209
rect 1743 4205 1744 4209
rect 1738 4204 1744 4205
rect 1934 4208 1940 4209
rect 1934 4204 1935 4208
rect 1939 4204 1940 4208
rect 110 4203 116 4204
rect 112 4139 114 4203
rect 788 4139 790 4204
rect 924 4139 926 4204
rect 1060 4139 1062 4204
rect 1196 4139 1198 4204
rect 1332 4139 1334 4204
rect 1468 4139 1470 4204
rect 1604 4139 1606 4204
rect 1740 4139 1742 4204
rect 1934 4203 1940 4204
rect 1936 4139 1938 4203
rect 1976 4190 1978 4213
rect 1974 4189 1980 4190
rect 2568 4189 2570 4213
rect 2704 4189 2706 4213
rect 2840 4189 2842 4213
rect 2976 4189 2978 4213
rect 3800 4190 3802 4213
rect 3798 4189 3804 4190
rect 1974 4185 1975 4189
rect 1979 4185 1980 4189
rect 1974 4184 1980 4185
rect 2566 4188 2572 4189
rect 2566 4184 2567 4188
rect 2571 4184 2572 4188
rect 2566 4183 2572 4184
rect 2702 4188 2708 4189
rect 2702 4184 2703 4188
rect 2707 4184 2708 4188
rect 2702 4183 2708 4184
rect 2838 4188 2844 4189
rect 2838 4184 2839 4188
rect 2843 4184 2844 4188
rect 2838 4183 2844 4184
rect 2974 4188 2980 4189
rect 2974 4184 2975 4188
rect 2979 4184 2980 4188
rect 3798 4185 3799 4189
rect 3803 4185 3804 4189
rect 3798 4184 3804 4185
rect 2974 4183 2980 4184
rect 2538 4173 2544 4174
rect 1974 4172 1980 4173
rect 1974 4168 1975 4172
rect 1979 4168 1980 4172
rect 2538 4169 2539 4173
rect 2543 4169 2544 4173
rect 2538 4168 2544 4169
rect 2674 4173 2680 4174
rect 2674 4169 2675 4173
rect 2679 4169 2680 4173
rect 2674 4168 2680 4169
rect 2810 4173 2816 4174
rect 2810 4169 2811 4173
rect 2815 4169 2816 4173
rect 2810 4168 2816 4169
rect 2946 4173 2952 4174
rect 2946 4169 2947 4173
rect 2951 4169 2952 4173
rect 2946 4168 2952 4169
rect 3798 4172 3804 4173
rect 3798 4168 3799 4172
rect 3803 4168 3804 4172
rect 1974 4167 1980 4168
rect 111 4138 115 4139
rect 111 4133 115 4134
rect 731 4138 735 4139
rect 731 4133 735 4134
rect 787 4138 791 4139
rect 787 4133 791 4134
rect 867 4138 871 4139
rect 867 4133 871 4134
rect 923 4138 927 4139
rect 923 4133 927 4134
rect 1003 4138 1007 4139
rect 1003 4133 1007 4134
rect 1059 4138 1063 4139
rect 1059 4133 1063 4134
rect 1139 4138 1143 4139
rect 1139 4133 1143 4134
rect 1195 4138 1199 4139
rect 1195 4133 1199 4134
rect 1275 4138 1279 4139
rect 1275 4133 1279 4134
rect 1331 4138 1335 4139
rect 1331 4133 1335 4134
rect 1411 4138 1415 4139
rect 1411 4133 1415 4134
rect 1467 4138 1471 4139
rect 1467 4133 1471 4134
rect 1547 4138 1551 4139
rect 1547 4133 1551 4134
rect 1603 4138 1607 4139
rect 1603 4133 1607 4134
rect 1739 4138 1743 4139
rect 1739 4133 1743 4134
rect 1935 4138 1939 4139
rect 1935 4133 1939 4134
rect 112 4073 114 4133
rect 110 4072 116 4073
rect 732 4072 734 4133
rect 868 4072 870 4133
rect 1004 4072 1006 4133
rect 1140 4072 1142 4133
rect 1276 4072 1278 4133
rect 1412 4072 1414 4133
rect 1548 4072 1550 4133
rect 1936 4073 1938 4133
rect 1976 4087 1978 4167
rect 2540 4087 2542 4168
rect 2676 4087 2678 4168
rect 2812 4087 2814 4168
rect 2948 4087 2950 4168
rect 3798 4167 3804 4168
rect 3840 4167 3842 4226
rect 3888 4167 3890 4227
rect 4072 4167 4074 4227
rect 4280 4167 4282 4227
rect 4504 4167 4506 4227
rect 4744 4167 4746 4227
rect 5000 4167 5002 4227
rect 5264 4167 5266 4227
rect 5528 4167 5530 4227
rect 5662 4226 5668 4227
rect 5664 4167 5666 4226
rect 3800 4087 3802 4167
rect 3839 4166 3843 4167
rect 3839 4161 3843 4162
rect 3887 4166 3891 4167
rect 3887 4161 3891 4162
rect 4071 4166 4075 4167
rect 4071 4161 4075 4162
rect 4279 4166 4283 4167
rect 4279 4161 4283 4162
rect 4415 4166 4419 4167
rect 4415 4161 4419 4162
rect 4503 4166 4507 4167
rect 4503 4161 4507 4162
rect 4743 4166 4747 4167
rect 4743 4161 4747 4162
rect 4975 4166 4979 4167
rect 4975 4161 4979 4162
rect 4999 4166 5003 4167
rect 4999 4161 5003 4162
rect 5263 4166 5267 4167
rect 5263 4161 5267 4162
rect 5527 4166 5531 4167
rect 5527 4161 5531 4162
rect 5543 4166 5547 4167
rect 5543 4161 5547 4162
rect 5663 4166 5667 4167
rect 5663 4161 5667 4162
rect 3840 4138 3842 4161
rect 3838 4137 3844 4138
rect 3888 4137 3890 4161
rect 4416 4137 4418 4161
rect 4976 4137 4978 4161
rect 5544 4137 5546 4161
rect 5664 4138 5666 4161
rect 5662 4137 5668 4138
rect 3838 4133 3839 4137
rect 3843 4133 3844 4137
rect 3838 4132 3844 4133
rect 3886 4136 3892 4137
rect 3886 4132 3887 4136
rect 3891 4132 3892 4136
rect 3886 4131 3892 4132
rect 4414 4136 4420 4137
rect 4414 4132 4415 4136
rect 4419 4132 4420 4136
rect 4414 4131 4420 4132
rect 4974 4136 4980 4137
rect 4974 4132 4975 4136
rect 4979 4132 4980 4136
rect 4974 4131 4980 4132
rect 5542 4136 5548 4137
rect 5542 4132 5543 4136
rect 5547 4132 5548 4136
rect 5662 4133 5663 4137
rect 5667 4133 5668 4137
rect 5662 4132 5668 4133
rect 5542 4131 5548 4132
rect 3858 4121 3864 4122
rect 3838 4120 3844 4121
rect 3838 4116 3839 4120
rect 3843 4116 3844 4120
rect 3858 4117 3859 4121
rect 3863 4117 3864 4121
rect 3858 4116 3864 4117
rect 4386 4121 4392 4122
rect 4386 4117 4387 4121
rect 4391 4117 4392 4121
rect 4386 4116 4392 4117
rect 4946 4121 4952 4122
rect 4946 4117 4947 4121
rect 4951 4117 4952 4121
rect 4946 4116 4952 4117
rect 5514 4121 5520 4122
rect 5514 4117 5515 4121
rect 5519 4117 5520 4121
rect 5514 4116 5520 4117
rect 5662 4120 5668 4121
rect 5662 4116 5663 4120
rect 5667 4116 5668 4120
rect 3838 4115 3844 4116
rect 1975 4086 1979 4087
rect 1975 4081 1979 4082
rect 2291 4086 2295 4087
rect 2291 4081 2295 4082
rect 2427 4086 2431 4087
rect 2427 4081 2431 4082
rect 2539 4086 2543 4087
rect 2539 4081 2543 4082
rect 2563 4086 2567 4087
rect 2563 4081 2567 4082
rect 2675 4086 2679 4087
rect 2675 4081 2679 4082
rect 2699 4086 2703 4087
rect 2699 4081 2703 4082
rect 2811 4086 2815 4087
rect 2811 4081 2815 4082
rect 2835 4086 2839 4087
rect 2835 4081 2839 4082
rect 2947 4086 2951 4087
rect 2947 4081 2951 4082
rect 3799 4086 3803 4087
rect 3799 4081 3803 4082
rect 1934 4072 1940 4073
rect 110 4068 111 4072
rect 115 4068 116 4072
rect 110 4067 116 4068
rect 730 4071 736 4072
rect 730 4067 731 4071
rect 735 4067 736 4071
rect 730 4066 736 4067
rect 866 4071 872 4072
rect 866 4067 867 4071
rect 871 4067 872 4071
rect 866 4066 872 4067
rect 1002 4071 1008 4072
rect 1002 4067 1003 4071
rect 1007 4067 1008 4071
rect 1002 4066 1008 4067
rect 1138 4071 1144 4072
rect 1138 4067 1139 4071
rect 1143 4067 1144 4071
rect 1138 4066 1144 4067
rect 1274 4071 1280 4072
rect 1274 4067 1275 4071
rect 1279 4067 1280 4071
rect 1274 4066 1280 4067
rect 1410 4071 1416 4072
rect 1410 4067 1411 4071
rect 1415 4067 1416 4071
rect 1410 4066 1416 4067
rect 1546 4071 1552 4072
rect 1546 4067 1547 4071
rect 1551 4067 1552 4071
rect 1934 4068 1935 4072
rect 1939 4068 1940 4072
rect 1934 4067 1940 4068
rect 1546 4066 1552 4067
rect 758 4056 764 4057
rect 110 4055 116 4056
rect 110 4051 111 4055
rect 115 4051 116 4055
rect 758 4052 759 4056
rect 763 4052 764 4056
rect 758 4051 764 4052
rect 894 4056 900 4057
rect 894 4052 895 4056
rect 899 4052 900 4056
rect 894 4051 900 4052
rect 1030 4056 1036 4057
rect 1030 4052 1031 4056
rect 1035 4052 1036 4056
rect 1030 4051 1036 4052
rect 1166 4056 1172 4057
rect 1166 4052 1167 4056
rect 1171 4052 1172 4056
rect 1166 4051 1172 4052
rect 1302 4056 1308 4057
rect 1302 4052 1303 4056
rect 1307 4052 1308 4056
rect 1302 4051 1308 4052
rect 1438 4056 1444 4057
rect 1438 4052 1439 4056
rect 1443 4052 1444 4056
rect 1438 4051 1444 4052
rect 1574 4056 1580 4057
rect 1574 4052 1575 4056
rect 1579 4052 1580 4056
rect 1574 4051 1580 4052
rect 1934 4055 1940 4056
rect 1934 4051 1935 4055
rect 1939 4051 1940 4055
rect 110 4050 116 4051
rect 112 4003 114 4050
rect 760 4003 762 4051
rect 896 4003 898 4051
rect 1032 4003 1034 4051
rect 1168 4003 1170 4051
rect 1304 4003 1306 4051
rect 1440 4003 1442 4051
rect 1576 4003 1578 4051
rect 1934 4050 1940 4051
rect 1936 4003 1938 4050
rect 1976 4021 1978 4081
rect 1974 4020 1980 4021
rect 2292 4020 2294 4081
rect 2428 4020 2430 4081
rect 2564 4020 2566 4081
rect 2700 4020 2702 4081
rect 2836 4020 2838 4081
rect 3800 4021 3802 4081
rect 3840 4055 3842 4115
rect 3860 4055 3862 4116
rect 4388 4055 4390 4116
rect 4948 4055 4950 4116
rect 5516 4055 5518 4116
rect 5662 4115 5668 4116
rect 5664 4055 5666 4115
rect 3839 4054 3843 4055
rect 3839 4049 3843 4050
rect 3859 4054 3863 4055
rect 3859 4049 3863 4050
rect 4003 4054 4007 4055
rect 4003 4049 4007 4050
rect 4171 4054 4175 4055
rect 4171 4049 4175 4050
rect 4339 4054 4343 4055
rect 4339 4049 4343 4050
rect 4387 4054 4391 4055
rect 4387 4049 4391 4050
rect 4499 4054 4503 4055
rect 4499 4049 4503 4050
rect 4651 4054 4655 4055
rect 4651 4049 4655 4050
rect 4803 4054 4807 4055
rect 4803 4049 4807 4050
rect 4947 4054 4951 4055
rect 4947 4049 4951 4050
rect 5091 4054 5095 4055
rect 5091 4049 5095 4050
rect 5235 4054 5239 4055
rect 5235 4049 5239 4050
rect 5379 4054 5383 4055
rect 5379 4049 5383 4050
rect 5515 4054 5519 4055
rect 5515 4049 5519 4050
rect 5663 4054 5667 4055
rect 5663 4049 5667 4050
rect 3798 4020 3804 4021
rect 1974 4016 1975 4020
rect 1979 4016 1980 4020
rect 1974 4015 1980 4016
rect 2290 4019 2296 4020
rect 2290 4015 2291 4019
rect 2295 4015 2296 4019
rect 2290 4014 2296 4015
rect 2426 4019 2432 4020
rect 2426 4015 2427 4019
rect 2431 4015 2432 4019
rect 2426 4014 2432 4015
rect 2562 4019 2568 4020
rect 2562 4015 2563 4019
rect 2567 4015 2568 4019
rect 2562 4014 2568 4015
rect 2698 4019 2704 4020
rect 2698 4015 2699 4019
rect 2703 4015 2704 4019
rect 2698 4014 2704 4015
rect 2834 4019 2840 4020
rect 2834 4015 2835 4019
rect 2839 4015 2840 4019
rect 3798 4016 3799 4020
rect 3803 4016 3804 4020
rect 3798 4015 3804 4016
rect 2834 4014 2840 4015
rect 2318 4004 2324 4005
rect 1974 4003 1980 4004
rect 111 4002 115 4003
rect 111 3997 115 3998
rect 511 4002 515 4003
rect 511 3997 515 3998
rect 663 4002 667 4003
rect 663 3997 667 3998
rect 759 4002 763 4003
rect 759 3997 763 3998
rect 823 4002 827 4003
rect 823 3997 827 3998
rect 895 4002 899 4003
rect 895 3997 899 3998
rect 983 4002 987 4003
rect 983 3997 987 3998
rect 1031 4002 1035 4003
rect 1031 3997 1035 3998
rect 1151 4002 1155 4003
rect 1151 3997 1155 3998
rect 1167 4002 1171 4003
rect 1167 3997 1171 3998
rect 1303 4002 1307 4003
rect 1303 3997 1307 3998
rect 1319 4002 1323 4003
rect 1319 3997 1323 3998
rect 1439 4002 1443 4003
rect 1439 3997 1443 3998
rect 1575 4002 1579 4003
rect 1575 3997 1579 3998
rect 1935 4002 1939 4003
rect 1974 3999 1975 4003
rect 1979 3999 1980 4003
rect 2318 4000 2319 4004
rect 2323 4000 2324 4004
rect 2318 3999 2324 4000
rect 2454 4004 2460 4005
rect 2454 4000 2455 4004
rect 2459 4000 2460 4004
rect 2454 3999 2460 4000
rect 2590 4004 2596 4005
rect 2590 4000 2591 4004
rect 2595 4000 2596 4004
rect 2590 3999 2596 4000
rect 2726 4004 2732 4005
rect 2726 4000 2727 4004
rect 2731 4000 2732 4004
rect 2726 3999 2732 4000
rect 2862 4004 2868 4005
rect 2862 4000 2863 4004
rect 2867 4000 2868 4004
rect 2862 3999 2868 4000
rect 3798 4003 3804 4004
rect 3798 3999 3799 4003
rect 3803 3999 3804 4003
rect 1974 3998 1980 3999
rect 1935 3997 1939 3998
rect 112 3974 114 3997
rect 110 3973 116 3974
rect 512 3973 514 3997
rect 664 3973 666 3997
rect 824 3973 826 3997
rect 984 3973 986 3997
rect 1152 3973 1154 3997
rect 1320 3973 1322 3997
rect 1936 3974 1938 3997
rect 1934 3973 1940 3974
rect 110 3969 111 3973
rect 115 3969 116 3973
rect 110 3968 116 3969
rect 510 3972 516 3973
rect 510 3968 511 3972
rect 515 3968 516 3972
rect 510 3967 516 3968
rect 662 3972 668 3973
rect 662 3968 663 3972
rect 667 3968 668 3972
rect 662 3967 668 3968
rect 822 3972 828 3973
rect 822 3968 823 3972
rect 827 3968 828 3972
rect 822 3967 828 3968
rect 982 3972 988 3973
rect 982 3968 983 3972
rect 987 3968 988 3972
rect 982 3967 988 3968
rect 1150 3972 1156 3973
rect 1150 3968 1151 3972
rect 1155 3968 1156 3972
rect 1150 3967 1156 3968
rect 1318 3972 1324 3973
rect 1318 3968 1319 3972
rect 1323 3968 1324 3972
rect 1934 3969 1935 3973
rect 1939 3969 1940 3973
rect 1976 3971 1978 3998
rect 2320 3971 2322 3999
rect 2456 3971 2458 3999
rect 2592 3971 2594 3999
rect 2728 3971 2730 3999
rect 2864 3971 2866 3999
rect 3798 3998 3804 3999
rect 3800 3971 3802 3998
rect 3840 3989 3842 4049
rect 3838 3988 3844 3989
rect 3860 3988 3862 4049
rect 4004 3988 4006 4049
rect 4172 3988 4174 4049
rect 4340 3988 4342 4049
rect 4500 3988 4502 4049
rect 4652 3988 4654 4049
rect 4804 3988 4806 4049
rect 4948 3988 4950 4049
rect 5092 3988 5094 4049
rect 5236 3988 5238 4049
rect 5380 3988 5382 4049
rect 5516 3988 5518 4049
rect 5664 3989 5666 4049
rect 5662 3988 5668 3989
rect 3838 3984 3839 3988
rect 3843 3984 3844 3988
rect 3838 3983 3844 3984
rect 3858 3987 3864 3988
rect 3858 3983 3859 3987
rect 3863 3983 3864 3987
rect 3858 3982 3864 3983
rect 4002 3987 4008 3988
rect 4002 3983 4003 3987
rect 4007 3983 4008 3987
rect 4002 3982 4008 3983
rect 4170 3987 4176 3988
rect 4170 3983 4171 3987
rect 4175 3983 4176 3987
rect 4170 3982 4176 3983
rect 4338 3987 4344 3988
rect 4338 3983 4339 3987
rect 4343 3983 4344 3987
rect 4338 3982 4344 3983
rect 4498 3987 4504 3988
rect 4498 3983 4499 3987
rect 4503 3983 4504 3987
rect 4498 3982 4504 3983
rect 4650 3987 4656 3988
rect 4650 3983 4651 3987
rect 4655 3983 4656 3987
rect 4650 3982 4656 3983
rect 4802 3987 4808 3988
rect 4802 3983 4803 3987
rect 4807 3983 4808 3987
rect 4802 3982 4808 3983
rect 4946 3987 4952 3988
rect 4946 3983 4947 3987
rect 4951 3983 4952 3987
rect 4946 3982 4952 3983
rect 5090 3987 5096 3988
rect 5090 3983 5091 3987
rect 5095 3983 5096 3987
rect 5090 3982 5096 3983
rect 5234 3987 5240 3988
rect 5234 3983 5235 3987
rect 5239 3983 5240 3987
rect 5234 3982 5240 3983
rect 5378 3987 5384 3988
rect 5378 3983 5379 3987
rect 5383 3983 5384 3987
rect 5378 3982 5384 3983
rect 5514 3987 5520 3988
rect 5514 3983 5515 3987
rect 5519 3983 5520 3987
rect 5662 3984 5663 3988
rect 5667 3984 5668 3988
rect 5662 3983 5668 3984
rect 5514 3982 5520 3983
rect 3886 3972 3892 3973
rect 3838 3971 3844 3972
rect 1934 3968 1940 3969
rect 1975 3970 1979 3971
rect 1318 3967 1324 3968
rect 1975 3965 1979 3966
rect 2119 3970 2123 3971
rect 2119 3965 2123 3966
rect 2319 3970 2323 3971
rect 2319 3965 2323 3966
rect 2327 3970 2331 3971
rect 2327 3965 2331 3966
rect 2455 3970 2459 3971
rect 2455 3965 2459 3966
rect 2535 3970 2539 3971
rect 2535 3965 2539 3966
rect 2591 3970 2595 3971
rect 2591 3965 2595 3966
rect 2727 3970 2731 3971
rect 2727 3965 2731 3966
rect 2743 3970 2747 3971
rect 2743 3965 2747 3966
rect 2863 3970 2867 3971
rect 2863 3965 2867 3966
rect 2943 3970 2947 3971
rect 2943 3965 2947 3966
rect 3135 3970 3139 3971
rect 3135 3965 3139 3966
rect 3319 3970 3323 3971
rect 3319 3965 3323 3966
rect 3511 3970 3515 3971
rect 3511 3965 3515 3966
rect 3679 3970 3683 3971
rect 3679 3965 3683 3966
rect 3799 3970 3803 3971
rect 3838 3967 3839 3971
rect 3843 3967 3844 3971
rect 3886 3968 3887 3972
rect 3891 3968 3892 3972
rect 3886 3967 3892 3968
rect 4030 3972 4036 3973
rect 4030 3968 4031 3972
rect 4035 3968 4036 3972
rect 4030 3967 4036 3968
rect 4198 3972 4204 3973
rect 4198 3968 4199 3972
rect 4203 3968 4204 3972
rect 4198 3967 4204 3968
rect 4366 3972 4372 3973
rect 4366 3968 4367 3972
rect 4371 3968 4372 3972
rect 4366 3967 4372 3968
rect 4526 3972 4532 3973
rect 4526 3968 4527 3972
rect 4531 3968 4532 3972
rect 4526 3967 4532 3968
rect 4678 3972 4684 3973
rect 4678 3968 4679 3972
rect 4683 3968 4684 3972
rect 4678 3967 4684 3968
rect 4830 3972 4836 3973
rect 4830 3968 4831 3972
rect 4835 3968 4836 3972
rect 4830 3967 4836 3968
rect 4974 3972 4980 3973
rect 4974 3968 4975 3972
rect 4979 3968 4980 3972
rect 4974 3967 4980 3968
rect 5118 3972 5124 3973
rect 5118 3968 5119 3972
rect 5123 3968 5124 3972
rect 5118 3967 5124 3968
rect 5262 3972 5268 3973
rect 5262 3968 5263 3972
rect 5267 3968 5268 3972
rect 5262 3967 5268 3968
rect 5406 3972 5412 3973
rect 5406 3968 5407 3972
rect 5411 3968 5412 3972
rect 5406 3967 5412 3968
rect 5542 3972 5548 3973
rect 5542 3968 5543 3972
rect 5547 3968 5548 3972
rect 5542 3967 5548 3968
rect 5662 3971 5668 3972
rect 5662 3967 5663 3971
rect 5667 3967 5668 3971
rect 3838 3966 3844 3967
rect 3799 3965 3803 3966
rect 482 3957 488 3958
rect 110 3956 116 3957
rect 110 3952 111 3956
rect 115 3952 116 3956
rect 482 3953 483 3957
rect 487 3953 488 3957
rect 482 3952 488 3953
rect 634 3957 640 3958
rect 634 3953 635 3957
rect 639 3953 640 3957
rect 634 3952 640 3953
rect 794 3957 800 3958
rect 794 3953 795 3957
rect 799 3953 800 3957
rect 794 3952 800 3953
rect 954 3957 960 3958
rect 954 3953 955 3957
rect 959 3953 960 3957
rect 954 3952 960 3953
rect 1122 3957 1128 3958
rect 1122 3953 1123 3957
rect 1127 3953 1128 3957
rect 1122 3952 1128 3953
rect 1290 3957 1296 3958
rect 1290 3953 1291 3957
rect 1295 3953 1296 3957
rect 1290 3952 1296 3953
rect 1934 3956 1940 3957
rect 1934 3952 1935 3956
rect 1939 3952 1940 3956
rect 110 3951 116 3952
rect 112 3863 114 3951
rect 484 3863 486 3952
rect 636 3863 638 3952
rect 796 3863 798 3952
rect 956 3863 958 3952
rect 1124 3863 1126 3952
rect 1292 3863 1294 3952
rect 1934 3951 1940 3952
rect 1936 3863 1938 3951
rect 1976 3942 1978 3965
rect 1974 3941 1980 3942
rect 2120 3941 2122 3965
rect 2328 3941 2330 3965
rect 2536 3941 2538 3965
rect 2744 3941 2746 3965
rect 2944 3941 2946 3965
rect 3136 3941 3138 3965
rect 3320 3941 3322 3965
rect 3512 3941 3514 3965
rect 3680 3941 3682 3965
rect 3800 3942 3802 3965
rect 3798 3941 3804 3942
rect 1974 3937 1975 3941
rect 1979 3937 1980 3941
rect 1974 3936 1980 3937
rect 2118 3940 2124 3941
rect 2118 3936 2119 3940
rect 2123 3936 2124 3940
rect 2118 3935 2124 3936
rect 2326 3940 2332 3941
rect 2326 3936 2327 3940
rect 2331 3936 2332 3940
rect 2326 3935 2332 3936
rect 2534 3940 2540 3941
rect 2534 3936 2535 3940
rect 2539 3936 2540 3940
rect 2534 3935 2540 3936
rect 2742 3940 2748 3941
rect 2742 3936 2743 3940
rect 2747 3936 2748 3940
rect 2742 3935 2748 3936
rect 2942 3940 2948 3941
rect 2942 3936 2943 3940
rect 2947 3936 2948 3940
rect 2942 3935 2948 3936
rect 3134 3940 3140 3941
rect 3134 3936 3135 3940
rect 3139 3936 3140 3940
rect 3134 3935 3140 3936
rect 3318 3940 3324 3941
rect 3318 3936 3319 3940
rect 3323 3936 3324 3940
rect 3318 3935 3324 3936
rect 3510 3940 3516 3941
rect 3510 3936 3511 3940
rect 3515 3936 3516 3940
rect 3510 3935 3516 3936
rect 3678 3940 3684 3941
rect 3678 3936 3679 3940
rect 3683 3936 3684 3940
rect 3798 3937 3799 3941
rect 3803 3937 3804 3941
rect 3798 3936 3804 3937
rect 3678 3935 3684 3936
rect 2090 3925 2096 3926
rect 1974 3924 1980 3925
rect 1974 3920 1975 3924
rect 1979 3920 1980 3924
rect 2090 3921 2091 3925
rect 2095 3921 2096 3925
rect 2090 3920 2096 3921
rect 2298 3925 2304 3926
rect 2298 3921 2299 3925
rect 2303 3921 2304 3925
rect 2298 3920 2304 3921
rect 2506 3925 2512 3926
rect 2506 3921 2507 3925
rect 2511 3921 2512 3925
rect 2506 3920 2512 3921
rect 2714 3925 2720 3926
rect 2714 3921 2715 3925
rect 2719 3921 2720 3925
rect 2714 3920 2720 3921
rect 2914 3925 2920 3926
rect 2914 3921 2915 3925
rect 2919 3921 2920 3925
rect 2914 3920 2920 3921
rect 3106 3925 3112 3926
rect 3106 3921 3107 3925
rect 3111 3921 3112 3925
rect 3106 3920 3112 3921
rect 3290 3925 3296 3926
rect 3290 3921 3291 3925
rect 3295 3921 3296 3925
rect 3290 3920 3296 3921
rect 3482 3925 3488 3926
rect 3482 3921 3483 3925
rect 3487 3921 3488 3925
rect 3482 3920 3488 3921
rect 3650 3925 3656 3926
rect 3650 3921 3651 3925
rect 3655 3921 3656 3925
rect 3650 3920 3656 3921
rect 3798 3924 3804 3925
rect 3798 3920 3799 3924
rect 3803 3920 3804 3924
rect 1974 3919 1980 3920
rect 111 3862 115 3863
rect 111 3857 115 3858
rect 131 3862 135 3863
rect 131 3857 135 3858
rect 307 3862 311 3863
rect 307 3857 311 3858
rect 483 3862 487 3863
rect 483 3857 487 3858
rect 515 3862 519 3863
rect 515 3857 519 3858
rect 635 3862 639 3863
rect 635 3857 639 3858
rect 723 3862 727 3863
rect 723 3857 727 3858
rect 795 3862 799 3863
rect 795 3857 799 3858
rect 939 3862 943 3863
rect 939 3857 943 3858
rect 955 3862 959 3863
rect 955 3857 959 3858
rect 1123 3862 1127 3863
rect 1123 3857 1127 3858
rect 1163 3862 1167 3863
rect 1163 3857 1167 3858
rect 1291 3862 1295 3863
rect 1291 3857 1295 3858
rect 1935 3862 1939 3863
rect 1935 3857 1939 3858
rect 112 3797 114 3857
rect 110 3796 116 3797
rect 132 3796 134 3857
rect 308 3796 310 3857
rect 516 3796 518 3857
rect 724 3796 726 3857
rect 940 3796 942 3857
rect 1164 3796 1166 3857
rect 1936 3797 1938 3857
rect 1976 3847 1978 3919
rect 2092 3847 2094 3920
rect 2300 3847 2302 3920
rect 2508 3847 2510 3920
rect 2716 3847 2718 3920
rect 2916 3847 2918 3920
rect 3108 3847 3110 3920
rect 3292 3847 3294 3920
rect 3484 3847 3486 3920
rect 3652 3847 3654 3920
rect 3798 3919 3804 3920
rect 3840 3919 3842 3966
rect 3888 3919 3890 3967
rect 4032 3919 4034 3967
rect 4200 3919 4202 3967
rect 4368 3919 4370 3967
rect 4528 3919 4530 3967
rect 4680 3919 4682 3967
rect 4832 3919 4834 3967
rect 4976 3919 4978 3967
rect 5120 3919 5122 3967
rect 5264 3919 5266 3967
rect 5408 3919 5410 3967
rect 5544 3919 5546 3967
rect 5662 3966 5668 3967
rect 5664 3919 5666 3966
rect 3800 3847 3802 3919
rect 3839 3918 3843 3919
rect 3839 3913 3843 3914
rect 3887 3918 3891 3919
rect 3887 3913 3891 3914
rect 4031 3918 4035 3919
rect 4031 3913 4035 3914
rect 4199 3918 4203 3919
rect 4199 3913 4203 3914
rect 4367 3918 4371 3919
rect 4367 3913 4371 3914
rect 4383 3918 4387 3919
rect 4383 3913 4387 3914
rect 4527 3918 4531 3919
rect 4527 3913 4531 3914
rect 4599 3918 4603 3919
rect 4599 3913 4603 3914
rect 4679 3918 4683 3919
rect 4679 3913 4683 3914
rect 4823 3918 4827 3919
rect 4823 3913 4827 3914
rect 4831 3918 4835 3919
rect 4831 3913 4835 3914
rect 4975 3918 4979 3919
rect 4975 3913 4979 3914
rect 5063 3918 5067 3919
rect 5063 3913 5067 3914
rect 5119 3918 5123 3919
rect 5119 3913 5123 3914
rect 5263 3918 5267 3919
rect 5263 3913 5267 3914
rect 5311 3918 5315 3919
rect 5311 3913 5315 3914
rect 5407 3918 5411 3919
rect 5407 3913 5411 3914
rect 5543 3918 5547 3919
rect 5543 3913 5547 3914
rect 5663 3918 5667 3919
rect 5663 3913 5667 3914
rect 3840 3890 3842 3913
rect 3838 3889 3844 3890
rect 4384 3889 4386 3913
rect 4600 3889 4602 3913
rect 4824 3889 4826 3913
rect 5064 3889 5066 3913
rect 5312 3889 5314 3913
rect 5544 3889 5546 3913
rect 5664 3890 5666 3913
rect 5662 3889 5668 3890
rect 3838 3885 3839 3889
rect 3843 3885 3844 3889
rect 3838 3884 3844 3885
rect 4382 3888 4388 3889
rect 4382 3884 4383 3888
rect 4387 3884 4388 3888
rect 4382 3883 4388 3884
rect 4598 3888 4604 3889
rect 4598 3884 4599 3888
rect 4603 3884 4604 3888
rect 4598 3883 4604 3884
rect 4822 3888 4828 3889
rect 4822 3884 4823 3888
rect 4827 3884 4828 3888
rect 4822 3883 4828 3884
rect 5062 3888 5068 3889
rect 5062 3884 5063 3888
rect 5067 3884 5068 3888
rect 5062 3883 5068 3884
rect 5310 3888 5316 3889
rect 5310 3884 5311 3888
rect 5315 3884 5316 3888
rect 5310 3883 5316 3884
rect 5542 3888 5548 3889
rect 5542 3884 5543 3888
rect 5547 3884 5548 3888
rect 5662 3885 5663 3889
rect 5667 3885 5668 3889
rect 5662 3884 5668 3885
rect 5542 3883 5548 3884
rect 4354 3873 4360 3874
rect 3838 3872 3844 3873
rect 3838 3868 3839 3872
rect 3843 3868 3844 3872
rect 4354 3869 4355 3873
rect 4359 3869 4360 3873
rect 4354 3868 4360 3869
rect 4570 3873 4576 3874
rect 4570 3869 4571 3873
rect 4575 3869 4576 3873
rect 4570 3868 4576 3869
rect 4794 3873 4800 3874
rect 4794 3869 4795 3873
rect 4799 3869 4800 3873
rect 4794 3868 4800 3869
rect 5034 3873 5040 3874
rect 5034 3869 5035 3873
rect 5039 3869 5040 3873
rect 5034 3868 5040 3869
rect 5282 3873 5288 3874
rect 5282 3869 5283 3873
rect 5287 3869 5288 3873
rect 5282 3868 5288 3869
rect 5514 3873 5520 3874
rect 5514 3869 5515 3873
rect 5519 3869 5520 3873
rect 5514 3868 5520 3869
rect 5662 3872 5668 3873
rect 5662 3868 5663 3872
rect 5667 3868 5668 3872
rect 3838 3867 3844 3868
rect 1975 3846 1979 3847
rect 1975 3841 1979 3842
rect 2091 3846 2095 3847
rect 2091 3841 2095 3842
rect 2139 3846 2143 3847
rect 2139 3841 2143 3842
rect 2299 3846 2303 3847
rect 2299 3841 2303 3842
rect 2371 3846 2375 3847
rect 2371 3841 2375 3842
rect 2507 3846 2511 3847
rect 2507 3841 2511 3842
rect 2587 3846 2591 3847
rect 2587 3841 2591 3842
rect 2715 3846 2719 3847
rect 2715 3841 2719 3842
rect 2795 3846 2799 3847
rect 2795 3841 2799 3842
rect 2915 3846 2919 3847
rect 2915 3841 2919 3842
rect 2995 3846 2999 3847
rect 2995 3841 2999 3842
rect 3107 3846 3111 3847
rect 3107 3841 3111 3842
rect 3195 3846 3199 3847
rect 3195 3841 3199 3842
rect 3291 3846 3295 3847
rect 3291 3841 3295 3842
rect 3403 3846 3407 3847
rect 3403 3841 3407 3842
rect 3483 3846 3487 3847
rect 3483 3841 3487 3842
rect 3651 3846 3655 3847
rect 3651 3841 3655 3842
rect 3799 3846 3803 3847
rect 3799 3841 3803 3842
rect 1934 3796 1940 3797
rect 110 3792 111 3796
rect 115 3792 116 3796
rect 110 3791 116 3792
rect 130 3795 136 3796
rect 130 3791 131 3795
rect 135 3791 136 3795
rect 130 3790 136 3791
rect 306 3795 312 3796
rect 306 3791 307 3795
rect 311 3791 312 3795
rect 306 3790 312 3791
rect 514 3795 520 3796
rect 514 3791 515 3795
rect 519 3791 520 3795
rect 514 3790 520 3791
rect 722 3795 728 3796
rect 722 3791 723 3795
rect 727 3791 728 3795
rect 722 3790 728 3791
rect 938 3795 944 3796
rect 938 3791 939 3795
rect 943 3791 944 3795
rect 938 3790 944 3791
rect 1162 3795 1168 3796
rect 1162 3791 1163 3795
rect 1167 3791 1168 3795
rect 1934 3792 1935 3796
rect 1939 3792 1940 3796
rect 1934 3791 1940 3792
rect 1162 3790 1168 3791
rect 1976 3781 1978 3841
rect 158 3780 164 3781
rect 110 3779 116 3780
rect 110 3775 111 3779
rect 115 3775 116 3779
rect 158 3776 159 3780
rect 163 3776 164 3780
rect 158 3775 164 3776
rect 334 3780 340 3781
rect 334 3776 335 3780
rect 339 3776 340 3780
rect 334 3775 340 3776
rect 542 3780 548 3781
rect 542 3776 543 3780
rect 547 3776 548 3780
rect 542 3775 548 3776
rect 750 3780 756 3781
rect 750 3776 751 3780
rect 755 3776 756 3780
rect 750 3775 756 3776
rect 966 3780 972 3781
rect 966 3776 967 3780
rect 971 3776 972 3780
rect 966 3775 972 3776
rect 1190 3780 1196 3781
rect 1974 3780 1980 3781
rect 2140 3780 2142 3841
rect 2372 3780 2374 3841
rect 2588 3780 2590 3841
rect 2796 3780 2798 3841
rect 2996 3780 2998 3841
rect 3196 3780 3198 3841
rect 3404 3780 3406 3841
rect 3800 3781 3802 3841
rect 3840 3791 3842 3867
rect 4356 3791 4358 3868
rect 4572 3791 4574 3868
rect 4796 3791 4798 3868
rect 5036 3791 5038 3868
rect 5284 3791 5286 3868
rect 5516 3791 5518 3868
rect 5662 3867 5668 3868
rect 5664 3791 5666 3867
rect 3839 3790 3843 3791
rect 3839 3785 3843 3786
rect 3995 3790 3999 3791
rect 3995 3785 3999 3786
rect 4203 3790 4207 3791
rect 4203 3785 4207 3786
rect 4355 3790 4359 3791
rect 4355 3785 4359 3786
rect 4435 3790 4439 3791
rect 4435 3785 4439 3786
rect 4571 3790 4575 3791
rect 4571 3785 4575 3786
rect 4691 3790 4695 3791
rect 4691 3785 4695 3786
rect 4795 3790 4799 3791
rect 4795 3785 4799 3786
rect 4963 3790 4967 3791
rect 4963 3785 4967 3786
rect 5035 3790 5039 3791
rect 5035 3785 5039 3786
rect 5251 3790 5255 3791
rect 5251 3785 5255 3786
rect 5283 3790 5287 3791
rect 5283 3785 5287 3786
rect 5515 3790 5519 3791
rect 5515 3785 5519 3786
rect 5663 3790 5667 3791
rect 5663 3785 5667 3786
rect 3798 3780 3804 3781
rect 1190 3776 1191 3780
rect 1195 3776 1196 3780
rect 1190 3775 1196 3776
rect 1934 3779 1940 3780
rect 1934 3775 1935 3779
rect 1939 3775 1940 3779
rect 1974 3776 1975 3780
rect 1979 3776 1980 3780
rect 1974 3775 1980 3776
rect 2138 3779 2144 3780
rect 2138 3775 2139 3779
rect 2143 3775 2144 3779
rect 110 3774 116 3775
rect 112 3751 114 3774
rect 160 3751 162 3775
rect 336 3751 338 3775
rect 544 3751 546 3775
rect 752 3751 754 3775
rect 968 3751 970 3775
rect 1192 3751 1194 3775
rect 1934 3774 1940 3775
rect 2138 3774 2144 3775
rect 2370 3779 2376 3780
rect 2370 3775 2371 3779
rect 2375 3775 2376 3779
rect 2370 3774 2376 3775
rect 2586 3779 2592 3780
rect 2586 3775 2587 3779
rect 2591 3775 2592 3779
rect 2586 3774 2592 3775
rect 2794 3779 2800 3780
rect 2794 3775 2795 3779
rect 2799 3775 2800 3779
rect 2794 3774 2800 3775
rect 2994 3779 3000 3780
rect 2994 3775 2995 3779
rect 2999 3775 3000 3779
rect 2994 3774 3000 3775
rect 3194 3779 3200 3780
rect 3194 3775 3195 3779
rect 3199 3775 3200 3779
rect 3194 3774 3200 3775
rect 3402 3779 3408 3780
rect 3402 3775 3403 3779
rect 3407 3775 3408 3779
rect 3798 3776 3799 3780
rect 3803 3776 3804 3780
rect 3798 3775 3804 3776
rect 3402 3774 3408 3775
rect 1936 3751 1938 3774
rect 2166 3764 2172 3765
rect 1974 3763 1980 3764
rect 1974 3759 1975 3763
rect 1979 3759 1980 3763
rect 2166 3760 2167 3764
rect 2171 3760 2172 3764
rect 2166 3759 2172 3760
rect 2398 3764 2404 3765
rect 2398 3760 2399 3764
rect 2403 3760 2404 3764
rect 2398 3759 2404 3760
rect 2614 3764 2620 3765
rect 2614 3760 2615 3764
rect 2619 3760 2620 3764
rect 2614 3759 2620 3760
rect 2822 3764 2828 3765
rect 2822 3760 2823 3764
rect 2827 3760 2828 3764
rect 2822 3759 2828 3760
rect 3022 3764 3028 3765
rect 3022 3760 3023 3764
rect 3027 3760 3028 3764
rect 3022 3759 3028 3760
rect 3222 3764 3228 3765
rect 3222 3760 3223 3764
rect 3227 3760 3228 3764
rect 3222 3759 3228 3760
rect 3430 3764 3436 3765
rect 3430 3760 3431 3764
rect 3435 3760 3436 3764
rect 3430 3759 3436 3760
rect 3798 3763 3804 3764
rect 3798 3759 3799 3763
rect 3803 3759 3804 3763
rect 1974 3758 1980 3759
rect 111 3750 115 3751
rect 111 3745 115 3746
rect 159 3750 163 3751
rect 159 3745 163 3746
rect 335 3750 339 3751
rect 335 3745 339 3746
rect 527 3750 531 3751
rect 527 3745 531 3746
rect 543 3750 547 3751
rect 543 3745 547 3746
rect 711 3750 715 3751
rect 711 3745 715 3746
rect 751 3750 755 3751
rect 751 3745 755 3746
rect 887 3750 891 3751
rect 887 3745 891 3746
rect 967 3750 971 3751
rect 967 3745 971 3746
rect 1055 3750 1059 3751
rect 1055 3745 1059 3746
rect 1191 3750 1195 3751
rect 1191 3745 1195 3746
rect 1215 3750 1219 3751
rect 1215 3745 1219 3746
rect 1367 3750 1371 3751
rect 1367 3745 1371 3746
rect 1519 3750 1523 3751
rect 1519 3745 1523 3746
rect 1679 3750 1683 3751
rect 1679 3745 1683 3746
rect 1815 3750 1819 3751
rect 1815 3745 1819 3746
rect 1935 3750 1939 3751
rect 1935 3745 1939 3746
rect 112 3722 114 3745
rect 110 3721 116 3722
rect 160 3721 162 3745
rect 336 3721 338 3745
rect 528 3721 530 3745
rect 712 3721 714 3745
rect 888 3721 890 3745
rect 1056 3721 1058 3745
rect 1216 3721 1218 3745
rect 1368 3721 1370 3745
rect 1520 3721 1522 3745
rect 1680 3721 1682 3745
rect 1816 3721 1818 3745
rect 1936 3722 1938 3745
rect 1976 3731 1978 3758
rect 2168 3731 2170 3759
rect 2400 3731 2402 3759
rect 2616 3731 2618 3759
rect 2824 3731 2826 3759
rect 3024 3731 3026 3759
rect 3224 3731 3226 3759
rect 3432 3731 3434 3759
rect 3798 3758 3804 3759
rect 3800 3731 3802 3758
rect 1975 3730 1979 3731
rect 1975 3725 1979 3726
rect 2167 3730 2171 3731
rect 2167 3725 2171 3726
rect 2279 3730 2283 3731
rect 2279 3725 2283 3726
rect 2399 3730 2403 3731
rect 2399 3725 2403 3726
rect 2479 3730 2483 3731
rect 2479 3725 2483 3726
rect 2615 3730 2619 3731
rect 2615 3725 2619 3726
rect 2679 3730 2683 3731
rect 2679 3725 2683 3726
rect 2823 3730 2827 3731
rect 2823 3725 2827 3726
rect 2879 3730 2883 3731
rect 2879 3725 2883 3726
rect 3023 3730 3027 3731
rect 3023 3725 3027 3726
rect 3079 3730 3083 3731
rect 3079 3725 3083 3726
rect 3223 3730 3227 3731
rect 3223 3725 3227 3726
rect 3279 3730 3283 3731
rect 3279 3725 3283 3726
rect 3431 3730 3435 3731
rect 3431 3725 3435 3726
rect 3799 3730 3803 3731
rect 3799 3725 3803 3726
rect 3840 3725 3842 3785
rect 1934 3721 1940 3722
rect 110 3717 111 3721
rect 115 3717 116 3721
rect 110 3716 116 3717
rect 158 3720 164 3721
rect 158 3716 159 3720
rect 163 3716 164 3720
rect 158 3715 164 3716
rect 334 3720 340 3721
rect 334 3716 335 3720
rect 339 3716 340 3720
rect 334 3715 340 3716
rect 526 3720 532 3721
rect 526 3716 527 3720
rect 531 3716 532 3720
rect 526 3715 532 3716
rect 710 3720 716 3721
rect 710 3716 711 3720
rect 715 3716 716 3720
rect 710 3715 716 3716
rect 886 3720 892 3721
rect 886 3716 887 3720
rect 891 3716 892 3720
rect 886 3715 892 3716
rect 1054 3720 1060 3721
rect 1054 3716 1055 3720
rect 1059 3716 1060 3720
rect 1054 3715 1060 3716
rect 1214 3720 1220 3721
rect 1214 3716 1215 3720
rect 1219 3716 1220 3720
rect 1214 3715 1220 3716
rect 1366 3720 1372 3721
rect 1366 3716 1367 3720
rect 1371 3716 1372 3720
rect 1366 3715 1372 3716
rect 1518 3720 1524 3721
rect 1518 3716 1519 3720
rect 1523 3716 1524 3720
rect 1518 3715 1524 3716
rect 1678 3720 1684 3721
rect 1678 3716 1679 3720
rect 1683 3716 1684 3720
rect 1678 3715 1684 3716
rect 1814 3720 1820 3721
rect 1814 3716 1815 3720
rect 1819 3716 1820 3720
rect 1934 3717 1935 3721
rect 1939 3717 1940 3721
rect 1934 3716 1940 3717
rect 1814 3715 1820 3716
rect 130 3705 136 3706
rect 110 3704 116 3705
rect 110 3700 111 3704
rect 115 3700 116 3704
rect 130 3701 131 3705
rect 135 3701 136 3705
rect 130 3700 136 3701
rect 306 3705 312 3706
rect 306 3701 307 3705
rect 311 3701 312 3705
rect 306 3700 312 3701
rect 498 3705 504 3706
rect 498 3701 499 3705
rect 503 3701 504 3705
rect 498 3700 504 3701
rect 682 3705 688 3706
rect 682 3701 683 3705
rect 687 3701 688 3705
rect 682 3700 688 3701
rect 858 3705 864 3706
rect 858 3701 859 3705
rect 863 3701 864 3705
rect 858 3700 864 3701
rect 1026 3705 1032 3706
rect 1026 3701 1027 3705
rect 1031 3701 1032 3705
rect 1026 3700 1032 3701
rect 1186 3705 1192 3706
rect 1186 3701 1187 3705
rect 1191 3701 1192 3705
rect 1186 3700 1192 3701
rect 1338 3705 1344 3706
rect 1338 3701 1339 3705
rect 1343 3701 1344 3705
rect 1338 3700 1344 3701
rect 1490 3705 1496 3706
rect 1490 3701 1491 3705
rect 1495 3701 1496 3705
rect 1490 3700 1496 3701
rect 1650 3705 1656 3706
rect 1650 3701 1651 3705
rect 1655 3701 1656 3705
rect 1650 3700 1656 3701
rect 1786 3705 1792 3706
rect 1786 3701 1787 3705
rect 1791 3701 1792 3705
rect 1786 3700 1792 3701
rect 1934 3704 1940 3705
rect 1934 3700 1935 3704
rect 1939 3700 1940 3704
rect 1976 3702 1978 3725
rect 110 3699 116 3700
rect 112 3627 114 3699
rect 132 3627 134 3700
rect 308 3627 310 3700
rect 500 3627 502 3700
rect 684 3627 686 3700
rect 860 3627 862 3700
rect 1028 3627 1030 3700
rect 1188 3627 1190 3700
rect 1340 3627 1342 3700
rect 1492 3627 1494 3700
rect 1652 3627 1654 3700
rect 1788 3627 1790 3700
rect 1934 3699 1940 3700
rect 1974 3701 1980 3702
rect 2280 3701 2282 3725
rect 2480 3701 2482 3725
rect 2680 3701 2682 3725
rect 2880 3701 2882 3725
rect 3080 3701 3082 3725
rect 3280 3701 3282 3725
rect 3800 3702 3802 3725
rect 3838 3724 3844 3725
rect 3996 3724 3998 3785
rect 4204 3724 4206 3785
rect 4436 3724 4438 3785
rect 4692 3724 4694 3785
rect 4964 3724 4966 3785
rect 5252 3724 5254 3785
rect 5516 3724 5518 3785
rect 5664 3725 5666 3785
rect 5662 3724 5668 3725
rect 3838 3720 3839 3724
rect 3843 3720 3844 3724
rect 3838 3719 3844 3720
rect 3994 3723 4000 3724
rect 3994 3719 3995 3723
rect 3999 3719 4000 3723
rect 3994 3718 4000 3719
rect 4202 3723 4208 3724
rect 4202 3719 4203 3723
rect 4207 3719 4208 3723
rect 4202 3718 4208 3719
rect 4434 3723 4440 3724
rect 4434 3719 4435 3723
rect 4439 3719 4440 3723
rect 4434 3718 4440 3719
rect 4690 3723 4696 3724
rect 4690 3719 4691 3723
rect 4695 3719 4696 3723
rect 4690 3718 4696 3719
rect 4962 3723 4968 3724
rect 4962 3719 4963 3723
rect 4967 3719 4968 3723
rect 4962 3718 4968 3719
rect 5250 3723 5256 3724
rect 5250 3719 5251 3723
rect 5255 3719 5256 3723
rect 5250 3718 5256 3719
rect 5514 3723 5520 3724
rect 5514 3719 5515 3723
rect 5519 3719 5520 3723
rect 5662 3720 5663 3724
rect 5667 3720 5668 3724
rect 5662 3719 5668 3720
rect 5514 3718 5520 3719
rect 4022 3708 4028 3709
rect 3838 3707 3844 3708
rect 3838 3703 3839 3707
rect 3843 3703 3844 3707
rect 4022 3704 4023 3708
rect 4027 3704 4028 3708
rect 4022 3703 4028 3704
rect 4230 3708 4236 3709
rect 4230 3704 4231 3708
rect 4235 3704 4236 3708
rect 4230 3703 4236 3704
rect 4462 3708 4468 3709
rect 4462 3704 4463 3708
rect 4467 3704 4468 3708
rect 4462 3703 4468 3704
rect 4718 3708 4724 3709
rect 4718 3704 4719 3708
rect 4723 3704 4724 3708
rect 4718 3703 4724 3704
rect 4990 3708 4996 3709
rect 4990 3704 4991 3708
rect 4995 3704 4996 3708
rect 4990 3703 4996 3704
rect 5278 3708 5284 3709
rect 5278 3704 5279 3708
rect 5283 3704 5284 3708
rect 5278 3703 5284 3704
rect 5542 3708 5548 3709
rect 5542 3704 5543 3708
rect 5547 3704 5548 3708
rect 5542 3703 5548 3704
rect 5662 3707 5668 3708
rect 5662 3703 5663 3707
rect 5667 3703 5668 3707
rect 3838 3702 3844 3703
rect 3798 3701 3804 3702
rect 1936 3627 1938 3699
rect 1974 3697 1975 3701
rect 1979 3697 1980 3701
rect 1974 3696 1980 3697
rect 2278 3700 2284 3701
rect 2278 3696 2279 3700
rect 2283 3696 2284 3700
rect 2278 3695 2284 3696
rect 2478 3700 2484 3701
rect 2478 3696 2479 3700
rect 2483 3696 2484 3700
rect 2478 3695 2484 3696
rect 2678 3700 2684 3701
rect 2678 3696 2679 3700
rect 2683 3696 2684 3700
rect 2678 3695 2684 3696
rect 2878 3700 2884 3701
rect 2878 3696 2879 3700
rect 2883 3696 2884 3700
rect 2878 3695 2884 3696
rect 3078 3700 3084 3701
rect 3078 3696 3079 3700
rect 3083 3696 3084 3700
rect 3078 3695 3084 3696
rect 3278 3700 3284 3701
rect 3278 3696 3279 3700
rect 3283 3696 3284 3700
rect 3798 3697 3799 3701
rect 3803 3697 3804 3701
rect 3798 3696 3804 3697
rect 3278 3695 3284 3696
rect 2250 3685 2256 3686
rect 1974 3684 1980 3685
rect 1974 3680 1975 3684
rect 1979 3680 1980 3684
rect 2250 3681 2251 3685
rect 2255 3681 2256 3685
rect 2250 3680 2256 3681
rect 2450 3685 2456 3686
rect 2450 3681 2451 3685
rect 2455 3681 2456 3685
rect 2450 3680 2456 3681
rect 2650 3685 2656 3686
rect 2650 3681 2651 3685
rect 2655 3681 2656 3685
rect 2650 3680 2656 3681
rect 2850 3685 2856 3686
rect 2850 3681 2851 3685
rect 2855 3681 2856 3685
rect 2850 3680 2856 3681
rect 3050 3685 3056 3686
rect 3050 3681 3051 3685
rect 3055 3681 3056 3685
rect 3050 3680 3056 3681
rect 3250 3685 3256 3686
rect 3250 3681 3251 3685
rect 3255 3681 3256 3685
rect 3250 3680 3256 3681
rect 3798 3684 3804 3685
rect 3798 3680 3799 3684
rect 3803 3680 3804 3684
rect 1974 3679 1980 3680
rect 111 3626 115 3627
rect 111 3621 115 3622
rect 131 3626 135 3627
rect 131 3621 135 3622
rect 147 3626 151 3627
rect 147 3621 151 3622
rect 307 3626 311 3627
rect 307 3621 311 3622
rect 355 3626 359 3627
rect 355 3621 359 3622
rect 499 3626 503 3627
rect 499 3621 503 3622
rect 571 3626 575 3627
rect 571 3621 575 3622
rect 683 3626 687 3627
rect 683 3621 687 3622
rect 803 3626 807 3627
rect 803 3621 807 3622
rect 859 3626 863 3627
rect 859 3621 863 3622
rect 1027 3626 1031 3627
rect 1027 3621 1031 3622
rect 1043 3626 1047 3627
rect 1043 3621 1047 3622
rect 1187 3626 1191 3627
rect 1187 3621 1191 3622
rect 1291 3626 1295 3627
rect 1291 3621 1295 3622
rect 1339 3626 1343 3627
rect 1339 3621 1343 3622
rect 1491 3626 1495 3627
rect 1491 3621 1495 3622
rect 1547 3626 1551 3627
rect 1547 3621 1551 3622
rect 1651 3626 1655 3627
rect 1651 3621 1655 3622
rect 1787 3626 1791 3627
rect 1787 3621 1791 3622
rect 1935 3626 1939 3627
rect 1935 3621 1939 3622
rect 112 3561 114 3621
rect 110 3560 116 3561
rect 148 3560 150 3621
rect 356 3560 358 3621
rect 572 3560 574 3621
rect 804 3560 806 3621
rect 1044 3560 1046 3621
rect 1292 3560 1294 3621
rect 1548 3560 1550 3621
rect 1788 3560 1790 3621
rect 1936 3561 1938 3621
rect 1976 3607 1978 3679
rect 2252 3607 2254 3680
rect 2452 3607 2454 3680
rect 2652 3607 2654 3680
rect 2852 3607 2854 3680
rect 3052 3607 3054 3680
rect 3252 3607 3254 3680
rect 3798 3679 3804 3680
rect 3800 3607 3802 3679
rect 3840 3651 3842 3702
rect 4024 3651 4026 3703
rect 4232 3651 4234 3703
rect 4464 3651 4466 3703
rect 4720 3651 4722 3703
rect 4992 3651 4994 3703
rect 5280 3651 5282 3703
rect 5544 3651 5546 3703
rect 5662 3702 5668 3703
rect 5664 3651 5666 3702
rect 3839 3650 3843 3651
rect 3839 3645 3843 3646
rect 4023 3650 4027 3651
rect 4023 3645 4027 3646
rect 4215 3650 4219 3651
rect 4215 3645 4219 3646
rect 4231 3650 4235 3651
rect 4231 3645 4235 3646
rect 4399 3650 4403 3651
rect 4399 3645 4403 3646
rect 4463 3650 4467 3651
rect 4463 3645 4467 3646
rect 4607 3650 4611 3651
rect 4607 3645 4611 3646
rect 4719 3650 4723 3651
rect 4719 3645 4723 3646
rect 4831 3650 4835 3651
rect 4831 3645 4835 3646
rect 4991 3650 4995 3651
rect 4991 3645 4995 3646
rect 5071 3650 5075 3651
rect 5071 3645 5075 3646
rect 5279 3650 5283 3651
rect 5279 3645 5283 3646
rect 5319 3650 5323 3651
rect 5319 3645 5323 3646
rect 5543 3650 5547 3651
rect 5543 3645 5547 3646
rect 5663 3650 5667 3651
rect 5663 3645 5667 3646
rect 3840 3622 3842 3645
rect 3838 3621 3844 3622
rect 4216 3621 4218 3645
rect 4400 3621 4402 3645
rect 4608 3621 4610 3645
rect 4832 3621 4834 3645
rect 5072 3621 5074 3645
rect 5320 3621 5322 3645
rect 5544 3621 5546 3645
rect 5664 3622 5666 3645
rect 5662 3621 5668 3622
rect 3838 3617 3839 3621
rect 3843 3617 3844 3621
rect 3838 3616 3844 3617
rect 4214 3620 4220 3621
rect 4214 3616 4215 3620
rect 4219 3616 4220 3620
rect 4214 3615 4220 3616
rect 4398 3620 4404 3621
rect 4398 3616 4399 3620
rect 4403 3616 4404 3620
rect 4398 3615 4404 3616
rect 4606 3620 4612 3621
rect 4606 3616 4607 3620
rect 4611 3616 4612 3620
rect 4606 3615 4612 3616
rect 4830 3620 4836 3621
rect 4830 3616 4831 3620
rect 4835 3616 4836 3620
rect 4830 3615 4836 3616
rect 5070 3620 5076 3621
rect 5070 3616 5071 3620
rect 5075 3616 5076 3620
rect 5070 3615 5076 3616
rect 5318 3620 5324 3621
rect 5318 3616 5319 3620
rect 5323 3616 5324 3620
rect 5318 3615 5324 3616
rect 5542 3620 5548 3621
rect 5542 3616 5543 3620
rect 5547 3616 5548 3620
rect 5662 3617 5663 3621
rect 5667 3617 5668 3621
rect 5662 3616 5668 3617
rect 5542 3615 5548 3616
rect 1975 3606 1979 3607
rect 1975 3601 1979 3602
rect 1995 3606 1999 3607
rect 1995 3601 1999 3602
rect 2251 3606 2255 3607
rect 2251 3601 2255 3602
rect 2451 3606 2455 3607
rect 2451 3601 2455 3602
rect 2515 3606 2519 3607
rect 2515 3601 2519 3602
rect 2651 3606 2655 3607
rect 2651 3601 2655 3602
rect 2755 3606 2759 3607
rect 2755 3601 2759 3602
rect 2851 3606 2855 3607
rect 2851 3601 2855 3602
rect 2979 3606 2983 3607
rect 2979 3601 2983 3602
rect 3051 3606 3055 3607
rect 3051 3601 3055 3602
rect 3195 3606 3199 3607
rect 3195 3601 3199 3602
rect 3251 3606 3255 3607
rect 3251 3601 3255 3602
rect 3411 3606 3415 3607
rect 3411 3601 3415 3602
rect 3627 3606 3631 3607
rect 3627 3601 3631 3602
rect 3799 3606 3803 3607
rect 4186 3605 4192 3606
rect 3799 3601 3803 3602
rect 3838 3604 3844 3605
rect 1934 3560 1940 3561
rect 110 3556 111 3560
rect 115 3556 116 3560
rect 110 3555 116 3556
rect 146 3559 152 3560
rect 146 3555 147 3559
rect 151 3555 152 3559
rect 146 3554 152 3555
rect 354 3559 360 3560
rect 354 3555 355 3559
rect 359 3555 360 3559
rect 354 3554 360 3555
rect 570 3559 576 3560
rect 570 3555 571 3559
rect 575 3555 576 3559
rect 570 3554 576 3555
rect 802 3559 808 3560
rect 802 3555 803 3559
rect 807 3555 808 3559
rect 802 3554 808 3555
rect 1042 3559 1048 3560
rect 1042 3555 1043 3559
rect 1047 3555 1048 3559
rect 1042 3554 1048 3555
rect 1290 3559 1296 3560
rect 1290 3555 1291 3559
rect 1295 3555 1296 3559
rect 1290 3554 1296 3555
rect 1546 3559 1552 3560
rect 1546 3555 1547 3559
rect 1551 3555 1552 3559
rect 1546 3554 1552 3555
rect 1786 3559 1792 3560
rect 1786 3555 1787 3559
rect 1791 3555 1792 3559
rect 1934 3556 1935 3560
rect 1939 3556 1940 3560
rect 1934 3555 1940 3556
rect 1786 3554 1792 3555
rect 174 3544 180 3545
rect 110 3543 116 3544
rect 110 3539 111 3543
rect 115 3539 116 3543
rect 174 3540 175 3544
rect 179 3540 180 3544
rect 174 3539 180 3540
rect 382 3544 388 3545
rect 382 3540 383 3544
rect 387 3540 388 3544
rect 382 3539 388 3540
rect 598 3544 604 3545
rect 598 3540 599 3544
rect 603 3540 604 3544
rect 598 3539 604 3540
rect 830 3544 836 3545
rect 830 3540 831 3544
rect 835 3540 836 3544
rect 830 3539 836 3540
rect 1070 3544 1076 3545
rect 1070 3540 1071 3544
rect 1075 3540 1076 3544
rect 1070 3539 1076 3540
rect 1318 3544 1324 3545
rect 1318 3540 1319 3544
rect 1323 3540 1324 3544
rect 1318 3539 1324 3540
rect 1574 3544 1580 3545
rect 1574 3540 1575 3544
rect 1579 3540 1580 3544
rect 1574 3539 1580 3540
rect 1814 3544 1820 3545
rect 1814 3540 1815 3544
rect 1819 3540 1820 3544
rect 1814 3539 1820 3540
rect 1934 3543 1940 3544
rect 1934 3539 1935 3543
rect 1939 3539 1940 3543
rect 1976 3541 1978 3601
rect 110 3538 116 3539
rect 112 3491 114 3538
rect 176 3491 178 3539
rect 384 3491 386 3539
rect 600 3491 602 3539
rect 832 3491 834 3539
rect 1072 3491 1074 3539
rect 1320 3491 1322 3539
rect 1576 3491 1578 3539
rect 1816 3491 1818 3539
rect 1934 3538 1940 3539
rect 1974 3540 1980 3541
rect 1996 3540 1998 3601
rect 2252 3540 2254 3601
rect 2516 3540 2518 3601
rect 2756 3540 2758 3601
rect 2980 3540 2982 3601
rect 3196 3540 3198 3601
rect 3412 3540 3414 3601
rect 3628 3540 3630 3601
rect 3800 3541 3802 3601
rect 3838 3600 3839 3604
rect 3843 3600 3844 3604
rect 4186 3601 4187 3605
rect 4191 3601 4192 3605
rect 4186 3600 4192 3601
rect 4370 3605 4376 3606
rect 4370 3601 4371 3605
rect 4375 3601 4376 3605
rect 4370 3600 4376 3601
rect 4578 3605 4584 3606
rect 4578 3601 4579 3605
rect 4583 3601 4584 3605
rect 4578 3600 4584 3601
rect 4802 3605 4808 3606
rect 4802 3601 4803 3605
rect 4807 3601 4808 3605
rect 4802 3600 4808 3601
rect 5042 3605 5048 3606
rect 5042 3601 5043 3605
rect 5047 3601 5048 3605
rect 5042 3600 5048 3601
rect 5290 3605 5296 3606
rect 5290 3601 5291 3605
rect 5295 3601 5296 3605
rect 5290 3600 5296 3601
rect 5514 3605 5520 3606
rect 5514 3601 5515 3605
rect 5519 3601 5520 3605
rect 5514 3600 5520 3601
rect 5662 3604 5668 3605
rect 5662 3600 5663 3604
rect 5667 3600 5668 3604
rect 3838 3599 3844 3600
rect 3798 3540 3804 3541
rect 1936 3491 1938 3538
rect 1974 3536 1975 3540
rect 1979 3536 1980 3540
rect 1974 3535 1980 3536
rect 1994 3539 2000 3540
rect 1994 3535 1995 3539
rect 1999 3535 2000 3539
rect 1994 3534 2000 3535
rect 2250 3539 2256 3540
rect 2250 3535 2251 3539
rect 2255 3535 2256 3539
rect 2250 3534 2256 3535
rect 2514 3539 2520 3540
rect 2514 3535 2515 3539
rect 2519 3535 2520 3539
rect 2514 3534 2520 3535
rect 2754 3539 2760 3540
rect 2754 3535 2755 3539
rect 2759 3535 2760 3539
rect 2754 3534 2760 3535
rect 2978 3539 2984 3540
rect 2978 3535 2979 3539
rect 2983 3535 2984 3539
rect 2978 3534 2984 3535
rect 3194 3539 3200 3540
rect 3194 3535 3195 3539
rect 3199 3535 3200 3539
rect 3194 3534 3200 3535
rect 3410 3539 3416 3540
rect 3410 3535 3411 3539
rect 3415 3535 3416 3539
rect 3410 3534 3416 3535
rect 3626 3539 3632 3540
rect 3626 3535 3627 3539
rect 3631 3535 3632 3539
rect 3798 3536 3799 3540
rect 3803 3536 3804 3540
rect 3798 3535 3804 3536
rect 3626 3534 3632 3535
rect 2022 3524 2028 3525
rect 1974 3523 1980 3524
rect 1974 3519 1975 3523
rect 1979 3519 1980 3523
rect 2022 3520 2023 3524
rect 2027 3520 2028 3524
rect 2022 3519 2028 3520
rect 2278 3524 2284 3525
rect 2278 3520 2279 3524
rect 2283 3520 2284 3524
rect 2278 3519 2284 3520
rect 2542 3524 2548 3525
rect 2542 3520 2543 3524
rect 2547 3520 2548 3524
rect 2542 3519 2548 3520
rect 2782 3524 2788 3525
rect 2782 3520 2783 3524
rect 2787 3520 2788 3524
rect 2782 3519 2788 3520
rect 3006 3524 3012 3525
rect 3006 3520 3007 3524
rect 3011 3520 3012 3524
rect 3006 3519 3012 3520
rect 3222 3524 3228 3525
rect 3222 3520 3223 3524
rect 3227 3520 3228 3524
rect 3222 3519 3228 3520
rect 3438 3524 3444 3525
rect 3438 3520 3439 3524
rect 3443 3520 3444 3524
rect 3438 3519 3444 3520
rect 3654 3524 3660 3525
rect 3654 3520 3655 3524
rect 3659 3520 3660 3524
rect 3654 3519 3660 3520
rect 3798 3523 3804 3524
rect 3798 3519 3799 3523
rect 3803 3519 3804 3523
rect 1974 3518 1980 3519
rect 111 3490 115 3491
rect 111 3485 115 3486
rect 175 3490 179 3491
rect 175 3485 179 3486
rect 303 3490 307 3491
rect 303 3485 307 3486
rect 383 3490 387 3491
rect 383 3485 387 3486
rect 447 3490 451 3491
rect 447 3485 451 3486
rect 599 3490 603 3491
rect 599 3485 603 3486
rect 759 3490 763 3491
rect 759 3485 763 3486
rect 831 3490 835 3491
rect 831 3485 835 3486
rect 935 3490 939 3491
rect 935 3485 939 3486
rect 1071 3490 1075 3491
rect 1071 3485 1075 3486
rect 1111 3490 1115 3491
rect 1111 3485 1115 3486
rect 1295 3490 1299 3491
rect 1295 3485 1299 3486
rect 1319 3490 1323 3491
rect 1319 3485 1323 3486
rect 1487 3490 1491 3491
rect 1487 3485 1491 3486
rect 1575 3490 1579 3491
rect 1575 3485 1579 3486
rect 1815 3490 1819 3491
rect 1815 3485 1819 3486
rect 1935 3490 1939 3491
rect 1976 3487 1978 3518
rect 2024 3487 2026 3519
rect 2280 3487 2282 3519
rect 2544 3487 2546 3519
rect 2784 3487 2786 3519
rect 3008 3487 3010 3519
rect 3224 3487 3226 3519
rect 3440 3487 3442 3519
rect 3656 3487 3658 3519
rect 3798 3518 3804 3519
rect 3800 3487 3802 3518
rect 3840 3515 3842 3599
rect 4188 3515 4190 3600
rect 4372 3515 4374 3600
rect 4580 3515 4582 3600
rect 4804 3515 4806 3600
rect 5044 3515 5046 3600
rect 5292 3515 5294 3600
rect 5516 3515 5518 3600
rect 5662 3599 5668 3600
rect 5664 3515 5666 3599
rect 3839 3514 3843 3515
rect 3839 3509 3843 3510
rect 4187 3514 4191 3515
rect 4187 3509 4191 3510
rect 4371 3514 4375 3515
rect 4371 3509 4375 3510
rect 4531 3514 4535 3515
rect 4531 3509 4535 3510
rect 4579 3514 4583 3515
rect 4579 3509 4583 3510
rect 4683 3514 4687 3515
rect 4683 3509 4687 3510
rect 4803 3514 4807 3515
rect 4803 3509 4807 3510
rect 4843 3514 4847 3515
rect 4843 3509 4847 3510
rect 5003 3514 5007 3515
rect 5003 3509 5007 3510
rect 5043 3514 5047 3515
rect 5043 3509 5047 3510
rect 5171 3514 5175 3515
rect 5171 3509 5175 3510
rect 5291 3514 5295 3515
rect 5291 3509 5295 3510
rect 5347 3514 5351 3515
rect 5347 3509 5351 3510
rect 5515 3514 5519 3515
rect 5515 3509 5519 3510
rect 5663 3514 5667 3515
rect 5663 3509 5667 3510
rect 1935 3485 1939 3486
rect 1975 3486 1979 3487
rect 112 3462 114 3485
rect 110 3461 116 3462
rect 304 3461 306 3485
rect 448 3461 450 3485
rect 600 3461 602 3485
rect 760 3461 762 3485
rect 936 3461 938 3485
rect 1112 3461 1114 3485
rect 1296 3461 1298 3485
rect 1488 3461 1490 3485
rect 1936 3462 1938 3485
rect 1975 3481 1979 3482
rect 2023 3486 2027 3487
rect 2023 3481 2027 3482
rect 2191 3486 2195 3487
rect 2191 3481 2195 3482
rect 2279 3486 2283 3487
rect 2279 3481 2283 3482
rect 2399 3486 2403 3487
rect 2399 3481 2403 3482
rect 2543 3486 2547 3487
rect 2543 3481 2547 3482
rect 2615 3486 2619 3487
rect 2615 3481 2619 3482
rect 2783 3486 2787 3487
rect 2783 3481 2787 3482
rect 2831 3486 2835 3487
rect 2831 3481 2835 3482
rect 3007 3486 3011 3487
rect 3007 3481 3011 3482
rect 3047 3486 3051 3487
rect 3047 3481 3051 3482
rect 3223 3486 3227 3487
rect 3223 3481 3227 3482
rect 3263 3486 3267 3487
rect 3263 3481 3267 3482
rect 3439 3486 3443 3487
rect 3439 3481 3443 3482
rect 3479 3486 3483 3487
rect 3479 3481 3483 3482
rect 3655 3486 3659 3487
rect 3655 3481 3659 3482
rect 3679 3486 3683 3487
rect 3679 3481 3683 3482
rect 3799 3486 3803 3487
rect 3799 3481 3803 3482
rect 1934 3461 1940 3462
rect 110 3457 111 3461
rect 115 3457 116 3461
rect 110 3456 116 3457
rect 302 3460 308 3461
rect 302 3456 303 3460
rect 307 3456 308 3460
rect 302 3455 308 3456
rect 446 3460 452 3461
rect 446 3456 447 3460
rect 451 3456 452 3460
rect 446 3455 452 3456
rect 598 3460 604 3461
rect 598 3456 599 3460
rect 603 3456 604 3460
rect 598 3455 604 3456
rect 758 3460 764 3461
rect 758 3456 759 3460
rect 763 3456 764 3460
rect 758 3455 764 3456
rect 934 3460 940 3461
rect 934 3456 935 3460
rect 939 3456 940 3460
rect 934 3455 940 3456
rect 1110 3460 1116 3461
rect 1110 3456 1111 3460
rect 1115 3456 1116 3460
rect 1110 3455 1116 3456
rect 1294 3460 1300 3461
rect 1294 3456 1295 3460
rect 1299 3456 1300 3460
rect 1294 3455 1300 3456
rect 1486 3460 1492 3461
rect 1486 3456 1487 3460
rect 1491 3456 1492 3460
rect 1934 3457 1935 3461
rect 1939 3457 1940 3461
rect 1976 3458 1978 3481
rect 1934 3456 1940 3457
rect 1974 3457 1980 3458
rect 2024 3457 2026 3481
rect 2192 3457 2194 3481
rect 2400 3457 2402 3481
rect 2616 3457 2618 3481
rect 2832 3457 2834 3481
rect 3048 3457 3050 3481
rect 3264 3457 3266 3481
rect 3480 3457 3482 3481
rect 3680 3457 3682 3481
rect 3800 3458 3802 3481
rect 3798 3457 3804 3458
rect 1486 3455 1492 3456
rect 1974 3453 1975 3457
rect 1979 3453 1980 3457
rect 1974 3452 1980 3453
rect 2022 3456 2028 3457
rect 2022 3452 2023 3456
rect 2027 3452 2028 3456
rect 2022 3451 2028 3452
rect 2190 3456 2196 3457
rect 2190 3452 2191 3456
rect 2195 3452 2196 3456
rect 2190 3451 2196 3452
rect 2398 3456 2404 3457
rect 2398 3452 2399 3456
rect 2403 3452 2404 3456
rect 2398 3451 2404 3452
rect 2614 3456 2620 3457
rect 2614 3452 2615 3456
rect 2619 3452 2620 3456
rect 2614 3451 2620 3452
rect 2830 3456 2836 3457
rect 2830 3452 2831 3456
rect 2835 3452 2836 3456
rect 2830 3451 2836 3452
rect 3046 3456 3052 3457
rect 3046 3452 3047 3456
rect 3051 3452 3052 3456
rect 3046 3451 3052 3452
rect 3262 3456 3268 3457
rect 3262 3452 3263 3456
rect 3267 3452 3268 3456
rect 3262 3451 3268 3452
rect 3478 3456 3484 3457
rect 3478 3452 3479 3456
rect 3483 3452 3484 3456
rect 3478 3451 3484 3452
rect 3678 3456 3684 3457
rect 3678 3452 3679 3456
rect 3683 3452 3684 3456
rect 3798 3453 3799 3457
rect 3803 3453 3804 3457
rect 3798 3452 3804 3453
rect 3678 3451 3684 3452
rect 3840 3449 3842 3509
rect 3838 3448 3844 3449
rect 4532 3448 4534 3509
rect 4684 3448 4686 3509
rect 4844 3448 4846 3509
rect 5004 3448 5006 3509
rect 5172 3448 5174 3509
rect 5348 3448 5350 3509
rect 5516 3448 5518 3509
rect 5664 3449 5666 3509
rect 5662 3448 5668 3449
rect 274 3445 280 3446
rect 110 3444 116 3445
rect 110 3440 111 3444
rect 115 3440 116 3444
rect 274 3441 275 3445
rect 279 3441 280 3445
rect 274 3440 280 3441
rect 418 3445 424 3446
rect 418 3441 419 3445
rect 423 3441 424 3445
rect 418 3440 424 3441
rect 570 3445 576 3446
rect 570 3441 571 3445
rect 575 3441 576 3445
rect 570 3440 576 3441
rect 730 3445 736 3446
rect 730 3441 731 3445
rect 735 3441 736 3445
rect 730 3440 736 3441
rect 906 3445 912 3446
rect 906 3441 907 3445
rect 911 3441 912 3445
rect 906 3440 912 3441
rect 1082 3445 1088 3446
rect 1082 3441 1083 3445
rect 1087 3441 1088 3445
rect 1082 3440 1088 3441
rect 1266 3445 1272 3446
rect 1266 3441 1267 3445
rect 1271 3441 1272 3445
rect 1266 3440 1272 3441
rect 1458 3445 1464 3446
rect 1458 3441 1459 3445
rect 1463 3441 1464 3445
rect 1458 3440 1464 3441
rect 1934 3444 1940 3445
rect 1934 3440 1935 3444
rect 1939 3440 1940 3444
rect 3838 3444 3839 3448
rect 3843 3444 3844 3448
rect 3838 3443 3844 3444
rect 4530 3447 4536 3448
rect 4530 3443 4531 3447
rect 4535 3443 4536 3447
rect 4530 3442 4536 3443
rect 4682 3447 4688 3448
rect 4682 3443 4683 3447
rect 4687 3443 4688 3447
rect 4682 3442 4688 3443
rect 4842 3447 4848 3448
rect 4842 3443 4843 3447
rect 4847 3443 4848 3447
rect 4842 3442 4848 3443
rect 5002 3447 5008 3448
rect 5002 3443 5003 3447
rect 5007 3443 5008 3447
rect 5002 3442 5008 3443
rect 5170 3447 5176 3448
rect 5170 3443 5171 3447
rect 5175 3443 5176 3447
rect 5170 3442 5176 3443
rect 5346 3447 5352 3448
rect 5346 3443 5347 3447
rect 5351 3443 5352 3447
rect 5346 3442 5352 3443
rect 5514 3447 5520 3448
rect 5514 3443 5515 3447
rect 5519 3443 5520 3447
rect 5662 3444 5663 3448
rect 5667 3444 5668 3448
rect 5662 3443 5668 3444
rect 5514 3442 5520 3443
rect 1994 3441 2000 3442
rect 110 3439 116 3440
rect 112 3363 114 3439
rect 276 3363 278 3440
rect 420 3363 422 3440
rect 572 3363 574 3440
rect 732 3363 734 3440
rect 908 3363 910 3440
rect 1084 3363 1086 3440
rect 1268 3363 1270 3440
rect 1460 3363 1462 3440
rect 1934 3439 1940 3440
rect 1974 3440 1980 3441
rect 1936 3363 1938 3439
rect 1974 3436 1975 3440
rect 1979 3436 1980 3440
rect 1994 3437 1995 3441
rect 1999 3437 2000 3441
rect 1994 3436 2000 3437
rect 2162 3441 2168 3442
rect 2162 3437 2163 3441
rect 2167 3437 2168 3441
rect 2162 3436 2168 3437
rect 2370 3441 2376 3442
rect 2370 3437 2371 3441
rect 2375 3437 2376 3441
rect 2370 3436 2376 3437
rect 2586 3441 2592 3442
rect 2586 3437 2587 3441
rect 2591 3437 2592 3441
rect 2586 3436 2592 3437
rect 2802 3441 2808 3442
rect 2802 3437 2803 3441
rect 2807 3437 2808 3441
rect 2802 3436 2808 3437
rect 3018 3441 3024 3442
rect 3018 3437 3019 3441
rect 3023 3437 3024 3441
rect 3018 3436 3024 3437
rect 3234 3441 3240 3442
rect 3234 3437 3235 3441
rect 3239 3437 3240 3441
rect 3234 3436 3240 3437
rect 3450 3441 3456 3442
rect 3450 3437 3451 3441
rect 3455 3437 3456 3441
rect 3450 3436 3456 3437
rect 3650 3441 3656 3442
rect 3650 3437 3651 3441
rect 3655 3437 3656 3441
rect 3650 3436 3656 3437
rect 3798 3440 3804 3441
rect 3798 3436 3799 3440
rect 3803 3436 3804 3440
rect 1974 3435 1980 3436
rect 111 3362 115 3363
rect 111 3357 115 3358
rect 275 3362 279 3363
rect 275 3357 279 3358
rect 419 3362 423 3363
rect 419 3357 423 3358
rect 467 3362 471 3363
rect 467 3357 471 3358
rect 571 3362 575 3363
rect 571 3357 575 3358
rect 667 3362 671 3363
rect 667 3357 671 3358
rect 731 3362 735 3363
rect 731 3357 735 3358
rect 875 3362 879 3363
rect 875 3357 879 3358
rect 907 3362 911 3363
rect 907 3357 911 3358
rect 1083 3362 1087 3363
rect 1083 3357 1087 3358
rect 1091 3362 1095 3363
rect 1091 3357 1095 3358
rect 1267 3362 1271 3363
rect 1267 3357 1271 3358
rect 1315 3362 1319 3363
rect 1315 3357 1319 3358
rect 1459 3362 1463 3363
rect 1459 3357 1463 3358
rect 1935 3362 1939 3363
rect 1935 3357 1939 3358
rect 112 3297 114 3357
rect 110 3296 116 3297
rect 468 3296 470 3357
rect 668 3296 670 3357
rect 876 3296 878 3357
rect 1092 3296 1094 3357
rect 1316 3296 1318 3357
rect 1936 3297 1938 3357
rect 1976 3335 1978 3435
rect 1996 3335 1998 3436
rect 2164 3335 2166 3436
rect 2372 3335 2374 3436
rect 2588 3335 2590 3436
rect 2804 3335 2806 3436
rect 3020 3335 3022 3436
rect 3236 3335 3238 3436
rect 3452 3335 3454 3436
rect 3652 3335 3654 3436
rect 3798 3435 3804 3436
rect 3800 3335 3802 3435
rect 4558 3432 4564 3433
rect 3838 3431 3844 3432
rect 3838 3427 3839 3431
rect 3843 3427 3844 3431
rect 4558 3428 4559 3432
rect 4563 3428 4564 3432
rect 4558 3427 4564 3428
rect 4710 3432 4716 3433
rect 4710 3428 4711 3432
rect 4715 3428 4716 3432
rect 4710 3427 4716 3428
rect 4870 3432 4876 3433
rect 4870 3428 4871 3432
rect 4875 3428 4876 3432
rect 4870 3427 4876 3428
rect 5030 3432 5036 3433
rect 5030 3428 5031 3432
rect 5035 3428 5036 3432
rect 5030 3427 5036 3428
rect 5198 3432 5204 3433
rect 5198 3428 5199 3432
rect 5203 3428 5204 3432
rect 5198 3427 5204 3428
rect 5374 3432 5380 3433
rect 5374 3428 5375 3432
rect 5379 3428 5380 3432
rect 5374 3427 5380 3428
rect 5542 3432 5548 3433
rect 5542 3428 5543 3432
rect 5547 3428 5548 3432
rect 5542 3427 5548 3428
rect 5662 3431 5668 3432
rect 5662 3427 5663 3431
rect 5667 3427 5668 3431
rect 3838 3426 3844 3427
rect 3840 3399 3842 3426
rect 4560 3399 4562 3427
rect 4712 3399 4714 3427
rect 4872 3399 4874 3427
rect 5032 3399 5034 3427
rect 5200 3399 5202 3427
rect 5376 3399 5378 3427
rect 5544 3399 5546 3427
rect 5662 3426 5668 3427
rect 5664 3399 5666 3426
rect 3839 3398 3843 3399
rect 3839 3393 3843 3394
rect 3887 3398 3891 3399
rect 3887 3393 3891 3394
rect 4151 3398 4155 3399
rect 4151 3393 4155 3394
rect 4423 3398 4427 3399
rect 4423 3393 4427 3394
rect 4559 3398 4563 3399
rect 4559 3393 4563 3394
rect 4671 3398 4675 3399
rect 4671 3393 4675 3394
rect 4711 3398 4715 3399
rect 4711 3393 4715 3394
rect 4871 3398 4875 3399
rect 4871 3393 4875 3394
rect 4895 3398 4899 3399
rect 4895 3393 4899 3394
rect 5031 3398 5035 3399
rect 5031 3393 5035 3394
rect 5111 3398 5115 3399
rect 5111 3393 5115 3394
rect 5199 3398 5203 3399
rect 5199 3393 5203 3394
rect 5327 3398 5331 3399
rect 5327 3393 5331 3394
rect 5375 3398 5379 3399
rect 5375 3393 5379 3394
rect 5543 3398 5547 3399
rect 5543 3393 5547 3394
rect 5663 3398 5667 3399
rect 5663 3393 5667 3394
rect 3840 3370 3842 3393
rect 3838 3369 3844 3370
rect 3888 3369 3890 3393
rect 4152 3369 4154 3393
rect 4424 3369 4426 3393
rect 4672 3369 4674 3393
rect 4896 3369 4898 3393
rect 5112 3369 5114 3393
rect 5328 3369 5330 3393
rect 5544 3369 5546 3393
rect 5664 3370 5666 3393
rect 5662 3369 5668 3370
rect 3838 3365 3839 3369
rect 3843 3365 3844 3369
rect 3838 3364 3844 3365
rect 3886 3368 3892 3369
rect 3886 3364 3887 3368
rect 3891 3364 3892 3368
rect 3886 3363 3892 3364
rect 4150 3368 4156 3369
rect 4150 3364 4151 3368
rect 4155 3364 4156 3368
rect 4150 3363 4156 3364
rect 4422 3368 4428 3369
rect 4422 3364 4423 3368
rect 4427 3364 4428 3368
rect 4422 3363 4428 3364
rect 4670 3368 4676 3369
rect 4670 3364 4671 3368
rect 4675 3364 4676 3368
rect 4670 3363 4676 3364
rect 4894 3368 4900 3369
rect 4894 3364 4895 3368
rect 4899 3364 4900 3368
rect 4894 3363 4900 3364
rect 5110 3368 5116 3369
rect 5110 3364 5111 3368
rect 5115 3364 5116 3368
rect 5110 3363 5116 3364
rect 5326 3368 5332 3369
rect 5326 3364 5327 3368
rect 5331 3364 5332 3368
rect 5326 3363 5332 3364
rect 5542 3368 5548 3369
rect 5542 3364 5543 3368
rect 5547 3364 5548 3368
rect 5662 3365 5663 3369
rect 5667 3365 5668 3369
rect 5662 3364 5668 3365
rect 5542 3363 5548 3364
rect 3858 3353 3864 3354
rect 3838 3352 3844 3353
rect 3838 3348 3839 3352
rect 3843 3348 3844 3352
rect 3858 3349 3859 3353
rect 3863 3349 3864 3353
rect 3858 3348 3864 3349
rect 4122 3353 4128 3354
rect 4122 3349 4123 3353
rect 4127 3349 4128 3353
rect 4122 3348 4128 3349
rect 4394 3353 4400 3354
rect 4394 3349 4395 3353
rect 4399 3349 4400 3353
rect 4394 3348 4400 3349
rect 4642 3353 4648 3354
rect 4642 3349 4643 3353
rect 4647 3349 4648 3353
rect 4642 3348 4648 3349
rect 4866 3353 4872 3354
rect 4866 3349 4867 3353
rect 4871 3349 4872 3353
rect 4866 3348 4872 3349
rect 5082 3353 5088 3354
rect 5082 3349 5083 3353
rect 5087 3349 5088 3353
rect 5082 3348 5088 3349
rect 5298 3353 5304 3354
rect 5298 3349 5299 3353
rect 5303 3349 5304 3353
rect 5298 3348 5304 3349
rect 5514 3353 5520 3354
rect 5514 3349 5515 3353
rect 5519 3349 5520 3353
rect 5514 3348 5520 3349
rect 5662 3352 5668 3353
rect 5662 3348 5663 3352
rect 5667 3348 5668 3352
rect 3838 3347 3844 3348
rect 1975 3334 1979 3335
rect 1975 3329 1979 3330
rect 1995 3334 1999 3335
rect 1995 3329 1999 3330
rect 2163 3334 2167 3335
rect 2163 3329 2167 3330
rect 2195 3334 2199 3335
rect 2195 3329 2199 3330
rect 2371 3334 2375 3335
rect 2371 3329 2375 3330
rect 2411 3334 2415 3335
rect 2411 3329 2415 3330
rect 2587 3334 2591 3335
rect 2587 3329 2591 3330
rect 2619 3334 2623 3335
rect 2619 3329 2623 3330
rect 2803 3334 2807 3335
rect 2803 3329 2807 3330
rect 2811 3334 2815 3335
rect 2811 3329 2815 3330
rect 3003 3334 3007 3335
rect 3003 3329 3007 3330
rect 3019 3334 3023 3335
rect 3019 3329 3023 3330
rect 3187 3334 3191 3335
rect 3187 3329 3191 3330
rect 3235 3334 3239 3335
rect 3235 3329 3239 3330
rect 3371 3334 3375 3335
rect 3371 3329 3375 3330
rect 3451 3334 3455 3335
rect 3451 3329 3455 3330
rect 3555 3334 3559 3335
rect 3555 3329 3559 3330
rect 3651 3334 3655 3335
rect 3651 3329 3655 3330
rect 3799 3334 3803 3335
rect 3799 3329 3803 3330
rect 1934 3296 1940 3297
rect 110 3292 111 3296
rect 115 3292 116 3296
rect 110 3291 116 3292
rect 466 3295 472 3296
rect 466 3291 467 3295
rect 471 3291 472 3295
rect 466 3290 472 3291
rect 666 3295 672 3296
rect 666 3291 667 3295
rect 671 3291 672 3295
rect 666 3290 672 3291
rect 874 3295 880 3296
rect 874 3291 875 3295
rect 879 3291 880 3295
rect 874 3290 880 3291
rect 1090 3295 1096 3296
rect 1090 3291 1091 3295
rect 1095 3291 1096 3295
rect 1090 3290 1096 3291
rect 1314 3295 1320 3296
rect 1314 3291 1315 3295
rect 1319 3291 1320 3295
rect 1934 3292 1935 3296
rect 1939 3292 1940 3296
rect 1934 3291 1940 3292
rect 1314 3290 1320 3291
rect 494 3280 500 3281
rect 110 3279 116 3280
rect 110 3275 111 3279
rect 115 3275 116 3279
rect 494 3276 495 3280
rect 499 3276 500 3280
rect 494 3275 500 3276
rect 694 3280 700 3281
rect 694 3276 695 3280
rect 699 3276 700 3280
rect 694 3275 700 3276
rect 902 3280 908 3281
rect 902 3276 903 3280
rect 907 3276 908 3280
rect 902 3275 908 3276
rect 1118 3280 1124 3281
rect 1118 3276 1119 3280
rect 1123 3276 1124 3280
rect 1118 3275 1124 3276
rect 1342 3280 1348 3281
rect 1342 3276 1343 3280
rect 1347 3276 1348 3280
rect 1342 3275 1348 3276
rect 1934 3279 1940 3280
rect 1934 3275 1935 3279
rect 1939 3275 1940 3279
rect 110 3274 116 3275
rect 112 3251 114 3274
rect 496 3251 498 3275
rect 696 3251 698 3275
rect 904 3251 906 3275
rect 1120 3251 1122 3275
rect 1344 3251 1346 3275
rect 1934 3274 1940 3275
rect 1936 3251 1938 3274
rect 1976 3269 1978 3329
rect 1974 3268 1980 3269
rect 1996 3268 1998 3329
rect 2196 3268 2198 3329
rect 2412 3268 2414 3329
rect 2620 3268 2622 3329
rect 2812 3268 2814 3329
rect 3004 3268 3006 3329
rect 3188 3268 3190 3329
rect 3372 3268 3374 3329
rect 3556 3268 3558 3329
rect 3800 3269 3802 3329
rect 3840 3287 3842 3347
rect 3860 3287 3862 3348
rect 4124 3287 4126 3348
rect 4396 3287 4398 3348
rect 4644 3287 4646 3348
rect 4868 3287 4870 3348
rect 5084 3287 5086 3348
rect 5300 3287 5302 3348
rect 5516 3287 5518 3348
rect 5662 3347 5668 3348
rect 5664 3287 5666 3347
rect 3839 3286 3843 3287
rect 3839 3281 3843 3282
rect 3859 3286 3863 3287
rect 3859 3281 3863 3282
rect 4099 3286 4103 3287
rect 4099 3281 4103 3282
rect 4123 3286 4127 3287
rect 4123 3281 4127 3282
rect 4347 3286 4351 3287
rect 4347 3281 4351 3282
rect 4395 3286 4399 3287
rect 4395 3281 4399 3282
rect 4579 3286 4583 3287
rect 4579 3281 4583 3282
rect 4643 3286 4647 3287
rect 4643 3281 4647 3282
rect 4787 3286 4791 3287
rect 4787 3281 4791 3282
rect 4867 3286 4871 3287
rect 4867 3281 4871 3282
rect 4987 3286 4991 3287
rect 4987 3281 4991 3282
rect 5083 3286 5087 3287
rect 5083 3281 5087 3282
rect 5171 3286 5175 3287
rect 5171 3281 5175 3282
rect 5299 3286 5303 3287
rect 5299 3281 5303 3282
rect 5355 3286 5359 3287
rect 5355 3281 5359 3282
rect 5515 3286 5519 3287
rect 5515 3281 5519 3282
rect 5663 3286 5667 3287
rect 5663 3281 5667 3282
rect 3798 3268 3804 3269
rect 1974 3264 1975 3268
rect 1979 3264 1980 3268
rect 1974 3263 1980 3264
rect 1994 3267 2000 3268
rect 1994 3263 1995 3267
rect 1999 3263 2000 3267
rect 1994 3262 2000 3263
rect 2194 3267 2200 3268
rect 2194 3263 2195 3267
rect 2199 3263 2200 3267
rect 2194 3262 2200 3263
rect 2410 3267 2416 3268
rect 2410 3263 2411 3267
rect 2415 3263 2416 3267
rect 2410 3262 2416 3263
rect 2618 3267 2624 3268
rect 2618 3263 2619 3267
rect 2623 3263 2624 3267
rect 2618 3262 2624 3263
rect 2810 3267 2816 3268
rect 2810 3263 2811 3267
rect 2815 3263 2816 3267
rect 2810 3262 2816 3263
rect 3002 3267 3008 3268
rect 3002 3263 3003 3267
rect 3007 3263 3008 3267
rect 3002 3262 3008 3263
rect 3186 3267 3192 3268
rect 3186 3263 3187 3267
rect 3191 3263 3192 3267
rect 3186 3262 3192 3263
rect 3370 3267 3376 3268
rect 3370 3263 3371 3267
rect 3375 3263 3376 3267
rect 3370 3262 3376 3263
rect 3554 3267 3560 3268
rect 3554 3263 3555 3267
rect 3559 3263 3560 3267
rect 3798 3264 3799 3268
rect 3803 3264 3804 3268
rect 3798 3263 3804 3264
rect 3554 3262 3560 3263
rect 2022 3252 2028 3253
rect 1974 3251 1980 3252
rect 111 3250 115 3251
rect 111 3245 115 3246
rect 495 3250 499 3251
rect 495 3245 499 3246
rect 535 3250 539 3251
rect 535 3245 539 3246
rect 695 3250 699 3251
rect 695 3245 699 3246
rect 727 3250 731 3251
rect 727 3245 731 3246
rect 903 3250 907 3251
rect 903 3245 907 3246
rect 919 3250 923 3251
rect 919 3245 923 3246
rect 1111 3250 1115 3251
rect 1111 3245 1115 3246
rect 1119 3250 1123 3251
rect 1119 3245 1123 3246
rect 1295 3250 1299 3251
rect 1295 3245 1299 3246
rect 1343 3250 1347 3251
rect 1343 3245 1347 3246
rect 1471 3250 1475 3251
rect 1471 3245 1475 3246
rect 1655 3250 1659 3251
rect 1655 3245 1659 3246
rect 1815 3250 1819 3251
rect 1815 3245 1819 3246
rect 1935 3250 1939 3251
rect 1974 3247 1975 3251
rect 1979 3247 1980 3251
rect 2022 3248 2023 3252
rect 2027 3248 2028 3252
rect 2022 3247 2028 3248
rect 2222 3252 2228 3253
rect 2222 3248 2223 3252
rect 2227 3248 2228 3252
rect 2222 3247 2228 3248
rect 2438 3252 2444 3253
rect 2438 3248 2439 3252
rect 2443 3248 2444 3252
rect 2438 3247 2444 3248
rect 2646 3252 2652 3253
rect 2646 3248 2647 3252
rect 2651 3248 2652 3252
rect 2646 3247 2652 3248
rect 2838 3252 2844 3253
rect 2838 3248 2839 3252
rect 2843 3248 2844 3252
rect 2838 3247 2844 3248
rect 3030 3252 3036 3253
rect 3030 3248 3031 3252
rect 3035 3248 3036 3252
rect 3030 3247 3036 3248
rect 3214 3252 3220 3253
rect 3214 3248 3215 3252
rect 3219 3248 3220 3252
rect 3214 3247 3220 3248
rect 3398 3252 3404 3253
rect 3398 3248 3399 3252
rect 3403 3248 3404 3252
rect 3398 3247 3404 3248
rect 3582 3252 3588 3253
rect 3582 3248 3583 3252
rect 3587 3248 3588 3252
rect 3582 3247 3588 3248
rect 3798 3251 3804 3252
rect 3798 3247 3799 3251
rect 3803 3247 3804 3251
rect 1974 3246 1980 3247
rect 1935 3245 1939 3246
rect 112 3222 114 3245
rect 110 3221 116 3222
rect 536 3221 538 3245
rect 728 3221 730 3245
rect 920 3221 922 3245
rect 1112 3221 1114 3245
rect 1296 3221 1298 3245
rect 1472 3221 1474 3245
rect 1656 3221 1658 3245
rect 1816 3221 1818 3245
rect 1936 3222 1938 3245
rect 1976 3223 1978 3246
rect 2024 3223 2026 3247
rect 2224 3223 2226 3247
rect 2440 3223 2442 3247
rect 2648 3223 2650 3247
rect 2840 3223 2842 3247
rect 3032 3223 3034 3247
rect 3216 3223 3218 3247
rect 3400 3223 3402 3247
rect 3584 3223 3586 3247
rect 3798 3246 3804 3247
rect 3800 3223 3802 3246
rect 1975 3222 1979 3223
rect 1934 3221 1940 3222
rect 110 3217 111 3221
rect 115 3217 116 3221
rect 110 3216 116 3217
rect 534 3220 540 3221
rect 534 3216 535 3220
rect 539 3216 540 3220
rect 534 3215 540 3216
rect 726 3220 732 3221
rect 726 3216 727 3220
rect 731 3216 732 3220
rect 726 3215 732 3216
rect 918 3220 924 3221
rect 918 3216 919 3220
rect 923 3216 924 3220
rect 918 3215 924 3216
rect 1110 3220 1116 3221
rect 1110 3216 1111 3220
rect 1115 3216 1116 3220
rect 1110 3215 1116 3216
rect 1294 3220 1300 3221
rect 1294 3216 1295 3220
rect 1299 3216 1300 3220
rect 1294 3215 1300 3216
rect 1470 3220 1476 3221
rect 1470 3216 1471 3220
rect 1475 3216 1476 3220
rect 1470 3215 1476 3216
rect 1654 3220 1660 3221
rect 1654 3216 1655 3220
rect 1659 3216 1660 3220
rect 1654 3215 1660 3216
rect 1814 3220 1820 3221
rect 1814 3216 1815 3220
rect 1819 3216 1820 3220
rect 1934 3217 1935 3221
rect 1939 3217 1940 3221
rect 1975 3217 1979 3218
rect 2023 3222 2027 3223
rect 2023 3217 2027 3218
rect 2223 3222 2227 3223
rect 2223 3217 2227 3218
rect 2439 3222 2443 3223
rect 2439 3217 2443 3218
rect 2463 3222 2467 3223
rect 2463 3217 2467 3218
rect 2647 3222 2651 3223
rect 2647 3217 2651 3218
rect 2663 3222 2667 3223
rect 2663 3217 2667 3218
rect 2839 3222 2843 3223
rect 2839 3217 2843 3218
rect 2863 3222 2867 3223
rect 2863 3217 2867 3218
rect 3031 3222 3035 3223
rect 3031 3217 3035 3218
rect 3055 3222 3059 3223
rect 3055 3217 3059 3218
rect 3215 3222 3219 3223
rect 3215 3217 3219 3218
rect 3239 3222 3243 3223
rect 3239 3217 3243 3218
rect 3399 3222 3403 3223
rect 3399 3217 3403 3218
rect 3431 3222 3435 3223
rect 3431 3217 3435 3218
rect 3583 3222 3587 3223
rect 3583 3217 3587 3218
rect 3623 3222 3627 3223
rect 3623 3217 3627 3218
rect 3799 3222 3803 3223
rect 3840 3221 3842 3281
rect 3799 3217 3803 3218
rect 3838 3220 3844 3221
rect 3860 3220 3862 3281
rect 4100 3220 4102 3281
rect 4348 3220 4350 3281
rect 4580 3220 4582 3281
rect 4788 3220 4790 3281
rect 4988 3220 4990 3281
rect 5172 3220 5174 3281
rect 5356 3220 5358 3281
rect 5516 3220 5518 3281
rect 5664 3221 5666 3281
rect 5662 3220 5668 3221
rect 1934 3216 1940 3217
rect 1814 3215 1820 3216
rect 506 3205 512 3206
rect 110 3204 116 3205
rect 110 3200 111 3204
rect 115 3200 116 3204
rect 506 3201 507 3205
rect 511 3201 512 3205
rect 506 3200 512 3201
rect 698 3205 704 3206
rect 698 3201 699 3205
rect 703 3201 704 3205
rect 698 3200 704 3201
rect 890 3205 896 3206
rect 890 3201 891 3205
rect 895 3201 896 3205
rect 890 3200 896 3201
rect 1082 3205 1088 3206
rect 1082 3201 1083 3205
rect 1087 3201 1088 3205
rect 1082 3200 1088 3201
rect 1266 3205 1272 3206
rect 1266 3201 1267 3205
rect 1271 3201 1272 3205
rect 1266 3200 1272 3201
rect 1442 3205 1448 3206
rect 1442 3201 1443 3205
rect 1447 3201 1448 3205
rect 1442 3200 1448 3201
rect 1626 3205 1632 3206
rect 1626 3201 1627 3205
rect 1631 3201 1632 3205
rect 1626 3200 1632 3201
rect 1786 3205 1792 3206
rect 1786 3201 1787 3205
rect 1791 3201 1792 3205
rect 1786 3200 1792 3201
rect 1934 3204 1940 3205
rect 1934 3200 1935 3204
rect 1939 3200 1940 3204
rect 110 3199 116 3200
rect 112 3131 114 3199
rect 508 3131 510 3200
rect 700 3131 702 3200
rect 892 3131 894 3200
rect 1084 3131 1086 3200
rect 1268 3131 1270 3200
rect 1444 3131 1446 3200
rect 1628 3131 1630 3200
rect 1788 3131 1790 3200
rect 1934 3199 1940 3200
rect 1936 3131 1938 3199
rect 1976 3194 1978 3217
rect 1974 3193 1980 3194
rect 2464 3193 2466 3217
rect 2664 3193 2666 3217
rect 2864 3193 2866 3217
rect 3056 3193 3058 3217
rect 3240 3193 3242 3217
rect 3432 3193 3434 3217
rect 3624 3193 3626 3217
rect 3800 3194 3802 3217
rect 3838 3216 3839 3220
rect 3843 3216 3844 3220
rect 3838 3215 3844 3216
rect 3858 3219 3864 3220
rect 3858 3215 3859 3219
rect 3863 3215 3864 3219
rect 3858 3214 3864 3215
rect 4098 3219 4104 3220
rect 4098 3215 4099 3219
rect 4103 3215 4104 3219
rect 4098 3214 4104 3215
rect 4346 3219 4352 3220
rect 4346 3215 4347 3219
rect 4351 3215 4352 3219
rect 4346 3214 4352 3215
rect 4578 3219 4584 3220
rect 4578 3215 4579 3219
rect 4583 3215 4584 3219
rect 4578 3214 4584 3215
rect 4786 3219 4792 3220
rect 4786 3215 4787 3219
rect 4791 3215 4792 3219
rect 4786 3214 4792 3215
rect 4986 3219 4992 3220
rect 4986 3215 4987 3219
rect 4991 3215 4992 3219
rect 4986 3214 4992 3215
rect 5170 3219 5176 3220
rect 5170 3215 5171 3219
rect 5175 3215 5176 3219
rect 5170 3214 5176 3215
rect 5354 3219 5360 3220
rect 5354 3215 5355 3219
rect 5359 3215 5360 3219
rect 5354 3214 5360 3215
rect 5514 3219 5520 3220
rect 5514 3215 5515 3219
rect 5519 3215 5520 3219
rect 5662 3216 5663 3220
rect 5667 3216 5668 3220
rect 5662 3215 5668 3216
rect 5514 3214 5520 3215
rect 3886 3204 3892 3205
rect 3838 3203 3844 3204
rect 3838 3199 3839 3203
rect 3843 3199 3844 3203
rect 3886 3200 3887 3204
rect 3891 3200 3892 3204
rect 3886 3199 3892 3200
rect 4126 3204 4132 3205
rect 4126 3200 4127 3204
rect 4131 3200 4132 3204
rect 4126 3199 4132 3200
rect 4374 3204 4380 3205
rect 4374 3200 4375 3204
rect 4379 3200 4380 3204
rect 4374 3199 4380 3200
rect 4606 3204 4612 3205
rect 4606 3200 4607 3204
rect 4611 3200 4612 3204
rect 4606 3199 4612 3200
rect 4814 3204 4820 3205
rect 4814 3200 4815 3204
rect 4819 3200 4820 3204
rect 4814 3199 4820 3200
rect 5014 3204 5020 3205
rect 5014 3200 5015 3204
rect 5019 3200 5020 3204
rect 5014 3199 5020 3200
rect 5198 3204 5204 3205
rect 5198 3200 5199 3204
rect 5203 3200 5204 3204
rect 5198 3199 5204 3200
rect 5382 3204 5388 3205
rect 5382 3200 5383 3204
rect 5387 3200 5388 3204
rect 5382 3199 5388 3200
rect 5542 3204 5548 3205
rect 5542 3200 5543 3204
rect 5547 3200 5548 3204
rect 5542 3199 5548 3200
rect 5662 3203 5668 3204
rect 5662 3199 5663 3203
rect 5667 3199 5668 3203
rect 3838 3198 3844 3199
rect 3798 3193 3804 3194
rect 1974 3189 1975 3193
rect 1979 3189 1980 3193
rect 1974 3188 1980 3189
rect 2462 3192 2468 3193
rect 2462 3188 2463 3192
rect 2467 3188 2468 3192
rect 2462 3187 2468 3188
rect 2662 3192 2668 3193
rect 2662 3188 2663 3192
rect 2667 3188 2668 3192
rect 2662 3187 2668 3188
rect 2862 3192 2868 3193
rect 2862 3188 2863 3192
rect 2867 3188 2868 3192
rect 2862 3187 2868 3188
rect 3054 3192 3060 3193
rect 3054 3188 3055 3192
rect 3059 3188 3060 3192
rect 3054 3187 3060 3188
rect 3238 3192 3244 3193
rect 3238 3188 3239 3192
rect 3243 3188 3244 3192
rect 3238 3187 3244 3188
rect 3430 3192 3436 3193
rect 3430 3188 3431 3192
rect 3435 3188 3436 3192
rect 3430 3187 3436 3188
rect 3622 3192 3628 3193
rect 3622 3188 3623 3192
rect 3627 3188 3628 3192
rect 3798 3189 3799 3193
rect 3803 3189 3804 3193
rect 3798 3188 3804 3189
rect 3622 3187 3628 3188
rect 2434 3177 2440 3178
rect 1974 3176 1980 3177
rect 1974 3172 1975 3176
rect 1979 3172 1980 3176
rect 2434 3173 2435 3177
rect 2439 3173 2440 3177
rect 2434 3172 2440 3173
rect 2634 3177 2640 3178
rect 2634 3173 2635 3177
rect 2639 3173 2640 3177
rect 2634 3172 2640 3173
rect 2834 3177 2840 3178
rect 2834 3173 2835 3177
rect 2839 3173 2840 3177
rect 2834 3172 2840 3173
rect 3026 3177 3032 3178
rect 3026 3173 3027 3177
rect 3031 3173 3032 3177
rect 3026 3172 3032 3173
rect 3210 3177 3216 3178
rect 3210 3173 3211 3177
rect 3215 3173 3216 3177
rect 3210 3172 3216 3173
rect 3402 3177 3408 3178
rect 3402 3173 3403 3177
rect 3407 3173 3408 3177
rect 3402 3172 3408 3173
rect 3594 3177 3600 3178
rect 3594 3173 3595 3177
rect 3599 3173 3600 3177
rect 3594 3172 3600 3173
rect 3798 3176 3804 3177
rect 3798 3172 3799 3176
rect 3803 3172 3804 3176
rect 1974 3171 1980 3172
rect 111 3130 115 3131
rect 111 3125 115 3126
rect 427 3130 431 3131
rect 427 3125 431 3126
rect 507 3130 511 3131
rect 507 3125 511 3126
rect 563 3130 567 3131
rect 563 3125 567 3126
rect 699 3130 703 3131
rect 699 3125 703 3126
rect 835 3130 839 3131
rect 835 3125 839 3126
rect 891 3130 895 3131
rect 891 3125 895 3126
rect 971 3130 975 3131
rect 971 3125 975 3126
rect 1083 3130 1087 3131
rect 1083 3125 1087 3126
rect 1107 3130 1111 3131
rect 1107 3125 1111 3126
rect 1243 3130 1247 3131
rect 1243 3125 1247 3126
rect 1267 3130 1271 3131
rect 1267 3125 1271 3126
rect 1379 3130 1383 3131
rect 1379 3125 1383 3126
rect 1443 3130 1447 3131
rect 1443 3125 1447 3126
rect 1515 3130 1519 3131
rect 1515 3125 1519 3126
rect 1627 3130 1631 3131
rect 1627 3125 1631 3126
rect 1651 3130 1655 3131
rect 1651 3125 1655 3126
rect 1787 3130 1791 3131
rect 1787 3125 1791 3126
rect 1935 3130 1939 3131
rect 1935 3125 1939 3126
rect 112 3065 114 3125
rect 110 3064 116 3065
rect 428 3064 430 3125
rect 564 3064 566 3125
rect 700 3064 702 3125
rect 836 3064 838 3125
rect 972 3064 974 3125
rect 1108 3064 1110 3125
rect 1244 3064 1246 3125
rect 1380 3064 1382 3125
rect 1516 3064 1518 3125
rect 1652 3064 1654 3125
rect 1788 3064 1790 3125
rect 1936 3065 1938 3125
rect 1976 3099 1978 3171
rect 2436 3099 2438 3172
rect 2636 3099 2638 3172
rect 2836 3099 2838 3172
rect 3028 3099 3030 3172
rect 3212 3099 3214 3172
rect 3404 3099 3406 3172
rect 3596 3099 3598 3172
rect 3798 3171 3804 3172
rect 3800 3099 3802 3171
rect 3840 3159 3842 3198
rect 3888 3159 3890 3199
rect 4128 3159 4130 3199
rect 4376 3159 4378 3199
rect 4608 3159 4610 3199
rect 4816 3159 4818 3199
rect 5016 3159 5018 3199
rect 5200 3159 5202 3199
rect 5384 3159 5386 3199
rect 5544 3159 5546 3199
rect 5662 3198 5668 3199
rect 5664 3159 5666 3198
rect 3839 3158 3843 3159
rect 3839 3153 3843 3154
rect 3887 3158 3891 3159
rect 3887 3153 3891 3154
rect 3903 3158 3907 3159
rect 3903 3153 3907 3154
rect 4127 3158 4131 3159
rect 4127 3153 4131 3154
rect 4135 3158 4139 3159
rect 4135 3153 4139 3154
rect 4359 3158 4363 3159
rect 4359 3153 4363 3154
rect 4375 3158 4379 3159
rect 4375 3153 4379 3154
rect 4583 3158 4587 3159
rect 4583 3153 4587 3154
rect 4607 3158 4611 3159
rect 4607 3153 4611 3154
rect 4807 3158 4811 3159
rect 4807 3153 4811 3154
rect 4815 3158 4819 3159
rect 4815 3153 4819 3154
rect 5015 3158 5019 3159
rect 5015 3153 5019 3154
rect 5031 3158 5035 3159
rect 5031 3153 5035 3154
rect 5199 3158 5203 3159
rect 5199 3153 5203 3154
rect 5383 3158 5387 3159
rect 5383 3153 5387 3154
rect 5543 3158 5547 3159
rect 5543 3153 5547 3154
rect 5663 3158 5667 3159
rect 5663 3153 5667 3154
rect 3840 3130 3842 3153
rect 3838 3129 3844 3130
rect 3904 3129 3906 3153
rect 4136 3129 4138 3153
rect 4360 3129 4362 3153
rect 4584 3129 4586 3153
rect 4808 3129 4810 3153
rect 5032 3129 5034 3153
rect 5664 3130 5666 3153
rect 5662 3129 5668 3130
rect 3838 3125 3839 3129
rect 3843 3125 3844 3129
rect 3838 3124 3844 3125
rect 3902 3128 3908 3129
rect 3902 3124 3903 3128
rect 3907 3124 3908 3128
rect 3902 3123 3908 3124
rect 4134 3128 4140 3129
rect 4134 3124 4135 3128
rect 4139 3124 4140 3128
rect 4134 3123 4140 3124
rect 4358 3128 4364 3129
rect 4358 3124 4359 3128
rect 4363 3124 4364 3128
rect 4358 3123 4364 3124
rect 4582 3128 4588 3129
rect 4582 3124 4583 3128
rect 4587 3124 4588 3128
rect 4582 3123 4588 3124
rect 4806 3128 4812 3129
rect 4806 3124 4807 3128
rect 4811 3124 4812 3128
rect 4806 3123 4812 3124
rect 5030 3128 5036 3129
rect 5030 3124 5031 3128
rect 5035 3124 5036 3128
rect 5662 3125 5663 3129
rect 5667 3125 5668 3129
rect 5662 3124 5668 3125
rect 5030 3123 5036 3124
rect 3874 3113 3880 3114
rect 3838 3112 3844 3113
rect 3838 3108 3839 3112
rect 3843 3108 3844 3112
rect 3874 3109 3875 3113
rect 3879 3109 3880 3113
rect 3874 3108 3880 3109
rect 4106 3113 4112 3114
rect 4106 3109 4107 3113
rect 4111 3109 4112 3113
rect 4106 3108 4112 3109
rect 4330 3113 4336 3114
rect 4330 3109 4331 3113
rect 4335 3109 4336 3113
rect 4330 3108 4336 3109
rect 4554 3113 4560 3114
rect 4554 3109 4555 3113
rect 4559 3109 4560 3113
rect 4554 3108 4560 3109
rect 4778 3113 4784 3114
rect 4778 3109 4779 3113
rect 4783 3109 4784 3113
rect 4778 3108 4784 3109
rect 5002 3113 5008 3114
rect 5002 3109 5003 3113
rect 5007 3109 5008 3113
rect 5002 3108 5008 3109
rect 5662 3112 5668 3113
rect 5662 3108 5663 3112
rect 5667 3108 5668 3112
rect 3838 3107 3844 3108
rect 1975 3098 1979 3099
rect 1975 3093 1979 3094
rect 2331 3098 2335 3099
rect 2331 3093 2335 3094
rect 2435 3098 2439 3099
rect 2435 3093 2439 3094
rect 2555 3098 2559 3099
rect 2555 3093 2559 3094
rect 2635 3098 2639 3099
rect 2635 3093 2639 3094
rect 2779 3098 2783 3099
rect 2779 3093 2783 3094
rect 2835 3098 2839 3099
rect 2835 3093 2839 3094
rect 3003 3098 3007 3099
rect 3003 3093 3007 3094
rect 3027 3098 3031 3099
rect 3027 3093 3031 3094
rect 3211 3098 3215 3099
rect 3211 3093 3215 3094
rect 3235 3098 3239 3099
rect 3235 3093 3239 3094
rect 3403 3098 3407 3099
rect 3403 3093 3407 3094
rect 3467 3098 3471 3099
rect 3467 3093 3471 3094
rect 3595 3098 3599 3099
rect 3595 3093 3599 3094
rect 3799 3098 3803 3099
rect 3799 3093 3803 3094
rect 1934 3064 1940 3065
rect 110 3060 111 3064
rect 115 3060 116 3064
rect 110 3059 116 3060
rect 426 3063 432 3064
rect 426 3059 427 3063
rect 431 3059 432 3063
rect 426 3058 432 3059
rect 562 3063 568 3064
rect 562 3059 563 3063
rect 567 3059 568 3063
rect 562 3058 568 3059
rect 698 3063 704 3064
rect 698 3059 699 3063
rect 703 3059 704 3063
rect 698 3058 704 3059
rect 834 3063 840 3064
rect 834 3059 835 3063
rect 839 3059 840 3063
rect 834 3058 840 3059
rect 970 3063 976 3064
rect 970 3059 971 3063
rect 975 3059 976 3063
rect 970 3058 976 3059
rect 1106 3063 1112 3064
rect 1106 3059 1107 3063
rect 1111 3059 1112 3063
rect 1106 3058 1112 3059
rect 1242 3063 1248 3064
rect 1242 3059 1243 3063
rect 1247 3059 1248 3063
rect 1242 3058 1248 3059
rect 1378 3063 1384 3064
rect 1378 3059 1379 3063
rect 1383 3059 1384 3063
rect 1378 3058 1384 3059
rect 1514 3063 1520 3064
rect 1514 3059 1515 3063
rect 1519 3059 1520 3063
rect 1514 3058 1520 3059
rect 1650 3063 1656 3064
rect 1650 3059 1651 3063
rect 1655 3059 1656 3063
rect 1650 3058 1656 3059
rect 1786 3063 1792 3064
rect 1786 3059 1787 3063
rect 1791 3059 1792 3063
rect 1934 3060 1935 3064
rect 1939 3060 1940 3064
rect 1934 3059 1940 3060
rect 1786 3058 1792 3059
rect 454 3048 460 3049
rect 110 3047 116 3048
rect 110 3043 111 3047
rect 115 3043 116 3047
rect 454 3044 455 3048
rect 459 3044 460 3048
rect 454 3043 460 3044
rect 590 3048 596 3049
rect 590 3044 591 3048
rect 595 3044 596 3048
rect 590 3043 596 3044
rect 726 3048 732 3049
rect 726 3044 727 3048
rect 731 3044 732 3048
rect 726 3043 732 3044
rect 862 3048 868 3049
rect 862 3044 863 3048
rect 867 3044 868 3048
rect 862 3043 868 3044
rect 998 3048 1004 3049
rect 998 3044 999 3048
rect 1003 3044 1004 3048
rect 998 3043 1004 3044
rect 1134 3048 1140 3049
rect 1134 3044 1135 3048
rect 1139 3044 1140 3048
rect 1134 3043 1140 3044
rect 1270 3048 1276 3049
rect 1270 3044 1271 3048
rect 1275 3044 1276 3048
rect 1270 3043 1276 3044
rect 1406 3048 1412 3049
rect 1406 3044 1407 3048
rect 1411 3044 1412 3048
rect 1406 3043 1412 3044
rect 1542 3048 1548 3049
rect 1542 3044 1543 3048
rect 1547 3044 1548 3048
rect 1542 3043 1548 3044
rect 1678 3048 1684 3049
rect 1678 3044 1679 3048
rect 1683 3044 1684 3048
rect 1678 3043 1684 3044
rect 1814 3048 1820 3049
rect 1814 3044 1815 3048
rect 1819 3044 1820 3048
rect 1814 3043 1820 3044
rect 1934 3047 1940 3048
rect 1934 3043 1935 3047
rect 1939 3043 1940 3047
rect 110 3042 116 3043
rect 112 2991 114 3042
rect 456 2991 458 3043
rect 592 2991 594 3043
rect 728 2991 730 3043
rect 864 2991 866 3043
rect 1000 2991 1002 3043
rect 1136 2991 1138 3043
rect 1272 2991 1274 3043
rect 1408 2991 1410 3043
rect 1544 2991 1546 3043
rect 1680 2991 1682 3043
rect 1816 2991 1818 3043
rect 1934 3042 1940 3043
rect 1936 2991 1938 3042
rect 1976 3033 1978 3093
rect 1974 3032 1980 3033
rect 2332 3032 2334 3093
rect 2556 3032 2558 3093
rect 2780 3032 2782 3093
rect 3004 3032 3006 3093
rect 3236 3032 3238 3093
rect 3468 3032 3470 3093
rect 3800 3033 3802 3093
rect 3840 3047 3842 3107
rect 3876 3047 3878 3108
rect 4108 3047 4110 3108
rect 4332 3047 4334 3108
rect 4556 3047 4558 3108
rect 4780 3047 4782 3108
rect 5004 3047 5006 3108
rect 5662 3107 5668 3108
rect 5664 3047 5666 3107
rect 3839 3046 3843 3047
rect 3839 3041 3843 3042
rect 3875 3046 3879 3047
rect 3875 3041 3879 3042
rect 3907 3046 3911 3047
rect 3907 3041 3911 3042
rect 4075 3046 4079 3047
rect 4075 3041 4079 3042
rect 4107 3046 4111 3047
rect 4107 3041 4111 3042
rect 4243 3046 4247 3047
rect 4243 3041 4247 3042
rect 4331 3046 4335 3047
rect 4331 3041 4335 3042
rect 4411 3046 4415 3047
rect 4411 3041 4415 3042
rect 4555 3046 4559 3047
rect 4555 3041 4559 3042
rect 4579 3046 4583 3047
rect 4579 3041 4583 3042
rect 4755 3046 4759 3047
rect 4755 3041 4759 3042
rect 4779 3046 4783 3047
rect 4779 3041 4783 3042
rect 5003 3046 5007 3047
rect 5003 3041 5007 3042
rect 5663 3046 5667 3047
rect 5663 3041 5667 3042
rect 3798 3032 3804 3033
rect 1974 3028 1975 3032
rect 1979 3028 1980 3032
rect 1974 3027 1980 3028
rect 2330 3031 2336 3032
rect 2330 3027 2331 3031
rect 2335 3027 2336 3031
rect 2330 3026 2336 3027
rect 2554 3031 2560 3032
rect 2554 3027 2555 3031
rect 2559 3027 2560 3031
rect 2554 3026 2560 3027
rect 2778 3031 2784 3032
rect 2778 3027 2779 3031
rect 2783 3027 2784 3031
rect 2778 3026 2784 3027
rect 3002 3031 3008 3032
rect 3002 3027 3003 3031
rect 3007 3027 3008 3031
rect 3002 3026 3008 3027
rect 3234 3031 3240 3032
rect 3234 3027 3235 3031
rect 3239 3027 3240 3031
rect 3234 3026 3240 3027
rect 3466 3031 3472 3032
rect 3466 3027 3467 3031
rect 3471 3027 3472 3031
rect 3798 3028 3799 3032
rect 3803 3028 3804 3032
rect 3798 3027 3804 3028
rect 3466 3026 3472 3027
rect 2358 3016 2364 3017
rect 1974 3015 1980 3016
rect 1974 3011 1975 3015
rect 1979 3011 1980 3015
rect 2358 3012 2359 3016
rect 2363 3012 2364 3016
rect 2358 3011 2364 3012
rect 2582 3016 2588 3017
rect 2582 3012 2583 3016
rect 2587 3012 2588 3016
rect 2582 3011 2588 3012
rect 2806 3016 2812 3017
rect 2806 3012 2807 3016
rect 2811 3012 2812 3016
rect 2806 3011 2812 3012
rect 3030 3016 3036 3017
rect 3030 3012 3031 3016
rect 3035 3012 3036 3016
rect 3030 3011 3036 3012
rect 3262 3016 3268 3017
rect 3262 3012 3263 3016
rect 3267 3012 3268 3016
rect 3262 3011 3268 3012
rect 3494 3016 3500 3017
rect 3494 3012 3495 3016
rect 3499 3012 3500 3016
rect 3494 3011 3500 3012
rect 3798 3015 3804 3016
rect 3798 3011 3799 3015
rect 3803 3011 3804 3015
rect 1974 3010 1980 3011
rect 111 2990 115 2991
rect 111 2985 115 2986
rect 199 2990 203 2991
rect 199 2985 203 2986
rect 455 2990 459 2991
rect 455 2985 459 2986
rect 511 2990 515 2991
rect 511 2985 515 2986
rect 591 2990 595 2991
rect 591 2985 595 2986
rect 727 2990 731 2991
rect 727 2985 731 2986
rect 815 2990 819 2991
rect 815 2985 819 2986
rect 863 2990 867 2991
rect 863 2985 867 2986
rect 999 2990 1003 2991
rect 999 2985 1003 2986
rect 1111 2990 1115 2991
rect 1111 2985 1115 2986
rect 1135 2990 1139 2991
rect 1135 2985 1139 2986
rect 1271 2990 1275 2991
rect 1271 2985 1275 2986
rect 1407 2990 1411 2991
rect 1407 2985 1411 2986
rect 1415 2990 1419 2991
rect 1415 2985 1419 2986
rect 1543 2990 1547 2991
rect 1543 2985 1547 2986
rect 1679 2990 1683 2991
rect 1679 2985 1683 2986
rect 1719 2990 1723 2991
rect 1719 2985 1723 2986
rect 1815 2990 1819 2991
rect 1815 2985 1819 2986
rect 1935 2990 1939 2991
rect 1935 2985 1939 2986
rect 112 2962 114 2985
rect 110 2961 116 2962
rect 200 2961 202 2985
rect 512 2961 514 2985
rect 816 2961 818 2985
rect 1112 2961 1114 2985
rect 1416 2961 1418 2985
rect 1720 2961 1722 2985
rect 1936 2962 1938 2985
rect 1976 2975 1978 3010
rect 2360 2975 2362 3011
rect 2584 2975 2586 3011
rect 2808 2975 2810 3011
rect 3032 2975 3034 3011
rect 3264 2975 3266 3011
rect 3496 2975 3498 3011
rect 3798 3010 3804 3011
rect 3800 2975 3802 3010
rect 3840 2981 3842 3041
rect 3838 2980 3844 2981
rect 3908 2980 3910 3041
rect 4076 2980 4078 3041
rect 4244 2980 4246 3041
rect 4412 2980 4414 3041
rect 4580 2980 4582 3041
rect 4756 2980 4758 3041
rect 5664 2981 5666 3041
rect 5662 2980 5668 2981
rect 3838 2976 3839 2980
rect 3843 2976 3844 2980
rect 3838 2975 3844 2976
rect 3906 2979 3912 2980
rect 3906 2975 3907 2979
rect 3911 2975 3912 2979
rect 1975 2974 1979 2975
rect 1975 2969 1979 2970
rect 2143 2974 2147 2975
rect 2143 2969 2147 2970
rect 2343 2974 2347 2975
rect 2343 2969 2347 2970
rect 2359 2974 2363 2975
rect 2359 2969 2363 2970
rect 2543 2974 2547 2975
rect 2543 2969 2547 2970
rect 2583 2974 2587 2975
rect 2583 2969 2587 2970
rect 2743 2974 2747 2975
rect 2743 2969 2747 2970
rect 2807 2974 2811 2975
rect 2807 2969 2811 2970
rect 2935 2974 2939 2975
rect 2935 2969 2939 2970
rect 3031 2974 3035 2975
rect 3031 2969 3035 2970
rect 3135 2974 3139 2975
rect 3135 2969 3139 2970
rect 3263 2974 3267 2975
rect 3263 2969 3267 2970
rect 3335 2974 3339 2975
rect 3335 2969 3339 2970
rect 3495 2974 3499 2975
rect 3495 2969 3499 2970
rect 3799 2974 3803 2975
rect 3906 2974 3912 2975
rect 4074 2979 4080 2980
rect 4074 2975 4075 2979
rect 4079 2975 4080 2979
rect 4074 2974 4080 2975
rect 4242 2979 4248 2980
rect 4242 2975 4243 2979
rect 4247 2975 4248 2979
rect 4242 2974 4248 2975
rect 4410 2979 4416 2980
rect 4410 2975 4411 2979
rect 4415 2975 4416 2979
rect 4410 2974 4416 2975
rect 4578 2979 4584 2980
rect 4578 2975 4579 2979
rect 4583 2975 4584 2979
rect 4578 2974 4584 2975
rect 4754 2979 4760 2980
rect 4754 2975 4755 2979
rect 4759 2975 4760 2979
rect 5662 2976 5663 2980
rect 5667 2976 5668 2980
rect 5662 2975 5668 2976
rect 4754 2974 4760 2975
rect 3799 2969 3803 2970
rect 1934 2961 1940 2962
rect 110 2957 111 2961
rect 115 2957 116 2961
rect 110 2956 116 2957
rect 198 2960 204 2961
rect 198 2956 199 2960
rect 203 2956 204 2960
rect 198 2955 204 2956
rect 510 2960 516 2961
rect 510 2956 511 2960
rect 515 2956 516 2960
rect 510 2955 516 2956
rect 814 2960 820 2961
rect 814 2956 815 2960
rect 819 2956 820 2960
rect 814 2955 820 2956
rect 1110 2960 1116 2961
rect 1110 2956 1111 2960
rect 1115 2956 1116 2960
rect 1110 2955 1116 2956
rect 1414 2960 1420 2961
rect 1414 2956 1415 2960
rect 1419 2956 1420 2960
rect 1414 2955 1420 2956
rect 1718 2960 1724 2961
rect 1718 2956 1719 2960
rect 1723 2956 1724 2960
rect 1934 2957 1935 2961
rect 1939 2957 1940 2961
rect 1934 2956 1940 2957
rect 1718 2955 1724 2956
rect 1976 2946 1978 2969
rect 170 2945 176 2946
rect 110 2944 116 2945
rect 110 2940 111 2944
rect 115 2940 116 2944
rect 170 2941 171 2945
rect 175 2941 176 2945
rect 170 2940 176 2941
rect 482 2945 488 2946
rect 482 2941 483 2945
rect 487 2941 488 2945
rect 482 2940 488 2941
rect 786 2945 792 2946
rect 786 2941 787 2945
rect 791 2941 792 2945
rect 786 2940 792 2941
rect 1082 2945 1088 2946
rect 1082 2941 1083 2945
rect 1087 2941 1088 2945
rect 1082 2940 1088 2941
rect 1386 2945 1392 2946
rect 1386 2941 1387 2945
rect 1391 2941 1392 2945
rect 1386 2940 1392 2941
rect 1690 2945 1696 2946
rect 1974 2945 1980 2946
rect 2144 2945 2146 2969
rect 2344 2945 2346 2969
rect 2544 2945 2546 2969
rect 2744 2945 2746 2969
rect 2936 2945 2938 2969
rect 3136 2945 3138 2969
rect 3336 2945 3338 2969
rect 3800 2946 3802 2969
rect 3934 2964 3940 2965
rect 3838 2963 3844 2964
rect 3838 2959 3839 2963
rect 3843 2959 3844 2963
rect 3934 2960 3935 2964
rect 3939 2960 3940 2964
rect 3934 2959 3940 2960
rect 4102 2964 4108 2965
rect 4102 2960 4103 2964
rect 4107 2960 4108 2964
rect 4102 2959 4108 2960
rect 4270 2964 4276 2965
rect 4270 2960 4271 2964
rect 4275 2960 4276 2964
rect 4270 2959 4276 2960
rect 4438 2964 4444 2965
rect 4438 2960 4439 2964
rect 4443 2960 4444 2964
rect 4438 2959 4444 2960
rect 4606 2964 4612 2965
rect 4606 2960 4607 2964
rect 4611 2960 4612 2964
rect 4606 2959 4612 2960
rect 4782 2964 4788 2965
rect 4782 2960 4783 2964
rect 4787 2960 4788 2964
rect 4782 2959 4788 2960
rect 5662 2963 5668 2964
rect 5662 2959 5663 2963
rect 5667 2959 5668 2963
rect 3838 2958 3844 2959
rect 3798 2945 3804 2946
rect 1690 2941 1691 2945
rect 1695 2941 1696 2945
rect 1690 2940 1696 2941
rect 1934 2944 1940 2945
rect 1934 2940 1935 2944
rect 1939 2940 1940 2944
rect 1974 2941 1975 2945
rect 1979 2941 1980 2945
rect 1974 2940 1980 2941
rect 2142 2944 2148 2945
rect 2142 2940 2143 2944
rect 2147 2940 2148 2944
rect 110 2939 116 2940
rect 112 2879 114 2939
rect 172 2879 174 2940
rect 484 2879 486 2940
rect 788 2879 790 2940
rect 1084 2879 1086 2940
rect 1388 2879 1390 2940
rect 1692 2879 1694 2940
rect 1934 2939 1940 2940
rect 2142 2939 2148 2940
rect 2342 2944 2348 2945
rect 2342 2940 2343 2944
rect 2347 2940 2348 2944
rect 2342 2939 2348 2940
rect 2542 2944 2548 2945
rect 2542 2940 2543 2944
rect 2547 2940 2548 2944
rect 2542 2939 2548 2940
rect 2742 2944 2748 2945
rect 2742 2940 2743 2944
rect 2747 2940 2748 2944
rect 2742 2939 2748 2940
rect 2934 2944 2940 2945
rect 2934 2940 2935 2944
rect 2939 2940 2940 2944
rect 2934 2939 2940 2940
rect 3134 2944 3140 2945
rect 3134 2940 3135 2944
rect 3139 2940 3140 2944
rect 3134 2939 3140 2940
rect 3334 2944 3340 2945
rect 3334 2940 3335 2944
rect 3339 2940 3340 2944
rect 3798 2941 3799 2945
rect 3803 2941 3804 2945
rect 3798 2940 3804 2941
rect 3334 2939 3340 2940
rect 1936 2879 1938 2939
rect 3840 2931 3842 2958
rect 3936 2931 3938 2959
rect 4104 2931 4106 2959
rect 4272 2931 4274 2959
rect 4440 2931 4442 2959
rect 4608 2931 4610 2959
rect 4784 2931 4786 2959
rect 5662 2958 5668 2959
rect 5664 2931 5666 2958
rect 3839 2930 3843 2931
rect 2114 2929 2120 2930
rect 1974 2928 1980 2929
rect 1974 2924 1975 2928
rect 1979 2924 1980 2928
rect 2114 2925 2115 2929
rect 2119 2925 2120 2929
rect 2114 2924 2120 2925
rect 2314 2929 2320 2930
rect 2314 2925 2315 2929
rect 2319 2925 2320 2929
rect 2314 2924 2320 2925
rect 2514 2929 2520 2930
rect 2514 2925 2515 2929
rect 2519 2925 2520 2929
rect 2514 2924 2520 2925
rect 2714 2929 2720 2930
rect 2714 2925 2715 2929
rect 2719 2925 2720 2929
rect 2714 2924 2720 2925
rect 2906 2929 2912 2930
rect 2906 2925 2907 2929
rect 2911 2925 2912 2929
rect 2906 2924 2912 2925
rect 3106 2929 3112 2930
rect 3106 2925 3107 2929
rect 3111 2925 3112 2929
rect 3106 2924 3112 2925
rect 3306 2929 3312 2930
rect 3306 2925 3307 2929
rect 3311 2925 3312 2929
rect 3306 2924 3312 2925
rect 3798 2928 3804 2929
rect 3798 2924 3799 2928
rect 3803 2924 3804 2928
rect 3839 2925 3843 2926
rect 3895 2930 3899 2931
rect 3895 2925 3899 2926
rect 3935 2930 3939 2931
rect 3935 2925 3939 2926
rect 4031 2930 4035 2931
rect 4031 2925 4035 2926
rect 4103 2930 4107 2931
rect 4103 2925 4107 2926
rect 4167 2930 4171 2931
rect 4167 2925 4171 2926
rect 4271 2930 4275 2931
rect 4271 2925 4275 2926
rect 4303 2930 4307 2931
rect 4303 2925 4307 2926
rect 4439 2930 4443 2931
rect 4439 2925 4443 2926
rect 4575 2930 4579 2931
rect 4575 2925 4579 2926
rect 4607 2930 4611 2931
rect 4607 2925 4611 2926
rect 4783 2930 4787 2931
rect 4783 2925 4787 2926
rect 5663 2930 5667 2931
rect 5663 2925 5667 2926
rect 1974 2923 1980 2924
rect 111 2878 115 2879
rect 111 2873 115 2874
rect 131 2878 135 2879
rect 131 2873 135 2874
rect 171 2878 175 2879
rect 171 2873 175 2874
rect 307 2878 311 2879
rect 307 2873 311 2874
rect 483 2878 487 2879
rect 483 2873 487 2874
rect 523 2878 527 2879
rect 523 2873 527 2874
rect 763 2878 767 2879
rect 763 2873 767 2874
rect 787 2878 791 2879
rect 787 2873 791 2874
rect 1011 2878 1015 2879
rect 1011 2873 1015 2874
rect 1083 2878 1087 2879
rect 1083 2873 1087 2874
rect 1275 2878 1279 2879
rect 1275 2873 1279 2874
rect 1387 2878 1391 2879
rect 1387 2873 1391 2874
rect 1539 2878 1543 2879
rect 1539 2873 1543 2874
rect 1691 2878 1695 2879
rect 1691 2873 1695 2874
rect 1935 2878 1939 2879
rect 1935 2873 1939 2874
rect 112 2813 114 2873
rect 110 2812 116 2813
rect 132 2812 134 2873
rect 308 2812 310 2873
rect 524 2812 526 2873
rect 764 2812 766 2873
rect 1012 2812 1014 2873
rect 1276 2812 1278 2873
rect 1540 2812 1542 2873
rect 1936 2813 1938 2873
rect 1976 2855 1978 2923
rect 2116 2855 2118 2924
rect 2316 2855 2318 2924
rect 2516 2855 2518 2924
rect 2716 2855 2718 2924
rect 2908 2855 2910 2924
rect 3108 2855 3110 2924
rect 3308 2855 3310 2924
rect 3798 2923 3804 2924
rect 3800 2855 3802 2923
rect 3840 2902 3842 2925
rect 3838 2901 3844 2902
rect 3896 2901 3898 2925
rect 4032 2901 4034 2925
rect 4168 2901 4170 2925
rect 4304 2901 4306 2925
rect 4440 2901 4442 2925
rect 4576 2901 4578 2925
rect 5664 2902 5666 2925
rect 5662 2901 5668 2902
rect 3838 2897 3839 2901
rect 3843 2897 3844 2901
rect 3838 2896 3844 2897
rect 3894 2900 3900 2901
rect 3894 2896 3895 2900
rect 3899 2896 3900 2900
rect 3894 2895 3900 2896
rect 4030 2900 4036 2901
rect 4030 2896 4031 2900
rect 4035 2896 4036 2900
rect 4030 2895 4036 2896
rect 4166 2900 4172 2901
rect 4166 2896 4167 2900
rect 4171 2896 4172 2900
rect 4166 2895 4172 2896
rect 4302 2900 4308 2901
rect 4302 2896 4303 2900
rect 4307 2896 4308 2900
rect 4302 2895 4308 2896
rect 4438 2900 4444 2901
rect 4438 2896 4439 2900
rect 4443 2896 4444 2900
rect 4438 2895 4444 2896
rect 4574 2900 4580 2901
rect 4574 2896 4575 2900
rect 4579 2896 4580 2900
rect 5662 2897 5663 2901
rect 5667 2897 5668 2901
rect 5662 2896 5668 2897
rect 4574 2895 4580 2896
rect 3866 2885 3872 2886
rect 3838 2884 3844 2885
rect 3838 2880 3839 2884
rect 3843 2880 3844 2884
rect 3866 2881 3867 2885
rect 3871 2881 3872 2885
rect 3866 2880 3872 2881
rect 4002 2885 4008 2886
rect 4002 2881 4003 2885
rect 4007 2881 4008 2885
rect 4002 2880 4008 2881
rect 4138 2885 4144 2886
rect 4138 2881 4139 2885
rect 4143 2881 4144 2885
rect 4138 2880 4144 2881
rect 4274 2885 4280 2886
rect 4274 2881 4275 2885
rect 4279 2881 4280 2885
rect 4274 2880 4280 2881
rect 4410 2885 4416 2886
rect 4410 2881 4411 2885
rect 4415 2881 4416 2885
rect 4410 2880 4416 2881
rect 4546 2885 4552 2886
rect 4546 2881 4547 2885
rect 4551 2881 4552 2885
rect 4546 2880 4552 2881
rect 5662 2884 5668 2885
rect 5662 2880 5663 2884
rect 5667 2880 5668 2884
rect 3838 2879 3844 2880
rect 1975 2854 1979 2855
rect 1975 2849 1979 2850
rect 2011 2854 2015 2855
rect 2011 2849 2015 2850
rect 2115 2854 2119 2855
rect 2115 2849 2119 2850
rect 2259 2854 2263 2855
rect 2259 2849 2263 2850
rect 2315 2854 2319 2855
rect 2315 2849 2319 2850
rect 2507 2854 2511 2855
rect 2507 2849 2511 2850
rect 2515 2854 2519 2855
rect 2515 2849 2519 2850
rect 2715 2854 2719 2855
rect 2715 2849 2719 2850
rect 2755 2854 2759 2855
rect 2755 2849 2759 2850
rect 2907 2854 2911 2855
rect 2907 2849 2911 2850
rect 3003 2854 3007 2855
rect 3003 2849 3007 2850
rect 3107 2854 3111 2855
rect 3107 2849 3111 2850
rect 3307 2854 3311 2855
rect 3307 2849 3311 2850
rect 3799 2854 3803 2855
rect 3799 2849 3803 2850
rect 1934 2812 1940 2813
rect 110 2808 111 2812
rect 115 2808 116 2812
rect 110 2807 116 2808
rect 130 2811 136 2812
rect 130 2807 131 2811
rect 135 2807 136 2811
rect 130 2806 136 2807
rect 306 2811 312 2812
rect 306 2807 307 2811
rect 311 2807 312 2811
rect 306 2806 312 2807
rect 522 2811 528 2812
rect 522 2807 523 2811
rect 527 2807 528 2811
rect 522 2806 528 2807
rect 762 2811 768 2812
rect 762 2807 763 2811
rect 767 2807 768 2811
rect 762 2806 768 2807
rect 1010 2811 1016 2812
rect 1010 2807 1011 2811
rect 1015 2807 1016 2811
rect 1010 2806 1016 2807
rect 1274 2811 1280 2812
rect 1274 2807 1275 2811
rect 1279 2807 1280 2811
rect 1274 2806 1280 2807
rect 1538 2811 1544 2812
rect 1538 2807 1539 2811
rect 1543 2807 1544 2811
rect 1934 2808 1935 2812
rect 1939 2808 1940 2812
rect 1934 2807 1940 2808
rect 1538 2806 1544 2807
rect 158 2796 164 2797
rect 110 2795 116 2796
rect 110 2791 111 2795
rect 115 2791 116 2795
rect 158 2792 159 2796
rect 163 2792 164 2796
rect 158 2791 164 2792
rect 334 2796 340 2797
rect 334 2792 335 2796
rect 339 2792 340 2796
rect 334 2791 340 2792
rect 550 2796 556 2797
rect 550 2792 551 2796
rect 555 2792 556 2796
rect 550 2791 556 2792
rect 790 2796 796 2797
rect 790 2792 791 2796
rect 795 2792 796 2796
rect 790 2791 796 2792
rect 1038 2796 1044 2797
rect 1038 2792 1039 2796
rect 1043 2792 1044 2796
rect 1038 2791 1044 2792
rect 1302 2796 1308 2797
rect 1302 2792 1303 2796
rect 1307 2792 1308 2796
rect 1302 2791 1308 2792
rect 1566 2796 1572 2797
rect 1566 2792 1567 2796
rect 1571 2792 1572 2796
rect 1566 2791 1572 2792
rect 1934 2795 1940 2796
rect 1934 2791 1935 2795
rect 1939 2791 1940 2795
rect 110 2790 116 2791
rect 112 2763 114 2790
rect 160 2763 162 2791
rect 336 2763 338 2791
rect 552 2763 554 2791
rect 792 2763 794 2791
rect 1040 2763 1042 2791
rect 1304 2763 1306 2791
rect 1568 2763 1570 2791
rect 1934 2790 1940 2791
rect 1936 2763 1938 2790
rect 1976 2789 1978 2849
rect 1974 2788 1980 2789
rect 2012 2788 2014 2849
rect 2260 2788 2262 2849
rect 2508 2788 2510 2849
rect 2756 2788 2758 2849
rect 3004 2788 3006 2849
rect 3800 2789 3802 2849
rect 3840 2811 3842 2879
rect 3868 2811 3870 2880
rect 4004 2811 4006 2880
rect 4140 2811 4142 2880
rect 4276 2811 4278 2880
rect 4412 2811 4414 2880
rect 4548 2811 4550 2880
rect 5662 2879 5668 2880
rect 5664 2811 5666 2879
rect 3839 2810 3843 2811
rect 3839 2805 3843 2806
rect 3859 2810 3863 2811
rect 3859 2805 3863 2806
rect 3867 2810 3871 2811
rect 3867 2805 3871 2806
rect 3995 2810 3999 2811
rect 3995 2805 3999 2806
rect 4003 2810 4007 2811
rect 4003 2805 4007 2806
rect 4131 2810 4135 2811
rect 4131 2805 4135 2806
rect 4139 2810 4143 2811
rect 4139 2805 4143 2806
rect 4267 2810 4271 2811
rect 4267 2805 4271 2806
rect 4275 2810 4279 2811
rect 4275 2805 4279 2806
rect 4403 2810 4407 2811
rect 4403 2805 4407 2806
rect 4411 2810 4415 2811
rect 4411 2805 4415 2806
rect 4539 2810 4543 2811
rect 4539 2805 4543 2806
rect 4547 2810 4551 2811
rect 4547 2805 4551 2806
rect 4675 2810 4679 2811
rect 4675 2805 4679 2806
rect 4811 2810 4815 2811
rect 4811 2805 4815 2806
rect 5663 2810 5667 2811
rect 5663 2805 5667 2806
rect 3798 2788 3804 2789
rect 1974 2784 1975 2788
rect 1979 2784 1980 2788
rect 1974 2783 1980 2784
rect 2010 2787 2016 2788
rect 2010 2783 2011 2787
rect 2015 2783 2016 2787
rect 2010 2782 2016 2783
rect 2258 2787 2264 2788
rect 2258 2783 2259 2787
rect 2263 2783 2264 2787
rect 2258 2782 2264 2783
rect 2506 2787 2512 2788
rect 2506 2783 2507 2787
rect 2511 2783 2512 2787
rect 2506 2782 2512 2783
rect 2754 2787 2760 2788
rect 2754 2783 2755 2787
rect 2759 2783 2760 2787
rect 2754 2782 2760 2783
rect 3002 2787 3008 2788
rect 3002 2783 3003 2787
rect 3007 2783 3008 2787
rect 3798 2784 3799 2788
rect 3803 2784 3804 2788
rect 3798 2783 3804 2784
rect 3002 2782 3008 2783
rect 2038 2772 2044 2773
rect 1974 2771 1980 2772
rect 1974 2767 1975 2771
rect 1979 2767 1980 2771
rect 2038 2768 2039 2772
rect 2043 2768 2044 2772
rect 2038 2767 2044 2768
rect 2286 2772 2292 2773
rect 2286 2768 2287 2772
rect 2291 2768 2292 2772
rect 2286 2767 2292 2768
rect 2534 2772 2540 2773
rect 2534 2768 2535 2772
rect 2539 2768 2540 2772
rect 2534 2767 2540 2768
rect 2782 2772 2788 2773
rect 2782 2768 2783 2772
rect 2787 2768 2788 2772
rect 2782 2767 2788 2768
rect 3030 2772 3036 2773
rect 3030 2768 3031 2772
rect 3035 2768 3036 2772
rect 3030 2767 3036 2768
rect 3798 2771 3804 2772
rect 3798 2767 3799 2771
rect 3803 2767 3804 2771
rect 1974 2766 1980 2767
rect 111 2762 115 2763
rect 111 2757 115 2758
rect 159 2762 163 2763
rect 159 2757 163 2758
rect 279 2762 283 2763
rect 279 2757 283 2758
rect 335 2762 339 2763
rect 335 2757 339 2758
rect 455 2762 459 2763
rect 455 2757 459 2758
rect 551 2762 555 2763
rect 551 2757 555 2758
rect 647 2762 651 2763
rect 647 2757 651 2758
rect 791 2762 795 2763
rect 791 2757 795 2758
rect 855 2762 859 2763
rect 855 2757 859 2758
rect 1039 2762 1043 2763
rect 1039 2757 1043 2758
rect 1079 2762 1083 2763
rect 1079 2757 1083 2758
rect 1303 2762 1307 2763
rect 1303 2757 1307 2758
rect 1311 2762 1315 2763
rect 1311 2757 1315 2758
rect 1551 2762 1555 2763
rect 1551 2757 1555 2758
rect 1567 2762 1571 2763
rect 1567 2757 1571 2758
rect 1799 2762 1803 2763
rect 1799 2757 1803 2758
rect 1935 2762 1939 2763
rect 1935 2757 1939 2758
rect 112 2734 114 2757
rect 110 2733 116 2734
rect 280 2733 282 2757
rect 456 2733 458 2757
rect 648 2733 650 2757
rect 856 2733 858 2757
rect 1080 2733 1082 2757
rect 1312 2733 1314 2757
rect 1552 2733 1554 2757
rect 1800 2733 1802 2757
rect 1936 2734 1938 2757
rect 1976 2739 1978 2766
rect 2040 2739 2042 2767
rect 2288 2739 2290 2767
rect 2536 2739 2538 2767
rect 2784 2739 2786 2767
rect 3032 2739 3034 2767
rect 3798 2766 3804 2767
rect 3800 2739 3802 2766
rect 3840 2745 3842 2805
rect 3838 2744 3844 2745
rect 3860 2744 3862 2805
rect 3996 2744 3998 2805
rect 4132 2744 4134 2805
rect 4268 2744 4270 2805
rect 4404 2744 4406 2805
rect 4540 2744 4542 2805
rect 4676 2744 4678 2805
rect 4812 2744 4814 2805
rect 5664 2745 5666 2805
rect 5662 2744 5668 2745
rect 3838 2740 3839 2744
rect 3843 2740 3844 2744
rect 3838 2739 3844 2740
rect 3858 2743 3864 2744
rect 3858 2739 3859 2743
rect 3863 2739 3864 2743
rect 1975 2738 1979 2739
rect 1934 2733 1940 2734
rect 1975 2733 1979 2734
rect 2023 2738 2027 2739
rect 2023 2733 2027 2734
rect 2039 2738 2043 2739
rect 2039 2733 2043 2734
rect 2247 2738 2251 2739
rect 2247 2733 2251 2734
rect 2287 2738 2291 2739
rect 2287 2733 2291 2734
rect 2503 2738 2507 2739
rect 2503 2733 2507 2734
rect 2535 2738 2539 2739
rect 2535 2733 2539 2734
rect 2759 2738 2763 2739
rect 2759 2733 2763 2734
rect 2783 2738 2787 2739
rect 2783 2733 2787 2734
rect 3015 2738 3019 2739
rect 3015 2733 3019 2734
rect 3031 2738 3035 2739
rect 3031 2733 3035 2734
rect 3799 2738 3803 2739
rect 3858 2738 3864 2739
rect 3994 2743 4000 2744
rect 3994 2739 3995 2743
rect 3999 2739 4000 2743
rect 3994 2738 4000 2739
rect 4130 2743 4136 2744
rect 4130 2739 4131 2743
rect 4135 2739 4136 2743
rect 4130 2738 4136 2739
rect 4266 2743 4272 2744
rect 4266 2739 4267 2743
rect 4271 2739 4272 2743
rect 4266 2738 4272 2739
rect 4402 2743 4408 2744
rect 4402 2739 4403 2743
rect 4407 2739 4408 2743
rect 4402 2738 4408 2739
rect 4538 2743 4544 2744
rect 4538 2739 4539 2743
rect 4543 2739 4544 2743
rect 4538 2738 4544 2739
rect 4674 2743 4680 2744
rect 4674 2739 4675 2743
rect 4679 2739 4680 2743
rect 4674 2738 4680 2739
rect 4810 2743 4816 2744
rect 4810 2739 4811 2743
rect 4815 2739 4816 2743
rect 5662 2740 5663 2744
rect 5667 2740 5668 2744
rect 5662 2739 5668 2740
rect 4810 2738 4816 2739
rect 3799 2733 3803 2734
rect 110 2729 111 2733
rect 115 2729 116 2733
rect 110 2728 116 2729
rect 278 2732 284 2733
rect 278 2728 279 2732
rect 283 2728 284 2732
rect 278 2727 284 2728
rect 454 2732 460 2733
rect 454 2728 455 2732
rect 459 2728 460 2732
rect 454 2727 460 2728
rect 646 2732 652 2733
rect 646 2728 647 2732
rect 651 2728 652 2732
rect 646 2727 652 2728
rect 854 2732 860 2733
rect 854 2728 855 2732
rect 859 2728 860 2732
rect 854 2727 860 2728
rect 1078 2732 1084 2733
rect 1078 2728 1079 2732
rect 1083 2728 1084 2732
rect 1078 2727 1084 2728
rect 1310 2732 1316 2733
rect 1310 2728 1311 2732
rect 1315 2728 1316 2732
rect 1310 2727 1316 2728
rect 1550 2732 1556 2733
rect 1550 2728 1551 2732
rect 1555 2728 1556 2732
rect 1550 2727 1556 2728
rect 1798 2732 1804 2733
rect 1798 2728 1799 2732
rect 1803 2728 1804 2732
rect 1934 2729 1935 2733
rect 1939 2729 1940 2733
rect 1934 2728 1940 2729
rect 1798 2727 1804 2728
rect 250 2717 256 2718
rect 110 2716 116 2717
rect 110 2712 111 2716
rect 115 2712 116 2716
rect 250 2713 251 2717
rect 255 2713 256 2717
rect 250 2712 256 2713
rect 426 2717 432 2718
rect 426 2713 427 2717
rect 431 2713 432 2717
rect 426 2712 432 2713
rect 618 2717 624 2718
rect 618 2713 619 2717
rect 623 2713 624 2717
rect 618 2712 624 2713
rect 826 2717 832 2718
rect 826 2713 827 2717
rect 831 2713 832 2717
rect 826 2712 832 2713
rect 1050 2717 1056 2718
rect 1050 2713 1051 2717
rect 1055 2713 1056 2717
rect 1050 2712 1056 2713
rect 1282 2717 1288 2718
rect 1282 2713 1283 2717
rect 1287 2713 1288 2717
rect 1282 2712 1288 2713
rect 1522 2717 1528 2718
rect 1522 2713 1523 2717
rect 1527 2713 1528 2717
rect 1522 2712 1528 2713
rect 1770 2717 1776 2718
rect 1770 2713 1771 2717
rect 1775 2713 1776 2717
rect 1770 2712 1776 2713
rect 1934 2716 1940 2717
rect 1934 2712 1935 2716
rect 1939 2712 1940 2716
rect 110 2711 116 2712
rect 112 2651 114 2711
rect 252 2651 254 2712
rect 428 2651 430 2712
rect 620 2651 622 2712
rect 828 2651 830 2712
rect 1052 2651 1054 2712
rect 1284 2651 1286 2712
rect 1524 2651 1526 2712
rect 1772 2651 1774 2712
rect 1934 2711 1940 2712
rect 1936 2651 1938 2711
rect 1976 2710 1978 2733
rect 1974 2709 1980 2710
rect 2024 2709 2026 2733
rect 2248 2709 2250 2733
rect 2504 2709 2506 2733
rect 2760 2709 2762 2733
rect 3016 2709 3018 2733
rect 3800 2710 3802 2733
rect 3886 2728 3892 2729
rect 3838 2727 3844 2728
rect 3838 2723 3839 2727
rect 3843 2723 3844 2727
rect 3886 2724 3887 2728
rect 3891 2724 3892 2728
rect 3886 2723 3892 2724
rect 4022 2728 4028 2729
rect 4022 2724 4023 2728
rect 4027 2724 4028 2728
rect 4022 2723 4028 2724
rect 4158 2728 4164 2729
rect 4158 2724 4159 2728
rect 4163 2724 4164 2728
rect 4158 2723 4164 2724
rect 4294 2728 4300 2729
rect 4294 2724 4295 2728
rect 4299 2724 4300 2728
rect 4294 2723 4300 2724
rect 4430 2728 4436 2729
rect 4430 2724 4431 2728
rect 4435 2724 4436 2728
rect 4430 2723 4436 2724
rect 4566 2728 4572 2729
rect 4566 2724 4567 2728
rect 4571 2724 4572 2728
rect 4566 2723 4572 2724
rect 4702 2728 4708 2729
rect 4702 2724 4703 2728
rect 4707 2724 4708 2728
rect 4702 2723 4708 2724
rect 4838 2728 4844 2729
rect 4838 2724 4839 2728
rect 4843 2724 4844 2728
rect 4838 2723 4844 2724
rect 5662 2727 5668 2728
rect 5662 2723 5663 2727
rect 5667 2723 5668 2727
rect 3838 2722 3844 2723
rect 3798 2709 3804 2710
rect 1974 2705 1975 2709
rect 1979 2705 1980 2709
rect 1974 2704 1980 2705
rect 2022 2708 2028 2709
rect 2022 2704 2023 2708
rect 2027 2704 2028 2708
rect 2022 2703 2028 2704
rect 2246 2708 2252 2709
rect 2246 2704 2247 2708
rect 2251 2704 2252 2708
rect 2246 2703 2252 2704
rect 2502 2708 2508 2709
rect 2502 2704 2503 2708
rect 2507 2704 2508 2708
rect 2502 2703 2508 2704
rect 2758 2708 2764 2709
rect 2758 2704 2759 2708
rect 2763 2704 2764 2708
rect 2758 2703 2764 2704
rect 3014 2708 3020 2709
rect 3014 2704 3015 2708
rect 3019 2704 3020 2708
rect 3798 2705 3799 2709
rect 3803 2705 3804 2709
rect 3798 2704 3804 2705
rect 3014 2703 3020 2704
rect 3840 2699 3842 2722
rect 3888 2699 3890 2723
rect 4024 2699 4026 2723
rect 4160 2699 4162 2723
rect 4296 2699 4298 2723
rect 4432 2699 4434 2723
rect 4568 2699 4570 2723
rect 4704 2699 4706 2723
rect 4840 2699 4842 2723
rect 5662 2722 5668 2723
rect 5664 2699 5666 2722
rect 3839 2698 3843 2699
rect 1994 2693 2000 2694
rect 1974 2692 1980 2693
rect 1974 2688 1975 2692
rect 1979 2688 1980 2692
rect 1994 2689 1995 2693
rect 1999 2689 2000 2693
rect 1994 2688 2000 2689
rect 2218 2693 2224 2694
rect 2218 2689 2219 2693
rect 2223 2689 2224 2693
rect 2218 2688 2224 2689
rect 2474 2693 2480 2694
rect 2474 2689 2475 2693
rect 2479 2689 2480 2693
rect 2474 2688 2480 2689
rect 2730 2693 2736 2694
rect 2730 2689 2731 2693
rect 2735 2689 2736 2693
rect 2730 2688 2736 2689
rect 2986 2693 2992 2694
rect 3839 2693 3843 2694
rect 3887 2698 3891 2699
rect 3887 2693 3891 2694
rect 3959 2698 3963 2699
rect 3959 2693 3963 2694
rect 4023 2698 4027 2699
rect 4023 2693 4027 2694
rect 4159 2698 4163 2699
rect 4159 2693 4163 2694
rect 4255 2698 4259 2699
rect 4255 2693 4259 2694
rect 4295 2698 4299 2699
rect 4295 2693 4299 2694
rect 4431 2698 4435 2699
rect 4431 2693 4435 2694
rect 4543 2698 4547 2699
rect 4543 2693 4547 2694
rect 4567 2698 4571 2699
rect 4567 2693 4571 2694
rect 4703 2698 4707 2699
rect 4703 2693 4707 2694
rect 4823 2698 4827 2699
rect 4823 2693 4827 2694
rect 4839 2698 4843 2699
rect 4839 2693 4843 2694
rect 5111 2698 5115 2699
rect 5111 2693 5115 2694
rect 5399 2698 5403 2699
rect 5399 2693 5403 2694
rect 5663 2698 5667 2699
rect 5663 2693 5667 2694
rect 2986 2689 2987 2693
rect 2991 2689 2992 2693
rect 2986 2688 2992 2689
rect 3798 2692 3804 2693
rect 3798 2688 3799 2692
rect 3803 2688 3804 2692
rect 1974 2687 1980 2688
rect 111 2650 115 2651
rect 111 2645 115 2646
rect 251 2650 255 2651
rect 251 2645 255 2646
rect 427 2650 431 2651
rect 427 2645 431 2646
rect 571 2650 575 2651
rect 571 2645 575 2646
rect 619 2650 623 2651
rect 619 2645 623 2646
rect 731 2650 735 2651
rect 731 2645 735 2646
rect 827 2650 831 2651
rect 827 2645 831 2646
rect 891 2650 895 2651
rect 891 2645 895 2646
rect 1043 2650 1047 2651
rect 1043 2645 1047 2646
rect 1051 2650 1055 2651
rect 1051 2645 1055 2646
rect 1195 2650 1199 2651
rect 1195 2645 1199 2646
rect 1283 2650 1287 2651
rect 1283 2645 1287 2646
rect 1355 2650 1359 2651
rect 1355 2645 1359 2646
rect 1515 2650 1519 2651
rect 1515 2645 1519 2646
rect 1523 2650 1527 2651
rect 1523 2645 1527 2646
rect 1675 2650 1679 2651
rect 1675 2645 1679 2646
rect 1771 2650 1775 2651
rect 1771 2645 1775 2646
rect 1935 2650 1939 2651
rect 1935 2645 1939 2646
rect 112 2585 114 2645
rect 110 2584 116 2585
rect 572 2584 574 2645
rect 732 2584 734 2645
rect 892 2584 894 2645
rect 1044 2584 1046 2645
rect 1196 2584 1198 2645
rect 1356 2584 1358 2645
rect 1516 2584 1518 2645
rect 1676 2584 1678 2645
rect 1936 2585 1938 2645
rect 1976 2615 1978 2687
rect 1996 2615 1998 2688
rect 2220 2615 2222 2688
rect 2476 2615 2478 2688
rect 2732 2615 2734 2688
rect 2988 2615 2990 2688
rect 3798 2687 3804 2688
rect 3800 2615 3802 2687
rect 3840 2670 3842 2693
rect 3838 2669 3844 2670
rect 3960 2669 3962 2693
rect 4256 2669 4258 2693
rect 4544 2669 4546 2693
rect 4824 2669 4826 2693
rect 5112 2669 5114 2693
rect 5400 2669 5402 2693
rect 5664 2670 5666 2693
rect 5662 2669 5668 2670
rect 3838 2665 3839 2669
rect 3843 2665 3844 2669
rect 3838 2664 3844 2665
rect 3958 2668 3964 2669
rect 3958 2664 3959 2668
rect 3963 2664 3964 2668
rect 3958 2663 3964 2664
rect 4254 2668 4260 2669
rect 4254 2664 4255 2668
rect 4259 2664 4260 2668
rect 4254 2663 4260 2664
rect 4542 2668 4548 2669
rect 4542 2664 4543 2668
rect 4547 2664 4548 2668
rect 4542 2663 4548 2664
rect 4822 2668 4828 2669
rect 4822 2664 4823 2668
rect 4827 2664 4828 2668
rect 4822 2663 4828 2664
rect 5110 2668 5116 2669
rect 5110 2664 5111 2668
rect 5115 2664 5116 2668
rect 5110 2663 5116 2664
rect 5398 2668 5404 2669
rect 5398 2664 5399 2668
rect 5403 2664 5404 2668
rect 5662 2665 5663 2669
rect 5667 2665 5668 2669
rect 5662 2664 5668 2665
rect 5398 2663 5404 2664
rect 3930 2653 3936 2654
rect 3838 2652 3844 2653
rect 3838 2648 3839 2652
rect 3843 2648 3844 2652
rect 3930 2649 3931 2653
rect 3935 2649 3936 2653
rect 3930 2648 3936 2649
rect 4226 2653 4232 2654
rect 4226 2649 4227 2653
rect 4231 2649 4232 2653
rect 4226 2648 4232 2649
rect 4514 2653 4520 2654
rect 4514 2649 4515 2653
rect 4519 2649 4520 2653
rect 4514 2648 4520 2649
rect 4794 2653 4800 2654
rect 4794 2649 4795 2653
rect 4799 2649 4800 2653
rect 4794 2648 4800 2649
rect 5082 2653 5088 2654
rect 5082 2649 5083 2653
rect 5087 2649 5088 2653
rect 5082 2648 5088 2649
rect 5370 2653 5376 2654
rect 5370 2649 5371 2653
rect 5375 2649 5376 2653
rect 5370 2648 5376 2649
rect 5662 2652 5668 2653
rect 5662 2648 5663 2652
rect 5667 2648 5668 2652
rect 3838 2647 3844 2648
rect 1975 2614 1979 2615
rect 1975 2609 1979 2610
rect 1995 2614 1999 2615
rect 1995 2609 1999 2610
rect 2219 2614 2223 2615
rect 2219 2609 2223 2610
rect 2475 2614 2479 2615
rect 2475 2609 2479 2610
rect 2555 2614 2559 2615
rect 2555 2609 2559 2610
rect 2691 2614 2695 2615
rect 2691 2609 2695 2610
rect 2731 2614 2735 2615
rect 2731 2609 2735 2610
rect 2827 2614 2831 2615
rect 2827 2609 2831 2610
rect 2963 2614 2967 2615
rect 2963 2609 2967 2610
rect 2987 2614 2991 2615
rect 2987 2609 2991 2610
rect 3099 2614 3103 2615
rect 3099 2609 3103 2610
rect 3799 2614 3803 2615
rect 3799 2609 3803 2610
rect 1934 2584 1940 2585
rect 110 2580 111 2584
rect 115 2580 116 2584
rect 110 2579 116 2580
rect 570 2583 576 2584
rect 570 2579 571 2583
rect 575 2579 576 2583
rect 570 2578 576 2579
rect 730 2583 736 2584
rect 730 2579 731 2583
rect 735 2579 736 2583
rect 730 2578 736 2579
rect 890 2583 896 2584
rect 890 2579 891 2583
rect 895 2579 896 2583
rect 890 2578 896 2579
rect 1042 2583 1048 2584
rect 1042 2579 1043 2583
rect 1047 2579 1048 2583
rect 1042 2578 1048 2579
rect 1194 2583 1200 2584
rect 1194 2579 1195 2583
rect 1199 2579 1200 2583
rect 1194 2578 1200 2579
rect 1354 2583 1360 2584
rect 1354 2579 1355 2583
rect 1359 2579 1360 2583
rect 1354 2578 1360 2579
rect 1514 2583 1520 2584
rect 1514 2579 1515 2583
rect 1519 2579 1520 2583
rect 1514 2578 1520 2579
rect 1674 2583 1680 2584
rect 1674 2579 1675 2583
rect 1679 2579 1680 2583
rect 1934 2580 1935 2584
rect 1939 2580 1940 2584
rect 1934 2579 1940 2580
rect 1674 2578 1680 2579
rect 598 2568 604 2569
rect 110 2567 116 2568
rect 110 2563 111 2567
rect 115 2563 116 2567
rect 598 2564 599 2568
rect 603 2564 604 2568
rect 598 2563 604 2564
rect 758 2568 764 2569
rect 758 2564 759 2568
rect 763 2564 764 2568
rect 758 2563 764 2564
rect 918 2568 924 2569
rect 918 2564 919 2568
rect 923 2564 924 2568
rect 918 2563 924 2564
rect 1070 2568 1076 2569
rect 1070 2564 1071 2568
rect 1075 2564 1076 2568
rect 1070 2563 1076 2564
rect 1222 2568 1228 2569
rect 1222 2564 1223 2568
rect 1227 2564 1228 2568
rect 1222 2563 1228 2564
rect 1382 2568 1388 2569
rect 1382 2564 1383 2568
rect 1387 2564 1388 2568
rect 1382 2563 1388 2564
rect 1542 2568 1548 2569
rect 1542 2564 1543 2568
rect 1547 2564 1548 2568
rect 1542 2563 1548 2564
rect 1702 2568 1708 2569
rect 1702 2564 1703 2568
rect 1707 2564 1708 2568
rect 1702 2563 1708 2564
rect 1934 2567 1940 2568
rect 1934 2563 1935 2567
rect 1939 2563 1940 2567
rect 110 2562 116 2563
rect 112 2539 114 2562
rect 600 2539 602 2563
rect 760 2539 762 2563
rect 920 2539 922 2563
rect 1072 2539 1074 2563
rect 1224 2539 1226 2563
rect 1384 2539 1386 2563
rect 1544 2539 1546 2563
rect 1704 2539 1706 2563
rect 1934 2562 1940 2563
rect 1936 2539 1938 2562
rect 1976 2549 1978 2609
rect 1974 2548 1980 2549
rect 2556 2548 2558 2609
rect 2692 2548 2694 2609
rect 2828 2548 2830 2609
rect 2964 2548 2966 2609
rect 3100 2548 3102 2609
rect 3800 2549 3802 2609
rect 3840 2587 3842 2647
rect 3932 2587 3934 2648
rect 4228 2587 4230 2648
rect 4516 2587 4518 2648
rect 4796 2587 4798 2648
rect 5084 2587 5086 2648
rect 5372 2587 5374 2648
rect 5662 2647 5668 2648
rect 5664 2587 5666 2647
rect 3839 2586 3843 2587
rect 3839 2581 3843 2582
rect 3859 2586 3863 2587
rect 3859 2581 3863 2582
rect 3931 2586 3935 2587
rect 3931 2581 3935 2582
rect 4083 2586 4087 2587
rect 4083 2581 4087 2582
rect 4227 2586 4231 2587
rect 4227 2581 4231 2582
rect 4331 2586 4335 2587
rect 4331 2581 4335 2582
rect 4515 2586 4519 2587
rect 4515 2581 4519 2582
rect 4579 2586 4583 2587
rect 4579 2581 4583 2582
rect 4795 2586 4799 2587
rect 4795 2581 4799 2582
rect 4827 2586 4831 2587
rect 4827 2581 4831 2582
rect 5075 2586 5079 2587
rect 5075 2581 5079 2582
rect 5083 2586 5087 2587
rect 5083 2581 5087 2582
rect 5323 2586 5327 2587
rect 5323 2581 5327 2582
rect 5371 2586 5375 2587
rect 5371 2581 5375 2582
rect 5663 2586 5667 2587
rect 5663 2581 5667 2582
rect 3798 2548 3804 2549
rect 1974 2544 1975 2548
rect 1979 2544 1980 2548
rect 1974 2543 1980 2544
rect 2554 2547 2560 2548
rect 2554 2543 2555 2547
rect 2559 2543 2560 2547
rect 2554 2542 2560 2543
rect 2690 2547 2696 2548
rect 2690 2543 2691 2547
rect 2695 2543 2696 2547
rect 2690 2542 2696 2543
rect 2826 2547 2832 2548
rect 2826 2543 2827 2547
rect 2831 2543 2832 2547
rect 2826 2542 2832 2543
rect 2962 2547 2968 2548
rect 2962 2543 2963 2547
rect 2967 2543 2968 2547
rect 2962 2542 2968 2543
rect 3098 2547 3104 2548
rect 3098 2543 3099 2547
rect 3103 2543 3104 2547
rect 3798 2544 3799 2548
rect 3803 2544 3804 2548
rect 3798 2543 3804 2544
rect 3098 2542 3104 2543
rect 111 2538 115 2539
rect 111 2533 115 2534
rect 383 2538 387 2539
rect 383 2533 387 2534
rect 599 2538 603 2539
rect 599 2533 603 2534
rect 759 2538 763 2539
rect 759 2533 763 2534
rect 815 2538 819 2539
rect 815 2533 819 2534
rect 919 2538 923 2539
rect 919 2533 923 2534
rect 1023 2538 1027 2539
rect 1023 2533 1027 2534
rect 1071 2538 1075 2539
rect 1071 2533 1075 2534
rect 1223 2538 1227 2539
rect 1223 2533 1227 2534
rect 1231 2538 1235 2539
rect 1231 2533 1235 2534
rect 1383 2538 1387 2539
rect 1383 2533 1387 2534
rect 1431 2538 1435 2539
rect 1431 2533 1435 2534
rect 1543 2538 1547 2539
rect 1543 2533 1547 2534
rect 1631 2538 1635 2539
rect 1631 2533 1635 2534
rect 1703 2538 1707 2539
rect 1703 2533 1707 2534
rect 1815 2538 1819 2539
rect 1815 2533 1819 2534
rect 1935 2538 1939 2539
rect 1935 2533 1939 2534
rect 112 2510 114 2533
rect 110 2509 116 2510
rect 384 2509 386 2533
rect 600 2509 602 2533
rect 816 2509 818 2533
rect 1024 2509 1026 2533
rect 1232 2509 1234 2533
rect 1432 2509 1434 2533
rect 1632 2509 1634 2533
rect 1816 2509 1818 2533
rect 1936 2510 1938 2533
rect 2582 2532 2588 2533
rect 1974 2531 1980 2532
rect 1974 2527 1975 2531
rect 1979 2527 1980 2531
rect 2582 2528 2583 2532
rect 2587 2528 2588 2532
rect 2582 2527 2588 2528
rect 2718 2532 2724 2533
rect 2718 2528 2719 2532
rect 2723 2528 2724 2532
rect 2718 2527 2724 2528
rect 2854 2532 2860 2533
rect 2854 2528 2855 2532
rect 2859 2528 2860 2532
rect 2854 2527 2860 2528
rect 2990 2532 2996 2533
rect 2990 2528 2991 2532
rect 2995 2528 2996 2532
rect 2990 2527 2996 2528
rect 3126 2532 3132 2533
rect 3126 2528 3127 2532
rect 3131 2528 3132 2532
rect 3126 2527 3132 2528
rect 3798 2531 3804 2532
rect 3798 2527 3799 2531
rect 3803 2527 3804 2531
rect 1974 2526 1980 2527
rect 1934 2509 1940 2510
rect 110 2505 111 2509
rect 115 2505 116 2509
rect 110 2504 116 2505
rect 382 2508 388 2509
rect 382 2504 383 2508
rect 387 2504 388 2508
rect 382 2503 388 2504
rect 598 2508 604 2509
rect 598 2504 599 2508
rect 603 2504 604 2508
rect 598 2503 604 2504
rect 814 2508 820 2509
rect 814 2504 815 2508
rect 819 2504 820 2508
rect 814 2503 820 2504
rect 1022 2508 1028 2509
rect 1022 2504 1023 2508
rect 1027 2504 1028 2508
rect 1022 2503 1028 2504
rect 1230 2508 1236 2509
rect 1230 2504 1231 2508
rect 1235 2504 1236 2508
rect 1230 2503 1236 2504
rect 1430 2508 1436 2509
rect 1430 2504 1431 2508
rect 1435 2504 1436 2508
rect 1430 2503 1436 2504
rect 1630 2508 1636 2509
rect 1630 2504 1631 2508
rect 1635 2504 1636 2508
rect 1630 2503 1636 2504
rect 1814 2508 1820 2509
rect 1814 2504 1815 2508
rect 1819 2504 1820 2508
rect 1934 2505 1935 2509
rect 1939 2505 1940 2509
rect 1934 2504 1940 2505
rect 1814 2503 1820 2504
rect 354 2493 360 2494
rect 110 2492 116 2493
rect 110 2488 111 2492
rect 115 2488 116 2492
rect 354 2489 355 2493
rect 359 2489 360 2493
rect 354 2488 360 2489
rect 570 2493 576 2494
rect 570 2489 571 2493
rect 575 2489 576 2493
rect 570 2488 576 2489
rect 786 2493 792 2494
rect 786 2489 787 2493
rect 791 2489 792 2493
rect 786 2488 792 2489
rect 994 2493 1000 2494
rect 994 2489 995 2493
rect 999 2489 1000 2493
rect 994 2488 1000 2489
rect 1202 2493 1208 2494
rect 1202 2489 1203 2493
rect 1207 2489 1208 2493
rect 1202 2488 1208 2489
rect 1402 2493 1408 2494
rect 1402 2489 1403 2493
rect 1407 2489 1408 2493
rect 1402 2488 1408 2489
rect 1602 2493 1608 2494
rect 1602 2489 1603 2493
rect 1607 2489 1608 2493
rect 1602 2488 1608 2489
rect 1786 2493 1792 2494
rect 1786 2489 1787 2493
rect 1791 2489 1792 2493
rect 1786 2488 1792 2489
rect 1934 2492 1940 2493
rect 1934 2488 1935 2492
rect 1939 2488 1940 2492
rect 110 2487 116 2488
rect 112 2423 114 2487
rect 356 2423 358 2488
rect 572 2423 574 2488
rect 788 2423 790 2488
rect 996 2423 998 2488
rect 1204 2423 1206 2488
rect 1404 2423 1406 2488
rect 1604 2423 1606 2488
rect 1788 2423 1790 2488
rect 1934 2487 1940 2488
rect 1936 2423 1938 2487
rect 1976 2479 1978 2526
rect 2584 2479 2586 2527
rect 2720 2479 2722 2527
rect 2856 2479 2858 2527
rect 2992 2479 2994 2527
rect 3128 2479 3130 2527
rect 3798 2526 3804 2527
rect 3800 2479 3802 2526
rect 3840 2521 3842 2581
rect 3838 2520 3844 2521
rect 3860 2520 3862 2581
rect 4084 2520 4086 2581
rect 4332 2520 4334 2581
rect 4580 2520 4582 2581
rect 4828 2520 4830 2581
rect 5076 2520 5078 2581
rect 5324 2520 5326 2581
rect 5664 2521 5666 2581
rect 5662 2520 5668 2521
rect 3838 2516 3839 2520
rect 3843 2516 3844 2520
rect 3838 2515 3844 2516
rect 3858 2519 3864 2520
rect 3858 2515 3859 2519
rect 3863 2515 3864 2519
rect 3858 2514 3864 2515
rect 4082 2519 4088 2520
rect 4082 2515 4083 2519
rect 4087 2515 4088 2519
rect 4082 2514 4088 2515
rect 4330 2519 4336 2520
rect 4330 2515 4331 2519
rect 4335 2515 4336 2519
rect 4330 2514 4336 2515
rect 4578 2519 4584 2520
rect 4578 2515 4579 2519
rect 4583 2515 4584 2519
rect 4578 2514 4584 2515
rect 4826 2519 4832 2520
rect 4826 2515 4827 2519
rect 4831 2515 4832 2519
rect 4826 2514 4832 2515
rect 5074 2519 5080 2520
rect 5074 2515 5075 2519
rect 5079 2515 5080 2519
rect 5074 2514 5080 2515
rect 5322 2519 5328 2520
rect 5322 2515 5323 2519
rect 5327 2515 5328 2519
rect 5662 2516 5663 2520
rect 5667 2516 5668 2520
rect 5662 2515 5668 2516
rect 5322 2514 5328 2515
rect 3886 2504 3892 2505
rect 3838 2503 3844 2504
rect 3838 2499 3839 2503
rect 3843 2499 3844 2503
rect 3886 2500 3887 2504
rect 3891 2500 3892 2504
rect 3886 2499 3892 2500
rect 4110 2504 4116 2505
rect 4110 2500 4111 2504
rect 4115 2500 4116 2504
rect 4110 2499 4116 2500
rect 4358 2504 4364 2505
rect 4358 2500 4359 2504
rect 4363 2500 4364 2504
rect 4358 2499 4364 2500
rect 4606 2504 4612 2505
rect 4606 2500 4607 2504
rect 4611 2500 4612 2504
rect 4606 2499 4612 2500
rect 4854 2504 4860 2505
rect 4854 2500 4855 2504
rect 4859 2500 4860 2504
rect 4854 2499 4860 2500
rect 5102 2504 5108 2505
rect 5102 2500 5103 2504
rect 5107 2500 5108 2504
rect 5102 2499 5108 2500
rect 5350 2504 5356 2505
rect 5350 2500 5351 2504
rect 5355 2500 5356 2504
rect 5350 2499 5356 2500
rect 5662 2503 5668 2504
rect 5662 2499 5663 2503
rect 5667 2499 5668 2503
rect 3838 2498 3844 2499
rect 1975 2478 1979 2479
rect 1975 2473 1979 2474
rect 2023 2478 2027 2479
rect 2023 2473 2027 2474
rect 2223 2478 2227 2479
rect 2223 2473 2227 2474
rect 2447 2478 2451 2479
rect 2447 2473 2451 2474
rect 2583 2478 2587 2479
rect 2583 2473 2587 2474
rect 2679 2478 2683 2479
rect 2679 2473 2683 2474
rect 2719 2478 2723 2479
rect 2719 2473 2723 2474
rect 2855 2478 2859 2479
rect 2855 2473 2859 2474
rect 2927 2478 2931 2479
rect 2927 2473 2931 2474
rect 2991 2478 2995 2479
rect 2991 2473 2995 2474
rect 3127 2478 3131 2479
rect 3127 2473 3131 2474
rect 3183 2478 3187 2479
rect 3183 2473 3187 2474
rect 3439 2478 3443 2479
rect 3439 2473 3443 2474
rect 3679 2478 3683 2479
rect 3679 2473 3683 2474
rect 3799 2478 3803 2479
rect 3799 2473 3803 2474
rect 1976 2450 1978 2473
rect 1974 2449 1980 2450
rect 2024 2449 2026 2473
rect 2224 2449 2226 2473
rect 2448 2449 2450 2473
rect 2680 2449 2682 2473
rect 2928 2449 2930 2473
rect 3184 2449 3186 2473
rect 3440 2449 3442 2473
rect 3680 2449 3682 2473
rect 3800 2450 3802 2473
rect 3840 2471 3842 2498
rect 3888 2471 3890 2499
rect 4112 2471 4114 2499
rect 4360 2471 4362 2499
rect 4608 2471 4610 2499
rect 4856 2471 4858 2499
rect 5104 2471 5106 2499
rect 5352 2471 5354 2499
rect 5662 2498 5668 2499
rect 5664 2471 5666 2498
rect 3839 2470 3843 2471
rect 3839 2465 3843 2466
rect 3887 2470 3891 2471
rect 3887 2465 3891 2466
rect 4087 2470 4091 2471
rect 4087 2465 4091 2466
rect 4111 2470 4115 2471
rect 4111 2465 4115 2466
rect 4327 2470 4331 2471
rect 4327 2465 4331 2466
rect 4359 2470 4363 2471
rect 4359 2465 4363 2466
rect 4583 2470 4587 2471
rect 4583 2465 4587 2466
rect 4607 2470 4611 2471
rect 4607 2465 4611 2466
rect 4847 2470 4851 2471
rect 4847 2465 4851 2466
rect 4855 2470 4859 2471
rect 4855 2465 4859 2466
rect 5103 2470 5107 2471
rect 5103 2465 5107 2466
rect 5119 2470 5123 2471
rect 5119 2465 5123 2466
rect 5351 2470 5355 2471
rect 5351 2465 5355 2466
rect 5399 2470 5403 2471
rect 5399 2465 5403 2466
rect 5663 2470 5667 2471
rect 5663 2465 5667 2466
rect 3798 2449 3804 2450
rect 1974 2445 1975 2449
rect 1979 2445 1980 2449
rect 1974 2444 1980 2445
rect 2022 2448 2028 2449
rect 2022 2444 2023 2448
rect 2027 2444 2028 2448
rect 2022 2443 2028 2444
rect 2222 2448 2228 2449
rect 2222 2444 2223 2448
rect 2227 2444 2228 2448
rect 2222 2443 2228 2444
rect 2446 2448 2452 2449
rect 2446 2444 2447 2448
rect 2451 2444 2452 2448
rect 2446 2443 2452 2444
rect 2678 2448 2684 2449
rect 2678 2444 2679 2448
rect 2683 2444 2684 2448
rect 2678 2443 2684 2444
rect 2926 2448 2932 2449
rect 2926 2444 2927 2448
rect 2931 2444 2932 2448
rect 2926 2443 2932 2444
rect 3182 2448 3188 2449
rect 3182 2444 3183 2448
rect 3187 2444 3188 2448
rect 3182 2443 3188 2444
rect 3438 2448 3444 2449
rect 3438 2444 3439 2448
rect 3443 2444 3444 2448
rect 3438 2443 3444 2444
rect 3678 2448 3684 2449
rect 3678 2444 3679 2448
rect 3683 2444 3684 2448
rect 3798 2445 3799 2449
rect 3803 2445 3804 2449
rect 3798 2444 3804 2445
rect 3678 2443 3684 2444
rect 3840 2442 3842 2465
rect 3838 2441 3844 2442
rect 3888 2441 3890 2465
rect 4088 2441 4090 2465
rect 4328 2441 4330 2465
rect 4584 2441 4586 2465
rect 4848 2441 4850 2465
rect 5120 2441 5122 2465
rect 5400 2441 5402 2465
rect 5664 2442 5666 2465
rect 5662 2441 5668 2442
rect 3838 2437 3839 2441
rect 3843 2437 3844 2441
rect 3838 2436 3844 2437
rect 3886 2440 3892 2441
rect 3886 2436 3887 2440
rect 3891 2436 3892 2440
rect 3886 2435 3892 2436
rect 4086 2440 4092 2441
rect 4086 2436 4087 2440
rect 4091 2436 4092 2440
rect 4086 2435 4092 2436
rect 4326 2440 4332 2441
rect 4326 2436 4327 2440
rect 4331 2436 4332 2440
rect 4326 2435 4332 2436
rect 4582 2440 4588 2441
rect 4582 2436 4583 2440
rect 4587 2436 4588 2440
rect 4582 2435 4588 2436
rect 4846 2440 4852 2441
rect 4846 2436 4847 2440
rect 4851 2436 4852 2440
rect 4846 2435 4852 2436
rect 5118 2440 5124 2441
rect 5118 2436 5119 2440
rect 5123 2436 5124 2440
rect 5118 2435 5124 2436
rect 5398 2440 5404 2441
rect 5398 2436 5399 2440
rect 5403 2436 5404 2440
rect 5662 2437 5663 2441
rect 5667 2437 5668 2441
rect 5662 2436 5668 2437
rect 5398 2435 5404 2436
rect 1994 2433 2000 2434
rect 1974 2432 1980 2433
rect 1974 2428 1975 2432
rect 1979 2428 1980 2432
rect 1994 2429 1995 2433
rect 1999 2429 2000 2433
rect 1994 2428 2000 2429
rect 2194 2433 2200 2434
rect 2194 2429 2195 2433
rect 2199 2429 2200 2433
rect 2194 2428 2200 2429
rect 2418 2433 2424 2434
rect 2418 2429 2419 2433
rect 2423 2429 2424 2433
rect 2418 2428 2424 2429
rect 2650 2433 2656 2434
rect 2650 2429 2651 2433
rect 2655 2429 2656 2433
rect 2650 2428 2656 2429
rect 2898 2433 2904 2434
rect 2898 2429 2899 2433
rect 2903 2429 2904 2433
rect 2898 2428 2904 2429
rect 3154 2433 3160 2434
rect 3154 2429 3155 2433
rect 3159 2429 3160 2433
rect 3154 2428 3160 2429
rect 3410 2433 3416 2434
rect 3410 2429 3411 2433
rect 3415 2429 3416 2433
rect 3410 2428 3416 2429
rect 3650 2433 3656 2434
rect 3650 2429 3651 2433
rect 3655 2429 3656 2433
rect 3650 2428 3656 2429
rect 3798 2432 3804 2433
rect 3798 2428 3799 2432
rect 3803 2428 3804 2432
rect 1974 2427 1980 2428
rect 111 2422 115 2423
rect 111 2417 115 2418
rect 227 2422 231 2423
rect 227 2417 231 2418
rect 355 2422 359 2423
rect 355 2417 359 2418
rect 523 2422 527 2423
rect 523 2417 527 2418
rect 571 2422 575 2423
rect 571 2417 575 2418
rect 787 2422 791 2423
rect 787 2417 791 2418
rect 835 2422 839 2423
rect 835 2417 839 2418
rect 995 2422 999 2423
rect 995 2417 999 2418
rect 1155 2422 1159 2423
rect 1155 2417 1159 2418
rect 1203 2422 1207 2423
rect 1203 2417 1207 2418
rect 1403 2422 1407 2423
rect 1403 2417 1407 2418
rect 1483 2422 1487 2423
rect 1483 2417 1487 2418
rect 1603 2422 1607 2423
rect 1603 2417 1607 2418
rect 1787 2422 1791 2423
rect 1787 2417 1791 2418
rect 1935 2422 1939 2423
rect 1935 2417 1939 2418
rect 112 2357 114 2417
rect 110 2356 116 2357
rect 228 2356 230 2417
rect 524 2356 526 2417
rect 836 2356 838 2417
rect 1156 2356 1158 2417
rect 1484 2356 1486 2417
rect 1788 2356 1790 2417
rect 1936 2357 1938 2417
rect 1976 2359 1978 2427
rect 1996 2359 1998 2428
rect 2196 2359 2198 2428
rect 2420 2359 2422 2428
rect 2652 2359 2654 2428
rect 2900 2359 2902 2428
rect 3156 2359 3158 2428
rect 3412 2359 3414 2428
rect 3652 2359 3654 2428
rect 3798 2427 3804 2428
rect 3800 2359 3802 2427
rect 3858 2425 3864 2426
rect 3838 2424 3844 2425
rect 3838 2420 3839 2424
rect 3843 2420 3844 2424
rect 3858 2421 3859 2425
rect 3863 2421 3864 2425
rect 3858 2420 3864 2421
rect 4058 2425 4064 2426
rect 4058 2421 4059 2425
rect 4063 2421 4064 2425
rect 4058 2420 4064 2421
rect 4298 2425 4304 2426
rect 4298 2421 4299 2425
rect 4303 2421 4304 2425
rect 4298 2420 4304 2421
rect 4554 2425 4560 2426
rect 4554 2421 4555 2425
rect 4559 2421 4560 2425
rect 4554 2420 4560 2421
rect 4818 2425 4824 2426
rect 4818 2421 4819 2425
rect 4823 2421 4824 2425
rect 4818 2420 4824 2421
rect 5090 2425 5096 2426
rect 5090 2421 5091 2425
rect 5095 2421 5096 2425
rect 5090 2420 5096 2421
rect 5370 2425 5376 2426
rect 5370 2421 5371 2425
rect 5375 2421 5376 2425
rect 5370 2420 5376 2421
rect 5662 2424 5668 2425
rect 5662 2420 5663 2424
rect 5667 2420 5668 2424
rect 3838 2419 3844 2420
rect 1975 2358 1979 2359
rect 1934 2356 1940 2357
rect 110 2352 111 2356
rect 115 2352 116 2356
rect 110 2351 116 2352
rect 226 2355 232 2356
rect 226 2351 227 2355
rect 231 2351 232 2355
rect 226 2350 232 2351
rect 522 2355 528 2356
rect 522 2351 523 2355
rect 527 2351 528 2355
rect 522 2350 528 2351
rect 834 2355 840 2356
rect 834 2351 835 2355
rect 839 2351 840 2355
rect 834 2350 840 2351
rect 1154 2355 1160 2356
rect 1154 2351 1155 2355
rect 1159 2351 1160 2355
rect 1154 2350 1160 2351
rect 1482 2355 1488 2356
rect 1482 2351 1483 2355
rect 1487 2351 1488 2355
rect 1482 2350 1488 2351
rect 1786 2355 1792 2356
rect 1786 2351 1787 2355
rect 1791 2351 1792 2355
rect 1934 2352 1935 2356
rect 1939 2352 1940 2356
rect 1975 2353 1979 2354
rect 1995 2358 1999 2359
rect 1995 2353 1999 2354
rect 2155 2358 2159 2359
rect 2155 2353 2159 2354
rect 2195 2358 2199 2359
rect 2195 2353 2199 2354
rect 2347 2358 2351 2359
rect 2347 2353 2351 2354
rect 2419 2358 2423 2359
rect 2419 2353 2423 2354
rect 2539 2358 2543 2359
rect 2539 2353 2543 2354
rect 2651 2358 2655 2359
rect 2651 2353 2655 2354
rect 2731 2358 2735 2359
rect 2731 2353 2735 2354
rect 2899 2358 2903 2359
rect 2899 2353 2903 2354
rect 2923 2358 2927 2359
rect 2923 2353 2927 2354
rect 3115 2358 3119 2359
rect 3115 2353 3119 2354
rect 3155 2358 3159 2359
rect 3155 2353 3159 2354
rect 3299 2358 3303 2359
rect 3299 2353 3303 2354
rect 3411 2358 3415 2359
rect 3411 2353 3415 2354
rect 3483 2358 3487 2359
rect 3483 2353 3487 2354
rect 3651 2358 3655 2359
rect 3651 2353 3655 2354
rect 3799 2358 3803 2359
rect 3799 2353 3803 2354
rect 1934 2351 1940 2352
rect 1786 2350 1792 2351
rect 254 2340 260 2341
rect 110 2339 116 2340
rect 110 2335 111 2339
rect 115 2335 116 2339
rect 254 2336 255 2340
rect 259 2336 260 2340
rect 254 2335 260 2336
rect 550 2340 556 2341
rect 550 2336 551 2340
rect 555 2336 556 2340
rect 550 2335 556 2336
rect 862 2340 868 2341
rect 862 2336 863 2340
rect 867 2336 868 2340
rect 862 2335 868 2336
rect 1182 2340 1188 2341
rect 1182 2336 1183 2340
rect 1187 2336 1188 2340
rect 1182 2335 1188 2336
rect 1510 2340 1516 2341
rect 1510 2336 1511 2340
rect 1515 2336 1516 2340
rect 1510 2335 1516 2336
rect 1814 2340 1820 2341
rect 1814 2336 1815 2340
rect 1819 2336 1820 2340
rect 1814 2335 1820 2336
rect 1934 2339 1940 2340
rect 1934 2335 1935 2339
rect 1939 2335 1940 2339
rect 110 2334 116 2335
rect 112 2295 114 2334
rect 256 2295 258 2335
rect 552 2295 554 2335
rect 864 2295 866 2335
rect 1184 2295 1186 2335
rect 1512 2295 1514 2335
rect 1816 2295 1818 2335
rect 1934 2334 1940 2335
rect 1936 2295 1938 2334
rect 111 2294 115 2295
rect 111 2289 115 2290
rect 159 2294 163 2295
rect 159 2289 163 2290
rect 255 2294 259 2295
rect 255 2289 259 2290
rect 367 2294 371 2295
rect 367 2289 371 2290
rect 551 2294 555 2295
rect 551 2289 555 2290
rect 599 2294 603 2295
rect 599 2289 603 2290
rect 831 2294 835 2295
rect 831 2289 835 2290
rect 863 2294 867 2295
rect 863 2289 867 2290
rect 1063 2294 1067 2295
rect 1063 2289 1067 2290
rect 1183 2294 1187 2295
rect 1183 2289 1187 2290
rect 1511 2294 1515 2295
rect 1511 2289 1515 2290
rect 1815 2294 1819 2295
rect 1815 2289 1819 2290
rect 1935 2294 1939 2295
rect 1976 2293 1978 2353
rect 1935 2289 1939 2290
rect 1974 2292 1980 2293
rect 1996 2292 1998 2353
rect 2156 2292 2158 2353
rect 2348 2292 2350 2353
rect 2540 2292 2542 2353
rect 2732 2292 2734 2353
rect 2924 2292 2926 2353
rect 3116 2292 3118 2353
rect 3300 2292 3302 2353
rect 3484 2292 3486 2353
rect 3652 2292 3654 2353
rect 3800 2293 3802 2353
rect 3840 2347 3842 2419
rect 3860 2347 3862 2420
rect 4060 2347 4062 2420
rect 4300 2347 4302 2420
rect 4556 2347 4558 2420
rect 4820 2347 4822 2420
rect 5092 2347 5094 2420
rect 5372 2347 5374 2420
rect 5662 2419 5668 2420
rect 5664 2347 5666 2419
rect 3839 2346 3843 2347
rect 3839 2341 3843 2342
rect 3859 2346 3863 2347
rect 3859 2341 3863 2342
rect 4059 2346 4063 2347
rect 4059 2341 4063 2342
rect 4299 2346 4303 2347
rect 4299 2341 4303 2342
rect 4443 2346 4447 2347
rect 4443 2341 4447 2342
rect 4555 2346 4559 2347
rect 4555 2341 4559 2342
rect 4611 2346 4615 2347
rect 4611 2341 4615 2342
rect 4787 2346 4791 2347
rect 4787 2341 4791 2342
rect 4819 2346 4823 2347
rect 4819 2341 4823 2342
rect 4963 2346 4967 2347
rect 4963 2341 4967 2342
rect 5091 2346 5095 2347
rect 5091 2341 5095 2342
rect 5147 2346 5151 2347
rect 5147 2341 5151 2342
rect 5339 2346 5343 2347
rect 5339 2341 5343 2342
rect 5371 2346 5375 2347
rect 5371 2341 5375 2342
rect 5515 2346 5519 2347
rect 5515 2341 5519 2342
rect 5663 2346 5667 2347
rect 5663 2341 5667 2342
rect 3798 2292 3804 2293
rect 112 2266 114 2289
rect 110 2265 116 2266
rect 160 2265 162 2289
rect 368 2265 370 2289
rect 600 2265 602 2289
rect 832 2265 834 2289
rect 1064 2265 1066 2289
rect 1936 2266 1938 2289
rect 1974 2288 1975 2292
rect 1979 2288 1980 2292
rect 1974 2287 1980 2288
rect 1994 2291 2000 2292
rect 1994 2287 1995 2291
rect 1999 2287 2000 2291
rect 1994 2286 2000 2287
rect 2154 2291 2160 2292
rect 2154 2287 2155 2291
rect 2159 2287 2160 2291
rect 2154 2286 2160 2287
rect 2346 2291 2352 2292
rect 2346 2287 2347 2291
rect 2351 2287 2352 2291
rect 2346 2286 2352 2287
rect 2538 2291 2544 2292
rect 2538 2287 2539 2291
rect 2543 2287 2544 2291
rect 2538 2286 2544 2287
rect 2730 2291 2736 2292
rect 2730 2287 2731 2291
rect 2735 2287 2736 2291
rect 2730 2286 2736 2287
rect 2922 2291 2928 2292
rect 2922 2287 2923 2291
rect 2927 2287 2928 2291
rect 2922 2286 2928 2287
rect 3114 2291 3120 2292
rect 3114 2287 3115 2291
rect 3119 2287 3120 2291
rect 3114 2286 3120 2287
rect 3298 2291 3304 2292
rect 3298 2287 3299 2291
rect 3303 2287 3304 2291
rect 3298 2286 3304 2287
rect 3482 2291 3488 2292
rect 3482 2287 3483 2291
rect 3487 2287 3488 2291
rect 3482 2286 3488 2287
rect 3650 2291 3656 2292
rect 3650 2287 3651 2291
rect 3655 2287 3656 2291
rect 3798 2288 3799 2292
rect 3803 2288 3804 2292
rect 3798 2287 3804 2288
rect 3650 2286 3656 2287
rect 3840 2281 3842 2341
rect 3838 2280 3844 2281
rect 4444 2280 4446 2341
rect 4612 2280 4614 2341
rect 4788 2280 4790 2341
rect 4964 2280 4966 2341
rect 5148 2280 5150 2341
rect 5340 2280 5342 2341
rect 5516 2280 5518 2341
rect 5664 2281 5666 2341
rect 5662 2280 5668 2281
rect 2022 2276 2028 2277
rect 1974 2275 1980 2276
rect 1974 2271 1975 2275
rect 1979 2271 1980 2275
rect 2022 2272 2023 2276
rect 2027 2272 2028 2276
rect 2022 2271 2028 2272
rect 2182 2276 2188 2277
rect 2182 2272 2183 2276
rect 2187 2272 2188 2276
rect 2182 2271 2188 2272
rect 2374 2276 2380 2277
rect 2374 2272 2375 2276
rect 2379 2272 2380 2276
rect 2374 2271 2380 2272
rect 2566 2276 2572 2277
rect 2566 2272 2567 2276
rect 2571 2272 2572 2276
rect 2566 2271 2572 2272
rect 2758 2276 2764 2277
rect 2758 2272 2759 2276
rect 2763 2272 2764 2276
rect 2758 2271 2764 2272
rect 2950 2276 2956 2277
rect 2950 2272 2951 2276
rect 2955 2272 2956 2276
rect 2950 2271 2956 2272
rect 3142 2276 3148 2277
rect 3142 2272 3143 2276
rect 3147 2272 3148 2276
rect 3142 2271 3148 2272
rect 3326 2276 3332 2277
rect 3326 2272 3327 2276
rect 3331 2272 3332 2276
rect 3326 2271 3332 2272
rect 3510 2276 3516 2277
rect 3510 2272 3511 2276
rect 3515 2272 3516 2276
rect 3510 2271 3516 2272
rect 3678 2276 3684 2277
rect 3838 2276 3839 2280
rect 3843 2276 3844 2280
rect 3678 2272 3679 2276
rect 3683 2272 3684 2276
rect 3678 2271 3684 2272
rect 3798 2275 3804 2276
rect 3838 2275 3844 2276
rect 4442 2279 4448 2280
rect 4442 2275 4443 2279
rect 4447 2275 4448 2279
rect 3798 2271 3799 2275
rect 3803 2271 3804 2275
rect 4442 2274 4448 2275
rect 4610 2279 4616 2280
rect 4610 2275 4611 2279
rect 4615 2275 4616 2279
rect 4610 2274 4616 2275
rect 4786 2279 4792 2280
rect 4786 2275 4787 2279
rect 4791 2275 4792 2279
rect 4786 2274 4792 2275
rect 4962 2279 4968 2280
rect 4962 2275 4963 2279
rect 4967 2275 4968 2279
rect 4962 2274 4968 2275
rect 5146 2279 5152 2280
rect 5146 2275 5147 2279
rect 5151 2275 5152 2279
rect 5146 2274 5152 2275
rect 5338 2279 5344 2280
rect 5338 2275 5339 2279
rect 5343 2275 5344 2279
rect 5338 2274 5344 2275
rect 5514 2279 5520 2280
rect 5514 2275 5515 2279
rect 5519 2275 5520 2279
rect 5662 2276 5663 2280
rect 5667 2276 5668 2280
rect 5662 2275 5668 2276
rect 5514 2274 5520 2275
rect 1974 2270 1980 2271
rect 1934 2265 1940 2266
rect 110 2261 111 2265
rect 115 2261 116 2265
rect 110 2260 116 2261
rect 158 2264 164 2265
rect 158 2260 159 2264
rect 163 2260 164 2264
rect 158 2259 164 2260
rect 366 2264 372 2265
rect 366 2260 367 2264
rect 371 2260 372 2264
rect 366 2259 372 2260
rect 598 2264 604 2265
rect 598 2260 599 2264
rect 603 2260 604 2264
rect 598 2259 604 2260
rect 830 2264 836 2265
rect 830 2260 831 2264
rect 835 2260 836 2264
rect 830 2259 836 2260
rect 1062 2264 1068 2265
rect 1062 2260 1063 2264
rect 1067 2260 1068 2264
rect 1934 2261 1935 2265
rect 1939 2261 1940 2265
rect 1934 2260 1940 2261
rect 1062 2259 1068 2260
rect 130 2249 136 2250
rect 110 2248 116 2249
rect 110 2244 111 2248
rect 115 2244 116 2248
rect 130 2245 131 2249
rect 135 2245 136 2249
rect 130 2244 136 2245
rect 338 2249 344 2250
rect 338 2245 339 2249
rect 343 2245 344 2249
rect 338 2244 344 2245
rect 570 2249 576 2250
rect 570 2245 571 2249
rect 575 2245 576 2249
rect 570 2244 576 2245
rect 802 2249 808 2250
rect 802 2245 803 2249
rect 807 2245 808 2249
rect 802 2244 808 2245
rect 1034 2249 1040 2250
rect 1034 2245 1035 2249
rect 1039 2245 1040 2249
rect 1034 2244 1040 2245
rect 1934 2248 1940 2249
rect 1934 2244 1935 2248
rect 1939 2244 1940 2248
rect 110 2243 116 2244
rect 112 2171 114 2243
rect 132 2171 134 2244
rect 340 2171 342 2244
rect 572 2171 574 2244
rect 804 2171 806 2244
rect 1036 2171 1038 2244
rect 1934 2243 1940 2244
rect 1936 2171 1938 2243
rect 1976 2239 1978 2270
rect 2024 2239 2026 2271
rect 2184 2239 2186 2271
rect 2376 2239 2378 2271
rect 2568 2239 2570 2271
rect 2760 2239 2762 2271
rect 2952 2239 2954 2271
rect 3144 2239 3146 2271
rect 3328 2239 3330 2271
rect 3512 2239 3514 2271
rect 3680 2239 3682 2271
rect 3798 2270 3804 2271
rect 3800 2239 3802 2270
rect 4470 2264 4476 2265
rect 3838 2263 3844 2264
rect 3838 2259 3839 2263
rect 3843 2259 3844 2263
rect 4470 2260 4471 2264
rect 4475 2260 4476 2264
rect 4470 2259 4476 2260
rect 4638 2264 4644 2265
rect 4638 2260 4639 2264
rect 4643 2260 4644 2264
rect 4638 2259 4644 2260
rect 4814 2264 4820 2265
rect 4814 2260 4815 2264
rect 4819 2260 4820 2264
rect 4814 2259 4820 2260
rect 4990 2264 4996 2265
rect 4990 2260 4991 2264
rect 4995 2260 4996 2264
rect 4990 2259 4996 2260
rect 5174 2264 5180 2265
rect 5174 2260 5175 2264
rect 5179 2260 5180 2264
rect 5174 2259 5180 2260
rect 5366 2264 5372 2265
rect 5366 2260 5367 2264
rect 5371 2260 5372 2264
rect 5366 2259 5372 2260
rect 5542 2264 5548 2265
rect 5542 2260 5543 2264
rect 5547 2260 5548 2264
rect 5542 2259 5548 2260
rect 5662 2263 5668 2264
rect 5662 2259 5663 2263
rect 5667 2259 5668 2263
rect 3838 2258 3844 2259
rect 1975 2238 1979 2239
rect 1975 2233 1979 2234
rect 2023 2238 2027 2239
rect 2023 2233 2027 2234
rect 2183 2238 2187 2239
rect 2183 2233 2187 2234
rect 2191 2238 2195 2239
rect 2191 2233 2195 2234
rect 2359 2238 2363 2239
rect 2359 2233 2363 2234
rect 2375 2238 2379 2239
rect 2375 2233 2379 2234
rect 2535 2238 2539 2239
rect 2535 2233 2539 2234
rect 2567 2238 2571 2239
rect 2567 2233 2571 2234
rect 2711 2238 2715 2239
rect 2711 2233 2715 2234
rect 2759 2238 2763 2239
rect 2759 2233 2763 2234
rect 2879 2238 2883 2239
rect 2879 2233 2883 2234
rect 2951 2238 2955 2239
rect 2951 2233 2955 2234
rect 3047 2238 3051 2239
rect 3047 2233 3051 2234
rect 3143 2238 3147 2239
rect 3143 2233 3147 2234
rect 3207 2238 3211 2239
rect 3207 2233 3211 2234
rect 3327 2238 3331 2239
rect 3327 2233 3331 2234
rect 3367 2238 3371 2239
rect 3367 2233 3371 2234
rect 3511 2238 3515 2239
rect 3511 2233 3515 2234
rect 3535 2238 3539 2239
rect 3535 2233 3539 2234
rect 3679 2238 3683 2239
rect 3679 2233 3683 2234
rect 3799 2238 3803 2239
rect 3799 2233 3803 2234
rect 1976 2210 1978 2233
rect 1974 2209 1980 2210
rect 2024 2209 2026 2233
rect 2192 2209 2194 2233
rect 2360 2209 2362 2233
rect 2536 2209 2538 2233
rect 2712 2209 2714 2233
rect 2880 2209 2882 2233
rect 3048 2209 3050 2233
rect 3208 2209 3210 2233
rect 3368 2209 3370 2233
rect 3536 2209 3538 2233
rect 3680 2209 3682 2233
rect 3800 2210 3802 2233
rect 3840 2223 3842 2258
rect 4472 2223 4474 2259
rect 4640 2223 4642 2259
rect 4816 2223 4818 2259
rect 4992 2223 4994 2259
rect 5176 2223 5178 2259
rect 5368 2223 5370 2259
rect 5544 2223 5546 2259
rect 5662 2258 5668 2259
rect 5664 2223 5666 2258
rect 3839 2222 3843 2223
rect 3839 2217 3843 2218
rect 4471 2222 4475 2223
rect 4471 2217 4475 2218
rect 4543 2222 4547 2223
rect 4543 2217 4547 2218
rect 4639 2222 4643 2223
rect 4639 2217 4643 2218
rect 4719 2222 4723 2223
rect 4719 2217 4723 2218
rect 4815 2222 4819 2223
rect 4815 2217 4819 2218
rect 4911 2222 4915 2223
rect 4911 2217 4915 2218
rect 4991 2222 4995 2223
rect 4991 2217 4995 2218
rect 5119 2222 5123 2223
rect 5119 2217 5123 2218
rect 5175 2222 5179 2223
rect 5175 2217 5179 2218
rect 5335 2222 5339 2223
rect 5335 2217 5339 2218
rect 5367 2222 5371 2223
rect 5367 2217 5371 2218
rect 5543 2222 5547 2223
rect 5543 2217 5547 2218
rect 5663 2222 5667 2223
rect 5663 2217 5667 2218
rect 3798 2209 3804 2210
rect 1974 2205 1975 2209
rect 1979 2205 1980 2209
rect 1974 2204 1980 2205
rect 2022 2208 2028 2209
rect 2022 2204 2023 2208
rect 2027 2204 2028 2208
rect 2022 2203 2028 2204
rect 2190 2208 2196 2209
rect 2190 2204 2191 2208
rect 2195 2204 2196 2208
rect 2190 2203 2196 2204
rect 2358 2208 2364 2209
rect 2358 2204 2359 2208
rect 2363 2204 2364 2208
rect 2358 2203 2364 2204
rect 2534 2208 2540 2209
rect 2534 2204 2535 2208
rect 2539 2204 2540 2208
rect 2534 2203 2540 2204
rect 2710 2208 2716 2209
rect 2710 2204 2711 2208
rect 2715 2204 2716 2208
rect 2710 2203 2716 2204
rect 2878 2208 2884 2209
rect 2878 2204 2879 2208
rect 2883 2204 2884 2208
rect 2878 2203 2884 2204
rect 3046 2208 3052 2209
rect 3046 2204 3047 2208
rect 3051 2204 3052 2208
rect 3046 2203 3052 2204
rect 3206 2208 3212 2209
rect 3206 2204 3207 2208
rect 3211 2204 3212 2208
rect 3206 2203 3212 2204
rect 3366 2208 3372 2209
rect 3366 2204 3367 2208
rect 3371 2204 3372 2208
rect 3366 2203 3372 2204
rect 3534 2208 3540 2209
rect 3534 2204 3535 2208
rect 3539 2204 3540 2208
rect 3534 2203 3540 2204
rect 3678 2208 3684 2209
rect 3678 2204 3679 2208
rect 3683 2204 3684 2208
rect 3798 2205 3799 2209
rect 3803 2205 3804 2209
rect 3798 2204 3804 2205
rect 3678 2203 3684 2204
rect 3840 2194 3842 2217
rect 1994 2193 2000 2194
rect 1974 2192 1980 2193
rect 1974 2188 1975 2192
rect 1979 2188 1980 2192
rect 1994 2189 1995 2193
rect 1999 2189 2000 2193
rect 1994 2188 2000 2189
rect 2162 2193 2168 2194
rect 2162 2189 2163 2193
rect 2167 2189 2168 2193
rect 2162 2188 2168 2189
rect 2330 2193 2336 2194
rect 2330 2189 2331 2193
rect 2335 2189 2336 2193
rect 2330 2188 2336 2189
rect 2506 2193 2512 2194
rect 2506 2189 2507 2193
rect 2511 2189 2512 2193
rect 2506 2188 2512 2189
rect 2682 2193 2688 2194
rect 2682 2189 2683 2193
rect 2687 2189 2688 2193
rect 2682 2188 2688 2189
rect 2850 2193 2856 2194
rect 2850 2189 2851 2193
rect 2855 2189 2856 2193
rect 2850 2188 2856 2189
rect 3018 2193 3024 2194
rect 3018 2189 3019 2193
rect 3023 2189 3024 2193
rect 3018 2188 3024 2189
rect 3178 2193 3184 2194
rect 3178 2189 3179 2193
rect 3183 2189 3184 2193
rect 3178 2188 3184 2189
rect 3338 2193 3344 2194
rect 3338 2189 3339 2193
rect 3343 2189 3344 2193
rect 3338 2188 3344 2189
rect 3506 2193 3512 2194
rect 3506 2189 3507 2193
rect 3511 2189 3512 2193
rect 3506 2188 3512 2189
rect 3650 2193 3656 2194
rect 3838 2193 3844 2194
rect 4544 2193 4546 2217
rect 4720 2193 4722 2217
rect 4912 2193 4914 2217
rect 5120 2193 5122 2217
rect 5336 2193 5338 2217
rect 5544 2193 5546 2217
rect 5664 2194 5666 2217
rect 5662 2193 5668 2194
rect 3650 2189 3651 2193
rect 3655 2189 3656 2193
rect 3650 2188 3656 2189
rect 3798 2192 3804 2193
rect 3798 2188 3799 2192
rect 3803 2188 3804 2192
rect 3838 2189 3839 2193
rect 3843 2189 3844 2193
rect 3838 2188 3844 2189
rect 4542 2192 4548 2193
rect 4542 2188 4543 2192
rect 4547 2188 4548 2192
rect 1974 2187 1980 2188
rect 111 2170 115 2171
rect 111 2165 115 2166
rect 131 2170 135 2171
rect 131 2165 135 2166
rect 339 2170 343 2171
rect 339 2165 343 2166
rect 347 2170 351 2171
rect 347 2165 351 2166
rect 571 2170 575 2171
rect 571 2165 575 2166
rect 595 2170 599 2171
rect 595 2165 599 2166
rect 803 2170 807 2171
rect 803 2165 807 2166
rect 835 2170 839 2171
rect 835 2165 839 2166
rect 1035 2170 1039 2171
rect 1035 2165 1039 2166
rect 1075 2170 1079 2171
rect 1075 2165 1079 2166
rect 1315 2170 1319 2171
rect 1315 2165 1319 2166
rect 1563 2170 1567 2171
rect 1563 2165 1567 2166
rect 1787 2170 1791 2171
rect 1787 2165 1791 2166
rect 1935 2170 1939 2171
rect 1935 2165 1939 2166
rect 112 2105 114 2165
rect 110 2104 116 2105
rect 132 2104 134 2165
rect 348 2104 350 2165
rect 596 2104 598 2165
rect 836 2104 838 2165
rect 1076 2104 1078 2165
rect 1316 2104 1318 2165
rect 1564 2104 1566 2165
rect 1788 2104 1790 2165
rect 1936 2105 1938 2165
rect 1976 2111 1978 2187
rect 1996 2111 1998 2188
rect 2164 2111 2166 2188
rect 2332 2111 2334 2188
rect 2508 2111 2510 2188
rect 2684 2111 2686 2188
rect 2852 2111 2854 2188
rect 3020 2111 3022 2188
rect 3180 2111 3182 2188
rect 3340 2111 3342 2188
rect 3508 2111 3510 2188
rect 3652 2111 3654 2188
rect 3798 2187 3804 2188
rect 4542 2187 4548 2188
rect 4718 2192 4724 2193
rect 4718 2188 4719 2192
rect 4723 2188 4724 2192
rect 4718 2187 4724 2188
rect 4910 2192 4916 2193
rect 4910 2188 4911 2192
rect 4915 2188 4916 2192
rect 4910 2187 4916 2188
rect 5118 2192 5124 2193
rect 5118 2188 5119 2192
rect 5123 2188 5124 2192
rect 5118 2187 5124 2188
rect 5334 2192 5340 2193
rect 5334 2188 5335 2192
rect 5339 2188 5340 2192
rect 5334 2187 5340 2188
rect 5542 2192 5548 2193
rect 5542 2188 5543 2192
rect 5547 2188 5548 2192
rect 5662 2189 5663 2193
rect 5667 2189 5668 2193
rect 5662 2188 5668 2189
rect 5542 2187 5548 2188
rect 3800 2111 3802 2187
rect 4514 2177 4520 2178
rect 3838 2176 3844 2177
rect 3838 2172 3839 2176
rect 3843 2172 3844 2176
rect 4514 2173 4515 2177
rect 4519 2173 4520 2177
rect 4514 2172 4520 2173
rect 4690 2177 4696 2178
rect 4690 2173 4691 2177
rect 4695 2173 4696 2177
rect 4690 2172 4696 2173
rect 4882 2177 4888 2178
rect 4882 2173 4883 2177
rect 4887 2173 4888 2177
rect 4882 2172 4888 2173
rect 5090 2177 5096 2178
rect 5090 2173 5091 2177
rect 5095 2173 5096 2177
rect 5090 2172 5096 2173
rect 5306 2177 5312 2178
rect 5306 2173 5307 2177
rect 5311 2173 5312 2177
rect 5306 2172 5312 2173
rect 5514 2177 5520 2178
rect 5514 2173 5515 2177
rect 5519 2173 5520 2177
rect 5514 2172 5520 2173
rect 5662 2176 5668 2177
rect 5662 2172 5663 2176
rect 5667 2172 5668 2176
rect 3838 2171 3844 2172
rect 3840 2111 3842 2171
rect 4516 2111 4518 2172
rect 4692 2111 4694 2172
rect 4884 2111 4886 2172
rect 5092 2111 5094 2172
rect 5308 2111 5310 2172
rect 5516 2111 5518 2172
rect 5662 2171 5668 2172
rect 5664 2111 5666 2171
rect 1975 2110 1979 2111
rect 1975 2105 1979 2106
rect 1995 2110 1999 2111
rect 1995 2105 1999 2106
rect 2163 2110 2167 2111
rect 2163 2105 2167 2106
rect 2331 2110 2335 2111
rect 2331 2105 2335 2106
rect 2507 2110 2511 2111
rect 2507 2105 2511 2106
rect 2683 2110 2687 2111
rect 2683 2105 2687 2106
rect 2851 2110 2855 2111
rect 2851 2105 2855 2106
rect 3019 2110 3023 2111
rect 3019 2105 3023 2106
rect 3107 2110 3111 2111
rect 3107 2105 3111 2106
rect 3179 2110 3183 2111
rect 3179 2105 3183 2106
rect 3243 2110 3247 2111
rect 3243 2105 3247 2106
rect 3339 2110 3343 2111
rect 3339 2105 3343 2106
rect 3379 2110 3383 2111
rect 3379 2105 3383 2106
rect 3507 2110 3511 2111
rect 3507 2105 3511 2106
rect 3515 2110 3519 2111
rect 3515 2105 3519 2106
rect 3651 2110 3655 2111
rect 3651 2105 3655 2106
rect 3799 2110 3803 2111
rect 3799 2105 3803 2106
rect 3839 2110 3843 2111
rect 3839 2105 3843 2106
rect 4515 2110 4519 2111
rect 4515 2105 4519 2106
rect 4635 2110 4639 2111
rect 4635 2105 4639 2106
rect 4691 2110 4695 2111
rect 4691 2105 4695 2106
rect 4771 2110 4775 2111
rect 4771 2105 4775 2106
rect 4883 2110 4887 2111
rect 4883 2105 4887 2106
rect 4907 2110 4911 2111
rect 4907 2105 4911 2106
rect 5043 2110 5047 2111
rect 5043 2105 5047 2106
rect 5091 2110 5095 2111
rect 5091 2105 5095 2106
rect 5179 2110 5183 2111
rect 5179 2105 5183 2106
rect 5307 2110 5311 2111
rect 5307 2105 5311 2106
rect 5515 2110 5519 2111
rect 5515 2105 5519 2106
rect 5663 2110 5667 2111
rect 5663 2105 5667 2106
rect 1934 2104 1940 2105
rect 110 2100 111 2104
rect 115 2100 116 2104
rect 110 2099 116 2100
rect 130 2103 136 2104
rect 130 2099 131 2103
rect 135 2099 136 2103
rect 130 2098 136 2099
rect 346 2103 352 2104
rect 346 2099 347 2103
rect 351 2099 352 2103
rect 346 2098 352 2099
rect 594 2103 600 2104
rect 594 2099 595 2103
rect 599 2099 600 2103
rect 594 2098 600 2099
rect 834 2103 840 2104
rect 834 2099 835 2103
rect 839 2099 840 2103
rect 834 2098 840 2099
rect 1074 2103 1080 2104
rect 1074 2099 1075 2103
rect 1079 2099 1080 2103
rect 1074 2098 1080 2099
rect 1314 2103 1320 2104
rect 1314 2099 1315 2103
rect 1319 2099 1320 2103
rect 1314 2098 1320 2099
rect 1562 2103 1568 2104
rect 1562 2099 1563 2103
rect 1567 2099 1568 2103
rect 1562 2098 1568 2099
rect 1786 2103 1792 2104
rect 1786 2099 1787 2103
rect 1791 2099 1792 2103
rect 1934 2100 1935 2104
rect 1939 2100 1940 2104
rect 1934 2099 1940 2100
rect 1786 2098 1792 2099
rect 158 2088 164 2089
rect 110 2087 116 2088
rect 110 2083 111 2087
rect 115 2083 116 2087
rect 158 2084 159 2088
rect 163 2084 164 2088
rect 158 2083 164 2084
rect 374 2088 380 2089
rect 374 2084 375 2088
rect 379 2084 380 2088
rect 374 2083 380 2084
rect 622 2088 628 2089
rect 622 2084 623 2088
rect 627 2084 628 2088
rect 622 2083 628 2084
rect 862 2088 868 2089
rect 862 2084 863 2088
rect 867 2084 868 2088
rect 862 2083 868 2084
rect 1102 2088 1108 2089
rect 1102 2084 1103 2088
rect 1107 2084 1108 2088
rect 1102 2083 1108 2084
rect 1342 2088 1348 2089
rect 1342 2084 1343 2088
rect 1347 2084 1348 2088
rect 1342 2083 1348 2084
rect 1590 2088 1596 2089
rect 1590 2084 1591 2088
rect 1595 2084 1596 2088
rect 1590 2083 1596 2084
rect 1814 2088 1820 2089
rect 1814 2084 1815 2088
rect 1819 2084 1820 2088
rect 1814 2083 1820 2084
rect 1934 2087 1940 2088
rect 1934 2083 1935 2087
rect 1939 2083 1940 2087
rect 110 2082 116 2083
rect 112 2055 114 2082
rect 160 2055 162 2083
rect 376 2055 378 2083
rect 624 2055 626 2083
rect 864 2055 866 2083
rect 1104 2055 1106 2083
rect 1344 2055 1346 2083
rect 1592 2055 1594 2083
rect 1816 2055 1818 2083
rect 1934 2082 1940 2083
rect 1936 2055 1938 2082
rect 111 2054 115 2055
rect 111 2049 115 2050
rect 159 2054 163 2055
rect 159 2049 163 2050
rect 271 2054 275 2055
rect 271 2049 275 2050
rect 375 2054 379 2055
rect 375 2049 379 2050
rect 407 2054 411 2055
rect 407 2049 411 2050
rect 543 2054 547 2055
rect 543 2049 547 2050
rect 623 2054 627 2055
rect 623 2049 627 2050
rect 687 2054 691 2055
rect 687 2049 691 2050
rect 831 2054 835 2055
rect 831 2049 835 2050
rect 863 2054 867 2055
rect 863 2049 867 2050
rect 975 2054 979 2055
rect 975 2049 979 2050
rect 1103 2054 1107 2055
rect 1103 2049 1107 2050
rect 1119 2054 1123 2055
rect 1119 2049 1123 2050
rect 1263 2054 1267 2055
rect 1263 2049 1267 2050
rect 1343 2054 1347 2055
rect 1343 2049 1347 2050
rect 1407 2054 1411 2055
rect 1407 2049 1411 2050
rect 1543 2054 1547 2055
rect 1543 2049 1547 2050
rect 1591 2054 1595 2055
rect 1591 2049 1595 2050
rect 1679 2054 1683 2055
rect 1679 2049 1683 2050
rect 1815 2054 1819 2055
rect 1815 2049 1819 2050
rect 1935 2054 1939 2055
rect 1935 2049 1939 2050
rect 112 2026 114 2049
rect 110 2025 116 2026
rect 272 2025 274 2049
rect 408 2025 410 2049
rect 544 2025 546 2049
rect 688 2025 690 2049
rect 832 2025 834 2049
rect 976 2025 978 2049
rect 1120 2025 1122 2049
rect 1264 2025 1266 2049
rect 1408 2025 1410 2049
rect 1544 2025 1546 2049
rect 1680 2025 1682 2049
rect 1816 2025 1818 2049
rect 1936 2026 1938 2049
rect 1976 2045 1978 2105
rect 1974 2044 1980 2045
rect 3108 2044 3110 2105
rect 3244 2044 3246 2105
rect 3380 2044 3382 2105
rect 3516 2044 3518 2105
rect 3652 2044 3654 2105
rect 3800 2045 3802 2105
rect 3840 2045 3842 2105
rect 3798 2044 3804 2045
rect 1974 2040 1975 2044
rect 1979 2040 1980 2044
rect 1974 2039 1980 2040
rect 3106 2043 3112 2044
rect 3106 2039 3107 2043
rect 3111 2039 3112 2043
rect 3106 2038 3112 2039
rect 3242 2043 3248 2044
rect 3242 2039 3243 2043
rect 3247 2039 3248 2043
rect 3242 2038 3248 2039
rect 3378 2043 3384 2044
rect 3378 2039 3379 2043
rect 3383 2039 3384 2043
rect 3378 2038 3384 2039
rect 3514 2043 3520 2044
rect 3514 2039 3515 2043
rect 3519 2039 3520 2043
rect 3514 2038 3520 2039
rect 3650 2043 3656 2044
rect 3650 2039 3651 2043
rect 3655 2039 3656 2043
rect 3798 2040 3799 2044
rect 3803 2040 3804 2044
rect 3798 2039 3804 2040
rect 3838 2044 3844 2045
rect 4636 2044 4638 2105
rect 4772 2044 4774 2105
rect 4908 2044 4910 2105
rect 5044 2044 5046 2105
rect 5180 2044 5182 2105
rect 5664 2045 5666 2105
rect 5662 2044 5668 2045
rect 3838 2040 3839 2044
rect 3843 2040 3844 2044
rect 3838 2039 3844 2040
rect 4634 2043 4640 2044
rect 4634 2039 4635 2043
rect 4639 2039 4640 2043
rect 3650 2038 3656 2039
rect 4634 2038 4640 2039
rect 4770 2043 4776 2044
rect 4770 2039 4771 2043
rect 4775 2039 4776 2043
rect 4770 2038 4776 2039
rect 4906 2043 4912 2044
rect 4906 2039 4907 2043
rect 4911 2039 4912 2043
rect 4906 2038 4912 2039
rect 5042 2043 5048 2044
rect 5042 2039 5043 2043
rect 5047 2039 5048 2043
rect 5042 2038 5048 2039
rect 5178 2043 5184 2044
rect 5178 2039 5179 2043
rect 5183 2039 5184 2043
rect 5662 2040 5663 2044
rect 5667 2040 5668 2044
rect 5662 2039 5668 2040
rect 5178 2038 5184 2039
rect 3134 2028 3140 2029
rect 1974 2027 1980 2028
rect 1934 2025 1940 2026
rect 110 2021 111 2025
rect 115 2021 116 2025
rect 110 2020 116 2021
rect 270 2024 276 2025
rect 270 2020 271 2024
rect 275 2020 276 2024
rect 270 2019 276 2020
rect 406 2024 412 2025
rect 406 2020 407 2024
rect 411 2020 412 2024
rect 406 2019 412 2020
rect 542 2024 548 2025
rect 542 2020 543 2024
rect 547 2020 548 2024
rect 542 2019 548 2020
rect 686 2024 692 2025
rect 686 2020 687 2024
rect 691 2020 692 2024
rect 686 2019 692 2020
rect 830 2024 836 2025
rect 830 2020 831 2024
rect 835 2020 836 2024
rect 830 2019 836 2020
rect 974 2024 980 2025
rect 974 2020 975 2024
rect 979 2020 980 2024
rect 974 2019 980 2020
rect 1118 2024 1124 2025
rect 1118 2020 1119 2024
rect 1123 2020 1124 2024
rect 1118 2019 1124 2020
rect 1262 2024 1268 2025
rect 1262 2020 1263 2024
rect 1267 2020 1268 2024
rect 1262 2019 1268 2020
rect 1406 2024 1412 2025
rect 1406 2020 1407 2024
rect 1411 2020 1412 2024
rect 1406 2019 1412 2020
rect 1542 2024 1548 2025
rect 1542 2020 1543 2024
rect 1547 2020 1548 2024
rect 1542 2019 1548 2020
rect 1678 2024 1684 2025
rect 1678 2020 1679 2024
rect 1683 2020 1684 2024
rect 1678 2019 1684 2020
rect 1814 2024 1820 2025
rect 1814 2020 1815 2024
rect 1819 2020 1820 2024
rect 1934 2021 1935 2025
rect 1939 2021 1940 2025
rect 1974 2023 1975 2027
rect 1979 2023 1980 2027
rect 3134 2024 3135 2028
rect 3139 2024 3140 2028
rect 3134 2023 3140 2024
rect 3270 2028 3276 2029
rect 3270 2024 3271 2028
rect 3275 2024 3276 2028
rect 3270 2023 3276 2024
rect 3406 2028 3412 2029
rect 3406 2024 3407 2028
rect 3411 2024 3412 2028
rect 3406 2023 3412 2024
rect 3542 2028 3548 2029
rect 3542 2024 3543 2028
rect 3547 2024 3548 2028
rect 3542 2023 3548 2024
rect 3678 2028 3684 2029
rect 4662 2028 4668 2029
rect 3678 2024 3679 2028
rect 3683 2024 3684 2028
rect 3678 2023 3684 2024
rect 3798 2027 3804 2028
rect 3798 2023 3799 2027
rect 3803 2023 3804 2027
rect 1974 2022 1980 2023
rect 1934 2020 1940 2021
rect 1814 2019 1820 2020
rect 242 2009 248 2010
rect 110 2008 116 2009
rect 110 2004 111 2008
rect 115 2004 116 2008
rect 242 2005 243 2009
rect 247 2005 248 2009
rect 242 2004 248 2005
rect 378 2009 384 2010
rect 378 2005 379 2009
rect 383 2005 384 2009
rect 378 2004 384 2005
rect 514 2009 520 2010
rect 514 2005 515 2009
rect 519 2005 520 2009
rect 514 2004 520 2005
rect 658 2009 664 2010
rect 658 2005 659 2009
rect 663 2005 664 2009
rect 658 2004 664 2005
rect 802 2009 808 2010
rect 802 2005 803 2009
rect 807 2005 808 2009
rect 802 2004 808 2005
rect 946 2009 952 2010
rect 946 2005 947 2009
rect 951 2005 952 2009
rect 946 2004 952 2005
rect 1090 2009 1096 2010
rect 1090 2005 1091 2009
rect 1095 2005 1096 2009
rect 1090 2004 1096 2005
rect 1234 2009 1240 2010
rect 1234 2005 1235 2009
rect 1239 2005 1240 2009
rect 1234 2004 1240 2005
rect 1378 2009 1384 2010
rect 1378 2005 1379 2009
rect 1383 2005 1384 2009
rect 1378 2004 1384 2005
rect 1514 2009 1520 2010
rect 1514 2005 1515 2009
rect 1519 2005 1520 2009
rect 1514 2004 1520 2005
rect 1650 2009 1656 2010
rect 1650 2005 1651 2009
rect 1655 2005 1656 2009
rect 1650 2004 1656 2005
rect 1786 2009 1792 2010
rect 1786 2005 1787 2009
rect 1791 2005 1792 2009
rect 1786 2004 1792 2005
rect 1934 2008 1940 2009
rect 1934 2004 1935 2008
rect 1939 2004 1940 2008
rect 110 2003 116 2004
rect 112 1939 114 2003
rect 244 1939 246 2004
rect 380 1939 382 2004
rect 516 1939 518 2004
rect 660 1939 662 2004
rect 804 1939 806 2004
rect 948 1939 950 2004
rect 1092 1939 1094 2004
rect 1236 1939 1238 2004
rect 1380 1939 1382 2004
rect 1516 1939 1518 2004
rect 1652 1939 1654 2004
rect 1788 1939 1790 2004
rect 1934 2003 1940 2004
rect 1936 1939 1938 2003
rect 1976 1999 1978 2022
rect 3136 1999 3138 2023
rect 3272 1999 3274 2023
rect 3408 1999 3410 2023
rect 3544 1999 3546 2023
rect 3680 1999 3682 2023
rect 3798 2022 3804 2023
rect 3838 2027 3844 2028
rect 3838 2023 3839 2027
rect 3843 2023 3844 2027
rect 4662 2024 4663 2028
rect 4667 2024 4668 2028
rect 4662 2023 4668 2024
rect 4798 2028 4804 2029
rect 4798 2024 4799 2028
rect 4803 2024 4804 2028
rect 4798 2023 4804 2024
rect 4934 2028 4940 2029
rect 4934 2024 4935 2028
rect 4939 2024 4940 2028
rect 4934 2023 4940 2024
rect 5070 2028 5076 2029
rect 5070 2024 5071 2028
rect 5075 2024 5076 2028
rect 5070 2023 5076 2024
rect 5206 2028 5212 2029
rect 5206 2024 5207 2028
rect 5211 2024 5212 2028
rect 5206 2023 5212 2024
rect 5662 2027 5668 2028
rect 5662 2023 5663 2027
rect 5667 2023 5668 2027
rect 3838 2022 3844 2023
rect 3800 1999 3802 2022
rect 3840 1999 3842 2022
rect 4664 1999 4666 2023
rect 4800 1999 4802 2023
rect 4936 1999 4938 2023
rect 5072 1999 5074 2023
rect 5208 1999 5210 2023
rect 5662 2022 5668 2023
rect 5664 1999 5666 2022
rect 1975 1998 1979 1999
rect 1975 1993 1979 1994
rect 3127 1998 3131 1999
rect 3127 1993 3131 1994
rect 3135 1998 3139 1999
rect 3135 1993 3139 1994
rect 3263 1998 3267 1999
rect 3263 1993 3267 1994
rect 3271 1998 3275 1999
rect 3271 1993 3275 1994
rect 3399 1998 3403 1999
rect 3399 1993 3403 1994
rect 3407 1998 3411 1999
rect 3407 1993 3411 1994
rect 3535 1998 3539 1999
rect 3535 1993 3539 1994
rect 3543 1998 3547 1999
rect 3543 1993 3547 1994
rect 3671 1998 3675 1999
rect 3671 1993 3675 1994
rect 3679 1998 3683 1999
rect 3679 1993 3683 1994
rect 3799 1998 3803 1999
rect 3799 1993 3803 1994
rect 3839 1998 3843 1999
rect 3839 1993 3843 1994
rect 4663 1998 4667 1999
rect 4663 1993 4667 1994
rect 4799 1998 4803 1999
rect 4799 1993 4803 1994
rect 4863 1998 4867 1999
rect 4863 1993 4867 1994
rect 4935 1998 4939 1999
rect 4935 1993 4939 1994
rect 4999 1998 5003 1999
rect 4999 1993 5003 1994
rect 5071 1998 5075 1999
rect 5071 1993 5075 1994
rect 5135 1998 5139 1999
rect 5135 1993 5139 1994
rect 5207 1998 5211 1999
rect 5207 1993 5211 1994
rect 5271 1998 5275 1999
rect 5271 1993 5275 1994
rect 5407 1998 5411 1999
rect 5407 1993 5411 1994
rect 5543 1998 5547 1999
rect 5543 1993 5547 1994
rect 5663 1998 5667 1999
rect 5663 1993 5667 1994
rect 1976 1970 1978 1993
rect 1974 1969 1980 1970
rect 3128 1969 3130 1993
rect 3264 1969 3266 1993
rect 3400 1969 3402 1993
rect 3536 1969 3538 1993
rect 3672 1969 3674 1993
rect 3800 1970 3802 1993
rect 3840 1970 3842 1993
rect 3798 1969 3804 1970
rect 1974 1965 1975 1969
rect 1979 1965 1980 1969
rect 1974 1964 1980 1965
rect 3126 1968 3132 1969
rect 3126 1964 3127 1968
rect 3131 1964 3132 1968
rect 3126 1963 3132 1964
rect 3262 1968 3268 1969
rect 3262 1964 3263 1968
rect 3267 1964 3268 1968
rect 3262 1963 3268 1964
rect 3398 1968 3404 1969
rect 3398 1964 3399 1968
rect 3403 1964 3404 1968
rect 3398 1963 3404 1964
rect 3534 1968 3540 1969
rect 3534 1964 3535 1968
rect 3539 1964 3540 1968
rect 3534 1963 3540 1964
rect 3670 1968 3676 1969
rect 3670 1964 3671 1968
rect 3675 1964 3676 1968
rect 3798 1965 3799 1969
rect 3803 1965 3804 1969
rect 3798 1964 3804 1965
rect 3838 1969 3844 1970
rect 4864 1969 4866 1993
rect 5000 1969 5002 1993
rect 5136 1969 5138 1993
rect 5272 1969 5274 1993
rect 5408 1969 5410 1993
rect 5544 1969 5546 1993
rect 5664 1970 5666 1993
rect 5662 1969 5668 1970
rect 3838 1965 3839 1969
rect 3843 1965 3844 1969
rect 3838 1964 3844 1965
rect 4862 1968 4868 1969
rect 4862 1964 4863 1968
rect 4867 1964 4868 1968
rect 3670 1963 3676 1964
rect 4862 1963 4868 1964
rect 4998 1968 5004 1969
rect 4998 1964 4999 1968
rect 5003 1964 5004 1968
rect 4998 1963 5004 1964
rect 5134 1968 5140 1969
rect 5134 1964 5135 1968
rect 5139 1964 5140 1968
rect 5134 1963 5140 1964
rect 5270 1968 5276 1969
rect 5270 1964 5271 1968
rect 5275 1964 5276 1968
rect 5270 1963 5276 1964
rect 5406 1968 5412 1969
rect 5406 1964 5407 1968
rect 5411 1964 5412 1968
rect 5406 1963 5412 1964
rect 5542 1968 5548 1969
rect 5542 1964 5543 1968
rect 5547 1964 5548 1968
rect 5662 1965 5663 1969
rect 5667 1965 5668 1969
rect 5662 1964 5668 1965
rect 5542 1963 5548 1964
rect 3098 1953 3104 1954
rect 1974 1952 1980 1953
rect 1974 1948 1975 1952
rect 1979 1948 1980 1952
rect 3098 1949 3099 1953
rect 3103 1949 3104 1953
rect 3098 1948 3104 1949
rect 3234 1953 3240 1954
rect 3234 1949 3235 1953
rect 3239 1949 3240 1953
rect 3234 1948 3240 1949
rect 3370 1953 3376 1954
rect 3370 1949 3371 1953
rect 3375 1949 3376 1953
rect 3370 1948 3376 1949
rect 3506 1953 3512 1954
rect 3506 1949 3507 1953
rect 3511 1949 3512 1953
rect 3506 1948 3512 1949
rect 3642 1953 3648 1954
rect 4834 1953 4840 1954
rect 3642 1949 3643 1953
rect 3647 1949 3648 1953
rect 3642 1948 3648 1949
rect 3798 1952 3804 1953
rect 3798 1948 3799 1952
rect 3803 1948 3804 1952
rect 1974 1947 1980 1948
rect 111 1938 115 1939
rect 111 1933 115 1934
rect 187 1938 191 1939
rect 187 1933 191 1934
rect 243 1938 247 1939
rect 243 1933 247 1934
rect 379 1938 383 1939
rect 379 1933 383 1934
rect 515 1938 519 1939
rect 515 1933 519 1934
rect 587 1938 591 1939
rect 587 1933 591 1934
rect 659 1938 663 1939
rect 659 1933 663 1934
rect 803 1938 807 1939
rect 803 1933 807 1934
rect 811 1938 815 1939
rect 811 1933 815 1934
rect 947 1938 951 1939
rect 947 1933 951 1934
rect 1051 1938 1055 1939
rect 1051 1933 1055 1934
rect 1091 1938 1095 1939
rect 1091 1933 1095 1934
rect 1235 1938 1239 1939
rect 1235 1933 1239 1934
rect 1299 1938 1303 1939
rect 1299 1933 1303 1934
rect 1379 1938 1383 1939
rect 1379 1933 1383 1934
rect 1515 1938 1519 1939
rect 1515 1933 1519 1934
rect 1555 1938 1559 1939
rect 1555 1933 1559 1934
rect 1651 1938 1655 1939
rect 1651 1933 1655 1934
rect 1787 1938 1791 1939
rect 1787 1933 1791 1934
rect 1935 1938 1939 1939
rect 1935 1933 1939 1934
rect 112 1873 114 1933
rect 110 1872 116 1873
rect 188 1872 190 1933
rect 380 1872 382 1933
rect 588 1872 590 1933
rect 812 1872 814 1933
rect 1052 1872 1054 1933
rect 1300 1872 1302 1933
rect 1556 1872 1558 1933
rect 1788 1872 1790 1933
rect 1936 1873 1938 1933
rect 1976 1875 1978 1947
rect 3100 1875 3102 1948
rect 3236 1875 3238 1948
rect 3372 1875 3374 1948
rect 3508 1875 3510 1948
rect 3644 1875 3646 1948
rect 3798 1947 3804 1948
rect 3838 1952 3844 1953
rect 3838 1948 3839 1952
rect 3843 1948 3844 1952
rect 4834 1949 4835 1953
rect 4839 1949 4840 1953
rect 4834 1948 4840 1949
rect 4970 1953 4976 1954
rect 4970 1949 4971 1953
rect 4975 1949 4976 1953
rect 4970 1948 4976 1949
rect 5106 1953 5112 1954
rect 5106 1949 5107 1953
rect 5111 1949 5112 1953
rect 5106 1948 5112 1949
rect 5242 1953 5248 1954
rect 5242 1949 5243 1953
rect 5247 1949 5248 1953
rect 5242 1948 5248 1949
rect 5378 1953 5384 1954
rect 5378 1949 5379 1953
rect 5383 1949 5384 1953
rect 5378 1948 5384 1949
rect 5514 1953 5520 1954
rect 5514 1949 5515 1953
rect 5519 1949 5520 1953
rect 5514 1948 5520 1949
rect 5662 1952 5668 1953
rect 5662 1948 5663 1952
rect 5667 1948 5668 1952
rect 3838 1947 3844 1948
rect 3800 1875 3802 1947
rect 3840 1875 3842 1947
rect 4836 1875 4838 1948
rect 4972 1875 4974 1948
rect 5108 1875 5110 1948
rect 5244 1875 5246 1948
rect 5380 1875 5382 1948
rect 5516 1875 5518 1948
rect 5662 1947 5668 1948
rect 5664 1875 5666 1947
rect 1975 1874 1979 1875
rect 1934 1872 1940 1873
rect 110 1868 111 1872
rect 115 1868 116 1872
rect 110 1867 116 1868
rect 186 1871 192 1872
rect 186 1867 187 1871
rect 191 1867 192 1871
rect 186 1866 192 1867
rect 378 1871 384 1872
rect 378 1867 379 1871
rect 383 1867 384 1871
rect 378 1866 384 1867
rect 586 1871 592 1872
rect 586 1867 587 1871
rect 591 1867 592 1871
rect 586 1866 592 1867
rect 810 1871 816 1872
rect 810 1867 811 1871
rect 815 1867 816 1871
rect 810 1866 816 1867
rect 1050 1871 1056 1872
rect 1050 1867 1051 1871
rect 1055 1867 1056 1871
rect 1050 1866 1056 1867
rect 1298 1871 1304 1872
rect 1298 1867 1299 1871
rect 1303 1867 1304 1871
rect 1298 1866 1304 1867
rect 1554 1871 1560 1872
rect 1554 1867 1555 1871
rect 1559 1867 1560 1871
rect 1554 1866 1560 1867
rect 1786 1871 1792 1872
rect 1786 1867 1787 1871
rect 1791 1867 1792 1871
rect 1934 1868 1935 1872
rect 1939 1868 1940 1872
rect 1975 1869 1979 1870
rect 1995 1874 1999 1875
rect 1995 1869 1999 1870
rect 2227 1874 2231 1875
rect 2227 1869 2231 1870
rect 2467 1874 2471 1875
rect 2467 1869 2471 1870
rect 2691 1874 2695 1875
rect 2691 1869 2695 1870
rect 2907 1874 2911 1875
rect 2907 1869 2911 1870
rect 3099 1874 3103 1875
rect 3099 1869 3103 1870
rect 3107 1874 3111 1875
rect 3107 1869 3111 1870
rect 3235 1874 3239 1875
rect 3235 1869 3239 1870
rect 3299 1874 3303 1875
rect 3299 1869 3303 1870
rect 3371 1874 3375 1875
rect 3371 1869 3375 1870
rect 3483 1874 3487 1875
rect 3483 1869 3487 1870
rect 3507 1874 3511 1875
rect 3507 1869 3511 1870
rect 3643 1874 3647 1875
rect 3643 1869 3647 1870
rect 3651 1874 3655 1875
rect 3651 1869 3655 1870
rect 3799 1874 3803 1875
rect 3799 1869 3803 1870
rect 3839 1874 3843 1875
rect 3839 1869 3843 1870
rect 4675 1874 4679 1875
rect 4675 1869 4679 1870
rect 4819 1874 4823 1875
rect 4819 1869 4823 1870
rect 4835 1874 4839 1875
rect 4835 1869 4839 1870
rect 4963 1874 4967 1875
rect 4963 1869 4967 1870
rect 4971 1874 4975 1875
rect 4971 1869 4975 1870
rect 5107 1874 5111 1875
rect 5107 1869 5111 1870
rect 5243 1874 5247 1875
rect 5243 1869 5247 1870
rect 5379 1874 5383 1875
rect 5379 1869 5383 1870
rect 5515 1874 5519 1875
rect 5515 1869 5519 1870
rect 5663 1874 5667 1875
rect 5663 1869 5667 1870
rect 1934 1867 1940 1868
rect 1786 1866 1792 1867
rect 214 1856 220 1857
rect 110 1855 116 1856
rect 110 1851 111 1855
rect 115 1851 116 1855
rect 214 1852 215 1856
rect 219 1852 220 1856
rect 214 1851 220 1852
rect 406 1856 412 1857
rect 406 1852 407 1856
rect 411 1852 412 1856
rect 406 1851 412 1852
rect 614 1856 620 1857
rect 614 1852 615 1856
rect 619 1852 620 1856
rect 614 1851 620 1852
rect 838 1856 844 1857
rect 838 1852 839 1856
rect 843 1852 844 1856
rect 838 1851 844 1852
rect 1078 1856 1084 1857
rect 1078 1852 1079 1856
rect 1083 1852 1084 1856
rect 1078 1851 1084 1852
rect 1326 1856 1332 1857
rect 1326 1852 1327 1856
rect 1331 1852 1332 1856
rect 1326 1851 1332 1852
rect 1582 1856 1588 1857
rect 1582 1852 1583 1856
rect 1587 1852 1588 1856
rect 1582 1851 1588 1852
rect 1814 1856 1820 1857
rect 1814 1852 1815 1856
rect 1819 1852 1820 1856
rect 1814 1851 1820 1852
rect 1934 1855 1940 1856
rect 1934 1851 1935 1855
rect 1939 1851 1940 1855
rect 110 1850 116 1851
rect 112 1819 114 1850
rect 216 1819 218 1851
rect 408 1819 410 1851
rect 616 1819 618 1851
rect 840 1819 842 1851
rect 1080 1819 1082 1851
rect 1328 1819 1330 1851
rect 1584 1819 1586 1851
rect 1816 1819 1818 1851
rect 1934 1850 1940 1851
rect 1936 1819 1938 1850
rect 111 1818 115 1819
rect 111 1813 115 1814
rect 159 1818 163 1819
rect 159 1813 163 1814
rect 215 1818 219 1819
rect 215 1813 219 1814
rect 375 1818 379 1819
rect 375 1813 379 1814
rect 407 1818 411 1819
rect 407 1813 411 1814
rect 591 1818 595 1819
rect 591 1813 595 1814
rect 615 1818 619 1819
rect 615 1813 619 1814
rect 799 1818 803 1819
rect 799 1813 803 1814
rect 839 1818 843 1819
rect 839 1813 843 1814
rect 999 1818 1003 1819
rect 999 1813 1003 1814
rect 1079 1818 1083 1819
rect 1079 1813 1083 1814
rect 1191 1818 1195 1819
rect 1191 1813 1195 1814
rect 1327 1818 1331 1819
rect 1327 1813 1331 1814
rect 1383 1818 1387 1819
rect 1383 1813 1387 1814
rect 1575 1818 1579 1819
rect 1575 1813 1579 1814
rect 1583 1818 1587 1819
rect 1583 1813 1587 1814
rect 1815 1818 1819 1819
rect 1815 1813 1819 1814
rect 1935 1818 1939 1819
rect 1935 1813 1939 1814
rect 112 1790 114 1813
rect 110 1789 116 1790
rect 160 1789 162 1813
rect 376 1789 378 1813
rect 592 1789 594 1813
rect 800 1789 802 1813
rect 1000 1789 1002 1813
rect 1192 1789 1194 1813
rect 1384 1789 1386 1813
rect 1576 1789 1578 1813
rect 1936 1790 1938 1813
rect 1976 1809 1978 1869
rect 1974 1808 1980 1809
rect 1996 1808 1998 1869
rect 2228 1808 2230 1869
rect 2468 1808 2470 1869
rect 2692 1808 2694 1869
rect 2908 1808 2910 1869
rect 3108 1808 3110 1869
rect 3300 1808 3302 1869
rect 3484 1808 3486 1869
rect 3652 1808 3654 1869
rect 3800 1809 3802 1869
rect 3840 1809 3842 1869
rect 3798 1808 3804 1809
rect 1974 1804 1975 1808
rect 1979 1804 1980 1808
rect 1974 1803 1980 1804
rect 1994 1807 2000 1808
rect 1994 1803 1995 1807
rect 1999 1803 2000 1807
rect 1994 1802 2000 1803
rect 2226 1807 2232 1808
rect 2226 1803 2227 1807
rect 2231 1803 2232 1807
rect 2226 1802 2232 1803
rect 2466 1807 2472 1808
rect 2466 1803 2467 1807
rect 2471 1803 2472 1807
rect 2466 1802 2472 1803
rect 2690 1807 2696 1808
rect 2690 1803 2691 1807
rect 2695 1803 2696 1807
rect 2690 1802 2696 1803
rect 2906 1807 2912 1808
rect 2906 1803 2907 1807
rect 2911 1803 2912 1807
rect 2906 1802 2912 1803
rect 3106 1807 3112 1808
rect 3106 1803 3107 1807
rect 3111 1803 3112 1807
rect 3106 1802 3112 1803
rect 3298 1807 3304 1808
rect 3298 1803 3299 1807
rect 3303 1803 3304 1807
rect 3298 1802 3304 1803
rect 3482 1807 3488 1808
rect 3482 1803 3483 1807
rect 3487 1803 3488 1807
rect 3482 1802 3488 1803
rect 3650 1807 3656 1808
rect 3650 1803 3651 1807
rect 3655 1803 3656 1807
rect 3798 1804 3799 1808
rect 3803 1804 3804 1808
rect 3798 1803 3804 1804
rect 3838 1808 3844 1809
rect 4676 1808 4678 1869
rect 4820 1808 4822 1869
rect 4964 1808 4966 1869
rect 5108 1808 5110 1869
rect 5244 1808 5246 1869
rect 5380 1808 5382 1869
rect 5516 1808 5518 1869
rect 5664 1809 5666 1869
rect 5662 1808 5668 1809
rect 3838 1804 3839 1808
rect 3843 1804 3844 1808
rect 3838 1803 3844 1804
rect 4674 1807 4680 1808
rect 4674 1803 4675 1807
rect 4679 1803 4680 1807
rect 3650 1802 3656 1803
rect 4674 1802 4680 1803
rect 4818 1807 4824 1808
rect 4818 1803 4819 1807
rect 4823 1803 4824 1807
rect 4818 1802 4824 1803
rect 4962 1807 4968 1808
rect 4962 1803 4963 1807
rect 4967 1803 4968 1807
rect 4962 1802 4968 1803
rect 5106 1807 5112 1808
rect 5106 1803 5107 1807
rect 5111 1803 5112 1807
rect 5106 1802 5112 1803
rect 5242 1807 5248 1808
rect 5242 1803 5243 1807
rect 5247 1803 5248 1807
rect 5242 1802 5248 1803
rect 5378 1807 5384 1808
rect 5378 1803 5379 1807
rect 5383 1803 5384 1807
rect 5378 1802 5384 1803
rect 5514 1807 5520 1808
rect 5514 1803 5515 1807
rect 5519 1803 5520 1807
rect 5662 1804 5663 1808
rect 5667 1804 5668 1808
rect 5662 1803 5668 1804
rect 5514 1802 5520 1803
rect 2022 1792 2028 1793
rect 1974 1791 1980 1792
rect 1934 1789 1940 1790
rect 110 1785 111 1789
rect 115 1785 116 1789
rect 110 1784 116 1785
rect 158 1788 164 1789
rect 158 1784 159 1788
rect 163 1784 164 1788
rect 158 1783 164 1784
rect 374 1788 380 1789
rect 374 1784 375 1788
rect 379 1784 380 1788
rect 374 1783 380 1784
rect 590 1788 596 1789
rect 590 1784 591 1788
rect 595 1784 596 1788
rect 590 1783 596 1784
rect 798 1788 804 1789
rect 798 1784 799 1788
rect 803 1784 804 1788
rect 798 1783 804 1784
rect 998 1788 1004 1789
rect 998 1784 999 1788
rect 1003 1784 1004 1788
rect 998 1783 1004 1784
rect 1190 1788 1196 1789
rect 1190 1784 1191 1788
rect 1195 1784 1196 1788
rect 1190 1783 1196 1784
rect 1382 1788 1388 1789
rect 1382 1784 1383 1788
rect 1387 1784 1388 1788
rect 1382 1783 1388 1784
rect 1574 1788 1580 1789
rect 1574 1784 1575 1788
rect 1579 1784 1580 1788
rect 1934 1785 1935 1789
rect 1939 1785 1940 1789
rect 1974 1787 1975 1791
rect 1979 1787 1980 1791
rect 2022 1788 2023 1792
rect 2027 1788 2028 1792
rect 2022 1787 2028 1788
rect 2254 1792 2260 1793
rect 2254 1788 2255 1792
rect 2259 1788 2260 1792
rect 2254 1787 2260 1788
rect 2494 1792 2500 1793
rect 2494 1788 2495 1792
rect 2499 1788 2500 1792
rect 2494 1787 2500 1788
rect 2718 1792 2724 1793
rect 2718 1788 2719 1792
rect 2723 1788 2724 1792
rect 2718 1787 2724 1788
rect 2934 1792 2940 1793
rect 2934 1788 2935 1792
rect 2939 1788 2940 1792
rect 2934 1787 2940 1788
rect 3134 1792 3140 1793
rect 3134 1788 3135 1792
rect 3139 1788 3140 1792
rect 3134 1787 3140 1788
rect 3326 1792 3332 1793
rect 3326 1788 3327 1792
rect 3331 1788 3332 1792
rect 3326 1787 3332 1788
rect 3510 1792 3516 1793
rect 3510 1788 3511 1792
rect 3515 1788 3516 1792
rect 3510 1787 3516 1788
rect 3678 1792 3684 1793
rect 4702 1792 4708 1793
rect 3678 1788 3679 1792
rect 3683 1788 3684 1792
rect 3678 1787 3684 1788
rect 3798 1791 3804 1792
rect 3798 1787 3799 1791
rect 3803 1787 3804 1791
rect 1974 1786 1980 1787
rect 1934 1784 1940 1785
rect 1574 1783 1580 1784
rect 130 1773 136 1774
rect 110 1772 116 1773
rect 110 1768 111 1772
rect 115 1768 116 1772
rect 130 1769 131 1773
rect 135 1769 136 1773
rect 130 1768 136 1769
rect 346 1773 352 1774
rect 346 1769 347 1773
rect 351 1769 352 1773
rect 346 1768 352 1769
rect 562 1773 568 1774
rect 562 1769 563 1773
rect 567 1769 568 1773
rect 562 1768 568 1769
rect 770 1773 776 1774
rect 770 1769 771 1773
rect 775 1769 776 1773
rect 770 1768 776 1769
rect 970 1773 976 1774
rect 970 1769 971 1773
rect 975 1769 976 1773
rect 970 1768 976 1769
rect 1162 1773 1168 1774
rect 1162 1769 1163 1773
rect 1167 1769 1168 1773
rect 1162 1768 1168 1769
rect 1354 1773 1360 1774
rect 1354 1769 1355 1773
rect 1359 1769 1360 1773
rect 1354 1768 1360 1769
rect 1546 1773 1552 1774
rect 1546 1769 1547 1773
rect 1551 1769 1552 1773
rect 1546 1768 1552 1769
rect 1934 1772 1940 1773
rect 1934 1768 1935 1772
rect 1939 1768 1940 1772
rect 110 1767 116 1768
rect 112 1683 114 1767
rect 132 1683 134 1768
rect 348 1683 350 1768
rect 564 1683 566 1768
rect 772 1683 774 1768
rect 972 1683 974 1768
rect 1164 1683 1166 1768
rect 1356 1683 1358 1768
rect 1548 1683 1550 1768
rect 1934 1767 1940 1768
rect 1936 1683 1938 1767
rect 1976 1755 1978 1786
rect 2024 1755 2026 1787
rect 2256 1755 2258 1787
rect 2496 1755 2498 1787
rect 2720 1755 2722 1787
rect 2936 1755 2938 1787
rect 3136 1755 3138 1787
rect 3328 1755 3330 1787
rect 3512 1755 3514 1787
rect 3680 1755 3682 1787
rect 3798 1786 3804 1787
rect 3838 1791 3844 1792
rect 3838 1787 3839 1791
rect 3843 1787 3844 1791
rect 4702 1788 4703 1792
rect 4707 1788 4708 1792
rect 4702 1787 4708 1788
rect 4846 1792 4852 1793
rect 4846 1788 4847 1792
rect 4851 1788 4852 1792
rect 4846 1787 4852 1788
rect 4990 1792 4996 1793
rect 4990 1788 4991 1792
rect 4995 1788 4996 1792
rect 4990 1787 4996 1788
rect 5134 1792 5140 1793
rect 5134 1788 5135 1792
rect 5139 1788 5140 1792
rect 5134 1787 5140 1788
rect 5270 1792 5276 1793
rect 5270 1788 5271 1792
rect 5275 1788 5276 1792
rect 5270 1787 5276 1788
rect 5406 1792 5412 1793
rect 5406 1788 5407 1792
rect 5411 1788 5412 1792
rect 5406 1787 5412 1788
rect 5542 1792 5548 1793
rect 5542 1788 5543 1792
rect 5547 1788 5548 1792
rect 5542 1787 5548 1788
rect 5662 1791 5668 1792
rect 5662 1787 5663 1791
rect 5667 1787 5668 1791
rect 3838 1786 3844 1787
rect 3800 1755 3802 1786
rect 1975 1754 1979 1755
rect 1975 1749 1979 1750
rect 2023 1754 2027 1755
rect 2023 1749 2027 1750
rect 2159 1754 2163 1755
rect 2159 1749 2163 1750
rect 2255 1754 2259 1755
rect 2255 1749 2259 1750
rect 2311 1754 2315 1755
rect 2311 1749 2315 1750
rect 2471 1754 2475 1755
rect 2471 1749 2475 1750
rect 2495 1754 2499 1755
rect 2495 1749 2499 1750
rect 2639 1754 2643 1755
rect 2639 1749 2643 1750
rect 2719 1754 2723 1755
rect 2719 1749 2723 1750
rect 2807 1754 2811 1755
rect 2807 1749 2811 1750
rect 2935 1754 2939 1755
rect 2935 1749 2939 1750
rect 2975 1754 2979 1755
rect 2975 1749 2979 1750
rect 3135 1754 3139 1755
rect 3135 1749 3139 1750
rect 3151 1754 3155 1755
rect 3151 1749 3155 1750
rect 3327 1754 3331 1755
rect 3327 1749 3331 1750
rect 3511 1754 3515 1755
rect 3511 1749 3515 1750
rect 3679 1754 3683 1755
rect 3679 1749 3683 1750
rect 3799 1754 3803 1755
rect 3799 1749 3803 1750
rect 1976 1726 1978 1749
rect 1974 1725 1980 1726
rect 2024 1725 2026 1749
rect 2160 1725 2162 1749
rect 2312 1725 2314 1749
rect 2472 1725 2474 1749
rect 2640 1725 2642 1749
rect 2808 1725 2810 1749
rect 2976 1725 2978 1749
rect 3152 1725 3154 1749
rect 3800 1726 3802 1749
rect 3840 1747 3842 1786
rect 4704 1747 4706 1787
rect 4848 1747 4850 1787
rect 4992 1747 4994 1787
rect 5136 1747 5138 1787
rect 5272 1747 5274 1787
rect 5408 1747 5410 1787
rect 5544 1747 5546 1787
rect 5662 1786 5668 1787
rect 5664 1747 5666 1786
rect 3839 1746 3843 1747
rect 3839 1741 3843 1742
rect 3887 1746 3891 1747
rect 3887 1741 3891 1742
rect 4079 1746 4083 1747
rect 4079 1741 4083 1742
rect 4303 1746 4307 1747
rect 4303 1741 4307 1742
rect 4535 1746 4539 1747
rect 4535 1741 4539 1742
rect 4703 1746 4707 1747
rect 4703 1741 4707 1742
rect 4775 1746 4779 1747
rect 4775 1741 4779 1742
rect 4847 1746 4851 1747
rect 4847 1741 4851 1742
rect 4991 1746 4995 1747
rect 4991 1741 4995 1742
rect 5023 1746 5027 1747
rect 5023 1741 5027 1742
rect 5135 1746 5139 1747
rect 5135 1741 5139 1742
rect 5271 1746 5275 1747
rect 5271 1741 5275 1742
rect 5279 1746 5283 1747
rect 5279 1741 5283 1742
rect 5407 1746 5411 1747
rect 5407 1741 5411 1742
rect 5535 1746 5539 1747
rect 5535 1741 5539 1742
rect 5543 1746 5547 1747
rect 5543 1741 5547 1742
rect 5663 1746 5667 1747
rect 5663 1741 5667 1742
rect 3798 1725 3804 1726
rect 1974 1721 1975 1725
rect 1979 1721 1980 1725
rect 1974 1720 1980 1721
rect 2022 1724 2028 1725
rect 2022 1720 2023 1724
rect 2027 1720 2028 1724
rect 2022 1719 2028 1720
rect 2158 1724 2164 1725
rect 2158 1720 2159 1724
rect 2163 1720 2164 1724
rect 2158 1719 2164 1720
rect 2310 1724 2316 1725
rect 2310 1720 2311 1724
rect 2315 1720 2316 1724
rect 2310 1719 2316 1720
rect 2470 1724 2476 1725
rect 2470 1720 2471 1724
rect 2475 1720 2476 1724
rect 2470 1719 2476 1720
rect 2638 1724 2644 1725
rect 2638 1720 2639 1724
rect 2643 1720 2644 1724
rect 2638 1719 2644 1720
rect 2806 1724 2812 1725
rect 2806 1720 2807 1724
rect 2811 1720 2812 1724
rect 2806 1719 2812 1720
rect 2974 1724 2980 1725
rect 2974 1720 2975 1724
rect 2979 1720 2980 1724
rect 2974 1719 2980 1720
rect 3150 1724 3156 1725
rect 3150 1720 3151 1724
rect 3155 1720 3156 1724
rect 3798 1721 3799 1725
rect 3803 1721 3804 1725
rect 3798 1720 3804 1721
rect 3150 1719 3156 1720
rect 3840 1718 3842 1741
rect 3838 1717 3844 1718
rect 3888 1717 3890 1741
rect 4080 1717 4082 1741
rect 4304 1717 4306 1741
rect 4536 1717 4538 1741
rect 4776 1717 4778 1741
rect 5024 1717 5026 1741
rect 5280 1717 5282 1741
rect 5536 1717 5538 1741
rect 5664 1718 5666 1741
rect 5662 1717 5668 1718
rect 3838 1713 3839 1717
rect 3843 1713 3844 1717
rect 3838 1712 3844 1713
rect 3886 1716 3892 1717
rect 3886 1712 3887 1716
rect 3891 1712 3892 1716
rect 3886 1711 3892 1712
rect 4078 1716 4084 1717
rect 4078 1712 4079 1716
rect 4083 1712 4084 1716
rect 4078 1711 4084 1712
rect 4302 1716 4308 1717
rect 4302 1712 4303 1716
rect 4307 1712 4308 1716
rect 4302 1711 4308 1712
rect 4534 1716 4540 1717
rect 4534 1712 4535 1716
rect 4539 1712 4540 1716
rect 4534 1711 4540 1712
rect 4774 1716 4780 1717
rect 4774 1712 4775 1716
rect 4779 1712 4780 1716
rect 4774 1711 4780 1712
rect 5022 1716 5028 1717
rect 5022 1712 5023 1716
rect 5027 1712 5028 1716
rect 5022 1711 5028 1712
rect 5278 1716 5284 1717
rect 5278 1712 5279 1716
rect 5283 1712 5284 1716
rect 5278 1711 5284 1712
rect 5534 1716 5540 1717
rect 5534 1712 5535 1716
rect 5539 1712 5540 1716
rect 5662 1713 5663 1717
rect 5667 1713 5668 1717
rect 5662 1712 5668 1713
rect 5534 1711 5540 1712
rect 1994 1709 2000 1710
rect 1974 1708 1980 1709
rect 1974 1704 1975 1708
rect 1979 1704 1980 1708
rect 1994 1705 1995 1709
rect 1999 1705 2000 1709
rect 1994 1704 2000 1705
rect 2130 1709 2136 1710
rect 2130 1705 2131 1709
rect 2135 1705 2136 1709
rect 2130 1704 2136 1705
rect 2282 1709 2288 1710
rect 2282 1705 2283 1709
rect 2287 1705 2288 1709
rect 2282 1704 2288 1705
rect 2442 1709 2448 1710
rect 2442 1705 2443 1709
rect 2447 1705 2448 1709
rect 2442 1704 2448 1705
rect 2610 1709 2616 1710
rect 2610 1705 2611 1709
rect 2615 1705 2616 1709
rect 2610 1704 2616 1705
rect 2778 1709 2784 1710
rect 2778 1705 2779 1709
rect 2783 1705 2784 1709
rect 2778 1704 2784 1705
rect 2946 1709 2952 1710
rect 2946 1705 2947 1709
rect 2951 1705 2952 1709
rect 2946 1704 2952 1705
rect 3122 1709 3128 1710
rect 3122 1705 3123 1709
rect 3127 1705 3128 1709
rect 3122 1704 3128 1705
rect 3798 1708 3804 1709
rect 3798 1704 3799 1708
rect 3803 1704 3804 1708
rect 1974 1703 1980 1704
rect 111 1682 115 1683
rect 111 1677 115 1678
rect 131 1682 135 1683
rect 131 1677 135 1678
rect 347 1682 351 1683
rect 347 1677 351 1678
rect 395 1682 399 1683
rect 395 1677 399 1678
rect 563 1682 567 1683
rect 563 1677 567 1678
rect 683 1682 687 1683
rect 683 1677 687 1678
rect 771 1682 775 1683
rect 771 1677 775 1678
rect 971 1682 975 1683
rect 971 1677 975 1678
rect 979 1682 983 1683
rect 979 1677 983 1678
rect 1163 1682 1167 1683
rect 1163 1677 1167 1678
rect 1275 1682 1279 1683
rect 1275 1677 1279 1678
rect 1355 1682 1359 1683
rect 1355 1677 1359 1678
rect 1547 1682 1551 1683
rect 1547 1677 1551 1678
rect 1935 1682 1939 1683
rect 1935 1677 1939 1678
rect 112 1617 114 1677
rect 110 1616 116 1617
rect 132 1616 134 1677
rect 396 1616 398 1677
rect 684 1616 686 1677
rect 980 1616 982 1677
rect 1276 1616 1278 1677
rect 1936 1617 1938 1677
rect 1976 1635 1978 1703
rect 1996 1635 1998 1704
rect 2132 1635 2134 1704
rect 2284 1635 2286 1704
rect 2444 1635 2446 1704
rect 2612 1635 2614 1704
rect 2780 1635 2782 1704
rect 2948 1635 2950 1704
rect 3124 1635 3126 1704
rect 3798 1703 3804 1704
rect 3800 1635 3802 1703
rect 3858 1701 3864 1702
rect 3838 1700 3844 1701
rect 3838 1696 3839 1700
rect 3843 1696 3844 1700
rect 3858 1697 3859 1701
rect 3863 1697 3864 1701
rect 3858 1696 3864 1697
rect 4050 1701 4056 1702
rect 4050 1697 4051 1701
rect 4055 1697 4056 1701
rect 4050 1696 4056 1697
rect 4274 1701 4280 1702
rect 4274 1697 4275 1701
rect 4279 1697 4280 1701
rect 4274 1696 4280 1697
rect 4506 1701 4512 1702
rect 4506 1697 4507 1701
rect 4511 1697 4512 1701
rect 4506 1696 4512 1697
rect 4746 1701 4752 1702
rect 4746 1697 4747 1701
rect 4751 1697 4752 1701
rect 4746 1696 4752 1697
rect 4994 1701 5000 1702
rect 4994 1697 4995 1701
rect 4999 1697 5000 1701
rect 4994 1696 5000 1697
rect 5250 1701 5256 1702
rect 5250 1697 5251 1701
rect 5255 1697 5256 1701
rect 5250 1696 5256 1697
rect 5506 1701 5512 1702
rect 5506 1697 5507 1701
rect 5511 1697 5512 1701
rect 5506 1696 5512 1697
rect 5662 1700 5668 1701
rect 5662 1696 5663 1700
rect 5667 1696 5668 1700
rect 3838 1695 3844 1696
rect 3840 1635 3842 1695
rect 3860 1635 3862 1696
rect 4052 1635 4054 1696
rect 4276 1635 4278 1696
rect 4508 1635 4510 1696
rect 4748 1635 4750 1696
rect 4996 1635 4998 1696
rect 5252 1635 5254 1696
rect 5508 1635 5510 1696
rect 5662 1695 5668 1696
rect 5664 1635 5666 1695
rect 1975 1634 1979 1635
rect 1975 1629 1979 1630
rect 1995 1634 1999 1635
rect 1995 1629 1999 1630
rect 2091 1634 2095 1635
rect 2091 1629 2095 1630
rect 2131 1634 2135 1635
rect 2131 1629 2135 1630
rect 2227 1634 2231 1635
rect 2227 1629 2231 1630
rect 2283 1634 2287 1635
rect 2283 1629 2287 1630
rect 2363 1634 2367 1635
rect 2363 1629 2367 1630
rect 2443 1634 2447 1635
rect 2443 1629 2447 1630
rect 2499 1634 2503 1635
rect 2499 1629 2503 1630
rect 2611 1634 2615 1635
rect 2611 1629 2615 1630
rect 2635 1634 2639 1635
rect 2635 1629 2639 1630
rect 2771 1634 2775 1635
rect 2771 1629 2775 1630
rect 2779 1634 2783 1635
rect 2779 1629 2783 1630
rect 2907 1634 2911 1635
rect 2907 1629 2911 1630
rect 2947 1634 2951 1635
rect 2947 1629 2951 1630
rect 3043 1634 3047 1635
rect 3043 1629 3047 1630
rect 3123 1634 3127 1635
rect 3123 1629 3127 1630
rect 3179 1634 3183 1635
rect 3179 1629 3183 1630
rect 3799 1634 3803 1635
rect 3799 1629 3803 1630
rect 3839 1634 3843 1635
rect 3839 1629 3843 1630
rect 3859 1634 3863 1635
rect 3859 1629 3863 1630
rect 3995 1634 3999 1635
rect 3995 1629 3999 1630
rect 4051 1634 4055 1635
rect 4051 1629 4055 1630
rect 4155 1634 4159 1635
rect 4155 1629 4159 1630
rect 4275 1634 4279 1635
rect 4275 1629 4279 1630
rect 4355 1634 4359 1635
rect 4355 1629 4359 1630
rect 4507 1634 4511 1635
rect 4507 1629 4511 1630
rect 4587 1634 4591 1635
rect 4587 1629 4591 1630
rect 4747 1634 4751 1635
rect 4747 1629 4751 1630
rect 4851 1634 4855 1635
rect 4851 1629 4855 1630
rect 4995 1634 4999 1635
rect 4995 1629 4999 1630
rect 5131 1634 5135 1635
rect 5131 1629 5135 1630
rect 5251 1634 5255 1635
rect 5251 1629 5255 1630
rect 5419 1634 5423 1635
rect 5419 1629 5423 1630
rect 5507 1634 5511 1635
rect 5507 1629 5511 1630
rect 5663 1634 5667 1635
rect 5663 1629 5667 1630
rect 1934 1616 1940 1617
rect 110 1612 111 1616
rect 115 1612 116 1616
rect 110 1611 116 1612
rect 130 1615 136 1616
rect 130 1611 131 1615
rect 135 1611 136 1615
rect 130 1610 136 1611
rect 394 1615 400 1616
rect 394 1611 395 1615
rect 399 1611 400 1615
rect 394 1610 400 1611
rect 682 1615 688 1616
rect 682 1611 683 1615
rect 687 1611 688 1615
rect 682 1610 688 1611
rect 978 1615 984 1616
rect 978 1611 979 1615
rect 983 1611 984 1615
rect 978 1610 984 1611
rect 1274 1615 1280 1616
rect 1274 1611 1275 1615
rect 1279 1611 1280 1615
rect 1934 1612 1935 1616
rect 1939 1612 1940 1616
rect 1934 1611 1940 1612
rect 1274 1610 1280 1611
rect 158 1600 164 1601
rect 110 1599 116 1600
rect 110 1595 111 1599
rect 115 1595 116 1599
rect 158 1596 159 1600
rect 163 1596 164 1600
rect 158 1595 164 1596
rect 422 1600 428 1601
rect 422 1596 423 1600
rect 427 1596 428 1600
rect 422 1595 428 1596
rect 710 1600 716 1601
rect 710 1596 711 1600
rect 715 1596 716 1600
rect 710 1595 716 1596
rect 1006 1600 1012 1601
rect 1006 1596 1007 1600
rect 1011 1596 1012 1600
rect 1006 1595 1012 1596
rect 1302 1600 1308 1601
rect 1302 1596 1303 1600
rect 1307 1596 1308 1600
rect 1302 1595 1308 1596
rect 1934 1599 1940 1600
rect 1934 1595 1935 1599
rect 1939 1595 1940 1599
rect 110 1594 116 1595
rect 112 1559 114 1594
rect 160 1559 162 1595
rect 424 1559 426 1595
rect 712 1559 714 1595
rect 1008 1559 1010 1595
rect 1304 1559 1306 1595
rect 1934 1594 1940 1595
rect 1936 1559 1938 1594
rect 1976 1569 1978 1629
rect 1974 1568 1980 1569
rect 2092 1568 2094 1629
rect 2228 1568 2230 1629
rect 2364 1568 2366 1629
rect 2500 1568 2502 1629
rect 2636 1568 2638 1629
rect 2772 1568 2774 1629
rect 2908 1568 2910 1629
rect 3044 1568 3046 1629
rect 3180 1568 3182 1629
rect 3800 1569 3802 1629
rect 3840 1569 3842 1629
rect 3798 1568 3804 1569
rect 1974 1564 1975 1568
rect 1979 1564 1980 1568
rect 1974 1563 1980 1564
rect 2090 1567 2096 1568
rect 2090 1563 2091 1567
rect 2095 1563 2096 1567
rect 2090 1562 2096 1563
rect 2226 1567 2232 1568
rect 2226 1563 2227 1567
rect 2231 1563 2232 1567
rect 2226 1562 2232 1563
rect 2362 1567 2368 1568
rect 2362 1563 2363 1567
rect 2367 1563 2368 1567
rect 2362 1562 2368 1563
rect 2498 1567 2504 1568
rect 2498 1563 2499 1567
rect 2503 1563 2504 1567
rect 2498 1562 2504 1563
rect 2634 1567 2640 1568
rect 2634 1563 2635 1567
rect 2639 1563 2640 1567
rect 2634 1562 2640 1563
rect 2770 1567 2776 1568
rect 2770 1563 2771 1567
rect 2775 1563 2776 1567
rect 2770 1562 2776 1563
rect 2906 1567 2912 1568
rect 2906 1563 2907 1567
rect 2911 1563 2912 1567
rect 2906 1562 2912 1563
rect 3042 1567 3048 1568
rect 3042 1563 3043 1567
rect 3047 1563 3048 1567
rect 3042 1562 3048 1563
rect 3178 1567 3184 1568
rect 3178 1563 3179 1567
rect 3183 1563 3184 1567
rect 3798 1564 3799 1568
rect 3803 1564 3804 1568
rect 3798 1563 3804 1564
rect 3838 1568 3844 1569
rect 3860 1568 3862 1629
rect 3996 1568 3998 1629
rect 4156 1568 4158 1629
rect 4356 1568 4358 1629
rect 4588 1568 4590 1629
rect 4852 1568 4854 1629
rect 5132 1568 5134 1629
rect 5420 1568 5422 1629
rect 5664 1569 5666 1629
rect 5662 1568 5668 1569
rect 3838 1564 3839 1568
rect 3843 1564 3844 1568
rect 3838 1563 3844 1564
rect 3858 1567 3864 1568
rect 3858 1563 3859 1567
rect 3863 1563 3864 1567
rect 3178 1562 3184 1563
rect 3858 1562 3864 1563
rect 3994 1567 4000 1568
rect 3994 1563 3995 1567
rect 3999 1563 4000 1567
rect 3994 1562 4000 1563
rect 4154 1567 4160 1568
rect 4154 1563 4155 1567
rect 4159 1563 4160 1567
rect 4154 1562 4160 1563
rect 4354 1567 4360 1568
rect 4354 1563 4355 1567
rect 4359 1563 4360 1567
rect 4354 1562 4360 1563
rect 4586 1567 4592 1568
rect 4586 1563 4587 1567
rect 4591 1563 4592 1567
rect 4586 1562 4592 1563
rect 4850 1567 4856 1568
rect 4850 1563 4851 1567
rect 4855 1563 4856 1567
rect 4850 1562 4856 1563
rect 5130 1567 5136 1568
rect 5130 1563 5131 1567
rect 5135 1563 5136 1567
rect 5130 1562 5136 1563
rect 5418 1567 5424 1568
rect 5418 1563 5419 1567
rect 5423 1563 5424 1567
rect 5662 1564 5663 1568
rect 5667 1564 5668 1568
rect 5662 1563 5668 1564
rect 5418 1562 5424 1563
rect 111 1558 115 1559
rect 111 1553 115 1554
rect 159 1558 163 1559
rect 159 1553 163 1554
rect 375 1558 379 1559
rect 375 1553 379 1554
rect 423 1558 427 1559
rect 423 1553 427 1554
rect 607 1558 611 1559
rect 607 1553 611 1554
rect 711 1558 715 1559
rect 711 1553 715 1554
rect 839 1558 843 1559
rect 839 1553 843 1554
rect 1007 1558 1011 1559
rect 1007 1553 1011 1554
rect 1071 1558 1075 1559
rect 1071 1553 1075 1554
rect 1303 1558 1307 1559
rect 1303 1553 1307 1554
rect 1935 1558 1939 1559
rect 1935 1553 1939 1554
rect 112 1530 114 1553
rect 110 1529 116 1530
rect 160 1529 162 1553
rect 376 1529 378 1553
rect 608 1529 610 1553
rect 840 1529 842 1553
rect 1072 1529 1074 1553
rect 1304 1529 1306 1553
rect 1936 1530 1938 1553
rect 2118 1552 2124 1553
rect 1974 1551 1980 1552
rect 1974 1547 1975 1551
rect 1979 1547 1980 1551
rect 2118 1548 2119 1552
rect 2123 1548 2124 1552
rect 2118 1547 2124 1548
rect 2254 1552 2260 1553
rect 2254 1548 2255 1552
rect 2259 1548 2260 1552
rect 2254 1547 2260 1548
rect 2390 1552 2396 1553
rect 2390 1548 2391 1552
rect 2395 1548 2396 1552
rect 2390 1547 2396 1548
rect 2526 1552 2532 1553
rect 2526 1548 2527 1552
rect 2531 1548 2532 1552
rect 2526 1547 2532 1548
rect 2662 1552 2668 1553
rect 2662 1548 2663 1552
rect 2667 1548 2668 1552
rect 2662 1547 2668 1548
rect 2798 1552 2804 1553
rect 2798 1548 2799 1552
rect 2803 1548 2804 1552
rect 2798 1547 2804 1548
rect 2934 1552 2940 1553
rect 2934 1548 2935 1552
rect 2939 1548 2940 1552
rect 2934 1547 2940 1548
rect 3070 1552 3076 1553
rect 3070 1548 3071 1552
rect 3075 1548 3076 1552
rect 3070 1547 3076 1548
rect 3206 1552 3212 1553
rect 3886 1552 3892 1553
rect 3206 1548 3207 1552
rect 3211 1548 3212 1552
rect 3206 1547 3212 1548
rect 3798 1551 3804 1552
rect 3798 1547 3799 1551
rect 3803 1547 3804 1551
rect 1974 1546 1980 1547
rect 1934 1529 1940 1530
rect 110 1525 111 1529
rect 115 1525 116 1529
rect 110 1524 116 1525
rect 158 1528 164 1529
rect 158 1524 159 1528
rect 163 1524 164 1528
rect 158 1523 164 1524
rect 374 1528 380 1529
rect 374 1524 375 1528
rect 379 1524 380 1528
rect 374 1523 380 1524
rect 606 1528 612 1529
rect 606 1524 607 1528
rect 611 1524 612 1528
rect 606 1523 612 1524
rect 838 1528 844 1529
rect 838 1524 839 1528
rect 843 1524 844 1528
rect 838 1523 844 1524
rect 1070 1528 1076 1529
rect 1070 1524 1071 1528
rect 1075 1524 1076 1528
rect 1070 1523 1076 1524
rect 1302 1528 1308 1529
rect 1302 1524 1303 1528
rect 1307 1524 1308 1528
rect 1934 1525 1935 1529
rect 1939 1525 1940 1529
rect 1934 1524 1940 1525
rect 1302 1523 1308 1524
rect 130 1513 136 1514
rect 110 1512 116 1513
rect 110 1508 111 1512
rect 115 1508 116 1512
rect 130 1509 131 1513
rect 135 1509 136 1513
rect 130 1508 136 1509
rect 346 1513 352 1514
rect 346 1509 347 1513
rect 351 1509 352 1513
rect 346 1508 352 1509
rect 578 1513 584 1514
rect 578 1509 579 1513
rect 583 1509 584 1513
rect 578 1508 584 1509
rect 810 1513 816 1514
rect 810 1509 811 1513
rect 815 1509 816 1513
rect 810 1508 816 1509
rect 1042 1513 1048 1514
rect 1042 1509 1043 1513
rect 1047 1509 1048 1513
rect 1042 1508 1048 1509
rect 1274 1513 1280 1514
rect 1274 1509 1275 1513
rect 1279 1509 1280 1513
rect 1274 1508 1280 1509
rect 1934 1512 1940 1513
rect 1934 1508 1935 1512
rect 1939 1508 1940 1512
rect 110 1507 116 1508
rect 112 1435 114 1507
rect 132 1435 134 1508
rect 348 1435 350 1508
rect 580 1435 582 1508
rect 812 1435 814 1508
rect 1044 1435 1046 1508
rect 1276 1435 1278 1508
rect 1934 1507 1940 1508
rect 1936 1435 1938 1507
rect 1976 1503 1978 1546
rect 2120 1503 2122 1547
rect 2256 1503 2258 1547
rect 2392 1503 2394 1547
rect 2528 1503 2530 1547
rect 2664 1503 2666 1547
rect 2800 1503 2802 1547
rect 2936 1503 2938 1547
rect 3072 1503 3074 1547
rect 3208 1503 3210 1547
rect 3798 1546 3804 1547
rect 3838 1551 3844 1552
rect 3838 1547 3839 1551
rect 3843 1547 3844 1551
rect 3886 1548 3887 1552
rect 3891 1548 3892 1552
rect 3886 1547 3892 1548
rect 4022 1552 4028 1553
rect 4022 1548 4023 1552
rect 4027 1548 4028 1552
rect 4022 1547 4028 1548
rect 4182 1552 4188 1553
rect 4182 1548 4183 1552
rect 4187 1548 4188 1552
rect 4182 1547 4188 1548
rect 4382 1552 4388 1553
rect 4382 1548 4383 1552
rect 4387 1548 4388 1552
rect 4382 1547 4388 1548
rect 4614 1552 4620 1553
rect 4614 1548 4615 1552
rect 4619 1548 4620 1552
rect 4614 1547 4620 1548
rect 4878 1552 4884 1553
rect 4878 1548 4879 1552
rect 4883 1548 4884 1552
rect 4878 1547 4884 1548
rect 5158 1552 5164 1553
rect 5158 1548 5159 1552
rect 5163 1548 5164 1552
rect 5158 1547 5164 1548
rect 5446 1552 5452 1553
rect 5446 1548 5447 1552
rect 5451 1548 5452 1552
rect 5446 1547 5452 1548
rect 5662 1551 5668 1552
rect 5662 1547 5663 1551
rect 5667 1547 5668 1551
rect 3838 1546 3844 1547
rect 3800 1503 3802 1546
rect 3840 1523 3842 1546
rect 3888 1523 3890 1547
rect 4024 1523 4026 1547
rect 4184 1523 4186 1547
rect 4384 1523 4386 1547
rect 4616 1523 4618 1547
rect 4880 1523 4882 1547
rect 5160 1523 5162 1547
rect 5448 1523 5450 1547
rect 5662 1546 5668 1547
rect 5664 1523 5666 1546
rect 3839 1522 3843 1523
rect 3839 1517 3843 1518
rect 3887 1522 3891 1523
rect 3887 1517 3891 1518
rect 4023 1522 4027 1523
rect 4023 1517 4027 1518
rect 4159 1522 4163 1523
rect 4159 1517 4163 1518
rect 4183 1522 4187 1523
rect 4183 1517 4187 1518
rect 4303 1522 4307 1523
rect 4303 1517 4307 1518
rect 4383 1522 4387 1523
rect 4383 1517 4387 1518
rect 4495 1522 4499 1523
rect 4495 1517 4499 1518
rect 4615 1522 4619 1523
rect 4615 1517 4619 1518
rect 4719 1522 4723 1523
rect 4719 1517 4723 1518
rect 4879 1522 4883 1523
rect 4879 1517 4883 1518
rect 4967 1522 4971 1523
rect 4967 1517 4971 1518
rect 5159 1522 5163 1523
rect 5159 1517 5163 1518
rect 5223 1522 5227 1523
rect 5223 1517 5227 1518
rect 5447 1522 5451 1523
rect 5447 1517 5451 1518
rect 5487 1522 5491 1523
rect 5487 1517 5491 1518
rect 5663 1522 5667 1523
rect 5663 1517 5667 1518
rect 1975 1502 1979 1503
rect 1975 1497 1979 1498
rect 2023 1502 2027 1503
rect 2023 1497 2027 1498
rect 2119 1502 2123 1503
rect 2119 1497 2123 1498
rect 2159 1502 2163 1503
rect 2159 1497 2163 1498
rect 2255 1502 2259 1503
rect 2255 1497 2259 1498
rect 2295 1502 2299 1503
rect 2295 1497 2299 1498
rect 2391 1502 2395 1503
rect 2391 1497 2395 1498
rect 2431 1502 2435 1503
rect 2431 1497 2435 1498
rect 2527 1502 2531 1503
rect 2527 1497 2531 1498
rect 2567 1502 2571 1503
rect 2567 1497 2571 1498
rect 2663 1502 2667 1503
rect 2663 1497 2667 1498
rect 2703 1502 2707 1503
rect 2703 1497 2707 1498
rect 2799 1502 2803 1503
rect 2799 1497 2803 1498
rect 2839 1502 2843 1503
rect 2839 1497 2843 1498
rect 2935 1502 2939 1503
rect 2935 1497 2939 1498
rect 2975 1502 2979 1503
rect 2975 1497 2979 1498
rect 3071 1502 3075 1503
rect 3071 1497 3075 1498
rect 3207 1502 3211 1503
rect 3207 1497 3211 1498
rect 3799 1502 3803 1503
rect 3799 1497 3803 1498
rect 1976 1474 1978 1497
rect 1974 1473 1980 1474
rect 2024 1473 2026 1497
rect 2160 1473 2162 1497
rect 2296 1473 2298 1497
rect 2432 1473 2434 1497
rect 2568 1473 2570 1497
rect 2704 1473 2706 1497
rect 2840 1473 2842 1497
rect 2976 1473 2978 1497
rect 3800 1474 3802 1497
rect 3840 1494 3842 1517
rect 3838 1493 3844 1494
rect 3888 1493 3890 1517
rect 4024 1493 4026 1517
rect 4160 1493 4162 1517
rect 4304 1493 4306 1517
rect 4496 1493 4498 1517
rect 4720 1493 4722 1517
rect 4968 1493 4970 1517
rect 5224 1493 5226 1517
rect 5488 1493 5490 1517
rect 5664 1494 5666 1517
rect 5662 1493 5668 1494
rect 3838 1489 3839 1493
rect 3843 1489 3844 1493
rect 3838 1488 3844 1489
rect 3886 1492 3892 1493
rect 3886 1488 3887 1492
rect 3891 1488 3892 1492
rect 3886 1487 3892 1488
rect 4022 1492 4028 1493
rect 4022 1488 4023 1492
rect 4027 1488 4028 1492
rect 4022 1487 4028 1488
rect 4158 1492 4164 1493
rect 4158 1488 4159 1492
rect 4163 1488 4164 1492
rect 4158 1487 4164 1488
rect 4302 1492 4308 1493
rect 4302 1488 4303 1492
rect 4307 1488 4308 1492
rect 4302 1487 4308 1488
rect 4494 1492 4500 1493
rect 4494 1488 4495 1492
rect 4499 1488 4500 1492
rect 4494 1487 4500 1488
rect 4718 1492 4724 1493
rect 4718 1488 4719 1492
rect 4723 1488 4724 1492
rect 4718 1487 4724 1488
rect 4966 1492 4972 1493
rect 4966 1488 4967 1492
rect 4971 1488 4972 1492
rect 4966 1487 4972 1488
rect 5222 1492 5228 1493
rect 5222 1488 5223 1492
rect 5227 1488 5228 1492
rect 5222 1487 5228 1488
rect 5486 1492 5492 1493
rect 5486 1488 5487 1492
rect 5491 1488 5492 1492
rect 5662 1489 5663 1493
rect 5667 1489 5668 1493
rect 5662 1488 5668 1489
rect 5486 1487 5492 1488
rect 3858 1477 3864 1478
rect 3838 1476 3844 1477
rect 3798 1473 3804 1474
rect 1974 1469 1975 1473
rect 1979 1469 1980 1473
rect 1974 1468 1980 1469
rect 2022 1472 2028 1473
rect 2022 1468 2023 1472
rect 2027 1468 2028 1472
rect 2022 1467 2028 1468
rect 2158 1472 2164 1473
rect 2158 1468 2159 1472
rect 2163 1468 2164 1472
rect 2158 1467 2164 1468
rect 2294 1472 2300 1473
rect 2294 1468 2295 1472
rect 2299 1468 2300 1472
rect 2294 1467 2300 1468
rect 2430 1472 2436 1473
rect 2430 1468 2431 1472
rect 2435 1468 2436 1472
rect 2430 1467 2436 1468
rect 2566 1472 2572 1473
rect 2566 1468 2567 1472
rect 2571 1468 2572 1472
rect 2566 1467 2572 1468
rect 2702 1472 2708 1473
rect 2702 1468 2703 1472
rect 2707 1468 2708 1472
rect 2702 1467 2708 1468
rect 2838 1472 2844 1473
rect 2838 1468 2839 1472
rect 2843 1468 2844 1472
rect 2838 1467 2844 1468
rect 2974 1472 2980 1473
rect 2974 1468 2975 1472
rect 2979 1468 2980 1472
rect 3798 1469 3799 1473
rect 3803 1469 3804 1473
rect 3838 1472 3839 1476
rect 3843 1472 3844 1476
rect 3858 1473 3859 1477
rect 3863 1473 3864 1477
rect 3858 1472 3864 1473
rect 3994 1477 4000 1478
rect 3994 1473 3995 1477
rect 3999 1473 4000 1477
rect 3994 1472 4000 1473
rect 4130 1477 4136 1478
rect 4130 1473 4131 1477
rect 4135 1473 4136 1477
rect 4130 1472 4136 1473
rect 4274 1477 4280 1478
rect 4274 1473 4275 1477
rect 4279 1473 4280 1477
rect 4274 1472 4280 1473
rect 4466 1477 4472 1478
rect 4466 1473 4467 1477
rect 4471 1473 4472 1477
rect 4466 1472 4472 1473
rect 4690 1477 4696 1478
rect 4690 1473 4691 1477
rect 4695 1473 4696 1477
rect 4690 1472 4696 1473
rect 4938 1477 4944 1478
rect 4938 1473 4939 1477
rect 4943 1473 4944 1477
rect 4938 1472 4944 1473
rect 5194 1477 5200 1478
rect 5194 1473 5195 1477
rect 5199 1473 5200 1477
rect 5194 1472 5200 1473
rect 5458 1477 5464 1478
rect 5458 1473 5459 1477
rect 5463 1473 5464 1477
rect 5458 1472 5464 1473
rect 5662 1476 5668 1477
rect 5662 1472 5663 1476
rect 5667 1472 5668 1476
rect 3838 1471 3844 1472
rect 3798 1468 3804 1469
rect 2974 1467 2980 1468
rect 1994 1457 2000 1458
rect 1974 1456 1980 1457
rect 1974 1452 1975 1456
rect 1979 1452 1980 1456
rect 1994 1453 1995 1457
rect 1999 1453 2000 1457
rect 1994 1452 2000 1453
rect 2130 1457 2136 1458
rect 2130 1453 2131 1457
rect 2135 1453 2136 1457
rect 2130 1452 2136 1453
rect 2266 1457 2272 1458
rect 2266 1453 2267 1457
rect 2271 1453 2272 1457
rect 2266 1452 2272 1453
rect 2402 1457 2408 1458
rect 2402 1453 2403 1457
rect 2407 1453 2408 1457
rect 2402 1452 2408 1453
rect 2538 1457 2544 1458
rect 2538 1453 2539 1457
rect 2543 1453 2544 1457
rect 2538 1452 2544 1453
rect 2674 1457 2680 1458
rect 2674 1453 2675 1457
rect 2679 1453 2680 1457
rect 2674 1452 2680 1453
rect 2810 1457 2816 1458
rect 2810 1453 2811 1457
rect 2815 1453 2816 1457
rect 2810 1452 2816 1453
rect 2946 1457 2952 1458
rect 2946 1453 2947 1457
rect 2951 1453 2952 1457
rect 2946 1452 2952 1453
rect 3798 1456 3804 1457
rect 3798 1452 3799 1456
rect 3803 1452 3804 1456
rect 1974 1451 1980 1452
rect 111 1434 115 1435
rect 111 1429 115 1430
rect 131 1434 135 1435
rect 131 1429 135 1430
rect 347 1434 351 1435
rect 347 1429 351 1430
rect 411 1434 415 1435
rect 411 1429 415 1430
rect 579 1434 583 1435
rect 579 1429 583 1430
rect 739 1434 743 1435
rect 739 1429 743 1430
rect 811 1434 815 1435
rect 811 1429 815 1430
rect 1043 1434 1047 1435
rect 1043 1429 1047 1430
rect 1091 1434 1095 1435
rect 1091 1429 1095 1430
rect 1275 1434 1279 1435
rect 1275 1429 1279 1430
rect 1451 1434 1455 1435
rect 1451 1429 1455 1430
rect 1787 1434 1791 1435
rect 1787 1429 1791 1430
rect 1935 1434 1939 1435
rect 1935 1429 1939 1430
rect 112 1369 114 1429
rect 110 1368 116 1369
rect 132 1368 134 1429
rect 412 1368 414 1429
rect 740 1368 742 1429
rect 1092 1368 1094 1429
rect 1452 1368 1454 1429
rect 1788 1368 1790 1429
rect 1936 1369 1938 1429
rect 1976 1383 1978 1451
rect 1996 1383 1998 1452
rect 2132 1383 2134 1452
rect 2268 1383 2270 1452
rect 2404 1383 2406 1452
rect 2540 1383 2542 1452
rect 2676 1383 2678 1452
rect 2812 1383 2814 1452
rect 2948 1383 2950 1452
rect 3798 1451 3804 1452
rect 3800 1383 3802 1451
rect 3840 1407 3842 1471
rect 3860 1407 3862 1472
rect 3996 1407 3998 1472
rect 4132 1407 4134 1472
rect 4276 1407 4278 1472
rect 4468 1407 4470 1472
rect 4692 1407 4694 1472
rect 4940 1407 4942 1472
rect 5196 1407 5198 1472
rect 5460 1407 5462 1472
rect 5662 1471 5668 1472
rect 5664 1407 5666 1471
rect 3839 1406 3843 1407
rect 3839 1401 3843 1402
rect 3859 1406 3863 1407
rect 3859 1401 3863 1402
rect 3995 1406 3999 1407
rect 3995 1401 3999 1402
rect 4059 1406 4063 1407
rect 4059 1401 4063 1402
rect 4131 1406 4135 1407
rect 4131 1401 4135 1402
rect 4275 1406 4279 1407
rect 4275 1401 4279 1402
rect 4307 1406 4311 1407
rect 4307 1401 4311 1402
rect 4467 1406 4471 1407
rect 4467 1401 4471 1402
rect 4579 1406 4583 1407
rect 4579 1401 4583 1402
rect 4691 1406 4695 1407
rect 4691 1401 4695 1402
rect 4875 1406 4879 1407
rect 4875 1401 4879 1402
rect 4939 1406 4943 1407
rect 4939 1401 4943 1402
rect 5187 1406 5191 1407
rect 5187 1401 5191 1402
rect 5195 1406 5199 1407
rect 5195 1401 5199 1402
rect 5459 1406 5463 1407
rect 5459 1401 5463 1402
rect 5499 1406 5503 1407
rect 5499 1401 5503 1402
rect 5663 1406 5667 1407
rect 5663 1401 5667 1402
rect 1975 1382 1979 1383
rect 1975 1377 1979 1378
rect 1995 1382 1999 1383
rect 1995 1377 1999 1378
rect 2131 1382 2135 1383
rect 2131 1377 2135 1378
rect 2267 1382 2271 1383
rect 2267 1377 2271 1378
rect 2275 1382 2279 1383
rect 2275 1377 2279 1378
rect 2403 1382 2407 1383
rect 2403 1377 2407 1378
rect 2539 1382 2543 1383
rect 2539 1377 2543 1378
rect 2563 1382 2567 1383
rect 2563 1377 2567 1378
rect 2675 1382 2679 1383
rect 2675 1377 2679 1378
rect 2811 1382 2815 1383
rect 2811 1377 2815 1378
rect 2843 1382 2847 1383
rect 2843 1377 2847 1378
rect 2947 1382 2951 1383
rect 2947 1377 2951 1378
rect 3123 1382 3127 1383
rect 3123 1377 3127 1378
rect 3395 1382 3399 1383
rect 3395 1377 3399 1378
rect 3651 1382 3655 1383
rect 3651 1377 3655 1378
rect 3799 1382 3803 1383
rect 3799 1377 3803 1378
rect 1934 1368 1940 1369
rect 110 1364 111 1368
rect 115 1364 116 1368
rect 110 1363 116 1364
rect 130 1367 136 1368
rect 130 1363 131 1367
rect 135 1363 136 1367
rect 130 1362 136 1363
rect 410 1367 416 1368
rect 410 1363 411 1367
rect 415 1363 416 1367
rect 410 1362 416 1363
rect 738 1367 744 1368
rect 738 1363 739 1367
rect 743 1363 744 1367
rect 738 1362 744 1363
rect 1090 1367 1096 1368
rect 1090 1363 1091 1367
rect 1095 1363 1096 1367
rect 1090 1362 1096 1363
rect 1450 1367 1456 1368
rect 1450 1363 1451 1367
rect 1455 1363 1456 1367
rect 1450 1362 1456 1363
rect 1786 1367 1792 1368
rect 1786 1363 1787 1367
rect 1791 1363 1792 1367
rect 1934 1364 1935 1368
rect 1939 1364 1940 1368
rect 1934 1363 1940 1364
rect 1786 1362 1792 1363
rect 158 1352 164 1353
rect 110 1351 116 1352
rect 110 1347 111 1351
rect 115 1347 116 1351
rect 158 1348 159 1352
rect 163 1348 164 1352
rect 158 1347 164 1348
rect 438 1352 444 1353
rect 438 1348 439 1352
rect 443 1348 444 1352
rect 438 1347 444 1348
rect 766 1352 772 1353
rect 766 1348 767 1352
rect 771 1348 772 1352
rect 766 1347 772 1348
rect 1118 1352 1124 1353
rect 1118 1348 1119 1352
rect 1123 1348 1124 1352
rect 1118 1347 1124 1348
rect 1478 1352 1484 1353
rect 1478 1348 1479 1352
rect 1483 1348 1484 1352
rect 1478 1347 1484 1348
rect 1814 1352 1820 1353
rect 1814 1348 1815 1352
rect 1819 1348 1820 1352
rect 1814 1347 1820 1348
rect 1934 1351 1940 1352
rect 1934 1347 1935 1351
rect 1939 1347 1940 1351
rect 110 1346 116 1347
rect 112 1323 114 1346
rect 160 1323 162 1347
rect 440 1323 442 1347
rect 768 1323 770 1347
rect 1120 1323 1122 1347
rect 1480 1323 1482 1347
rect 1816 1323 1818 1347
rect 1934 1346 1940 1347
rect 1936 1323 1938 1346
rect 111 1322 115 1323
rect 111 1317 115 1318
rect 159 1322 163 1323
rect 159 1317 163 1318
rect 359 1322 363 1323
rect 359 1317 363 1318
rect 439 1322 443 1323
rect 439 1317 443 1318
rect 575 1322 579 1323
rect 575 1317 579 1318
rect 767 1322 771 1323
rect 767 1317 771 1318
rect 775 1322 779 1323
rect 775 1317 779 1318
rect 967 1322 971 1323
rect 967 1317 971 1318
rect 1119 1322 1123 1323
rect 1119 1317 1123 1318
rect 1151 1322 1155 1323
rect 1151 1317 1155 1318
rect 1327 1322 1331 1323
rect 1327 1317 1331 1318
rect 1479 1322 1483 1323
rect 1479 1317 1483 1318
rect 1495 1322 1499 1323
rect 1495 1317 1499 1318
rect 1663 1322 1667 1323
rect 1663 1317 1667 1318
rect 1815 1322 1819 1323
rect 1815 1317 1819 1318
rect 1935 1322 1939 1323
rect 1935 1317 1939 1318
rect 1976 1317 1978 1377
rect 112 1294 114 1317
rect 110 1293 116 1294
rect 160 1293 162 1317
rect 360 1293 362 1317
rect 576 1293 578 1317
rect 776 1293 778 1317
rect 968 1293 970 1317
rect 1152 1293 1154 1317
rect 1328 1293 1330 1317
rect 1496 1293 1498 1317
rect 1664 1293 1666 1317
rect 1816 1293 1818 1317
rect 1936 1294 1938 1317
rect 1974 1316 1980 1317
rect 1996 1316 1998 1377
rect 2276 1316 2278 1377
rect 2564 1316 2566 1377
rect 2844 1316 2846 1377
rect 3124 1316 3126 1377
rect 3396 1316 3398 1377
rect 3652 1316 3654 1377
rect 3800 1317 3802 1377
rect 3840 1341 3842 1401
rect 3838 1340 3844 1341
rect 3860 1340 3862 1401
rect 4060 1340 4062 1401
rect 4308 1340 4310 1401
rect 4580 1340 4582 1401
rect 4876 1340 4878 1401
rect 5188 1340 5190 1401
rect 5500 1340 5502 1401
rect 5664 1341 5666 1401
rect 5662 1340 5668 1341
rect 3838 1336 3839 1340
rect 3843 1336 3844 1340
rect 3838 1335 3844 1336
rect 3858 1339 3864 1340
rect 3858 1335 3859 1339
rect 3863 1335 3864 1339
rect 3858 1334 3864 1335
rect 4058 1339 4064 1340
rect 4058 1335 4059 1339
rect 4063 1335 4064 1339
rect 4058 1334 4064 1335
rect 4306 1339 4312 1340
rect 4306 1335 4307 1339
rect 4311 1335 4312 1339
rect 4306 1334 4312 1335
rect 4578 1339 4584 1340
rect 4578 1335 4579 1339
rect 4583 1335 4584 1339
rect 4578 1334 4584 1335
rect 4874 1339 4880 1340
rect 4874 1335 4875 1339
rect 4879 1335 4880 1339
rect 4874 1334 4880 1335
rect 5186 1339 5192 1340
rect 5186 1335 5187 1339
rect 5191 1335 5192 1339
rect 5186 1334 5192 1335
rect 5498 1339 5504 1340
rect 5498 1335 5499 1339
rect 5503 1335 5504 1339
rect 5662 1336 5663 1340
rect 5667 1336 5668 1340
rect 5662 1335 5668 1336
rect 5498 1334 5504 1335
rect 3886 1324 3892 1325
rect 3838 1323 3844 1324
rect 3838 1319 3839 1323
rect 3843 1319 3844 1323
rect 3886 1320 3887 1324
rect 3891 1320 3892 1324
rect 3886 1319 3892 1320
rect 4086 1324 4092 1325
rect 4086 1320 4087 1324
rect 4091 1320 4092 1324
rect 4086 1319 4092 1320
rect 4334 1324 4340 1325
rect 4334 1320 4335 1324
rect 4339 1320 4340 1324
rect 4334 1319 4340 1320
rect 4606 1324 4612 1325
rect 4606 1320 4607 1324
rect 4611 1320 4612 1324
rect 4606 1319 4612 1320
rect 4902 1324 4908 1325
rect 4902 1320 4903 1324
rect 4907 1320 4908 1324
rect 4902 1319 4908 1320
rect 5214 1324 5220 1325
rect 5214 1320 5215 1324
rect 5219 1320 5220 1324
rect 5214 1319 5220 1320
rect 5526 1324 5532 1325
rect 5526 1320 5527 1324
rect 5531 1320 5532 1324
rect 5526 1319 5532 1320
rect 5662 1323 5668 1324
rect 5662 1319 5663 1323
rect 5667 1319 5668 1323
rect 3838 1318 3844 1319
rect 3798 1316 3804 1317
rect 1974 1312 1975 1316
rect 1979 1312 1980 1316
rect 1974 1311 1980 1312
rect 1994 1315 2000 1316
rect 1994 1311 1995 1315
rect 1999 1311 2000 1315
rect 1994 1310 2000 1311
rect 2274 1315 2280 1316
rect 2274 1311 2275 1315
rect 2279 1311 2280 1315
rect 2274 1310 2280 1311
rect 2562 1315 2568 1316
rect 2562 1311 2563 1315
rect 2567 1311 2568 1315
rect 2562 1310 2568 1311
rect 2842 1315 2848 1316
rect 2842 1311 2843 1315
rect 2847 1311 2848 1315
rect 2842 1310 2848 1311
rect 3122 1315 3128 1316
rect 3122 1311 3123 1315
rect 3127 1311 3128 1315
rect 3122 1310 3128 1311
rect 3394 1315 3400 1316
rect 3394 1311 3395 1315
rect 3399 1311 3400 1315
rect 3394 1310 3400 1311
rect 3650 1315 3656 1316
rect 3650 1311 3651 1315
rect 3655 1311 3656 1315
rect 3798 1312 3799 1316
rect 3803 1312 3804 1316
rect 3798 1311 3804 1312
rect 3650 1310 3656 1311
rect 2022 1300 2028 1301
rect 1974 1299 1980 1300
rect 1974 1295 1975 1299
rect 1979 1295 1980 1299
rect 2022 1296 2023 1300
rect 2027 1296 2028 1300
rect 2022 1295 2028 1296
rect 2302 1300 2308 1301
rect 2302 1296 2303 1300
rect 2307 1296 2308 1300
rect 2302 1295 2308 1296
rect 2590 1300 2596 1301
rect 2590 1296 2591 1300
rect 2595 1296 2596 1300
rect 2590 1295 2596 1296
rect 2870 1300 2876 1301
rect 2870 1296 2871 1300
rect 2875 1296 2876 1300
rect 2870 1295 2876 1296
rect 3150 1300 3156 1301
rect 3150 1296 3151 1300
rect 3155 1296 3156 1300
rect 3150 1295 3156 1296
rect 3422 1300 3428 1301
rect 3422 1296 3423 1300
rect 3427 1296 3428 1300
rect 3422 1295 3428 1296
rect 3678 1300 3684 1301
rect 3678 1296 3679 1300
rect 3683 1296 3684 1300
rect 3678 1295 3684 1296
rect 3798 1299 3804 1300
rect 3798 1295 3799 1299
rect 3803 1295 3804 1299
rect 1974 1294 1980 1295
rect 1934 1293 1940 1294
rect 110 1289 111 1293
rect 115 1289 116 1293
rect 110 1288 116 1289
rect 158 1292 164 1293
rect 158 1288 159 1292
rect 163 1288 164 1292
rect 158 1287 164 1288
rect 358 1292 364 1293
rect 358 1288 359 1292
rect 363 1288 364 1292
rect 358 1287 364 1288
rect 574 1292 580 1293
rect 574 1288 575 1292
rect 579 1288 580 1292
rect 574 1287 580 1288
rect 774 1292 780 1293
rect 774 1288 775 1292
rect 779 1288 780 1292
rect 774 1287 780 1288
rect 966 1292 972 1293
rect 966 1288 967 1292
rect 971 1288 972 1292
rect 966 1287 972 1288
rect 1150 1292 1156 1293
rect 1150 1288 1151 1292
rect 1155 1288 1156 1292
rect 1150 1287 1156 1288
rect 1326 1292 1332 1293
rect 1326 1288 1327 1292
rect 1331 1288 1332 1292
rect 1326 1287 1332 1288
rect 1494 1292 1500 1293
rect 1494 1288 1495 1292
rect 1499 1288 1500 1292
rect 1494 1287 1500 1288
rect 1662 1292 1668 1293
rect 1662 1288 1663 1292
rect 1667 1288 1668 1292
rect 1662 1287 1668 1288
rect 1814 1292 1820 1293
rect 1814 1288 1815 1292
rect 1819 1288 1820 1292
rect 1934 1289 1935 1293
rect 1939 1289 1940 1293
rect 1934 1288 1940 1289
rect 1814 1287 1820 1288
rect 130 1277 136 1278
rect 110 1276 116 1277
rect 110 1272 111 1276
rect 115 1272 116 1276
rect 130 1273 131 1277
rect 135 1273 136 1277
rect 130 1272 136 1273
rect 330 1277 336 1278
rect 330 1273 331 1277
rect 335 1273 336 1277
rect 330 1272 336 1273
rect 546 1277 552 1278
rect 546 1273 547 1277
rect 551 1273 552 1277
rect 546 1272 552 1273
rect 746 1277 752 1278
rect 746 1273 747 1277
rect 751 1273 752 1277
rect 746 1272 752 1273
rect 938 1277 944 1278
rect 938 1273 939 1277
rect 943 1273 944 1277
rect 938 1272 944 1273
rect 1122 1277 1128 1278
rect 1122 1273 1123 1277
rect 1127 1273 1128 1277
rect 1122 1272 1128 1273
rect 1298 1277 1304 1278
rect 1298 1273 1299 1277
rect 1303 1273 1304 1277
rect 1298 1272 1304 1273
rect 1466 1277 1472 1278
rect 1466 1273 1467 1277
rect 1471 1273 1472 1277
rect 1466 1272 1472 1273
rect 1634 1277 1640 1278
rect 1634 1273 1635 1277
rect 1639 1273 1640 1277
rect 1634 1272 1640 1273
rect 1786 1277 1792 1278
rect 1786 1273 1787 1277
rect 1791 1273 1792 1277
rect 1786 1272 1792 1273
rect 1934 1276 1940 1277
rect 1934 1272 1935 1276
rect 1939 1272 1940 1276
rect 110 1271 116 1272
rect 112 1199 114 1271
rect 132 1199 134 1272
rect 332 1199 334 1272
rect 548 1199 550 1272
rect 748 1199 750 1272
rect 940 1199 942 1272
rect 1124 1199 1126 1272
rect 1300 1199 1302 1272
rect 1468 1199 1470 1272
rect 1636 1199 1638 1272
rect 1788 1199 1790 1272
rect 1934 1271 1940 1272
rect 1936 1199 1938 1271
rect 1976 1247 1978 1294
rect 2024 1247 2026 1295
rect 2304 1247 2306 1295
rect 2592 1247 2594 1295
rect 2872 1247 2874 1295
rect 3152 1247 3154 1295
rect 3424 1247 3426 1295
rect 3680 1247 3682 1295
rect 3798 1294 3804 1295
rect 3800 1247 3802 1294
rect 3840 1287 3842 1318
rect 3888 1287 3890 1319
rect 4088 1287 4090 1319
rect 4336 1287 4338 1319
rect 4608 1287 4610 1319
rect 4904 1287 4906 1319
rect 5216 1287 5218 1319
rect 5528 1287 5530 1319
rect 5662 1318 5668 1319
rect 5664 1287 5666 1318
rect 3839 1286 3843 1287
rect 3839 1281 3843 1282
rect 3887 1286 3891 1287
rect 3887 1281 3891 1282
rect 4087 1286 4091 1287
rect 4087 1281 4091 1282
rect 4335 1286 4339 1287
rect 4335 1281 4339 1282
rect 4607 1286 4611 1287
rect 4607 1281 4611 1282
rect 4615 1286 4619 1287
rect 4615 1281 4619 1282
rect 4791 1286 4795 1287
rect 4791 1281 4795 1282
rect 4903 1286 4907 1287
rect 4903 1281 4907 1282
rect 4975 1286 4979 1287
rect 4975 1281 4979 1282
rect 5167 1286 5171 1287
rect 5167 1281 5171 1282
rect 5215 1286 5219 1287
rect 5215 1281 5219 1282
rect 5367 1286 5371 1287
rect 5367 1281 5371 1282
rect 5527 1286 5531 1287
rect 5527 1281 5531 1282
rect 5543 1286 5547 1287
rect 5543 1281 5547 1282
rect 5663 1286 5667 1287
rect 5663 1281 5667 1282
rect 3840 1258 3842 1281
rect 3838 1257 3844 1258
rect 4616 1257 4618 1281
rect 4792 1257 4794 1281
rect 4976 1257 4978 1281
rect 5168 1257 5170 1281
rect 5368 1257 5370 1281
rect 5544 1257 5546 1281
rect 5664 1258 5666 1281
rect 5662 1257 5668 1258
rect 3838 1253 3839 1257
rect 3843 1253 3844 1257
rect 3838 1252 3844 1253
rect 4614 1256 4620 1257
rect 4614 1252 4615 1256
rect 4619 1252 4620 1256
rect 4614 1251 4620 1252
rect 4790 1256 4796 1257
rect 4790 1252 4791 1256
rect 4795 1252 4796 1256
rect 4790 1251 4796 1252
rect 4974 1256 4980 1257
rect 4974 1252 4975 1256
rect 4979 1252 4980 1256
rect 4974 1251 4980 1252
rect 5166 1256 5172 1257
rect 5166 1252 5167 1256
rect 5171 1252 5172 1256
rect 5166 1251 5172 1252
rect 5366 1256 5372 1257
rect 5366 1252 5367 1256
rect 5371 1252 5372 1256
rect 5366 1251 5372 1252
rect 5542 1256 5548 1257
rect 5542 1252 5543 1256
rect 5547 1252 5548 1256
rect 5662 1253 5663 1257
rect 5667 1253 5668 1257
rect 5662 1252 5668 1253
rect 5542 1251 5548 1252
rect 1975 1246 1979 1247
rect 1975 1241 1979 1242
rect 2023 1246 2027 1247
rect 2023 1241 2027 1242
rect 2303 1246 2307 1247
rect 2303 1241 2307 1242
rect 2591 1246 2595 1247
rect 2591 1241 2595 1242
rect 2655 1246 2659 1247
rect 2655 1241 2659 1242
rect 2831 1246 2835 1247
rect 2831 1241 2835 1242
rect 2871 1246 2875 1247
rect 2871 1241 2875 1242
rect 3007 1246 3011 1247
rect 3007 1241 3011 1242
rect 3151 1246 3155 1247
rect 3151 1241 3155 1242
rect 3183 1246 3187 1247
rect 3183 1241 3187 1242
rect 3359 1246 3363 1247
rect 3359 1241 3363 1242
rect 3423 1246 3427 1247
rect 3423 1241 3427 1242
rect 3543 1246 3547 1247
rect 3543 1241 3547 1242
rect 3679 1246 3683 1247
rect 3679 1241 3683 1242
rect 3799 1246 3803 1247
rect 3799 1241 3803 1242
rect 4586 1241 4592 1242
rect 1976 1218 1978 1241
rect 1974 1217 1980 1218
rect 2656 1217 2658 1241
rect 2832 1217 2834 1241
rect 3008 1217 3010 1241
rect 3184 1217 3186 1241
rect 3360 1217 3362 1241
rect 3544 1217 3546 1241
rect 3800 1218 3802 1241
rect 3838 1240 3844 1241
rect 3838 1236 3839 1240
rect 3843 1236 3844 1240
rect 4586 1237 4587 1241
rect 4591 1237 4592 1241
rect 4586 1236 4592 1237
rect 4762 1241 4768 1242
rect 4762 1237 4763 1241
rect 4767 1237 4768 1241
rect 4762 1236 4768 1237
rect 4946 1241 4952 1242
rect 4946 1237 4947 1241
rect 4951 1237 4952 1241
rect 4946 1236 4952 1237
rect 5138 1241 5144 1242
rect 5138 1237 5139 1241
rect 5143 1237 5144 1241
rect 5138 1236 5144 1237
rect 5338 1241 5344 1242
rect 5338 1237 5339 1241
rect 5343 1237 5344 1241
rect 5338 1236 5344 1237
rect 5514 1241 5520 1242
rect 5514 1237 5515 1241
rect 5519 1237 5520 1241
rect 5514 1236 5520 1237
rect 5662 1240 5668 1241
rect 5662 1236 5663 1240
rect 5667 1236 5668 1240
rect 3838 1235 3844 1236
rect 3798 1217 3804 1218
rect 1974 1213 1975 1217
rect 1979 1213 1980 1217
rect 1974 1212 1980 1213
rect 2654 1216 2660 1217
rect 2654 1212 2655 1216
rect 2659 1212 2660 1216
rect 2654 1211 2660 1212
rect 2830 1216 2836 1217
rect 2830 1212 2831 1216
rect 2835 1212 2836 1216
rect 2830 1211 2836 1212
rect 3006 1216 3012 1217
rect 3006 1212 3007 1216
rect 3011 1212 3012 1216
rect 3006 1211 3012 1212
rect 3182 1216 3188 1217
rect 3182 1212 3183 1216
rect 3187 1212 3188 1216
rect 3182 1211 3188 1212
rect 3358 1216 3364 1217
rect 3358 1212 3359 1216
rect 3363 1212 3364 1216
rect 3358 1211 3364 1212
rect 3542 1216 3548 1217
rect 3542 1212 3543 1216
rect 3547 1212 3548 1216
rect 3798 1213 3799 1217
rect 3803 1213 3804 1217
rect 3798 1212 3804 1213
rect 3542 1211 3548 1212
rect 2626 1201 2632 1202
rect 1974 1200 1980 1201
rect 111 1198 115 1199
rect 111 1193 115 1194
rect 131 1198 135 1199
rect 131 1193 135 1194
rect 291 1198 295 1199
rect 291 1193 295 1194
rect 331 1198 335 1199
rect 331 1193 335 1194
rect 475 1198 479 1199
rect 475 1193 479 1194
rect 547 1198 551 1199
rect 547 1193 551 1194
rect 659 1198 663 1199
rect 659 1193 663 1194
rect 747 1198 751 1199
rect 747 1193 751 1194
rect 835 1198 839 1199
rect 835 1193 839 1194
rect 939 1198 943 1199
rect 939 1193 943 1194
rect 1003 1198 1007 1199
rect 1003 1193 1007 1194
rect 1123 1198 1127 1199
rect 1123 1193 1127 1194
rect 1171 1198 1175 1199
rect 1171 1193 1175 1194
rect 1299 1198 1303 1199
rect 1299 1193 1303 1194
rect 1331 1198 1335 1199
rect 1331 1193 1335 1194
rect 1467 1198 1471 1199
rect 1467 1193 1471 1194
rect 1491 1198 1495 1199
rect 1491 1193 1495 1194
rect 1635 1198 1639 1199
rect 1635 1193 1639 1194
rect 1651 1198 1655 1199
rect 1651 1193 1655 1194
rect 1787 1198 1791 1199
rect 1787 1193 1791 1194
rect 1935 1198 1939 1199
rect 1974 1196 1975 1200
rect 1979 1196 1980 1200
rect 2626 1197 2627 1201
rect 2631 1197 2632 1201
rect 2626 1196 2632 1197
rect 2802 1201 2808 1202
rect 2802 1197 2803 1201
rect 2807 1197 2808 1201
rect 2802 1196 2808 1197
rect 2978 1201 2984 1202
rect 2978 1197 2979 1201
rect 2983 1197 2984 1201
rect 2978 1196 2984 1197
rect 3154 1201 3160 1202
rect 3154 1197 3155 1201
rect 3159 1197 3160 1201
rect 3154 1196 3160 1197
rect 3330 1201 3336 1202
rect 3330 1197 3331 1201
rect 3335 1197 3336 1201
rect 3330 1196 3336 1197
rect 3514 1201 3520 1202
rect 3514 1197 3515 1201
rect 3519 1197 3520 1201
rect 3514 1196 3520 1197
rect 3798 1200 3804 1201
rect 3798 1196 3799 1200
rect 3803 1196 3804 1200
rect 1974 1195 1980 1196
rect 1935 1193 1939 1194
rect 112 1133 114 1193
rect 110 1132 116 1133
rect 132 1132 134 1193
rect 292 1132 294 1193
rect 476 1132 478 1193
rect 660 1132 662 1193
rect 836 1132 838 1193
rect 1004 1132 1006 1193
rect 1172 1132 1174 1193
rect 1332 1132 1334 1193
rect 1492 1132 1494 1193
rect 1652 1132 1654 1193
rect 1788 1132 1790 1193
rect 1936 1133 1938 1193
rect 1934 1132 1940 1133
rect 110 1128 111 1132
rect 115 1128 116 1132
rect 110 1127 116 1128
rect 130 1131 136 1132
rect 130 1127 131 1131
rect 135 1127 136 1131
rect 130 1126 136 1127
rect 290 1131 296 1132
rect 290 1127 291 1131
rect 295 1127 296 1131
rect 290 1126 296 1127
rect 474 1131 480 1132
rect 474 1127 475 1131
rect 479 1127 480 1131
rect 474 1126 480 1127
rect 658 1131 664 1132
rect 658 1127 659 1131
rect 663 1127 664 1131
rect 658 1126 664 1127
rect 834 1131 840 1132
rect 834 1127 835 1131
rect 839 1127 840 1131
rect 834 1126 840 1127
rect 1002 1131 1008 1132
rect 1002 1127 1003 1131
rect 1007 1127 1008 1131
rect 1002 1126 1008 1127
rect 1170 1131 1176 1132
rect 1170 1127 1171 1131
rect 1175 1127 1176 1131
rect 1170 1126 1176 1127
rect 1330 1131 1336 1132
rect 1330 1127 1331 1131
rect 1335 1127 1336 1131
rect 1330 1126 1336 1127
rect 1490 1131 1496 1132
rect 1490 1127 1491 1131
rect 1495 1127 1496 1131
rect 1490 1126 1496 1127
rect 1650 1131 1656 1132
rect 1650 1127 1651 1131
rect 1655 1127 1656 1131
rect 1650 1126 1656 1127
rect 1786 1131 1792 1132
rect 1786 1127 1787 1131
rect 1791 1127 1792 1131
rect 1934 1128 1935 1132
rect 1939 1128 1940 1132
rect 1934 1127 1940 1128
rect 1786 1126 1792 1127
rect 1976 1119 1978 1195
rect 2628 1119 2630 1196
rect 2804 1119 2806 1196
rect 2980 1119 2982 1196
rect 3156 1119 3158 1196
rect 3332 1119 3334 1196
rect 3516 1119 3518 1196
rect 3798 1195 3804 1196
rect 3800 1119 3802 1195
rect 3840 1171 3842 1235
rect 4588 1171 4590 1236
rect 4764 1171 4766 1236
rect 4948 1171 4950 1236
rect 5140 1171 5142 1236
rect 5340 1171 5342 1236
rect 5516 1171 5518 1236
rect 5662 1235 5668 1236
rect 5664 1171 5666 1235
rect 3839 1170 3843 1171
rect 3839 1165 3843 1166
rect 4587 1170 4591 1171
rect 4587 1165 4591 1166
rect 4763 1170 4767 1171
rect 4763 1165 4767 1166
rect 4835 1170 4839 1171
rect 4835 1165 4839 1166
rect 4947 1170 4951 1171
rect 4947 1165 4951 1166
rect 4971 1170 4975 1171
rect 4971 1165 4975 1166
rect 5107 1170 5111 1171
rect 5107 1165 5111 1166
rect 5139 1170 5143 1171
rect 5139 1165 5143 1166
rect 5243 1170 5247 1171
rect 5243 1165 5247 1166
rect 5339 1170 5343 1171
rect 5339 1165 5343 1166
rect 5379 1170 5383 1171
rect 5379 1165 5383 1166
rect 5515 1170 5519 1171
rect 5515 1165 5519 1166
rect 5663 1170 5667 1171
rect 5663 1165 5667 1166
rect 1975 1118 1979 1119
rect 158 1116 164 1117
rect 110 1115 116 1116
rect 110 1111 111 1115
rect 115 1111 116 1115
rect 158 1112 159 1116
rect 163 1112 164 1116
rect 158 1111 164 1112
rect 318 1116 324 1117
rect 318 1112 319 1116
rect 323 1112 324 1116
rect 318 1111 324 1112
rect 502 1116 508 1117
rect 502 1112 503 1116
rect 507 1112 508 1116
rect 502 1111 508 1112
rect 686 1116 692 1117
rect 686 1112 687 1116
rect 691 1112 692 1116
rect 686 1111 692 1112
rect 862 1116 868 1117
rect 862 1112 863 1116
rect 867 1112 868 1116
rect 862 1111 868 1112
rect 1030 1116 1036 1117
rect 1030 1112 1031 1116
rect 1035 1112 1036 1116
rect 1030 1111 1036 1112
rect 1198 1116 1204 1117
rect 1198 1112 1199 1116
rect 1203 1112 1204 1116
rect 1198 1111 1204 1112
rect 1358 1116 1364 1117
rect 1358 1112 1359 1116
rect 1363 1112 1364 1116
rect 1358 1111 1364 1112
rect 1518 1116 1524 1117
rect 1518 1112 1519 1116
rect 1523 1112 1524 1116
rect 1518 1111 1524 1112
rect 1678 1116 1684 1117
rect 1678 1112 1679 1116
rect 1683 1112 1684 1116
rect 1678 1111 1684 1112
rect 1814 1116 1820 1117
rect 1814 1112 1815 1116
rect 1819 1112 1820 1116
rect 1814 1111 1820 1112
rect 1934 1115 1940 1116
rect 1934 1111 1935 1115
rect 1939 1111 1940 1115
rect 1975 1113 1979 1114
rect 1995 1118 1999 1119
rect 1995 1113 1999 1114
rect 2171 1118 2175 1119
rect 2171 1113 2175 1114
rect 2363 1118 2367 1119
rect 2363 1113 2367 1114
rect 2547 1118 2551 1119
rect 2547 1113 2551 1114
rect 2627 1118 2631 1119
rect 2627 1113 2631 1114
rect 2723 1118 2727 1119
rect 2723 1113 2727 1114
rect 2803 1118 2807 1119
rect 2803 1113 2807 1114
rect 2891 1118 2895 1119
rect 2891 1113 2895 1114
rect 2979 1118 2983 1119
rect 2979 1113 2983 1114
rect 3059 1118 3063 1119
rect 3059 1113 3063 1114
rect 3155 1118 3159 1119
rect 3155 1113 3159 1114
rect 3219 1118 3223 1119
rect 3219 1113 3223 1114
rect 3331 1118 3335 1119
rect 3331 1113 3335 1114
rect 3387 1118 3391 1119
rect 3387 1113 3391 1114
rect 3515 1118 3519 1119
rect 3515 1113 3519 1114
rect 3799 1118 3803 1119
rect 3799 1113 3803 1114
rect 110 1110 116 1111
rect 112 1075 114 1110
rect 160 1075 162 1111
rect 320 1075 322 1111
rect 504 1075 506 1111
rect 688 1075 690 1111
rect 864 1075 866 1111
rect 1032 1075 1034 1111
rect 1200 1075 1202 1111
rect 1360 1075 1362 1111
rect 1520 1075 1522 1111
rect 1680 1075 1682 1111
rect 1816 1075 1818 1111
rect 1934 1110 1940 1111
rect 1936 1075 1938 1110
rect 111 1074 115 1075
rect 111 1069 115 1070
rect 159 1074 163 1075
rect 159 1069 163 1070
rect 175 1074 179 1075
rect 175 1069 179 1070
rect 319 1074 323 1075
rect 319 1069 323 1070
rect 431 1074 435 1075
rect 431 1069 435 1070
rect 503 1074 507 1075
rect 503 1069 507 1070
rect 687 1074 691 1075
rect 687 1069 691 1070
rect 863 1074 867 1075
rect 863 1069 867 1070
rect 951 1074 955 1075
rect 951 1069 955 1070
rect 1031 1074 1035 1075
rect 1031 1069 1035 1070
rect 1199 1074 1203 1075
rect 1199 1069 1203 1070
rect 1215 1074 1219 1075
rect 1215 1069 1219 1070
rect 1359 1074 1363 1075
rect 1359 1069 1363 1070
rect 1519 1074 1523 1075
rect 1519 1069 1523 1070
rect 1679 1074 1683 1075
rect 1679 1069 1683 1070
rect 1815 1074 1819 1075
rect 1815 1069 1819 1070
rect 1935 1074 1939 1075
rect 1935 1069 1939 1070
rect 112 1046 114 1069
rect 110 1045 116 1046
rect 176 1045 178 1069
rect 432 1045 434 1069
rect 688 1045 690 1069
rect 952 1045 954 1069
rect 1216 1045 1218 1069
rect 1936 1046 1938 1069
rect 1976 1053 1978 1113
rect 1974 1052 1980 1053
rect 1996 1052 1998 1113
rect 2172 1052 2174 1113
rect 2364 1052 2366 1113
rect 2548 1052 2550 1113
rect 2724 1052 2726 1113
rect 2892 1052 2894 1113
rect 3060 1052 3062 1113
rect 3220 1052 3222 1113
rect 3388 1052 3390 1113
rect 3800 1053 3802 1113
rect 3840 1105 3842 1165
rect 3838 1104 3844 1105
rect 4836 1104 4838 1165
rect 4972 1104 4974 1165
rect 5108 1104 5110 1165
rect 5244 1104 5246 1165
rect 5380 1104 5382 1165
rect 5516 1104 5518 1165
rect 5664 1105 5666 1165
rect 5662 1104 5668 1105
rect 3838 1100 3839 1104
rect 3843 1100 3844 1104
rect 3838 1099 3844 1100
rect 4834 1103 4840 1104
rect 4834 1099 4835 1103
rect 4839 1099 4840 1103
rect 4834 1098 4840 1099
rect 4970 1103 4976 1104
rect 4970 1099 4971 1103
rect 4975 1099 4976 1103
rect 4970 1098 4976 1099
rect 5106 1103 5112 1104
rect 5106 1099 5107 1103
rect 5111 1099 5112 1103
rect 5106 1098 5112 1099
rect 5242 1103 5248 1104
rect 5242 1099 5243 1103
rect 5247 1099 5248 1103
rect 5242 1098 5248 1099
rect 5378 1103 5384 1104
rect 5378 1099 5379 1103
rect 5383 1099 5384 1103
rect 5378 1098 5384 1099
rect 5514 1103 5520 1104
rect 5514 1099 5515 1103
rect 5519 1099 5520 1103
rect 5662 1100 5663 1104
rect 5667 1100 5668 1104
rect 5662 1099 5668 1100
rect 5514 1098 5520 1099
rect 4862 1088 4868 1089
rect 3838 1087 3844 1088
rect 3838 1083 3839 1087
rect 3843 1083 3844 1087
rect 4862 1084 4863 1088
rect 4867 1084 4868 1088
rect 4862 1083 4868 1084
rect 4998 1088 5004 1089
rect 4998 1084 4999 1088
rect 5003 1084 5004 1088
rect 4998 1083 5004 1084
rect 5134 1088 5140 1089
rect 5134 1084 5135 1088
rect 5139 1084 5140 1088
rect 5134 1083 5140 1084
rect 5270 1088 5276 1089
rect 5270 1084 5271 1088
rect 5275 1084 5276 1088
rect 5270 1083 5276 1084
rect 5406 1088 5412 1089
rect 5406 1084 5407 1088
rect 5411 1084 5412 1088
rect 5406 1083 5412 1084
rect 5542 1088 5548 1089
rect 5542 1084 5543 1088
rect 5547 1084 5548 1088
rect 5542 1083 5548 1084
rect 5662 1087 5668 1088
rect 5662 1083 5663 1087
rect 5667 1083 5668 1087
rect 3838 1082 3844 1083
rect 3840 1055 3842 1082
rect 4864 1055 4866 1083
rect 5000 1055 5002 1083
rect 5136 1055 5138 1083
rect 5272 1055 5274 1083
rect 5408 1055 5410 1083
rect 5544 1055 5546 1083
rect 5662 1082 5668 1083
rect 5664 1055 5666 1082
rect 3839 1054 3843 1055
rect 3798 1052 3804 1053
rect 1974 1048 1975 1052
rect 1979 1048 1980 1052
rect 1974 1047 1980 1048
rect 1994 1051 2000 1052
rect 1994 1047 1995 1051
rect 1999 1047 2000 1051
rect 1994 1046 2000 1047
rect 2170 1051 2176 1052
rect 2170 1047 2171 1051
rect 2175 1047 2176 1051
rect 2170 1046 2176 1047
rect 2362 1051 2368 1052
rect 2362 1047 2363 1051
rect 2367 1047 2368 1051
rect 2362 1046 2368 1047
rect 2546 1051 2552 1052
rect 2546 1047 2547 1051
rect 2551 1047 2552 1051
rect 2546 1046 2552 1047
rect 2722 1051 2728 1052
rect 2722 1047 2723 1051
rect 2727 1047 2728 1051
rect 2722 1046 2728 1047
rect 2890 1051 2896 1052
rect 2890 1047 2891 1051
rect 2895 1047 2896 1051
rect 2890 1046 2896 1047
rect 3058 1051 3064 1052
rect 3058 1047 3059 1051
rect 3063 1047 3064 1051
rect 3058 1046 3064 1047
rect 3218 1051 3224 1052
rect 3218 1047 3219 1051
rect 3223 1047 3224 1051
rect 3218 1046 3224 1047
rect 3386 1051 3392 1052
rect 3386 1047 3387 1051
rect 3391 1047 3392 1051
rect 3798 1048 3799 1052
rect 3803 1048 3804 1052
rect 3839 1049 3843 1050
rect 4807 1054 4811 1055
rect 4807 1049 4811 1050
rect 4863 1054 4867 1055
rect 4863 1049 4867 1050
rect 4943 1054 4947 1055
rect 4943 1049 4947 1050
rect 4999 1054 5003 1055
rect 4999 1049 5003 1050
rect 5079 1054 5083 1055
rect 5079 1049 5083 1050
rect 5135 1054 5139 1055
rect 5135 1049 5139 1050
rect 5215 1054 5219 1055
rect 5215 1049 5219 1050
rect 5271 1054 5275 1055
rect 5271 1049 5275 1050
rect 5351 1054 5355 1055
rect 5351 1049 5355 1050
rect 5407 1054 5411 1055
rect 5407 1049 5411 1050
rect 5487 1054 5491 1055
rect 5487 1049 5491 1050
rect 5543 1054 5547 1055
rect 5543 1049 5547 1050
rect 5663 1054 5667 1055
rect 5663 1049 5667 1050
rect 3798 1047 3804 1048
rect 3386 1046 3392 1047
rect 1934 1045 1940 1046
rect 110 1041 111 1045
rect 115 1041 116 1045
rect 110 1040 116 1041
rect 174 1044 180 1045
rect 174 1040 175 1044
rect 179 1040 180 1044
rect 174 1039 180 1040
rect 430 1044 436 1045
rect 430 1040 431 1044
rect 435 1040 436 1044
rect 430 1039 436 1040
rect 686 1044 692 1045
rect 686 1040 687 1044
rect 691 1040 692 1044
rect 686 1039 692 1040
rect 950 1044 956 1045
rect 950 1040 951 1044
rect 955 1040 956 1044
rect 950 1039 956 1040
rect 1214 1044 1220 1045
rect 1214 1040 1215 1044
rect 1219 1040 1220 1044
rect 1934 1041 1935 1045
rect 1939 1041 1940 1045
rect 1934 1040 1940 1041
rect 1214 1039 1220 1040
rect 2022 1036 2028 1037
rect 1974 1035 1980 1036
rect 1974 1031 1975 1035
rect 1979 1031 1980 1035
rect 2022 1032 2023 1036
rect 2027 1032 2028 1036
rect 2022 1031 2028 1032
rect 2198 1036 2204 1037
rect 2198 1032 2199 1036
rect 2203 1032 2204 1036
rect 2198 1031 2204 1032
rect 2390 1036 2396 1037
rect 2390 1032 2391 1036
rect 2395 1032 2396 1036
rect 2390 1031 2396 1032
rect 2574 1036 2580 1037
rect 2574 1032 2575 1036
rect 2579 1032 2580 1036
rect 2574 1031 2580 1032
rect 2750 1036 2756 1037
rect 2750 1032 2751 1036
rect 2755 1032 2756 1036
rect 2750 1031 2756 1032
rect 2918 1036 2924 1037
rect 2918 1032 2919 1036
rect 2923 1032 2924 1036
rect 2918 1031 2924 1032
rect 3086 1036 3092 1037
rect 3086 1032 3087 1036
rect 3091 1032 3092 1036
rect 3086 1031 3092 1032
rect 3246 1036 3252 1037
rect 3246 1032 3247 1036
rect 3251 1032 3252 1036
rect 3246 1031 3252 1032
rect 3414 1036 3420 1037
rect 3414 1032 3415 1036
rect 3419 1032 3420 1036
rect 3414 1031 3420 1032
rect 3798 1035 3804 1036
rect 3798 1031 3799 1035
rect 3803 1031 3804 1035
rect 1974 1030 1980 1031
rect 146 1029 152 1030
rect 110 1028 116 1029
rect 110 1024 111 1028
rect 115 1024 116 1028
rect 146 1025 147 1029
rect 151 1025 152 1029
rect 146 1024 152 1025
rect 402 1029 408 1030
rect 402 1025 403 1029
rect 407 1025 408 1029
rect 402 1024 408 1025
rect 658 1029 664 1030
rect 658 1025 659 1029
rect 663 1025 664 1029
rect 658 1024 664 1025
rect 922 1029 928 1030
rect 922 1025 923 1029
rect 927 1025 928 1029
rect 922 1024 928 1025
rect 1186 1029 1192 1030
rect 1186 1025 1187 1029
rect 1191 1025 1192 1029
rect 1186 1024 1192 1025
rect 1934 1028 1940 1029
rect 1934 1024 1935 1028
rect 1939 1024 1940 1028
rect 110 1023 116 1024
rect 112 951 114 1023
rect 148 951 150 1024
rect 404 951 406 1024
rect 660 951 662 1024
rect 924 951 926 1024
rect 1188 951 1190 1024
rect 1934 1023 1940 1024
rect 1936 951 1938 1023
rect 1976 1007 1978 1030
rect 2024 1007 2026 1031
rect 2200 1007 2202 1031
rect 2392 1007 2394 1031
rect 2576 1007 2578 1031
rect 2752 1007 2754 1031
rect 2920 1007 2922 1031
rect 3088 1007 3090 1031
rect 3248 1007 3250 1031
rect 3416 1007 3418 1031
rect 3798 1030 3804 1031
rect 3800 1007 3802 1030
rect 3840 1026 3842 1049
rect 3838 1025 3844 1026
rect 4808 1025 4810 1049
rect 4944 1025 4946 1049
rect 5080 1025 5082 1049
rect 5216 1025 5218 1049
rect 5352 1025 5354 1049
rect 5488 1025 5490 1049
rect 5664 1026 5666 1049
rect 5662 1025 5668 1026
rect 3838 1021 3839 1025
rect 3843 1021 3844 1025
rect 3838 1020 3844 1021
rect 4806 1024 4812 1025
rect 4806 1020 4807 1024
rect 4811 1020 4812 1024
rect 4806 1019 4812 1020
rect 4942 1024 4948 1025
rect 4942 1020 4943 1024
rect 4947 1020 4948 1024
rect 4942 1019 4948 1020
rect 5078 1024 5084 1025
rect 5078 1020 5079 1024
rect 5083 1020 5084 1024
rect 5078 1019 5084 1020
rect 5214 1024 5220 1025
rect 5214 1020 5215 1024
rect 5219 1020 5220 1024
rect 5214 1019 5220 1020
rect 5350 1024 5356 1025
rect 5350 1020 5351 1024
rect 5355 1020 5356 1024
rect 5350 1019 5356 1020
rect 5486 1024 5492 1025
rect 5486 1020 5487 1024
rect 5491 1020 5492 1024
rect 5662 1021 5663 1025
rect 5667 1021 5668 1025
rect 5662 1020 5668 1021
rect 5486 1019 5492 1020
rect 4778 1009 4784 1010
rect 3838 1008 3844 1009
rect 1975 1006 1979 1007
rect 1975 1001 1979 1002
rect 2023 1006 2027 1007
rect 2023 1001 2027 1002
rect 2191 1006 2195 1007
rect 2191 1001 2195 1002
rect 2199 1006 2203 1007
rect 2199 1001 2203 1002
rect 2375 1006 2379 1007
rect 2375 1001 2379 1002
rect 2391 1006 2395 1007
rect 2391 1001 2395 1002
rect 2567 1006 2571 1007
rect 2567 1001 2571 1002
rect 2575 1006 2579 1007
rect 2575 1001 2579 1002
rect 2751 1006 2755 1007
rect 2751 1001 2755 1002
rect 2759 1006 2763 1007
rect 2759 1001 2763 1002
rect 2919 1006 2923 1007
rect 2919 1001 2923 1002
rect 2943 1006 2947 1007
rect 2943 1001 2947 1002
rect 3087 1006 3091 1007
rect 3087 1001 3091 1002
rect 3127 1006 3131 1007
rect 3127 1001 3131 1002
rect 3247 1006 3251 1007
rect 3247 1001 3251 1002
rect 3311 1006 3315 1007
rect 3311 1001 3315 1002
rect 3415 1006 3419 1007
rect 3415 1001 3419 1002
rect 3495 1006 3499 1007
rect 3495 1001 3499 1002
rect 3679 1006 3683 1007
rect 3679 1001 3683 1002
rect 3799 1006 3803 1007
rect 3838 1004 3839 1008
rect 3843 1004 3844 1008
rect 4778 1005 4779 1009
rect 4783 1005 4784 1009
rect 4778 1004 4784 1005
rect 4914 1009 4920 1010
rect 4914 1005 4915 1009
rect 4919 1005 4920 1009
rect 4914 1004 4920 1005
rect 5050 1009 5056 1010
rect 5050 1005 5051 1009
rect 5055 1005 5056 1009
rect 5050 1004 5056 1005
rect 5186 1009 5192 1010
rect 5186 1005 5187 1009
rect 5191 1005 5192 1009
rect 5186 1004 5192 1005
rect 5322 1009 5328 1010
rect 5322 1005 5323 1009
rect 5327 1005 5328 1009
rect 5322 1004 5328 1005
rect 5458 1009 5464 1010
rect 5458 1005 5459 1009
rect 5463 1005 5464 1009
rect 5458 1004 5464 1005
rect 5662 1008 5668 1009
rect 5662 1004 5663 1008
rect 5667 1004 5668 1008
rect 3838 1003 3844 1004
rect 3799 1001 3803 1002
rect 1976 978 1978 1001
rect 1974 977 1980 978
rect 2024 977 2026 1001
rect 2192 977 2194 1001
rect 2376 977 2378 1001
rect 2568 977 2570 1001
rect 2760 977 2762 1001
rect 2944 977 2946 1001
rect 3128 977 3130 1001
rect 3312 977 3314 1001
rect 3496 977 3498 1001
rect 3680 977 3682 1001
rect 3800 978 3802 1001
rect 3798 977 3804 978
rect 1974 973 1975 977
rect 1979 973 1980 977
rect 1974 972 1980 973
rect 2022 976 2028 977
rect 2022 972 2023 976
rect 2027 972 2028 976
rect 2022 971 2028 972
rect 2190 976 2196 977
rect 2190 972 2191 976
rect 2195 972 2196 976
rect 2190 971 2196 972
rect 2374 976 2380 977
rect 2374 972 2375 976
rect 2379 972 2380 976
rect 2374 971 2380 972
rect 2566 976 2572 977
rect 2566 972 2567 976
rect 2571 972 2572 976
rect 2566 971 2572 972
rect 2758 976 2764 977
rect 2758 972 2759 976
rect 2763 972 2764 976
rect 2758 971 2764 972
rect 2942 976 2948 977
rect 2942 972 2943 976
rect 2947 972 2948 976
rect 2942 971 2948 972
rect 3126 976 3132 977
rect 3126 972 3127 976
rect 3131 972 3132 976
rect 3126 971 3132 972
rect 3310 976 3316 977
rect 3310 972 3311 976
rect 3315 972 3316 976
rect 3310 971 3316 972
rect 3494 976 3500 977
rect 3494 972 3495 976
rect 3499 972 3500 976
rect 3494 971 3500 972
rect 3678 976 3684 977
rect 3678 972 3679 976
rect 3683 972 3684 976
rect 3798 973 3799 977
rect 3803 973 3804 977
rect 3798 972 3804 973
rect 3678 971 3684 972
rect 1994 961 2000 962
rect 1974 960 1980 961
rect 1974 956 1975 960
rect 1979 956 1980 960
rect 1994 957 1995 961
rect 1999 957 2000 961
rect 1994 956 2000 957
rect 2162 961 2168 962
rect 2162 957 2163 961
rect 2167 957 2168 961
rect 2162 956 2168 957
rect 2346 961 2352 962
rect 2346 957 2347 961
rect 2351 957 2352 961
rect 2346 956 2352 957
rect 2538 961 2544 962
rect 2538 957 2539 961
rect 2543 957 2544 961
rect 2538 956 2544 957
rect 2730 961 2736 962
rect 2730 957 2731 961
rect 2735 957 2736 961
rect 2730 956 2736 957
rect 2914 961 2920 962
rect 2914 957 2915 961
rect 2919 957 2920 961
rect 2914 956 2920 957
rect 3098 961 3104 962
rect 3098 957 3099 961
rect 3103 957 3104 961
rect 3098 956 3104 957
rect 3282 961 3288 962
rect 3282 957 3283 961
rect 3287 957 3288 961
rect 3282 956 3288 957
rect 3466 961 3472 962
rect 3466 957 3467 961
rect 3471 957 3472 961
rect 3466 956 3472 957
rect 3650 961 3656 962
rect 3650 957 3651 961
rect 3655 957 3656 961
rect 3650 956 3656 957
rect 3798 960 3804 961
rect 3798 956 3799 960
rect 3803 956 3804 960
rect 1974 955 1980 956
rect 111 950 115 951
rect 111 945 115 946
rect 147 950 151 951
rect 147 945 151 946
rect 235 950 239 951
rect 235 945 239 946
rect 403 950 407 951
rect 403 945 407 946
rect 459 950 463 951
rect 459 945 463 946
rect 659 950 663 951
rect 659 945 663 946
rect 683 950 687 951
rect 683 945 687 946
rect 907 950 911 951
rect 907 945 911 946
rect 923 950 927 951
rect 923 945 927 946
rect 1131 950 1135 951
rect 1131 945 1135 946
rect 1187 950 1191 951
rect 1187 945 1191 946
rect 1363 950 1367 951
rect 1363 945 1367 946
rect 1935 950 1939 951
rect 1935 945 1939 946
rect 112 885 114 945
rect 110 884 116 885
rect 236 884 238 945
rect 460 884 462 945
rect 684 884 686 945
rect 908 884 910 945
rect 1132 884 1134 945
rect 1364 884 1366 945
rect 1936 885 1938 945
rect 1976 891 1978 955
rect 1996 891 1998 956
rect 2164 891 2166 956
rect 2348 891 2350 956
rect 2540 891 2542 956
rect 2732 891 2734 956
rect 2916 891 2918 956
rect 3100 891 3102 956
rect 3284 891 3286 956
rect 3468 891 3470 956
rect 3652 891 3654 956
rect 3798 955 3804 956
rect 3800 891 3802 955
rect 3840 939 3842 1003
rect 4780 939 4782 1004
rect 4916 939 4918 1004
rect 5052 939 5054 1004
rect 5188 939 5190 1004
rect 5324 939 5326 1004
rect 5460 939 5462 1004
rect 5662 1003 5668 1004
rect 5664 939 5666 1003
rect 3839 938 3843 939
rect 3839 933 3843 934
rect 3859 938 3863 939
rect 3859 933 3863 934
rect 3995 938 3999 939
rect 3995 933 3999 934
rect 4171 938 4175 939
rect 4171 933 4175 934
rect 4387 938 4391 939
rect 4387 933 4391 934
rect 4643 938 4647 939
rect 4643 933 4647 934
rect 4779 938 4783 939
rect 4779 933 4783 934
rect 4915 938 4919 939
rect 4915 933 4919 934
rect 4931 938 4935 939
rect 4931 933 4935 934
rect 5051 938 5055 939
rect 5051 933 5055 934
rect 5187 938 5191 939
rect 5187 933 5191 934
rect 5235 938 5239 939
rect 5235 933 5239 934
rect 5323 938 5327 939
rect 5323 933 5327 934
rect 5459 938 5463 939
rect 5459 933 5463 934
rect 5515 938 5519 939
rect 5515 933 5519 934
rect 5663 938 5667 939
rect 5663 933 5667 934
rect 1975 890 1979 891
rect 1975 885 1979 886
rect 1995 890 1999 891
rect 1995 885 1999 886
rect 2163 890 2167 891
rect 2163 885 2167 886
rect 2179 890 2183 891
rect 2179 885 2183 886
rect 2347 890 2351 891
rect 2347 885 2351 886
rect 2403 890 2407 891
rect 2403 885 2407 886
rect 2539 890 2543 891
rect 2539 885 2543 886
rect 2675 890 2679 891
rect 2675 885 2679 886
rect 2731 890 2735 891
rect 2731 885 2735 886
rect 2915 890 2919 891
rect 2915 885 2919 886
rect 2987 890 2991 891
rect 2987 885 2991 886
rect 3099 890 3103 891
rect 3099 885 3103 886
rect 3283 890 3287 891
rect 3283 885 3287 886
rect 3323 890 3327 891
rect 3323 885 3327 886
rect 3467 890 3471 891
rect 3467 885 3471 886
rect 3651 890 3655 891
rect 3651 885 3655 886
rect 3799 890 3803 891
rect 3799 885 3803 886
rect 1934 884 1940 885
rect 110 880 111 884
rect 115 880 116 884
rect 110 879 116 880
rect 234 883 240 884
rect 234 879 235 883
rect 239 879 240 883
rect 234 878 240 879
rect 458 883 464 884
rect 458 879 459 883
rect 463 879 464 883
rect 458 878 464 879
rect 682 883 688 884
rect 682 879 683 883
rect 687 879 688 883
rect 682 878 688 879
rect 906 883 912 884
rect 906 879 907 883
rect 911 879 912 883
rect 906 878 912 879
rect 1130 883 1136 884
rect 1130 879 1131 883
rect 1135 879 1136 883
rect 1130 878 1136 879
rect 1362 883 1368 884
rect 1362 879 1363 883
rect 1367 879 1368 883
rect 1934 880 1935 884
rect 1939 880 1940 884
rect 1934 879 1940 880
rect 1362 878 1368 879
rect 262 868 268 869
rect 110 867 116 868
rect 110 863 111 867
rect 115 863 116 867
rect 262 864 263 868
rect 267 864 268 868
rect 262 863 268 864
rect 486 868 492 869
rect 486 864 487 868
rect 491 864 492 868
rect 486 863 492 864
rect 710 868 716 869
rect 710 864 711 868
rect 715 864 716 868
rect 710 863 716 864
rect 934 868 940 869
rect 934 864 935 868
rect 939 864 940 868
rect 934 863 940 864
rect 1158 868 1164 869
rect 1158 864 1159 868
rect 1163 864 1164 868
rect 1158 863 1164 864
rect 1390 868 1396 869
rect 1390 864 1391 868
rect 1395 864 1396 868
rect 1390 863 1396 864
rect 1934 867 1940 868
rect 1934 863 1935 867
rect 1939 863 1940 867
rect 110 862 116 863
rect 112 823 114 862
rect 264 823 266 863
rect 488 823 490 863
rect 712 823 714 863
rect 936 823 938 863
rect 1160 823 1162 863
rect 1392 823 1394 863
rect 1934 862 1940 863
rect 1936 823 1938 862
rect 1976 825 1978 885
rect 1974 824 1980 825
rect 1996 824 1998 885
rect 2180 824 2182 885
rect 2404 824 2406 885
rect 2676 824 2678 885
rect 2988 824 2990 885
rect 3324 824 3326 885
rect 3652 824 3654 885
rect 3800 825 3802 885
rect 3840 873 3842 933
rect 3838 872 3844 873
rect 3860 872 3862 933
rect 3996 872 3998 933
rect 4172 872 4174 933
rect 4388 872 4390 933
rect 4644 872 4646 933
rect 4932 872 4934 933
rect 5236 872 5238 933
rect 5516 872 5518 933
rect 5664 873 5666 933
rect 5662 872 5668 873
rect 3838 868 3839 872
rect 3843 868 3844 872
rect 3838 867 3844 868
rect 3858 871 3864 872
rect 3858 867 3859 871
rect 3863 867 3864 871
rect 3858 866 3864 867
rect 3994 871 4000 872
rect 3994 867 3995 871
rect 3999 867 4000 871
rect 3994 866 4000 867
rect 4170 871 4176 872
rect 4170 867 4171 871
rect 4175 867 4176 871
rect 4170 866 4176 867
rect 4386 871 4392 872
rect 4386 867 4387 871
rect 4391 867 4392 871
rect 4386 866 4392 867
rect 4642 871 4648 872
rect 4642 867 4643 871
rect 4647 867 4648 871
rect 4642 866 4648 867
rect 4930 871 4936 872
rect 4930 867 4931 871
rect 4935 867 4936 871
rect 4930 866 4936 867
rect 5234 871 5240 872
rect 5234 867 5235 871
rect 5239 867 5240 871
rect 5234 866 5240 867
rect 5514 871 5520 872
rect 5514 867 5515 871
rect 5519 867 5520 871
rect 5662 868 5663 872
rect 5667 868 5668 872
rect 5662 867 5668 868
rect 5514 866 5520 867
rect 3886 856 3892 857
rect 3838 855 3844 856
rect 3838 851 3839 855
rect 3843 851 3844 855
rect 3886 852 3887 856
rect 3891 852 3892 856
rect 3886 851 3892 852
rect 4022 856 4028 857
rect 4022 852 4023 856
rect 4027 852 4028 856
rect 4022 851 4028 852
rect 4198 856 4204 857
rect 4198 852 4199 856
rect 4203 852 4204 856
rect 4198 851 4204 852
rect 4414 856 4420 857
rect 4414 852 4415 856
rect 4419 852 4420 856
rect 4414 851 4420 852
rect 4670 856 4676 857
rect 4670 852 4671 856
rect 4675 852 4676 856
rect 4670 851 4676 852
rect 4958 856 4964 857
rect 4958 852 4959 856
rect 4963 852 4964 856
rect 4958 851 4964 852
rect 5262 856 5268 857
rect 5262 852 5263 856
rect 5267 852 5268 856
rect 5262 851 5268 852
rect 5542 856 5548 857
rect 5542 852 5543 856
rect 5547 852 5548 856
rect 5542 851 5548 852
rect 5662 855 5668 856
rect 5662 851 5663 855
rect 5667 851 5668 855
rect 3838 850 3844 851
rect 3840 827 3842 850
rect 3888 827 3890 851
rect 4024 827 4026 851
rect 4200 827 4202 851
rect 4416 827 4418 851
rect 4672 827 4674 851
rect 4960 827 4962 851
rect 5264 827 5266 851
rect 5544 827 5546 851
rect 5662 850 5668 851
rect 5664 827 5666 850
rect 3839 826 3843 827
rect 3798 824 3804 825
rect 111 822 115 823
rect 111 817 115 818
rect 175 822 179 823
rect 175 817 179 818
rect 263 822 267 823
rect 263 817 267 818
rect 431 822 435 823
rect 431 817 435 818
rect 487 822 491 823
rect 487 817 491 818
rect 671 822 675 823
rect 671 817 675 818
rect 711 822 715 823
rect 711 817 715 818
rect 903 822 907 823
rect 903 817 907 818
rect 935 822 939 823
rect 935 817 939 818
rect 1127 822 1131 823
rect 1127 817 1131 818
rect 1159 822 1163 823
rect 1159 817 1163 818
rect 1351 822 1355 823
rect 1351 817 1355 818
rect 1391 822 1395 823
rect 1391 817 1395 818
rect 1575 822 1579 823
rect 1575 817 1579 818
rect 1935 822 1939 823
rect 1974 820 1975 824
rect 1979 820 1980 824
rect 1974 819 1980 820
rect 1994 823 2000 824
rect 1994 819 1995 823
rect 1999 819 2000 823
rect 1994 818 2000 819
rect 2178 823 2184 824
rect 2178 819 2179 823
rect 2183 819 2184 823
rect 2178 818 2184 819
rect 2402 823 2408 824
rect 2402 819 2403 823
rect 2407 819 2408 823
rect 2402 818 2408 819
rect 2674 823 2680 824
rect 2674 819 2675 823
rect 2679 819 2680 823
rect 2674 818 2680 819
rect 2986 823 2992 824
rect 2986 819 2987 823
rect 2991 819 2992 823
rect 2986 818 2992 819
rect 3322 823 3328 824
rect 3322 819 3323 823
rect 3327 819 3328 823
rect 3322 818 3328 819
rect 3650 823 3656 824
rect 3650 819 3651 823
rect 3655 819 3656 823
rect 3798 820 3799 824
rect 3803 820 3804 824
rect 3839 821 3843 822
rect 3887 826 3891 827
rect 3887 821 3891 822
rect 4023 826 4027 827
rect 4023 821 4027 822
rect 4159 826 4163 827
rect 4159 821 4163 822
rect 4199 826 4203 827
rect 4199 821 4203 822
rect 4295 826 4299 827
rect 4295 821 4299 822
rect 4415 826 4419 827
rect 4415 821 4419 822
rect 4431 826 4435 827
rect 4431 821 4435 822
rect 4567 826 4571 827
rect 4567 821 4571 822
rect 4671 826 4675 827
rect 4671 821 4675 822
rect 4719 826 4723 827
rect 4719 821 4723 822
rect 4895 826 4899 827
rect 4895 821 4899 822
rect 4959 826 4963 827
rect 4959 821 4963 822
rect 5087 826 5091 827
rect 5087 821 5091 822
rect 5263 826 5267 827
rect 5263 821 5267 822
rect 5287 826 5291 827
rect 5287 821 5291 822
rect 5487 826 5491 827
rect 5487 821 5491 822
rect 5543 826 5547 827
rect 5543 821 5547 822
rect 5663 826 5667 827
rect 5663 821 5667 822
rect 3798 819 3804 820
rect 3650 818 3656 819
rect 1935 817 1939 818
rect 112 794 114 817
rect 110 793 116 794
rect 176 793 178 817
rect 432 793 434 817
rect 672 793 674 817
rect 904 793 906 817
rect 1128 793 1130 817
rect 1352 793 1354 817
rect 1576 793 1578 817
rect 1936 794 1938 817
rect 2022 808 2028 809
rect 1974 807 1980 808
rect 1974 803 1975 807
rect 1979 803 1980 807
rect 2022 804 2023 808
rect 2027 804 2028 808
rect 2022 803 2028 804
rect 2206 808 2212 809
rect 2206 804 2207 808
rect 2211 804 2212 808
rect 2206 803 2212 804
rect 2430 808 2436 809
rect 2430 804 2431 808
rect 2435 804 2436 808
rect 2430 803 2436 804
rect 2702 808 2708 809
rect 2702 804 2703 808
rect 2707 804 2708 808
rect 2702 803 2708 804
rect 3014 808 3020 809
rect 3014 804 3015 808
rect 3019 804 3020 808
rect 3014 803 3020 804
rect 3350 808 3356 809
rect 3350 804 3351 808
rect 3355 804 3356 808
rect 3350 803 3356 804
rect 3678 808 3684 809
rect 3678 804 3679 808
rect 3683 804 3684 808
rect 3678 803 3684 804
rect 3798 807 3804 808
rect 3798 803 3799 807
rect 3803 803 3804 807
rect 1974 802 1980 803
rect 1934 793 1940 794
rect 110 789 111 793
rect 115 789 116 793
rect 110 788 116 789
rect 174 792 180 793
rect 174 788 175 792
rect 179 788 180 792
rect 174 787 180 788
rect 430 792 436 793
rect 430 788 431 792
rect 435 788 436 792
rect 430 787 436 788
rect 670 792 676 793
rect 670 788 671 792
rect 675 788 676 792
rect 670 787 676 788
rect 902 792 908 793
rect 902 788 903 792
rect 907 788 908 792
rect 902 787 908 788
rect 1126 792 1132 793
rect 1126 788 1127 792
rect 1131 788 1132 792
rect 1126 787 1132 788
rect 1350 792 1356 793
rect 1350 788 1351 792
rect 1355 788 1356 792
rect 1350 787 1356 788
rect 1574 792 1580 793
rect 1574 788 1575 792
rect 1579 788 1580 792
rect 1934 789 1935 793
rect 1939 789 1940 793
rect 1934 788 1940 789
rect 1574 787 1580 788
rect 146 777 152 778
rect 110 776 116 777
rect 110 772 111 776
rect 115 772 116 776
rect 146 773 147 777
rect 151 773 152 777
rect 146 772 152 773
rect 402 777 408 778
rect 402 773 403 777
rect 407 773 408 777
rect 402 772 408 773
rect 642 777 648 778
rect 642 773 643 777
rect 647 773 648 777
rect 642 772 648 773
rect 874 777 880 778
rect 874 773 875 777
rect 879 773 880 777
rect 874 772 880 773
rect 1098 777 1104 778
rect 1098 773 1099 777
rect 1103 773 1104 777
rect 1098 772 1104 773
rect 1322 777 1328 778
rect 1322 773 1323 777
rect 1327 773 1328 777
rect 1322 772 1328 773
rect 1546 777 1552 778
rect 1546 773 1547 777
rect 1551 773 1552 777
rect 1546 772 1552 773
rect 1934 776 1940 777
rect 1934 772 1935 776
rect 1939 772 1940 776
rect 110 771 116 772
rect 112 711 114 771
rect 148 711 150 772
rect 404 711 406 772
rect 644 711 646 772
rect 876 711 878 772
rect 1100 711 1102 772
rect 1324 711 1326 772
rect 1548 711 1550 772
rect 1934 771 1940 772
rect 1936 711 1938 771
rect 111 710 115 711
rect 111 705 115 706
rect 131 710 135 711
rect 131 705 135 706
rect 147 710 151 711
rect 147 705 151 706
rect 315 710 319 711
rect 315 705 319 706
rect 403 710 407 711
rect 403 705 407 706
rect 523 710 527 711
rect 523 705 527 706
rect 643 710 647 711
rect 643 705 647 706
rect 723 710 727 711
rect 723 705 727 706
rect 875 710 879 711
rect 875 705 879 706
rect 907 710 911 711
rect 907 705 911 706
rect 1083 710 1087 711
rect 1083 705 1087 706
rect 1099 710 1103 711
rect 1099 705 1103 706
rect 1259 710 1263 711
rect 1259 705 1263 706
rect 1323 710 1327 711
rect 1323 705 1327 706
rect 1427 710 1431 711
rect 1427 705 1431 706
rect 1547 710 1551 711
rect 1547 705 1551 706
rect 1595 710 1599 711
rect 1595 705 1599 706
rect 1771 710 1775 711
rect 1771 705 1775 706
rect 1935 710 1939 711
rect 1935 705 1939 706
rect 112 645 114 705
rect 110 644 116 645
rect 132 644 134 705
rect 316 644 318 705
rect 524 644 526 705
rect 724 644 726 705
rect 908 644 910 705
rect 1084 644 1086 705
rect 1260 644 1262 705
rect 1428 644 1430 705
rect 1596 644 1598 705
rect 1772 644 1774 705
rect 1936 645 1938 705
rect 1934 644 1940 645
rect 110 640 111 644
rect 115 640 116 644
rect 110 639 116 640
rect 130 643 136 644
rect 130 639 131 643
rect 135 639 136 643
rect 130 638 136 639
rect 314 643 320 644
rect 314 639 315 643
rect 319 639 320 643
rect 314 638 320 639
rect 522 643 528 644
rect 522 639 523 643
rect 527 639 528 643
rect 522 638 528 639
rect 722 643 728 644
rect 722 639 723 643
rect 727 639 728 643
rect 722 638 728 639
rect 906 643 912 644
rect 906 639 907 643
rect 911 639 912 643
rect 906 638 912 639
rect 1082 643 1088 644
rect 1082 639 1083 643
rect 1087 639 1088 643
rect 1082 638 1088 639
rect 1258 643 1264 644
rect 1258 639 1259 643
rect 1263 639 1264 643
rect 1258 638 1264 639
rect 1426 643 1432 644
rect 1426 639 1427 643
rect 1431 639 1432 643
rect 1426 638 1432 639
rect 1594 643 1600 644
rect 1594 639 1595 643
rect 1599 639 1600 643
rect 1594 638 1600 639
rect 1770 643 1776 644
rect 1770 639 1771 643
rect 1775 639 1776 643
rect 1934 640 1935 644
rect 1939 640 1940 644
rect 1934 639 1940 640
rect 1770 638 1776 639
rect 158 628 164 629
rect 110 627 116 628
rect 110 623 111 627
rect 115 623 116 627
rect 158 624 159 628
rect 163 624 164 628
rect 158 623 164 624
rect 342 628 348 629
rect 342 624 343 628
rect 347 624 348 628
rect 342 623 348 624
rect 550 628 556 629
rect 550 624 551 628
rect 555 624 556 628
rect 550 623 556 624
rect 750 628 756 629
rect 750 624 751 628
rect 755 624 756 628
rect 750 623 756 624
rect 934 628 940 629
rect 934 624 935 628
rect 939 624 940 628
rect 934 623 940 624
rect 1110 628 1116 629
rect 1110 624 1111 628
rect 1115 624 1116 628
rect 1110 623 1116 624
rect 1286 628 1292 629
rect 1286 624 1287 628
rect 1291 624 1292 628
rect 1286 623 1292 624
rect 1454 628 1460 629
rect 1454 624 1455 628
rect 1459 624 1460 628
rect 1454 623 1460 624
rect 1622 628 1628 629
rect 1622 624 1623 628
rect 1627 624 1628 628
rect 1622 623 1628 624
rect 1798 628 1804 629
rect 1798 624 1799 628
rect 1803 624 1804 628
rect 1798 623 1804 624
rect 1934 627 1940 628
rect 1934 623 1935 627
rect 1939 623 1940 627
rect 110 622 116 623
rect 112 599 114 622
rect 160 599 162 623
rect 344 599 346 623
rect 552 599 554 623
rect 752 599 754 623
rect 936 599 938 623
rect 1112 599 1114 623
rect 1288 599 1290 623
rect 1456 599 1458 623
rect 1624 599 1626 623
rect 1800 599 1802 623
rect 1934 622 1940 623
rect 1936 599 1938 622
rect 111 598 115 599
rect 111 593 115 594
rect 159 598 163 599
rect 159 593 163 594
rect 343 598 347 599
rect 343 593 347 594
rect 375 598 379 599
rect 375 593 379 594
rect 551 598 555 599
rect 551 593 555 594
rect 599 598 603 599
rect 599 593 603 594
rect 751 598 755 599
rect 751 593 755 594
rect 807 598 811 599
rect 807 593 811 594
rect 935 598 939 599
rect 935 593 939 594
rect 999 598 1003 599
rect 999 593 1003 594
rect 1111 598 1115 599
rect 1111 593 1115 594
rect 1175 598 1179 599
rect 1175 593 1179 594
rect 1287 598 1291 599
rect 1287 593 1291 594
rect 1343 598 1347 599
rect 1343 593 1347 594
rect 1455 598 1459 599
rect 1455 593 1459 594
rect 1511 598 1515 599
rect 1511 593 1515 594
rect 1623 598 1627 599
rect 1623 593 1627 594
rect 1671 598 1675 599
rect 1671 593 1675 594
rect 1799 598 1803 599
rect 1799 593 1803 594
rect 1815 598 1819 599
rect 1815 593 1819 594
rect 1935 598 1939 599
rect 1935 593 1939 594
rect 112 570 114 593
rect 110 569 116 570
rect 160 569 162 593
rect 376 569 378 593
rect 600 569 602 593
rect 808 569 810 593
rect 1000 569 1002 593
rect 1176 569 1178 593
rect 1344 569 1346 593
rect 1512 569 1514 593
rect 1672 569 1674 593
rect 1816 569 1818 593
rect 1936 570 1938 593
rect 1976 579 1978 802
rect 2024 579 2026 803
rect 2208 579 2210 803
rect 2432 579 2434 803
rect 2704 579 2706 803
rect 3016 579 3018 803
rect 3352 579 3354 803
rect 3680 579 3682 803
rect 3798 802 3804 803
rect 3800 579 3802 802
rect 3840 798 3842 821
rect 3838 797 3844 798
rect 3888 797 3890 821
rect 4024 797 4026 821
rect 4160 797 4162 821
rect 4296 797 4298 821
rect 4432 797 4434 821
rect 4568 797 4570 821
rect 4720 797 4722 821
rect 4896 797 4898 821
rect 5088 797 5090 821
rect 5288 797 5290 821
rect 5488 797 5490 821
rect 5664 798 5666 821
rect 5662 797 5668 798
rect 3838 793 3839 797
rect 3843 793 3844 797
rect 3838 792 3844 793
rect 3886 796 3892 797
rect 3886 792 3887 796
rect 3891 792 3892 796
rect 3886 791 3892 792
rect 4022 796 4028 797
rect 4022 792 4023 796
rect 4027 792 4028 796
rect 4022 791 4028 792
rect 4158 796 4164 797
rect 4158 792 4159 796
rect 4163 792 4164 796
rect 4158 791 4164 792
rect 4294 796 4300 797
rect 4294 792 4295 796
rect 4299 792 4300 796
rect 4294 791 4300 792
rect 4430 796 4436 797
rect 4430 792 4431 796
rect 4435 792 4436 796
rect 4430 791 4436 792
rect 4566 796 4572 797
rect 4566 792 4567 796
rect 4571 792 4572 796
rect 4566 791 4572 792
rect 4718 796 4724 797
rect 4718 792 4719 796
rect 4723 792 4724 796
rect 4718 791 4724 792
rect 4894 796 4900 797
rect 4894 792 4895 796
rect 4899 792 4900 796
rect 4894 791 4900 792
rect 5086 796 5092 797
rect 5086 792 5087 796
rect 5091 792 5092 796
rect 5086 791 5092 792
rect 5286 796 5292 797
rect 5286 792 5287 796
rect 5291 792 5292 796
rect 5286 791 5292 792
rect 5486 796 5492 797
rect 5486 792 5487 796
rect 5491 792 5492 796
rect 5662 793 5663 797
rect 5667 793 5668 797
rect 5662 792 5668 793
rect 5486 791 5492 792
rect 3858 781 3864 782
rect 3838 780 3844 781
rect 3838 776 3839 780
rect 3843 776 3844 780
rect 3858 777 3859 781
rect 3863 777 3864 781
rect 3858 776 3864 777
rect 3994 781 4000 782
rect 3994 777 3995 781
rect 3999 777 4000 781
rect 3994 776 4000 777
rect 4130 781 4136 782
rect 4130 777 4131 781
rect 4135 777 4136 781
rect 4130 776 4136 777
rect 4266 781 4272 782
rect 4266 777 4267 781
rect 4271 777 4272 781
rect 4266 776 4272 777
rect 4402 781 4408 782
rect 4402 777 4403 781
rect 4407 777 4408 781
rect 4402 776 4408 777
rect 4538 781 4544 782
rect 4538 777 4539 781
rect 4543 777 4544 781
rect 4538 776 4544 777
rect 4690 781 4696 782
rect 4690 777 4691 781
rect 4695 777 4696 781
rect 4690 776 4696 777
rect 4866 781 4872 782
rect 4866 777 4867 781
rect 4871 777 4872 781
rect 4866 776 4872 777
rect 5058 781 5064 782
rect 5058 777 5059 781
rect 5063 777 5064 781
rect 5058 776 5064 777
rect 5258 781 5264 782
rect 5258 777 5259 781
rect 5263 777 5264 781
rect 5258 776 5264 777
rect 5458 781 5464 782
rect 5458 777 5459 781
rect 5463 777 5464 781
rect 5458 776 5464 777
rect 5662 780 5668 781
rect 5662 776 5663 780
rect 5667 776 5668 780
rect 3838 775 3844 776
rect 3840 711 3842 775
rect 3860 711 3862 776
rect 3996 711 3998 776
rect 4132 711 4134 776
rect 4268 711 4270 776
rect 4404 711 4406 776
rect 4540 711 4542 776
rect 4692 711 4694 776
rect 4868 711 4870 776
rect 5060 711 5062 776
rect 5260 711 5262 776
rect 5460 711 5462 776
rect 5662 775 5668 776
rect 5664 711 5666 775
rect 3839 710 3843 711
rect 3839 705 3843 706
rect 3859 710 3863 711
rect 3859 705 3863 706
rect 3995 710 3999 711
rect 3995 705 3999 706
rect 4131 710 4135 711
rect 4131 705 4135 706
rect 4267 710 4271 711
rect 4267 705 4271 706
rect 4403 710 4407 711
rect 4403 705 4407 706
rect 4539 710 4543 711
rect 4539 705 4543 706
rect 4691 710 4695 711
rect 4691 705 4695 706
rect 4699 710 4703 711
rect 4699 705 4703 706
rect 4867 710 4871 711
rect 4867 705 4871 706
rect 4891 710 4895 711
rect 4891 705 4895 706
rect 5059 710 5063 711
rect 5059 705 5063 706
rect 5099 710 5103 711
rect 5099 705 5103 706
rect 5259 710 5263 711
rect 5259 705 5263 706
rect 5315 710 5319 711
rect 5315 705 5319 706
rect 5459 710 5463 711
rect 5459 705 5463 706
rect 5515 710 5519 711
rect 5515 705 5519 706
rect 5663 710 5667 711
rect 5663 705 5667 706
rect 3840 645 3842 705
rect 3838 644 3844 645
rect 3860 644 3862 705
rect 3996 644 3998 705
rect 4132 644 4134 705
rect 4268 644 4270 705
rect 4404 644 4406 705
rect 4540 644 4542 705
rect 4700 644 4702 705
rect 4892 644 4894 705
rect 5100 644 5102 705
rect 5316 644 5318 705
rect 5516 644 5518 705
rect 5664 645 5666 705
rect 5662 644 5668 645
rect 3838 640 3839 644
rect 3843 640 3844 644
rect 3838 639 3844 640
rect 3858 643 3864 644
rect 3858 639 3859 643
rect 3863 639 3864 643
rect 3858 638 3864 639
rect 3994 643 4000 644
rect 3994 639 3995 643
rect 3999 639 4000 643
rect 3994 638 4000 639
rect 4130 643 4136 644
rect 4130 639 4131 643
rect 4135 639 4136 643
rect 4130 638 4136 639
rect 4266 643 4272 644
rect 4266 639 4267 643
rect 4271 639 4272 643
rect 4266 638 4272 639
rect 4402 643 4408 644
rect 4402 639 4403 643
rect 4407 639 4408 643
rect 4402 638 4408 639
rect 4538 643 4544 644
rect 4538 639 4539 643
rect 4543 639 4544 643
rect 4538 638 4544 639
rect 4698 643 4704 644
rect 4698 639 4699 643
rect 4703 639 4704 643
rect 4698 638 4704 639
rect 4890 643 4896 644
rect 4890 639 4891 643
rect 4895 639 4896 643
rect 4890 638 4896 639
rect 5098 643 5104 644
rect 5098 639 5099 643
rect 5103 639 5104 643
rect 5098 638 5104 639
rect 5314 643 5320 644
rect 5314 639 5315 643
rect 5319 639 5320 643
rect 5314 638 5320 639
rect 5514 643 5520 644
rect 5514 639 5515 643
rect 5519 639 5520 643
rect 5662 640 5663 644
rect 5667 640 5668 644
rect 5662 639 5668 640
rect 5514 638 5520 639
rect 3886 628 3892 629
rect 3838 627 3844 628
rect 3838 623 3839 627
rect 3843 623 3844 627
rect 3886 624 3887 628
rect 3891 624 3892 628
rect 3886 623 3892 624
rect 4022 628 4028 629
rect 4022 624 4023 628
rect 4027 624 4028 628
rect 4022 623 4028 624
rect 4158 628 4164 629
rect 4158 624 4159 628
rect 4163 624 4164 628
rect 4158 623 4164 624
rect 4294 628 4300 629
rect 4294 624 4295 628
rect 4299 624 4300 628
rect 4294 623 4300 624
rect 4430 628 4436 629
rect 4430 624 4431 628
rect 4435 624 4436 628
rect 4430 623 4436 624
rect 4566 628 4572 629
rect 4566 624 4567 628
rect 4571 624 4572 628
rect 4566 623 4572 624
rect 4726 628 4732 629
rect 4726 624 4727 628
rect 4731 624 4732 628
rect 4726 623 4732 624
rect 4918 628 4924 629
rect 4918 624 4919 628
rect 4923 624 4924 628
rect 4918 623 4924 624
rect 5126 628 5132 629
rect 5126 624 5127 628
rect 5131 624 5132 628
rect 5126 623 5132 624
rect 5342 628 5348 629
rect 5342 624 5343 628
rect 5347 624 5348 628
rect 5342 623 5348 624
rect 5542 628 5548 629
rect 5542 624 5543 628
rect 5547 624 5548 628
rect 5542 623 5548 624
rect 5662 627 5668 628
rect 5662 623 5663 627
rect 5667 623 5668 627
rect 3838 622 3844 623
rect 3840 599 3842 622
rect 3888 599 3890 623
rect 4024 599 4026 623
rect 4160 599 4162 623
rect 4296 599 4298 623
rect 4432 599 4434 623
rect 4568 599 4570 623
rect 4728 599 4730 623
rect 4920 599 4922 623
rect 5128 599 5130 623
rect 5344 599 5346 623
rect 5544 599 5546 623
rect 5662 622 5668 623
rect 5664 599 5666 622
rect 3839 598 3843 599
rect 3839 593 3843 594
rect 3887 598 3891 599
rect 3887 593 3891 594
rect 4023 598 4027 599
rect 4023 593 4027 594
rect 4071 598 4075 599
rect 4071 593 4075 594
rect 4159 598 4163 599
rect 4159 593 4163 594
rect 4295 598 4299 599
rect 4295 593 4299 594
rect 4311 598 4315 599
rect 4311 593 4315 594
rect 4431 598 4435 599
rect 4431 593 4435 594
rect 4567 598 4571 599
rect 4567 593 4571 594
rect 4575 598 4579 599
rect 4575 593 4579 594
rect 4727 598 4731 599
rect 4727 593 4731 594
rect 4855 598 4859 599
rect 4855 593 4859 594
rect 4919 598 4923 599
rect 4919 593 4923 594
rect 5127 598 5131 599
rect 5127 593 5131 594
rect 5151 598 5155 599
rect 5151 593 5155 594
rect 5343 598 5347 599
rect 5343 593 5347 594
rect 5447 598 5451 599
rect 5447 593 5451 594
rect 5543 598 5547 599
rect 5543 593 5547 594
rect 5663 598 5667 599
rect 5663 593 5667 594
rect 1975 578 1979 579
rect 1975 573 1979 574
rect 2023 578 2027 579
rect 2023 573 2027 574
rect 2207 578 2211 579
rect 2207 573 2211 574
rect 2431 578 2435 579
rect 2431 573 2435 574
rect 2703 578 2707 579
rect 2703 573 2707 574
rect 3015 578 3019 579
rect 3015 573 3019 574
rect 3135 578 3139 579
rect 3135 573 3139 574
rect 3271 578 3275 579
rect 3271 573 3275 574
rect 3351 578 3355 579
rect 3351 573 3355 574
rect 3407 578 3411 579
rect 3407 573 3411 574
rect 3543 578 3547 579
rect 3543 573 3547 574
rect 3679 578 3683 579
rect 3679 573 3683 574
rect 3799 578 3803 579
rect 3799 573 3803 574
rect 1934 569 1940 570
rect 110 565 111 569
rect 115 565 116 569
rect 110 564 116 565
rect 158 568 164 569
rect 158 564 159 568
rect 163 564 164 568
rect 158 563 164 564
rect 374 568 380 569
rect 374 564 375 568
rect 379 564 380 568
rect 374 563 380 564
rect 598 568 604 569
rect 598 564 599 568
rect 603 564 604 568
rect 598 563 604 564
rect 806 568 812 569
rect 806 564 807 568
rect 811 564 812 568
rect 806 563 812 564
rect 998 568 1004 569
rect 998 564 999 568
rect 1003 564 1004 568
rect 998 563 1004 564
rect 1174 568 1180 569
rect 1174 564 1175 568
rect 1179 564 1180 568
rect 1174 563 1180 564
rect 1342 568 1348 569
rect 1342 564 1343 568
rect 1347 564 1348 568
rect 1342 563 1348 564
rect 1510 568 1516 569
rect 1510 564 1511 568
rect 1515 564 1516 568
rect 1510 563 1516 564
rect 1670 568 1676 569
rect 1670 564 1671 568
rect 1675 564 1676 568
rect 1670 563 1676 564
rect 1814 568 1820 569
rect 1814 564 1815 568
rect 1819 564 1820 568
rect 1934 565 1935 569
rect 1939 565 1940 569
rect 1934 564 1940 565
rect 1814 563 1820 564
rect 130 553 136 554
rect 110 552 116 553
rect 110 548 111 552
rect 115 548 116 552
rect 130 549 131 553
rect 135 549 136 553
rect 130 548 136 549
rect 346 553 352 554
rect 346 549 347 553
rect 351 549 352 553
rect 346 548 352 549
rect 570 553 576 554
rect 570 549 571 553
rect 575 549 576 553
rect 570 548 576 549
rect 778 553 784 554
rect 778 549 779 553
rect 783 549 784 553
rect 778 548 784 549
rect 970 553 976 554
rect 970 549 971 553
rect 975 549 976 553
rect 970 548 976 549
rect 1146 553 1152 554
rect 1146 549 1147 553
rect 1151 549 1152 553
rect 1146 548 1152 549
rect 1314 553 1320 554
rect 1314 549 1315 553
rect 1319 549 1320 553
rect 1314 548 1320 549
rect 1482 553 1488 554
rect 1482 549 1483 553
rect 1487 549 1488 553
rect 1482 548 1488 549
rect 1642 553 1648 554
rect 1642 549 1643 553
rect 1647 549 1648 553
rect 1642 548 1648 549
rect 1786 553 1792 554
rect 1786 549 1787 553
rect 1791 549 1792 553
rect 1786 548 1792 549
rect 1934 552 1940 553
rect 1934 548 1935 552
rect 1939 548 1940 552
rect 1976 550 1978 573
rect 110 547 116 548
rect 112 487 114 547
rect 132 487 134 548
rect 348 487 350 548
rect 572 487 574 548
rect 780 487 782 548
rect 972 487 974 548
rect 1148 487 1150 548
rect 1316 487 1318 548
rect 1484 487 1486 548
rect 1644 487 1646 548
rect 1788 487 1790 548
rect 1934 547 1940 548
rect 1974 549 1980 550
rect 3136 549 3138 573
rect 3272 549 3274 573
rect 3408 549 3410 573
rect 3544 549 3546 573
rect 3680 549 3682 573
rect 3800 550 3802 573
rect 3840 570 3842 593
rect 3838 569 3844 570
rect 3888 569 3890 593
rect 4072 569 4074 593
rect 4312 569 4314 593
rect 4576 569 4578 593
rect 4856 569 4858 593
rect 5152 569 5154 593
rect 5448 569 5450 593
rect 5664 570 5666 593
rect 5662 569 5668 570
rect 3838 565 3839 569
rect 3843 565 3844 569
rect 3838 564 3844 565
rect 3886 568 3892 569
rect 3886 564 3887 568
rect 3891 564 3892 568
rect 3886 563 3892 564
rect 4070 568 4076 569
rect 4070 564 4071 568
rect 4075 564 4076 568
rect 4070 563 4076 564
rect 4310 568 4316 569
rect 4310 564 4311 568
rect 4315 564 4316 568
rect 4310 563 4316 564
rect 4574 568 4580 569
rect 4574 564 4575 568
rect 4579 564 4580 568
rect 4574 563 4580 564
rect 4854 568 4860 569
rect 4854 564 4855 568
rect 4859 564 4860 568
rect 4854 563 4860 564
rect 5150 568 5156 569
rect 5150 564 5151 568
rect 5155 564 5156 568
rect 5150 563 5156 564
rect 5446 568 5452 569
rect 5446 564 5447 568
rect 5451 564 5452 568
rect 5662 565 5663 569
rect 5667 565 5668 569
rect 5662 564 5668 565
rect 5446 563 5452 564
rect 3858 553 3864 554
rect 3838 552 3844 553
rect 3798 549 3804 550
rect 1936 487 1938 547
rect 1974 545 1975 549
rect 1979 545 1980 549
rect 1974 544 1980 545
rect 3134 548 3140 549
rect 3134 544 3135 548
rect 3139 544 3140 548
rect 3134 543 3140 544
rect 3270 548 3276 549
rect 3270 544 3271 548
rect 3275 544 3276 548
rect 3270 543 3276 544
rect 3406 548 3412 549
rect 3406 544 3407 548
rect 3411 544 3412 548
rect 3406 543 3412 544
rect 3542 548 3548 549
rect 3542 544 3543 548
rect 3547 544 3548 548
rect 3542 543 3548 544
rect 3678 548 3684 549
rect 3678 544 3679 548
rect 3683 544 3684 548
rect 3798 545 3799 549
rect 3803 545 3804 549
rect 3838 548 3839 552
rect 3843 548 3844 552
rect 3858 549 3859 553
rect 3863 549 3864 553
rect 3858 548 3864 549
rect 4042 553 4048 554
rect 4042 549 4043 553
rect 4047 549 4048 553
rect 4042 548 4048 549
rect 4282 553 4288 554
rect 4282 549 4283 553
rect 4287 549 4288 553
rect 4282 548 4288 549
rect 4546 553 4552 554
rect 4546 549 4547 553
rect 4551 549 4552 553
rect 4546 548 4552 549
rect 4826 553 4832 554
rect 4826 549 4827 553
rect 4831 549 4832 553
rect 4826 548 4832 549
rect 5122 553 5128 554
rect 5122 549 5123 553
rect 5127 549 5128 553
rect 5122 548 5128 549
rect 5418 553 5424 554
rect 5418 549 5419 553
rect 5423 549 5424 553
rect 5418 548 5424 549
rect 5662 552 5668 553
rect 5662 548 5663 552
rect 5667 548 5668 552
rect 3838 547 3844 548
rect 3798 544 3804 545
rect 3678 543 3684 544
rect 3106 533 3112 534
rect 1974 532 1980 533
rect 1974 528 1975 532
rect 1979 528 1980 532
rect 3106 529 3107 533
rect 3111 529 3112 533
rect 3106 528 3112 529
rect 3242 533 3248 534
rect 3242 529 3243 533
rect 3247 529 3248 533
rect 3242 528 3248 529
rect 3378 533 3384 534
rect 3378 529 3379 533
rect 3383 529 3384 533
rect 3378 528 3384 529
rect 3514 533 3520 534
rect 3514 529 3515 533
rect 3519 529 3520 533
rect 3514 528 3520 529
rect 3650 533 3656 534
rect 3650 529 3651 533
rect 3655 529 3656 533
rect 3650 528 3656 529
rect 3798 532 3804 533
rect 3798 528 3799 532
rect 3803 528 3804 532
rect 1974 527 1980 528
rect 111 486 115 487
rect 111 481 115 482
rect 131 486 135 487
rect 131 481 135 482
rect 155 486 159 487
rect 155 481 159 482
rect 347 486 351 487
rect 347 481 351 482
rect 483 486 487 487
rect 483 481 487 482
rect 571 486 575 487
rect 571 481 575 482
rect 779 486 783 487
rect 779 481 783 482
rect 811 486 815 487
rect 811 481 815 482
rect 971 486 975 487
rect 971 481 975 482
rect 1139 486 1143 487
rect 1139 481 1143 482
rect 1147 486 1151 487
rect 1147 481 1151 482
rect 1315 486 1319 487
rect 1315 481 1319 482
rect 1475 486 1479 487
rect 1475 481 1479 482
rect 1483 486 1487 487
rect 1483 481 1487 482
rect 1643 486 1647 487
rect 1643 481 1647 482
rect 1787 486 1791 487
rect 1787 481 1791 482
rect 1935 486 1939 487
rect 1935 481 1939 482
rect 112 421 114 481
rect 110 420 116 421
rect 156 420 158 481
rect 484 420 486 481
rect 812 420 814 481
rect 1140 420 1142 481
rect 1476 420 1478 481
rect 1788 420 1790 481
rect 1936 421 1938 481
rect 1976 467 1978 527
rect 3108 467 3110 528
rect 3244 467 3246 528
rect 3380 467 3382 528
rect 3516 467 3518 528
rect 3652 467 3654 528
rect 3798 527 3804 528
rect 3800 467 3802 527
rect 3840 475 3842 547
rect 3860 475 3862 548
rect 4044 475 4046 548
rect 4284 475 4286 548
rect 4548 475 4550 548
rect 4828 475 4830 548
rect 5124 475 5126 548
rect 5420 475 5422 548
rect 5662 547 5668 548
rect 5664 475 5666 547
rect 3839 474 3843 475
rect 3839 469 3843 470
rect 3859 474 3863 475
rect 3859 469 3863 470
rect 4043 474 4047 475
rect 4043 469 4047 470
rect 4283 474 4287 475
rect 4283 469 4287 470
rect 4451 474 4455 475
rect 4451 469 4455 470
rect 4547 474 4551 475
rect 4547 469 4551 470
rect 4643 474 4647 475
rect 4643 469 4647 470
rect 4827 474 4831 475
rect 4827 469 4831 470
rect 4843 474 4847 475
rect 4843 469 4847 470
rect 5051 474 5055 475
rect 5051 469 5055 470
rect 5123 474 5127 475
rect 5123 469 5127 470
rect 5267 474 5271 475
rect 5267 469 5271 470
rect 5419 474 5423 475
rect 5419 469 5423 470
rect 5483 474 5487 475
rect 5483 469 5487 470
rect 5663 474 5667 475
rect 5663 469 5667 470
rect 1975 466 1979 467
rect 1975 461 1979 462
rect 1995 466 1999 467
rect 1995 461 1999 462
rect 2203 466 2207 467
rect 2203 461 2207 462
rect 2427 466 2431 467
rect 2427 461 2431 462
rect 2651 466 2655 467
rect 2651 461 2655 462
rect 2859 466 2863 467
rect 2859 461 2863 462
rect 3067 466 3071 467
rect 3067 461 3071 462
rect 3107 466 3111 467
rect 3107 461 3111 462
rect 3243 466 3247 467
rect 3243 461 3247 462
rect 3267 466 3271 467
rect 3267 461 3271 462
rect 3379 466 3383 467
rect 3379 461 3383 462
rect 3467 466 3471 467
rect 3467 461 3471 462
rect 3515 466 3519 467
rect 3515 461 3519 462
rect 3651 466 3655 467
rect 3651 461 3655 462
rect 3799 466 3803 467
rect 3799 461 3803 462
rect 1934 420 1940 421
rect 110 416 111 420
rect 115 416 116 420
rect 110 415 116 416
rect 154 419 160 420
rect 154 415 155 419
rect 159 415 160 419
rect 154 414 160 415
rect 482 419 488 420
rect 482 415 483 419
rect 487 415 488 419
rect 482 414 488 415
rect 810 419 816 420
rect 810 415 811 419
rect 815 415 816 419
rect 810 414 816 415
rect 1138 419 1144 420
rect 1138 415 1139 419
rect 1143 415 1144 419
rect 1138 414 1144 415
rect 1474 419 1480 420
rect 1474 415 1475 419
rect 1479 415 1480 419
rect 1474 414 1480 415
rect 1786 419 1792 420
rect 1786 415 1787 419
rect 1791 415 1792 419
rect 1934 416 1935 420
rect 1939 416 1940 420
rect 1934 415 1940 416
rect 1786 414 1792 415
rect 182 404 188 405
rect 110 403 116 404
rect 110 399 111 403
rect 115 399 116 403
rect 182 400 183 404
rect 187 400 188 404
rect 182 399 188 400
rect 510 404 516 405
rect 510 400 511 404
rect 515 400 516 404
rect 510 399 516 400
rect 838 404 844 405
rect 838 400 839 404
rect 843 400 844 404
rect 838 399 844 400
rect 1166 404 1172 405
rect 1166 400 1167 404
rect 1171 400 1172 404
rect 1166 399 1172 400
rect 1502 404 1508 405
rect 1502 400 1503 404
rect 1507 400 1508 404
rect 1502 399 1508 400
rect 1814 404 1820 405
rect 1814 400 1815 404
rect 1819 400 1820 404
rect 1814 399 1820 400
rect 1934 403 1940 404
rect 1934 399 1935 403
rect 1939 399 1940 403
rect 1976 401 1978 461
rect 110 398 116 399
rect 112 363 114 398
rect 184 363 186 399
rect 512 363 514 399
rect 840 363 842 399
rect 1168 363 1170 399
rect 1504 363 1506 399
rect 1816 363 1818 399
rect 1934 398 1940 399
rect 1974 400 1980 401
rect 1996 400 1998 461
rect 2204 400 2206 461
rect 2428 400 2430 461
rect 2652 400 2654 461
rect 2860 400 2862 461
rect 3068 400 3070 461
rect 3268 400 3270 461
rect 3468 400 3470 461
rect 3652 400 3654 461
rect 3800 401 3802 461
rect 3840 409 3842 469
rect 3838 408 3844 409
rect 4452 408 4454 469
rect 4644 408 4646 469
rect 4844 408 4846 469
rect 5052 408 5054 469
rect 5268 408 5270 469
rect 5484 408 5486 469
rect 5664 409 5666 469
rect 5662 408 5668 409
rect 3838 404 3839 408
rect 3843 404 3844 408
rect 3838 403 3844 404
rect 4450 407 4456 408
rect 4450 403 4451 407
rect 4455 403 4456 407
rect 4450 402 4456 403
rect 4642 407 4648 408
rect 4642 403 4643 407
rect 4647 403 4648 407
rect 4642 402 4648 403
rect 4842 407 4848 408
rect 4842 403 4843 407
rect 4847 403 4848 407
rect 4842 402 4848 403
rect 5050 407 5056 408
rect 5050 403 5051 407
rect 5055 403 5056 407
rect 5050 402 5056 403
rect 5266 407 5272 408
rect 5266 403 5267 407
rect 5271 403 5272 407
rect 5266 402 5272 403
rect 5482 407 5488 408
rect 5482 403 5483 407
rect 5487 403 5488 407
rect 5662 404 5663 408
rect 5667 404 5668 408
rect 5662 403 5668 404
rect 5482 402 5488 403
rect 3798 400 3804 401
rect 1936 363 1938 398
rect 1974 396 1975 400
rect 1979 396 1980 400
rect 1974 395 1980 396
rect 1994 399 2000 400
rect 1994 395 1995 399
rect 1999 395 2000 399
rect 1994 394 2000 395
rect 2202 399 2208 400
rect 2202 395 2203 399
rect 2207 395 2208 399
rect 2202 394 2208 395
rect 2426 399 2432 400
rect 2426 395 2427 399
rect 2431 395 2432 399
rect 2426 394 2432 395
rect 2650 399 2656 400
rect 2650 395 2651 399
rect 2655 395 2656 399
rect 2650 394 2656 395
rect 2858 399 2864 400
rect 2858 395 2859 399
rect 2863 395 2864 399
rect 2858 394 2864 395
rect 3066 399 3072 400
rect 3066 395 3067 399
rect 3071 395 3072 399
rect 3066 394 3072 395
rect 3266 399 3272 400
rect 3266 395 3267 399
rect 3271 395 3272 399
rect 3266 394 3272 395
rect 3466 399 3472 400
rect 3466 395 3467 399
rect 3471 395 3472 399
rect 3466 394 3472 395
rect 3650 399 3656 400
rect 3650 395 3651 399
rect 3655 395 3656 399
rect 3798 396 3799 400
rect 3803 396 3804 400
rect 3798 395 3804 396
rect 3650 394 3656 395
rect 4478 392 4484 393
rect 3838 391 3844 392
rect 3838 387 3839 391
rect 3843 387 3844 391
rect 4478 388 4479 392
rect 4483 388 4484 392
rect 4478 387 4484 388
rect 4670 392 4676 393
rect 4670 388 4671 392
rect 4675 388 4676 392
rect 4670 387 4676 388
rect 4870 392 4876 393
rect 4870 388 4871 392
rect 4875 388 4876 392
rect 4870 387 4876 388
rect 5078 392 5084 393
rect 5078 388 5079 392
rect 5083 388 5084 392
rect 5078 387 5084 388
rect 5294 392 5300 393
rect 5294 388 5295 392
rect 5299 388 5300 392
rect 5294 387 5300 388
rect 5510 392 5516 393
rect 5510 388 5511 392
rect 5515 388 5516 392
rect 5510 387 5516 388
rect 5662 391 5668 392
rect 5662 387 5663 391
rect 5667 387 5668 391
rect 3838 386 3844 387
rect 2022 384 2028 385
rect 1974 383 1980 384
rect 1974 379 1975 383
rect 1979 379 1980 383
rect 2022 380 2023 384
rect 2027 380 2028 384
rect 2022 379 2028 380
rect 2230 384 2236 385
rect 2230 380 2231 384
rect 2235 380 2236 384
rect 2230 379 2236 380
rect 2454 384 2460 385
rect 2454 380 2455 384
rect 2459 380 2460 384
rect 2454 379 2460 380
rect 2678 384 2684 385
rect 2678 380 2679 384
rect 2683 380 2684 384
rect 2678 379 2684 380
rect 2886 384 2892 385
rect 2886 380 2887 384
rect 2891 380 2892 384
rect 2886 379 2892 380
rect 3094 384 3100 385
rect 3094 380 3095 384
rect 3099 380 3100 384
rect 3094 379 3100 380
rect 3294 384 3300 385
rect 3294 380 3295 384
rect 3299 380 3300 384
rect 3294 379 3300 380
rect 3494 384 3500 385
rect 3494 380 3495 384
rect 3499 380 3500 384
rect 3494 379 3500 380
rect 3678 384 3684 385
rect 3678 380 3679 384
rect 3683 380 3684 384
rect 3678 379 3684 380
rect 3798 383 3804 384
rect 3798 379 3799 383
rect 3803 379 3804 383
rect 1974 378 1980 379
rect 111 362 115 363
rect 111 357 115 358
rect 183 362 187 363
rect 183 357 187 358
rect 279 362 283 363
rect 279 357 283 358
rect 487 362 491 363
rect 487 357 491 358
rect 511 362 515 363
rect 511 357 515 358
rect 703 362 707 363
rect 703 357 707 358
rect 839 362 843 363
rect 839 357 843 358
rect 919 362 923 363
rect 919 357 923 358
rect 1135 362 1139 363
rect 1135 357 1139 358
rect 1167 362 1171 363
rect 1167 357 1171 358
rect 1503 362 1507 363
rect 1503 357 1507 358
rect 1815 362 1819 363
rect 1815 357 1819 358
rect 1935 362 1939 363
rect 1935 357 1939 358
rect 112 334 114 357
rect 110 333 116 334
rect 280 333 282 357
rect 488 333 490 357
rect 704 333 706 357
rect 920 333 922 357
rect 1136 333 1138 357
rect 1936 334 1938 357
rect 1976 339 1978 378
rect 2024 339 2026 379
rect 2232 339 2234 379
rect 2456 339 2458 379
rect 2680 339 2682 379
rect 2888 339 2890 379
rect 3096 339 3098 379
rect 3296 339 3298 379
rect 3496 339 3498 379
rect 3680 339 3682 379
rect 3798 378 3804 379
rect 3800 339 3802 378
rect 3840 359 3842 386
rect 4480 359 4482 387
rect 4672 359 4674 387
rect 4872 359 4874 387
rect 5080 359 5082 387
rect 5296 359 5298 387
rect 5512 359 5514 387
rect 5662 386 5668 387
rect 5664 359 5666 386
rect 3839 358 3843 359
rect 3839 353 3843 354
rect 4479 358 4483 359
rect 4479 353 4483 354
rect 4615 358 4619 359
rect 4615 353 4619 354
rect 4671 358 4675 359
rect 4671 353 4675 354
rect 4775 358 4779 359
rect 4775 353 4779 354
rect 4871 358 4875 359
rect 4871 353 4875 354
rect 4951 358 4955 359
rect 4951 353 4955 354
rect 5079 358 5083 359
rect 5079 353 5083 354
rect 5135 358 5139 359
rect 5135 353 5139 354
rect 5295 358 5299 359
rect 5295 353 5299 354
rect 5327 358 5331 359
rect 5327 353 5331 354
rect 5511 358 5515 359
rect 5511 353 5515 354
rect 5527 358 5531 359
rect 5527 353 5531 354
rect 5663 358 5667 359
rect 5663 353 5667 354
rect 1975 338 1979 339
rect 1934 333 1940 334
rect 1975 333 1979 334
rect 2023 338 2027 339
rect 2023 333 2027 334
rect 2159 338 2163 339
rect 2159 333 2163 334
rect 2231 338 2235 339
rect 2231 333 2235 334
rect 2295 338 2299 339
rect 2295 333 2299 334
rect 2431 338 2435 339
rect 2431 333 2435 334
rect 2455 338 2459 339
rect 2455 333 2459 334
rect 2567 338 2571 339
rect 2567 333 2571 334
rect 2679 338 2683 339
rect 2679 333 2683 334
rect 2703 338 2707 339
rect 2703 333 2707 334
rect 2839 338 2843 339
rect 2839 333 2843 334
rect 2887 338 2891 339
rect 2887 333 2891 334
rect 2975 338 2979 339
rect 2975 333 2979 334
rect 3095 338 3099 339
rect 3095 333 3099 334
rect 3111 338 3115 339
rect 3111 333 3115 334
rect 3247 338 3251 339
rect 3247 333 3251 334
rect 3295 338 3299 339
rect 3295 333 3299 334
rect 3383 338 3387 339
rect 3383 333 3387 334
rect 3495 338 3499 339
rect 3495 333 3499 334
rect 3519 338 3523 339
rect 3519 333 3523 334
rect 3655 338 3659 339
rect 3655 333 3659 334
rect 3679 338 3683 339
rect 3679 333 3683 334
rect 3799 338 3803 339
rect 3799 333 3803 334
rect 110 329 111 333
rect 115 329 116 333
rect 110 328 116 329
rect 278 332 284 333
rect 278 328 279 332
rect 283 328 284 332
rect 278 327 284 328
rect 486 332 492 333
rect 486 328 487 332
rect 491 328 492 332
rect 486 327 492 328
rect 702 332 708 333
rect 702 328 703 332
rect 707 328 708 332
rect 702 327 708 328
rect 918 332 924 333
rect 918 328 919 332
rect 923 328 924 332
rect 918 327 924 328
rect 1134 332 1140 333
rect 1134 328 1135 332
rect 1139 328 1140 332
rect 1934 329 1935 333
rect 1939 329 1940 333
rect 1934 328 1940 329
rect 1134 327 1140 328
rect 250 317 256 318
rect 110 316 116 317
rect 110 312 111 316
rect 115 312 116 316
rect 250 313 251 317
rect 255 313 256 317
rect 250 312 256 313
rect 458 317 464 318
rect 458 313 459 317
rect 463 313 464 317
rect 458 312 464 313
rect 674 317 680 318
rect 674 313 675 317
rect 679 313 680 317
rect 674 312 680 313
rect 890 317 896 318
rect 890 313 891 317
rect 895 313 896 317
rect 890 312 896 313
rect 1106 317 1112 318
rect 1106 313 1107 317
rect 1111 313 1112 317
rect 1106 312 1112 313
rect 1934 316 1940 317
rect 1934 312 1935 316
rect 1939 312 1940 316
rect 110 311 116 312
rect 112 211 114 311
rect 252 211 254 312
rect 460 211 462 312
rect 676 211 678 312
rect 892 211 894 312
rect 1108 211 1110 312
rect 1934 311 1940 312
rect 1936 211 1938 311
rect 1976 310 1978 333
rect 1974 309 1980 310
rect 2024 309 2026 333
rect 2160 309 2162 333
rect 2296 309 2298 333
rect 2432 309 2434 333
rect 2568 309 2570 333
rect 2704 309 2706 333
rect 2840 309 2842 333
rect 2976 309 2978 333
rect 3112 309 3114 333
rect 3248 309 3250 333
rect 3384 309 3386 333
rect 3520 309 3522 333
rect 3656 309 3658 333
rect 3800 310 3802 333
rect 3840 330 3842 353
rect 3838 329 3844 330
rect 4616 329 4618 353
rect 4776 329 4778 353
rect 4952 329 4954 353
rect 5136 329 5138 353
rect 5328 329 5330 353
rect 5528 329 5530 353
rect 5664 330 5666 353
rect 5662 329 5668 330
rect 3838 325 3839 329
rect 3843 325 3844 329
rect 3838 324 3844 325
rect 4614 328 4620 329
rect 4614 324 4615 328
rect 4619 324 4620 328
rect 4614 323 4620 324
rect 4774 328 4780 329
rect 4774 324 4775 328
rect 4779 324 4780 328
rect 4774 323 4780 324
rect 4950 328 4956 329
rect 4950 324 4951 328
rect 4955 324 4956 328
rect 4950 323 4956 324
rect 5134 328 5140 329
rect 5134 324 5135 328
rect 5139 324 5140 328
rect 5134 323 5140 324
rect 5326 328 5332 329
rect 5326 324 5327 328
rect 5331 324 5332 328
rect 5326 323 5332 324
rect 5526 328 5532 329
rect 5526 324 5527 328
rect 5531 324 5532 328
rect 5662 325 5663 329
rect 5667 325 5668 329
rect 5662 324 5668 325
rect 5526 323 5532 324
rect 4586 313 4592 314
rect 3838 312 3844 313
rect 3798 309 3804 310
rect 1974 305 1975 309
rect 1979 305 1980 309
rect 1974 304 1980 305
rect 2022 308 2028 309
rect 2022 304 2023 308
rect 2027 304 2028 308
rect 2022 303 2028 304
rect 2158 308 2164 309
rect 2158 304 2159 308
rect 2163 304 2164 308
rect 2158 303 2164 304
rect 2294 308 2300 309
rect 2294 304 2295 308
rect 2299 304 2300 308
rect 2294 303 2300 304
rect 2430 308 2436 309
rect 2430 304 2431 308
rect 2435 304 2436 308
rect 2430 303 2436 304
rect 2566 308 2572 309
rect 2566 304 2567 308
rect 2571 304 2572 308
rect 2566 303 2572 304
rect 2702 308 2708 309
rect 2702 304 2703 308
rect 2707 304 2708 308
rect 2702 303 2708 304
rect 2838 308 2844 309
rect 2838 304 2839 308
rect 2843 304 2844 308
rect 2838 303 2844 304
rect 2974 308 2980 309
rect 2974 304 2975 308
rect 2979 304 2980 308
rect 2974 303 2980 304
rect 3110 308 3116 309
rect 3110 304 3111 308
rect 3115 304 3116 308
rect 3110 303 3116 304
rect 3246 308 3252 309
rect 3246 304 3247 308
rect 3251 304 3252 308
rect 3246 303 3252 304
rect 3382 308 3388 309
rect 3382 304 3383 308
rect 3387 304 3388 308
rect 3382 303 3388 304
rect 3518 308 3524 309
rect 3518 304 3519 308
rect 3523 304 3524 308
rect 3518 303 3524 304
rect 3654 308 3660 309
rect 3654 304 3655 308
rect 3659 304 3660 308
rect 3798 305 3799 309
rect 3803 305 3804 309
rect 3838 308 3839 312
rect 3843 308 3844 312
rect 4586 309 4587 313
rect 4591 309 4592 313
rect 4586 308 4592 309
rect 4746 313 4752 314
rect 4746 309 4747 313
rect 4751 309 4752 313
rect 4746 308 4752 309
rect 4922 313 4928 314
rect 4922 309 4923 313
rect 4927 309 4928 313
rect 4922 308 4928 309
rect 5106 313 5112 314
rect 5106 309 5107 313
rect 5111 309 5112 313
rect 5106 308 5112 309
rect 5298 313 5304 314
rect 5298 309 5299 313
rect 5303 309 5304 313
rect 5298 308 5304 309
rect 5498 313 5504 314
rect 5498 309 5499 313
rect 5503 309 5504 313
rect 5498 308 5504 309
rect 5662 312 5668 313
rect 5662 308 5663 312
rect 5667 308 5668 312
rect 3838 307 3844 308
rect 3798 304 3804 305
rect 3654 303 3660 304
rect 1994 293 2000 294
rect 1974 292 1980 293
rect 1974 288 1975 292
rect 1979 288 1980 292
rect 1994 289 1995 293
rect 1999 289 2000 293
rect 1994 288 2000 289
rect 2130 293 2136 294
rect 2130 289 2131 293
rect 2135 289 2136 293
rect 2130 288 2136 289
rect 2266 293 2272 294
rect 2266 289 2267 293
rect 2271 289 2272 293
rect 2266 288 2272 289
rect 2402 293 2408 294
rect 2402 289 2403 293
rect 2407 289 2408 293
rect 2402 288 2408 289
rect 2538 293 2544 294
rect 2538 289 2539 293
rect 2543 289 2544 293
rect 2538 288 2544 289
rect 2674 293 2680 294
rect 2674 289 2675 293
rect 2679 289 2680 293
rect 2674 288 2680 289
rect 2810 293 2816 294
rect 2810 289 2811 293
rect 2815 289 2816 293
rect 2810 288 2816 289
rect 2946 293 2952 294
rect 2946 289 2947 293
rect 2951 289 2952 293
rect 2946 288 2952 289
rect 3082 293 3088 294
rect 3082 289 3083 293
rect 3087 289 3088 293
rect 3082 288 3088 289
rect 3218 293 3224 294
rect 3218 289 3219 293
rect 3223 289 3224 293
rect 3218 288 3224 289
rect 3354 293 3360 294
rect 3354 289 3355 293
rect 3359 289 3360 293
rect 3354 288 3360 289
rect 3490 293 3496 294
rect 3490 289 3491 293
rect 3495 289 3496 293
rect 3490 288 3496 289
rect 3626 293 3632 294
rect 3626 289 3627 293
rect 3631 289 3632 293
rect 3626 288 3632 289
rect 3798 292 3804 293
rect 3798 288 3799 292
rect 3803 288 3804 292
rect 1974 287 1980 288
rect 111 210 115 211
rect 111 205 115 206
rect 131 210 135 211
rect 131 205 135 206
rect 251 210 255 211
rect 251 205 255 206
rect 267 210 271 211
rect 267 205 271 206
rect 403 210 407 211
rect 403 205 407 206
rect 459 210 463 211
rect 459 205 463 206
rect 539 210 543 211
rect 539 205 543 206
rect 675 210 679 211
rect 675 205 679 206
rect 811 210 815 211
rect 811 205 815 206
rect 891 210 895 211
rect 891 205 895 206
rect 947 210 951 211
rect 947 205 951 206
rect 1083 210 1087 211
rect 1083 205 1087 206
rect 1107 210 1111 211
rect 1107 205 1111 206
rect 1935 210 1939 211
rect 1935 205 1939 206
rect 112 145 114 205
rect 110 144 116 145
rect 132 144 134 205
rect 268 144 270 205
rect 404 144 406 205
rect 540 144 542 205
rect 676 144 678 205
rect 812 144 814 205
rect 948 144 950 205
rect 1084 144 1086 205
rect 1936 145 1938 205
rect 1976 191 1978 287
rect 1996 191 1998 288
rect 2132 191 2134 288
rect 2268 191 2270 288
rect 2404 191 2406 288
rect 2540 191 2542 288
rect 2676 191 2678 288
rect 2812 191 2814 288
rect 2948 191 2950 288
rect 3084 191 3086 288
rect 3220 191 3222 288
rect 3356 191 3358 288
rect 3492 191 3494 288
rect 3628 191 3630 288
rect 3798 287 3804 288
rect 3800 191 3802 287
rect 3840 207 3842 307
rect 4588 207 4590 308
rect 4748 207 4750 308
rect 4924 207 4926 308
rect 5108 207 5110 308
rect 5300 207 5302 308
rect 5500 207 5502 308
rect 5662 307 5668 308
rect 5664 207 5666 307
rect 3839 206 3843 207
rect 3839 201 3843 202
rect 4291 206 4295 207
rect 4291 201 4295 202
rect 4427 206 4431 207
rect 4427 201 4431 202
rect 4563 206 4567 207
rect 4563 201 4567 202
rect 4587 206 4591 207
rect 4587 201 4591 202
rect 4699 206 4703 207
rect 4699 201 4703 202
rect 4747 206 4751 207
rect 4747 201 4751 202
rect 4835 206 4839 207
rect 4835 201 4839 202
rect 4923 206 4927 207
rect 4923 201 4927 202
rect 4971 206 4975 207
rect 4971 201 4975 202
rect 5107 206 5111 207
rect 5107 201 5111 202
rect 5243 206 5247 207
rect 5243 201 5247 202
rect 5299 206 5303 207
rect 5299 201 5303 202
rect 5379 206 5383 207
rect 5379 201 5383 202
rect 5499 206 5503 207
rect 5499 201 5503 202
rect 5515 206 5519 207
rect 5515 201 5519 202
rect 5663 206 5667 207
rect 5663 201 5667 202
rect 1975 190 1979 191
rect 1975 185 1979 186
rect 1995 190 1999 191
rect 1995 185 1999 186
rect 2131 190 2135 191
rect 2131 185 2135 186
rect 2267 190 2271 191
rect 2267 185 2271 186
rect 2403 190 2407 191
rect 2403 185 2407 186
rect 2539 190 2543 191
rect 2539 185 2543 186
rect 2675 190 2679 191
rect 2675 185 2679 186
rect 2811 190 2815 191
rect 2811 185 2815 186
rect 2947 190 2951 191
rect 2947 185 2951 186
rect 3083 190 3087 191
rect 3083 185 3087 186
rect 3219 190 3223 191
rect 3219 185 3223 186
rect 3355 190 3359 191
rect 3355 185 3359 186
rect 3491 190 3495 191
rect 3491 185 3495 186
rect 3627 190 3631 191
rect 3627 185 3631 186
rect 3799 190 3803 191
rect 3799 185 3803 186
rect 1934 144 1940 145
rect 110 140 111 144
rect 115 140 116 144
rect 110 139 116 140
rect 130 143 136 144
rect 130 139 131 143
rect 135 139 136 143
rect 130 138 136 139
rect 266 143 272 144
rect 266 139 267 143
rect 271 139 272 143
rect 266 138 272 139
rect 402 143 408 144
rect 402 139 403 143
rect 407 139 408 143
rect 402 138 408 139
rect 538 143 544 144
rect 538 139 539 143
rect 543 139 544 143
rect 538 138 544 139
rect 674 143 680 144
rect 674 139 675 143
rect 679 139 680 143
rect 674 138 680 139
rect 810 143 816 144
rect 810 139 811 143
rect 815 139 816 143
rect 810 138 816 139
rect 946 143 952 144
rect 946 139 947 143
rect 951 139 952 143
rect 946 138 952 139
rect 1082 143 1088 144
rect 1082 139 1083 143
rect 1087 139 1088 143
rect 1934 140 1935 144
rect 1939 140 1940 144
rect 1934 139 1940 140
rect 1082 138 1088 139
rect 158 128 164 129
rect 110 127 116 128
rect 110 123 111 127
rect 115 123 116 127
rect 158 124 159 128
rect 163 124 164 128
rect 158 123 164 124
rect 294 128 300 129
rect 294 124 295 128
rect 299 124 300 128
rect 294 123 300 124
rect 430 128 436 129
rect 430 124 431 128
rect 435 124 436 128
rect 430 123 436 124
rect 566 128 572 129
rect 566 124 567 128
rect 571 124 572 128
rect 566 123 572 124
rect 702 128 708 129
rect 702 124 703 128
rect 707 124 708 128
rect 702 123 708 124
rect 838 128 844 129
rect 838 124 839 128
rect 843 124 844 128
rect 838 123 844 124
rect 974 128 980 129
rect 974 124 975 128
rect 979 124 980 128
rect 974 123 980 124
rect 1110 128 1116 129
rect 1110 124 1111 128
rect 1115 124 1116 128
rect 1110 123 1116 124
rect 1934 127 1940 128
rect 1934 123 1935 127
rect 1939 123 1940 127
rect 1976 125 1978 185
rect 110 122 116 123
rect 112 99 114 122
rect 160 99 162 123
rect 296 99 298 123
rect 432 99 434 123
rect 568 99 570 123
rect 704 99 706 123
rect 840 99 842 123
rect 976 99 978 123
rect 1112 99 1114 123
rect 1934 122 1940 123
rect 1974 124 1980 125
rect 1996 124 1998 185
rect 2132 124 2134 185
rect 2268 124 2270 185
rect 2404 124 2406 185
rect 2540 124 2542 185
rect 2676 124 2678 185
rect 2812 124 2814 185
rect 2948 124 2950 185
rect 3084 124 3086 185
rect 3220 124 3222 185
rect 3356 124 3358 185
rect 3492 124 3494 185
rect 3628 124 3630 185
rect 3800 125 3802 185
rect 3840 141 3842 201
rect 3838 140 3844 141
rect 4292 140 4294 201
rect 4428 140 4430 201
rect 4564 140 4566 201
rect 4700 140 4702 201
rect 4836 140 4838 201
rect 4972 140 4974 201
rect 5108 140 5110 201
rect 5244 140 5246 201
rect 5380 140 5382 201
rect 5516 140 5518 201
rect 5664 141 5666 201
rect 5662 140 5668 141
rect 3838 136 3839 140
rect 3843 136 3844 140
rect 3838 135 3844 136
rect 4290 139 4296 140
rect 4290 135 4291 139
rect 4295 135 4296 139
rect 4290 134 4296 135
rect 4426 139 4432 140
rect 4426 135 4427 139
rect 4431 135 4432 139
rect 4426 134 4432 135
rect 4562 139 4568 140
rect 4562 135 4563 139
rect 4567 135 4568 139
rect 4562 134 4568 135
rect 4698 139 4704 140
rect 4698 135 4699 139
rect 4703 135 4704 139
rect 4698 134 4704 135
rect 4834 139 4840 140
rect 4834 135 4835 139
rect 4839 135 4840 139
rect 4834 134 4840 135
rect 4970 139 4976 140
rect 4970 135 4971 139
rect 4975 135 4976 139
rect 4970 134 4976 135
rect 5106 139 5112 140
rect 5106 135 5107 139
rect 5111 135 5112 139
rect 5106 134 5112 135
rect 5242 139 5248 140
rect 5242 135 5243 139
rect 5247 135 5248 139
rect 5242 134 5248 135
rect 5378 139 5384 140
rect 5378 135 5379 139
rect 5383 135 5384 139
rect 5378 134 5384 135
rect 5514 139 5520 140
rect 5514 135 5515 139
rect 5519 135 5520 139
rect 5662 136 5663 140
rect 5667 136 5668 140
rect 5662 135 5668 136
rect 5514 134 5520 135
rect 3798 124 3804 125
rect 4318 124 4324 125
rect 1936 99 1938 122
rect 1974 120 1975 124
rect 1979 120 1980 124
rect 1974 119 1980 120
rect 1994 123 2000 124
rect 1994 119 1995 123
rect 1999 119 2000 123
rect 1994 118 2000 119
rect 2130 123 2136 124
rect 2130 119 2131 123
rect 2135 119 2136 123
rect 2130 118 2136 119
rect 2266 123 2272 124
rect 2266 119 2267 123
rect 2271 119 2272 123
rect 2266 118 2272 119
rect 2402 123 2408 124
rect 2402 119 2403 123
rect 2407 119 2408 123
rect 2402 118 2408 119
rect 2538 123 2544 124
rect 2538 119 2539 123
rect 2543 119 2544 123
rect 2538 118 2544 119
rect 2674 123 2680 124
rect 2674 119 2675 123
rect 2679 119 2680 123
rect 2674 118 2680 119
rect 2810 123 2816 124
rect 2810 119 2811 123
rect 2815 119 2816 123
rect 2810 118 2816 119
rect 2946 123 2952 124
rect 2946 119 2947 123
rect 2951 119 2952 123
rect 2946 118 2952 119
rect 3082 123 3088 124
rect 3082 119 3083 123
rect 3087 119 3088 123
rect 3082 118 3088 119
rect 3218 123 3224 124
rect 3218 119 3219 123
rect 3223 119 3224 123
rect 3218 118 3224 119
rect 3354 123 3360 124
rect 3354 119 3355 123
rect 3359 119 3360 123
rect 3354 118 3360 119
rect 3490 123 3496 124
rect 3490 119 3491 123
rect 3495 119 3496 123
rect 3490 118 3496 119
rect 3626 123 3632 124
rect 3626 119 3627 123
rect 3631 119 3632 123
rect 3798 120 3799 124
rect 3803 120 3804 124
rect 3798 119 3804 120
rect 3838 123 3844 124
rect 3838 119 3839 123
rect 3843 119 3844 123
rect 4318 120 4319 124
rect 4323 120 4324 124
rect 4318 119 4324 120
rect 4454 124 4460 125
rect 4454 120 4455 124
rect 4459 120 4460 124
rect 4454 119 4460 120
rect 4590 124 4596 125
rect 4590 120 4591 124
rect 4595 120 4596 124
rect 4590 119 4596 120
rect 4726 124 4732 125
rect 4726 120 4727 124
rect 4731 120 4732 124
rect 4726 119 4732 120
rect 4862 124 4868 125
rect 4862 120 4863 124
rect 4867 120 4868 124
rect 4862 119 4868 120
rect 4998 124 5004 125
rect 4998 120 4999 124
rect 5003 120 5004 124
rect 4998 119 5004 120
rect 5134 124 5140 125
rect 5134 120 5135 124
rect 5139 120 5140 124
rect 5134 119 5140 120
rect 5270 124 5276 125
rect 5270 120 5271 124
rect 5275 120 5276 124
rect 5270 119 5276 120
rect 5406 124 5412 125
rect 5406 120 5407 124
rect 5411 120 5412 124
rect 5406 119 5412 120
rect 5542 124 5548 125
rect 5542 120 5543 124
rect 5547 120 5548 124
rect 5542 119 5548 120
rect 5662 123 5668 124
rect 5662 119 5663 123
rect 5667 119 5668 123
rect 3626 118 3632 119
rect 3838 118 3844 119
rect 2022 108 2028 109
rect 1974 107 1980 108
rect 1974 103 1975 107
rect 1979 103 1980 107
rect 2022 104 2023 108
rect 2027 104 2028 108
rect 2022 103 2028 104
rect 2158 108 2164 109
rect 2158 104 2159 108
rect 2163 104 2164 108
rect 2158 103 2164 104
rect 2294 108 2300 109
rect 2294 104 2295 108
rect 2299 104 2300 108
rect 2294 103 2300 104
rect 2430 108 2436 109
rect 2430 104 2431 108
rect 2435 104 2436 108
rect 2430 103 2436 104
rect 2566 108 2572 109
rect 2566 104 2567 108
rect 2571 104 2572 108
rect 2566 103 2572 104
rect 2702 108 2708 109
rect 2702 104 2703 108
rect 2707 104 2708 108
rect 2702 103 2708 104
rect 2838 108 2844 109
rect 2838 104 2839 108
rect 2843 104 2844 108
rect 2838 103 2844 104
rect 2974 108 2980 109
rect 2974 104 2975 108
rect 2979 104 2980 108
rect 2974 103 2980 104
rect 3110 108 3116 109
rect 3110 104 3111 108
rect 3115 104 3116 108
rect 3110 103 3116 104
rect 3246 108 3252 109
rect 3246 104 3247 108
rect 3251 104 3252 108
rect 3246 103 3252 104
rect 3382 108 3388 109
rect 3382 104 3383 108
rect 3387 104 3388 108
rect 3382 103 3388 104
rect 3518 108 3524 109
rect 3518 104 3519 108
rect 3523 104 3524 108
rect 3518 103 3524 104
rect 3654 108 3660 109
rect 3654 104 3655 108
rect 3659 104 3660 108
rect 3654 103 3660 104
rect 3798 107 3804 108
rect 3798 103 3799 107
rect 3803 103 3804 107
rect 1974 102 1980 103
rect 111 98 115 99
rect 111 93 115 94
rect 159 98 163 99
rect 159 93 163 94
rect 295 98 299 99
rect 295 93 299 94
rect 431 98 435 99
rect 431 93 435 94
rect 567 98 571 99
rect 567 93 571 94
rect 703 98 707 99
rect 703 93 707 94
rect 839 98 843 99
rect 839 93 843 94
rect 975 98 979 99
rect 975 93 979 94
rect 1111 98 1115 99
rect 1111 93 1115 94
rect 1935 98 1939 99
rect 1935 93 1939 94
rect 1976 79 1978 102
rect 2024 79 2026 103
rect 2160 79 2162 103
rect 2296 79 2298 103
rect 2432 79 2434 103
rect 2568 79 2570 103
rect 2704 79 2706 103
rect 2840 79 2842 103
rect 2976 79 2978 103
rect 3112 79 3114 103
rect 3248 79 3250 103
rect 3384 79 3386 103
rect 3520 79 3522 103
rect 3656 79 3658 103
rect 3798 102 3804 103
rect 3800 79 3802 102
rect 3840 95 3842 118
rect 4320 95 4322 119
rect 4456 95 4458 119
rect 4592 95 4594 119
rect 4728 95 4730 119
rect 4864 95 4866 119
rect 5000 95 5002 119
rect 5136 95 5138 119
rect 5272 95 5274 119
rect 5408 95 5410 119
rect 5544 95 5546 119
rect 5662 118 5668 119
rect 5664 95 5666 118
rect 3839 94 3843 95
rect 3839 89 3843 90
rect 4319 94 4323 95
rect 4319 89 4323 90
rect 4455 94 4459 95
rect 4455 89 4459 90
rect 4591 94 4595 95
rect 4591 89 4595 90
rect 4727 94 4731 95
rect 4727 89 4731 90
rect 4863 94 4867 95
rect 4863 89 4867 90
rect 4999 94 5003 95
rect 4999 89 5003 90
rect 5135 94 5139 95
rect 5135 89 5139 90
rect 5271 94 5275 95
rect 5271 89 5275 90
rect 5407 94 5411 95
rect 5407 89 5411 90
rect 5543 94 5547 95
rect 5543 89 5547 90
rect 5663 94 5667 95
rect 5663 89 5667 90
rect 1975 78 1979 79
rect 1975 73 1979 74
rect 2023 78 2027 79
rect 2023 73 2027 74
rect 2159 78 2163 79
rect 2159 73 2163 74
rect 2295 78 2299 79
rect 2295 73 2299 74
rect 2431 78 2435 79
rect 2431 73 2435 74
rect 2567 78 2571 79
rect 2567 73 2571 74
rect 2703 78 2707 79
rect 2703 73 2707 74
rect 2839 78 2843 79
rect 2839 73 2843 74
rect 2975 78 2979 79
rect 2975 73 2979 74
rect 3111 78 3115 79
rect 3111 73 3115 74
rect 3247 78 3251 79
rect 3247 73 3251 74
rect 3383 78 3387 79
rect 3383 73 3387 74
rect 3519 78 3523 79
rect 3519 73 3523 74
rect 3655 78 3659 79
rect 3655 73 3659 74
rect 3799 78 3803 79
rect 3799 73 3803 74
<< m4c >>
rect 111 5754 115 5758
rect 159 5754 163 5758
rect 295 5754 299 5758
rect 1935 5754 1939 5758
rect 1975 5654 1979 5658
rect 2023 5654 2027 5658
rect 2183 5654 2187 5658
rect 2367 5654 2371 5658
rect 2551 5654 2555 5658
rect 2727 5654 2731 5658
rect 2895 5654 2899 5658
rect 3063 5654 3067 5658
rect 3223 5654 3227 5658
rect 3383 5654 3387 5658
rect 3543 5654 3547 5658
rect 3679 5654 3683 5658
rect 3799 5654 3803 5658
rect 111 5642 115 5646
rect 131 5642 135 5646
rect 267 5642 271 5646
rect 275 5642 279 5646
rect 475 5642 479 5646
rect 699 5642 703 5646
rect 955 5642 959 5646
rect 1227 5642 1231 5646
rect 1515 5642 1519 5646
rect 1787 5642 1791 5646
rect 1935 5642 1939 5646
rect 3839 5650 3843 5654
rect 4335 5650 4339 5654
rect 4471 5650 4475 5654
rect 4607 5650 4611 5654
rect 4743 5650 4747 5654
rect 4879 5650 4883 5654
rect 5015 5650 5019 5654
rect 5663 5650 5667 5654
rect 1975 5542 1979 5546
rect 1995 5542 1999 5546
rect 2139 5542 2143 5546
rect 2155 5542 2159 5546
rect 2339 5542 2343 5546
rect 2355 5542 2359 5546
rect 2523 5542 2527 5546
rect 2563 5542 2567 5546
rect 2699 5542 2703 5546
rect 2755 5542 2759 5546
rect 2867 5542 2871 5546
rect 2939 5542 2943 5546
rect 3035 5542 3039 5546
rect 3115 5542 3119 5546
rect 3195 5542 3199 5546
rect 3291 5542 3295 5546
rect 3355 5542 3359 5546
rect 3467 5542 3471 5546
rect 3515 5542 3519 5546
rect 3643 5542 3647 5546
rect 3651 5542 3655 5546
rect 3799 5542 3803 5546
rect 111 5530 115 5534
rect 159 5530 163 5534
rect 279 5530 283 5534
rect 303 5530 307 5534
rect 503 5530 507 5534
rect 519 5530 523 5534
rect 727 5530 731 5534
rect 767 5530 771 5534
rect 983 5530 987 5534
rect 1015 5530 1019 5534
rect 1255 5530 1259 5534
rect 1263 5530 1267 5534
rect 1511 5530 1515 5534
rect 1543 5530 1547 5534
rect 1767 5530 1771 5534
rect 1815 5530 1819 5534
rect 1935 5530 1939 5534
rect 3839 5538 3843 5542
rect 4251 5538 4255 5542
rect 4307 5538 4311 5542
rect 4403 5538 4407 5542
rect 4443 5538 4447 5542
rect 4555 5538 4559 5542
rect 4579 5538 4583 5542
rect 4707 5538 4711 5542
rect 4715 5538 4719 5542
rect 4851 5538 4855 5542
rect 4859 5538 4863 5542
rect 4987 5538 4991 5542
rect 5019 5538 5023 5542
rect 5663 5538 5667 5542
rect 111 5418 115 5422
rect 251 5418 255 5422
rect 411 5418 415 5422
rect 491 5418 495 5422
rect 611 5418 615 5422
rect 739 5418 743 5422
rect 819 5418 823 5422
rect 987 5418 991 5422
rect 1035 5418 1039 5422
rect 1235 5418 1239 5422
rect 1259 5418 1263 5422
rect 1483 5418 1487 5422
rect 1491 5418 1495 5422
rect 1739 5418 1743 5422
rect 1935 5418 1939 5422
rect 1975 5422 1979 5426
rect 2167 5422 2171 5426
rect 2311 5422 2315 5426
rect 2383 5422 2387 5426
rect 2511 5422 2515 5426
rect 2591 5422 2595 5426
rect 2703 5422 2707 5426
rect 2783 5422 2787 5426
rect 2887 5422 2891 5426
rect 2967 5422 2971 5426
rect 3071 5422 3075 5426
rect 3143 5422 3147 5426
rect 3247 5422 3251 5426
rect 3319 5422 3323 5426
rect 3423 5422 3427 5426
rect 3495 5422 3499 5426
rect 3607 5422 3611 5426
rect 3671 5422 3675 5426
rect 3799 5422 3803 5426
rect 3839 5406 3843 5410
rect 4279 5406 4283 5410
rect 4431 5406 4435 5410
rect 4487 5406 4491 5410
rect 4583 5406 4587 5410
rect 4695 5406 4699 5410
rect 4735 5406 4739 5410
rect 4887 5406 4891 5410
rect 4911 5406 4915 5410
rect 5047 5406 5051 5410
rect 5127 5406 5131 5410
rect 5663 5406 5667 5410
rect 111 5306 115 5310
rect 439 5306 443 5310
rect 591 5306 595 5310
rect 639 5306 643 5310
rect 727 5306 731 5310
rect 847 5306 851 5310
rect 863 5306 867 5310
rect 999 5306 1003 5310
rect 1063 5306 1067 5310
rect 1135 5306 1139 5310
rect 1271 5306 1275 5310
rect 1287 5306 1291 5310
rect 1407 5306 1411 5310
rect 1519 5306 1523 5310
rect 1543 5306 1547 5310
rect 1935 5306 1939 5310
rect 1975 5310 1979 5314
rect 2195 5310 2199 5314
rect 2283 5310 2287 5314
rect 2339 5310 2343 5314
rect 2483 5310 2487 5314
rect 2491 5310 2495 5314
rect 2651 5310 2655 5314
rect 2675 5310 2679 5314
rect 2819 5310 2823 5314
rect 2859 5310 2863 5314
rect 3003 5310 3007 5314
rect 3043 5310 3047 5314
rect 3187 5310 3191 5314
rect 3219 5310 3223 5314
rect 3379 5310 3383 5314
rect 3395 5310 3399 5314
rect 3579 5310 3583 5314
rect 3799 5310 3803 5314
rect 3839 5278 3843 5282
rect 4251 5278 4255 5282
rect 4459 5278 4463 5282
rect 4483 5278 4487 5282
rect 4667 5278 4671 5282
rect 4715 5278 4719 5282
rect 4883 5278 4887 5282
rect 4947 5278 4951 5282
rect 5099 5278 5103 5282
rect 5187 5278 5191 5282
rect 5663 5278 5667 5282
rect 1975 5198 1979 5202
rect 2023 5198 2027 5202
rect 2159 5198 2163 5202
rect 2223 5198 2227 5202
rect 2327 5198 2331 5202
rect 2367 5198 2371 5202
rect 2511 5198 2515 5202
rect 2519 5198 2523 5202
rect 2679 5198 2683 5202
rect 2695 5198 2699 5202
rect 2847 5198 2851 5202
rect 2887 5198 2891 5202
rect 3031 5198 3035 5202
rect 3087 5198 3091 5202
rect 3215 5198 3219 5202
rect 3287 5198 3291 5202
rect 3407 5198 3411 5202
rect 3495 5198 3499 5202
rect 3607 5198 3611 5202
rect 3679 5198 3683 5202
rect 3799 5198 3803 5202
rect 111 5090 115 5094
rect 347 5090 351 5094
rect 483 5090 487 5094
rect 563 5090 567 5094
rect 619 5090 623 5094
rect 699 5090 703 5094
rect 755 5090 759 5094
rect 835 5090 839 5094
rect 891 5090 895 5094
rect 971 5090 975 5094
rect 1035 5090 1039 5094
rect 1107 5090 1111 5094
rect 1187 5090 1191 5094
rect 1243 5090 1247 5094
rect 1339 5090 1343 5094
rect 1379 5090 1383 5094
rect 1491 5090 1495 5094
rect 1515 5090 1519 5094
rect 1651 5090 1655 5094
rect 1787 5090 1791 5094
rect 1935 5090 1939 5094
rect 3839 5138 3843 5142
rect 3887 5138 3891 5142
rect 4135 5138 4139 5142
rect 4279 5138 4283 5142
rect 4407 5138 4411 5142
rect 4511 5138 4515 5142
rect 4679 5138 4683 5142
rect 4743 5138 4747 5142
rect 4959 5138 4963 5142
rect 4975 5138 4979 5142
rect 5215 5138 5219 5142
rect 5239 5138 5243 5142
rect 5663 5138 5667 5142
rect 1975 5086 1979 5090
rect 1995 5086 1999 5090
rect 2131 5086 2135 5090
rect 2299 5086 2303 5090
rect 2483 5086 2487 5090
rect 2531 5086 2535 5090
rect 2667 5086 2671 5090
rect 2859 5086 2863 5090
rect 3059 5086 3063 5090
rect 3099 5086 3103 5090
rect 3259 5086 3263 5090
rect 3467 5086 3471 5090
rect 3651 5086 3655 5090
rect 3799 5086 3803 5090
rect 3839 5014 3843 5018
rect 3859 5014 3863 5018
rect 4019 5014 4023 5018
rect 4107 5014 4111 5018
rect 4211 5014 4215 5018
rect 4379 5014 4383 5018
rect 4411 5014 4415 5018
rect 4627 5014 4631 5018
rect 4651 5014 4655 5018
rect 4843 5014 4847 5018
rect 4931 5014 4935 5018
rect 5067 5014 5071 5018
rect 5211 5014 5215 5018
rect 5299 5014 5303 5018
rect 5663 5014 5667 5018
rect 111 4978 115 4982
rect 159 4978 163 4982
rect 343 4978 347 4982
rect 375 4978 379 4982
rect 511 4978 515 4982
rect 551 4978 555 4982
rect 647 4978 651 4982
rect 751 4978 755 4982
rect 783 4978 787 4982
rect 919 4978 923 4982
rect 943 4978 947 4982
rect 1063 4978 1067 4982
rect 1127 4978 1131 4982
rect 1215 4978 1219 4982
rect 1311 4978 1315 4982
rect 1367 4978 1371 4982
rect 1487 4978 1491 4982
rect 1519 4978 1523 4982
rect 1663 4978 1667 4982
rect 1679 4978 1683 4982
rect 1815 4978 1819 4982
rect 1935 4978 1939 4982
rect 1975 4942 1979 4946
rect 2023 4942 2027 4946
rect 2559 4942 2563 4946
rect 2871 4942 2875 4946
rect 3007 4942 3011 4946
rect 3127 4942 3131 4946
rect 3679 4942 3683 4946
rect 3799 4942 3803 4946
rect 111 4858 115 4862
rect 131 4858 135 4862
rect 267 4858 271 4862
rect 315 4858 319 4862
rect 403 4858 407 4862
rect 523 4858 527 4862
rect 539 4858 543 4862
rect 675 4858 679 4862
rect 723 4858 727 4862
rect 915 4858 919 4862
rect 1099 4858 1103 4862
rect 1283 4858 1287 4862
rect 1459 4858 1463 4862
rect 1635 4858 1639 4862
rect 1787 4858 1791 4862
rect 1935 4858 1939 4862
rect 3839 4882 3843 4886
rect 3887 4882 3891 4886
rect 4047 4882 4051 4886
rect 4071 4882 4075 4886
rect 4239 4882 4243 4886
rect 4287 4882 4291 4886
rect 4439 4882 4443 4886
rect 4511 4882 4515 4886
rect 4655 4882 4659 4886
rect 4735 4882 4739 4886
rect 4871 4882 4875 4886
rect 4959 4882 4963 4886
rect 5095 4882 5099 4886
rect 5183 4882 5187 4886
rect 5327 4882 5331 4886
rect 5407 4882 5411 4886
rect 5663 4882 5667 4886
rect 1975 4806 1979 4810
rect 1995 4806 1999 4810
rect 2155 4806 2159 4810
rect 2347 4806 2351 4810
rect 2539 4806 2543 4810
rect 2731 4806 2735 4810
rect 2843 4806 2847 4810
rect 2931 4806 2935 4810
rect 2979 4806 2983 4810
rect 3131 4806 3135 4810
rect 3799 4806 3803 4810
rect 3839 4766 3843 4770
rect 3859 4766 3863 4770
rect 3915 4766 3919 4770
rect 4043 4766 4047 4770
rect 4187 4766 4191 4770
rect 4259 4766 4263 4770
rect 4467 4766 4471 4770
rect 4483 4766 4487 4770
rect 4707 4766 4711 4770
rect 4763 4766 4767 4770
rect 4931 4766 4935 4770
rect 5067 4766 5071 4770
rect 5155 4766 5159 4770
rect 5371 4766 5375 4770
rect 5379 4766 5383 4770
rect 5663 4766 5667 4770
rect 111 4738 115 4742
rect 159 4738 163 4742
rect 295 4738 299 4742
rect 343 4738 347 4742
rect 431 4738 435 4742
rect 567 4738 571 4742
rect 703 4738 707 4742
rect 807 4738 811 4742
rect 1055 4738 1059 4742
rect 1311 4738 1315 4742
rect 1575 4738 1579 4742
rect 1815 4738 1819 4742
rect 1935 4738 1939 4742
rect 1975 4690 1979 4694
rect 2023 4690 2027 4694
rect 2183 4690 2187 4694
rect 2239 4690 2243 4694
rect 2375 4690 2379 4694
rect 2471 4690 2475 4694
rect 2567 4690 2571 4694
rect 2695 4690 2699 4694
rect 2759 4690 2763 4694
rect 2919 4690 2923 4694
rect 2959 4690 2963 4694
rect 3143 4690 3147 4694
rect 3159 4690 3163 4694
rect 3367 4690 3371 4694
rect 3799 4690 3803 4694
rect 3839 4654 3843 4658
rect 3943 4654 3947 4658
rect 4063 4654 4067 4658
rect 4215 4654 4219 4658
rect 4327 4654 4331 4658
rect 4495 4654 4499 4658
rect 4599 4654 4603 4658
rect 4791 4654 4795 4658
rect 4871 4654 4875 4658
rect 5095 4654 5099 4658
rect 5151 4654 5155 4658
rect 5399 4654 5403 4658
rect 5439 4654 5443 4658
rect 5663 4654 5667 4658
rect 111 4610 115 4614
rect 131 4610 135 4614
rect 171 4610 175 4614
rect 315 4610 319 4614
rect 395 4610 399 4614
rect 539 4610 543 4614
rect 643 4610 647 4614
rect 779 4610 783 4614
rect 907 4610 911 4614
rect 1027 4610 1031 4614
rect 1195 4610 1199 4614
rect 1283 4610 1287 4614
rect 1491 4610 1495 4614
rect 1547 4610 1551 4614
rect 1787 4610 1791 4614
rect 1935 4610 1939 4614
rect 1975 4574 1979 4578
rect 1995 4574 1999 4578
rect 2099 4574 2103 4578
rect 2211 4574 2215 4578
rect 2347 4574 2351 4578
rect 2443 4574 2447 4578
rect 2579 4574 2583 4578
rect 2667 4574 2671 4578
rect 2795 4574 2799 4578
rect 2891 4574 2895 4578
rect 3003 4574 3007 4578
rect 3115 4574 3119 4578
rect 3203 4574 3207 4578
rect 3339 4574 3343 4578
rect 3403 4574 3407 4578
rect 3611 4574 3615 4578
rect 3799 4574 3803 4578
rect 3839 4542 3843 4546
rect 4035 4542 4039 4546
rect 4179 4542 4183 4546
rect 4299 4542 4303 4546
rect 4411 4542 4415 4546
rect 4571 4542 4575 4546
rect 4659 4542 4663 4546
rect 4843 4542 4847 4546
rect 4915 4542 4919 4546
rect 5123 4542 5127 4546
rect 5179 4542 5183 4546
rect 5411 4542 5415 4546
rect 5443 4542 5447 4546
rect 5663 4542 5667 4546
rect 111 4494 115 4498
rect 199 4494 203 4498
rect 423 4494 427 4498
rect 447 4494 451 4498
rect 655 4494 659 4498
rect 671 4494 675 4498
rect 887 4494 891 4498
rect 935 4494 939 4498
rect 1143 4494 1147 4498
rect 1223 4494 1227 4498
rect 1407 4494 1411 4498
rect 1519 4494 1523 4498
rect 1679 4494 1683 4498
rect 1815 4494 1819 4498
rect 1935 4494 1939 4498
rect 1975 4454 1979 4458
rect 2127 4454 2131 4458
rect 2231 4454 2235 4458
rect 2375 4454 2379 4458
rect 2447 4454 2451 4458
rect 2607 4454 2611 4458
rect 2663 4454 2667 4458
rect 2823 4454 2827 4458
rect 2871 4454 2875 4458
rect 3031 4454 3035 4458
rect 3079 4454 3083 4458
rect 3231 4454 3235 4458
rect 3287 4454 3291 4458
rect 3431 4454 3435 4458
rect 3495 4454 3499 4458
rect 3639 4454 3643 4458
rect 3679 4454 3683 4458
rect 3799 4454 3803 4458
rect 3839 4422 3843 4426
rect 4207 4422 4211 4426
rect 4359 4422 4363 4426
rect 4439 4422 4443 4426
rect 4519 4422 4523 4426
rect 4687 4422 4691 4426
rect 4879 4422 4883 4426
rect 4943 4422 4947 4426
rect 5079 4422 5083 4426
rect 5207 4422 5211 4426
rect 5287 4422 5291 4426
rect 5471 4422 5475 4426
rect 5503 4422 5507 4426
rect 5663 4422 5667 4426
rect 111 4378 115 4382
rect 419 4378 423 4382
rect 627 4378 631 4382
rect 667 4378 671 4382
rect 811 4378 815 4382
rect 859 4378 863 4382
rect 963 4378 967 4382
rect 1115 4378 1119 4382
rect 1123 4378 1127 4382
rect 1291 4378 1295 4382
rect 1379 4378 1383 4382
rect 1467 4378 1471 4382
rect 1651 4378 1655 4382
rect 1935 4378 1939 4382
rect 1975 4334 1979 4338
rect 2203 4334 2207 4338
rect 2307 4334 2311 4338
rect 2419 4334 2423 4338
rect 2459 4334 2463 4338
rect 2627 4334 2631 4338
rect 2635 4334 2639 4338
rect 2811 4334 2815 4338
rect 2843 4334 2847 4338
rect 3011 4334 3015 4338
rect 3051 4334 3055 4338
rect 3227 4334 3231 4338
rect 3259 4334 3263 4338
rect 3451 4334 3455 4338
rect 3467 4334 3471 4338
rect 3651 4334 3655 4338
rect 3799 4334 3803 4338
rect 3839 4310 3843 4314
rect 3859 4310 3863 4314
rect 4043 4310 4047 4314
rect 4251 4310 4255 4314
rect 4331 4310 4335 4314
rect 4475 4310 4479 4314
rect 4491 4310 4495 4314
rect 4659 4310 4663 4314
rect 4715 4310 4719 4314
rect 4851 4310 4855 4314
rect 4971 4310 4975 4314
rect 5051 4310 5055 4314
rect 5235 4310 5239 4314
rect 5259 4310 5263 4314
rect 5475 4310 5479 4314
rect 5499 4310 5503 4314
rect 5663 4310 5667 4314
rect 111 4250 115 4254
rect 695 4250 699 4254
rect 815 4250 819 4254
rect 839 4250 843 4254
rect 951 4250 955 4254
rect 991 4250 995 4254
rect 1087 4250 1091 4254
rect 1151 4250 1155 4254
rect 1223 4250 1227 4254
rect 1319 4250 1323 4254
rect 1359 4250 1363 4254
rect 1495 4250 1499 4254
rect 1631 4250 1635 4254
rect 1679 4250 1683 4254
rect 1767 4250 1771 4254
rect 1935 4250 1939 4254
rect 1975 4214 1979 4218
rect 2335 4214 2339 4218
rect 2487 4214 2491 4218
rect 2567 4214 2571 4218
rect 2655 4214 2659 4218
rect 2703 4214 2707 4218
rect 2839 4214 2843 4218
rect 2975 4214 2979 4218
rect 3039 4214 3043 4218
rect 3255 4214 3259 4218
rect 3479 4214 3483 4218
rect 3679 4214 3683 4218
rect 3799 4214 3803 4218
rect 111 4134 115 4138
rect 731 4134 735 4138
rect 787 4134 791 4138
rect 867 4134 871 4138
rect 923 4134 927 4138
rect 1003 4134 1007 4138
rect 1059 4134 1063 4138
rect 1139 4134 1143 4138
rect 1195 4134 1199 4138
rect 1275 4134 1279 4138
rect 1331 4134 1335 4138
rect 1411 4134 1415 4138
rect 1467 4134 1471 4138
rect 1547 4134 1551 4138
rect 1603 4134 1607 4138
rect 1739 4134 1743 4138
rect 1935 4134 1939 4138
rect 3839 4162 3843 4166
rect 3887 4162 3891 4166
rect 4071 4162 4075 4166
rect 4279 4162 4283 4166
rect 4415 4162 4419 4166
rect 4503 4162 4507 4166
rect 4743 4162 4747 4166
rect 4975 4162 4979 4166
rect 4999 4162 5003 4166
rect 5263 4162 5267 4166
rect 5527 4162 5531 4166
rect 5543 4162 5547 4166
rect 5663 4162 5667 4166
rect 1975 4082 1979 4086
rect 2291 4082 2295 4086
rect 2427 4082 2431 4086
rect 2539 4082 2543 4086
rect 2563 4082 2567 4086
rect 2675 4082 2679 4086
rect 2699 4082 2703 4086
rect 2811 4082 2815 4086
rect 2835 4082 2839 4086
rect 2947 4082 2951 4086
rect 3799 4082 3803 4086
rect 3839 4050 3843 4054
rect 3859 4050 3863 4054
rect 4003 4050 4007 4054
rect 4171 4050 4175 4054
rect 4339 4050 4343 4054
rect 4387 4050 4391 4054
rect 4499 4050 4503 4054
rect 4651 4050 4655 4054
rect 4803 4050 4807 4054
rect 4947 4050 4951 4054
rect 5091 4050 5095 4054
rect 5235 4050 5239 4054
rect 5379 4050 5383 4054
rect 5515 4050 5519 4054
rect 5663 4050 5667 4054
rect 111 3998 115 4002
rect 511 3998 515 4002
rect 663 3998 667 4002
rect 759 3998 763 4002
rect 823 3998 827 4002
rect 895 3998 899 4002
rect 983 3998 987 4002
rect 1031 3998 1035 4002
rect 1151 3998 1155 4002
rect 1167 3998 1171 4002
rect 1303 3998 1307 4002
rect 1319 3998 1323 4002
rect 1439 3998 1443 4002
rect 1575 3998 1579 4002
rect 1935 3998 1939 4002
rect 1975 3966 1979 3970
rect 2119 3966 2123 3970
rect 2319 3966 2323 3970
rect 2327 3966 2331 3970
rect 2455 3966 2459 3970
rect 2535 3966 2539 3970
rect 2591 3966 2595 3970
rect 2727 3966 2731 3970
rect 2743 3966 2747 3970
rect 2863 3966 2867 3970
rect 2943 3966 2947 3970
rect 3135 3966 3139 3970
rect 3319 3966 3323 3970
rect 3511 3966 3515 3970
rect 3679 3966 3683 3970
rect 3799 3966 3803 3970
rect 111 3858 115 3862
rect 131 3858 135 3862
rect 307 3858 311 3862
rect 483 3858 487 3862
rect 515 3858 519 3862
rect 635 3858 639 3862
rect 723 3858 727 3862
rect 795 3858 799 3862
rect 939 3858 943 3862
rect 955 3858 959 3862
rect 1123 3858 1127 3862
rect 1163 3858 1167 3862
rect 1291 3858 1295 3862
rect 1935 3858 1939 3862
rect 3839 3914 3843 3918
rect 3887 3914 3891 3918
rect 4031 3914 4035 3918
rect 4199 3914 4203 3918
rect 4367 3914 4371 3918
rect 4383 3914 4387 3918
rect 4527 3914 4531 3918
rect 4599 3914 4603 3918
rect 4679 3914 4683 3918
rect 4823 3914 4827 3918
rect 4831 3914 4835 3918
rect 4975 3914 4979 3918
rect 5063 3914 5067 3918
rect 5119 3914 5123 3918
rect 5263 3914 5267 3918
rect 5311 3914 5315 3918
rect 5407 3914 5411 3918
rect 5543 3914 5547 3918
rect 5663 3914 5667 3918
rect 1975 3842 1979 3846
rect 2091 3842 2095 3846
rect 2139 3842 2143 3846
rect 2299 3842 2303 3846
rect 2371 3842 2375 3846
rect 2507 3842 2511 3846
rect 2587 3842 2591 3846
rect 2715 3842 2719 3846
rect 2795 3842 2799 3846
rect 2915 3842 2919 3846
rect 2995 3842 2999 3846
rect 3107 3842 3111 3846
rect 3195 3842 3199 3846
rect 3291 3842 3295 3846
rect 3403 3842 3407 3846
rect 3483 3842 3487 3846
rect 3651 3842 3655 3846
rect 3799 3842 3803 3846
rect 3839 3786 3843 3790
rect 3995 3786 3999 3790
rect 4203 3786 4207 3790
rect 4355 3786 4359 3790
rect 4435 3786 4439 3790
rect 4571 3786 4575 3790
rect 4691 3786 4695 3790
rect 4795 3786 4799 3790
rect 4963 3786 4967 3790
rect 5035 3786 5039 3790
rect 5251 3786 5255 3790
rect 5283 3786 5287 3790
rect 5515 3786 5519 3790
rect 5663 3786 5667 3790
rect 111 3746 115 3750
rect 159 3746 163 3750
rect 335 3746 339 3750
rect 527 3746 531 3750
rect 543 3746 547 3750
rect 711 3746 715 3750
rect 751 3746 755 3750
rect 887 3746 891 3750
rect 967 3746 971 3750
rect 1055 3746 1059 3750
rect 1191 3746 1195 3750
rect 1215 3746 1219 3750
rect 1367 3746 1371 3750
rect 1519 3746 1523 3750
rect 1679 3746 1683 3750
rect 1815 3746 1819 3750
rect 1935 3746 1939 3750
rect 1975 3726 1979 3730
rect 2167 3726 2171 3730
rect 2279 3726 2283 3730
rect 2399 3726 2403 3730
rect 2479 3726 2483 3730
rect 2615 3726 2619 3730
rect 2679 3726 2683 3730
rect 2823 3726 2827 3730
rect 2879 3726 2883 3730
rect 3023 3726 3027 3730
rect 3079 3726 3083 3730
rect 3223 3726 3227 3730
rect 3279 3726 3283 3730
rect 3431 3726 3435 3730
rect 3799 3726 3803 3730
rect 111 3622 115 3626
rect 131 3622 135 3626
rect 147 3622 151 3626
rect 307 3622 311 3626
rect 355 3622 359 3626
rect 499 3622 503 3626
rect 571 3622 575 3626
rect 683 3622 687 3626
rect 803 3622 807 3626
rect 859 3622 863 3626
rect 1027 3622 1031 3626
rect 1043 3622 1047 3626
rect 1187 3622 1191 3626
rect 1291 3622 1295 3626
rect 1339 3622 1343 3626
rect 1491 3622 1495 3626
rect 1547 3622 1551 3626
rect 1651 3622 1655 3626
rect 1787 3622 1791 3626
rect 1935 3622 1939 3626
rect 3839 3646 3843 3650
rect 4023 3646 4027 3650
rect 4215 3646 4219 3650
rect 4231 3646 4235 3650
rect 4399 3646 4403 3650
rect 4463 3646 4467 3650
rect 4607 3646 4611 3650
rect 4719 3646 4723 3650
rect 4831 3646 4835 3650
rect 4991 3646 4995 3650
rect 5071 3646 5075 3650
rect 5279 3646 5283 3650
rect 5319 3646 5323 3650
rect 5543 3646 5547 3650
rect 5663 3646 5667 3650
rect 1975 3602 1979 3606
rect 1995 3602 1999 3606
rect 2251 3602 2255 3606
rect 2451 3602 2455 3606
rect 2515 3602 2519 3606
rect 2651 3602 2655 3606
rect 2755 3602 2759 3606
rect 2851 3602 2855 3606
rect 2979 3602 2983 3606
rect 3051 3602 3055 3606
rect 3195 3602 3199 3606
rect 3251 3602 3255 3606
rect 3411 3602 3415 3606
rect 3627 3602 3631 3606
rect 3799 3602 3803 3606
rect 111 3486 115 3490
rect 175 3486 179 3490
rect 303 3486 307 3490
rect 383 3486 387 3490
rect 447 3486 451 3490
rect 599 3486 603 3490
rect 759 3486 763 3490
rect 831 3486 835 3490
rect 935 3486 939 3490
rect 1071 3486 1075 3490
rect 1111 3486 1115 3490
rect 1295 3486 1299 3490
rect 1319 3486 1323 3490
rect 1487 3486 1491 3490
rect 1575 3486 1579 3490
rect 1815 3486 1819 3490
rect 1935 3486 1939 3490
rect 3839 3510 3843 3514
rect 4187 3510 4191 3514
rect 4371 3510 4375 3514
rect 4531 3510 4535 3514
rect 4579 3510 4583 3514
rect 4683 3510 4687 3514
rect 4803 3510 4807 3514
rect 4843 3510 4847 3514
rect 5003 3510 5007 3514
rect 5043 3510 5047 3514
rect 5171 3510 5175 3514
rect 5291 3510 5295 3514
rect 5347 3510 5351 3514
rect 5515 3510 5519 3514
rect 5663 3510 5667 3514
rect 1975 3482 1979 3486
rect 2023 3482 2027 3486
rect 2191 3482 2195 3486
rect 2279 3482 2283 3486
rect 2399 3482 2403 3486
rect 2543 3482 2547 3486
rect 2615 3482 2619 3486
rect 2783 3482 2787 3486
rect 2831 3482 2835 3486
rect 3007 3482 3011 3486
rect 3047 3482 3051 3486
rect 3223 3482 3227 3486
rect 3263 3482 3267 3486
rect 3439 3482 3443 3486
rect 3479 3482 3483 3486
rect 3655 3482 3659 3486
rect 3679 3482 3683 3486
rect 3799 3482 3803 3486
rect 111 3358 115 3362
rect 275 3358 279 3362
rect 419 3358 423 3362
rect 467 3358 471 3362
rect 571 3358 575 3362
rect 667 3358 671 3362
rect 731 3358 735 3362
rect 875 3358 879 3362
rect 907 3358 911 3362
rect 1083 3358 1087 3362
rect 1091 3358 1095 3362
rect 1267 3358 1271 3362
rect 1315 3358 1319 3362
rect 1459 3358 1463 3362
rect 1935 3358 1939 3362
rect 3839 3394 3843 3398
rect 3887 3394 3891 3398
rect 4151 3394 4155 3398
rect 4423 3394 4427 3398
rect 4559 3394 4563 3398
rect 4671 3394 4675 3398
rect 4711 3394 4715 3398
rect 4871 3394 4875 3398
rect 4895 3394 4899 3398
rect 5031 3394 5035 3398
rect 5111 3394 5115 3398
rect 5199 3394 5203 3398
rect 5327 3394 5331 3398
rect 5375 3394 5379 3398
rect 5543 3394 5547 3398
rect 5663 3394 5667 3398
rect 1975 3330 1979 3334
rect 1995 3330 1999 3334
rect 2163 3330 2167 3334
rect 2195 3330 2199 3334
rect 2371 3330 2375 3334
rect 2411 3330 2415 3334
rect 2587 3330 2591 3334
rect 2619 3330 2623 3334
rect 2803 3330 2807 3334
rect 2811 3330 2815 3334
rect 3003 3330 3007 3334
rect 3019 3330 3023 3334
rect 3187 3330 3191 3334
rect 3235 3330 3239 3334
rect 3371 3330 3375 3334
rect 3451 3330 3455 3334
rect 3555 3330 3559 3334
rect 3651 3330 3655 3334
rect 3799 3330 3803 3334
rect 3839 3282 3843 3286
rect 3859 3282 3863 3286
rect 4099 3282 4103 3286
rect 4123 3282 4127 3286
rect 4347 3282 4351 3286
rect 4395 3282 4399 3286
rect 4579 3282 4583 3286
rect 4643 3282 4647 3286
rect 4787 3282 4791 3286
rect 4867 3282 4871 3286
rect 4987 3282 4991 3286
rect 5083 3282 5087 3286
rect 5171 3282 5175 3286
rect 5299 3282 5303 3286
rect 5355 3282 5359 3286
rect 5515 3282 5519 3286
rect 5663 3282 5667 3286
rect 111 3246 115 3250
rect 495 3246 499 3250
rect 535 3246 539 3250
rect 695 3246 699 3250
rect 727 3246 731 3250
rect 903 3246 907 3250
rect 919 3246 923 3250
rect 1111 3246 1115 3250
rect 1119 3246 1123 3250
rect 1295 3246 1299 3250
rect 1343 3246 1347 3250
rect 1471 3246 1475 3250
rect 1655 3246 1659 3250
rect 1815 3246 1819 3250
rect 1935 3246 1939 3250
rect 1975 3218 1979 3222
rect 2023 3218 2027 3222
rect 2223 3218 2227 3222
rect 2439 3218 2443 3222
rect 2463 3218 2467 3222
rect 2647 3218 2651 3222
rect 2663 3218 2667 3222
rect 2839 3218 2843 3222
rect 2863 3218 2867 3222
rect 3031 3218 3035 3222
rect 3055 3218 3059 3222
rect 3215 3218 3219 3222
rect 3239 3218 3243 3222
rect 3399 3218 3403 3222
rect 3431 3218 3435 3222
rect 3583 3218 3587 3222
rect 3623 3218 3627 3222
rect 3799 3218 3803 3222
rect 111 3126 115 3130
rect 427 3126 431 3130
rect 507 3126 511 3130
rect 563 3126 567 3130
rect 699 3126 703 3130
rect 835 3126 839 3130
rect 891 3126 895 3130
rect 971 3126 975 3130
rect 1083 3126 1087 3130
rect 1107 3126 1111 3130
rect 1243 3126 1247 3130
rect 1267 3126 1271 3130
rect 1379 3126 1383 3130
rect 1443 3126 1447 3130
rect 1515 3126 1519 3130
rect 1627 3126 1631 3130
rect 1651 3126 1655 3130
rect 1787 3126 1791 3130
rect 1935 3126 1939 3130
rect 3839 3154 3843 3158
rect 3887 3154 3891 3158
rect 3903 3154 3907 3158
rect 4127 3154 4131 3158
rect 4135 3154 4139 3158
rect 4359 3154 4363 3158
rect 4375 3154 4379 3158
rect 4583 3154 4587 3158
rect 4607 3154 4611 3158
rect 4807 3154 4811 3158
rect 4815 3154 4819 3158
rect 5015 3154 5019 3158
rect 5031 3154 5035 3158
rect 5199 3154 5203 3158
rect 5383 3154 5387 3158
rect 5543 3154 5547 3158
rect 5663 3154 5667 3158
rect 1975 3094 1979 3098
rect 2331 3094 2335 3098
rect 2435 3094 2439 3098
rect 2555 3094 2559 3098
rect 2635 3094 2639 3098
rect 2779 3094 2783 3098
rect 2835 3094 2839 3098
rect 3003 3094 3007 3098
rect 3027 3094 3031 3098
rect 3211 3094 3215 3098
rect 3235 3094 3239 3098
rect 3403 3094 3407 3098
rect 3467 3094 3471 3098
rect 3595 3094 3599 3098
rect 3799 3094 3803 3098
rect 3839 3042 3843 3046
rect 3875 3042 3879 3046
rect 3907 3042 3911 3046
rect 4075 3042 4079 3046
rect 4107 3042 4111 3046
rect 4243 3042 4247 3046
rect 4331 3042 4335 3046
rect 4411 3042 4415 3046
rect 4555 3042 4559 3046
rect 4579 3042 4583 3046
rect 4755 3042 4759 3046
rect 4779 3042 4783 3046
rect 5003 3042 5007 3046
rect 5663 3042 5667 3046
rect 111 2986 115 2990
rect 199 2986 203 2990
rect 455 2986 459 2990
rect 511 2986 515 2990
rect 591 2986 595 2990
rect 727 2986 731 2990
rect 815 2986 819 2990
rect 863 2986 867 2990
rect 999 2986 1003 2990
rect 1111 2986 1115 2990
rect 1135 2986 1139 2990
rect 1271 2986 1275 2990
rect 1407 2986 1411 2990
rect 1415 2986 1419 2990
rect 1543 2986 1547 2990
rect 1679 2986 1683 2990
rect 1719 2986 1723 2990
rect 1815 2986 1819 2990
rect 1935 2986 1939 2990
rect 1975 2970 1979 2974
rect 2143 2970 2147 2974
rect 2343 2970 2347 2974
rect 2359 2970 2363 2974
rect 2543 2970 2547 2974
rect 2583 2970 2587 2974
rect 2743 2970 2747 2974
rect 2807 2970 2811 2974
rect 2935 2970 2939 2974
rect 3031 2970 3035 2974
rect 3135 2970 3139 2974
rect 3263 2970 3267 2974
rect 3335 2970 3339 2974
rect 3495 2970 3499 2974
rect 3799 2970 3803 2974
rect 3839 2926 3843 2930
rect 3895 2926 3899 2930
rect 3935 2926 3939 2930
rect 4031 2926 4035 2930
rect 4103 2926 4107 2930
rect 4167 2926 4171 2930
rect 4271 2926 4275 2930
rect 4303 2926 4307 2930
rect 4439 2926 4443 2930
rect 4575 2926 4579 2930
rect 4607 2926 4611 2930
rect 4783 2926 4787 2930
rect 5663 2926 5667 2930
rect 111 2874 115 2878
rect 131 2874 135 2878
rect 171 2874 175 2878
rect 307 2874 311 2878
rect 483 2874 487 2878
rect 523 2874 527 2878
rect 763 2874 767 2878
rect 787 2874 791 2878
rect 1011 2874 1015 2878
rect 1083 2874 1087 2878
rect 1275 2874 1279 2878
rect 1387 2874 1391 2878
rect 1539 2874 1543 2878
rect 1691 2874 1695 2878
rect 1935 2874 1939 2878
rect 1975 2850 1979 2854
rect 2011 2850 2015 2854
rect 2115 2850 2119 2854
rect 2259 2850 2263 2854
rect 2315 2850 2319 2854
rect 2507 2850 2511 2854
rect 2515 2850 2519 2854
rect 2715 2850 2719 2854
rect 2755 2850 2759 2854
rect 2907 2850 2911 2854
rect 3003 2850 3007 2854
rect 3107 2850 3111 2854
rect 3307 2850 3311 2854
rect 3799 2850 3803 2854
rect 3839 2806 3843 2810
rect 3859 2806 3863 2810
rect 3867 2806 3871 2810
rect 3995 2806 3999 2810
rect 4003 2806 4007 2810
rect 4131 2806 4135 2810
rect 4139 2806 4143 2810
rect 4267 2806 4271 2810
rect 4275 2806 4279 2810
rect 4403 2806 4407 2810
rect 4411 2806 4415 2810
rect 4539 2806 4543 2810
rect 4547 2806 4551 2810
rect 4675 2806 4679 2810
rect 4811 2806 4815 2810
rect 5663 2806 5667 2810
rect 111 2758 115 2762
rect 159 2758 163 2762
rect 279 2758 283 2762
rect 335 2758 339 2762
rect 455 2758 459 2762
rect 551 2758 555 2762
rect 647 2758 651 2762
rect 791 2758 795 2762
rect 855 2758 859 2762
rect 1039 2758 1043 2762
rect 1079 2758 1083 2762
rect 1303 2758 1307 2762
rect 1311 2758 1315 2762
rect 1551 2758 1555 2762
rect 1567 2758 1571 2762
rect 1799 2758 1803 2762
rect 1935 2758 1939 2762
rect 1975 2734 1979 2738
rect 2023 2734 2027 2738
rect 2039 2734 2043 2738
rect 2247 2734 2251 2738
rect 2287 2734 2291 2738
rect 2503 2734 2507 2738
rect 2535 2734 2539 2738
rect 2759 2734 2763 2738
rect 2783 2734 2787 2738
rect 3015 2734 3019 2738
rect 3031 2734 3035 2738
rect 3799 2734 3803 2738
rect 3839 2694 3843 2698
rect 3887 2694 3891 2698
rect 3959 2694 3963 2698
rect 4023 2694 4027 2698
rect 4159 2694 4163 2698
rect 4255 2694 4259 2698
rect 4295 2694 4299 2698
rect 4431 2694 4435 2698
rect 4543 2694 4547 2698
rect 4567 2694 4571 2698
rect 4703 2694 4707 2698
rect 4823 2694 4827 2698
rect 4839 2694 4843 2698
rect 5111 2694 5115 2698
rect 5399 2694 5403 2698
rect 5663 2694 5667 2698
rect 111 2646 115 2650
rect 251 2646 255 2650
rect 427 2646 431 2650
rect 571 2646 575 2650
rect 619 2646 623 2650
rect 731 2646 735 2650
rect 827 2646 831 2650
rect 891 2646 895 2650
rect 1043 2646 1047 2650
rect 1051 2646 1055 2650
rect 1195 2646 1199 2650
rect 1283 2646 1287 2650
rect 1355 2646 1359 2650
rect 1515 2646 1519 2650
rect 1523 2646 1527 2650
rect 1675 2646 1679 2650
rect 1771 2646 1775 2650
rect 1935 2646 1939 2650
rect 1975 2610 1979 2614
rect 1995 2610 1999 2614
rect 2219 2610 2223 2614
rect 2475 2610 2479 2614
rect 2555 2610 2559 2614
rect 2691 2610 2695 2614
rect 2731 2610 2735 2614
rect 2827 2610 2831 2614
rect 2963 2610 2967 2614
rect 2987 2610 2991 2614
rect 3099 2610 3103 2614
rect 3799 2610 3803 2614
rect 3839 2582 3843 2586
rect 3859 2582 3863 2586
rect 3931 2582 3935 2586
rect 4083 2582 4087 2586
rect 4227 2582 4231 2586
rect 4331 2582 4335 2586
rect 4515 2582 4519 2586
rect 4579 2582 4583 2586
rect 4795 2582 4799 2586
rect 4827 2582 4831 2586
rect 5075 2582 5079 2586
rect 5083 2582 5087 2586
rect 5323 2582 5327 2586
rect 5371 2582 5375 2586
rect 5663 2582 5667 2586
rect 111 2534 115 2538
rect 383 2534 387 2538
rect 599 2534 603 2538
rect 759 2534 763 2538
rect 815 2534 819 2538
rect 919 2534 923 2538
rect 1023 2534 1027 2538
rect 1071 2534 1075 2538
rect 1223 2534 1227 2538
rect 1231 2534 1235 2538
rect 1383 2534 1387 2538
rect 1431 2534 1435 2538
rect 1543 2534 1547 2538
rect 1631 2534 1635 2538
rect 1703 2534 1707 2538
rect 1815 2534 1819 2538
rect 1935 2534 1939 2538
rect 1975 2474 1979 2478
rect 2023 2474 2027 2478
rect 2223 2474 2227 2478
rect 2447 2474 2451 2478
rect 2583 2474 2587 2478
rect 2679 2474 2683 2478
rect 2719 2474 2723 2478
rect 2855 2474 2859 2478
rect 2927 2474 2931 2478
rect 2991 2474 2995 2478
rect 3127 2474 3131 2478
rect 3183 2474 3187 2478
rect 3439 2474 3443 2478
rect 3679 2474 3683 2478
rect 3799 2474 3803 2478
rect 3839 2466 3843 2470
rect 3887 2466 3891 2470
rect 4087 2466 4091 2470
rect 4111 2466 4115 2470
rect 4327 2466 4331 2470
rect 4359 2466 4363 2470
rect 4583 2466 4587 2470
rect 4607 2466 4611 2470
rect 4847 2466 4851 2470
rect 4855 2466 4859 2470
rect 5103 2466 5107 2470
rect 5119 2466 5123 2470
rect 5351 2466 5355 2470
rect 5399 2466 5403 2470
rect 5663 2466 5667 2470
rect 111 2418 115 2422
rect 227 2418 231 2422
rect 355 2418 359 2422
rect 523 2418 527 2422
rect 571 2418 575 2422
rect 787 2418 791 2422
rect 835 2418 839 2422
rect 995 2418 999 2422
rect 1155 2418 1159 2422
rect 1203 2418 1207 2422
rect 1403 2418 1407 2422
rect 1483 2418 1487 2422
rect 1603 2418 1607 2422
rect 1787 2418 1791 2422
rect 1935 2418 1939 2422
rect 1975 2354 1979 2358
rect 1995 2354 1999 2358
rect 2155 2354 2159 2358
rect 2195 2354 2199 2358
rect 2347 2354 2351 2358
rect 2419 2354 2423 2358
rect 2539 2354 2543 2358
rect 2651 2354 2655 2358
rect 2731 2354 2735 2358
rect 2899 2354 2903 2358
rect 2923 2354 2927 2358
rect 3115 2354 3119 2358
rect 3155 2354 3159 2358
rect 3299 2354 3303 2358
rect 3411 2354 3415 2358
rect 3483 2354 3487 2358
rect 3651 2354 3655 2358
rect 3799 2354 3803 2358
rect 111 2290 115 2294
rect 159 2290 163 2294
rect 255 2290 259 2294
rect 367 2290 371 2294
rect 551 2290 555 2294
rect 599 2290 603 2294
rect 831 2290 835 2294
rect 863 2290 867 2294
rect 1063 2290 1067 2294
rect 1183 2290 1187 2294
rect 1511 2290 1515 2294
rect 1815 2290 1819 2294
rect 1935 2290 1939 2294
rect 3839 2342 3843 2346
rect 3859 2342 3863 2346
rect 4059 2342 4063 2346
rect 4299 2342 4303 2346
rect 4443 2342 4447 2346
rect 4555 2342 4559 2346
rect 4611 2342 4615 2346
rect 4787 2342 4791 2346
rect 4819 2342 4823 2346
rect 4963 2342 4967 2346
rect 5091 2342 5095 2346
rect 5147 2342 5151 2346
rect 5339 2342 5343 2346
rect 5371 2342 5375 2346
rect 5515 2342 5519 2346
rect 5663 2342 5667 2346
rect 1975 2234 1979 2238
rect 2023 2234 2027 2238
rect 2183 2234 2187 2238
rect 2191 2234 2195 2238
rect 2359 2234 2363 2238
rect 2375 2234 2379 2238
rect 2535 2234 2539 2238
rect 2567 2234 2571 2238
rect 2711 2234 2715 2238
rect 2759 2234 2763 2238
rect 2879 2234 2883 2238
rect 2951 2234 2955 2238
rect 3047 2234 3051 2238
rect 3143 2234 3147 2238
rect 3207 2234 3211 2238
rect 3327 2234 3331 2238
rect 3367 2234 3371 2238
rect 3511 2234 3515 2238
rect 3535 2234 3539 2238
rect 3679 2234 3683 2238
rect 3799 2234 3803 2238
rect 3839 2218 3843 2222
rect 4471 2218 4475 2222
rect 4543 2218 4547 2222
rect 4639 2218 4643 2222
rect 4719 2218 4723 2222
rect 4815 2218 4819 2222
rect 4911 2218 4915 2222
rect 4991 2218 4995 2222
rect 5119 2218 5123 2222
rect 5175 2218 5179 2222
rect 5335 2218 5339 2222
rect 5367 2218 5371 2222
rect 5543 2218 5547 2222
rect 5663 2218 5667 2222
rect 111 2166 115 2170
rect 131 2166 135 2170
rect 339 2166 343 2170
rect 347 2166 351 2170
rect 571 2166 575 2170
rect 595 2166 599 2170
rect 803 2166 807 2170
rect 835 2166 839 2170
rect 1035 2166 1039 2170
rect 1075 2166 1079 2170
rect 1315 2166 1319 2170
rect 1563 2166 1567 2170
rect 1787 2166 1791 2170
rect 1935 2166 1939 2170
rect 1975 2106 1979 2110
rect 1995 2106 1999 2110
rect 2163 2106 2167 2110
rect 2331 2106 2335 2110
rect 2507 2106 2511 2110
rect 2683 2106 2687 2110
rect 2851 2106 2855 2110
rect 3019 2106 3023 2110
rect 3107 2106 3111 2110
rect 3179 2106 3183 2110
rect 3243 2106 3247 2110
rect 3339 2106 3343 2110
rect 3379 2106 3383 2110
rect 3507 2106 3511 2110
rect 3515 2106 3519 2110
rect 3651 2106 3655 2110
rect 3799 2106 3803 2110
rect 3839 2106 3843 2110
rect 4515 2106 4519 2110
rect 4635 2106 4639 2110
rect 4691 2106 4695 2110
rect 4771 2106 4775 2110
rect 4883 2106 4887 2110
rect 4907 2106 4911 2110
rect 5043 2106 5047 2110
rect 5091 2106 5095 2110
rect 5179 2106 5183 2110
rect 5307 2106 5311 2110
rect 5515 2106 5519 2110
rect 5663 2106 5667 2110
rect 111 2050 115 2054
rect 159 2050 163 2054
rect 271 2050 275 2054
rect 375 2050 379 2054
rect 407 2050 411 2054
rect 543 2050 547 2054
rect 623 2050 627 2054
rect 687 2050 691 2054
rect 831 2050 835 2054
rect 863 2050 867 2054
rect 975 2050 979 2054
rect 1103 2050 1107 2054
rect 1119 2050 1123 2054
rect 1263 2050 1267 2054
rect 1343 2050 1347 2054
rect 1407 2050 1411 2054
rect 1543 2050 1547 2054
rect 1591 2050 1595 2054
rect 1679 2050 1683 2054
rect 1815 2050 1819 2054
rect 1935 2050 1939 2054
rect 1975 1994 1979 1998
rect 3127 1994 3131 1998
rect 3135 1994 3139 1998
rect 3263 1994 3267 1998
rect 3271 1994 3275 1998
rect 3399 1994 3403 1998
rect 3407 1994 3411 1998
rect 3535 1994 3539 1998
rect 3543 1994 3547 1998
rect 3671 1994 3675 1998
rect 3679 1994 3683 1998
rect 3799 1994 3803 1998
rect 3839 1994 3843 1998
rect 4663 1994 4667 1998
rect 4799 1994 4803 1998
rect 4863 1994 4867 1998
rect 4935 1994 4939 1998
rect 4999 1994 5003 1998
rect 5071 1994 5075 1998
rect 5135 1994 5139 1998
rect 5207 1994 5211 1998
rect 5271 1994 5275 1998
rect 5407 1994 5411 1998
rect 5543 1994 5547 1998
rect 5663 1994 5667 1998
rect 111 1934 115 1938
rect 187 1934 191 1938
rect 243 1934 247 1938
rect 379 1934 383 1938
rect 515 1934 519 1938
rect 587 1934 591 1938
rect 659 1934 663 1938
rect 803 1934 807 1938
rect 811 1934 815 1938
rect 947 1934 951 1938
rect 1051 1934 1055 1938
rect 1091 1934 1095 1938
rect 1235 1934 1239 1938
rect 1299 1934 1303 1938
rect 1379 1934 1383 1938
rect 1515 1934 1519 1938
rect 1555 1934 1559 1938
rect 1651 1934 1655 1938
rect 1787 1934 1791 1938
rect 1935 1934 1939 1938
rect 1975 1870 1979 1874
rect 1995 1870 1999 1874
rect 2227 1870 2231 1874
rect 2467 1870 2471 1874
rect 2691 1870 2695 1874
rect 2907 1870 2911 1874
rect 3099 1870 3103 1874
rect 3107 1870 3111 1874
rect 3235 1870 3239 1874
rect 3299 1870 3303 1874
rect 3371 1870 3375 1874
rect 3483 1870 3487 1874
rect 3507 1870 3511 1874
rect 3643 1870 3647 1874
rect 3651 1870 3655 1874
rect 3799 1870 3803 1874
rect 3839 1870 3843 1874
rect 4675 1870 4679 1874
rect 4819 1870 4823 1874
rect 4835 1870 4839 1874
rect 4963 1870 4967 1874
rect 4971 1870 4975 1874
rect 5107 1870 5111 1874
rect 5243 1870 5247 1874
rect 5379 1870 5383 1874
rect 5515 1870 5519 1874
rect 5663 1870 5667 1874
rect 111 1814 115 1818
rect 159 1814 163 1818
rect 215 1814 219 1818
rect 375 1814 379 1818
rect 407 1814 411 1818
rect 591 1814 595 1818
rect 615 1814 619 1818
rect 799 1814 803 1818
rect 839 1814 843 1818
rect 999 1814 1003 1818
rect 1079 1814 1083 1818
rect 1191 1814 1195 1818
rect 1327 1814 1331 1818
rect 1383 1814 1387 1818
rect 1575 1814 1579 1818
rect 1583 1814 1587 1818
rect 1815 1814 1819 1818
rect 1935 1814 1939 1818
rect 1975 1750 1979 1754
rect 2023 1750 2027 1754
rect 2159 1750 2163 1754
rect 2255 1750 2259 1754
rect 2311 1750 2315 1754
rect 2471 1750 2475 1754
rect 2495 1750 2499 1754
rect 2639 1750 2643 1754
rect 2719 1750 2723 1754
rect 2807 1750 2811 1754
rect 2935 1750 2939 1754
rect 2975 1750 2979 1754
rect 3135 1750 3139 1754
rect 3151 1750 3155 1754
rect 3327 1750 3331 1754
rect 3511 1750 3515 1754
rect 3679 1750 3683 1754
rect 3799 1750 3803 1754
rect 3839 1742 3843 1746
rect 3887 1742 3891 1746
rect 4079 1742 4083 1746
rect 4303 1742 4307 1746
rect 4535 1742 4539 1746
rect 4703 1742 4707 1746
rect 4775 1742 4779 1746
rect 4847 1742 4851 1746
rect 4991 1742 4995 1746
rect 5023 1742 5027 1746
rect 5135 1742 5139 1746
rect 5271 1742 5275 1746
rect 5279 1742 5283 1746
rect 5407 1742 5411 1746
rect 5535 1742 5539 1746
rect 5543 1742 5547 1746
rect 5663 1742 5667 1746
rect 111 1678 115 1682
rect 131 1678 135 1682
rect 347 1678 351 1682
rect 395 1678 399 1682
rect 563 1678 567 1682
rect 683 1678 687 1682
rect 771 1678 775 1682
rect 971 1678 975 1682
rect 979 1678 983 1682
rect 1163 1678 1167 1682
rect 1275 1678 1279 1682
rect 1355 1678 1359 1682
rect 1547 1678 1551 1682
rect 1935 1678 1939 1682
rect 1975 1630 1979 1634
rect 1995 1630 1999 1634
rect 2091 1630 2095 1634
rect 2131 1630 2135 1634
rect 2227 1630 2231 1634
rect 2283 1630 2287 1634
rect 2363 1630 2367 1634
rect 2443 1630 2447 1634
rect 2499 1630 2503 1634
rect 2611 1630 2615 1634
rect 2635 1630 2639 1634
rect 2771 1630 2775 1634
rect 2779 1630 2783 1634
rect 2907 1630 2911 1634
rect 2947 1630 2951 1634
rect 3043 1630 3047 1634
rect 3123 1630 3127 1634
rect 3179 1630 3183 1634
rect 3799 1630 3803 1634
rect 3839 1630 3843 1634
rect 3859 1630 3863 1634
rect 3995 1630 3999 1634
rect 4051 1630 4055 1634
rect 4155 1630 4159 1634
rect 4275 1630 4279 1634
rect 4355 1630 4359 1634
rect 4507 1630 4511 1634
rect 4587 1630 4591 1634
rect 4747 1630 4751 1634
rect 4851 1630 4855 1634
rect 4995 1630 4999 1634
rect 5131 1630 5135 1634
rect 5251 1630 5255 1634
rect 5419 1630 5423 1634
rect 5507 1630 5511 1634
rect 5663 1630 5667 1634
rect 111 1554 115 1558
rect 159 1554 163 1558
rect 375 1554 379 1558
rect 423 1554 427 1558
rect 607 1554 611 1558
rect 711 1554 715 1558
rect 839 1554 843 1558
rect 1007 1554 1011 1558
rect 1071 1554 1075 1558
rect 1303 1554 1307 1558
rect 1935 1554 1939 1558
rect 3839 1518 3843 1522
rect 3887 1518 3891 1522
rect 4023 1518 4027 1522
rect 4159 1518 4163 1522
rect 4183 1518 4187 1522
rect 4303 1518 4307 1522
rect 4383 1518 4387 1522
rect 4495 1518 4499 1522
rect 4615 1518 4619 1522
rect 4719 1518 4723 1522
rect 4879 1518 4883 1522
rect 4967 1518 4971 1522
rect 5159 1518 5163 1522
rect 5223 1518 5227 1522
rect 5447 1518 5451 1522
rect 5487 1518 5491 1522
rect 5663 1518 5667 1522
rect 1975 1498 1979 1502
rect 2023 1498 2027 1502
rect 2119 1498 2123 1502
rect 2159 1498 2163 1502
rect 2255 1498 2259 1502
rect 2295 1498 2299 1502
rect 2391 1498 2395 1502
rect 2431 1498 2435 1502
rect 2527 1498 2531 1502
rect 2567 1498 2571 1502
rect 2663 1498 2667 1502
rect 2703 1498 2707 1502
rect 2799 1498 2803 1502
rect 2839 1498 2843 1502
rect 2935 1498 2939 1502
rect 2975 1498 2979 1502
rect 3071 1498 3075 1502
rect 3207 1498 3211 1502
rect 3799 1498 3803 1502
rect 111 1430 115 1434
rect 131 1430 135 1434
rect 347 1430 351 1434
rect 411 1430 415 1434
rect 579 1430 583 1434
rect 739 1430 743 1434
rect 811 1430 815 1434
rect 1043 1430 1047 1434
rect 1091 1430 1095 1434
rect 1275 1430 1279 1434
rect 1451 1430 1455 1434
rect 1787 1430 1791 1434
rect 1935 1430 1939 1434
rect 3839 1402 3843 1406
rect 3859 1402 3863 1406
rect 3995 1402 3999 1406
rect 4059 1402 4063 1406
rect 4131 1402 4135 1406
rect 4275 1402 4279 1406
rect 4307 1402 4311 1406
rect 4467 1402 4471 1406
rect 4579 1402 4583 1406
rect 4691 1402 4695 1406
rect 4875 1402 4879 1406
rect 4939 1402 4943 1406
rect 5187 1402 5191 1406
rect 5195 1402 5199 1406
rect 5459 1402 5463 1406
rect 5499 1402 5503 1406
rect 5663 1402 5667 1406
rect 1975 1378 1979 1382
rect 1995 1378 1999 1382
rect 2131 1378 2135 1382
rect 2267 1378 2271 1382
rect 2275 1378 2279 1382
rect 2403 1378 2407 1382
rect 2539 1378 2543 1382
rect 2563 1378 2567 1382
rect 2675 1378 2679 1382
rect 2811 1378 2815 1382
rect 2843 1378 2847 1382
rect 2947 1378 2951 1382
rect 3123 1378 3127 1382
rect 3395 1378 3399 1382
rect 3651 1378 3655 1382
rect 3799 1378 3803 1382
rect 111 1318 115 1322
rect 159 1318 163 1322
rect 359 1318 363 1322
rect 439 1318 443 1322
rect 575 1318 579 1322
rect 767 1318 771 1322
rect 775 1318 779 1322
rect 967 1318 971 1322
rect 1119 1318 1123 1322
rect 1151 1318 1155 1322
rect 1327 1318 1331 1322
rect 1479 1318 1483 1322
rect 1495 1318 1499 1322
rect 1663 1318 1667 1322
rect 1815 1318 1819 1322
rect 1935 1318 1939 1322
rect 3839 1282 3843 1286
rect 3887 1282 3891 1286
rect 4087 1282 4091 1286
rect 4335 1282 4339 1286
rect 4607 1282 4611 1286
rect 4615 1282 4619 1286
rect 4791 1282 4795 1286
rect 4903 1282 4907 1286
rect 4975 1282 4979 1286
rect 5167 1282 5171 1286
rect 5215 1282 5219 1286
rect 5367 1282 5371 1286
rect 5527 1282 5531 1286
rect 5543 1282 5547 1286
rect 5663 1282 5667 1286
rect 1975 1242 1979 1246
rect 2023 1242 2027 1246
rect 2303 1242 2307 1246
rect 2591 1242 2595 1246
rect 2655 1242 2659 1246
rect 2831 1242 2835 1246
rect 2871 1242 2875 1246
rect 3007 1242 3011 1246
rect 3151 1242 3155 1246
rect 3183 1242 3187 1246
rect 3359 1242 3363 1246
rect 3423 1242 3427 1246
rect 3543 1242 3547 1246
rect 3679 1242 3683 1246
rect 3799 1242 3803 1246
rect 111 1194 115 1198
rect 131 1194 135 1198
rect 291 1194 295 1198
rect 331 1194 335 1198
rect 475 1194 479 1198
rect 547 1194 551 1198
rect 659 1194 663 1198
rect 747 1194 751 1198
rect 835 1194 839 1198
rect 939 1194 943 1198
rect 1003 1194 1007 1198
rect 1123 1194 1127 1198
rect 1171 1194 1175 1198
rect 1299 1194 1303 1198
rect 1331 1194 1335 1198
rect 1467 1194 1471 1198
rect 1491 1194 1495 1198
rect 1635 1194 1639 1198
rect 1651 1194 1655 1198
rect 1787 1194 1791 1198
rect 1935 1194 1939 1198
rect 3839 1166 3843 1170
rect 4587 1166 4591 1170
rect 4763 1166 4767 1170
rect 4835 1166 4839 1170
rect 4947 1166 4951 1170
rect 4971 1166 4975 1170
rect 5107 1166 5111 1170
rect 5139 1166 5143 1170
rect 5243 1166 5247 1170
rect 5339 1166 5343 1170
rect 5379 1166 5383 1170
rect 5515 1166 5519 1170
rect 5663 1166 5667 1170
rect 1975 1114 1979 1118
rect 1995 1114 1999 1118
rect 2171 1114 2175 1118
rect 2363 1114 2367 1118
rect 2547 1114 2551 1118
rect 2627 1114 2631 1118
rect 2723 1114 2727 1118
rect 2803 1114 2807 1118
rect 2891 1114 2895 1118
rect 2979 1114 2983 1118
rect 3059 1114 3063 1118
rect 3155 1114 3159 1118
rect 3219 1114 3223 1118
rect 3331 1114 3335 1118
rect 3387 1114 3391 1118
rect 3515 1114 3519 1118
rect 3799 1114 3803 1118
rect 111 1070 115 1074
rect 159 1070 163 1074
rect 175 1070 179 1074
rect 319 1070 323 1074
rect 431 1070 435 1074
rect 503 1070 507 1074
rect 687 1070 691 1074
rect 863 1070 867 1074
rect 951 1070 955 1074
rect 1031 1070 1035 1074
rect 1199 1070 1203 1074
rect 1215 1070 1219 1074
rect 1359 1070 1363 1074
rect 1519 1070 1523 1074
rect 1679 1070 1683 1074
rect 1815 1070 1819 1074
rect 1935 1070 1939 1074
rect 3839 1050 3843 1054
rect 4807 1050 4811 1054
rect 4863 1050 4867 1054
rect 4943 1050 4947 1054
rect 4999 1050 5003 1054
rect 5079 1050 5083 1054
rect 5135 1050 5139 1054
rect 5215 1050 5219 1054
rect 5271 1050 5275 1054
rect 5351 1050 5355 1054
rect 5407 1050 5411 1054
rect 5487 1050 5491 1054
rect 5543 1050 5547 1054
rect 5663 1050 5667 1054
rect 1975 1002 1979 1006
rect 2023 1002 2027 1006
rect 2191 1002 2195 1006
rect 2199 1002 2203 1006
rect 2375 1002 2379 1006
rect 2391 1002 2395 1006
rect 2567 1002 2571 1006
rect 2575 1002 2579 1006
rect 2751 1002 2755 1006
rect 2759 1002 2763 1006
rect 2919 1002 2923 1006
rect 2943 1002 2947 1006
rect 3087 1002 3091 1006
rect 3127 1002 3131 1006
rect 3247 1002 3251 1006
rect 3311 1002 3315 1006
rect 3415 1002 3419 1006
rect 3495 1002 3499 1006
rect 3679 1002 3683 1006
rect 3799 1002 3803 1006
rect 111 946 115 950
rect 147 946 151 950
rect 235 946 239 950
rect 403 946 407 950
rect 459 946 463 950
rect 659 946 663 950
rect 683 946 687 950
rect 907 946 911 950
rect 923 946 927 950
rect 1131 946 1135 950
rect 1187 946 1191 950
rect 1363 946 1367 950
rect 1935 946 1939 950
rect 3839 934 3843 938
rect 3859 934 3863 938
rect 3995 934 3999 938
rect 4171 934 4175 938
rect 4387 934 4391 938
rect 4643 934 4647 938
rect 4779 934 4783 938
rect 4915 934 4919 938
rect 4931 934 4935 938
rect 5051 934 5055 938
rect 5187 934 5191 938
rect 5235 934 5239 938
rect 5323 934 5327 938
rect 5459 934 5463 938
rect 5515 934 5519 938
rect 5663 934 5667 938
rect 1975 886 1979 890
rect 1995 886 1999 890
rect 2163 886 2167 890
rect 2179 886 2183 890
rect 2347 886 2351 890
rect 2403 886 2407 890
rect 2539 886 2543 890
rect 2675 886 2679 890
rect 2731 886 2735 890
rect 2915 886 2919 890
rect 2987 886 2991 890
rect 3099 886 3103 890
rect 3283 886 3287 890
rect 3323 886 3327 890
rect 3467 886 3471 890
rect 3651 886 3655 890
rect 3799 886 3803 890
rect 111 818 115 822
rect 175 818 179 822
rect 263 818 267 822
rect 431 818 435 822
rect 487 818 491 822
rect 671 818 675 822
rect 711 818 715 822
rect 903 818 907 822
rect 935 818 939 822
rect 1127 818 1131 822
rect 1159 818 1163 822
rect 1351 818 1355 822
rect 1391 818 1395 822
rect 1575 818 1579 822
rect 1935 818 1939 822
rect 3839 822 3843 826
rect 3887 822 3891 826
rect 4023 822 4027 826
rect 4159 822 4163 826
rect 4199 822 4203 826
rect 4295 822 4299 826
rect 4415 822 4419 826
rect 4431 822 4435 826
rect 4567 822 4571 826
rect 4671 822 4675 826
rect 4719 822 4723 826
rect 4895 822 4899 826
rect 4959 822 4963 826
rect 5087 822 5091 826
rect 5263 822 5267 826
rect 5287 822 5291 826
rect 5487 822 5491 826
rect 5543 822 5547 826
rect 5663 822 5667 826
rect 111 706 115 710
rect 131 706 135 710
rect 147 706 151 710
rect 315 706 319 710
rect 403 706 407 710
rect 523 706 527 710
rect 643 706 647 710
rect 723 706 727 710
rect 875 706 879 710
rect 907 706 911 710
rect 1083 706 1087 710
rect 1099 706 1103 710
rect 1259 706 1263 710
rect 1323 706 1327 710
rect 1427 706 1431 710
rect 1547 706 1551 710
rect 1595 706 1599 710
rect 1771 706 1775 710
rect 1935 706 1939 710
rect 111 594 115 598
rect 159 594 163 598
rect 343 594 347 598
rect 375 594 379 598
rect 551 594 555 598
rect 599 594 603 598
rect 751 594 755 598
rect 807 594 811 598
rect 935 594 939 598
rect 999 594 1003 598
rect 1111 594 1115 598
rect 1175 594 1179 598
rect 1287 594 1291 598
rect 1343 594 1347 598
rect 1455 594 1459 598
rect 1511 594 1515 598
rect 1623 594 1627 598
rect 1671 594 1675 598
rect 1799 594 1803 598
rect 1815 594 1819 598
rect 1935 594 1939 598
rect 3839 706 3843 710
rect 3859 706 3863 710
rect 3995 706 3999 710
rect 4131 706 4135 710
rect 4267 706 4271 710
rect 4403 706 4407 710
rect 4539 706 4543 710
rect 4691 706 4695 710
rect 4699 706 4703 710
rect 4867 706 4871 710
rect 4891 706 4895 710
rect 5059 706 5063 710
rect 5099 706 5103 710
rect 5259 706 5263 710
rect 5315 706 5319 710
rect 5459 706 5463 710
rect 5515 706 5519 710
rect 5663 706 5667 710
rect 3839 594 3843 598
rect 3887 594 3891 598
rect 4023 594 4027 598
rect 4071 594 4075 598
rect 4159 594 4163 598
rect 4295 594 4299 598
rect 4311 594 4315 598
rect 4431 594 4435 598
rect 4567 594 4571 598
rect 4575 594 4579 598
rect 4727 594 4731 598
rect 4855 594 4859 598
rect 4919 594 4923 598
rect 5127 594 5131 598
rect 5151 594 5155 598
rect 5343 594 5347 598
rect 5447 594 5451 598
rect 5543 594 5547 598
rect 5663 594 5667 598
rect 1975 574 1979 578
rect 2023 574 2027 578
rect 2207 574 2211 578
rect 2431 574 2435 578
rect 2703 574 2707 578
rect 3015 574 3019 578
rect 3135 574 3139 578
rect 3271 574 3275 578
rect 3351 574 3355 578
rect 3407 574 3411 578
rect 3543 574 3547 578
rect 3679 574 3683 578
rect 3799 574 3803 578
rect 111 482 115 486
rect 131 482 135 486
rect 155 482 159 486
rect 347 482 351 486
rect 483 482 487 486
rect 571 482 575 486
rect 779 482 783 486
rect 811 482 815 486
rect 971 482 975 486
rect 1139 482 1143 486
rect 1147 482 1151 486
rect 1315 482 1319 486
rect 1475 482 1479 486
rect 1483 482 1487 486
rect 1643 482 1647 486
rect 1787 482 1791 486
rect 1935 482 1939 486
rect 3839 470 3843 474
rect 3859 470 3863 474
rect 4043 470 4047 474
rect 4283 470 4287 474
rect 4451 470 4455 474
rect 4547 470 4551 474
rect 4643 470 4647 474
rect 4827 470 4831 474
rect 4843 470 4847 474
rect 5051 470 5055 474
rect 5123 470 5127 474
rect 5267 470 5271 474
rect 5419 470 5423 474
rect 5483 470 5487 474
rect 5663 470 5667 474
rect 1975 462 1979 466
rect 1995 462 1999 466
rect 2203 462 2207 466
rect 2427 462 2431 466
rect 2651 462 2655 466
rect 2859 462 2863 466
rect 3067 462 3071 466
rect 3107 462 3111 466
rect 3243 462 3247 466
rect 3267 462 3271 466
rect 3379 462 3383 466
rect 3467 462 3471 466
rect 3515 462 3519 466
rect 3651 462 3655 466
rect 3799 462 3803 466
rect 111 358 115 362
rect 183 358 187 362
rect 279 358 283 362
rect 487 358 491 362
rect 511 358 515 362
rect 703 358 707 362
rect 839 358 843 362
rect 919 358 923 362
rect 1135 358 1139 362
rect 1167 358 1171 362
rect 1503 358 1507 362
rect 1815 358 1819 362
rect 1935 358 1939 362
rect 3839 354 3843 358
rect 4479 354 4483 358
rect 4615 354 4619 358
rect 4671 354 4675 358
rect 4775 354 4779 358
rect 4871 354 4875 358
rect 4951 354 4955 358
rect 5079 354 5083 358
rect 5135 354 5139 358
rect 5295 354 5299 358
rect 5327 354 5331 358
rect 5511 354 5515 358
rect 5527 354 5531 358
rect 5663 354 5667 358
rect 1975 334 1979 338
rect 2023 334 2027 338
rect 2159 334 2163 338
rect 2231 334 2235 338
rect 2295 334 2299 338
rect 2431 334 2435 338
rect 2455 334 2459 338
rect 2567 334 2571 338
rect 2679 334 2683 338
rect 2703 334 2707 338
rect 2839 334 2843 338
rect 2887 334 2891 338
rect 2975 334 2979 338
rect 3095 334 3099 338
rect 3111 334 3115 338
rect 3247 334 3251 338
rect 3295 334 3299 338
rect 3383 334 3387 338
rect 3495 334 3499 338
rect 3519 334 3523 338
rect 3655 334 3659 338
rect 3679 334 3683 338
rect 3799 334 3803 338
rect 111 206 115 210
rect 131 206 135 210
rect 251 206 255 210
rect 267 206 271 210
rect 403 206 407 210
rect 459 206 463 210
rect 539 206 543 210
rect 675 206 679 210
rect 811 206 815 210
rect 891 206 895 210
rect 947 206 951 210
rect 1083 206 1087 210
rect 1107 206 1111 210
rect 1935 206 1939 210
rect 3839 202 3843 206
rect 4291 202 4295 206
rect 4427 202 4431 206
rect 4563 202 4567 206
rect 4587 202 4591 206
rect 4699 202 4703 206
rect 4747 202 4751 206
rect 4835 202 4839 206
rect 4923 202 4927 206
rect 4971 202 4975 206
rect 5107 202 5111 206
rect 5243 202 5247 206
rect 5299 202 5303 206
rect 5379 202 5383 206
rect 5499 202 5503 206
rect 5515 202 5519 206
rect 5663 202 5667 206
rect 1975 186 1979 190
rect 1995 186 1999 190
rect 2131 186 2135 190
rect 2267 186 2271 190
rect 2403 186 2407 190
rect 2539 186 2543 190
rect 2675 186 2679 190
rect 2811 186 2815 190
rect 2947 186 2951 190
rect 3083 186 3087 190
rect 3219 186 3223 190
rect 3355 186 3359 190
rect 3491 186 3495 190
rect 3627 186 3631 190
rect 3799 186 3803 190
rect 111 94 115 98
rect 159 94 163 98
rect 295 94 299 98
rect 431 94 435 98
rect 567 94 571 98
rect 703 94 707 98
rect 839 94 843 98
rect 975 94 979 98
rect 1111 94 1115 98
rect 1935 94 1939 98
rect 3839 90 3843 94
rect 4319 90 4323 94
rect 4455 90 4459 94
rect 4591 90 4595 94
rect 4727 90 4731 94
rect 4863 90 4867 94
rect 4999 90 5003 94
rect 5135 90 5139 94
rect 5271 90 5275 94
rect 5407 90 5411 94
rect 5543 90 5547 94
rect 5663 90 5667 94
rect 1975 74 1979 78
rect 2023 74 2027 78
rect 2159 74 2163 78
rect 2295 74 2299 78
rect 2431 74 2435 78
rect 2567 74 2571 78
rect 2703 74 2707 78
rect 2839 74 2843 78
rect 2975 74 2979 78
rect 3111 74 3115 78
rect 3247 74 3251 78
rect 3383 74 3387 78
rect 3519 74 3523 78
rect 3655 74 3659 78
rect 3799 74 3803 78
<< m4 >>
rect 84 5753 85 5759
rect 91 5758 1947 5759
rect 91 5754 111 5758
rect 115 5754 159 5758
rect 163 5754 295 5758
rect 299 5754 1935 5758
rect 1939 5754 1947 5758
rect 91 5753 1947 5754
rect 1953 5753 1954 5759
rect 1946 5653 1947 5659
rect 1953 5658 3811 5659
rect 1953 5654 1975 5658
rect 1979 5654 2023 5658
rect 2027 5654 2183 5658
rect 2187 5654 2367 5658
rect 2371 5654 2551 5658
rect 2555 5654 2727 5658
rect 2731 5654 2895 5658
rect 2899 5654 3063 5658
rect 3067 5654 3223 5658
rect 3227 5654 3383 5658
rect 3387 5654 3543 5658
rect 3547 5654 3679 5658
rect 3683 5654 3799 5658
rect 3803 5654 3811 5658
rect 1953 5653 3811 5654
rect 3817 5655 3818 5659
rect 3817 5654 5702 5655
rect 3817 5653 3839 5654
rect 3810 5650 3839 5653
rect 3843 5650 4335 5654
rect 4339 5650 4471 5654
rect 4475 5650 4607 5654
rect 4611 5650 4743 5654
rect 4747 5650 4879 5654
rect 4883 5650 5015 5654
rect 5019 5650 5663 5654
rect 5667 5650 5702 5654
rect 3810 5649 5702 5650
rect 96 5641 97 5647
rect 103 5646 1959 5647
rect 103 5642 111 5646
rect 115 5642 131 5646
rect 135 5642 267 5646
rect 271 5642 275 5646
rect 279 5642 475 5646
rect 479 5642 699 5646
rect 703 5642 955 5646
rect 959 5642 1227 5646
rect 1231 5642 1515 5646
rect 1519 5642 1787 5646
rect 1791 5642 1935 5646
rect 1939 5642 1959 5646
rect 103 5641 1959 5642
rect 1965 5641 1966 5647
rect 1958 5541 1959 5547
rect 1965 5546 3823 5547
rect 1965 5542 1975 5546
rect 1979 5542 1995 5546
rect 1999 5542 2139 5546
rect 2143 5542 2155 5546
rect 2159 5542 2339 5546
rect 2343 5542 2355 5546
rect 2359 5542 2523 5546
rect 2527 5542 2563 5546
rect 2567 5542 2699 5546
rect 2703 5542 2755 5546
rect 2759 5542 2867 5546
rect 2871 5542 2939 5546
rect 2943 5542 3035 5546
rect 3039 5542 3115 5546
rect 3119 5542 3195 5546
rect 3199 5542 3291 5546
rect 3295 5542 3355 5546
rect 3359 5542 3467 5546
rect 3471 5542 3515 5546
rect 3519 5542 3643 5546
rect 3647 5542 3651 5546
rect 3655 5542 3799 5546
rect 3803 5542 3823 5546
rect 1965 5541 3823 5542
rect 3829 5543 3830 5547
rect 3829 5542 5714 5543
rect 3829 5541 3839 5542
rect 3822 5538 3839 5541
rect 3843 5538 4251 5542
rect 4255 5538 4307 5542
rect 4311 5538 4403 5542
rect 4407 5538 4443 5542
rect 4447 5538 4555 5542
rect 4559 5538 4579 5542
rect 4583 5538 4707 5542
rect 4711 5538 4715 5542
rect 4719 5538 4851 5542
rect 4855 5538 4859 5542
rect 4863 5538 4987 5542
rect 4991 5538 5019 5542
rect 5023 5538 5663 5542
rect 5667 5538 5714 5542
rect 3822 5537 5714 5538
rect 84 5529 85 5535
rect 91 5534 1947 5535
rect 91 5530 111 5534
rect 115 5530 159 5534
rect 163 5530 279 5534
rect 283 5530 303 5534
rect 307 5530 503 5534
rect 507 5530 519 5534
rect 523 5530 727 5534
rect 731 5530 767 5534
rect 771 5530 983 5534
rect 987 5530 1015 5534
rect 1019 5530 1255 5534
rect 1259 5530 1263 5534
rect 1267 5530 1511 5534
rect 1515 5530 1543 5534
rect 1547 5530 1767 5534
rect 1771 5530 1815 5534
rect 1819 5530 1935 5534
rect 1939 5530 1947 5534
rect 91 5529 1947 5530
rect 1953 5529 1954 5535
rect 1946 5427 1947 5433
rect 1953 5427 1978 5433
rect 1972 5426 3811 5427
rect 96 5417 97 5423
rect 103 5422 1959 5423
rect 103 5418 111 5422
rect 115 5418 251 5422
rect 255 5418 411 5422
rect 415 5418 491 5422
rect 495 5418 611 5422
rect 615 5418 739 5422
rect 743 5418 819 5422
rect 823 5418 987 5422
rect 991 5418 1035 5422
rect 1039 5418 1235 5422
rect 1239 5418 1259 5422
rect 1263 5418 1483 5422
rect 1487 5418 1491 5422
rect 1495 5418 1739 5422
rect 1743 5418 1935 5422
rect 1939 5418 1959 5422
rect 103 5417 1959 5418
rect 1965 5417 1966 5423
rect 1972 5422 1975 5426
rect 1979 5422 2167 5426
rect 2171 5422 2311 5426
rect 2315 5422 2383 5426
rect 2387 5422 2511 5426
rect 2515 5422 2591 5426
rect 2595 5422 2703 5426
rect 2707 5422 2783 5426
rect 2787 5422 2887 5426
rect 2891 5422 2967 5426
rect 2971 5422 3071 5426
rect 3075 5422 3143 5426
rect 3147 5422 3247 5426
rect 3251 5422 3319 5426
rect 3323 5422 3423 5426
rect 3427 5422 3495 5426
rect 3499 5422 3607 5426
rect 3611 5422 3671 5426
rect 3675 5422 3799 5426
rect 3803 5422 3811 5426
rect 1972 5421 3811 5422
rect 3817 5421 3818 5427
rect 3810 5405 3811 5411
rect 3817 5410 5695 5411
rect 3817 5406 3839 5410
rect 3843 5406 4279 5410
rect 4283 5406 4431 5410
rect 4435 5406 4487 5410
rect 4491 5406 4583 5410
rect 4587 5406 4695 5410
rect 4699 5406 4735 5410
rect 4739 5406 4887 5410
rect 4891 5406 4911 5410
rect 4915 5406 5047 5410
rect 5051 5406 5127 5410
rect 5131 5406 5663 5410
rect 5667 5406 5695 5410
rect 3817 5405 5695 5406
rect 5701 5405 5702 5411
rect 84 5305 85 5311
rect 91 5310 1947 5311
rect 91 5306 111 5310
rect 115 5306 439 5310
rect 443 5306 591 5310
rect 595 5306 639 5310
rect 643 5306 727 5310
rect 731 5306 847 5310
rect 851 5306 863 5310
rect 867 5306 999 5310
rect 1003 5306 1063 5310
rect 1067 5306 1135 5310
rect 1139 5306 1271 5310
rect 1275 5306 1287 5310
rect 1291 5306 1407 5310
rect 1411 5306 1519 5310
rect 1523 5306 1543 5310
rect 1547 5306 1935 5310
rect 1939 5306 1947 5310
rect 91 5305 1947 5306
rect 1953 5305 1954 5311
rect 1958 5309 1959 5315
rect 1965 5314 3823 5315
rect 1965 5310 1975 5314
rect 1979 5310 2195 5314
rect 2199 5310 2283 5314
rect 2287 5310 2339 5314
rect 2343 5310 2483 5314
rect 2487 5310 2491 5314
rect 2495 5310 2651 5314
rect 2655 5310 2675 5314
rect 2679 5310 2819 5314
rect 2823 5310 2859 5314
rect 2863 5310 3003 5314
rect 3007 5310 3043 5314
rect 3047 5310 3187 5314
rect 3191 5310 3219 5314
rect 3223 5310 3379 5314
rect 3383 5310 3395 5314
rect 3399 5310 3579 5314
rect 3583 5310 3799 5314
rect 3803 5310 3823 5314
rect 1965 5309 3823 5310
rect 3829 5309 3830 5315
rect 3822 5277 3823 5283
rect 3829 5282 5707 5283
rect 3829 5278 3839 5282
rect 3843 5278 4251 5282
rect 4255 5278 4459 5282
rect 4463 5278 4483 5282
rect 4487 5278 4667 5282
rect 4671 5278 4715 5282
rect 4719 5278 4883 5282
rect 4887 5278 4947 5282
rect 4951 5278 5099 5282
rect 5103 5278 5187 5282
rect 5191 5278 5663 5282
rect 5667 5278 5707 5282
rect 3829 5277 5707 5278
rect 5713 5277 5714 5283
rect 1946 5197 1947 5203
rect 1953 5202 3811 5203
rect 1953 5198 1975 5202
rect 1979 5198 2023 5202
rect 2027 5198 2159 5202
rect 2163 5198 2223 5202
rect 2227 5198 2327 5202
rect 2331 5198 2367 5202
rect 2371 5198 2511 5202
rect 2515 5198 2519 5202
rect 2523 5198 2679 5202
rect 2683 5198 2695 5202
rect 2699 5198 2847 5202
rect 2851 5198 2887 5202
rect 2891 5198 3031 5202
rect 3035 5198 3087 5202
rect 3091 5198 3215 5202
rect 3219 5198 3287 5202
rect 3291 5198 3407 5202
rect 3411 5198 3495 5202
rect 3499 5198 3607 5202
rect 3611 5198 3679 5202
rect 3683 5198 3799 5202
rect 3803 5198 3811 5202
rect 1953 5197 3811 5198
rect 3817 5197 3818 5203
rect 3810 5137 3811 5143
rect 3817 5142 5695 5143
rect 3817 5138 3839 5142
rect 3843 5138 3887 5142
rect 3891 5138 4135 5142
rect 4139 5138 4279 5142
rect 4283 5138 4407 5142
rect 4411 5138 4511 5142
rect 4515 5138 4679 5142
rect 4683 5138 4743 5142
rect 4747 5138 4959 5142
rect 4963 5138 4975 5142
rect 4979 5138 5215 5142
rect 5219 5138 5239 5142
rect 5243 5138 5663 5142
rect 5667 5138 5695 5142
rect 3817 5137 5695 5138
rect 5701 5137 5702 5143
rect 96 5089 97 5095
rect 103 5094 1959 5095
rect 103 5090 111 5094
rect 115 5090 347 5094
rect 351 5090 483 5094
rect 487 5090 563 5094
rect 567 5090 619 5094
rect 623 5090 699 5094
rect 703 5090 755 5094
rect 759 5090 835 5094
rect 839 5090 891 5094
rect 895 5090 971 5094
rect 975 5090 1035 5094
rect 1039 5090 1107 5094
rect 1111 5090 1187 5094
rect 1191 5090 1243 5094
rect 1247 5090 1339 5094
rect 1343 5090 1379 5094
rect 1383 5090 1491 5094
rect 1495 5090 1515 5094
rect 1519 5090 1651 5094
rect 1655 5090 1787 5094
rect 1791 5090 1935 5094
rect 1939 5090 1959 5094
rect 103 5089 1959 5090
rect 1965 5091 1966 5095
rect 1965 5090 3830 5091
rect 1965 5089 1975 5090
rect 1958 5086 1975 5089
rect 1979 5086 1995 5090
rect 1999 5086 2131 5090
rect 2135 5086 2299 5090
rect 2303 5086 2483 5090
rect 2487 5086 2531 5090
rect 2535 5086 2667 5090
rect 2671 5086 2859 5090
rect 2863 5086 3059 5090
rect 3063 5086 3099 5090
rect 3103 5086 3259 5090
rect 3263 5086 3467 5090
rect 3471 5086 3651 5090
rect 3655 5086 3799 5090
rect 3803 5086 3830 5090
rect 1958 5085 3830 5086
rect 3822 5013 3823 5019
rect 3829 5018 5707 5019
rect 3829 5014 3839 5018
rect 3843 5014 3859 5018
rect 3863 5014 4019 5018
rect 4023 5014 4107 5018
rect 4111 5014 4211 5018
rect 4215 5014 4379 5018
rect 4383 5014 4411 5018
rect 4415 5014 4627 5018
rect 4631 5014 4651 5018
rect 4655 5014 4843 5018
rect 4847 5014 4931 5018
rect 4935 5014 5067 5018
rect 5071 5014 5211 5018
rect 5215 5014 5299 5018
rect 5303 5014 5663 5018
rect 5667 5014 5707 5018
rect 3829 5013 5707 5014
rect 5713 5013 5714 5019
rect 84 4977 85 4983
rect 91 4982 1947 4983
rect 91 4978 111 4982
rect 115 4978 159 4982
rect 163 4978 343 4982
rect 347 4978 375 4982
rect 379 4978 511 4982
rect 515 4978 551 4982
rect 555 4978 647 4982
rect 651 4978 751 4982
rect 755 4978 783 4982
rect 787 4978 919 4982
rect 923 4978 943 4982
rect 947 4978 1063 4982
rect 1067 4978 1127 4982
rect 1131 4978 1215 4982
rect 1219 4978 1311 4982
rect 1315 4978 1367 4982
rect 1371 4978 1487 4982
rect 1491 4978 1519 4982
rect 1523 4978 1663 4982
rect 1667 4978 1679 4982
rect 1683 4978 1815 4982
rect 1819 4978 1935 4982
rect 1939 4978 1947 4982
rect 91 4977 1947 4978
rect 1953 4977 1954 4983
rect 1946 4941 1947 4947
rect 1953 4946 3811 4947
rect 1953 4942 1975 4946
rect 1979 4942 2023 4946
rect 2027 4942 2559 4946
rect 2563 4942 2871 4946
rect 2875 4942 3007 4946
rect 3011 4942 3127 4946
rect 3131 4942 3679 4946
rect 3683 4942 3799 4946
rect 3803 4942 3811 4946
rect 1953 4941 3811 4942
rect 3817 4941 3818 4947
rect 3810 4881 3811 4887
rect 3817 4886 5695 4887
rect 3817 4882 3839 4886
rect 3843 4882 3887 4886
rect 3891 4882 4047 4886
rect 4051 4882 4071 4886
rect 4075 4882 4239 4886
rect 4243 4882 4287 4886
rect 4291 4882 4439 4886
rect 4443 4882 4511 4886
rect 4515 4882 4655 4886
rect 4659 4882 4735 4886
rect 4739 4882 4871 4886
rect 4875 4882 4959 4886
rect 4963 4882 5095 4886
rect 5099 4882 5183 4886
rect 5187 4882 5327 4886
rect 5331 4882 5407 4886
rect 5411 4882 5663 4886
rect 5667 4882 5695 4886
rect 3817 4881 5695 4882
rect 5701 4881 5702 4887
rect 96 4857 97 4863
rect 103 4862 1959 4863
rect 103 4858 111 4862
rect 115 4858 131 4862
rect 135 4858 267 4862
rect 271 4858 315 4862
rect 319 4858 403 4862
rect 407 4858 523 4862
rect 527 4858 539 4862
rect 543 4858 675 4862
rect 679 4858 723 4862
rect 727 4858 915 4862
rect 919 4858 1099 4862
rect 1103 4858 1283 4862
rect 1287 4858 1459 4862
rect 1463 4858 1635 4862
rect 1639 4858 1787 4862
rect 1791 4858 1935 4862
rect 1939 4858 1959 4862
rect 103 4857 1959 4858
rect 1965 4857 1966 4863
rect 1958 4805 1959 4811
rect 1965 4810 3823 4811
rect 1965 4806 1975 4810
rect 1979 4806 1995 4810
rect 1999 4806 2155 4810
rect 2159 4806 2347 4810
rect 2351 4806 2539 4810
rect 2543 4806 2731 4810
rect 2735 4806 2843 4810
rect 2847 4806 2931 4810
rect 2935 4806 2979 4810
rect 2983 4806 3131 4810
rect 3135 4806 3799 4810
rect 3803 4806 3823 4810
rect 1965 4805 3823 4806
rect 3829 4805 3830 4811
rect 3822 4765 3823 4771
rect 3829 4770 5707 4771
rect 3829 4766 3839 4770
rect 3843 4766 3859 4770
rect 3863 4766 3915 4770
rect 3919 4766 4043 4770
rect 4047 4766 4187 4770
rect 4191 4766 4259 4770
rect 4263 4766 4467 4770
rect 4471 4766 4483 4770
rect 4487 4766 4707 4770
rect 4711 4766 4763 4770
rect 4767 4766 4931 4770
rect 4935 4766 5067 4770
rect 5071 4766 5155 4770
rect 5159 4766 5371 4770
rect 5375 4766 5379 4770
rect 5383 4766 5663 4770
rect 5667 4766 5707 4770
rect 3829 4765 5707 4766
rect 5713 4765 5714 4771
rect 84 4737 85 4743
rect 91 4742 1947 4743
rect 91 4738 111 4742
rect 115 4738 159 4742
rect 163 4738 295 4742
rect 299 4738 343 4742
rect 347 4738 431 4742
rect 435 4738 567 4742
rect 571 4738 703 4742
rect 707 4738 807 4742
rect 811 4738 1055 4742
rect 1059 4738 1311 4742
rect 1315 4738 1575 4742
rect 1579 4738 1815 4742
rect 1819 4738 1935 4742
rect 1939 4738 1947 4742
rect 91 4737 1947 4738
rect 1953 4737 1954 4743
rect 1946 4689 1947 4695
rect 1953 4694 3811 4695
rect 1953 4690 1975 4694
rect 1979 4690 2023 4694
rect 2027 4690 2183 4694
rect 2187 4690 2239 4694
rect 2243 4690 2375 4694
rect 2379 4690 2471 4694
rect 2475 4690 2567 4694
rect 2571 4690 2695 4694
rect 2699 4690 2759 4694
rect 2763 4690 2919 4694
rect 2923 4690 2959 4694
rect 2963 4690 3143 4694
rect 3147 4690 3159 4694
rect 3163 4690 3367 4694
rect 3371 4690 3799 4694
rect 3803 4690 3811 4694
rect 1953 4689 3811 4690
rect 3817 4689 3818 4695
rect 3810 4653 3811 4659
rect 3817 4658 5695 4659
rect 3817 4654 3839 4658
rect 3843 4654 3943 4658
rect 3947 4654 4063 4658
rect 4067 4654 4215 4658
rect 4219 4654 4327 4658
rect 4331 4654 4495 4658
rect 4499 4654 4599 4658
rect 4603 4654 4791 4658
rect 4795 4654 4871 4658
rect 4875 4654 5095 4658
rect 5099 4654 5151 4658
rect 5155 4654 5399 4658
rect 5403 4654 5439 4658
rect 5443 4654 5663 4658
rect 5667 4654 5695 4658
rect 3817 4653 5695 4654
rect 5701 4653 5702 4659
rect 96 4609 97 4615
rect 103 4614 1959 4615
rect 103 4610 111 4614
rect 115 4610 131 4614
rect 135 4610 171 4614
rect 175 4610 315 4614
rect 319 4610 395 4614
rect 399 4610 539 4614
rect 543 4610 643 4614
rect 647 4610 779 4614
rect 783 4610 907 4614
rect 911 4610 1027 4614
rect 1031 4610 1195 4614
rect 1199 4610 1283 4614
rect 1287 4610 1491 4614
rect 1495 4610 1547 4614
rect 1551 4610 1787 4614
rect 1791 4610 1935 4614
rect 1939 4610 1959 4614
rect 103 4609 1959 4610
rect 1965 4609 1966 4615
rect 1958 4573 1959 4579
rect 1965 4578 3823 4579
rect 1965 4574 1975 4578
rect 1979 4574 1995 4578
rect 1999 4574 2099 4578
rect 2103 4574 2211 4578
rect 2215 4574 2347 4578
rect 2351 4574 2443 4578
rect 2447 4574 2579 4578
rect 2583 4574 2667 4578
rect 2671 4574 2795 4578
rect 2799 4574 2891 4578
rect 2895 4574 3003 4578
rect 3007 4574 3115 4578
rect 3119 4574 3203 4578
rect 3207 4574 3339 4578
rect 3343 4574 3403 4578
rect 3407 4574 3611 4578
rect 3615 4574 3799 4578
rect 3803 4574 3823 4578
rect 1965 4573 3823 4574
rect 3829 4573 3830 4579
rect 3822 4541 3823 4547
rect 3829 4546 5707 4547
rect 3829 4542 3839 4546
rect 3843 4542 4035 4546
rect 4039 4542 4179 4546
rect 4183 4542 4299 4546
rect 4303 4542 4411 4546
rect 4415 4542 4571 4546
rect 4575 4542 4659 4546
rect 4663 4542 4843 4546
rect 4847 4542 4915 4546
rect 4919 4542 5123 4546
rect 5127 4542 5179 4546
rect 5183 4542 5411 4546
rect 5415 4542 5443 4546
rect 5447 4542 5663 4546
rect 5667 4542 5707 4546
rect 3829 4541 5707 4542
rect 5713 4541 5714 4547
rect 84 4493 85 4499
rect 91 4498 1947 4499
rect 91 4494 111 4498
rect 115 4494 199 4498
rect 203 4494 423 4498
rect 427 4494 447 4498
rect 451 4494 655 4498
rect 659 4494 671 4498
rect 675 4494 887 4498
rect 891 4494 935 4498
rect 939 4494 1143 4498
rect 1147 4494 1223 4498
rect 1227 4494 1407 4498
rect 1411 4494 1519 4498
rect 1523 4494 1679 4498
rect 1683 4494 1815 4498
rect 1819 4494 1935 4498
rect 1939 4494 1947 4498
rect 91 4493 1947 4494
rect 1953 4493 1954 4499
rect 1946 4453 1947 4459
rect 1953 4458 3811 4459
rect 1953 4454 1975 4458
rect 1979 4454 2127 4458
rect 2131 4454 2231 4458
rect 2235 4454 2375 4458
rect 2379 4454 2447 4458
rect 2451 4454 2607 4458
rect 2611 4454 2663 4458
rect 2667 4454 2823 4458
rect 2827 4454 2871 4458
rect 2875 4454 3031 4458
rect 3035 4454 3079 4458
rect 3083 4454 3231 4458
rect 3235 4454 3287 4458
rect 3291 4454 3431 4458
rect 3435 4454 3495 4458
rect 3499 4454 3639 4458
rect 3643 4454 3679 4458
rect 3683 4454 3799 4458
rect 3803 4454 3811 4458
rect 1953 4453 3811 4454
rect 3817 4453 3818 4459
rect 3810 4421 3811 4427
rect 3817 4426 5695 4427
rect 3817 4422 3839 4426
rect 3843 4422 4207 4426
rect 4211 4422 4359 4426
rect 4363 4422 4439 4426
rect 4443 4422 4519 4426
rect 4523 4422 4687 4426
rect 4691 4422 4879 4426
rect 4883 4422 4943 4426
rect 4947 4422 5079 4426
rect 5083 4422 5207 4426
rect 5211 4422 5287 4426
rect 5291 4422 5471 4426
rect 5475 4422 5503 4426
rect 5507 4422 5663 4426
rect 5667 4422 5695 4426
rect 3817 4421 5695 4422
rect 5701 4421 5702 4427
rect 96 4377 97 4383
rect 103 4382 1959 4383
rect 103 4378 111 4382
rect 115 4378 419 4382
rect 423 4378 627 4382
rect 631 4378 667 4382
rect 671 4378 811 4382
rect 815 4378 859 4382
rect 863 4378 963 4382
rect 967 4378 1115 4382
rect 1119 4378 1123 4382
rect 1127 4378 1291 4382
rect 1295 4378 1379 4382
rect 1383 4378 1467 4382
rect 1471 4378 1651 4382
rect 1655 4378 1935 4382
rect 1939 4378 1959 4382
rect 103 4377 1959 4378
rect 1965 4377 1966 4383
rect 1958 4333 1959 4339
rect 1965 4338 3823 4339
rect 1965 4334 1975 4338
rect 1979 4334 2203 4338
rect 2207 4334 2307 4338
rect 2311 4334 2419 4338
rect 2423 4334 2459 4338
rect 2463 4334 2627 4338
rect 2631 4334 2635 4338
rect 2639 4334 2811 4338
rect 2815 4334 2843 4338
rect 2847 4334 3011 4338
rect 3015 4334 3051 4338
rect 3055 4334 3227 4338
rect 3231 4334 3259 4338
rect 3263 4334 3451 4338
rect 3455 4334 3467 4338
rect 3471 4334 3651 4338
rect 3655 4334 3799 4338
rect 3803 4334 3823 4338
rect 1965 4333 3823 4334
rect 3829 4333 3830 4339
rect 3822 4309 3823 4315
rect 3829 4314 5707 4315
rect 3829 4310 3839 4314
rect 3843 4310 3859 4314
rect 3863 4310 4043 4314
rect 4047 4310 4251 4314
rect 4255 4310 4331 4314
rect 4335 4310 4475 4314
rect 4479 4310 4491 4314
rect 4495 4310 4659 4314
rect 4663 4310 4715 4314
rect 4719 4310 4851 4314
rect 4855 4310 4971 4314
rect 4975 4310 5051 4314
rect 5055 4310 5235 4314
rect 5239 4310 5259 4314
rect 5263 4310 5475 4314
rect 5479 4310 5499 4314
rect 5503 4310 5663 4314
rect 5667 4310 5707 4314
rect 3829 4309 5707 4310
rect 5713 4309 5714 4315
rect 84 4249 85 4255
rect 91 4254 1947 4255
rect 91 4250 111 4254
rect 115 4250 695 4254
rect 699 4250 815 4254
rect 819 4250 839 4254
rect 843 4250 951 4254
rect 955 4250 991 4254
rect 995 4250 1087 4254
rect 1091 4250 1151 4254
rect 1155 4250 1223 4254
rect 1227 4250 1319 4254
rect 1323 4250 1359 4254
rect 1363 4250 1495 4254
rect 1499 4250 1631 4254
rect 1635 4250 1679 4254
rect 1683 4250 1767 4254
rect 1771 4250 1935 4254
rect 1939 4250 1947 4254
rect 91 4249 1947 4250
rect 1953 4249 1954 4255
rect 1946 4213 1947 4219
rect 1953 4218 3811 4219
rect 1953 4214 1975 4218
rect 1979 4214 2335 4218
rect 2339 4214 2487 4218
rect 2491 4214 2567 4218
rect 2571 4214 2655 4218
rect 2659 4214 2703 4218
rect 2707 4214 2839 4218
rect 2843 4214 2975 4218
rect 2979 4214 3039 4218
rect 3043 4214 3255 4218
rect 3259 4214 3479 4218
rect 3483 4214 3679 4218
rect 3683 4214 3799 4218
rect 3803 4214 3811 4218
rect 1953 4213 3811 4214
rect 3817 4213 3818 4219
rect 3810 4161 3811 4167
rect 3817 4166 5695 4167
rect 3817 4162 3839 4166
rect 3843 4162 3887 4166
rect 3891 4162 4071 4166
rect 4075 4162 4279 4166
rect 4283 4162 4415 4166
rect 4419 4162 4503 4166
rect 4507 4162 4743 4166
rect 4747 4162 4975 4166
rect 4979 4162 4999 4166
rect 5003 4162 5263 4166
rect 5267 4162 5527 4166
rect 5531 4162 5543 4166
rect 5547 4162 5663 4166
rect 5667 4162 5695 4166
rect 3817 4161 5695 4162
rect 5701 4161 5702 4167
rect 96 4133 97 4139
rect 103 4138 1959 4139
rect 103 4134 111 4138
rect 115 4134 731 4138
rect 735 4134 787 4138
rect 791 4134 867 4138
rect 871 4134 923 4138
rect 927 4134 1003 4138
rect 1007 4134 1059 4138
rect 1063 4134 1139 4138
rect 1143 4134 1195 4138
rect 1199 4134 1275 4138
rect 1279 4134 1331 4138
rect 1335 4134 1411 4138
rect 1415 4134 1467 4138
rect 1471 4134 1547 4138
rect 1551 4134 1603 4138
rect 1607 4134 1739 4138
rect 1743 4134 1935 4138
rect 1939 4134 1959 4138
rect 103 4133 1959 4134
rect 1965 4133 1966 4139
rect 1958 4081 1959 4087
rect 1965 4086 3823 4087
rect 1965 4082 1975 4086
rect 1979 4082 2291 4086
rect 2295 4082 2427 4086
rect 2431 4082 2539 4086
rect 2543 4082 2563 4086
rect 2567 4082 2675 4086
rect 2679 4082 2699 4086
rect 2703 4082 2811 4086
rect 2815 4082 2835 4086
rect 2839 4082 2947 4086
rect 2951 4082 3799 4086
rect 3803 4082 3823 4086
rect 1965 4081 3823 4082
rect 3829 4081 3830 4087
rect 3822 4049 3823 4055
rect 3829 4054 5707 4055
rect 3829 4050 3839 4054
rect 3843 4050 3859 4054
rect 3863 4050 4003 4054
rect 4007 4050 4171 4054
rect 4175 4050 4339 4054
rect 4343 4050 4387 4054
rect 4391 4050 4499 4054
rect 4503 4050 4651 4054
rect 4655 4050 4803 4054
rect 4807 4050 4947 4054
rect 4951 4050 5091 4054
rect 5095 4050 5235 4054
rect 5239 4050 5379 4054
rect 5383 4050 5515 4054
rect 5519 4050 5663 4054
rect 5667 4050 5707 4054
rect 3829 4049 5707 4050
rect 5713 4049 5714 4055
rect 84 3997 85 4003
rect 91 4002 1947 4003
rect 91 3998 111 4002
rect 115 3998 511 4002
rect 515 3998 663 4002
rect 667 3998 759 4002
rect 763 3998 823 4002
rect 827 3998 895 4002
rect 899 3998 983 4002
rect 987 3998 1031 4002
rect 1035 3998 1151 4002
rect 1155 3998 1167 4002
rect 1171 3998 1303 4002
rect 1307 3998 1319 4002
rect 1323 3998 1439 4002
rect 1443 3998 1575 4002
rect 1579 3998 1935 4002
rect 1939 3998 1947 4002
rect 91 3997 1947 3998
rect 1953 3997 1954 4003
rect 1946 3965 1947 3971
rect 1953 3970 3811 3971
rect 1953 3966 1975 3970
rect 1979 3966 2119 3970
rect 2123 3966 2319 3970
rect 2323 3966 2327 3970
rect 2331 3966 2455 3970
rect 2459 3966 2535 3970
rect 2539 3966 2591 3970
rect 2595 3966 2727 3970
rect 2731 3966 2743 3970
rect 2747 3966 2863 3970
rect 2867 3966 2943 3970
rect 2947 3966 3135 3970
rect 3139 3966 3319 3970
rect 3323 3966 3511 3970
rect 3515 3966 3679 3970
rect 3683 3966 3799 3970
rect 3803 3966 3811 3970
rect 1953 3965 3811 3966
rect 3817 3965 3818 3971
rect 3810 3913 3811 3919
rect 3817 3918 5695 3919
rect 3817 3914 3839 3918
rect 3843 3914 3887 3918
rect 3891 3914 4031 3918
rect 4035 3914 4199 3918
rect 4203 3914 4367 3918
rect 4371 3914 4383 3918
rect 4387 3914 4527 3918
rect 4531 3914 4599 3918
rect 4603 3914 4679 3918
rect 4683 3914 4823 3918
rect 4827 3914 4831 3918
rect 4835 3914 4975 3918
rect 4979 3914 5063 3918
rect 5067 3914 5119 3918
rect 5123 3914 5263 3918
rect 5267 3914 5311 3918
rect 5315 3914 5407 3918
rect 5411 3914 5543 3918
rect 5547 3914 5663 3918
rect 5667 3914 5695 3918
rect 3817 3913 5695 3914
rect 5701 3913 5702 3919
rect 96 3857 97 3863
rect 103 3862 1959 3863
rect 103 3858 111 3862
rect 115 3858 131 3862
rect 135 3858 307 3862
rect 311 3858 483 3862
rect 487 3858 515 3862
rect 519 3858 635 3862
rect 639 3858 723 3862
rect 727 3858 795 3862
rect 799 3858 939 3862
rect 943 3858 955 3862
rect 959 3858 1123 3862
rect 1127 3858 1163 3862
rect 1167 3858 1291 3862
rect 1295 3858 1935 3862
rect 1939 3858 1959 3862
rect 103 3857 1959 3858
rect 1965 3857 1966 3863
rect 1958 3841 1959 3847
rect 1965 3846 3823 3847
rect 1965 3842 1975 3846
rect 1979 3842 2091 3846
rect 2095 3842 2139 3846
rect 2143 3842 2299 3846
rect 2303 3842 2371 3846
rect 2375 3842 2507 3846
rect 2511 3842 2587 3846
rect 2591 3842 2715 3846
rect 2719 3842 2795 3846
rect 2799 3842 2915 3846
rect 2919 3842 2995 3846
rect 2999 3842 3107 3846
rect 3111 3842 3195 3846
rect 3199 3842 3291 3846
rect 3295 3842 3403 3846
rect 3407 3842 3483 3846
rect 3487 3842 3651 3846
rect 3655 3842 3799 3846
rect 3803 3842 3823 3846
rect 1965 3841 3823 3842
rect 3829 3841 3830 3847
rect 3822 3785 3823 3791
rect 3829 3790 5707 3791
rect 3829 3786 3839 3790
rect 3843 3786 3995 3790
rect 3999 3786 4203 3790
rect 4207 3786 4355 3790
rect 4359 3786 4435 3790
rect 4439 3786 4571 3790
rect 4575 3786 4691 3790
rect 4695 3786 4795 3790
rect 4799 3786 4963 3790
rect 4967 3786 5035 3790
rect 5039 3786 5251 3790
rect 5255 3786 5283 3790
rect 5287 3786 5515 3790
rect 5519 3786 5663 3790
rect 5667 3786 5707 3790
rect 3829 3785 5707 3786
rect 5713 3785 5714 3791
rect 84 3745 85 3751
rect 91 3750 1947 3751
rect 91 3746 111 3750
rect 115 3746 159 3750
rect 163 3746 335 3750
rect 339 3746 527 3750
rect 531 3746 543 3750
rect 547 3746 711 3750
rect 715 3746 751 3750
rect 755 3746 887 3750
rect 891 3746 967 3750
rect 971 3746 1055 3750
rect 1059 3746 1191 3750
rect 1195 3746 1215 3750
rect 1219 3746 1367 3750
rect 1371 3746 1519 3750
rect 1523 3746 1679 3750
rect 1683 3746 1815 3750
rect 1819 3746 1935 3750
rect 1939 3746 1947 3750
rect 91 3745 1947 3746
rect 1953 3745 1954 3751
rect 1946 3725 1947 3731
rect 1953 3730 3811 3731
rect 1953 3726 1975 3730
rect 1979 3726 2167 3730
rect 2171 3726 2279 3730
rect 2283 3726 2399 3730
rect 2403 3726 2479 3730
rect 2483 3726 2615 3730
rect 2619 3726 2679 3730
rect 2683 3726 2823 3730
rect 2827 3726 2879 3730
rect 2883 3726 3023 3730
rect 3027 3726 3079 3730
rect 3083 3726 3223 3730
rect 3227 3726 3279 3730
rect 3283 3726 3431 3730
rect 3435 3726 3799 3730
rect 3803 3726 3811 3730
rect 1953 3725 3811 3726
rect 3817 3725 3818 3731
rect 3810 3645 3811 3651
rect 3817 3650 5695 3651
rect 3817 3646 3839 3650
rect 3843 3646 4023 3650
rect 4027 3646 4215 3650
rect 4219 3646 4231 3650
rect 4235 3646 4399 3650
rect 4403 3646 4463 3650
rect 4467 3646 4607 3650
rect 4611 3646 4719 3650
rect 4723 3646 4831 3650
rect 4835 3646 4991 3650
rect 4995 3646 5071 3650
rect 5075 3646 5279 3650
rect 5283 3646 5319 3650
rect 5323 3646 5543 3650
rect 5547 3646 5663 3650
rect 5667 3646 5695 3650
rect 3817 3645 5695 3646
rect 5701 3645 5702 3651
rect 96 3621 97 3627
rect 103 3626 1959 3627
rect 103 3622 111 3626
rect 115 3622 131 3626
rect 135 3622 147 3626
rect 151 3622 307 3626
rect 311 3622 355 3626
rect 359 3622 499 3626
rect 503 3622 571 3626
rect 575 3622 683 3626
rect 687 3622 803 3626
rect 807 3622 859 3626
rect 863 3622 1027 3626
rect 1031 3622 1043 3626
rect 1047 3622 1187 3626
rect 1191 3622 1291 3626
rect 1295 3622 1339 3626
rect 1343 3622 1491 3626
rect 1495 3622 1547 3626
rect 1551 3622 1651 3626
rect 1655 3622 1787 3626
rect 1791 3622 1935 3626
rect 1939 3622 1959 3626
rect 103 3621 1959 3622
rect 1965 3621 1966 3627
rect 1958 3601 1959 3607
rect 1965 3606 3823 3607
rect 1965 3602 1975 3606
rect 1979 3602 1995 3606
rect 1999 3602 2251 3606
rect 2255 3602 2451 3606
rect 2455 3602 2515 3606
rect 2519 3602 2651 3606
rect 2655 3602 2755 3606
rect 2759 3602 2851 3606
rect 2855 3602 2979 3606
rect 2983 3602 3051 3606
rect 3055 3602 3195 3606
rect 3199 3602 3251 3606
rect 3255 3602 3411 3606
rect 3415 3602 3627 3606
rect 3631 3602 3799 3606
rect 3803 3602 3823 3606
rect 1965 3601 3823 3602
rect 3829 3601 3830 3607
rect 3822 3509 3823 3515
rect 3829 3514 5707 3515
rect 3829 3510 3839 3514
rect 3843 3510 4187 3514
rect 4191 3510 4371 3514
rect 4375 3510 4531 3514
rect 4535 3510 4579 3514
rect 4583 3510 4683 3514
rect 4687 3510 4803 3514
rect 4807 3510 4843 3514
rect 4847 3510 5003 3514
rect 5007 3510 5043 3514
rect 5047 3510 5171 3514
rect 5175 3510 5291 3514
rect 5295 3510 5347 3514
rect 5351 3510 5515 3514
rect 5519 3510 5663 3514
rect 5667 3510 5707 3514
rect 3829 3509 5707 3510
rect 5713 3509 5714 3515
rect 84 3485 85 3491
rect 91 3490 1947 3491
rect 91 3486 111 3490
rect 115 3486 175 3490
rect 179 3486 303 3490
rect 307 3486 383 3490
rect 387 3486 447 3490
rect 451 3486 599 3490
rect 603 3486 759 3490
rect 763 3486 831 3490
rect 835 3486 935 3490
rect 939 3486 1071 3490
rect 1075 3486 1111 3490
rect 1115 3486 1295 3490
rect 1299 3486 1319 3490
rect 1323 3486 1487 3490
rect 1491 3486 1575 3490
rect 1579 3486 1815 3490
rect 1819 3486 1935 3490
rect 1939 3486 1947 3490
rect 91 3485 1947 3486
rect 1953 3487 1954 3491
rect 1953 3486 3818 3487
rect 1953 3485 1975 3486
rect 1946 3482 1975 3485
rect 1979 3482 2023 3486
rect 2027 3482 2191 3486
rect 2195 3482 2279 3486
rect 2283 3482 2399 3486
rect 2403 3482 2543 3486
rect 2547 3482 2615 3486
rect 2619 3482 2783 3486
rect 2787 3482 2831 3486
rect 2835 3482 3007 3486
rect 3011 3482 3047 3486
rect 3051 3482 3223 3486
rect 3227 3482 3263 3486
rect 3267 3482 3439 3486
rect 3443 3482 3479 3486
rect 3483 3482 3655 3486
rect 3659 3482 3679 3486
rect 3683 3482 3799 3486
rect 3803 3482 3818 3486
rect 1946 3481 3818 3482
rect 3810 3393 3811 3399
rect 3817 3398 5695 3399
rect 3817 3394 3839 3398
rect 3843 3394 3887 3398
rect 3891 3394 4151 3398
rect 4155 3394 4423 3398
rect 4427 3394 4559 3398
rect 4563 3394 4671 3398
rect 4675 3394 4711 3398
rect 4715 3394 4871 3398
rect 4875 3394 4895 3398
rect 4899 3394 5031 3398
rect 5035 3394 5111 3398
rect 5115 3394 5199 3398
rect 5203 3394 5327 3398
rect 5331 3394 5375 3398
rect 5379 3394 5543 3398
rect 5547 3394 5663 3398
rect 5667 3394 5695 3398
rect 3817 3393 5695 3394
rect 5701 3393 5702 3399
rect 96 3357 97 3363
rect 103 3362 1959 3363
rect 103 3358 111 3362
rect 115 3358 275 3362
rect 279 3358 419 3362
rect 423 3358 467 3362
rect 471 3358 571 3362
rect 575 3358 667 3362
rect 671 3358 731 3362
rect 735 3358 875 3362
rect 879 3358 907 3362
rect 911 3358 1083 3362
rect 1087 3358 1091 3362
rect 1095 3358 1267 3362
rect 1271 3358 1315 3362
rect 1319 3358 1459 3362
rect 1463 3358 1935 3362
rect 1939 3358 1959 3362
rect 103 3357 1959 3358
rect 1965 3357 1966 3363
rect 1958 3329 1959 3335
rect 1965 3334 3823 3335
rect 1965 3330 1975 3334
rect 1979 3330 1995 3334
rect 1999 3330 2163 3334
rect 2167 3330 2195 3334
rect 2199 3330 2371 3334
rect 2375 3330 2411 3334
rect 2415 3330 2587 3334
rect 2591 3330 2619 3334
rect 2623 3330 2803 3334
rect 2807 3330 2811 3334
rect 2815 3330 3003 3334
rect 3007 3330 3019 3334
rect 3023 3330 3187 3334
rect 3191 3330 3235 3334
rect 3239 3330 3371 3334
rect 3375 3330 3451 3334
rect 3455 3330 3555 3334
rect 3559 3330 3651 3334
rect 3655 3330 3799 3334
rect 3803 3330 3823 3334
rect 1965 3329 3823 3330
rect 3829 3329 3830 3335
rect 3822 3281 3823 3287
rect 3829 3286 5707 3287
rect 3829 3282 3839 3286
rect 3843 3282 3859 3286
rect 3863 3282 4099 3286
rect 4103 3282 4123 3286
rect 4127 3282 4347 3286
rect 4351 3282 4395 3286
rect 4399 3282 4579 3286
rect 4583 3282 4643 3286
rect 4647 3282 4787 3286
rect 4791 3282 4867 3286
rect 4871 3282 4987 3286
rect 4991 3282 5083 3286
rect 5087 3282 5171 3286
rect 5175 3282 5299 3286
rect 5303 3282 5355 3286
rect 5359 3282 5515 3286
rect 5519 3282 5663 3286
rect 5667 3282 5707 3286
rect 3829 3281 5707 3282
rect 5713 3281 5714 3287
rect 84 3245 85 3251
rect 91 3250 1947 3251
rect 91 3246 111 3250
rect 115 3246 495 3250
rect 499 3246 535 3250
rect 539 3246 695 3250
rect 699 3246 727 3250
rect 731 3246 903 3250
rect 907 3246 919 3250
rect 923 3246 1111 3250
rect 1115 3246 1119 3250
rect 1123 3246 1295 3250
rect 1299 3246 1343 3250
rect 1347 3246 1471 3250
rect 1475 3246 1655 3250
rect 1659 3246 1815 3250
rect 1819 3246 1935 3250
rect 1939 3246 1947 3250
rect 91 3245 1947 3246
rect 1953 3245 1954 3251
rect 1946 3217 1947 3223
rect 1953 3222 3811 3223
rect 1953 3218 1975 3222
rect 1979 3218 2023 3222
rect 2027 3218 2223 3222
rect 2227 3218 2439 3222
rect 2443 3218 2463 3222
rect 2467 3218 2647 3222
rect 2651 3218 2663 3222
rect 2667 3218 2839 3222
rect 2843 3218 2863 3222
rect 2867 3218 3031 3222
rect 3035 3218 3055 3222
rect 3059 3218 3215 3222
rect 3219 3218 3239 3222
rect 3243 3218 3399 3222
rect 3403 3218 3431 3222
rect 3435 3218 3583 3222
rect 3587 3218 3623 3222
rect 3627 3218 3799 3222
rect 3803 3218 3811 3222
rect 1953 3217 3811 3218
rect 3817 3217 3818 3223
rect 3810 3153 3811 3159
rect 3817 3158 5695 3159
rect 3817 3154 3839 3158
rect 3843 3154 3887 3158
rect 3891 3154 3903 3158
rect 3907 3154 4127 3158
rect 4131 3154 4135 3158
rect 4139 3154 4359 3158
rect 4363 3154 4375 3158
rect 4379 3154 4583 3158
rect 4587 3154 4607 3158
rect 4611 3154 4807 3158
rect 4811 3154 4815 3158
rect 4819 3154 5015 3158
rect 5019 3154 5031 3158
rect 5035 3154 5199 3158
rect 5203 3154 5383 3158
rect 5387 3154 5543 3158
rect 5547 3154 5663 3158
rect 5667 3154 5695 3158
rect 3817 3153 5695 3154
rect 5701 3153 5702 3159
rect 96 3125 97 3131
rect 103 3130 1959 3131
rect 103 3126 111 3130
rect 115 3126 427 3130
rect 431 3126 507 3130
rect 511 3126 563 3130
rect 567 3126 699 3130
rect 703 3126 835 3130
rect 839 3126 891 3130
rect 895 3126 971 3130
rect 975 3126 1083 3130
rect 1087 3126 1107 3130
rect 1111 3126 1243 3130
rect 1247 3126 1267 3130
rect 1271 3126 1379 3130
rect 1383 3126 1443 3130
rect 1447 3126 1515 3130
rect 1519 3126 1627 3130
rect 1631 3126 1651 3130
rect 1655 3126 1787 3130
rect 1791 3126 1935 3130
rect 1939 3126 1959 3130
rect 103 3125 1959 3126
rect 1965 3125 1966 3131
rect 1958 3093 1959 3099
rect 1965 3098 3823 3099
rect 1965 3094 1975 3098
rect 1979 3094 2331 3098
rect 2335 3094 2435 3098
rect 2439 3094 2555 3098
rect 2559 3094 2635 3098
rect 2639 3094 2779 3098
rect 2783 3094 2835 3098
rect 2839 3094 3003 3098
rect 3007 3094 3027 3098
rect 3031 3094 3211 3098
rect 3215 3094 3235 3098
rect 3239 3094 3403 3098
rect 3407 3094 3467 3098
rect 3471 3094 3595 3098
rect 3599 3094 3799 3098
rect 3803 3094 3823 3098
rect 1965 3093 3823 3094
rect 3829 3093 3830 3099
rect 3822 3041 3823 3047
rect 3829 3046 5707 3047
rect 3829 3042 3839 3046
rect 3843 3042 3875 3046
rect 3879 3042 3907 3046
rect 3911 3042 4075 3046
rect 4079 3042 4107 3046
rect 4111 3042 4243 3046
rect 4247 3042 4331 3046
rect 4335 3042 4411 3046
rect 4415 3042 4555 3046
rect 4559 3042 4579 3046
rect 4583 3042 4755 3046
rect 4759 3042 4779 3046
rect 4783 3042 5003 3046
rect 5007 3042 5663 3046
rect 5667 3042 5707 3046
rect 3829 3041 5707 3042
rect 5713 3041 5714 3047
rect 84 2985 85 2991
rect 91 2990 1947 2991
rect 91 2986 111 2990
rect 115 2986 199 2990
rect 203 2986 455 2990
rect 459 2986 511 2990
rect 515 2986 591 2990
rect 595 2986 727 2990
rect 731 2986 815 2990
rect 819 2986 863 2990
rect 867 2986 999 2990
rect 1003 2986 1111 2990
rect 1115 2986 1135 2990
rect 1139 2986 1271 2990
rect 1275 2986 1407 2990
rect 1411 2986 1415 2990
rect 1419 2986 1543 2990
rect 1547 2986 1679 2990
rect 1683 2986 1719 2990
rect 1723 2986 1815 2990
rect 1819 2986 1935 2990
rect 1939 2986 1947 2990
rect 91 2985 1947 2986
rect 1953 2985 1954 2991
rect 1946 2969 1947 2975
rect 1953 2974 3811 2975
rect 1953 2970 1975 2974
rect 1979 2970 2143 2974
rect 2147 2970 2343 2974
rect 2347 2970 2359 2974
rect 2363 2970 2543 2974
rect 2547 2970 2583 2974
rect 2587 2970 2743 2974
rect 2747 2970 2807 2974
rect 2811 2970 2935 2974
rect 2939 2970 3031 2974
rect 3035 2970 3135 2974
rect 3139 2970 3263 2974
rect 3267 2970 3335 2974
rect 3339 2970 3495 2974
rect 3499 2970 3799 2974
rect 3803 2970 3811 2974
rect 1953 2969 3811 2970
rect 3817 2969 3818 2975
rect 3810 2925 3811 2931
rect 3817 2930 5695 2931
rect 3817 2926 3839 2930
rect 3843 2926 3895 2930
rect 3899 2926 3935 2930
rect 3939 2926 4031 2930
rect 4035 2926 4103 2930
rect 4107 2926 4167 2930
rect 4171 2926 4271 2930
rect 4275 2926 4303 2930
rect 4307 2926 4439 2930
rect 4443 2926 4575 2930
rect 4579 2926 4607 2930
rect 4611 2926 4783 2930
rect 4787 2926 5663 2930
rect 5667 2926 5695 2930
rect 3817 2925 5695 2926
rect 5701 2925 5702 2931
rect 96 2873 97 2879
rect 103 2878 1959 2879
rect 103 2874 111 2878
rect 115 2874 131 2878
rect 135 2874 171 2878
rect 175 2874 307 2878
rect 311 2874 483 2878
rect 487 2874 523 2878
rect 527 2874 763 2878
rect 767 2874 787 2878
rect 791 2874 1011 2878
rect 1015 2874 1083 2878
rect 1087 2874 1275 2878
rect 1279 2874 1387 2878
rect 1391 2874 1539 2878
rect 1543 2874 1691 2878
rect 1695 2874 1935 2878
rect 1939 2874 1959 2878
rect 103 2873 1959 2874
rect 1965 2873 1966 2879
rect 1958 2849 1959 2855
rect 1965 2854 3823 2855
rect 1965 2850 1975 2854
rect 1979 2850 2011 2854
rect 2015 2850 2115 2854
rect 2119 2850 2259 2854
rect 2263 2850 2315 2854
rect 2319 2850 2507 2854
rect 2511 2850 2515 2854
rect 2519 2850 2715 2854
rect 2719 2850 2755 2854
rect 2759 2850 2907 2854
rect 2911 2850 3003 2854
rect 3007 2850 3107 2854
rect 3111 2850 3307 2854
rect 3311 2850 3799 2854
rect 3803 2850 3823 2854
rect 1965 2849 3823 2850
rect 3829 2849 3830 2855
rect 3822 2805 3823 2811
rect 3829 2810 5707 2811
rect 3829 2806 3839 2810
rect 3843 2806 3859 2810
rect 3863 2806 3867 2810
rect 3871 2806 3995 2810
rect 3999 2806 4003 2810
rect 4007 2806 4131 2810
rect 4135 2806 4139 2810
rect 4143 2806 4267 2810
rect 4271 2806 4275 2810
rect 4279 2806 4403 2810
rect 4407 2806 4411 2810
rect 4415 2806 4539 2810
rect 4543 2806 4547 2810
rect 4551 2806 4675 2810
rect 4679 2806 4811 2810
rect 4815 2806 5663 2810
rect 5667 2806 5707 2810
rect 3829 2805 5707 2806
rect 5713 2805 5714 2811
rect 84 2757 85 2763
rect 91 2762 1947 2763
rect 91 2758 111 2762
rect 115 2758 159 2762
rect 163 2758 279 2762
rect 283 2758 335 2762
rect 339 2758 455 2762
rect 459 2758 551 2762
rect 555 2758 647 2762
rect 651 2758 791 2762
rect 795 2758 855 2762
rect 859 2758 1039 2762
rect 1043 2758 1079 2762
rect 1083 2758 1303 2762
rect 1307 2758 1311 2762
rect 1315 2758 1551 2762
rect 1555 2758 1567 2762
rect 1571 2758 1799 2762
rect 1803 2758 1935 2762
rect 1939 2758 1947 2762
rect 91 2757 1947 2758
rect 1953 2757 1954 2763
rect 1946 2733 1947 2739
rect 1953 2738 3811 2739
rect 1953 2734 1975 2738
rect 1979 2734 2023 2738
rect 2027 2734 2039 2738
rect 2043 2734 2247 2738
rect 2251 2734 2287 2738
rect 2291 2734 2503 2738
rect 2507 2734 2535 2738
rect 2539 2734 2759 2738
rect 2763 2734 2783 2738
rect 2787 2734 3015 2738
rect 3019 2734 3031 2738
rect 3035 2734 3799 2738
rect 3803 2734 3811 2738
rect 1953 2733 3811 2734
rect 3817 2733 3818 2739
rect 3810 2693 3811 2699
rect 3817 2698 5695 2699
rect 3817 2694 3839 2698
rect 3843 2694 3887 2698
rect 3891 2694 3959 2698
rect 3963 2694 4023 2698
rect 4027 2694 4159 2698
rect 4163 2694 4255 2698
rect 4259 2694 4295 2698
rect 4299 2694 4431 2698
rect 4435 2694 4543 2698
rect 4547 2694 4567 2698
rect 4571 2694 4703 2698
rect 4707 2694 4823 2698
rect 4827 2694 4839 2698
rect 4843 2694 5111 2698
rect 5115 2694 5399 2698
rect 5403 2694 5663 2698
rect 5667 2694 5695 2698
rect 3817 2693 5695 2694
rect 5701 2693 5702 2699
rect 96 2645 97 2651
rect 103 2650 1959 2651
rect 103 2646 111 2650
rect 115 2646 251 2650
rect 255 2646 427 2650
rect 431 2646 571 2650
rect 575 2646 619 2650
rect 623 2646 731 2650
rect 735 2646 827 2650
rect 831 2646 891 2650
rect 895 2646 1043 2650
rect 1047 2646 1051 2650
rect 1055 2646 1195 2650
rect 1199 2646 1283 2650
rect 1287 2646 1355 2650
rect 1359 2646 1515 2650
rect 1519 2646 1523 2650
rect 1527 2646 1675 2650
rect 1679 2646 1771 2650
rect 1775 2646 1935 2650
rect 1939 2646 1959 2650
rect 103 2645 1959 2646
rect 1965 2645 1966 2651
rect 1958 2609 1959 2615
rect 1965 2614 3823 2615
rect 1965 2610 1975 2614
rect 1979 2610 1995 2614
rect 1999 2610 2219 2614
rect 2223 2610 2475 2614
rect 2479 2610 2555 2614
rect 2559 2610 2691 2614
rect 2695 2610 2731 2614
rect 2735 2610 2827 2614
rect 2831 2610 2963 2614
rect 2967 2610 2987 2614
rect 2991 2610 3099 2614
rect 3103 2610 3799 2614
rect 3803 2610 3823 2614
rect 1965 2609 3823 2610
rect 3829 2609 3830 2615
rect 3822 2581 3823 2587
rect 3829 2586 5707 2587
rect 3829 2582 3839 2586
rect 3843 2582 3859 2586
rect 3863 2582 3931 2586
rect 3935 2582 4083 2586
rect 4087 2582 4227 2586
rect 4231 2582 4331 2586
rect 4335 2582 4515 2586
rect 4519 2582 4579 2586
rect 4583 2582 4795 2586
rect 4799 2582 4827 2586
rect 4831 2582 5075 2586
rect 5079 2582 5083 2586
rect 5087 2582 5323 2586
rect 5327 2582 5371 2586
rect 5375 2582 5663 2586
rect 5667 2582 5707 2586
rect 3829 2581 5707 2582
rect 5713 2581 5714 2587
rect 84 2533 85 2539
rect 91 2538 1947 2539
rect 91 2534 111 2538
rect 115 2534 383 2538
rect 387 2534 599 2538
rect 603 2534 759 2538
rect 763 2534 815 2538
rect 819 2534 919 2538
rect 923 2534 1023 2538
rect 1027 2534 1071 2538
rect 1075 2534 1223 2538
rect 1227 2534 1231 2538
rect 1235 2534 1383 2538
rect 1387 2534 1431 2538
rect 1435 2534 1543 2538
rect 1547 2534 1631 2538
rect 1635 2534 1703 2538
rect 1707 2534 1815 2538
rect 1819 2534 1935 2538
rect 1939 2534 1947 2538
rect 91 2533 1947 2534
rect 1953 2533 1954 2539
rect 1946 2473 1947 2479
rect 1953 2478 3811 2479
rect 1953 2474 1975 2478
rect 1979 2474 2023 2478
rect 2027 2474 2223 2478
rect 2227 2474 2447 2478
rect 2451 2474 2583 2478
rect 2587 2474 2679 2478
rect 2683 2474 2719 2478
rect 2723 2474 2855 2478
rect 2859 2474 2927 2478
rect 2931 2474 2991 2478
rect 2995 2474 3127 2478
rect 3131 2474 3183 2478
rect 3187 2474 3439 2478
rect 3443 2474 3679 2478
rect 3683 2474 3799 2478
rect 3803 2474 3811 2478
rect 1953 2473 3811 2474
rect 3817 2473 3818 2479
rect 3810 2471 3818 2473
rect 3810 2465 3811 2471
rect 3817 2470 5695 2471
rect 3817 2466 3839 2470
rect 3843 2466 3887 2470
rect 3891 2466 4087 2470
rect 4091 2466 4111 2470
rect 4115 2466 4327 2470
rect 4331 2466 4359 2470
rect 4363 2466 4583 2470
rect 4587 2466 4607 2470
rect 4611 2466 4847 2470
rect 4851 2466 4855 2470
rect 4859 2466 5103 2470
rect 5107 2466 5119 2470
rect 5123 2466 5351 2470
rect 5355 2466 5399 2470
rect 5403 2466 5663 2470
rect 5667 2466 5695 2470
rect 3817 2465 5695 2466
rect 5701 2465 5702 2471
rect 96 2417 97 2423
rect 103 2422 1959 2423
rect 103 2418 111 2422
rect 115 2418 227 2422
rect 231 2418 355 2422
rect 359 2418 523 2422
rect 527 2418 571 2422
rect 575 2418 787 2422
rect 791 2418 835 2422
rect 839 2418 995 2422
rect 999 2418 1155 2422
rect 1159 2418 1203 2422
rect 1207 2418 1403 2422
rect 1407 2418 1483 2422
rect 1487 2418 1603 2422
rect 1607 2418 1787 2422
rect 1791 2418 1935 2422
rect 1939 2418 1959 2422
rect 103 2417 1959 2418
rect 1965 2417 1966 2423
rect 1958 2353 1959 2359
rect 1965 2358 3823 2359
rect 1965 2354 1975 2358
rect 1979 2354 1995 2358
rect 1999 2354 2155 2358
rect 2159 2354 2195 2358
rect 2199 2354 2347 2358
rect 2351 2354 2419 2358
rect 2423 2354 2539 2358
rect 2543 2354 2651 2358
rect 2655 2354 2731 2358
rect 2735 2354 2899 2358
rect 2903 2354 2923 2358
rect 2927 2354 3115 2358
rect 3119 2354 3155 2358
rect 3159 2354 3299 2358
rect 3303 2354 3411 2358
rect 3415 2354 3483 2358
rect 3487 2354 3651 2358
rect 3655 2354 3799 2358
rect 3803 2354 3823 2358
rect 1965 2353 3823 2354
rect 3829 2353 3830 2359
rect 3822 2341 3823 2347
rect 3829 2346 5707 2347
rect 3829 2342 3839 2346
rect 3843 2342 3859 2346
rect 3863 2342 4059 2346
rect 4063 2342 4299 2346
rect 4303 2342 4443 2346
rect 4447 2342 4555 2346
rect 4559 2342 4611 2346
rect 4615 2342 4787 2346
rect 4791 2342 4819 2346
rect 4823 2342 4963 2346
rect 4967 2342 5091 2346
rect 5095 2342 5147 2346
rect 5151 2342 5339 2346
rect 5343 2342 5371 2346
rect 5375 2342 5515 2346
rect 5519 2342 5663 2346
rect 5667 2342 5707 2346
rect 3829 2341 5707 2342
rect 5713 2341 5714 2347
rect 84 2289 85 2295
rect 91 2294 1947 2295
rect 91 2290 111 2294
rect 115 2290 159 2294
rect 163 2290 255 2294
rect 259 2290 367 2294
rect 371 2290 551 2294
rect 555 2290 599 2294
rect 603 2290 831 2294
rect 835 2290 863 2294
rect 867 2290 1063 2294
rect 1067 2290 1183 2294
rect 1187 2290 1511 2294
rect 1515 2290 1815 2294
rect 1819 2290 1935 2294
rect 1939 2290 1947 2294
rect 91 2289 1947 2290
rect 1953 2289 1954 2295
rect 1946 2233 1947 2239
rect 1953 2238 3811 2239
rect 1953 2234 1975 2238
rect 1979 2234 2023 2238
rect 2027 2234 2183 2238
rect 2187 2234 2191 2238
rect 2195 2234 2359 2238
rect 2363 2234 2375 2238
rect 2379 2234 2535 2238
rect 2539 2234 2567 2238
rect 2571 2234 2711 2238
rect 2715 2234 2759 2238
rect 2763 2234 2879 2238
rect 2883 2234 2951 2238
rect 2955 2234 3047 2238
rect 3051 2234 3143 2238
rect 3147 2234 3207 2238
rect 3211 2234 3327 2238
rect 3331 2234 3367 2238
rect 3371 2234 3511 2238
rect 3515 2234 3535 2238
rect 3539 2234 3679 2238
rect 3683 2234 3799 2238
rect 3803 2234 3811 2238
rect 1953 2233 3811 2234
rect 3817 2233 3818 2239
rect 3810 2217 3811 2223
rect 3817 2222 5695 2223
rect 3817 2218 3839 2222
rect 3843 2218 4471 2222
rect 4475 2218 4543 2222
rect 4547 2218 4639 2222
rect 4643 2218 4719 2222
rect 4723 2218 4815 2222
rect 4819 2218 4911 2222
rect 4915 2218 4991 2222
rect 4995 2218 5119 2222
rect 5123 2218 5175 2222
rect 5179 2218 5335 2222
rect 5339 2218 5367 2222
rect 5371 2218 5543 2222
rect 5547 2218 5663 2222
rect 5667 2218 5695 2222
rect 3817 2217 5695 2218
rect 5701 2217 5702 2223
rect 96 2165 97 2171
rect 103 2170 1959 2171
rect 103 2166 111 2170
rect 115 2166 131 2170
rect 135 2166 339 2170
rect 343 2166 347 2170
rect 351 2166 571 2170
rect 575 2166 595 2170
rect 599 2166 803 2170
rect 807 2166 835 2170
rect 839 2166 1035 2170
rect 1039 2166 1075 2170
rect 1079 2166 1315 2170
rect 1319 2166 1563 2170
rect 1567 2166 1787 2170
rect 1791 2166 1935 2170
rect 1939 2166 1959 2170
rect 103 2165 1959 2166
rect 1965 2165 1966 2171
rect 1958 2105 1959 2111
rect 1965 2110 3823 2111
rect 1965 2106 1975 2110
rect 1979 2106 1995 2110
rect 1999 2106 2163 2110
rect 2167 2106 2331 2110
rect 2335 2106 2507 2110
rect 2511 2106 2683 2110
rect 2687 2106 2851 2110
rect 2855 2106 3019 2110
rect 3023 2106 3107 2110
rect 3111 2106 3179 2110
rect 3183 2106 3243 2110
rect 3247 2106 3339 2110
rect 3343 2106 3379 2110
rect 3383 2106 3507 2110
rect 3511 2106 3515 2110
rect 3519 2106 3651 2110
rect 3655 2106 3799 2110
rect 3803 2106 3823 2110
rect 1965 2105 3823 2106
rect 3829 2110 5714 2111
rect 3829 2106 3839 2110
rect 3843 2106 4515 2110
rect 4519 2106 4635 2110
rect 4639 2106 4691 2110
rect 4695 2106 4771 2110
rect 4775 2106 4883 2110
rect 4887 2106 4907 2110
rect 4911 2106 5043 2110
rect 5047 2106 5091 2110
rect 5095 2106 5179 2110
rect 5183 2106 5307 2110
rect 5311 2106 5515 2110
rect 5519 2106 5663 2110
rect 5667 2106 5714 2110
rect 3829 2105 5714 2106
rect 84 2049 85 2055
rect 91 2054 1947 2055
rect 91 2050 111 2054
rect 115 2050 159 2054
rect 163 2050 271 2054
rect 275 2050 375 2054
rect 379 2050 407 2054
rect 411 2050 543 2054
rect 547 2050 623 2054
rect 627 2050 687 2054
rect 691 2050 831 2054
rect 835 2050 863 2054
rect 867 2050 975 2054
rect 979 2050 1103 2054
rect 1107 2050 1119 2054
rect 1123 2050 1263 2054
rect 1267 2050 1343 2054
rect 1347 2050 1407 2054
rect 1411 2050 1543 2054
rect 1547 2050 1591 2054
rect 1595 2050 1679 2054
rect 1683 2050 1815 2054
rect 1819 2050 1935 2054
rect 1939 2050 1947 2054
rect 91 2049 1947 2050
rect 1953 2049 1954 2055
rect 1946 1993 1947 1999
rect 1953 1998 3811 1999
rect 1953 1994 1975 1998
rect 1979 1994 3127 1998
rect 3131 1994 3135 1998
rect 3139 1994 3263 1998
rect 3267 1994 3271 1998
rect 3275 1994 3399 1998
rect 3403 1994 3407 1998
rect 3411 1994 3535 1998
rect 3539 1994 3543 1998
rect 3547 1994 3671 1998
rect 3675 1994 3679 1998
rect 3683 1994 3799 1998
rect 3803 1994 3811 1998
rect 1953 1993 3811 1994
rect 3817 1998 5702 1999
rect 3817 1994 3839 1998
rect 3843 1994 4663 1998
rect 4667 1994 4799 1998
rect 4803 1994 4863 1998
rect 4867 1994 4935 1998
rect 4939 1994 4999 1998
rect 5003 1994 5071 1998
rect 5075 1994 5135 1998
rect 5139 1994 5207 1998
rect 5211 1994 5271 1998
rect 5275 1994 5407 1998
rect 5411 1994 5543 1998
rect 5547 1994 5663 1998
rect 5667 1994 5702 1998
rect 3817 1993 5702 1994
rect 96 1933 97 1939
rect 103 1938 1959 1939
rect 103 1934 111 1938
rect 115 1934 187 1938
rect 191 1934 243 1938
rect 247 1934 379 1938
rect 383 1934 515 1938
rect 519 1934 587 1938
rect 591 1934 659 1938
rect 663 1934 803 1938
rect 807 1934 811 1938
rect 815 1934 947 1938
rect 951 1934 1051 1938
rect 1055 1934 1091 1938
rect 1095 1934 1235 1938
rect 1239 1934 1299 1938
rect 1303 1934 1379 1938
rect 1383 1934 1515 1938
rect 1519 1934 1555 1938
rect 1559 1934 1651 1938
rect 1655 1934 1787 1938
rect 1791 1934 1935 1938
rect 1939 1934 1959 1938
rect 103 1933 1959 1934
rect 1965 1933 1966 1939
rect 1958 1869 1959 1875
rect 1965 1874 3823 1875
rect 1965 1870 1975 1874
rect 1979 1870 1995 1874
rect 1999 1870 2227 1874
rect 2231 1870 2467 1874
rect 2471 1870 2691 1874
rect 2695 1870 2907 1874
rect 2911 1870 3099 1874
rect 3103 1870 3107 1874
rect 3111 1870 3235 1874
rect 3239 1870 3299 1874
rect 3303 1870 3371 1874
rect 3375 1870 3483 1874
rect 3487 1870 3507 1874
rect 3511 1870 3643 1874
rect 3647 1870 3651 1874
rect 3655 1870 3799 1874
rect 3803 1870 3823 1874
rect 1965 1869 3823 1870
rect 3829 1874 5714 1875
rect 3829 1870 3839 1874
rect 3843 1870 4675 1874
rect 4679 1870 4819 1874
rect 4823 1870 4835 1874
rect 4839 1870 4963 1874
rect 4967 1870 4971 1874
rect 4975 1870 5107 1874
rect 5111 1870 5243 1874
rect 5247 1870 5379 1874
rect 5383 1870 5515 1874
rect 5519 1870 5663 1874
rect 5667 1870 5714 1874
rect 3829 1869 5714 1870
rect 84 1813 85 1819
rect 91 1818 1947 1819
rect 91 1814 111 1818
rect 115 1814 159 1818
rect 163 1814 215 1818
rect 219 1814 375 1818
rect 379 1814 407 1818
rect 411 1814 591 1818
rect 595 1814 615 1818
rect 619 1814 799 1818
rect 803 1814 839 1818
rect 843 1814 999 1818
rect 1003 1814 1079 1818
rect 1083 1814 1191 1818
rect 1195 1814 1327 1818
rect 1331 1814 1383 1818
rect 1387 1814 1575 1818
rect 1579 1814 1583 1818
rect 1587 1814 1815 1818
rect 1819 1814 1935 1818
rect 1939 1814 1947 1818
rect 91 1813 1947 1814
rect 1953 1813 1954 1819
rect 1946 1749 1947 1755
rect 1953 1754 3811 1755
rect 1953 1750 1975 1754
rect 1979 1750 2023 1754
rect 2027 1750 2159 1754
rect 2163 1750 2255 1754
rect 2259 1750 2311 1754
rect 2315 1750 2471 1754
rect 2475 1750 2495 1754
rect 2499 1750 2639 1754
rect 2643 1750 2719 1754
rect 2723 1750 2807 1754
rect 2811 1750 2935 1754
rect 2939 1750 2975 1754
rect 2979 1750 3135 1754
rect 3139 1750 3151 1754
rect 3155 1750 3327 1754
rect 3331 1750 3511 1754
rect 3515 1750 3679 1754
rect 3683 1750 3799 1754
rect 3803 1750 3811 1754
rect 1953 1749 3811 1750
rect 3817 1749 3818 1755
rect 3810 1747 3818 1749
rect 3810 1741 3811 1747
rect 3817 1746 5695 1747
rect 3817 1742 3839 1746
rect 3843 1742 3887 1746
rect 3891 1742 4079 1746
rect 4083 1742 4303 1746
rect 4307 1742 4535 1746
rect 4539 1742 4703 1746
rect 4707 1742 4775 1746
rect 4779 1742 4847 1746
rect 4851 1742 4991 1746
rect 4995 1742 5023 1746
rect 5027 1742 5135 1746
rect 5139 1742 5271 1746
rect 5275 1742 5279 1746
rect 5283 1742 5407 1746
rect 5411 1742 5535 1746
rect 5539 1742 5543 1746
rect 5547 1742 5663 1746
rect 5667 1742 5695 1746
rect 3817 1741 5695 1742
rect 5701 1741 5702 1747
rect 96 1677 97 1683
rect 103 1682 1959 1683
rect 103 1678 111 1682
rect 115 1678 131 1682
rect 135 1678 347 1682
rect 351 1678 395 1682
rect 399 1678 563 1682
rect 567 1678 683 1682
rect 687 1678 771 1682
rect 775 1678 971 1682
rect 975 1678 979 1682
rect 983 1678 1163 1682
rect 1167 1678 1275 1682
rect 1279 1678 1355 1682
rect 1359 1678 1547 1682
rect 1551 1678 1935 1682
rect 1939 1678 1959 1682
rect 103 1677 1959 1678
rect 1965 1677 1966 1683
rect 1958 1629 1959 1635
rect 1965 1634 3823 1635
rect 1965 1630 1975 1634
rect 1979 1630 1995 1634
rect 1999 1630 2091 1634
rect 2095 1630 2131 1634
rect 2135 1630 2227 1634
rect 2231 1630 2283 1634
rect 2287 1630 2363 1634
rect 2367 1630 2443 1634
rect 2447 1630 2499 1634
rect 2503 1630 2611 1634
rect 2615 1630 2635 1634
rect 2639 1630 2771 1634
rect 2775 1630 2779 1634
rect 2783 1630 2907 1634
rect 2911 1630 2947 1634
rect 2951 1630 3043 1634
rect 3047 1630 3123 1634
rect 3127 1630 3179 1634
rect 3183 1630 3799 1634
rect 3803 1630 3823 1634
rect 1965 1629 3823 1630
rect 3829 1634 5714 1635
rect 3829 1630 3839 1634
rect 3843 1630 3859 1634
rect 3863 1630 3995 1634
rect 3999 1630 4051 1634
rect 4055 1630 4155 1634
rect 4159 1630 4275 1634
rect 4279 1630 4355 1634
rect 4359 1630 4507 1634
rect 4511 1630 4587 1634
rect 4591 1630 4747 1634
rect 4751 1630 4851 1634
rect 4855 1630 4995 1634
rect 4999 1630 5131 1634
rect 5135 1630 5251 1634
rect 5255 1630 5419 1634
rect 5423 1630 5507 1634
rect 5511 1630 5663 1634
rect 5667 1630 5714 1634
rect 3829 1629 5714 1630
rect 84 1553 85 1559
rect 91 1558 1947 1559
rect 91 1554 111 1558
rect 115 1554 159 1558
rect 163 1554 375 1558
rect 379 1554 423 1558
rect 427 1554 607 1558
rect 611 1554 711 1558
rect 715 1554 839 1558
rect 843 1554 1007 1558
rect 1011 1554 1071 1558
rect 1075 1554 1303 1558
rect 1307 1554 1935 1558
rect 1939 1554 1947 1558
rect 91 1553 1947 1554
rect 1953 1553 1954 1559
rect 3810 1517 3811 1523
rect 3817 1522 5695 1523
rect 3817 1518 3839 1522
rect 3843 1518 3887 1522
rect 3891 1518 4023 1522
rect 4027 1518 4159 1522
rect 4163 1518 4183 1522
rect 4187 1518 4303 1522
rect 4307 1518 4383 1522
rect 4387 1518 4495 1522
rect 4499 1518 4615 1522
rect 4619 1518 4719 1522
rect 4723 1518 4879 1522
rect 4883 1518 4967 1522
rect 4971 1518 5159 1522
rect 5163 1518 5223 1522
rect 5227 1518 5447 1522
rect 5451 1518 5487 1522
rect 5491 1518 5663 1522
rect 5667 1518 5695 1522
rect 3817 1517 5695 1518
rect 5701 1517 5702 1523
rect 1946 1497 1947 1503
rect 1953 1502 3811 1503
rect 1953 1498 1975 1502
rect 1979 1498 2023 1502
rect 2027 1498 2119 1502
rect 2123 1498 2159 1502
rect 2163 1498 2255 1502
rect 2259 1498 2295 1502
rect 2299 1498 2391 1502
rect 2395 1498 2431 1502
rect 2435 1498 2527 1502
rect 2531 1498 2567 1502
rect 2571 1498 2663 1502
rect 2667 1498 2703 1502
rect 2707 1498 2799 1502
rect 2803 1498 2839 1502
rect 2843 1498 2935 1502
rect 2939 1498 2975 1502
rect 2979 1498 3071 1502
rect 3075 1498 3207 1502
rect 3211 1498 3799 1502
rect 3803 1498 3811 1502
rect 1953 1497 3811 1498
rect 3817 1497 3818 1503
rect 96 1429 97 1435
rect 103 1434 1959 1435
rect 103 1430 111 1434
rect 115 1430 131 1434
rect 135 1430 347 1434
rect 351 1430 411 1434
rect 415 1430 579 1434
rect 583 1430 739 1434
rect 743 1430 811 1434
rect 815 1430 1043 1434
rect 1047 1430 1091 1434
rect 1095 1430 1275 1434
rect 1279 1430 1451 1434
rect 1455 1430 1787 1434
rect 1791 1430 1935 1434
rect 1939 1430 1959 1434
rect 103 1429 1959 1430
rect 1965 1429 1966 1435
rect 3822 1401 3823 1407
rect 3829 1406 5707 1407
rect 3829 1402 3839 1406
rect 3843 1402 3859 1406
rect 3863 1402 3995 1406
rect 3999 1402 4059 1406
rect 4063 1402 4131 1406
rect 4135 1402 4275 1406
rect 4279 1402 4307 1406
rect 4311 1402 4467 1406
rect 4471 1402 4579 1406
rect 4583 1402 4691 1406
rect 4695 1402 4875 1406
rect 4879 1402 4939 1406
rect 4943 1402 5187 1406
rect 5191 1402 5195 1406
rect 5199 1402 5459 1406
rect 5463 1402 5499 1406
rect 5503 1402 5663 1406
rect 5667 1402 5707 1406
rect 3829 1401 5707 1402
rect 5713 1401 5714 1407
rect 1958 1377 1959 1383
rect 1965 1382 3823 1383
rect 1965 1378 1975 1382
rect 1979 1378 1995 1382
rect 1999 1378 2131 1382
rect 2135 1378 2267 1382
rect 2271 1378 2275 1382
rect 2279 1378 2403 1382
rect 2407 1378 2539 1382
rect 2543 1378 2563 1382
rect 2567 1378 2675 1382
rect 2679 1378 2811 1382
rect 2815 1378 2843 1382
rect 2847 1378 2947 1382
rect 2951 1378 3123 1382
rect 3127 1378 3395 1382
rect 3399 1378 3651 1382
rect 3655 1378 3799 1382
rect 3803 1378 3823 1382
rect 1965 1377 3823 1378
rect 3829 1377 3830 1383
rect 84 1317 85 1323
rect 91 1322 1947 1323
rect 91 1318 111 1322
rect 115 1318 159 1322
rect 163 1318 359 1322
rect 363 1318 439 1322
rect 443 1318 575 1322
rect 579 1318 767 1322
rect 771 1318 775 1322
rect 779 1318 967 1322
rect 971 1318 1119 1322
rect 1123 1318 1151 1322
rect 1155 1318 1327 1322
rect 1331 1318 1479 1322
rect 1483 1318 1495 1322
rect 1499 1318 1663 1322
rect 1667 1318 1815 1322
rect 1819 1318 1935 1322
rect 1939 1318 1947 1322
rect 91 1317 1947 1318
rect 1953 1317 1954 1323
rect 3810 1281 3811 1287
rect 3817 1286 5695 1287
rect 3817 1282 3839 1286
rect 3843 1282 3887 1286
rect 3891 1282 4087 1286
rect 4091 1282 4335 1286
rect 4339 1282 4607 1286
rect 4611 1282 4615 1286
rect 4619 1282 4791 1286
rect 4795 1282 4903 1286
rect 4907 1282 4975 1286
rect 4979 1282 5167 1286
rect 5171 1282 5215 1286
rect 5219 1282 5367 1286
rect 5371 1282 5527 1286
rect 5531 1282 5543 1286
rect 5547 1282 5663 1286
rect 5667 1282 5695 1286
rect 3817 1281 5695 1282
rect 5701 1281 5702 1287
rect 1946 1241 1947 1247
rect 1953 1246 3811 1247
rect 1953 1242 1975 1246
rect 1979 1242 2023 1246
rect 2027 1242 2303 1246
rect 2307 1242 2591 1246
rect 2595 1242 2655 1246
rect 2659 1242 2831 1246
rect 2835 1242 2871 1246
rect 2875 1242 3007 1246
rect 3011 1242 3151 1246
rect 3155 1242 3183 1246
rect 3187 1242 3359 1246
rect 3363 1242 3423 1246
rect 3427 1242 3543 1246
rect 3547 1242 3679 1246
rect 3683 1242 3799 1246
rect 3803 1242 3811 1246
rect 1953 1241 3811 1242
rect 3817 1241 3818 1247
rect 96 1193 97 1199
rect 103 1198 1959 1199
rect 103 1194 111 1198
rect 115 1194 131 1198
rect 135 1194 291 1198
rect 295 1194 331 1198
rect 335 1194 475 1198
rect 479 1194 547 1198
rect 551 1194 659 1198
rect 663 1194 747 1198
rect 751 1194 835 1198
rect 839 1194 939 1198
rect 943 1194 1003 1198
rect 1007 1194 1123 1198
rect 1127 1194 1171 1198
rect 1175 1194 1299 1198
rect 1303 1194 1331 1198
rect 1335 1194 1467 1198
rect 1471 1194 1491 1198
rect 1495 1194 1635 1198
rect 1639 1194 1651 1198
rect 1655 1194 1787 1198
rect 1791 1194 1935 1198
rect 1939 1194 1959 1198
rect 103 1193 1959 1194
rect 1965 1193 1966 1199
rect 3822 1165 3823 1171
rect 3829 1170 5707 1171
rect 3829 1166 3839 1170
rect 3843 1166 4587 1170
rect 4591 1166 4763 1170
rect 4767 1166 4835 1170
rect 4839 1166 4947 1170
rect 4951 1166 4971 1170
rect 4975 1166 5107 1170
rect 5111 1166 5139 1170
rect 5143 1166 5243 1170
rect 5247 1166 5339 1170
rect 5343 1166 5379 1170
rect 5383 1166 5515 1170
rect 5519 1166 5663 1170
rect 5667 1166 5707 1170
rect 3829 1165 5707 1166
rect 5713 1165 5714 1171
rect 1958 1113 1959 1119
rect 1965 1118 3823 1119
rect 1965 1114 1975 1118
rect 1979 1114 1995 1118
rect 1999 1114 2171 1118
rect 2175 1114 2363 1118
rect 2367 1114 2547 1118
rect 2551 1114 2627 1118
rect 2631 1114 2723 1118
rect 2727 1114 2803 1118
rect 2807 1114 2891 1118
rect 2895 1114 2979 1118
rect 2983 1114 3059 1118
rect 3063 1114 3155 1118
rect 3159 1114 3219 1118
rect 3223 1114 3331 1118
rect 3335 1114 3387 1118
rect 3391 1114 3515 1118
rect 3519 1114 3799 1118
rect 3803 1114 3823 1118
rect 1965 1113 3823 1114
rect 3829 1113 3830 1119
rect 84 1069 85 1075
rect 91 1074 1947 1075
rect 91 1070 111 1074
rect 115 1070 159 1074
rect 163 1070 175 1074
rect 179 1070 319 1074
rect 323 1070 431 1074
rect 435 1070 503 1074
rect 507 1070 687 1074
rect 691 1070 863 1074
rect 867 1070 951 1074
rect 955 1070 1031 1074
rect 1035 1070 1199 1074
rect 1203 1070 1215 1074
rect 1219 1070 1359 1074
rect 1363 1070 1519 1074
rect 1523 1070 1679 1074
rect 1683 1070 1815 1074
rect 1819 1070 1935 1074
rect 1939 1070 1947 1074
rect 91 1069 1947 1070
rect 1953 1069 1954 1075
rect 3810 1049 3811 1055
rect 3817 1054 5695 1055
rect 3817 1050 3839 1054
rect 3843 1050 4807 1054
rect 4811 1050 4863 1054
rect 4867 1050 4943 1054
rect 4947 1050 4999 1054
rect 5003 1050 5079 1054
rect 5083 1050 5135 1054
rect 5139 1050 5215 1054
rect 5219 1050 5271 1054
rect 5275 1050 5351 1054
rect 5355 1050 5407 1054
rect 5411 1050 5487 1054
rect 5491 1050 5543 1054
rect 5547 1050 5663 1054
rect 5667 1050 5695 1054
rect 3817 1049 5695 1050
rect 5701 1049 5702 1055
rect 1946 1001 1947 1007
rect 1953 1006 3811 1007
rect 1953 1002 1975 1006
rect 1979 1002 2023 1006
rect 2027 1002 2191 1006
rect 2195 1002 2199 1006
rect 2203 1002 2375 1006
rect 2379 1002 2391 1006
rect 2395 1002 2567 1006
rect 2571 1002 2575 1006
rect 2579 1002 2751 1006
rect 2755 1002 2759 1006
rect 2763 1002 2919 1006
rect 2923 1002 2943 1006
rect 2947 1002 3087 1006
rect 3091 1002 3127 1006
rect 3131 1002 3247 1006
rect 3251 1002 3311 1006
rect 3315 1002 3415 1006
rect 3419 1002 3495 1006
rect 3499 1002 3679 1006
rect 3683 1002 3799 1006
rect 3803 1002 3811 1006
rect 1953 1001 3811 1002
rect 3817 1001 3818 1007
rect 96 945 97 951
rect 103 950 1959 951
rect 103 946 111 950
rect 115 946 147 950
rect 151 946 235 950
rect 239 946 403 950
rect 407 946 459 950
rect 463 946 659 950
rect 663 946 683 950
rect 687 946 907 950
rect 911 946 923 950
rect 927 946 1131 950
rect 1135 946 1187 950
rect 1191 946 1363 950
rect 1367 946 1935 950
rect 1939 946 1959 950
rect 103 945 1959 946
rect 1965 945 1966 951
rect 3822 933 3823 939
rect 3829 938 5707 939
rect 3829 934 3839 938
rect 3843 934 3859 938
rect 3863 934 3995 938
rect 3999 934 4171 938
rect 4175 934 4387 938
rect 4391 934 4643 938
rect 4647 934 4779 938
rect 4783 934 4915 938
rect 4919 934 4931 938
rect 4935 934 5051 938
rect 5055 934 5187 938
rect 5191 934 5235 938
rect 5239 934 5323 938
rect 5327 934 5459 938
rect 5463 934 5515 938
rect 5519 934 5663 938
rect 5667 934 5707 938
rect 3829 933 5707 934
rect 5713 933 5714 939
rect 1958 885 1959 891
rect 1965 890 3823 891
rect 1965 886 1975 890
rect 1979 886 1995 890
rect 1999 886 2163 890
rect 2167 886 2179 890
rect 2183 886 2347 890
rect 2351 886 2403 890
rect 2407 886 2539 890
rect 2543 886 2675 890
rect 2679 886 2731 890
rect 2735 886 2915 890
rect 2919 886 2987 890
rect 2991 886 3099 890
rect 3103 886 3283 890
rect 3287 886 3323 890
rect 3327 886 3467 890
rect 3471 886 3651 890
rect 3655 886 3799 890
rect 3803 886 3823 890
rect 1965 885 3823 886
rect 3829 885 3830 891
rect 84 817 85 823
rect 91 822 1947 823
rect 91 818 111 822
rect 115 818 175 822
rect 179 818 263 822
rect 267 818 431 822
rect 435 818 487 822
rect 491 818 671 822
rect 675 818 711 822
rect 715 818 903 822
rect 907 818 935 822
rect 939 818 1127 822
rect 1131 818 1159 822
rect 1163 818 1351 822
rect 1355 818 1391 822
rect 1395 818 1575 822
rect 1579 818 1935 822
rect 1939 818 1947 822
rect 91 817 1947 818
rect 1953 817 1954 823
rect 3810 821 3811 827
rect 3817 826 5695 827
rect 3817 822 3839 826
rect 3843 822 3887 826
rect 3891 822 4023 826
rect 4027 822 4159 826
rect 4163 822 4199 826
rect 4203 822 4295 826
rect 4299 822 4415 826
rect 4419 822 4431 826
rect 4435 822 4567 826
rect 4571 822 4671 826
rect 4675 822 4719 826
rect 4723 822 4895 826
rect 4899 822 4959 826
rect 4963 822 5087 826
rect 5091 822 5263 826
rect 5267 822 5287 826
rect 5291 822 5487 826
rect 5491 822 5543 826
rect 5547 822 5663 826
rect 5667 822 5695 826
rect 3817 821 5695 822
rect 5701 821 5702 827
rect 96 705 97 711
rect 103 710 1959 711
rect 103 706 111 710
rect 115 706 131 710
rect 135 706 147 710
rect 151 706 315 710
rect 319 706 403 710
rect 407 706 523 710
rect 527 706 643 710
rect 647 706 723 710
rect 727 706 875 710
rect 879 706 907 710
rect 911 706 1083 710
rect 1087 706 1099 710
rect 1103 706 1259 710
rect 1263 706 1323 710
rect 1327 706 1427 710
rect 1431 706 1547 710
rect 1551 706 1595 710
rect 1599 706 1771 710
rect 1775 706 1935 710
rect 1939 706 1959 710
rect 103 705 1959 706
rect 1965 705 1966 711
rect 3822 705 3823 711
rect 3829 710 5707 711
rect 3829 706 3839 710
rect 3843 706 3859 710
rect 3863 706 3995 710
rect 3999 706 4131 710
rect 4135 706 4267 710
rect 4271 706 4403 710
rect 4407 706 4539 710
rect 4543 706 4691 710
rect 4695 706 4699 710
rect 4703 706 4867 710
rect 4871 706 4891 710
rect 4895 706 5059 710
rect 5063 706 5099 710
rect 5103 706 5259 710
rect 5263 706 5315 710
rect 5319 706 5459 710
rect 5463 706 5515 710
rect 5519 706 5663 710
rect 5667 706 5707 710
rect 3829 705 5707 706
rect 5713 705 5714 711
rect 84 593 85 599
rect 91 598 1947 599
rect 91 594 111 598
rect 115 594 159 598
rect 163 594 343 598
rect 347 594 375 598
rect 379 594 551 598
rect 555 594 599 598
rect 603 594 751 598
rect 755 594 807 598
rect 811 594 935 598
rect 939 594 999 598
rect 1003 594 1111 598
rect 1115 594 1175 598
rect 1179 594 1287 598
rect 1291 594 1343 598
rect 1347 594 1455 598
rect 1459 594 1511 598
rect 1515 594 1623 598
rect 1627 594 1671 598
rect 1675 594 1799 598
rect 1803 594 1815 598
rect 1819 594 1935 598
rect 1939 594 1947 598
rect 91 593 1947 594
rect 1953 593 1954 599
rect 3810 593 3811 599
rect 3817 598 5695 599
rect 3817 594 3839 598
rect 3843 594 3887 598
rect 3891 594 4023 598
rect 4027 594 4071 598
rect 4075 594 4159 598
rect 4163 594 4295 598
rect 4299 594 4311 598
rect 4315 594 4431 598
rect 4435 594 4567 598
rect 4571 594 4575 598
rect 4579 594 4727 598
rect 4731 594 4855 598
rect 4859 594 4919 598
rect 4923 594 5127 598
rect 5131 594 5151 598
rect 5155 594 5343 598
rect 5347 594 5447 598
rect 5451 594 5543 598
rect 5547 594 5663 598
rect 5667 594 5695 598
rect 3817 593 5695 594
rect 5701 593 5702 599
rect 1946 573 1947 579
rect 1953 578 3811 579
rect 1953 574 1975 578
rect 1979 574 2023 578
rect 2027 574 2207 578
rect 2211 574 2431 578
rect 2435 574 2703 578
rect 2707 574 3015 578
rect 3019 574 3135 578
rect 3139 574 3271 578
rect 3275 574 3351 578
rect 3355 574 3407 578
rect 3411 574 3543 578
rect 3547 574 3679 578
rect 3683 574 3799 578
rect 3803 574 3811 578
rect 1953 573 3811 574
rect 3817 573 3818 579
rect 96 481 97 487
rect 103 486 1959 487
rect 103 482 111 486
rect 115 482 131 486
rect 135 482 155 486
rect 159 482 347 486
rect 351 482 483 486
rect 487 482 571 486
rect 575 482 779 486
rect 783 482 811 486
rect 815 482 971 486
rect 975 482 1139 486
rect 1143 482 1147 486
rect 1151 482 1315 486
rect 1319 482 1475 486
rect 1479 482 1483 486
rect 1487 482 1643 486
rect 1647 482 1787 486
rect 1791 482 1935 486
rect 1939 482 1959 486
rect 103 481 1959 482
rect 1965 481 1966 487
rect 3822 469 3823 475
rect 3829 474 5707 475
rect 3829 470 3839 474
rect 3843 470 3859 474
rect 3863 470 4043 474
rect 4047 470 4283 474
rect 4287 470 4451 474
rect 4455 470 4547 474
rect 4551 470 4643 474
rect 4647 470 4827 474
rect 4831 470 4843 474
rect 4847 470 5051 474
rect 5055 470 5123 474
rect 5127 470 5267 474
rect 5271 470 5419 474
rect 5423 470 5483 474
rect 5487 470 5663 474
rect 5667 470 5707 474
rect 3829 469 5707 470
rect 5713 469 5714 475
rect 3822 467 3830 469
rect 1958 461 1959 467
rect 1965 466 3823 467
rect 1965 462 1975 466
rect 1979 462 1995 466
rect 1999 462 2203 466
rect 2207 462 2427 466
rect 2431 462 2651 466
rect 2655 462 2859 466
rect 2863 462 3067 466
rect 3071 462 3107 466
rect 3111 462 3243 466
rect 3247 462 3267 466
rect 3271 462 3379 466
rect 3383 462 3467 466
rect 3471 462 3515 466
rect 3519 462 3651 466
rect 3655 462 3799 466
rect 3803 462 3823 466
rect 1965 461 3823 462
rect 3829 461 3830 467
rect 84 357 85 363
rect 91 362 1947 363
rect 91 358 111 362
rect 115 358 183 362
rect 187 358 279 362
rect 283 358 487 362
rect 491 358 511 362
rect 515 358 703 362
rect 707 358 839 362
rect 843 358 919 362
rect 923 358 1135 362
rect 1139 358 1167 362
rect 1171 358 1503 362
rect 1507 358 1815 362
rect 1819 358 1935 362
rect 1939 358 1947 362
rect 91 357 1947 358
rect 1953 357 1954 363
rect 3810 353 3811 359
rect 3817 358 5695 359
rect 3817 354 3839 358
rect 3843 354 4479 358
rect 4483 354 4615 358
rect 4619 354 4671 358
rect 4675 354 4775 358
rect 4779 354 4871 358
rect 4875 354 4951 358
rect 4955 354 5079 358
rect 5083 354 5135 358
rect 5139 354 5295 358
rect 5299 354 5327 358
rect 5331 354 5511 358
rect 5515 354 5527 358
rect 5531 354 5663 358
rect 5667 354 5695 358
rect 3817 353 5695 354
rect 5701 353 5702 359
rect 1946 333 1947 339
rect 1953 338 3811 339
rect 1953 334 1975 338
rect 1979 334 2023 338
rect 2027 334 2159 338
rect 2163 334 2231 338
rect 2235 334 2295 338
rect 2299 334 2431 338
rect 2435 334 2455 338
rect 2459 334 2567 338
rect 2571 334 2679 338
rect 2683 334 2703 338
rect 2707 334 2839 338
rect 2843 334 2887 338
rect 2891 334 2975 338
rect 2979 334 3095 338
rect 3099 334 3111 338
rect 3115 334 3247 338
rect 3251 334 3295 338
rect 3299 334 3383 338
rect 3387 334 3495 338
rect 3499 334 3519 338
rect 3523 334 3655 338
rect 3659 334 3679 338
rect 3683 334 3799 338
rect 3803 334 3811 338
rect 1953 333 3811 334
rect 3817 333 3818 339
rect 96 205 97 211
rect 103 210 1959 211
rect 103 206 111 210
rect 115 206 131 210
rect 135 206 251 210
rect 255 206 267 210
rect 271 206 403 210
rect 407 206 459 210
rect 463 206 539 210
rect 543 206 675 210
rect 679 206 811 210
rect 815 206 891 210
rect 895 206 947 210
rect 951 206 1083 210
rect 1087 206 1107 210
rect 1111 206 1935 210
rect 1939 206 1959 210
rect 103 205 1959 206
rect 1965 205 1966 211
rect 3822 201 3823 207
rect 3829 206 5707 207
rect 3829 202 3839 206
rect 3843 202 4291 206
rect 4295 202 4427 206
rect 4431 202 4563 206
rect 4567 202 4587 206
rect 4591 202 4699 206
rect 4703 202 4747 206
rect 4751 202 4835 206
rect 4839 202 4923 206
rect 4927 202 4971 206
rect 4975 202 5107 206
rect 5111 202 5243 206
rect 5247 202 5299 206
rect 5303 202 5379 206
rect 5383 202 5499 206
rect 5503 202 5515 206
rect 5519 202 5663 206
rect 5667 202 5707 206
rect 3829 201 5707 202
rect 5713 201 5714 207
rect 1958 185 1959 191
rect 1965 190 3823 191
rect 1965 186 1975 190
rect 1979 186 1995 190
rect 1999 186 2131 190
rect 2135 186 2267 190
rect 2271 186 2403 190
rect 2407 186 2539 190
rect 2543 186 2675 190
rect 2679 186 2811 190
rect 2815 186 2947 190
rect 2951 186 3083 190
rect 3087 186 3219 190
rect 3223 186 3355 190
rect 3359 186 3491 190
rect 3495 186 3627 190
rect 3631 186 3799 190
rect 3803 186 3823 190
rect 1965 185 3823 186
rect 3829 185 3830 191
rect 84 93 85 99
rect 91 98 1947 99
rect 91 94 111 98
rect 115 94 159 98
rect 163 94 295 98
rect 299 94 431 98
rect 435 94 567 98
rect 571 94 703 98
rect 707 94 839 98
rect 843 94 975 98
rect 979 94 1111 98
rect 1115 94 1935 98
rect 1939 94 1947 98
rect 91 93 1947 94
rect 1953 93 1954 99
rect 3810 89 3811 95
rect 3817 94 5695 95
rect 3817 90 3839 94
rect 3843 90 4319 94
rect 4323 90 4455 94
rect 4459 90 4591 94
rect 4595 90 4727 94
rect 4731 90 4863 94
rect 4867 90 4999 94
rect 5003 90 5135 94
rect 5139 90 5271 94
rect 5275 90 5407 94
rect 5411 90 5543 94
rect 5547 90 5663 94
rect 5667 90 5695 94
rect 3817 89 5695 90
rect 5701 89 5702 95
rect 1946 73 1947 79
rect 1953 78 3811 79
rect 1953 74 1975 78
rect 1979 74 2023 78
rect 2027 74 2159 78
rect 2163 74 2295 78
rect 2299 74 2431 78
rect 2435 74 2567 78
rect 2571 74 2703 78
rect 2707 74 2839 78
rect 2843 74 2975 78
rect 2979 74 3111 78
rect 3115 74 3247 78
rect 3251 74 3383 78
rect 3387 74 3519 78
rect 3523 74 3655 78
rect 3659 74 3799 78
rect 3803 74 3811 78
rect 1953 73 3811 74
rect 3817 73 3818 79
<< m5c >>
rect 85 5753 91 5759
rect 1947 5753 1953 5759
rect 1947 5653 1953 5659
rect 3811 5653 3817 5659
rect 97 5641 103 5647
rect 1959 5641 1965 5647
rect 1959 5541 1965 5547
rect 3823 5541 3829 5547
rect 85 5529 91 5535
rect 1947 5529 1953 5535
rect 1947 5427 1953 5433
rect 97 5417 103 5423
rect 1959 5417 1965 5423
rect 3811 5421 3817 5427
rect 3811 5405 3817 5411
rect 5695 5405 5701 5411
rect 85 5305 91 5311
rect 1947 5305 1953 5311
rect 1959 5309 1965 5315
rect 3823 5309 3829 5315
rect 3823 5277 3829 5283
rect 5707 5277 5713 5283
rect 1947 5197 1953 5203
rect 3811 5197 3817 5203
rect 3811 5137 3817 5143
rect 5695 5137 5701 5143
rect 97 5089 103 5095
rect 1959 5089 1965 5095
rect 3823 5013 3829 5019
rect 5707 5013 5713 5019
rect 85 4977 91 4983
rect 1947 4977 1953 4983
rect 1947 4941 1953 4947
rect 3811 4941 3817 4947
rect 3811 4881 3817 4887
rect 5695 4881 5701 4887
rect 97 4857 103 4863
rect 1959 4857 1965 4863
rect 1959 4805 1965 4811
rect 3823 4805 3829 4811
rect 3823 4765 3829 4771
rect 5707 4765 5713 4771
rect 85 4737 91 4743
rect 1947 4737 1953 4743
rect 1947 4689 1953 4695
rect 3811 4689 3817 4695
rect 3811 4653 3817 4659
rect 5695 4653 5701 4659
rect 97 4609 103 4615
rect 1959 4609 1965 4615
rect 1959 4573 1965 4579
rect 3823 4573 3829 4579
rect 3823 4541 3829 4547
rect 5707 4541 5713 4547
rect 85 4493 91 4499
rect 1947 4493 1953 4499
rect 1947 4453 1953 4459
rect 3811 4453 3817 4459
rect 3811 4421 3817 4427
rect 5695 4421 5701 4427
rect 97 4377 103 4383
rect 1959 4377 1965 4383
rect 1959 4333 1965 4339
rect 3823 4333 3829 4339
rect 3823 4309 3829 4315
rect 5707 4309 5713 4315
rect 85 4249 91 4255
rect 1947 4249 1953 4255
rect 1947 4213 1953 4219
rect 3811 4213 3817 4219
rect 3811 4161 3817 4167
rect 5695 4161 5701 4167
rect 97 4133 103 4139
rect 1959 4133 1965 4139
rect 1959 4081 1965 4087
rect 3823 4081 3829 4087
rect 3823 4049 3829 4055
rect 5707 4049 5713 4055
rect 85 3997 91 4003
rect 1947 3997 1953 4003
rect 1947 3965 1953 3971
rect 3811 3965 3817 3971
rect 3811 3913 3817 3919
rect 5695 3913 5701 3919
rect 97 3857 103 3863
rect 1959 3857 1965 3863
rect 1959 3841 1965 3847
rect 3823 3841 3829 3847
rect 3823 3785 3829 3791
rect 5707 3785 5713 3791
rect 85 3745 91 3751
rect 1947 3745 1953 3751
rect 1947 3725 1953 3731
rect 3811 3725 3817 3731
rect 3811 3645 3817 3651
rect 5695 3645 5701 3651
rect 97 3621 103 3627
rect 1959 3621 1965 3627
rect 1959 3601 1965 3607
rect 3823 3601 3829 3607
rect 3823 3509 3829 3515
rect 5707 3509 5713 3515
rect 85 3485 91 3491
rect 1947 3485 1953 3491
rect 3811 3393 3817 3399
rect 5695 3393 5701 3399
rect 97 3357 103 3363
rect 1959 3357 1965 3363
rect 1959 3329 1965 3335
rect 3823 3329 3829 3335
rect 3823 3281 3829 3287
rect 5707 3281 5713 3287
rect 85 3245 91 3251
rect 1947 3245 1953 3251
rect 1947 3217 1953 3223
rect 3811 3217 3817 3223
rect 3811 3153 3817 3159
rect 5695 3153 5701 3159
rect 97 3125 103 3131
rect 1959 3125 1965 3131
rect 1959 3093 1965 3099
rect 3823 3093 3829 3099
rect 3823 3041 3829 3047
rect 5707 3041 5713 3047
rect 85 2985 91 2991
rect 1947 2985 1953 2991
rect 1947 2969 1953 2975
rect 3811 2969 3817 2975
rect 3811 2925 3817 2931
rect 5695 2925 5701 2931
rect 97 2873 103 2879
rect 1959 2873 1965 2879
rect 1959 2849 1965 2855
rect 3823 2849 3829 2855
rect 3823 2805 3829 2811
rect 5707 2805 5713 2811
rect 85 2757 91 2763
rect 1947 2757 1953 2763
rect 1947 2733 1953 2739
rect 3811 2733 3817 2739
rect 3811 2693 3817 2699
rect 5695 2693 5701 2699
rect 97 2645 103 2651
rect 1959 2645 1965 2651
rect 1959 2609 1965 2615
rect 3823 2609 3829 2615
rect 3823 2581 3829 2587
rect 5707 2581 5713 2587
rect 85 2533 91 2539
rect 1947 2533 1953 2539
rect 1947 2473 1953 2479
rect 3811 2473 3817 2479
rect 3811 2465 3817 2471
rect 5695 2465 5701 2471
rect 97 2417 103 2423
rect 1959 2417 1965 2423
rect 1959 2353 1965 2359
rect 3823 2353 3829 2359
rect 3823 2341 3829 2347
rect 5707 2341 5713 2347
rect 85 2289 91 2295
rect 1947 2289 1953 2295
rect 1947 2233 1953 2239
rect 3811 2233 3817 2239
rect 3811 2217 3817 2223
rect 5695 2217 5701 2223
rect 97 2165 103 2171
rect 1959 2165 1965 2171
rect 1959 2105 1965 2111
rect 3823 2105 3829 2111
rect 85 2049 91 2055
rect 1947 2049 1953 2055
rect 1947 1993 1953 1999
rect 3811 1993 3817 1999
rect 97 1933 103 1939
rect 1959 1933 1965 1939
rect 1959 1869 1965 1875
rect 3823 1869 3829 1875
rect 85 1813 91 1819
rect 1947 1813 1953 1819
rect 1947 1749 1953 1755
rect 3811 1749 3817 1755
rect 3811 1741 3817 1747
rect 5695 1741 5701 1747
rect 97 1677 103 1683
rect 1959 1677 1965 1683
rect 1959 1629 1965 1635
rect 3823 1629 3829 1635
rect 85 1553 91 1559
rect 1947 1553 1953 1559
rect 3811 1517 3817 1523
rect 5695 1517 5701 1523
rect 1947 1497 1953 1503
rect 3811 1497 3817 1503
rect 97 1429 103 1435
rect 1959 1429 1965 1435
rect 3823 1401 3829 1407
rect 5707 1401 5713 1407
rect 1959 1377 1965 1383
rect 3823 1377 3829 1383
rect 85 1317 91 1323
rect 1947 1317 1953 1323
rect 3811 1281 3817 1287
rect 5695 1281 5701 1287
rect 1947 1241 1953 1247
rect 3811 1241 3817 1247
rect 97 1193 103 1199
rect 1959 1193 1965 1199
rect 3823 1165 3829 1171
rect 5707 1165 5713 1171
rect 1959 1113 1965 1119
rect 3823 1113 3829 1119
rect 85 1069 91 1075
rect 1947 1069 1953 1075
rect 3811 1049 3817 1055
rect 5695 1049 5701 1055
rect 1947 1001 1953 1007
rect 3811 1001 3817 1007
rect 97 945 103 951
rect 1959 945 1965 951
rect 3823 933 3829 939
rect 5707 933 5713 939
rect 1959 885 1965 891
rect 3823 885 3829 891
rect 85 817 91 823
rect 1947 817 1953 823
rect 3811 821 3817 827
rect 5695 821 5701 827
rect 97 705 103 711
rect 1959 705 1965 711
rect 3823 705 3829 711
rect 5707 705 5713 711
rect 85 593 91 599
rect 1947 593 1953 599
rect 3811 593 3817 599
rect 5695 593 5701 599
rect 1947 573 1953 579
rect 3811 573 3817 579
rect 97 481 103 487
rect 1959 481 1965 487
rect 3823 469 3829 475
rect 5707 469 5713 475
rect 1959 461 1965 467
rect 3823 461 3829 467
rect 85 357 91 363
rect 1947 357 1953 363
rect 3811 353 3817 359
rect 5695 353 5701 359
rect 1947 333 1953 339
rect 3811 333 3817 339
rect 97 205 103 211
rect 1959 205 1965 211
rect 3823 201 3829 207
rect 5707 201 5713 207
rect 1959 185 1965 191
rect 3823 185 3829 191
rect 85 93 91 99
rect 1947 93 1953 99
rect 3811 89 3817 95
rect 5695 89 5701 95
rect 1947 73 1953 79
rect 3811 73 3817 79
<< m5 >>
rect 84 5759 92 5760
rect 84 5753 85 5759
rect 91 5753 92 5759
rect 84 5535 92 5753
rect 84 5529 85 5535
rect 91 5529 92 5535
rect 84 5311 92 5529
rect 84 5305 85 5311
rect 91 5305 92 5311
rect 84 4983 92 5305
rect 84 4977 85 4983
rect 91 4977 92 4983
rect 84 4743 92 4977
rect 84 4737 85 4743
rect 91 4737 92 4743
rect 84 4499 92 4737
rect 84 4493 85 4499
rect 91 4493 92 4499
rect 84 4255 92 4493
rect 84 4249 85 4255
rect 91 4249 92 4255
rect 84 4003 92 4249
rect 84 3997 85 4003
rect 91 3997 92 4003
rect 84 3751 92 3997
rect 84 3745 85 3751
rect 91 3745 92 3751
rect 84 3491 92 3745
rect 84 3485 85 3491
rect 91 3485 92 3491
rect 84 3251 92 3485
rect 84 3245 85 3251
rect 91 3245 92 3251
rect 84 2991 92 3245
rect 84 2985 85 2991
rect 91 2985 92 2991
rect 84 2763 92 2985
rect 84 2757 85 2763
rect 91 2757 92 2763
rect 84 2539 92 2757
rect 84 2533 85 2539
rect 91 2533 92 2539
rect 84 2295 92 2533
rect 84 2289 85 2295
rect 91 2289 92 2295
rect 84 2055 92 2289
rect 84 2049 85 2055
rect 91 2049 92 2055
rect 84 1819 92 2049
rect 84 1813 85 1819
rect 91 1813 92 1819
rect 84 1559 92 1813
rect 84 1553 85 1559
rect 91 1553 92 1559
rect 84 1323 92 1553
rect 84 1317 85 1323
rect 91 1317 92 1323
rect 84 1075 92 1317
rect 84 1069 85 1075
rect 91 1069 92 1075
rect 84 823 92 1069
rect 84 817 85 823
rect 91 817 92 823
rect 84 599 92 817
rect 84 593 85 599
rect 91 593 92 599
rect 84 363 92 593
rect 84 357 85 363
rect 91 357 92 363
rect 84 99 92 357
rect 84 93 85 99
rect 91 93 92 99
rect 84 72 92 93
rect 96 5647 104 5760
rect 96 5641 97 5647
rect 103 5641 104 5647
rect 96 5423 104 5641
rect 96 5417 97 5423
rect 103 5417 104 5423
rect 96 5095 104 5417
rect 96 5089 97 5095
rect 103 5089 104 5095
rect 96 4863 104 5089
rect 96 4857 97 4863
rect 103 4857 104 4863
rect 96 4615 104 4857
rect 96 4609 97 4615
rect 103 4609 104 4615
rect 96 4383 104 4609
rect 96 4377 97 4383
rect 103 4377 104 4383
rect 96 4139 104 4377
rect 96 4133 97 4139
rect 103 4133 104 4139
rect 96 3863 104 4133
rect 96 3857 97 3863
rect 103 3857 104 3863
rect 96 3627 104 3857
rect 96 3621 97 3627
rect 103 3621 104 3627
rect 96 3363 104 3621
rect 96 3357 97 3363
rect 103 3357 104 3363
rect 96 3131 104 3357
rect 96 3125 97 3131
rect 103 3125 104 3131
rect 96 2879 104 3125
rect 96 2873 97 2879
rect 103 2873 104 2879
rect 96 2651 104 2873
rect 96 2645 97 2651
rect 103 2645 104 2651
rect 96 2423 104 2645
rect 96 2417 97 2423
rect 103 2417 104 2423
rect 96 2171 104 2417
rect 96 2165 97 2171
rect 103 2165 104 2171
rect 96 1939 104 2165
rect 96 1933 97 1939
rect 103 1933 104 1939
rect 96 1683 104 1933
rect 96 1677 97 1683
rect 103 1677 104 1683
rect 96 1435 104 1677
rect 96 1429 97 1435
rect 103 1429 104 1435
rect 96 1199 104 1429
rect 96 1193 97 1199
rect 103 1193 104 1199
rect 96 951 104 1193
rect 96 945 97 951
rect 103 945 104 951
rect 96 711 104 945
rect 96 705 97 711
rect 103 705 104 711
rect 96 487 104 705
rect 96 481 97 487
rect 103 481 104 487
rect 96 211 104 481
rect 96 205 97 211
rect 103 205 104 211
rect 96 72 104 205
rect 1946 5759 1954 5760
rect 1946 5753 1947 5759
rect 1953 5753 1954 5759
rect 1946 5659 1954 5753
rect 1946 5653 1947 5659
rect 1953 5653 1954 5659
rect 1946 5535 1954 5653
rect 1946 5529 1947 5535
rect 1953 5529 1954 5535
rect 1946 5433 1954 5529
rect 1946 5427 1947 5433
rect 1953 5427 1954 5433
rect 1946 5311 1954 5427
rect 1946 5305 1947 5311
rect 1953 5305 1954 5311
rect 1946 5203 1954 5305
rect 1946 5197 1947 5203
rect 1953 5197 1954 5203
rect 1946 4983 1954 5197
rect 1946 4977 1947 4983
rect 1953 4977 1954 4983
rect 1946 4947 1954 4977
rect 1946 4941 1947 4947
rect 1953 4941 1954 4947
rect 1946 4743 1954 4941
rect 1946 4737 1947 4743
rect 1953 4737 1954 4743
rect 1946 4695 1954 4737
rect 1946 4689 1947 4695
rect 1953 4689 1954 4695
rect 1946 4499 1954 4689
rect 1946 4493 1947 4499
rect 1953 4493 1954 4499
rect 1946 4459 1954 4493
rect 1946 4453 1947 4459
rect 1953 4453 1954 4459
rect 1946 4255 1954 4453
rect 1946 4249 1947 4255
rect 1953 4249 1954 4255
rect 1946 4219 1954 4249
rect 1946 4213 1947 4219
rect 1953 4213 1954 4219
rect 1946 4003 1954 4213
rect 1946 3997 1947 4003
rect 1953 3997 1954 4003
rect 1946 3971 1954 3997
rect 1946 3965 1947 3971
rect 1953 3965 1954 3971
rect 1946 3751 1954 3965
rect 1946 3745 1947 3751
rect 1953 3745 1954 3751
rect 1946 3731 1954 3745
rect 1946 3725 1947 3731
rect 1953 3725 1954 3731
rect 1946 3491 1954 3725
rect 1946 3485 1947 3491
rect 1953 3485 1954 3491
rect 1946 3251 1954 3485
rect 1946 3245 1947 3251
rect 1953 3245 1954 3251
rect 1946 3223 1954 3245
rect 1946 3217 1947 3223
rect 1953 3217 1954 3223
rect 1946 2991 1954 3217
rect 1946 2985 1947 2991
rect 1953 2985 1954 2991
rect 1946 2975 1954 2985
rect 1946 2969 1947 2975
rect 1953 2969 1954 2975
rect 1946 2763 1954 2969
rect 1946 2757 1947 2763
rect 1953 2757 1954 2763
rect 1946 2739 1954 2757
rect 1946 2733 1947 2739
rect 1953 2733 1954 2739
rect 1946 2539 1954 2733
rect 1946 2533 1947 2539
rect 1953 2533 1954 2539
rect 1946 2479 1954 2533
rect 1946 2473 1947 2479
rect 1953 2473 1954 2479
rect 1946 2295 1954 2473
rect 1946 2289 1947 2295
rect 1953 2289 1954 2295
rect 1946 2239 1954 2289
rect 1946 2233 1947 2239
rect 1953 2233 1954 2239
rect 1946 2055 1954 2233
rect 1946 2049 1947 2055
rect 1953 2049 1954 2055
rect 1946 1999 1954 2049
rect 1946 1993 1947 1999
rect 1953 1993 1954 1999
rect 1946 1819 1954 1993
rect 1946 1813 1947 1819
rect 1953 1813 1954 1819
rect 1946 1755 1954 1813
rect 1946 1749 1947 1755
rect 1953 1749 1954 1755
rect 1946 1559 1954 1749
rect 1946 1553 1947 1559
rect 1953 1553 1954 1559
rect 1946 1503 1954 1553
rect 1946 1497 1947 1503
rect 1953 1497 1954 1503
rect 1946 1323 1954 1497
rect 1946 1317 1947 1323
rect 1953 1317 1954 1323
rect 1946 1247 1954 1317
rect 1946 1241 1947 1247
rect 1953 1241 1954 1247
rect 1946 1075 1954 1241
rect 1946 1069 1947 1075
rect 1953 1069 1954 1075
rect 1946 1007 1954 1069
rect 1946 1001 1947 1007
rect 1953 1001 1954 1007
rect 1946 823 1954 1001
rect 1946 817 1947 823
rect 1953 817 1954 823
rect 1946 599 1954 817
rect 1946 593 1947 599
rect 1953 593 1954 599
rect 1946 579 1954 593
rect 1946 573 1947 579
rect 1953 573 1954 579
rect 1946 363 1954 573
rect 1946 357 1947 363
rect 1953 357 1954 363
rect 1946 339 1954 357
rect 1946 333 1947 339
rect 1953 333 1954 339
rect 1946 99 1954 333
rect 1946 93 1947 99
rect 1953 93 1954 99
rect 1946 79 1954 93
rect 1946 73 1947 79
rect 1953 73 1954 79
rect 1946 72 1954 73
rect 1958 5647 1966 5760
rect 1958 5641 1959 5647
rect 1965 5641 1966 5647
rect 1958 5547 1966 5641
rect 1958 5541 1959 5547
rect 1965 5541 1966 5547
rect 1958 5423 1966 5541
rect 1958 5417 1959 5423
rect 1965 5417 1966 5423
rect 1958 5315 1966 5417
rect 1958 5309 1959 5315
rect 1965 5309 1966 5315
rect 1958 5095 1966 5309
rect 1958 5089 1959 5095
rect 1965 5089 1966 5095
rect 1958 4863 1966 5089
rect 1958 4857 1959 4863
rect 1965 4857 1966 4863
rect 1958 4811 1966 4857
rect 1958 4805 1959 4811
rect 1965 4805 1966 4811
rect 1958 4615 1966 4805
rect 1958 4609 1959 4615
rect 1965 4609 1966 4615
rect 1958 4579 1966 4609
rect 1958 4573 1959 4579
rect 1965 4573 1966 4579
rect 1958 4383 1966 4573
rect 1958 4377 1959 4383
rect 1965 4377 1966 4383
rect 1958 4339 1966 4377
rect 1958 4333 1959 4339
rect 1965 4333 1966 4339
rect 1958 4139 1966 4333
rect 1958 4133 1959 4139
rect 1965 4133 1966 4139
rect 1958 4087 1966 4133
rect 1958 4081 1959 4087
rect 1965 4081 1966 4087
rect 1958 3863 1966 4081
rect 1958 3857 1959 3863
rect 1965 3857 1966 3863
rect 1958 3847 1966 3857
rect 1958 3841 1959 3847
rect 1965 3841 1966 3847
rect 1958 3627 1966 3841
rect 1958 3621 1959 3627
rect 1965 3621 1966 3627
rect 1958 3607 1966 3621
rect 1958 3601 1959 3607
rect 1965 3601 1966 3607
rect 1958 3363 1966 3601
rect 1958 3357 1959 3363
rect 1965 3357 1966 3363
rect 1958 3335 1966 3357
rect 1958 3329 1959 3335
rect 1965 3329 1966 3335
rect 1958 3131 1966 3329
rect 1958 3125 1959 3131
rect 1965 3125 1966 3131
rect 1958 3099 1966 3125
rect 1958 3093 1959 3099
rect 1965 3093 1966 3099
rect 1958 2879 1966 3093
rect 1958 2873 1959 2879
rect 1965 2873 1966 2879
rect 1958 2855 1966 2873
rect 1958 2849 1959 2855
rect 1965 2849 1966 2855
rect 1958 2651 1966 2849
rect 1958 2645 1959 2651
rect 1965 2645 1966 2651
rect 1958 2615 1966 2645
rect 1958 2609 1959 2615
rect 1965 2609 1966 2615
rect 1958 2423 1966 2609
rect 1958 2417 1959 2423
rect 1965 2417 1966 2423
rect 1958 2359 1966 2417
rect 1958 2353 1959 2359
rect 1965 2353 1966 2359
rect 1958 2171 1966 2353
rect 1958 2165 1959 2171
rect 1965 2165 1966 2171
rect 1958 2111 1966 2165
rect 1958 2105 1959 2111
rect 1965 2105 1966 2111
rect 1958 1939 1966 2105
rect 1958 1933 1959 1939
rect 1965 1933 1966 1939
rect 1958 1875 1966 1933
rect 1958 1869 1959 1875
rect 1965 1869 1966 1875
rect 1958 1683 1966 1869
rect 1958 1677 1959 1683
rect 1965 1677 1966 1683
rect 1958 1635 1966 1677
rect 1958 1629 1959 1635
rect 1965 1629 1966 1635
rect 1958 1435 1966 1629
rect 1958 1429 1959 1435
rect 1965 1429 1966 1435
rect 1958 1383 1966 1429
rect 1958 1377 1959 1383
rect 1965 1377 1966 1383
rect 1958 1199 1966 1377
rect 1958 1193 1959 1199
rect 1965 1193 1966 1199
rect 1958 1119 1966 1193
rect 1958 1113 1959 1119
rect 1965 1113 1966 1119
rect 1958 951 1966 1113
rect 1958 945 1959 951
rect 1965 945 1966 951
rect 1958 891 1966 945
rect 1958 885 1959 891
rect 1965 885 1966 891
rect 1958 711 1966 885
rect 1958 705 1959 711
rect 1965 705 1966 711
rect 1958 487 1966 705
rect 1958 481 1959 487
rect 1965 481 1966 487
rect 1958 467 1966 481
rect 1958 461 1959 467
rect 1965 461 1966 467
rect 1958 211 1966 461
rect 1958 205 1959 211
rect 1965 205 1966 211
rect 1958 191 1966 205
rect 1958 185 1959 191
rect 1965 185 1966 191
rect 1958 72 1966 185
rect 3810 5659 3818 5760
rect 3810 5653 3811 5659
rect 3817 5653 3818 5659
rect 3810 5427 3818 5653
rect 3810 5421 3811 5427
rect 3817 5421 3818 5427
rect 3810 5411 3818 5421
rect 3810 5405 3811 5411
rect 3817 5405 3818 5411
rect 3810 5203 3818 5405
rect 3810 5197 3811 5203
rect 3817 5197 3818 5203
rect 3810 5143 3818 5197
rect 3810 5137 3811 5143
rect 3817 5137 3818 5143
rect 3810 4947 3818 5137
rect 3810 4941 3811 4947
rect 3817 4941 3818 4947
rect 3810 4887 3818 4941
rect 3810 4881 3811 4887
rect 3817 4881 3818 4887
rect 3810 4695 3818 4881
rect 3810 4689 3811 4695
rect 3817 4689 3818 4695
rect 3810 4659 3818 4689
rect 3810 4653 3811 4659
rect 3817 4653 3818 4659
rect 3810 4459 3818 4653
rect 3810 4453 3811 4459
rect 3817 4453 3818 4459
rect 3810 4427 3818 4453
rect 3810 4421 3811 4427
rect 3817 4421 3818 4427
rect 3810 4219 3818 4421
rect 3810 4213 3811 4219
rect 3817 4213 3818 4219
rect 3810 4167 3818 4213
rect 3810 4161 3811 4167
rect 3817 4161 3818 4167
rect 3810 3971 3818 4161
rect 3810 3965 3811 3971
rect 3817 3965 3818 3971
rect 3810 3919 3818 3965
rect 3810 3913 3811 3919
rect 3817 3913 3818 3919
rect 3810 3731 3818 3913
rect 3810 3725 3811 3731
rect 3817 3725 3818 3731
rect 3810 3651 3818 3725
rect 3810 3645 3811 3651
rect 3817 3645 3818 3651
rect 3810 3399 3818 3645
rect 3810 3393 3811 3399
rect 3817 3393 3818 3399
rect 3810 3223 3818 3393
rect 3810 3217 3811 3223
rect 3817 3217 3818 3223
rect 3810 3159 3818 3217
rect 3810 3153 3811 3159
rect 3817 3153 3818 3159
rect 3810 2975 3818 3153
rect 3810 2969 3811 2975
rect 3817 2969 3818 2975
rect 3810 2931 3818 2969
rect 3810 2925 3811 2931
rect 3817 2925 3818 2931
rect 3810 2739 3818 2925
rect 3810 2733 3811 2739
rect 3817 2733 3818 2739
rect 3810 2699 3818 2733
rect 3810 2693 3811 2699
rect 3817 2693 3818 2699
rect 3810 2479 3818 2693
rect 3810 2473 3811 2479
rect 3817 2473 3818 2479
rect 3810 2471 3818 2473
rect 3810 2465 3811 2471
rect 3817 2465 3818 2471
rect 3810 2239 3818 2465
rect 3810 2233 3811 2239
rect 3817 2233 3818 2239
rect 3810 2223 3818 2233
rect 3810 2217 3811 2223
rect 3817 2217 3818 2223
rect 3810 1999 3818 2217
rect 3810 1993 3811 1999
rect 3817 1993 3818 1999
rect 3810 1755 3818 1993
rect 3810 1749 3811 1755
rect 3817 1749 3818 1755
rect 3810 1747 3818 1749
rect 3810 1741 3811 1747
rect 3817 1741 3818 1747
rect 3810 1523 3818 1741
rect 3810 1517 3811 1523
rect 3817 1517 3818 1523
rect 3810 1503 3818 1517
rect 3810 1497 3811 1503
rect 3817 1497 3818 1503
rect 3810 1287 3818 1497
rect 3810 1281 3811 1287
rect 3817 1281 3818 1287
rect 3810 1247 3818 1281
rect 3810 1241 3811 1247
rect 3817 1241 3818 1247
rect 3810 1055 3818 1241
rect 3810 1049 3811 1055
rect 3817 1049 3818 1055
rect 3810 1007 3818 1049
rect 3810 1001 3811 1007
rect 3817 1001 3818 1007
rect 3810 827 3818 1001
rect 3810 821 3811 827
rect 3817 821 3818 827
rect 3810 599 3818 821
rect 3810 593 3811 599
rect 3817 593 3818 599
rect 3810 579 3818 593
rect 3810 573 3811 579
rect 3817 573 3818 579
rect 3810 359 3818 573
rect 3810 353 3811 359
rect 3817 353 3818 359
rect 3810 339 3818 353
rect 3810 333 3811 339
rect 3817 333 3818 339
rect 3810 95 3818 333
rect 3810 89 3811 95
rect 3817 89 3818 95
rect 3810 79 3818 89
rect 3810 73 3811 79
rect 3817 73 3818 79
rect 3810 72 3818 73
rect 3822 5547 3830 5760
rect 3822 5541 3823 5547
rect 3829 5541 3830 5547
rect 3822 5315 3830 5541
rect 3822 5309 3823 5315
rect 3829 5309 3830 5315
rect 3822 5283 3830 5309
rect 3822 5277 3823 5283
rect 3829 5277 3830 5283
rect 3822 5019 3830 5277
rect 3822 5013 3823 5019
rect 3829 5013 3830 5019
rect 3822 4811 3830 5013
rect 3822 4805 3823 4811
rect 3829 4805 3830 4811
rect 3822 4771 3830 4805
rect 3822 4765 3823 4771
rect 3829 4765 3830 4771
rect 3822 4579 3830 4765
rect 3822 4573 3823 4579
rect 3829 4573 3830 4579
rect 3822 4547 3830 4573
rect 3822 4541 3823 4547
rect 3829 4541 3830 4547
rect 3822 4339 3830 4541
rect 3822 4333 3823 4339
rect 3829 4333 3830 4339
rect 3822 4315 3830 4333
rect 3822 4309 3823 4315
rect 3829 4309 3830 4315
rect 3822 4087 3830 4309
rect 3822 4081 3823 4087
rect 3829 4081 3830 4087
rect 3822 4055 3830 4081
rect 3822 4049 3823 4055
rect 3829 4049 3830 4055
rect 3822 3847 3830 4049
rect 3822 3841 3823 3847
rect 3829 3841 3830 3847
rect 3822 3791 3830 3841
rect 3822 3785 3823 3791
rect 3829 3785 3830 3791
rect 3822 3607 3830 3785
rect 3822 3601 3823 3607
rect 3829 3601 3830 3607
rect 3822 3515 3830 3601
rect 3822 3509 3823 3515
rect 3829 3509 3830 3515
rect 3822 3335 3830 3509
rect 3822 3329 3823 3335
rect 3829 3329 3830 3335
rect 3822 3287 3830 3329
rect 3822 3281 3823 3287
rect 3829 3281 3830 3287
rect 3822 3099 3830 3281
rect 3822 3093 3823 3099
rect 3829 3093 3830 3099
rect 3822 3047 3830 3093
rect 3822 3041 3823 3047
rect 3829 3041 3830 3047
rect 3822 2855 3830 3041
rect 3822 2849 3823 2855
rect 3829 2849 3830 2855
rect 3822 2811 3830 2849
rect 3822 2805 3823 2811
rect 3829 2805 3830 2811
rect 3822 2615 3830 2805
rect 3822 2609 3823 2615
rect 3829 2609 3830 2615
rect 3822 2587 3830 2609
rect 3822 2581 3823 2587
rect 3829 2581 3830 2587
rect 3822 2359 3830 2581
rect 3822 2353 3823 2359
rect 3829 2353 3830 2359
rect 3822 2347 3830 2353
rect 3822 2341 3823 2347
rect 3829 2341 3830 2347
rect 3822 2111 3830 2341
rect 3822 2105 3823 2111
rect 3829 2105 3830 2111
rect 3822 1875 3830 2105
rect 3822 1869 3823 1875
rect 3829 1869 3830 1875
rect 3822 1635 3830 1869
rect 3822 1629 3823 1635
rect 3829 1629 3830 1635
rect 3822 1407 3830 1629
rect 3822 1401 3823 1407
rect 3829 1401 3830 1407
rect 3822 1383 3830 1401
rect 3822 1377 3823 1383
rect 3829 1377 3830 1383
rect 3822 1171 3830 1377
rect 3822 1165 3823 1171
rect 3829 1165 3830 1171
rect 3822 1119 3830 1165
rect 3822 1113 3823 1119
rect 3829 1113 3830 1119
rect 3822 939 3830 1113
rect 3822 933 3823 939
rect 3829 933 3830 939
rect 3822 891 3830 933
rect 3822 885 3823 891
rect 3829 885 3830 891
rect 3822 711 3830 885
rect 3822 705 3823 711
rect 3829 705 3830 711
rect 3822 475 3830 705
rect 3822 469 3823 475
rect 3829 469 3830 475
rect 3822 467 3830 469
rect 3822 461 3823 467
rect 3829 461 3830 467
rect 3822 207 3830 461
rect 3822 201 3823 207
rect 3829 201 3830 207
rect 3822 191 3830 201
rect 3822 185 3823 191
rect 3829 185 3830 191
rect 3822 72 3830 185
rect 5694 5411 5702 5760
rect 5694 5405 5695 5411
rect 5701 5405 5702 5411
rect 5694 5143 5702 5405
rect 5694 5137 5695 5143
rect 5701 5137 5702 5143
rect 5694 4887 5702 5137
rect 5694 4881 5695 4887
rect 5701 4881 5702 4887
rect 5694 4659 5702 4881
rect 5694 4653 5695 4659
rect 5701 4653 5702 4659
rect 5694 4427 5702 4653
rect 5694 4421 5695 4427
rect 5701 4421 5702 4427
rect 5694 4167 5702 4421
rect 5694 4161 5695 4167
rect 5701 4161 5702 4167
rect 5694 3919 5702 4161
rect 5694 3913 5695 3919
rect 5701 3913 5702 3919
rect 5694 3651 5702 3913
rect 5694 3645 5695 3651
rect 5701 3645 5702 3651
rect 5694 3399 5702 3645
rect 5694 3393 5695 3399
rect 5701 3393 5702 3399
rect 5694 3159 5702 3393
rect 5694 3153 5695 3159
rect 5701 3153 5702 3159
rect 5694 2931 5702 3153
rect 5694 2925 5695 2931
rect 5701 2925 5702 2931
rect 5694 2699 5702 2925
rect 5694 2693 5695 2699
rect 5701 2693 5702 2699
rect 5694 2471 5702 2693
rect 5694 2465 5695 2471
rect 5701 2465 5702 2471
rect 5694 2223 5702 2465
rect 5694 2217 5695 2223
rect 5701 2217 5702 2223
rect 5694 1747 5702 2217
rect 5694 1741 5695 1747
rect 5701 1741 5702 1747
rect 5694 1523 5702 1741
rect 5694 1517 5695 1523
rect 5701 1517 5702 1523
rect 5694 1287 5702 1517
rect 5694 1281 5695 1287
rect 5701 1281 5702 1287
rect 5694 1055 5702 1281
rect 5694 1049 5695 1055
rect 5701 1049 5702 1055
rect 5694 827 5702 1049
rect 5694 821 5695 827
rect 5701 821 5702 827
rect 5694 599 5702 821
rect 5694 593 5695 599
rect 5701 593 5702 599
rect 5694 359 5702 593
rect 5694 353 5695 359
rect 5701 353 5702 359
rect 5694 95 5702 353
rect 5694 89 5695 95
rect 5701 89 5702 95
rect 5694 72 5702 89
rect 5706 5283 5714 5760
rect 5706 5277 5707 5283
rect 5713 5277 5714 5283
rect 5706 5019 5714 5277
rect 5706 5013 5707 5019
rect 5713 5013 5714 5019
rect 5706 4771 5714 5013
rect 5706 4765 5707 4771
rect 5713 4765 5714 4771
rect 5706 4547 5714 4765
rect 5706 4541 5707 4547
rect 5713 4541 5714 4547
rect 5706 4315 5714 4541
rect 5706 4309 5707 4315
rect 5713 4309 5714 4315
rect 5706 4055 5714 4309
rect 5706 4049 5707 4055
rect 5713 4049 5714 4055
rect 5706 3791 5714 4049
rect 5706 3785 5707 3791
rect 5713 3785 5714 3791
rect 5706 3515 5714 3785
rect 5706 3509 5707 3515
rect 5713 3509 5714 3515
rect 5706 3287 5714 3509
rect 5706 3281 5707 3287
rect 5713 3281 5714 3287
rect 5706 3047 5714 3281
rect 5706 3041 5707 3047
rect 5713 3041 5714 3047
rect 5706 2811 5714 3041
rect 5706 2805 5707 2811
rect 5713 2805 5714 2811
rect 5706 2587 5714 2805
rect 5706 2581 5707 2587
rect 5713 2581 5714 2587
rect 5706 2347 5714 2581
rect 5706 2341 5707 2347
rect 5713 2341 5714 2347
rect 5706 1407 5714 2341
rect 5706 1401 5707 1407
rect 5713 1401 5714 1407
rect 5706 1171 5714 1401
rect 5706 1165 5707 1171
rect 5713 1165 5714 1171
rect 5706 939 5714 1165
rect 5706 933 5707 939
rect 5713 933 5714 939
rect 5706 711 5714 933
rect 5706 705 5707 711
rect 5713 705 5714 711
rect 5706 475 5714 705
rect 5706 469 5707 475
rect 5713 469 5714 475
rect 5706 207 5714 469
rect 5706 201 5707 207
rect 5713 201 5714 207
rect 5706 72 5714 201
use circuitwell  npwells
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use circuitppnp  ppnps
timestamp 0
transform 1 0 80 0 1 72
box 0 0 1 1
use welltap_svt  __well_tap__271
timestamp 1731220412
transform 1 0 5656 0 -1 5628
box 7 3 12 24
use welltap_svt  __well_tap__270
timestamp 1731220412
transform 1 0 3832 0 -1 5628
box 7 3 12 24
use welltap_svt  __well_tap__269
timestamp 1731220412
transform 1 0 5656 0 1 5452
box 7 3 12 24
use welltap_svt  __well_tap__268
timestamp 1731220412
transform 1 0 3832 0 1 5452
box 7 3 12 24
use welltap_svt  __well_tap__267
timestamp 1731220412
transform 1 0 5656 0 -1 5384
box 7 3 12 24
use welltap_svt  __well_tap__266
timestamp 1731220412
transform 1 0 3832 0 -1 5384
box 7 3 12 24
use welltap_svt  __well_tap__265
timestamp 1731220412
transform 1 0 5656 0 1 5192
box 7 3 12 24
use welltap_svt  __well_tap__264
timestamp 1731220412
transform 1 0 3832 0 1 5192
box 7 3 12 24
use welltap_svt  __well_tap__263
timestamp 1731220412
transform 1 0 5656 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__262
timestamp 1731220412
transform 1 0 3832 0 -1 5116
box 7 3 12 24
use welltap_svt  __well_tap__261
timestamp 1731220412
transform 1 0 5656 0 1 4928
box 7 3 12 24
use welltap_svt  __well_tap__260
timestamp 1731220412
transform 1 0 3832 0 1 4928
box 7 3 12 24
use welltap_svt  __well_tap__259
timestamp 1731220412
transform 1 0 5656 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__258
timestamp 1731220412
transform 1 0 3832 0 -1 4860
box 7 3 12 24
use welltap_svt  __well_tap__257
timestamp 1731220412
transform 1 0 5656 0 1 4680
box 7 3 12 24
use welltap_svt  __well_tap__256
timestamp 1731220412
transform 1 0 3832 0 1 4680
box 7 3 12 24
use welltap_svt  __well_tap__255
timestamp 1731220412
transform 1 0 5656 0 -1 4632
box 7 3 12 24
use welltap_svt  __well_tap__254
timestamp 1731220412
transform 1 0 3832 0 -1 4632
box 7 3 12 24
use welltap_svt  __well_tap__253
timestamp 1731220412
transform 1 0 5656 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__252
timestamp 1731220412
transform 1 0 3832 0 1 4456
box 7 3 12 24
use welltap_svt  __well_tap__251
timestamp 1731220412
transform 1 0 5656 0 -1 4400
box 7 3 12 24
use welltap_svt  __well_tap__250
timestamp 1731220412
transform 1 0 3832 0 -1 4400
box 7 3 12 24
use welltap_svt  __well_tap__249
timestamp 1731220412
transform 1 0 5656 0 1 4224
box 7 3 12 24
use welltap_svt  __well_tap__248
timestamp 1731220412
transform 1 0 3832 0 1 4224
box 7 3 12 24
use welltap_svt  __well_tap__247
timestamp 1731220412
transform 1 0 5656 0 -1 4140
box 7 3 12 24
use welltap_svt  __well_tap__246
timestamp 1731220412
transform 1 0 3832 0 -1 4140
box 7 3 12 24
use welltap_svt  __well_tap__245
timestamp 1731220412
transform 1 0 5656 0 1 3964
box 7 3 12 24
use welltap_svt  __well_tap__244
timestamp 1731220412
transform 1 0 3832 0 1 3964
box 7 3 12 24
use welltap_svt  __well_tap__243
timestamp 1731220412
transform 1 0 5656 0 -1 3892
box 7 3 12 24
use welltap_svt  __well_tap__242
timestamp 1731220412
transform 1 0 3832 0 -1 3892
box 7 3 12 24
use welltap_svt  __well_tap__241
timestamp 1731220412
transform 1 0 5656 0 1 3700
box 7 3 12 24
use welltap_svt  __well_tap__240
timestamp 1731220412
transform 1 0 3832 0 1 3700
box 7 3 12 24
use welltap_svt  __well_tap__239
timestamp 1731220412
transform 1 0 5656 0 -1 3624
box 7 3 12 24
use welltap_svt  __well_tap__238
timestamp 1731220412
transform 1 0 3832 0 -1 3624
box 7 3 12 24
use welltap_svt  __well_tap__237
timestamp 1731220412
transform 1 0 5656 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__236
timestamp 1731220412
transform 1 0 3832 0 1 3424
box 7 3 12 24
use welltap_svt  __well_tap__235
timestamp 1731220412
transform 1 0 5656 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__234
timestamp 1731220412
transform 1 0 3832 0 -1 3372
box 7 3 12 24
use welltap_svt  __well_tap__233
timestamp 1731220412
transform 1 0 5656 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__232
timestamp 1731220412
transform 1 0 3832 0 1 3196
box 7 3 12 24
use welltap_svt  __well_tap__231
timestamp 1731220412
transform 1 0 5656 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__230
timestamp 1731220412
transform 1 0 3832 0 -1 3132
box 7 3 12 24
use welltap_svt  __well_tap__229
timestamp 1731220412
transform 1 0 5656 0 1 2956
box 7 3 12 24
use welltap_svt  __well_tap__228
timestamp 1731220412
transform 1 0 3832 0 1 2956
box 7 3 12 24
use welltap_svt  __well_tap__227
timestamp 1731220412
transform 1 0 5656 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__226
timestamp 1731220412
transform 1 0 3832 0 -1 2904
box 7 3 12 24
use welltap_svt  __well_tap__225
timestamp 1731220412
transform 1 0 5656 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__224
timestamp 1731220412
transform 1 0 3832 0 1 2720
box 7 3 12 24
use welltap_svt  __well_tap__223
timestamp 1731220412
transform 1 0 5656 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__222
timestamp 1731220412
transform 1 0 3832 0 -1 2672
box 7 3 12 24
use welltap_svt  __well_tap__221
timestamp 1731220412
transform 1 0 5656 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__220
timestamp 1731220412
transform 1 0 3832 0 1 2496
box 7 3 12 24
use welltap_svt  __well_tap__219
timestamp 1731220412
transform 1 0 5656 0 -1 2444
box 7 3 12 24
use welltap_svt  __well_tap__218
timestamp 1731220412
transform 1 0 3832 0 -1 2444
box 7 3 12 24
use welltap_svt  __well_tap__217
timestamp 1731220412
transform 1 0 5656 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__216
timestamp 1731220412
transform 1 0 3832 0 1 2256
box 7 3 12 24
use welltap_svt  __well_tap__215
timestamp 1731220412
transform 1 0 5656 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__214
timestamp 1731220412
transform 1 0 3832 0 -1 2196
box 7 3 12 24
use welltap_svt  __well_tap__213
timestamp 1731220412
transform 1 0 5656 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__212
timestamp 1731220412
transform 1 0 3832 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__211
timestamp 1731220412
transform 1 0 5656 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__210
timestamp 1731220412
transform 1 0 3832 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__209
timestamp 1731220412
transform 1 0 5656 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__208
timestamp 1731220412
transform 1 0 3832 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__207
timestamp 1731220412
transform 1 0 5656 0 -1 1720
box 7 3 12 24
use welltap_svt  __well_tap__206
timestamp 1731220412
transform 1 0 3832 0 -1 1720
box 7 3 12 24
use welltap_svt  __well_tap__205
timestamp 1731220412
transform 1 0 5656 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__204
timestamp 1731220412
transform 1 0 3832 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__203
timestamp 1731220412
transform 1 0 5656 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__202
timestamp 1731220412
transform 1 0 3832 0 -1 1496
box 7 3 12 24
use welltap_svt  __well_tap__201
timestamp 1731220412
transform 1 0 5656 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__200
timestamp 1731220412
transform 1 0 3832 0 1 1316
box 7 3 12 24
use welltap_svt  __well_tap__199
timestamp 1731220412
transform 1 0 5656 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__198
timestamp 1731220412
transform 1 0 3832 0 -1 1260
box 7 3 12 24
use welltap_svt  __well_tap__197
timestamp 1731220412
transform 1 0 5656 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__196
timestamp 1731220412
transform 1 0 3832 0 1 1080
box 7 3 12 24
use welltap_svt  __well_tap__195
timestamp 1731220412
transform 1 0 5656 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__194
timestamp 1731220412
transform 1 0 3832 0 -1 1028
box 7 3 12 24
use welltap_svt  __well_tap__193
timestamp 1731220412
transform 1 0 5656 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__192
timestamp 1731220412
transform 1 0 3832 0 1 848
box 7 3 12 24
use welltap_svt  __well_tap__191
timestamp 1731220412
transform 1 0 5656 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__190
timestamp 1731220412
transform 1 0 3832 0 -1 800
box 7 3 12 24
use welltap_svt  __well_tap__189
timestamp 1731220412
transform 1 0 5656 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__188
timestamp 1731220412
transform 1 0 3832 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__187
timestamp 1731220412
transform 1 0 5656 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__186
timestamp 1731220412
transform 1 0 3832 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__185
timestamp 1731220412
transform 1 0 5656 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__184
timestamp 1731220412
transform 1 0 3832 0 1 384
box 7 3 12 24
use welltap_svt  __well_tap__183
timestamp 1731220412
transform 1 0 5656 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__182
timestamp 1731220412
transform 1 0 3832 0 -1 332
box 7 3 12 24
use welltap_svt  __well_tap__181
timestamp 1731220412
transform 1 0 5656 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__180
timestamp 1731220412
transform 1 0 3832 0 1 116
box 7 3 12 24
use welltap_svt  __well_tap__179
timestamp 1731220412
transform 1 0 3792 0 -1 5632
box 7 3 12 24
use welltap_svt  __well_tap__178
timestamp 1731220412
transform 1 0 1968 0 -1 5632
box 7 3 12 24
use welltap_svt  __well_tap__177
timestamp 1731220412
transform 1 0 3792 0 1 5456
box 7 3 12 24
use welltap_svt  __well_tap__176
timestamp 1731220412
transform 1 0 1968 0 1 5456
box 7 3 12 24
use welltap_svt  __well_tap__175
timestamp 1731220412
transform 1 0 3792 0 -1 5400
box 7 3 12 24
use welltap_svt  __well_tap__174
timestamp 1731220412
transform 1 0 1968 0 -1 5400
box 7 3 12 24
use welltap_svt  __well_tap__173
timestamp 1731220412
transform 1 0 3792 0 1 5224
box 7 3 12 24
use welltap_svt  __well_tap__172
timestamp 1731220412
transform 1 0 1968 0 1 5224
box 7 3 12 24
use welltap_svt  __well_tap__171
timestamp 1731220412
transform 1 0 3792 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__170
timestamp 1731220412
transform 1 0 1968 0 -1 5176
box 7 3 12 24
use welltap_svt  __well_tap__169
timestamp 1731220412
transform 1 0 3792 0 1 5000
box 7 3 12 24
use welltap_svt  __well_tap__168
timestamp 1731220412
transform 1 0 1968 0 1 5000
box 7 3 12 24
use welltap_svt  __well_tap__167
timestamp 1731220412
transform 1 0 3792 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__166
timestamp 1731220412
transform 1 0 1968 0 -1 4920
box 7 3 12 24
use welltap_svt  __well_tap__165
timestamp 1731220412
transform 1 0 3792 0 1 4720
box 7 3 12 24
use welltap_svt  __well_tap__164
timestamp 1731220412
transform 1 0 1968 0 1 4720
box 7 3 12 24
use welltap_svt  __well_tap__163
timestamp 1731220412
transform 1 0 3792 0 -1 4668
box 7 3 12 24
use welltap_svt  __well_tap__162
timestamp 1731220412
transform 1 0 1968 0 -1 4668
box 7 3 12 24
use welltap_svt  __well_tap__161
timestamp 1731220412
transform 1 0 3792 0 1 4488
box 7 3 12 24
use welltap_svt  __well_tap__160
timestamp 1731220412
transform 1 0 1968 0 1 4488
box 7 3 12 24
use welltap_svt  __well_tap__159
timestamp 1731220412
transform 1 0 3792 0 -1 4432
box 7 3 12 24
use welltap_svt  __well_tap__158
timestamp 1731220412
transform 1 0 1968 0 -1 4432
box 7 3 12 24
use welltap_svt  __well_tap__157
timestamp 1731220412
transform 1 0 3792 0 1 4248
box 7 3 12 24
use welltap_svt  __well_tap__156
timestamp 1731220412
transform 1 0 1968 0 1 4248
box 7 3 12 24
use welltap_svt  __well_tap__155
timestamp 1731220412
transform 1 0 3792 0 -1 4192
box 7 3 12 24
use welltap_svt  __well_tap__154
timestamp 1731220412
transform 1 0 1968 0 -1 4192
box 7 3 12 24
use welltap_svt  __well_tap__153
timestamp 1731220412
transform 1 0 3792 0 1 3996
box 7 3 12 24
use welltap_svt  __well_tap__152
timestamp 1731220412
transform 1 0 1968 0 1 3996
box 7 3 12 24
use welltap_svt  __well_tap__151
timestamp 1731220412
transform 1 0 3792 0 -1 3944
box 7 3 12 24
use welltap_svt  __well_tap__150
timestamp 1731220412
transform 1 0 1968 0 -1 3944
box 7 3 12 24
use welltap_svt  __well_tap__149
timestamp 1731220412
transform 1 0 3792 0 1 3756
box 7 3 12 24
use welltap_svt  __well_tap__148
timestamp 1731220412
transform 1 0 1968 0 1 3756
box 7 3 12 24
use welltap_svt  __well_tap__147
timestamp 1731220412
transform 1 0 3792 0 -1 3704
box 7 3 12 24
use welltap_svt  __well_tap__146
timestamp 1731220412
transform 1 0 1968 0 -1 3704
box 7 3 12 24
use welltap_svt  __well_tap__145
timestamp 1731220412
transform 1 0 3792 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__144
timestamp 1731220412
transform 1 0 1968 0 1 3516
box 7 3 12 24
use welltap_svt  __well_tap__143
timestamp 1731220412
transform 1 0 3792 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__142
timestamp 1731220412
transform 1 0 1968 0 -1 3460
box 7 3 12 24
use welltap_svt  __well_tap__141
timestamp 1731220412
transform 1 0 3792 0 1 3244
box 7 3 12 24
use welltap_svt  __well_tap__140
timestamp 1731220412
transform 1 0 1968 0 1 3244
box 7 3 12 24
use welltap_svt  __well_tap__139
timestamp 1731220412
transform 1 0 3792 0 -1 3196
box 7 3 12 24
use welltap_svt  __well_tap__138
timestamp 1731220412
transform 1 0 1968 0 -1 3196
box 7 3 12 24
use welltap_svt  __well_tap__137
timestamp 1731220412
transform 1 0 3792 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__136
timestamp 1731220412
transform 1 0 1968 0 1 3008
box 7 3 12 24
use welltap_svt  __well_tap__135
timestamp 1731220412
transform 1 0 3792 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__134
timestamp 1731220412
transform 1 0 1968 0 -1 2948
box 7 3 12 24
use welltap_svt  __well_tap__133
timestamp 1731220412
transform 1 0 3792 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__132
timestamp 1731220412
transform 1 0 1968 0 1 2764
box 7 3 12 24
use welltap_svt  __well_tap__131
timestamp 1731220412
transform 1 0 3792 0 -1 2712
box 7 3 12 24
use welltap_svt  __well_tap__130
timestamp 1731220412
transform 1 0 1968 0 -1 2712
box 7 3 12 24
use welltap_svt  __well_tap__129
timestamp 1731220412
transform 1 0 3792 0 1 2524
box 7 3 12 24
use welltap_svt  __well_tap__128
timestamp 1731220412
transform 1 0 1968 0 1 2524
box 7 3 12 24
use welltap_svt  __well_tap__127
timestamp 1731220412
transform 1 0 3792 0 -1 2452
box 7 3 12 24
use welltap_svt  __well_tap__126
timestamp 1731220412
transform 1 0 1968 0 -1 2452
box 7 3 12 24
use welltap_svt  __well_tap__125
timestamp 1731220412
transform 1 0 3792 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__124
timestamp 1731220412
transform 1 0 1968 0 1 2268
box 7 3 12 24
use welltap_svt  __well_tap__123
timestamp 1731220412
transform 1 0 3792 0 -1 2212
box 7 3 12 24
use welltap_svt  __well_tap__122
timestamp 1731220412
transform 1 0 1968 0 -1 2212
box 7 3 12 24
use welltap_svt  __well_tap__121
timestamp 1731220412
transform 1 0 3792 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__120
timestamp 1731220412
transform 1 0 1968 0 1 2020
box 7 3 12 24
use welltap_svt  __well_tap__119
timestamp 1731220412
transform 1 0 3792 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__118
timestamp 1731220412
transform 1 0 1968 0 -1 1972
box 7 3 12 24
use welltap_svt  __well_tap__117
timestamp 1731220412
transform 1 0 3792 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__116
timestamp 1731220412
transform 1 0 1968 0 1 1784
box 7 3 12 24
use welltap_svt  __well_tap__115
timestamp 1731220412
transform 1 0 3792 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__114
timestamp 1731220412
transform 1 0 1968 0 -1 1728
box 7 3 12 24
use welltap_svt  __well_tap__113
timestamp 1731220412
transform 1 0 3792 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__112
timestamp 1731220412
transform 1 0 1968 0 1 1544
box 7 3 12 24
use welltap_svt  __well_tap__111
timestamp 1731220412
transform 1 0 3792 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__110
timestamp 1731220412
transform 1 0 1968 0 -1 1476
box 7 3 12 24
use welltap_svt  __well_tap__109
timestamp 1731220412
transform 1 0 3792 0 1 1292
box 7 3 12 24
use welltap_svt  __well_tap__108
timestamp 1731220412
transform 1 0 1968 0 1 1292
box 7 3 12 24
use welltap_svt  __well_tap__107
timestamp 1731220412
transform 1 0 3792 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__106
timestamp 1731220412
transform 1 0 1968 0 -1 1220
box 7 3 12 24
use welltap_svt  __well_tap__105
timestamp 1731220412
transform 1 0 3792 0 1 1028
box 7 3 12 24
use welltap_svt  __well_tap__104
timestamp 1731220412
transform 1 0 1968 0 1 1028
box 7 3 12 24
use welltap_svt  __well_tap__103
timestamp 1731220412
transform 1 0 3792 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__102
timestamp 1731220412
transform 1 0 1968 0 -1 980
box 7 3 12 24
use welltap_svt  __well_tap__101
timestamp 1731220412
transform 1 0 3792 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__100
timestamp 1731220412
transform 1 0 1968 0 1 800
box 7 3 12 24
use welltap_svt  __well_tap__99
timestamp 1731220412
transform 1 0 3792 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__98
timestamp 1731220412
transform 1 0 1968 0 -1 552
box 7 3 12 24
use welltap_svt  __well_tap__97
timestamp 1731220412
transform 1 0 3792 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__96
timestamp 1731220412
transform 1 0 1968 0 1 376
box 7 3 12 24
use welltap_svt  __well_tap__95
timestamp 1731220412
transform 1 0 3792 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__94
timestamp 1731220412
transform 1 0 1968 0 -1 312
box 7 3 12 24
use welltap_svt  __well_tap__93
timestamp 1731220412
transform 1 0 3792 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__92
timestamp 1731220412
transform 1 0 1968 0 1 100
box 7 3 12 24
use welltap_svt  __well_tap__91
timestamp 1731220412
transform 1 0 1928 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__90
timestamp 1731220412
transform 1 0 104 0 -1 5732
box 7 3 12 24
use welltap_svt  __well_tap__89
timestamp 1731220412
transform 1 0 1928 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__88
timestamp 1731220412
transform 1 0 104 0 1 5556
box 7 3 12 24
use welltap_svt  __well_tap__87
timestamp 1731220412
transform 1 0 1928 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__86
timestamp 1731220412
transform 1 0 104 0 -1 5508
box 7 3 12 24
use welltap_svt  __well_tap__85
timestamp 1731220412
transform 1 0 1928 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__84
timestamp 1731220412
transform 1 0 104 0 1 5332
box 7 3 12 24
use welltap_svt  __well_tap__83
timestamp 1731220412
transform 1 0 1928 0 -1 5284
box 7 3 12 24
use welltap_svt  __well_tap__82
timestamp 1731220412
transform 1 0 104 0 -1 5284
box 7 3 12 24
use welltap_svt  __well_tap__81
timestamp 1731220412
transform 1 0 1928 0 1 5004
box 7 3 12 24
use welltap_svt  __well_tap__80
timestamp 1731220412
transform 1 0 104 0 1 5004
box 7 3 12 24
use welltap_svt  __well_tap__79
timestamp 1731220412
transform 1 0 1928 0 -1 4956
box 7 3 12 24
use welltap_svt  __well_tap__78
timestamp 1731220412
transform 1 0 104 0 -1 4956
box 7 3 12 24
use welltap_svt  __well_tap__77
timestamp 1731220412
transform 1 0 1928 0 1 4772
box 7 3 12 24
use welltap_svt  __well_tap__76
timestamp 1731220412
transform 1 0 104 0 1 4772
box 7 3 12 24
use welltap_svt  __well_tap__75
timestamp 1731220412
transform 1 0 1928 0 -1 4716
box 7 3 12 24
use welltap_svt  __well_tap__74
timestamp 1731220412
transform 1 0 104 0 -1 4716
box 7 3 12 24
use welltap_svt  __well_tap__73
timestamp 1731220412
transform 1 0 1928 0 1 4524
box 7 3 12 24
use welltap_svt  __well_tap__72
timestamp 1731220412
transform 1 0 104 0 1 4524
box 7 3 12 24
use welltap_svt  __well_tap__71
timestamp 1731220412
transform 1 0 1928 0 -1 4472
box 7 3 12 24
use welltap_svt  __well_tap__70
timestamp 1731220412
transform 1 0 104 0 -1 4472
box 7 3 12 24
use welltap_svt  __well_tap__69
timestamp 1731220412
transform 1 0 1928 0 1 4292
box 7 3 12 24
use welltap_svt  __well_tap__68
timestamp 1731220412
transform 1 0 104 0 1 4292
box 7 3 12 24
use welltap_svt  __well_tap__67
timestamp 1731220412
transform 1 0 1928 0 -1 4228
box 7 3 12 24
use welltap_svt  __well_tap__66
timestamp 1731220412
transform 1 0 104 0 -1 4228
box 7 3 12 24
use welltap_svt  __well_tap__65
timestamp 1731220412
transform 1 0 1928 0 1 4048
box 7 3 12 24
use welltap_svt  __well_tap__64
timestamp 1731220412
transform 1 0 104 0 1 4048
box 7 3 12 24
use welltap_svt  __well_tap__63
timestamp 1731220412
transform 1 0 1928 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__62
timestamp 1731220412
transform 1 0 104 0 -1 3976
box 7 3 12 24
use welltap_svt  __well_tap__61
timestamp 1731220412
transform 1 0 1928 0 1 3772
box 7 3 12 24
use welltap_svt  __well_tap__60
timestamp 1731220412
transform 1 0 104 0 1 3772
box 7 3 12 24
use welltap_svt  __well_tap__59
timestamp 1731220412
transform 1 0 1928 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__58
timestamp 1731220412
transform 1 0 104 0 -1 3724
box 7 3 12 24
use welltap_svt  __well_tap__57
timestamp 1731220412
transform 1 0 1928 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__56
timestamp 1731220412
transform 1 0 104 0 1 3536
box 7 3 12 24
use welltap_svt  __well_tap__55
timestamp 1731220412
transform 1 0 1928 0 -1 3464
box 7 3 12 24
use welltap_svt  __well_tap__54
timestamp 1731220412
transform 1 0 104 0 -1 3464
box 7 3 12 24
use welltap_svt  __well_tap__53
timestamp 1731220412
transform 1 0 1928 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__52
timestamp 1731220412
transform 1 0 104 0 1 3272
box 7 3 12 24
use welltap_svt  __well_tap__51
timestamp 1731220412
transform 1 0 1928 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__50
timestamp 1731220412
transform 1 0 104 0 -1 3224
box 7 3 12 24
use welltap_svt  __well_tap__49
timestamp 1731220412
transform 1 0 1928 0 1 3040
box 7 3 12 24
use welltap_svt  __well_tap__48
timestamp 1731220412
transform 1 0 104 0 1 3040
box 7 3 12 24
use welltap_svt  __well_tap__47
timestamp 1731220412
transform 1 0 1928 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__46
timestamp 1731220412
transform 1 0 104 0 -1 2964
box 7 3 12 24
use welltap_svt  __well_tap__45
timestamp 1731220412
transform 1 0 1928 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__44
timestamp 1731220412
transform 1 0 104 0 1 2788
box 7 3 12 24
use welltap_svt  __well_tap__43
timestamp 1731220412
transform 1 0 1928 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__42
timestamp 1731220412
transform 1 0 104 0 -1 2736
box 7 3 12 24
use welltap_svt  __well_tap__41
timestamp 1731220412
transform 1 0 1928 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__40
timestamp 1731220412
transform 1 0 104 0 1 2560
box 7 3 12 24
use welltap_svt  __well_tap__39
timestamp 1731220412
transform 1 0 1928 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__38
timestamp 1731220412
transform 1 0 104 0 -1 2512
box 7 3 12 24
use welltap_svt  __well_tap__37
timestamp 1731220412
transform 1 0 1928 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__36
timestamp 1731220412
transform 1 0 104 0 1 2332
box 7 3 12 24
use welltap_svt  __well_tap__35
timestamp 1731220412
transform 1 0 1928 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__34
timestamp 1731220412
transform 1 0 104 0 -1 2268
box 7 3 12 24
use welltap_svt  __well_tap__33
timestamp 1731220412
transform 1 0 1928 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__32
timestamp 1731220412
transform 1 0 104 0 1 2080
box 7 3 12 24
use welltap_svt  __well_tap__31
timestamp 1731220412
transform 1 0 1928 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__30
timestamp 1731220412
transform 1 0 104 0 -1 2028
box 7 3 12 24
use welltap_svt  __well_tap__29
timestamp 1731220412
transform 1 0 1928 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__28
timestamp 1731220412
transform 1 0 104 0 1 1848
box 7 3 12 24
use welltap_svt  __well_tap__27
timestamp 1731220412
transform 1 0 1928 0 -1 1792
box 7 3 12 24
use welltap_svt  __well_tap__26
timestamp 1731220412
transform 1 0 104 0 -1 1792
box 7 3 12 24
use welltap_svt  __well_tap__25
timestamp 1731220412
transform 1 0 1928 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__24
timestamp 1731220412
transform 1 0 104 0 1 1592
box 7 3 12 24
use welltap_svt  __well_tap__23
timestamp 1731220412
transform 1 0 1928 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__22
timestamp 1731220412
transform 1 0 104 0 -1 1532
box 7 3 12 24
use welltap_svt  __well_tap__21
timestamp 1731220412
transform 1 0 1928 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__20
timestamp 1731220412
transform 1 0 104 0 1 1344
box 7 3 12 24
use welltap_svt  __well_tap__19
timestamp 1731220412
transform 1 0 1928 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__18
timestamp 1731220412
transform 1 0 104 0 -1 1296
box 7 3 12 24
use welltap_svt  __well_tap__17
timestamp 1731220412
transform 1 0 1928 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__16
timestamp 1731220412
transform 1 0 104 0 1 1108
box 7 3 12 24
use welltap_svt  __well_tap__15
timestamp 1731220412
transform 1 0 1928 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__14
timestamp 1731220412
transform 1 0 104 0 -1 1048
box 7 3 12 24
use welltap_svt  __well_tap__13
timestamp 1731220412
transform 1 0 1928 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__12
timestamp 1731220412
transform 1 0 104 0 1 860
box 7 3 12 24
use welltap_svt  __well_tap__11
timestamp 1731220412
transform 1 0 1928 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__10
timestamp 1731220412
transform 1 0 104 0 -1 796
box 7 3 12 24
use welltap_svt  __well_tap__9
timestamp 1731220412
transform 1 0 1928 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__8
timestamp 1731220412
transform 1 0 104 0 1 620
box 7 3 12 24
use welltap_svt  __well_tap__7
timestamp 1731220412
transform 1 0 1928 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__6
timestamp 1731220412
transform 1 0 104 0 -1 572
box 7 3 12 24
use welltap_svt  __well_tap__5
timestamp 1731220412
transform 1 0 1928 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__4
timestamp 1731220412
transform 1 0 104 0 1 396
box 7 3 12 24
use welltap_svt  __well_tap__3
timestamp 1731220412
transform 1 0 1928 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__2
timestamp 1731220412
transform 1 0 104 0 -1 336
box 7 3 12 24
use welltap_svt  __well_tap__1
timestamp 1731220412
transform 1 0 1928 0 1 120
box 7 3 12 24
use welltap_svt  __well_tap__0
timestamp 1731220412
transform 1 0 104 0 1 120
box 7 3 12 24
use _0_0std_0_0cells_0_0FAX1  tst_5999_6
timestamp 1731220412
transform 1 0 5376 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5998_6
timestamp 1731220412
transform 1 0 5512 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5997_6
timestamp 1731220412
transform 1 0 5496 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5996_6
timestamp 1731220412
transform 1 0 5480 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5995_6
timestamp 1731220412
transform 1 0 5416 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5994_6
timestamp 1731220412
transform 1 0 5264 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5993_6
timestamp 1731220412
transform 1 0 5240 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5992_6
timestamp 1731220412
transform 1 0 5104 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5991_6
timestamp 1731220412
transform 1 0 4968 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5990_6
timestamp 1731220412
transform 1 0 4832 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5989_6
timestamp 1731220412
transform 1 0 4696 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5988_6
timestamp 1731220412
transform 1 0 4560 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5987_6
timestamp 1731220412
transform 1 0 4424 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5986_6
timestamp 1731220412
transform 1 0 4288 0 1 92
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5985_6
timestamp 1731220412
transform 1 0 5296 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5984_6
timestamp 1731220412
transform 1 0 5104 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5983_6
timestamp 1731220412
transform 1 0 4920 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5982_6
timestamp 1731220412
transform 1 0 4744 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5981_6
timestamp 1731220412
transform 1 0 4584 0 -1 356
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5980_6
timestamp 1731220412
transform 1 0 5048 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5979_6
timestamp 1731220412
transform 1 0 4840 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5978_6
timestamp 1731220412
transform 1 0 4640 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5977_6
timestamp 1731220412
transform 1 0 4448 0 1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5976_6
timestamp 1731220412
transform 1 0 5120 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5975_6
timestamp 1731220412
transform 1 0 4824 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5974_6
timestamp 1731220412
transform 1 0 4544 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5973_6
timestamp 1731220412
transform 1 0 4280 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5972_6
timestamp 1731220412
transform 1 0 4040 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5971_6
timestamp 1731220412
transform 1 0 5312 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5970_6
timestamp 1731220412
transform 1 0 5096 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5969_6
timestamp 1731220412
transform 1 0 4888 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5968_6
timestamp 1731220412
transform 1 0 4696 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5967_6
timestamp 1731220412
transform 1 0 4536 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5966_6
timestamp 1731220412
transform 1 0 4536 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5965_6
timestamp 1731220412
transform 1 0 4400 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5964_6
timestamp 1731220412
transform 1 0 4264 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5963_6
timestamp 1731220412
transform 1 0 4128 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5962_6
timestamp 1731220412
transform 1 0 3992 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5961_6
timestamp 1731220412
transform 1 0 3992 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5960_6
timestamp 1731220412
transform 1 0 4168 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5959_6
timestamp 1731220412
transform 1 0 4688 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5958_6
timestamp 1731220412
transform 1 0 4864 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5957_6
timestamp 1731220412
transform 1 0 5256 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5956_6
timestamp 1731220412
transform 1 0 5056 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5955_6
timestamp 1731220412
transform 1 0 4928 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5954_6
timestamp 1731220412
transform 1 0 4640 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5953_6
timestamp 1731220412
transform 1 0 4384 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5952_6
timestamp 1731220412
transform 1 0 5232 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5951_6
timestamp 1731220412
transform 1 0 5048 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5950_6
timestamp 1731220412
transform 1 0 4912 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5949_6
timestamp 1731220412
transform 1 0 4776 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5948_6
timestamp 1731220412
transform 1 0 5184 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5947_6
timestamp 1731220412
transform 1 0 5320 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5946_6
timestamp 1731220412
transform 1 0 5376 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5945_6
timestamp 1731220412
transform 1 0 5240 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5944_6
timestamp 1731220412
transform 1 0 5104 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5943_6
timestamp 1731220412
transform 1 0 4968 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5942_6
timestamp 1731220412
transform 1 0 4832 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5941_6
timestamp 1731220412
transform 1 0 5136 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5940_6
timestamp 1731220412
transform 1 0 4944 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5939_6
timestamp 1731220412
transform 1 0 4760 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5938_6
timestamp 1731220412
transform 1 0 4584 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5937_6
timestamp 1731220412
transform 1 0 5184 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5936_6
timestamp 1731220412
transform 1 0 4872 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5935_6
timestamp 1731220412
transform 1 0 4576 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5934_6
timestamp 1731220412
transform 1 0 4304 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5933_6
timestamp 1731220412
transform 1 0 4056 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5932_6
timestamp 1731220412
transform 1 0 5192 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5931_6
timestamp 1731220412
transform 1 0 4936 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5930_6
timestamp 1731220412
transform 1 0 4688 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5929_6
timestamp 1731220412
transform 1 0 4464 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5928_6
timestamp 1731220412
transform 1 0 4352 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5927_6
timestamp 1731220412
transform 1 0 4272 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5926_6
timestamp 1731220412
transform 1 0 3992 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5925_6
timestamp 1731220412
transform 1 0 3856 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5924_6
timestamp 1731220412
transform 1 0 4584 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5923_6
timestamp 1731220412
transform 1 0 5128 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5922_6
timestamp 1731220412
transform 1 0 4848 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5921_6
timestamp 1731220412
transform 1 0 4744 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5920_6
timestamp 1731220412
transform 1 0 4504 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5919_6
timestamp 1731220412
transform 1 0 4272 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5918_6
timestamp 1731220412
transform 1 0 4992 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5917_6
timestamp 1731220412
transform 1 0 4960 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5916_6
timestamp 1731220412
transform 1 0 4816 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5915_6
timestamp 1731220412
transform 1 0 4672 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5914_6
timestamp 1731220412
transform 1 0 4832 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5913_6
timestamp 1731220412
transform 1 0 4968 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5912_6
timestamp 1731220412
transform 1 0 5104 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5911_6
timestamp 1731220412
transform 1 0 5176 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5910_6
timestamp 1731220412
transform 1 0 5240 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5909_6
timestamp 1731220412
transform 1 0 5376 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5908_6
timestamp 1731220412
transform 1 0 5240 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5907_6
timestamp 1731220412
transform 1 0 5104 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5906_6
timestamp 1731220412
transform 1 0 5248 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5905_6
timestamp 1731220412
transform 1 0 5416 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5904_6
timestamp 1731220412
transform 1 0 5336 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5903_6
timestamp 1731220412
transform 1 0 5456 0 -1 1052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5902_6
timestamp 1731220412
transform 1 0 5456 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5901_6
timestamp 1731220412
transform 1 0 5512 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5900_6
timestamp 1731220412
transform 1 0 5512 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5899_6
timestamp 1731220412
transform 1 0 5512 0 1 1056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5898_6
timestamp 1731220412
transform 1 0 5512 0 -1 1284
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5897_6
timestamp 1731220412
transform 1 0 5496 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5896_6
timestamp 1731220412
transform 1 0 5456 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5895_6
timestamp 1731220412
transform 1 0 5504 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5894_6
timestamp 1731220412
transform 1 0 5376 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5893_6
timestamp 1731220412
transform 1 0 5512 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5892_6
timestamp 1731220412
transform 1 0 5512 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5891_6
timestamp 1731220412
transform 1 0 5512 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5890_6
timestamp 1731220412
transform 1 0 5512 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5889_6
timestamp 1731220412
transform 1 0 5336 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5888_6
timestamp 1731220412
transform 1 0 5368 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5887_6
timestamp 1731220412
transform 1 0 5320 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5886_6
timestamp 1731220412
transform 1 0 5368 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5885_6
timestamp 1731220412
transform 1 0 5080 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5884_6
timestamp 1731220412
transform 1 0 4792 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5883_6
timestamp 1731220412
transform 1 0 4824 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5882_6
timestamp 1731220412
transform 1 0 5072 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5881_6
timestamp 1731220412
transform 1 0 5088 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5880_6
timestamp 1731220412
transform 1 0 4960 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5879_6
timestamp 1731220412
transform 1 0 5144 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5878_6
timestamp 1731220412
transform 1 0 5304 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5877_6
timestamp 1731220412
transform 1 0 5088 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5876_6
timestamp 1731220412
transform 1 0 5040 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5875_6
timestamp 1731220412
transform 1 0 4904 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5874_6
timestamp 1731220412
transform 1 0 4768 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5873_6
timestamp 1731220412
transform 1 0 4632 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5872_6
timestamp 1731220412
transform 1 0 4512 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5871_6
timestamp 1731220412
transform 1 0 4688 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5870_6
timestamp 1731220412
transform 1 0 4880 0 -1 2220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5869_6
timestamp 1731220412
transform 1 0 4784 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5868_6
timestamp 1731220412
transform 1 0 4608 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5867_6
timestamp 1731220412
transform 1 0 4440 0 1 2232
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5866_6
timestamp 1731220412
transform 1 0 4816 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5865_6
timestamp 1731220412
transform 1 0 4552 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5864_6
timestamp 1731220412
transform 1 0 4296 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5863_6
timestamp 1731220412
transform 1 0 4328 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5862_6
timestamp 1731220412
transform 1 0 4576 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5861_6
timestamp 1731220412
transform 1 0 4512 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5860_6
timestamp 1731220412
transform 1 0 4224 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5859_6
timestamp 1731220412
transform 1 0 4808 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5858_6
timestamp 1731220412
transform 1 0 4672 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5857_6
timestamp 1731220412
transform 1 0 4536 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5856_6
timestamp 1731220412
transform 1 0 4400 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5855_6
timestamp 1731220412
transform 1 0 4264 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5854_6
timestamp 1731220412
transform 1 0 4128 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5853_6
timestamp 1731220412
transform 1 0 4000 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5852_6
timestamp 1731220412
transform 1 0 4136 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5851_6
timestamp 1731220412
transform 1 0 4544 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5850_6
timestamp 1731220412
transform 1 0 4408 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5849_6
timestamp 1731220412
transform 1 0 4272 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5848_6
timestamp 1731220412
transform 1 0 4240 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5847_6
timestamp 1731220412
transform 1 0 4072 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5846_6
timestamp 1731220412
transform 1 0 4752 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5845_6
timestamp 1731220412
transform 1 0 4576 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5844_6
timestamp 1731220412
transform 1 0 4408 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5843_6
timestamp 1731220412
transform 1 0 4328 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5842_6
timestamp 1731220412
transform 1 0 4104 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5841_6
timestamp 1731220412
transform 1 0 5000 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5840_6
timestamp 1731220412
transform 1 0 4776 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5839_6
timestamp 1731220412
transform 1 0 4552 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5838_6
timestamp 1731220412
transform 1 0 4344 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5837_6
timestamp 1731220412
transform 1 0 4096 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5836_6
timestamp 1731220412
transform 1 0 4576 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5835_6
timestamp 1731220412
transform 1 0 4784 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5834_6
timestamp 1731220412
transform 1 0 4984 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5833_6
timestamp 1731220412
transform 1 0 5296 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5832_6
timestamp 1731220412
transform 1 0 5080 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5831_6
timestamp 1731220412
transform 1 0 4864 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5830_6
timestamp 1731220412
transform 1 0 4640 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5829_6
timestamp 1731220412
transform 1 0 4392 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5828_6
timestamp 1731220412
transform 1 0 5168 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5827_6
timestamp 1731220412
transform 1 0 5000 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5826_6
timestamp 1731220412
transform 1 0 4840 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5825_6
timestamp 1731220412
transform 1 0 4680 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5824_6
timestamp 1731220412
transform 1 0 4528 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5823_6
timestamp 1731220412
transform 1 0 5040 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5822_6
timestamp 1731220412
transform 1 0 4800 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5821_6
timestamp 1731220412
transform 1 0 4576 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5820_6
timestamp 1731220412
transform 1 0 4368 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5819_6
timestamp 1731220412
transform 1 0 4184 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5818_6
timestamp 1731220412
transform 1 0 4688 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5817_6
timestamp 1731220412
transform 1 0 4432 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5816_6
timestamp 1731220412
transform 1 0 4200 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5815_6
timestamp 1731220412
transform 1 0 3992 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5814_6
timestamp 1731220412
transform 1 0 4960 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5813_6
timestamp 1731220412
transform 1 0 5032 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5812_6
timestamp 1731220412
transform 1 0 4792 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5811_6
timestamp 1731220412
transform 1 0 4568 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5810_6
timestamp 1731220412
transform 1 0 4352 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5809_6
timestamp 1731220412
transform 1 0 4336 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5808_6
timestamp 1731220412
transform 1 0 4496 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5807_6
timestamp 1731220412
transform 1 0 4648 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5806_6
timestamp 1731220412
transform 1 0 4800 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5805_6
timestamp 1731220412
transform 1 0 4944 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5804_6
timestamp 1731220412
transform 1 0 5088 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5803_6
timestamp 1731220412
transform 1 0 5232 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5802_6
timestamp 1731220412
transform 1 0 5376 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5801_6
timestamp 1731220412
transform 1 0 5280 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5800_6
timestamp 1731220412
transform 1 0 5248 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5799_6
timestamp 1731220412
transform 1 0 5288 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5798_6
timestamp 1731220412
transform 1 0 5344 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5797_6
timestamp 1731220412
transform 1 0 5168 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5796_6
timestamp 1731220412
transform 1 0 5352 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5795_6
timestamp 1731220412
transform 1 0 5512 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5794_6
timestamp 1731220412
transform 1 0 5512 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5793_6
timestamp 1731220412
transform 1 0 5512 0 1 3400
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5792_6
timestamp 1731220412
transform 1 0 5512 0 -1 3648
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5791_6
timestamp 1731220412
transform 1 0 5512 0 1 3676
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5790_6
timestamp 1731220412
transform 1 0 5512 0 -1 3916
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5789_6
timestamp 1731220412
transform 1 0 5512 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5788_6
timestamp 1731220412
transform 1 0 5512 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5787_6
timestamp 1731220412
transform 1 0 5496 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5786_6
timestamp 1731220412
transform 1 0 5472 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5785_6
timestamp 1731220412
transform 1 0 5440 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5784_6
timestamp 1731220412
transform 1 0 5408 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5783_6
timestamp 1731220412
transform 1 0 5368 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5782_6
timestamp 1731220412
transform 1 0 5376 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5781_6
timestamp 1731220412
transform 1 0 5152 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5780_6
timestamp 1731220412
transform 1 0 5064 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5779_6
timestamp 1731220412
transform 1 0 5296 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5778_6
timestamp 1731220412
transform 1 0 5208 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5777_6
timestamp 1731220412
transform 1 0 4928 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5776_6
timestamp 1731220412
transform 1 0 4712 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5775_6
timestamp 1731220412
transform 1 0 4944 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5774_6
timestamp 1731220412
transform 1 0 5184 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5773_6
timestamp 1731220412
transform 1 0 5096 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5772_6
timestamp 1731220412
transform 1 0 4880 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5771_6
timestamp 1731220412
transform 1 0 4664 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5770_6
timestamp 1731220412
transform 1 0 4704 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5769_6
timestamp 1731220412
transform 1 0 4856 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5768_6
timestamp 1731220412
transform 1 0 5016 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5767_6
timestamp 1731220412
transform 1 0 4984 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5766_6
timestamp 1731220412
transform 1 0 4848 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5765_6
timestamp 1731220412
transform 1 0 4712 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5764_6
timestamp 1731220412
transform 1 0 4576 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5763_6
timestamp 1731220412
transform 1 0 4440 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5762_6
timestamp 1731220412
transform 1 0 4304 0 -1 5652
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5761_6
timestamp 1731220412
transform 1 0 4248 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5760_6
timestamp 1731220412
transform 1 0 4400 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5759_6
timestamp 1731220412
transform 1 0 4552 0 1 5428
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5758_6
timestamp 1731220412
transform 1 0 4456 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5757_6
timestamp 1731220412
transform 1 0 4248 0 -1 5408
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5756_6
timestamp 1731220412
transform 1 0 4248 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5755_6
timestamp 1731220412
transform 1 0 4480 0 1 5168
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5754_6
timestamp 1731220412
transform 1 0 4376 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5753_6
timestamp 1731220412
transform 1 0 4104 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5752_6
timestamp 1731220412
transform 1 0 4648 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5751_6
timestamp 1731220412
transform 1 0 4624 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5750_6
timestamp 1731220412
transform 1 0 4408 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5749_6
timestamp 1731220412
transform 1 0 4840 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5748_6
timestamp 1731220412
transform 1 0 4704 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5747_6
timestamp 1731220412
transform 1 0 4480 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5746_6
timestamp 1731220412
transform 1 0 4928 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5745_6
timestamp 1731220412
transform 1 0 5064 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5744_6
timestamp 1731220412
transform 1 0 4760 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5743_6
timestamp 1731220412
transform 1 0 4840 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5742_6
timestamp 1731220412
transform 1 0 5120 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5741_6
timestamp 1731220412
transform 1 0 5176 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5740_6
timestamp 1731220412
transform 1 0 4912 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5739_6
timestamp 1731220412
transform 1 0 4848 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5738_6
timestamp 1731220412
transform 1 0 5048 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5737_6
timestamp 1731220412
transform 1 0 5256 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5736_6
timestamp 1731220412
transform 1 0 5232 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5735_6
timestamp 1731220412
transform 1 0 4968 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5734_6
timestamp 1731220412
transform 1 0 4712 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5733_6
timestamp 1731220412
transform 1 0 4472 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5732_6
timestamp 1731220412
transform 1 0 4248 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5731_6
timestamp 1731220412
transform 1 0 4328 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5730_6
timestamp 1731220412
transform 1 0 4488 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5729_6
timestamp 1731220412
transform 1 0 4656 0 -1 4424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5728_6
timestamp 1731220412
transform 1 0 4656 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5727_6
timestamp 1731220412
transform 1 0 4408 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5726_6
timestamp 1731220412
transform 1 0 4176 0 1 4432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5725_6
timestamp 1731220412
transform 1 0 4032 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5724_6
timestamp 1731220412
transform 1 0 4296 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5723_6
timestamp 1731220412
transform 1 0 4568 0 -1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5722_6
timestamp 1731220412
transform 1 0 4464 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5721_6
timestamp 1731220412
transform 1 0 4184 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5720_6
timestamp 1731220412
transform 1 0 3912 0 1 4656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5719_6
timestamp 1731220412
transform 1 0 3856 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5718_6
timestamp 1731220412
transform 1 0 4040 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5717_6
timestamp 1731220412
transform 1 0 4256 0 -1 4884
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5716_6
timestamp 1731220412
transform 1 0 4208 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5715_6
timestamp 1731220412
transform 1 0 4016 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5714_6
timestamp 1731220412
transform 1 0 3856 0 1 4904
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5713_6
timestamp 1731220412
transform 1 0 3856 0 -1 5140
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5712_6
timestamp 1731220412
transform 1 0 3648 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5711_6
timestamp 1731220412
transform 1 0 3648 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5710_6
timestamp 1731220412
transform 1 0 3464 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5709_6
timestamp 1731220412
transform 1 0 3256 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5708_6
timestamp 1731220412
transform 1 0 3376 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5707_6
timestamp 1731220412
transform 1 0 3576 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5706_6
timestamp 1731220412
transform 1 0 3576 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5705_6
timestamp 1731220412
transform 1 0 3392 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5704_6
timestamp 1731220412
transform 1 0 3216 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5703_6
timestamp 1731220412
transform 1 0 3288 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5702_6
timestamp 1731220412
transform 1 0 3464 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5701_6
timestamp 1731220412
transform 1 0 3640 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5700_6
timestamp 1731220412
transform 1 0 3648 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5699_6
timestamp 1731220412
transform 1 0 3512 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5698_6
timestamp 1731220412
transform 1 0 3352 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5697_6
timestamp 1731220412
transform 1 0 3192 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5696_6
timestamp 1731220412
transform 1 0 3032 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5695_6
timestamp 1731220412
transform 1 0 2864 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5694_6
timestamp 1731220412
transform 1 0 2696 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5693_6
timestamp 1731220412
transform 1 0 2752 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5692_6
timestamp 1731220412
transform 1 0 2936 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5691_6
timestamp 1731220412
transform 1 0 3112 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5690_6
timestamp 1731220412
transform 1 0 3040 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5689_6
timestamp 1731220412
transform 1 0 2856 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5688_6
timestamp 1731220412
transform 1 0 3000 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5687_6
timestamp 1731220412
transform 1 0 3184 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5686_6
timestamp 1731220412
transform 1 0 3056 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5685_6
timestamp 1731220412
transform 1 0 2856 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5684_6
timestamp 1731220412
transform 1 0 2528 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5683_6
timestamp 1731220412
transform 1 0 3096 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5682_6
timestamp 1731220412
transform 1 0 2840 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5681_6
timestamp 1731220412
transform 1 0 2976 0 -1 4944
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5680_6
timestamp 1731220412
transform 1 0 3128 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5679_6
timestamp 1731220412
transform 1 0 2928 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5678_6
timestamp 1731220412
transform 1 0 2728 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5677_6
timestamp 1731220412
transform 1 0 2664 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5676_6
timestamp 1731220412
transform 1 0 2888 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5675_6
timestamp 1731220412
transform 1 0 3336 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5674_6
timestamp 1731220412
transform 1 0 3112 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5673_6
timestamp 1731220412
transform 1 0 3000 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5672_6
timestamp 1731220412
transform 1 0 2792 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5671_6
timestamp 1731220412
transform 1 0 3200 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5670_6
timestamp 1731220412
transform 1 0 3400 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5669_6
timestamp 1731220412
transform 1 0 3608 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5668_6
timestamp 1731220412
transform 1 0 3648 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5667_6
timestamp 1731220412
transform 1 0 3464 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5666_6
timestamp 1731220412
transform 1 0 3256 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5665_6
timestamp 1731220412
transform 1 0 3048 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5664_6
timestamp 1731220412
transform 1 0 3448 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5663_6
timestamp 1731220412
transform 1 0 3648 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5662_6
timestamp 1731220412
transform 1 0 3856 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5661_6
timestamp 1731220412
transform 1 0 4040 0 1 4200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5660_6
timestamp 1731220412
transform 1 0 3856 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5659_6
timestamp 1731220412
transform 1 0 4944 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5658_6
timestamp 1731220412
transform 1 0 4384 0 -1 4164
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5657_6
timestamp 1731220412
transform 1 0 4168 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5656_6
timestamp 1731220412
transform 1 0 4000 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5655_6
timestamp 1731220412
transform 1 0 3856 0 1 3940
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5654_6
timestamp 1731220412
transform 1 0 3648 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5653_6
timestamp 1731220412
transform 1 0 3480 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5652_6
timestamp 1731220412
transform 1 0 3288 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5651_6
timestamp 1731220412
transform 1 0 3104 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5650_6
timestamp 1731220412
transform 1 0 2912 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5649_6
timestamp 1731220412
transform 1 0 3400 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5648_6
timestamp 1731220412
transform 1 0 3192 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5647_6
timestamp 1731220412
transform 1 0 2992 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5646_6
timestamp 1731220412
transform 1 0 2792 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5645_6
timestamp 1731220412
transform 1 0 2584 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5644_6
timestamp 1731220412
transform 1 0 2448 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5643_6
timestamp 1731220412
transform 1 0 2648 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5642_6
timestamp 1731220412
transform 1 0 2848 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5641_6
timestamp 1731220412
transform 1 0 3248 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5640_6
timestamp 1731220412
transform 1 0 3048 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5639_6
timestamp 1731220412
transform 1 0 2976 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5638_6
timestamp 1731220412
transform 1 0 2752 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5637_6
timestamp 1731220412
transform 1 0 3192 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5636_6
timestamp 1731220412
transform 1 0 3408 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5635_6
timestamp 1731220412
transform 1 0 3624 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5634_6
timestamp 1731220412
transform 1 0 3448 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5633_6
timestamp 1731220412
transform 1 0 3232 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5632_6
timestamp 1731220412
transform 1 0 3016 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5631_6
timestamp 1731220412
transform 1 0 3648 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5630_6
timestamp 1731220412
transform 1 0 3856 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5629_6
timestamp 1731220412
transform 1 0 4120 0 -1 3396
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5628_6
timestamp 1731220412
transform 1 0 3856 0 1 3172
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5627_6
timestamp 1731220412
transform 1 0 3872 0 -1 3156
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5626_6
timestamp 1731220412
transform 1 0 3904 0 1 2932
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5625_6
timestamp 1731220412
transform 1 0 3864 0 -1 2928
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5624_6
timestamp 1731220412
transform 1 0 3856 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5623_6
timestamp 1731220412
transform 1 0 3992 0 1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5622_6
timestamp 1731220412
transform 1 0 3928 0 -1 2696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5621_6
timestamp 1731220412
transform 1 0 3856 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5620_6
timestamp 1731220412
transform 1 0 4080 0 1 2472
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5619_6
timestamp 1731220412
transform 1 0 4056 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5618_6
timestamp 1731220412
transform 1 0 3856 0 -1 2468
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5617_6
timestamp 1731220412
transform 1 0 3648 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5616_6
timestamp 1731220412
transform 1 0 3648 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5615_6
timestamp 1731220412
transform 1 0 3480 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5614_6
timestamp 1731220412
transform 1 0 3408 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5613_6
timestamp 1731220412
transform 1 0 3152 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5612_6
timestamp 1731220412
transform 1 0 2896 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5611_6
timestamp 1731220412
transform 1 0 2824 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5610_6
timestamp 1731220412
transform 1 0 2960 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5609_6
timestamp 1731220412
transform 1 0 3096 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5608_6
timestamp 1731220412
transform 1 0 2984 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5607_6
timestamp 1731220412
transform 1 0 2728 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5606_6
timestamp 1731220412
transform 1 0 2472 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5605_6
timestamp 1731220412
transform 1 0 2752 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5604_6
timestamp 1731220412
transform 1 0 3000 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5603_6
timestamp 1731220412
transform 1 0 2904 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5602_6
timestamp 1731220412
transform 1 0 3104 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5601_6
timestamp 1731220412
transform 1 0 3304 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5600_6
timestamp 1731220412
transform 1 0 3232 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5599_6
timestamp 1731220412
transform 1 0 3464 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5598_6
timestamp 1731220412
transform 1 0 3400 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5597_6
timestamp 1731220412
transform 1 0 3208 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5596_6
timestamp 1731220412
transform 1 0 3592 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5595_6
timestamp 1731220412
transform 1 0 3552 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5594_6
timestamp 1731220412
transform 1 0 3368 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5593_6
timestamp 1731220412
transform 1 0 3184 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5592_6
timestamp 1731220412
transform 1 0 3000 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5591_6
timestamp 1731220412
transform 1 0 2808 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5590_6
timestamp 1731220412
transform 1 0 2832 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5589_6
timestamp 1731220412
transform 1 0 3024 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5588_6
timestamp 1731220412
transform 1 0 3000 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5587_6
timestamp 1731220412
transform 1 0 2776 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5586_6
timestamp 1731220412
transform 1 0 2712 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5585_6
timestamp 1731220412
transform 1 0 2504 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5584_6
timestamp 1731220412
transform 1 0 2216 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5583_6
timestamp 1731220412
transform 1 0 2552 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5582_6
timestamp 1731220412
transform 1 0 2688 0 1 2500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5581_6
timestamp 1731220412
transform 1 0 2648 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5580_6
timestamp 1731220412
transform 1 0 2416 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5579_6
timestamp 1731220412
transform 1 0 2192 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5578_6
timestamp 1731220412
transform 1 0 2536 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5577_6
timestamp 1731220412
transform 1 0 2728 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5576_6
timestamp 1731220412
transform 1 0 2680 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5575_6
timestamp 1731220412
transform 1 0 2504 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5574_6
timestamp 1731220412
transform 1 0 2328 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5573_6
timestamp 1731220412
transform 1 0 2160 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5572_6
timestamp 1731220412
transform 1 0 1992 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5571_6
timestamp 1731220412
transform 1 0 2344 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5570_6
timestamp 1731220412
transform 1 0 2152 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5569_6
timestamp 1731220412
transform 1 0 1992 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5568_6
timestamp 1731220412
transform 1 0 1992 0 -1 2476
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5567_6
timestamp 1731220412
transform 1 0 1784 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5566_6
timestamp 1731220412
transform 1 0 1784 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5565_6
timestamp 1731220412
transform 1 0 1600 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5564_6
timestamp 1731220412
transform 1 0 1400 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5563_6
timestamp 1731220412
transform 1 0 1512 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5562_6
timestamp 1731220412
transform 1 0 1672 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5561_6
timestamp 1731220412
transform 1 0 1768 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5560_6
timestamp 1731220412
transform 1 0 1992 0 -1 2736
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5559_6
timestamp 1731220412
transform 1 0 2008 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5558_6
timestamp 1731220412
transform 1 0 2256 0 1 2740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5557_6
timestamp 1731220412
transform 1 0 2112 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5556_6
timestamp 1731220412
transform 1 0 2312 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5555_6
timestamp 1731220412
transform 1 0 2512 0 -1 2972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5554_6
timestamp 1731220412
transform 1 0 2552 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5553_6
timestamp 1731220412
transform 1 0 2328 0 1 2984
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5552_6
timestamp 1731220412
transform 1 0 2432 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5551_6
timestamp 1731220412
transform 1 0 2632 0 -1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5550_6
timestamp 1731220412
transform 1 0 2616 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5549_6
timestamp 1731220412
transform 1 0 2408 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5548_6
timestamp 1731220412
transform 1 0 2800 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5547_6
timestamp 1731220412
transform 1 0 2584 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5546_6
timestamp 1731220412
transform 1 0 2512 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5545_6
timestamp 1731220412
transform 1 0 2248 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5544_6
timestamp 1731220412
transform 1 0 2248 0 -1 3728
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5543_6
timestamp 1731220412
transform 1 0 2368 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5542_6
timestamp 1731220412
transform 1 0 2136 0 1 3732
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5541_6
timestamp 1731220412
transform 1 0 2088 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5540_6
timestamp 1731220412
transform 1 0 2296 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5539_6
timestamp 1731220412
transform 1 0 2712 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5538_6
timestamp 1731220412
transform 1 0 2504 0 -1 3968
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5537_6
timestamp 1731220412
transform 1 0 2424 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5536_6
timestamp 1731220412
transform 1 0 2288 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5535_6
timestamp 1731220412
transform 1 0 2832 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5534_6
timestamp 1731220412
transform 1 0 2696 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5533_6
timestamp 1731220412
transform 1 0 2560 0 1 3972
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5532_6
timestamp 1731220412
transform 1 0 2536 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5531_6
timestamp 1731220412
transform 1 0 2672 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5530_6
timestamp 1731220412
transform 1 0 2808 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5529_6
timestamp 1731220412
transform 1 0 2944 0 -1 4216
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5528_6
timestamp 1731220412
transform 1 0 3224 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5527_6
timestamp 1731220412
transform 1 0 3008 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5526_6
timestamp 1731220412
transform 1 0 2808 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5525_6
timestamp 1731220412
transform 1 0 2624 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5524_6
timestamp 1731220412
transform 1 0 2456 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5523_6
timestamp 1731220412
transform 1 0 2304 0 1 4224
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5522_6
timestamp 1731220412
transform 1 0 2840 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5521_6
timestamp 1731220412
transform 1 0 2632 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5520_6
timestamp 1731220412
transform 1 0 2416 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5519_6
timestamp 1731220412
transform 1 0 2200 0 -1 4456
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5518_6
timestamp 1731220412
transform 1 0 2096 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5517_6
timestamp 1731220412
transform 1 0 2344 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5516_6
timestamp 1731220412
transform 1 0 2576 0 1 4464
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5515_6
timestamp 1731220412
transform 1 0 2440 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5514_6
timestamp 1731220412
transform 1 0 2208 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5513_6
timestamp 1731220412
transform 1 0 1992 0 -1 4692
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5512_6
timestamp 1731220412
transform 1 0 2536 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5511_6
timestamp 1731220412
transform 1 0 2344 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5510_6
timestamp 1731220412
transform 1 0 2152 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5509_6
timestamp 1731220412
transform 1 0 1992 0 1 4696
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5508_6
timestamp 1731220412
transform 1 0 1784 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5507_6
timestamp 1731220412
transform 1 0 1544 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5506_6
timestamp 1731220412
transform 1 0 1280 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5505_6
timestamp 1731220412
transform 1 0 1488 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5504_6
timestamp 1731220412
transform 1 0 1784 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5503_6
timestamp 1731220412
transform 1 0 1648 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5502_6
timestamp 1731220412
transform 1 0 1648 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5501_6
timestamp 1731220412
transform 1 0 1464 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5500_6
timestamp 1731220412
transform 1 0 1464 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5499_6
timestamp 1731220412
transform 1 0 1736 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5498_6
timestamp 1731220412
transform 1 0 1600 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5497_6
timestamp 1731220412
transform 1 0 1544 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5496_6
timestamp 1731220412
transform 1 0 1408 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5495_6
timestamp 1731220412
transform 1 0 1272 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5494_6
timestamp 1731220412
transform 1 0 1288 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5493_6
timestamp 1731220412
transform 1 0 1120 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5492_6
timestamp 1731220412
transform 1 0 1160 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5491_6
timestamp 1731220412
transform 1 0 936 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5490_6
timestamp 1731220412
transform 1 0 1024 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5489_6
timestamp 1731220412
transform 1 0 1040 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5488_6
timestamp 1731220412
transform 1 0 1080 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5487_6
timestamp 1731220412
transform 1 0 904 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5486_6
timestamp 1731220412
transform 1 0 464 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5485_6
timestamp 1731220412
transform 1 0 504 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5484_6
timestamp 1731220412
transform 1 0 424 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5483_6
timestamp 1731220412
transform 1 0 168 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5482_6
timestamp 1731220412
transform 1 0 480 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5481_6
timestamp 1731220412
transform 1 0 784 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5480_6
timestamp 1731220412
transform 1 0 1008 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5479_6
timestamp 1731220412
transform 1 0 760 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5478_6
timestamp 1731220412
transform 1 0 520 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5477_6
timestamp 1731220412
transform 1 0 304 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5476_6
timestamp 1731220412
transform 1 0 128 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5475_6
timestamp 1731220412
transform 1 0 248 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5474_6
timestamp 1731220412
transform 1 0 424 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5473_6
timestamp 1731220412
transform 1 0 616 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5472_6
timestamp 1731220412
transform 1 0 824 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5471_6
timestamp 1731220412
transform 1 0 1048 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5470_6
timestamp 1731220412
transform 1 0 888 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5469_6
timestamp 1731220412
transform 1 0 728 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5468_6
timestamp 1731220412
transform 1 0 568 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5467_6
timestamp 1731220412
transform 1 0 784 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5466_6
timestamp 1731220412
transform 1 0 568 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5465_6
timestamp 1731220412
transform 1 0 352 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5464_6
timestamp 1731220412
transform 1 0 224 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5463_6
timestamp 1731220412
transform 1 0 520 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5462_6
timestamp 1731220412
transform 1 0 568 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5461_6
timestamp 1731220412
transform 1 0 336 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5460_6
timestamp 1731220412
transform 1 0 128 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5459_6
timestamp 1731220412
transform 1 0 128 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5458_6
timestamp 1731220412
transform 1 0 344 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5457_6
timestamp 1731220412
transform 1 0 592 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5456_6
timestamp 1731220412
transform 1 0 512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5455_6
timestamp 1731220412
transform 1 0 376 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5454_6
timestamp 1731220412
transform 1 0 240 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5453_6
timestamp 1731220412
transform 1 0 184 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5452_6
timestamp 1731220412
transform 1 0 376 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5451_6
timestamp 1731220412
transform 1 0 344 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5450_6
timestamp 1731220412
transform 1 0 128 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5449_6
timestamp 1731220412
transform 1 0 128 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5448_6
timestamp 1731220412
transform 1 0 128 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5447_6
timestamp 1731220412
transform 1 0 344 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5446_6
timestamp 1731220412
transform 1 0 128 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5445_6
timestamp 1731220412
transform 1 0 128 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5444_6
timestamp 1731220412
transform 1 0 128 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5443_6
timestamp 1731220412
transform 1 0 144 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5442_6
timestamp 1731220412
transform 1 0 400 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5441_6
timestamp 1731220412
transform 1 0 232 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5440_6
timestamp 1731220412
transform 1 0 144 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5439_6
timestamp 1731220412
transform 1 0 128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5438_6
timestamp 1731220412
transform 1 0 312 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5437_6
timestamp 1731220412
transform 1 0 344 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5436_6
timestamp 1731220412
transform 1 0 128 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5435_6
timestamp 1731220412
transform 1 0 152 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5434_6
timestamp 1731220412
transform 1 0 480 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5433_6
timestamp 1731220412
transform 1 0 456 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5432_6
timestamp 1731220412
transform 1 0 248 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5431_6
timestamp 1731220412
transform 1 0 264 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5430_6
timestamp 1731220412
transform 1 0 128 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5429_6
timestamp 1731220412
transform 1 0 400 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5428_6
timestamp 1731220412
transform 1 0 536 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5427_6
timestamp 1731220412
transform 1 0 672 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5426_6
timestamp 1731220412
transform 1 0 1080 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5425_6
timestamp 1731220412
transform 1 0 944 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5424_6
timestamp 1731220412
transform 1 0 808 0 1 96
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5423_6
timestamp 1731220412
transform 1 0 672 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5422_6
timestamp 1731220412
transform 1 0 1104 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5421_6
timestamp 1731220412
transform 1 0 888 0 -1 360
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5420_6
timestamp 1731220412
transform 1 0 808 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5419_6
timestamp 1731220412
transform 1 0 1472 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5418_6
timestamp 1731220412
transform 1 0 1136 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5417_6
timestamp 1731220412
transform 1 0 968 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5416_6
timestamp 1731220412
transform 1 0 776 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5415_6
timestamp 1731220412
transform 1 0 568 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5414_6
timestamp 1731220412
transform 1 0 520 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5413_6
timestamp 1731220412
transform 1 0 904 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5412_6
timestamp 1731220412
transform 1 0 720 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5411_6
timestamp 1731220412
transform 1 0 640 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5410_6
timestamp 1731220412
transform 1 0 400 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5409_6
timestamp 1731220412
transform 1 0 456 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5408_6
timestamp 1731220412
transform 1 0 680 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5407_6
timestamp 1731220412
transform 1 0 656 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5406_6
timestamp 1731220412
transform 1 0 656 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5405_6
timestamp 1731220412
transform 1 0 472 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5404_6
timestamp 1731220412
transform 1 0 288 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5403_6
timestamp 1731220412
transform 1 0 328 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5402_6
timestamp 1731220412
transform 1 0 544 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5401_6
timestamp 1731220412
transform 1 0 408 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5400_6
timestamp 1731220412
transform 1 0 736 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5399_6
timestamp 1731220412
transform 1 0 576 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5398_6
timestamp 1731220412
transform 1 0 808 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5397_6
timestamp 1731220412
transform 1 0 976 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5396_6
timestamp 1731220412
transform 1 0 1272 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5395_6
timestamp 1731220412
transform 1 0 1160 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5394_6
timestamp 1731220412
transform 1 0 968 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5393_6
timestamp 1731220412
transform 1 0 1352 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5392_6
timestamp 1731220412
transform 1 0 1544 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5391_6
timestamp 1731220412
transform 1 0 1552 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5390_6
timestamp 1731220412
transform 1 0 1296 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5389_6
timestamp 1731220412
transform 1 0 1232 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5388_6
timestamp 1731220412
transform 1 0 1088 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5387_6
timestamp 1731220412
transform 1 0 1512 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5386_6
timestamp 1731220412
transform 1 0 1376 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5385_6
timestamp 1731220412
transform 1 0 1312 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5384_6
timestamp 1731220412
transform 1 0 1560 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5383_6
timestamp 1731220412
transform 1 0 1784 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5382_6
timestamp 1731220412
transform 1 0 1648 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5381_6
timestamp 1731220412
transform 1 0 1784 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5380_6
timestamp 1731220412
transform 1 0 1784 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5379_6
timestamp 1731220412
transform 1 0 1992 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5378_6
timestamp 1731220412
transform 1 0 2224 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5377_6
timestamp 1731220412
transform 1 0 2464 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5376_6
timestamp 1731220412
transform 1 0 2280 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5375_6
timestamp 1731220412
transform 1 0 2128 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5374_6
timestamp 1731220412
transform 1 0 1992 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5373_6
timestamp 1731220412
transform 1 0 2440 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5372_6
timestamp 1731220412
transform 1 0 2608 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5371_6
timestamp 1731220412
transform 1 0 2768 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5370_6
timestamp 1731220412
transform 1 0 2632 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5369_6
timestamp 1731220412
transform 1 0 2496 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5368_6
timestamp 1731220412
transform 1 0 2360 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5367_6
timestamp 1731220412
transform 1 0 2224 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5366_6
timestamp 1731220412
transform 1 0 2088 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5365_6
timestamp 1731220412
transform 1 0 2536 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5364_6
timestamp 1731220412
transform 1 0 2400 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5363_6
timestamp 1731220412
transform 1 0 2264 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5362_6
timestamp 1731220412
transform 1 0 2128 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5361_6
timestamp 1731220412
transform 1 0 1992 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5360_6
timestamp 1731220412
transform 1 0 2272 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5359_6
timestamp 1731220412
transform 1 0 1992 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5358_6
timestamp 1731220412
transform 1 0 1784 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5357_6
timestamp 1731220412
transform 1 0 1784 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5356_6
timestamp 1731220412
transform 1 0 1632 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5355_6
timestamp 1731220412
transform 1 0 1464 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5354_6
timestamp 1731220412
transform 1 0 1296 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5353_6
timestamp 1731220412
transform 1 0 1120 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5352_6
timestamp 1731220412
transform 1 0 1168 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5351_6
timestamp 1731220412
transform 1 0 1328 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5350_6
timestamp 1731220412
transform 1 0 1488 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5349_6
timestamp 1731220412
transform 1 0 1648 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5348_6
timestamp 1731220412
transform 1 0 1784 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5347_6
timestamp 1731220412
transform 1 0 1992 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5346_6
timestamp 1731220412
transform 1 0 1992 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5345_6
timestamp 1731220412
transform 1 0 2160 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5344_6
timestamp 1731220412
transform 1 0 2344 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5343_6
timestamp 1731220412
transform 1 0 2176 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5342_6
timestamp 1731220412
transform 1 0 1992 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5341_6
timestamp 1731220412
transform 1 0 2400 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5340_6
timestamp 1731220412
transform 1 0 2672 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5339_6
timestamp 1731220412
transform 1 0 3320 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5338_6
timestamp 1731220412
transform 1 0 2984 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5337_6
timestamp 1731220412
transform 1 0 2728 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5336_6
timestamp 1731220412
transform 1 0 2536 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5335_6
timestamp 1731220412
transform 1 0 2360 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5334_6
timestamp 1731220412
transform 1 0 2168 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5333_6
timestamp 1731220412
transform 1 0 2800 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5332_6
timestamp 1731220412
transform 1 0 2624 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5331_6
timestamp 1731220412
transform 1 0 2560 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5330_6
timestamp 1731220412
transform 1 0 2840 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5329_6
timestamp 1731220412
transform 1 0 2808 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5328_6
timestamp 1731220412
transform 1 0 2672 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5327_6
timestamp 1731220412
transform 1 0 2944 0 -1 1500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5326_6
timestamp 1731220412
transform 1 0 3176 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5325_6
timestamp 1731220412
transform 1 0 3040 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5324_6
timestamp 1731220412
transform 1 0 2904 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5323_6
timestamp 1731220412
transform 1 0 2776 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5322_6
timestamp 1731220412
transform 1 0 3120 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5321_6
timestamp 1731220412
transform 1 0 2944 0 -1 1752
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5320_6
timestamp 1731220412
transform 1 0 2904 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5319_6
timestamp 1731220412
transform 1 0 2688 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5318_6
timestamp 1731220412
transform 1 0 3104 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5317_6
timestamp 1731220412
transform 1 0 3096 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5316_6
timestamp 1731220412
transform 1 0 3232 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5315_6
timestamp 1731220412
transform 1 0 3368 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5314_6
timestamp 1731220412
transform 1 0 3376 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5313_6
timestamp 1731220412
transform 1 0 3240 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5312_6
timestamp 1731220412
transform 1 0 3104 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5311_6
timestamp 1731220412
transform 1 0 3016 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5310_6
timestamp 1731220412
transform 1 0 2848 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5309_6
timestamp 1731220412
transform 1 0 3176 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5308_6
timestamp 1731220412
transform 1 0 3112 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5307_6
timestamp 1731220412
transform 1 0 2920 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5306_6
timestamp 1731220412
transform 1 0 3296 0 1 2244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5305_6
timestamp 1731220412
transform 1 0 3336 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5304_6
timestamp 1731220412
transform 1 0 3504 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5303_6
timestamp 1731220412
transform 1 0 3648 0 -1 2236
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5302_6
timestamp 1731220412
transform 1 0 3648 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5301_6
timestamp 1731220412
transform 1 0 3512 0 1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5300_6
timestamp 1731220412
transform 1 0 3640 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5299_6
timestamp 1731220412
transform 1 0 3504 0 -1 1996
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5298_6
timestamp 1731220412
transform 1 0 3480 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5297_6
timestamp 1731220412
transform 1 0 3296 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5296_6
timestamp 1731220412
transform 1 0 3648 0 1 1760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5295_6
timestamp 1731220412
transform 1 0 3856 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5294_6
timestamp 1731220412
transform 1 0 4048 0 -1 1744
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5293_6
timestamp 1731220412
transform 1 0 4152 0 1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5292_6
timestamp 1731220412
transform 1 0 4128 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5291_6
timestamp 1731220412
transform 1 0 3992 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5290_6
timestamp 1731220412
transform 1 0 3856 0 -1 1520
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5289_6
timestamp 1731220412
transform 1 0 3856 0 1 1292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5288_6
timestamp 1731220412
transform 1 0 3648 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5287_6
timestamp 1731220412
transform 1 0 3392 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5286_6
timestamp 1731220412
transform 1 0 3120 0 1 1268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5285_6
timestamp 1731220412
transform 1 0 3512 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5284_6
timestamp 1731220412
transform 1 0 3328 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5283_6
timestamp 1731220412
transform 1 0 3152 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5282_6
timestamp 1731220412
transform 1 0 2976 0 -1 1244
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5281_6
timestamp 1731220412
transform 1 0 3216 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5280_6
timestamp 1731220412
transform 1 0 3056 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5279_6
timestamp 1731220412
transform 1 0 2888 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5278_6
timestamp 1731220412
transform 1 0 2720 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5277_6
timestamp 1731220412
transform 1 0 2544 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5276_6
timestamp 1731220412
transform 1 0 3384 0 1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5275_6
timestamp 1731220412
transform 1 0 3280 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5274_6
timestamp 1731220412
transform 1 0 3096 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5273_6
timestamp 1731220412
transform 1 0 2912 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5272_6
timestamp 1731220412
transform 1 0 3464 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5271_6
timestamp 1731220412
transform 1 0 3648 0 -1 1004
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5270_6
timestamp 1731220412
transform 1 0 3648 0 1 776
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5269_6
timestamp 1731220412
transform 1 0 3856 0 1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5268_6
timestamp 1731220412
transform 1 0 3856 0 -1 824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5267_6
timestamp 1731220412
transform 1 0 3856 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5266_6
timestamp 1731220412
transform 1 0 4400 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5265_6
timestamp 1731220412
transform 1 0 4264 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5264_6
timestamp 1731220412
transform 1 0 4128 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5263_6
timestamp 1731220412
transform 1 0 3992 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5262_6
timestamp 1731220412
transform 1 0 3856 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5261_6
timestamp 1731220412
transform 1 0 3648 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5260_6
timestamp 1731220412
transform 1 0 3512 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5259_6
timestamp 1731220412
transform 1 0 3376 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5258_6
timestamp 1731220412
transform 1 0 3240 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5257_6
timestamp 1731220412
transform 1 0 3104 0 -1 576
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5256_6
timestamp 1731220412
transform 1 0 3648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5255_6
timestamp 1731220412
transform 1 0 3464 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5254_6
timestamp 1731220412
transform 1 0 3264 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5253_6
timestamp 1731220412
transform 1 0 3064 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5252_6
timestamp 1731220412
transform 1 0 2856 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5251_6
timestamp 1731220412
transform 1 0 3624 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5250_6
timestamp 1731220412
transform 1 0 3488 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5249_6
timestamp 1731220412
transform 1 0 3352 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5248_6
timestamp 1731220412
transform 1 0 3216 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5247_6
timestamp 1731220412
transform 1 0 3080 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5246_6
timestamp 1731220412
transform 1 0 2944 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5245_6
timestamp 1731220412
transform 1 0 3624 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5244_6
timestamp 1731220412
transform 1 0 3488 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5243_6
timestamp 1731220412
transform 1 0 3352 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5242_6
timestamp 1731220412
transform 1 0 3216 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5241_6
timestamp 1731220412
transform 1 0 3080 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5240_6
timestamp 1731220412
transform 1 0 2944 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5239_6
timestamp 1731220412
transform 1 0 2808 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5238_6
timestamp 1731220412
transform 1 0 2672 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5237_6
timestamp 1731220412
transform 1 0 2536 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5236_6
timestamp 1731220412
transform 1 0 2400 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5235_6
timestamp 1731220412
transform 1 0 2264 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5234_6
timestamp 1731220412
transform 1 0 2128 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5233_6
timestamp 1731220412
transform 1 0 1992 0 1 76
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5232_6
timestamp 1731220412
transform 1 0 2808 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5231_6
timestamp 1731220412
transform 1 0 2672 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5230_6
timestamp 1731220412
transform 1 0 2536 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5229_6
timestamp 1731220412
transform 1 0 2400 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5228_6
timestamp 1731220412
transform 1 0 2264 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5227_6
timestamp 1731220412
transform 1 0 2128 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5226_6
timestamp 1731220412
transform 1 0 1992 0 -1 336
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5225_6
timestamp 1731220412
transform 1 0 2648 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5224_6
timestamp 1731220412
transform 1 0 2424 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5223_6
timestamp 1731220412
transform 1 0 2200 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5222_6
timestamp 1731220412
transform 1 0 1992 0 1 352
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5221_6
timestamp 1731220412
transform 1 0 1784 0 1 372
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5220_6
timestamp 1731220412
transform 1 0 1784 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5219_6
timestamp 1731220412
transform 1 0 1640 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5218_6
timestamp 1731220412
transform 1 0 1480 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5217_6
timestamp 1731220412
transform 1 0 1312 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5216_6
timestamp 1731220412
transform 1 0 1144 0 -1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5215_6
timestamp 1731220412
transform 1 0 1768 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5214_6
timestamp 1731220412
transform 1 0 1592 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5213_6
timestamp 1731220412
transform 1 0 1424 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5212_6
timestamp 1731220412
transform 1 0 1256 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5211_6
timestamp 1731220412
transform 1 0 1080 0 1 596
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5210_6
timestamp 1731220412
transform 1 0 872 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5209_6
timestamp 1731220412
transform 1 0 1096 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5208_6
timestamp 1731220412
transform 1 0 1320 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5207_6
timestamp 1731220412
transform 1 0 1544 0 -1 820
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5206_6
timestamp 1731220412
transform 1 0 1360 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5205_6
timestamp 1731220412
transform 1 0 1128 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5204_6
timestamp 1731220412
transform 1 0 904 0 1 836
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5203_6
timestamp 1731220412
transform 1 0 920 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5202_6
timestamp 1731220412
transform 1 0 1184 0 -1 1072
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5201_6
timestamp 1731220412
transform 1 0 1000 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5200_6
timestamp 1731220412
transform 1 0 832 0 1 1084
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5199_6
timestamp 1731220412
transform 1 0 744 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5198_6
timestamp 1731220412
transform 1 0 936 0 -1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5197_6
timestamp 1731220412
transform 1 0 1088 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5196_6
timestamp 1731220412
transform 1 0 1448 0 1 1320
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5195_6
timestamp 1731220412
transform 1 0 1272 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5194_6
timestamp 1731220412
transform 1 0 1040 0 -1 1556
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5193_6
timestamp 1731220412
transform 1 0 680 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5192_6
timestamp 1731220412
transform 1 0 392 0 1 1568
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5191_6
timestamp 1731220412
transform 1 0 560 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5190_6
timestamp 1731220412
transform 1 0 768 0 -1 1816
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5189_6
timestamp 1731220412
transform 1 0 1048 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5188_6
timestamp 1731220412
transform 1 0 808 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5187_6
timestamp 1731220412
transform 1 0 584 0 1 1824
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5186_6
timestamp 1731220412
transform 1 0 656 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5185_6
timestamp 1731220412
transform 1 0 800 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5184_6
timestamp 1731220412
transform 1 0 944 0 -1 2052
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5183_6
timestamp 1731220412
transform 1 0 832 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5182_6
timestamp 1731220412
transform 1 0 1072 0 1 2056
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5181_6
timestamp 1731220412
transform 1 0 1032 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5180_6
timestamp 1731220412
transform 1 0 800 0 -1 2292
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5179_6
timestamp 1731220412
transform 1 0 832 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5178_6
timestamp 1731220412
transform 1 0 1152 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5177_6
timestamp 1731220412
transform 1 0 1480 0 1 2308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5176_6
timestamp 1731220412
transform 1 0 1200 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5175_6
timestamp 1731220412
transform 1 0 992 0 -1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5174_6
timestamp 1731220412
transform 1 0 1040 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5173_6
timestamp 1731220412
transform 1 0 1192 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5172_6
timestamp 1731220412
transform 1 0 1352 0 1 2536
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5171_6
timestamp 1731220412
transform 1 0 1280 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5170_6
timestamp 1731220412
transform 1 0 1520 0 -1 2760
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5169_6
timestamp 1731220412
transform 1 0 1536 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5168_6
timestamp 1731220412
transform 1 0 1272 0 1 2764
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5167_6
timestamp 1731220412
transform 1 0 1080 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5166_6
timestamp 1731220412
transform 1 0 1384 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5165_6
timestamp 1731220412
transform 1 0 1688 0 -1 2988
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5164_6
timestamp 1731220412
transform 1 0 1784 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5163_6
timestamp 1731220412
transform 1 0 1648 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5162_6
timestamp 1731220412
transform 1 0 1512 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5161_6
timestamp 1731220412
transform 1 0 1440 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5160_6
timestamp 1731220412
transform 1 0 1624 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5159_6
timestamp 1731220412
transform 1 0 1784 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5158_6
timestamp 1731220412
transform 1 0 1992 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5157_6
timestamp 1731220412
transform 1 0 2192 0 1 3220
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5156_6
timestamp 1731220412
transform 1 0 2368 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5155_6
timestamp 1731220412
transform 1 0 2160 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5154_6
timestamp 1731220412
transform 1 0 1992 0 -1 3484
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5153_6
timestamp 1731220412
transform 1 0 1992 0 1 3492
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5152_6
timestamp 1731220412
transform 1 0 1784 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5151_6
timestamp 1731220412
transform 1 0 1784 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5150_6
timestamp 1731220412
transform 1 0 1648 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5149_6
timestamp 1731220412
transform 1 0 1488 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5148_6
timestamp 1731220412
transform 1 0 1336 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5147_6
timestamp 1731220412
transform 1 0 1184 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5146_6
timestamp 1731220412
transform 1 0 856 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5145_6
timestamp 1731220412
transform 1 0 680 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5144_6
timestamp 1731220412
transform 1 0 1288 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5143_6
timestamp 1731220412
transform 1 0 1544 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5142_6
timestamp 1731220412
transform 1 0 1456 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5141_6
timestamp 1731220412
transform 1 0 1264 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5140_6
timestamp 1731220412
transform 1 0 1312 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5139_6
timestamp 1731220412
transform 1 0 1264 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5138_6
timestamp 1731220412
transform 1 0 1080 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5137_6
timestamp 1731220412
transform 1 0 1376 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5136_6
timestamp 1731220412
transform 1 0 1240 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5135_6
timestamp 1731220412
transform 1 0 1104 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5134_6
timestamp 1731220412
transform 1 0 968 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5133_6
timestamp 1731220412
transform 1 0 832 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5132_6
timestamp 1731220412
transform 1 0 696 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5131_6
timestamp 1731220412
transform 1 0 560 0 1 3016
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5130_6
timestamp 1731220412
transform 1 0 696 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5129_6
timestamp 1731220412
transform 1 0 888 0 -1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5128_6
timestamp 1731220412
transform 1 0 1088 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5127_6
timestamp 1731220412
transform 1 0 872 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5126_6
timestamp 1731220412
transform 1 0 664 0 1 3248
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5125_6
timestamp 1731220412
transform 1 0 728 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5124_6
timestamp 1731220412
transform 1 0 568 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5123_6
timestamp 1731220412
transform 1 0 416 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5122_6
timestamp 1731220412
transform 1 0 272 0 -1 3488
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5121_6
timestamp 1731220412
transform 1 0 800 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5120_6
timestamp 1731220412
transform 1 0 568 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5119_6
timestamp 1731220412
transform 1 0 352 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5118_6
timestamp 1731220412
transform 1 0 144 0 1 3512
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5117_6
timestamp 1731220412
transform 1 0 128 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5116_6
timestamp 1731220412
transform 1 0 496 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5115_6
timestamp 1731220412
transform 1 0 304 0 -1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5114_6
timestamp 1731220412
transform 1 0 304 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5113_6
timestamp 1731220412
transform 1 0 128 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5112_6
timestamp 1731220412
transform 1 0 512 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5111_6
timestamp 1731220412
transform 1 0 720 0 1 3748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5110_6
timestamp 1731220412
transform 1 0 632 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5109_6
timestamp 1731220412
transform 1 0 480 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5108_6
timestamp 1731220412
transform 1 0 952 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5107_6
timestamp 1731220412
transform 1 0 792 0 -1 4000
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5106_6
timestamp 1731220412
transform 1 0 728 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5105_6
timestamp 1731220412
transform 1 0 864 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5104_6
timestamp 1731220412
transform 1 0 1000 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5103_6
timestamp 1731220412
transform 1 0 1136 0 1 4024
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5102_6
timestamp 1731220412
transform 1 0 1328 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5101_6
timestamp 1731220412
transform 1 0 1192 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_5100_6
timestamp 1731220412
transform 1 0 1056 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_599_6
timestamp 1731220412
transform 1 0 920 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_598_6
timestamp 1731220412
transform 1 0 784 0 -1 4252
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_597_6
timestamp 1731220412
transform 1 0 1288 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_596_6
timestamp 1731220412
transform 1 0 1120 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_595_6
timestamp 1731220412
transform 1 0 960 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_594_6
timestamp 1731220412
transform 1 0 808 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_593_6
timestamp 1731220412
transform 1 0 664 0 1 4268
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_592_6
timestamp 1731220412
transform 1 0 1376 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_591_6
timestamp 1731220412
transform 1 0 1112 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_590_6
timestamp 1731220412
transform 1 0 856 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_589_6
timestamp 1731220412
transform 1 0 624 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_588_6
timestamp 1731220412
transform 1 0 416 0 -1 4496
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_587_6
timestamp 1731220412
transform 1 0 1192 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_586_6
timestamp 1731220412
transform 1 0 904 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_585_6
timestamp 1731220412
transform 1 0 640 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_584_6
timestamp 1731220412
transform 1 0 392 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_583_6
timestamp 1731220412
transform 1 0 168 0 1 4500
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_582_6
timestamp 1731220412
transform 1 0 1024 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_581_6
timestamp 1731220412
transform 1 0 776 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_580_6
timestamp 1731220412
transform 1 0 536 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_579_6
timestamp 1731220412
transform 1 0 312 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_578_6
timestamp 1731220412
transform 1 0 128 0 -1 4740
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_577_6
timestamp 1731220412
transform 1 0 672 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_576_6
timestamp 1731220412
transform 1 0 536 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_575_6
timestamp 1731220412
transform 1 0 400 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_574_6
timestamp 1731220412
transform 1 0 264 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_573_6
timestamp 1731220412
transform 1 0 128 0 1 4748
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_572_6
timestamp 1731220412
transform 1 0 128 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_571_6
timestamp 1731220412
transform 1 0 312 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_570_6
timestamp 1731220412
transform 1 0 720 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_569_6
timestamp 1731220412
transform 1 0 520 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_568_6
timestamp 1731220412
transform 1 0 480 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_567_6
timestamp 1731220412
transform 1 0 344 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_566_6
timestamp 1731220412
transform 1 0 616 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_565_6
timestamp 1731220412
transform 1 0 752 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_564_6
timestamp 1731220412
transform 1 0 888 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_563_6
timestamp 1731220412
transform 1 0 1032 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_562_6
timestamp 1731220412
transform 1 0 1336 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_561_6
timestamp 1731220412
transform 1 0 1184 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_560_6
timestamp 1731220412
transform 1 0 1096 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_559_6
timestamp 1731220412
transform 1 0 912 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_558_6
timestamp 1731220412
transform 1 0 1280 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_557_6
timestamp 1731220412
transform 1 0 1456 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_556_6
timestamp 1731220412
transform 1 0 1632 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_555_6
timestamp 1731220412
transform 1 0 1784 0 -1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_554_6
timestamp 1731220412
transform 1 0 1648 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_553_6
timestamp 1731220412
transform 1 0 1488 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_552_6
timestamp 1731220412
transform 1 0 1784 0 1 4980
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_551_6
timestamp 1731220412
transform 1 0 1992 0 1 4976
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_550_6
timestamp 1731220412
transform 1 0 1992 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_549_6
timestamp 1731220412
transform 1 0 2128 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_548_6
timestamp 1731220412
transform 1 0 2664 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_547_6
timestamp 1731220412
transform 1 0 2480 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_546_6
timestamp 1731220412
transform 1 0 2296 0 -1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_545_6
timestamp 1731220412
transform 1 0 2192 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_544_6
timestamp 1731220412
transform 1 0 2336 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_543_6
timestamp 1731220412
transform 1 0 2488 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_542_6
timestamp 1731220412
transform 1 0 2648 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_541_6
timestamp 1731220412
transform 1 0 2816 0 1 5200
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_540_6
timestamp 1731220412
transform 1 0 2672 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_539_6
timestamp 1731220412
transform 1 0 2480 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_538_6
timestamp 1731220412
transform 1 0 2280 0 -1 5424
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_537_6
timestamp 1731220412
transform 1 0 2136 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_536_6
timestamp 1731220412
transform 1 0 2352 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_535_6
timestamp 1731220412
transform 1 0 2560 0 1 5432
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_534_6
timestamp 1731220412
transform 1 0 2520 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_533_6
timestamp 1731220412
transform 1 0 2336 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_532_6
timestamp 1731220412
transform 1 0 2152 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_531_6
timestamp 1731220412
transform 1 0 1992 0 -1 5656
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_530_6
timestamp 1731220412
transform 1 0 1784 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_529_6
timestamp 1731220412
transform 1 0 1512 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_528_6
timestamp 1731220412
transform 1 0 1736 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_527_6
timestamp 1731220412
transform 1 0 1480 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_526_6
timestamp 1731220412
transform 1 0 1232 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_525_6
timestamp 1731220412
transform 1 0 1256 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_524_6
timestamp 1731220412
transform 1 0 1488 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_523_6
timestamp 1731220412
transform 1 0 1512 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_522_6
timestamp 1731220412
transform 1 0 1376 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_521_6
timestamp 1731220412
transform 1 0 1240 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_520_6
timestamp 1731220412
transform 1 0 1104 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_519_6
timestamp 1731220412
transform 1 0 968 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_518_6
timestamp 1731220412
transform 1 0 832 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_517_6
timestamp 1731220412
transform 1 0 696 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_516_6
timestamp 1731220412
transform 1 0 560 0 -1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_515_6
timestamp 1731220412
transform 1 0 1032 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_514_6
timestamp 1731220412
transform 1 0 816 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_513_6
timestamp 1731220412
transform 1 0 608 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_512_6
timestamp 1731220412
transform 1 0 408 0 1 5308
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_511_6
timestamp 1731220412
transform 1 0 984 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_510_6
timestamp 1731220412
transform 1 0 736 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_59_6
timestamp 1731220412
transform 1 0 488 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_58_6
timestamp 1731220412
transform 1 0 248 0 -1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_57_6
timestamp 1731220412
transform 1 0 1224 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_56_6
timestamp 1731220412
transform 1 0 952 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_55_6
timestamp 1731220412
transform 1 0 696 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_54_6
timestamp 1731220412
transform 1 0 472 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_53_6
timestamp 1731220412
transform 1 0 272 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_52_6
timestamp 1731220412
transform 1 0 128 0 1 5532
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_51_6
timestamp 1731220412
transform 1 0 264 0 -1 5756
box 3 5 132 108
use _0_0std_0_0cells_0_0FAX1  tst_50_6
timestamp 1731220412
transform 1 0 128 0 -1 5756
box 3 5 132 108
<< end >>
